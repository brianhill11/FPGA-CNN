`ifndef RELU_BACKWARD_TEST_H
`define RELU_BACKWARD_TEST_H
reg [31:0] test_input [32];
reg [31:0] test_output [32];
initial begin
test_input[0:7] = '{32'h4263335c, 32'h40c5e004, 32'hc10ecd76, 32'hc234574d, 32'h429a1ec3, 32'hc29511fd, 32'hc230bfa6, 32'hc1e3c527};
test_output[0:7] = '{32'h4263335c, 32'h40c5e004, 32'h0, 32'h0, 32'h429a1ec3, 32'h0, 32'h0, 32'h0};
//############ DEBUG ############
test_input[0:7] = '{56.8001540825, 6.1835958546, -8.92516122294, -45.0852558653, 77.0600843176, -74.5351342745, -44.1871555525, -28.4712667127};
test_output[0:7] = '{56.8001540825, 6.1835958546, 0.0, 0.0, 77.0600843176, 0.0, 0.0, 0.0};
//############ END DEBUG ############
test_input[8:15] = '{32'hc280a753, 32'hc25c7b16, 32'h42520628, 32'h42038adc, 32'h4222b446, 32'h42c5de86, 32'hc1ed95fd, 32'h421b111c};
test_output[8:15] = '{32'h0, 32'h0, 32'h42520628, 32'h42038adc, 32'h4222b446, 32'h42c5de86, 32'h0, 32'h421b111c};
//############ DEBUG ############
test_input[8:15] = '{-64.3268041602, -55.1202022642, 52.5060120241, 32.8856055463, 40.6760468799, 98.9346179465, -29.6982371814, 38.7667074041};
test_output[8:15] = '{0.0, 0.0, 52.5060120241, 32.8856055463, 40.6760468799, 98.9346179465, 0.0, 38.7667074041};
//############ END DEBUG ############
test_input[16:23] = '{32'hc2b2b41b, 32'hc2471971, 32'hc26dd5e7, 32'h42915f19, 32'h4141a352, 32'hc2badca7, 32'h42296ee1, 32'h422b4b22};
test_output[16:23] = '{32'h0, 32'h0, 32'h0, 32'h42915f19, 32'h4141a352, 32'h0, 32'h42296ee1, 32'h422b4b22};
//############ DEBUG ############
test_input[16:23] = '{-89.351770573, -49.7748457119, -59.4588905815, 72.6857383973, 12.1023729536, -93.430964206, 42.3582786439, 42.8233715083};
test_output[16:23] = '{0.0, 0.0, 0.0, 72.6857383973, 12.1023729536, 0.0, 42.3582786439, 42.8233715083};
//############ END DEBUG ############
test_input[24:31] = '{32'hc2a45faf, 32'h4291e787, 32'h429fc169, 32'h419d2b60, 32'h429dd114, 32'h42167cb7, 32'h42b8dd37, 32'h42c1dc63};
test_output[24:31] = '{32'h0, 32'h4291e787, 32'h429fc169, 32'h419d2b60, 32'h429dd114, 32'h42167cb7, 32'h42b8dd37, 32'h42c1dc63};
//############ DEBUG ############
test_input[24:31] = '{-82.1868785675, 72.9522020312, 79.8777514968, 19.646179283, 78.9083533943, 37.6217937454, 92.432059414, 96.930441973};
test_output[24:31] = '{0.0, 72.9522020312, 79.8777514968, 19.646179283, 78.9083533943, 37.6217937454, 92.432059414, 96.930441973};
//############ END DEBUG ############
end
`endif
