`ifndef RELU_BACKWARD_TEST_H
`define RELU_BACKWARD_TEST_H
reg [31:0] test_input [32000];
reg [31:0] test_output [32000];
initial begin
test_input[0:7] = '{32'h427561dc, 32'hc2beb6d0, 32'hc287dcdf, 32'hc2a7a63c, 32'h424af192, 32'h41b32f48, 32'h41d3d4d4, 32'h4292ba86};
test_output[0:7] = '{32'h427561dc, 32'h0, 32'h0, 32'h0, 32'h424af192, 32'h41b32f48, 32'h41d3d4d4, 32'h4292ba86};
test_input[8:15] = '{32'hc29f92a9, 32'h429d2ca8, 32'hc1d3c6bf, 32'h42bae5ad, 32'h428eb550, 32'hc14f9bd5, 32'h40d26ae2, 32'hc1408e4b};
test_output[8:15] = '{32'h0, 32'h429d2ca8, 32'h0, 32'h42bae5ad, 32'h428eb550, 32'h0, 32'h40d26ae2, 32'h0};
test_input[16:23] = '{32'h428a839c, 32'hc1c8d9c6, 32'h42b5f433, 32'h4287843f, 32'hc2a7e465, 32'hc23c2ec5, 32'hc2170bb7, 32'h425629be};
test_output[16:23] = '{32'h428a839c, 32'h0, 32'h42b5f433, 32'h4287843f, 32'h0, 32'h0, 32'h0, 32'h425629be};
test_input[24:31] = '{32'h4228fb5e, 32'hc21b3dc5, 32'h429b56ae, 32'h42a9bee7, 32'h42b6d548, 32'hc201700c, 32'h42b904c2, 32'h4207cc04};
test_output[24:31] = '{32'h4228fb5e, 32'h0, 32'h429b56ae, 32'h42a9bee7, 32'h42b6d548, 32'h0, 32'h42b904c2, 32'h4207cc04};
test_input[32:39] = '{32'hc23259db, 32'h41874451, 32'h42ac92d3, 32'hc2ba27a7, 32'hc0e55510, 32'hc2331e37, 32'h4103d44c, 32'hc2862d59};
test_output[32:39] = '{32'h0, 32'h41874451, 32'h42ac92d3, 32'h0, 32'h0, 32'h0, 32'h4103d44c, 32'h0};
test_input[40:47] = '{32'h42a9a72f, 32'hc1fea3a4, 32'hc137b233, 32'h4193229a, 32'hc2b1cd45, 32'hc191cdba, 32'hc2c76be7, 32'h42628ebf};
test_output[40:47] = '{32'h42a9a72f, 32'h0, 32'h0, 32'h4193229a, 32'h0, 32'h0, 32'h0, 32'h42628ebf};
test_input[48:55] = '{32'h420b3f55, 32'hc1ce4744, 32'hc27c3fe2, 32'h4105338c, 32'h42a12d37, 32'hc2657d8f, 32'hc2884200, 32'h42aaefa2};
test_output[48:55] = '{32'h420b3f55, 32'h0, 32'h0, 32'h4105338c, 32'h42a12d37, 32'h0, 32'h0, 32'h42aaefa2};
test_input[56:63] = '{32'hc20f040b, 32'hc2c3e79d, 32'hc27b1cdb, 32'h4225a21a, 32'hc2823de6, 32'h40d94ea4, 32'hc24ff943, 32'h421b756e};
test_output[56:63] = '{32'h0, 32'h0, 32'h0, 32'h4225a21a, 32'h0, 32'h40d94ea4, 32'h0, 32'h421b756e};
test_input[64:71] = '{32'hc2a51869, 32'hc255629b, 32'hc1ae5b26, 32'h42aa86ca, 32'hc2190f15, 32'h3ec257aa, 32'hc2986d46, 32'h4209f35c};
test_output[64:71] = '{32'h0, 32'h0, 32'h0, 32'h42aa86ca, 32'h0, 32'h3ec257aa, 32'h0, 32'h4209f35c};
test_input[72:79] = '{32'hc2bdd3c4, 32'h429400de, 32'h42acd882, 32'h4271c0cd, 32'hc06850b3, 32'h426e9fd1, 32'hc195a16c, 32'h42a8be3f};
test_output[72:79] = '{32'h0, 32'h429400de, 32'h42acd882, 32'h4271c0cd, 32'h0, 32'h426e9fd1, 32'h0, 32'h42a8be3f};
test_input[80:87] = '{32'h4266ebb0, 32'h429106af, 32'h425e1b87, 32'h428cc31d, 32'h42b79d8e, 32'h4209a932, 32'h418ea19f, 32'h42bec318};
test_output[80:87] = '{32'h4266ebb0, 32'h429106af, 32'h425e1b87, 32'h428cc31d, 32'h42b79d8e, 32'h4209a932, 32'h418ea19f, 32'h42bec318};
test_input[88:95] = '{32'h400cad6f, 32'h42201c3e, 32'h424d460a, 32'hc2189d98, 32'hc1208dd0, 32'hc1cbf0f6, 32'hc21dc708, 32'h422627d6};
test_output[88:95] = '{32'h400cad6f, 32'h42201c3e, 32'h424d460a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422627d6};
test_input[96:103] = '{32'hc28fd09a, 32'h41ac1b1d, 32'h427ad952, 32'h42963792, 32'hc24d8da0, 32'h42a6bdf9, 32'hc24a41da, 32'h42808008};
test_output[96:103] = '{32'h0, 32'h41ac1b1d, 32'h427ad952, 32'h42963792, 32'h0, 32'h42a6bdf9, 32'h0, 32'h42808008};
test_input[104:111] = '{32'hc27eec79, 32'hc25062d9, 32'h41bc98cd, 32'hc26407d8, 32'h41ba6995, 32'hc275b48b, 32'hc2a73c73, 32'hc28db6c8};
test_output[104:111] = '{32'h0, 32'h0, 32'h41bc98cd, 32'h0, 32'h41ba6995, 32'h0, 32'h0, 32'h0};
test_input[112:119] = '{32'h42b84886, 32'h4282725a, 32'hc0d2a430, 32'h4240c0e1, 32'hc1da459f, 32'hc2ad7f3b, 32'h42850190, 32'h4289312f};
test_output[112:119] = '{32'h42b84886, 32'h4282725a, 32'h0, 32'h4240c0e1, 32'h0, 32'h0, 32'h42850190, 32'h4289312f};
test_input[120:127] = '{32'hc2aa1759, 32'h4228d7f4, 32'hc236e8bd, 32'h42b1a633, 32'h42272b9d, 32'hc102602f, 32'h419d20a8, 32'hc2a24d7d};
test_output[120:127] = '{32'h0, 32'h4228d7f4, 32'h0, 32'h42b1a633, 32'h42272b9d, 32'h0, 32'h419d20a8, 32'h0};
test_input[128:135] = '{32'hc237ec74, 32'h429a6d4d, 32'h4245077a, 32'hc2adf33e, 32'h412cf001, 32'h427b8861, 32'h429bdea2, 32'hc2839681};
test_output[128:135] = '{32'h0, 32'h429a6d4d, 32'h4245077a, 32'h0, 32'h412cf001, 32'h427b8861, 32'h429bdea2, 32'h0};
test_input[136:143] = '{32'hc24d0ded, 32'hc179cc88, 32'h429c12bc, 32'hc0e4d8fa, 32'h418544df, 32'hc1c482fc, 32'h428180f4, 32'hc1c8d003};
test_output[136:143] = '{32'h0, 32'h0, 32'h429c12bc, 32'h0, 32'h418544df, 32'h0, 32'h428180f4, 32'h0};
test_input[144:151] = '{32'h420309a1, 32'hc0cccaba, 32'h42915813, 32'h4270c8db, 32'h42a3897f, 32'h414157fc, 32'h422845ce, 32'h4210dd06};
test_output[144:151] = '{32'h420309a1, 32'h0, 32'h42915813, 32'h4270c8db, 32'h42a3897f, 32'h414157fc, 32'h422845ce, 32'h4210dd06};
test_input[152:159] = '{32'hc139d918, 32'hc212fff2, 32'h42bbd94b, 32'h41a3b7ab, 32'hc283b6d8, 32'hc2b772a9, 32'hc1b090e3, 32'hc2a3a96b};
test_output[152:159] = '{32'h0, 32'h0, 32'h42bbd94b, 32'h41a3b7ab, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[160:167] = '{32'hc2715519, 32'hc2637139, 32'h42416f41, 32'hc1d21a61, 32'hc0ecccbb, 32'h424980b8, 32'hc1c461e6, 32'hc23c3147};
test_output[160:167] = '{32'h0, 32'h0, 32'h42416f41, 32'h0, 32'h0, 32'h424980b8, 32'h0, 32'h0};
test_input[168:175] = '{32'hc18161db, 32'hc292003c, 32'h415c6fda, 32'h4211cc56, 32'hc29c606b, 32'hc1f52e51, 32'hc2179cf1, 32'h421cdf03};
test_output[168:175] = '{32'h0, 32'h0, 32'h415c6fda, 32'h4211cc56, 32'h0, 32'h0, 32'h0, 32'h421cdf03};
test_input[176:183] = '{32'h41af212f, 32'h421d6e26, 32'h42858815, 32'h4149d0ec, 32'hc0eb46ee, 32'h420fb8b4, 32'hc17b1bc9, 32'h4269323c};
test_output[176:183] = '{32'h41af212f, 32'h421d6e26, 32'h42858815, 32'h4149d0ec, 32'h0, 32'h420fb8b4, 32'h0, 32'h4269323c};
test_input[184:191] = '{32'h426d4346, 32'h42ab5f8b, 32'hc2ac4b95, 32'h4262c223, 32'h41599c5b, 32'hc0893267, 32'h4126cf8d, 32'hc237f687};
test_output[184:191] = '{32'h426d4346, 32'h42ab5f8b, 32'h0, 32'h4262c223, 32'h41599c5b, 32'h0, 32'h4126cf8d, 32'h0};
test_input[192:199] = '{32'h424ba453, 32'h41f7e7bf, 32'h42c4100d, 32'hc280a5bf, 32'h42384f49, 32'h418c6fbb, 32'hc28f41b2, 32'hc2b15a7c};
test_output[192:199] = '{32'h424ba453, 32'h41f7e7bf, 32'h42c4100d, 32'h0, 32'h42384f49, 32'h418c6fbb, 32'h0, 32'h0};
test_input[200:207] = '{32'hc190f114, 32'hc20bbe04, 32'hc2b65cd5, 32'h414bf233, 32'hc298a11f, 32'hc200a23a, 32'h42ad76ff, 32'hc216aa8e};
test_output[200:207] = '{32'h0, 32'h0, 32'h0, 32'h414bf233, 32'h0, 32'h0, 32'h42ad76ff, 32'h0};
test_input[208:215] = '{32'hc1f89ae6, 32'hc2a2b009, 32'hc2c7fd0a, 32'hc276b888, 32'hc2abbe3c, 32'hc285c192, 32'h429a94ec, 32'h421e6ec3};
test_output[208:215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429a94ec, 32'h421e6ec3};
test_input[216:223] = '{32'hc239b7d9, 32'h42a884cc, 32'hc2c73a33, 32'hc2024790, 32'hc222d8dd, 32'hc2af2171, 32'h428954cf, 32'hc0db5429};
test_output[216:223] = '{32'h0, 32'h42a884cc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428954cf, 32'h0};
test_input[224:231] = '{32'hc26810f6, 32'hc26d69e4, 32'hc27d931f, 32'hc2b73e10, 32'hc297793d, 32'h427b7d26, 32'hc2bec260, 32'hc2aea242};
test_output[224:231] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427b7d26, 32'h0, 32'h0};
test_input[232:239] = '{32'hc213a2dd, 32'h4234016d, 32'hc269c705, 32'h424ee065, 32'hc19efbd3, 32'h4205fa2b, 32'h4239e52c, 32'h42acefec};
test_output[232:239] = '{32'h0, 32'h4234016d, 32'h0, 32'h424ee065, 32'h0, 32'h4205fa2b, 32'h4239e52c, 32'h42acefec};
test_input[240:247] = '{32'hc2aa0587, 32'h429d7722, 32'hc2c1c06f, 32'hc221b422, 32'h42028b6b, 32'hc28e5841, 32'h4222f132, 32'h42b9569a};
test_output[240:247] = '{32'h0, 32'h429d7722, 32'h0, 32'h0, 32'h42028b6b, 32'h0, 32'h4222f132, 32'h42b9569a};
test_input[248:255] = '{32'h41983d36, 32'hc2140d16, 32'h428de0f3, 32'hc1f0176f, 32'hc2849e5e, 32'h4273e58f, 32'hc209ae22, 32'h41888298};
test_output[248:255] = '{32'h41983d36, 32'h0, 32'h428de0f3, 32'h0, 32'h0, 32'h4273e58f, 32'h0, 32'h41888298};
test_input[256:263] = '{32'h4227c4ba, 32'h42308c17, 32'hc2aed4e2, 32'hc2442825, 32'h4296e4e8, 32'hc152f915, 32'h4202bd4d, 32'h428329b8};
test_output[256:263] = '{32'h4227c4ba, 32'h42308c17, 32'h0, 32'h0, 32'h4296e4e8, 32'h0, 32'h4202bd4d, 32'h428329b8};
test_input[264:271] = '{32'h41879c27, 32'hc28625fc, 32'hc25ef2a5, 32'h422f92ab, 32'hc0cef961, 32'h4181508f, 32'h4251bb0a, 32'h4033ccab};
test_output[264:271] = '{32'h41879c27, 32'h0, 32'h0, 32'h422f92ab, 32'h0, 32'h4181508f, 32'h4251bb0a, 32'h4033ccab};
test_input[272:279] = '{32'hc20f2f73, 32'h42353627, 32'hc252b78b, 32'hc1155fd2, 32'h42b877c4, 32'h41a3d2e4, 32'h42927a7e, 32'hc27565e3};
test_output[272:279] = '{32'h0, 32'h42353627, 32'h0, 32'h0, 32'h42b877c4, 32'h41a3d2e4, 32'h42927a7e, 32'h0};
test_input[280:287] = '{32'h428aec4d, 32'hc2853710, 32'h420d0e86, 32'hc27d101f, 32'hc287b92e, 32'hc2b96625, 32'hc13df1f2, 32'hc1ab3fe1};
test_output[280:287] = '{32'h428aec4d, 32'h0, 32'h420d0e86, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[288:295] = '{32'h422180b2, 32'hc2911f7f, 32'hc26cd355, 32'h4250f5af, 32'h41250146, 32'h4283ba5e, 32'hc2b20ab4, 32'h42b20d38};
test_output[288:295] = '{32'h422180b2, 32'h0, 32'h0, 32'h4250f5af, 32'h41250146, 32'h4283ba5e, 32'h0, 32'h42b20d38};
test_input[296:303] = '{32'hc2bf9b7c, 32'hc242d326, 32'hc29f7e48, 32'h4293ceb0, 32'hc2b4d6f1, 32'hc25ab0ab, 32'h4228c8ec, 32'hc27229ad};
test_output[296:303] = '{32'h0, 32'h0, 32'h0, 32'h4293ceb0, 32'h0, 32'h0, 32'h4228c8ec, 32'h0};
test_input[304:311] = '{32'h4281a814, 32'hbf9e38b4, 32'hc22f9656, 32'h41cfe3eb, 32'hc294cce8, 32'hc1d28feb, 32'h42354b5f, 32'h419c52b0};
test_output[304:311] = '{32'h4281a814, 32'h0, 32'h0, 32'h41cfe3eb, 32'h0, 32'h0, 32'h42354b5f, 32'h419c52b0};
test_input[312:319] = '{32'hc236a354, 32'h42a4c206, 32'hc20be874, 32'hc23ad3e1, 32'h3f03fda9, 32'h42c7ec49, 32'h42930644, 32'h4234e7a4};
test_output[312:319] = '{32'h0, 32'h42a4c206, 32'h0, 32'h0, 32'h3f03fda9, 32'h42c7ec49, 32'h42930644, 32'h4234e7a4};
test_input[320:327] = '{32'hc24935d0, 32'hc2317635, 32'h41f4a8bd, 32'h4188c678, 32'hc290d724, 32'hc1adc328, 32'hc28fca62, 32'hc2179dca};
test_output[320:327] = '{32'h0, 32'h0, 32'h41f4a8bd, 32'h4188c678, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[328:335] = '{32'h42b6d6e7, 32'hc1349e23, 32'hc2468c3e, 32'hc2445d61, 32'hc2c241f1, 32'hc2bed042, 32'h42c09964, 32'h41b27370};
test_output[328:335] = '{32'h42b6d6e7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c09964, 32'h41b27370};
test_input[336:343] = '{32'hc0d42297, 32'hc27f212e, 32'hc240ef10, 32'h4291227c, 32'h42af81e9, 32'h401e6951, 32'hc1745144, 32'h42b2c8d7};
test_output[336:343] = '{32'h0, 32'h0, 32'h0, 32'h4291227c, 32'h42af81e9, 32'h401e6951, 32'h0, 32'h42b2c8d7};
test_input[344:351] = '{32'h428bb156, 32'h42bd4c97, 32'h4280a45e, 32'hc229bd31, 32'h4188a73a, 32'h42ab4af9, 32'hc22d1c9a, 32'h421e3c70};
test_output[344:351] = '{32'h428bb156, 32'h42bd4c97, 32'h4280a45e, 32'h0, 32'h4188a73a, 32'h42ab4af9, 32'h0, 32'h421e3c70};
test_input[352:359] = '{32'h422d30d6, 32'hc2007dd4, 32'h40d900b1, 32'h42ad54e4, 32'h411a6e8e, 32'hc2af68a2, 32'h423c2b7e, 32'hc121cd3e};
test_output[352:359] = '{32'h422d30d6, 32'h0, 32'h40d900b1, 32'h42ad54e4, 32'h411a6e8e, 32'h0, 32'h423c2b7e, 32'h0};
test_input[360:367] = '{32'h424b1687, 32'h41afde98, 32'h3fa41177, 32'h4299606d, 32'h41a023b9, 32'hc212faa1, 32'hc183ba0c, 32'hc20d4bbd};
test_output[360:367] = '{32'h424b1687, 32'h41afde98, 32'h3fa41177, 32'h4299606d, 32'h41a023b9, 32'h0, 32'h0, 32'h0};
test_input[368:375] = '{32'h42bc93d0, 32'hc29e3247, 32'h419f7d5f, 32'h428276d4, 32'hc2567eb3, 32'h41e9f5a6, 32'hc194aeb7, 32'hc2974a3f};
test_output[368:375] = '{32'h42bc93d0, 32'h0, 32'h419f7d5f, 32'h428276d4, 32'h0, 32'h41e9f5a6, 32'h0, 32'h0};
test_input[376:383] = '{32'h429dc92f, 32'hbfec48a5, 32'hc234613a, 32'hc193dd2a, 32'hc25e00b4, 32'h4218b0db, 32'h42883786, 32'h41f171e8};
test_output[376:383] = '{32'h429dc92f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4218b0db, 32'h42883786, 32'h41f171e8};
test_input[384:391] = '{32'h41d41957, 32'hc0acf7c2, 32'h42ae8289, 32'h4251a571, 32'hc2852027, 32'h42a1ab26, 32'hc2aff654, 32'h42799981};
test_output[384:391] = '{32'h41d41957, 32'h0, 32'h42ae8289, 32'h4251a571, 32'h0, 32'h42a1ab26, 32'h0, 32'h42799981};
test_input[392:399] = '{32'hc2616c87, 32'hc2bb3671, 32'hc20b4b22, 32'hc2952327, 32'hc121710c, 32'hc27e1305, 32'h41125555, 32'hc207a0fc};
test_output[392:399] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41125555, 32'h0};
test_input[400:407] = '{32'hc18ed6ff, 32'hc0272e69, 32'hc237b6bf, 32'h42a083b5, 32'h42c799f4, 32'h429aa13d, 32'hc2a67d03, 32'hc26af031};
test_output[400:407] = '{32'h0, 32'h0, 32'h0, 32'h42a083b5, 32'h42c799f4, 32'h429aa13d, 32'h0, 32'h0};
test_input[408:415] = '{32'hc2638be1, 32'h428555c1, 32'h4204e5e1, 32'hc2602bfb, 32'h428e08b0, 32'hc27b4bb3, 32'hc2b2abee, 32'h40a249de};
test_output[408:415] = '{32'h0, 32'h428555c1, 32'h4204e5e1, 32'h0, 32'h428e08b0, 32'h0, 32'h0, 32'h40a249de};
test_input[416:423] = '{32'h42bab132, 32'h428081c3, 32'h41e06eaf, 32'h427590de, 32'hc29ddee8, 32'h4220b3ff, 32'hc2949686, 32'hc1698ea9};
test_output[416:423] = '{32'h42bab132, 32'h428081c3, 32'h41e06eaf, 32'h427590de, 32'h0, 32'h4220b3ff, 32'h0, 32'h0};
test_input[424:431] = '{32'hc2c4441e, 32'h420e669f, 32'h42a87222, 32'hc155ab21, 32'hc2b18658, 32'hc11b9dd4, 32'h42519cc8, 32'h42bc5795};
test_output[424:431] = '{32'h0, 32'h420e669f, 32'h42a87222, 32'h0, 32'h0, 32'h0, 32'h42519cc8, 32'h42bc5795};
test_input[432:439] = '{32'h42c01e25, 32'hc2224730, 32'h40ea2371, 32'hc0617b71, 32'h428cb4b2, 32'hc2838b6e, 32'hc10dbef2, 32'hc29ddfe9};
test_output[432:439] = '{32'h42c01e25, 32'h0, 32'h40ea2371, 32'h0, 32'h428cb4b2, 32'h0, 32'h0, 32'h0};
test_input[440:447] = '{32'hc1951568, 32'h42bd780d, 32'hc22111fb, 32'h42a5b193, 32'h42979900, 32'hc1d719bb, 32'h428cfb92, 32'hc1b8032c};
test_output[440:447] = '{32'h0, 32'h42bd780d, 32'h0, 32'h42a5b193, 32'h42979900, 32'h0, 32'h428cfb92, 32'h0};
test_input[448:455] = '{32'hc26d8afc, 32'h4228006e, 32'hc1db3cce, 32'h42419ea0, 32'hc293e128, 32'hc2629dfd, 32'h42bc1af5, 32'h420d93c2};
test_output[448:455] = '{32'h0, 32'h4228006e, 32'h0, 32'h42419ea0, 32'h0, 32'h0, 32'h42bc1af5, 32'h420d93c2};
test_input[456:463] = '{32'h41d0f846, 32'h4299814a, 32'h42b0b77c, 32'hc22b1e6b, 32'h419465b3, 32'h422b7881, 32'h42a27ae1, 32'hc208ece2};
test_output[456:463] = '{32'h41d0f846, 32'h4299814a, 32'h42b0b77c, 32'h0, 32'h419465b3, 32'h422b7881, 32'h42a27ae1, 32'h0};
test_input[464:471] = '{32'hc2477e88, 32'hc117c69d, 32'hc1683d9b, 32'hc11d2c59, 32'hc2408597, 32'hc276b26e, 32'hc21bb742, 32'h42222375};
test_output[464:471] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42222375};
test_input[472:479] = '{32'hc2168068, 32'h4258cfba, 32'h41e3649e, 32'hc26f167f, 32'h420b42c5, 32'hc2c5467a, 32'hc2baa9da, 32'hc0cf3f40};
test_output[472:479] = '{32'h0, 32'h4258cfba, 32'h41e3649e, 32'h0, 32'h420b42c5, 32'h0, 32'h0, 32'h0};
test_input[480:487] = '{32'h42a38fd4, 32'hc2414fc5, 32'hc285c700, 32'h4288bb81, 32'hc2c2cda6, 32'h425b93a9, 32'hc2bc1b81, 32'hc24083e4};
test_output[480:487] = '{32'h42a38fd4, 32'h0, 32'h0, 32'h4288bb81, 32'h0, 32'h425b93a9, 32'h0, 32'h0};
test_input[488:495] = '{32'hc2312ed6, 32'hc2612531, 32'hc18b86dd, 32'h42c4e024, 32'h42a9ef48, 32'hc2a8ccde, 32'hc2347cf9, 32'hc244d203};
test_output[488:495] = '{32'h0, 32'h0, 32'h0, 32'h42c4e024, 32'h42a9ef48, 32'h0, 32'h0, 32'h0};
test_input[496:503] = '{32'h42927740, 32'h424f2a05, 32'h42b4f47a, 32'hc28a2dfd, 32'h4291fe8b, 32'hc2869d4a, 32'h426c29ab, 32'hc24e8e9c};
test_output[496:503] = '{32'h42927740, 32'h424f2a05, 32'h42b4f47a, 32'h0, 32'h4291fe8b, 32'h0, 32'h426c29ab, 32'h0};
test_input[504:511] = '{32'h42c45a11, 32'h41c2b6e9, 32'hc2725d77, 32'h429cf738, 32'hc2afdb66, 32'h41d5d21f, 32'h426d378c, 32'hc2c04779};
test_output[504:511] = '{32'h42c45a11, 32'h41c2b6e9, 32'h0, 32'h429cf738, 32'h0, 32'h41d5d21f, 32'h426d378c, 32'h0};
test_input[512:519] = '{32'hc279b192, 32'hc20d17b1, 32'h41a38dd5, 32'hc1d418eb, 32'hc2a32623, 32'hc18ce81f, 32'h42a3ca3b, 32'h42742e4a};
test_output[512:519] = '{32'h0, 32'h0, 32'h41a38dd5, 32'h0, 32'h0, 32'h0, 32'h42a3ca3b, 32'h42742e4a};
test_input[520:527] = '{32'hc28a6731, 32'hc2bd9f3f, 32'h429c3dca, 32'h411d2d2b, 32'h42b47d1d, 32'h41881f7f, 32'hc1f50787, 32'hc2bf8301};
test_output[520:527] = '{32'h0, 32'h0, 32'h429c3dca, 32'h411d2d2b, 32'h42b47d1d, 32'h41881f7f, 32'h0, 32'h0};
test_input[528:535] = '{32'hc28711c9, 32'h426ebfbc, 32'hc2808a98, 32'hc1d2b2a5, 32'hc241a813, 32'h422257f5, 32'hc27eca54, 32'hc27a219d};
test_output[528:535] = '{32'h0, 32'h426ebfbc, 32'h0, 32'h0, 32'h0, 32'h422257f5, 32'h0, 32'h0};
test_input[536:543] = '{32'h42937a5a, 32'hc1e612fc, 32'hc1692383, 32'hc2af1e9a, 32'h40c3e4ef, 32'hc28046ac, 32'h42b55b07, 32'hc01348f9};
test_output[536:543] = '{32'h42937a5a, 32'h0, 32'h0, 32'h0, 32'h40c3e4ef, 32'h0, 32'h42b55b07, 32'h0};
test_input[544:551] = '{32'hc2a29c7f, 32'hc1da39ac, 32'h4187ed50, 32'hc28d364d, 32'hc25f7ac3, 32'h41c423c9, 32'h42ba0d49, 32'h422b9c88};
test_output[544:551] = '{32'h0, 32'h0, 32'h4187ed50, 32'h0, 32'h0, 32'h41c423c9, 32'h42ba0d49, 32'h422b9c88};
test_input[552:559] = '{32'h42aed984, 32'hc1f88e4b, 32'h42308a23, 32'hc2728d6a, 32'h42687600, 32'hc2a798f4, 32'hbf9b978a, 32'h4265e3e2};
test_output[552:559] = '{32'h42aed984, 32'h0, 32'h42308a23, 32'h0, 32'h42687600, 32'h0, 32'h0, 32'h4265e3e2};
test_input[560:567] = '{32'h40f036e8, 32'h428778c1, 32'hc19bc87f, 32'h4202daf4, 32'h426a9f00, 32'h422d76a8, 32'h424df74d, 32'hc2865677};
test_output[560:567] = '{32'h40f036e8, 32'h428778c1, 32'h0, 32'h4202daf4, 32'h426a9f00, 32'h422d76a8, 32'h424df74d, 32'h0};
test_input[568:575] = '{32'h425e9472, 32'hc2945992, 32'hc2841d21, 32'h4242da0f, 32'h42281606, 32'h42b6f92c, 32'hc2740cd8, 32'hc2c3e041};
test_output[568:575] = '{32'h425e9472, 32'h0, 32'h0, 32'h4242da0f, 32'h42281606, 32'h42b6f92c, 32'h0, 32'h0};
test_input[576:583] = '{32'h4238aa4a, 32'hc2a13ba6, 32'hbfbce48d, 32'hc196f715, 32'h421bea2b, 32'hc28edb77, 32'h4241f3d2, 32'h42bef33d};
test_output[576:583] = '{32'h4238aa4a, 32'h0, 32'h0, 32'h0, 32'h421bea2b, 32'h0, 32'h4241f3d2, 32'h42bef33d};
test_input[584:591] = '{32'h42c1e162, 32'h3fd58644, 32'h421d0295, 32'h423847a2, 32'h414568ae, 32'h404f7b29, 32'hc297e439, 32'hc008c591};
test_output[584:591] = '{32'h42c1e162, 32'h3fd58644, 32'h421d0295, 32'h423847a2, 32'h414568ae, 32'h404f7b29, 32'h0, 32'h0};
test_input[592:599] = '{32'h4205d90d, 32'h42248087, 32'h42bd521d, 32'hc0e9aaf7, 32'h426556f4, 32'hc2ac640e, 32'h4241b29b, 32'h42172ac3};
test_output[592:599] = '{32'h4205d90d, 32'h42248087, 32'h42bd521d, 32'h0, 32'h426556f4, 32'h0, 32'h4241b29b, 32'h42172ac3};
test_input[600:607] = '{32'hc2beba02, 32'hc24fbe0b, 32'hc215f723, 32'hc29ee8e3, 32'hc285b045, 32'h419c46b3, 32'h421e3f9d, 32'h4269985c};
test_output[600:607] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h419c46b3, 32'h421e3f9d, 32'h4269985c};
test_input[608:615] = '{32'h4029a611, 32'h423924a7, 32'h41616057, 32'hc1f3cf0b, 32'h42b61e93, 32'h425f0063, 32'h4280a6c0, 32'h41882efc};
test_output[608:615] = '{32'h4029a611, 32'h423924a7, 32'h41616057, 32'h0, 32'h42b61e93, 32'h425f0063, 32'h4280a6c0, 32'h41882efc};
test_input[616:623] = '{32'hc1ad84b2, 32'hc22d7eaa, 32'h4259f0fd, 32'hc2910d1f, 32'h419f0bce, 32'h414cc172, 32'hc10bd2b9, 32'hc2034628};
test_output[616:623] = '{32'h0, 32'h0, 32'h4259f0fd, 32'h0, 32'h419f0bce, 32'h414cc172, 32'h0, 32'h0};
test_input[624:631] = '{32'h426ef4a9, 32'h425ea4cf, 32'hbf6e9c38, 32'h42c2f924, 32'hc1db6258, 32'h428836fa, 32'h428d6f43, 32'h41851d38};
test_output[624:631] = '{32'h426ef4a9, 32'h425ea4cf, 32'h0, 32'h42c2f924, 32'h0, 32'h428836fa, 32'h428d6f43, 32'h41851d38};
test_input[632:639] = '{32'hc2428514, 32'h40c8fd06, 32'hc2bfc170, 32'h41aa0eea, 32'h423853a7, 32'hc0411a9a, 32'hc1e6da65, 32'h42a0aa21};
test_output[632:639] = '{32'h0, 32'h40c8fd06, 32'h0, 32'h41aa0eea, 32'h423853a7, 32'h0, 32'h0, 32'h42a0aa21};
test_input[640:647] = '{32'hc25365e0, 32'h4221bd91, 32'h3dc35b0f, 32'hc291e8de, 32'hc1eac60d, 32'hc144add8, 32'h426395fb, 32'h42b2a1a2};
test_output[640:647] = '{32'h0, 32'h4221bd91, 32'h3dc35b0f, 32'h0, 32'h0, 32'h0, 32'h426395fb, 32'h42b2a1a2};
test_input[648:655] = '{32'hc2c41788, 32'h3f5d5571, 32'h42c4b13f, 32'h4239b8f6, 32'h42c7232f, 32'h424990c7, 32'h419d8f8b, 32'hc1a35c3d};
test_output[648:655] = '{32'h0, 32'h3f5d5571, 32'h42c4b13f, 32'h4239b8f6, 32'h42c7232f, 32'h424990c7, 32'h419d8f8b, 32'h0};
test_input[656:663] = '{32'hc1a8952a, 32'h4240ee57, 32'hc23bfb21, 32'hc2bea1ef, 32'hc20e240f, 32'h42b2b90a, 32'hc14902a9, 32'hc196af1f};
test_output[656:663] = '{32'h0, 32'h4240ee57, 32'h0, 32'h0, 32'h0, 32'h42b2b90a, 32'h0, 32'h0};
test_input[664:671] = '{32'h4254cc55, 32'hc1ea24ed, 32'hc2bc0d16, 32'h42b97c8e, 32'h40b0829b, 32'h420ee6c7, 32'hc263146a, 32'h3fb95fbb};
test_output[664:671] = '{32'h4254cc55, 32'h0, 32'h0, 32'h42b97c8e, 32'h40b0829b, 32'h420ee6c7, 32'h0, 32'h3fb95fbb};
test_input[672:679] = '{32'hc1daf4a6, 32'h4287a8b7, 32'hc2990217, 32'hc27d2ff0, 32'h40e4514a, 32'h42a5b9d5, 32'h41eae1d4, 32'hc2b1d89d};
test_output[672:679] = '{32'h0, 32'h4287a8b7, 32'h0, 32'h0, 32'h40e4514a, 32'h42a5b9d5, 32'h41eae1d4, 32'h0};
test_input[680:687] = '{32'h4052ce6f, 32'h4231f557, 32'hbf16f86a, 32'h42c77678, 32'h42b184ab, 32'hc26596c9, 32'h42a23b03, 32'h42c007fd};
test_output[680:687] = '{32'h4052ce6f, 32'h4231f557, 32'h0, 32'h42c77678, 32'h42b184ab, 32'h0, 32'h42a23b03, 32'h42c007fd};
test_input[688:695] = '{32'hc182a06b, 32'hc264c589, 32'hc172075d, 32'hc21dfee2, 32'h42868220, 32'h4279bf42, 32'h428a19a4, 32'h410e2cfa};
test_output[688:695] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42868220, 32'h4279bf42, 32'h428a19a4, 32'h410e2cfa};
test_input[696:703] = '{32'hc28e859f, 32'hc206a207, 32'h42622a6d, 32'hc1a5e766, 32'h427e56e6, 32'hc2323477, 32'hc2aef37c, 32'hc28313aa};
test_output[696:703] = '{32'h0, 32'h0, 32'h42622a6d, 32'h0, 32'h427e56e6, 32'h0, 32'h0, 32'h0};
test_input[704:711] = '{32'hc2382999, 32'hc1d6c316, 32'hc235c0e8, 32'h41b11d1c, 32'hc2b5597e, 32'h42b08e13, 32'h408ec426, 32'h41d823b1};
test_output[704:711] = '{32'h0, 32'h0, 32'h0, 32'h41b11d1c, 32'h0, 32'h42b08e13, 32'h408ec426, 32'h41d823b1};
test_input[712:719] = '{32'h422972b5, 32'h42135ae5, 32'h42740a9d, 32'hc203710f, 32'h42aced47, 32'h428ab0f1, 32'h428fb3f1, 32'h421f2d61};
test_output[712:719] = '{32'h422972b5, 32'h42135ae5, 32'h42740a9d, 32'h0, 32'h42aced47, 32'h428ab0f1, 32'h428fb3f1, 32'h421f2d61};
test_input[720:727] = '{32'hc28fcebe, 32'hc28b1058, 32'h4229c3c9, 32'hc2c5bc46, 32'h425a436c, 32'hc16b2a56, 32'h42a32e03, 32'hc20312bb};
test_output[720:727] = '{32'h0, 32'h0, 32'h4229c3c9, 32'h0, 32'h425a436c, 32'h0, 32'h42a32e03, 32'h0};
test_input[728:735] = '{32'h425215da, 32'hc2a26071, 32'h421883ec, 32'hc222db6d, 32'h4217387e, 32'hc10e6236, 32'h428de8bd, 32'hc04099df};
test_output[728:735] = '{32'h425215da, 32'h0, 32'h421883ec, 32'h0, 32'h4217387e, 32'h0, 32'h428de8bd, 32'h0};
test_input[736:743] = '{32'h40c37cbf, 32'hc234d440, 32'h4207caa6, 32'hc2894b09, 32'h42ab864d, 32'h41686f4f, 32'hc20c17d5, 32'hc2c1fb91};
test_output[736:743] = '{32'h40c37cbf, 32'h0, 32'h4207caa6, 32'h0, 32'h42ab864d, 32'h41686f4f, 32'h0, 32'h0};
test_input[744:751] = '{32'h42ba80e8, 32'h429430db, 32'hc244c74d, 32'hc21ca136, 32'h41390bf8, 32'h42bae464, 32'hc189c63b, 32'h429f01bd};
test_output[744:751] = '{32'h42ba80e8, 32'h429430db, 32'h0, 32'h0, 32'h41390bf8, 32'h42bae464, 32'h0, 32'h429f01bd};
test_input[752:759] = '{32'hc29911b8, 32'hc29bb685, 32'hbf9baa89, 32'hc0464a19, 32'hc28ddb1f, 32'h42c6a7a3, 32'hc0ac1a92, 32'h42276b39};
test_output[752:759] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c6a7a3, 32'h0, 32'h42276b39};
test_input[760:767] = '{32'hc28b0b23, 32'h424dacf2, 32'h42a1a7cf, 32'hc1be18fb, 32'h42474461, 32'hc28b3f4f, 32'hc2712d37, 32'hc2c65d72};
test_output[760:767] = '{32'h0, 32'h424dacf2, 32'h42a1a7cf, 32'h0, 32'h42474461, 32'h0, 32'h0, 32'h0};
test_input[768:775] = '{32'h4296453d, 32'h4299a875, 32'h42bb0e13, 32'hc232fafd, 32'h429526ae, 32'hc1a6dcfa, 32'h421b8f3c, 32'hc2c0a865};
test_output[768:775] = '{32'h4296453d, 32'h4299a875, 32'h42bb0e13, 32'h0, 32'h429526ae, 32'h0, 32'h421b8f3c, 32'h0};
test_input[776:783] = '{32'hc2acb373, 32'hc22a10b1, 32'h41635344, 32'h41a22fc0, 32'h421deb26, 32'hc2b9dc58, 32'h42930ab1, 32'h42989095};
test_output[776:783] = '{32'h0, 32'h0, 32'h41635344, 32'h41a22fc0, 32'h421deb26, 32'h0, 32'h42930ab1, 32'h42989095};
test_input[784:791] = '{32'h4219322e, 32'hc2a579e6, 32'hc20203db, 32'h41d22540, 32'h42029278, 32'h425321ce, 32'hc1ee7312, 32'hc2810886};
test_output[784:791] = '{32'h4219322e, 32'h0, 32'h0, 32'h41d22540, 32'h42029278, 32'h425321ce, 32'h0, 32'h0};
test_input[792:799] = '{32'h429ee607, 32'h3e549018, 32'hc1c7d7b0, 32'h42c45844, 32'hc0ddc50d, 32'hc2be31d4, 32'h416ba10b, 32'hc118d91b};
test_output[792:799] = '{32'h429ee607, 32'h3e549018, 32'h0, 32'h42c45844, 32'h0, 32'h0, 32'h416ba10b, 32'h0};
test_input[800:807] = '{32'h426139a7, 32'hc270101a, 32'h404fa37e, 32'h416b6f62, 32'hc2ba6543, 32'hc2081821, 32'h420b7e39, 32'h4261c55d};
test_output[800:807] = '{32'h426139a7, 32'h0, 32'h404fa37e, 32'h416b6f62, 32'h0, 32'h0, 32'h420b7e39, 32'h4261c55d};
test_input[808:815] = '{32'hc194d32a, 32'h42b89c2b, 32'h42b6e3f8, 32'hc219eb08, 32'hc0e43aae, 32'h425fd021, 32'h42a6ec79, 32'hc2363080};
test_output[808:815] = '{32'h0, 32'h42b89c2b, 32'h42b6e3f8, 32'h0, 32'h0, 32'h425fd021, 32'h42a6ec79, 32'h0};
test_input[816:823] = '{32'h42b2e5aa, 32'hc28cce31, 32'hc1c7d942, 32'h427b1cca, 32'h4276d319, 32'hc2b7989c, 32'h41806367, 32'h421b7916};
test_output[816:823] = '{32'h42b2e5aa, 32'h0, 32'h0, 32'h427b1cca, 32'h4276d319, 32'h0, 32'h41806367, 32'h421b7916};
test_input[824:831] = '{32'h421cc125, 32'hc294326d, 32'hc29c27a2, 32'h42acc455, 32'h42213a83, 32'hc1e7fcf0, 32'hc261e74e, 32'hc18e9185};
test_output[824:831] = '{32'h421cc125, 32'h0, 32'h0, 32'h42acc455, 32'h42213a83, 32'h0, 32'h0, 32'h0};
test_input[832:839] = '{32'h4290060b, 32'h413e2a9c, 32'hbffd7f17, 32'h42c2da02, 32'h429bcd0b, 32'h418ba1c0, 32'h41b09848, 32'h4281c02b};
test_output[832:839] = '{32'h4290060b, 32'h413e2a9c, 32'h0, 32'h42c2da02, 32'h429bcd0b, 32'h418ba1c0, 32'h41b09848, 32'h4281c02b};
test_input[840:847] = '{32'hc289012b, 32'hc2865dc8, 32'h429f05a1, 32'hc21c8ad7, 32'h42b3e400, 32'hc26e081f, 32'h420abab7, 32'h42a6da81};
test_output[840:847] = '{32'h0, 32'h0, 32'h429f05a1, 32'h0, 32'h42b3e400, 32'h0, 32'h420abab7, 32'h42a6da81};
test_input[848:855] = '{32'hc2c4899c, 32'hc2b3e336, 32'hc2441818, 32'h42a2aeb2, 32'h4217076f, 32'h426d9cb5, 32'h4014a398, 32'h418d4305};
test_output[848:855] = '{32'h0, 32'h0, 32'h0, 32'h42a2aeb2, 32'h4217076f, 32'h426d9cb5, 32'h4014a398, 32'h418d4305};
test_input[856:863] = '{32'h421aa289, 32'h4226cd96, 32'h4239d4de, 32'h42bbfb82, 32'hc27a6685, 32'hc2aa5390, 32'h42a1a2f6, 32'h428de796};
test_output[856:863] = '{32'h421aa289, 32'h4226cd96, 32'h4239d4de, 32'h42bbfb82, 32'h0, 32'h0, 32'h42a1a2f6, 32'h428de796};
test_input[864:871] = '{32'h428640a1, 32'h428608f7, 32'h41e6547c, 32'h423d27fa, 32'h42c5ecc0, 32'h410734ec, 32'h410c2bed, 32'h4183c769};
test_output[864:871] = '{32'h428640a1, 32'h428608f7, 32'h41e6547c, 32'h423d27fa, 32'h42c5ecc0, 32'h410734ec, 32'h410c2bed, 32'h4183c769};
test_input[872:879] = '{32'h420376ff, 32'h427d88d3, 32'h41e6501b, 32'h4227cfbd, 32'h41dcca4b, 32'h42a4886b, 32'h429fdf46, 32'h4292f6c4};
test_output[872:879] = '{32'h420376ff, 32'h427d88d3, 32'h41e6501b, 32'h4227cfbd, 32'h41dcca4b, 32'h42a4886b, 32'h429fdf46, 32'h4292f6c4};
test_input[880:887] = '{32'hc28883d7, 32'hc2c36a3d, 32'hc28f305e, 32'hc0793c20, 32'h429d6abe, 32'h42c24d9a, 32'h429a9d44, 32'hc234baa5};
test_output[880:887] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429d6abe, 32'h42c24d9a, 32'h429a9d44, 32'h0};
test_input[888:895] = '{32'h42c4bd0f, 32'h41ac8bbf, 32'hc2aaf7f5, 32'hbfbcadd8, 32'h41ea2c21, 32'h42bfea16, 32'hc2059bdf, 32'h41daee8b};
test_output[888:895] = '{32'h42c4bd0f, 32'h41ac8bbf, 32'h0, 32'h0, 32'h41ea2c21, 32'h42bfea16, 32'h0, 32'h41daee8b};
test_input[896:903] = '{32'hc2c3333e, 32'h42660621, 32'h42c43dd9, 32'h42c771bf, 32'h4272b6f4, 32'hc2be275b, 32'h4106b76f, 32'hc210f22c};
test_output[896:903] = '{32'h0, 32'h42660621, 32'h42c43dd9, 32'h42c771bf, 32'h4272b6f4, 32'h0, 32'h4106b76f, 32'h0};
test_input[904:911] = '{32'h4297e16d, 32'hc2bfeba7, 32'h4215dea7, 32'h42a5966e, 32'hc2af9931, 32'h3fdce752, 32'hc2339379, 32'h421134ee};
test_output[904:911] = '{32'h4297e16d, 32'h0, 32'h4215dea7, 32'h42a5966e, 32'h0, 32'h3fdce752, 32'h0, 32'h421134ee};
test_input[912:919] = '{32'h40ad8079, 32'hc142ca12, 32'h405f7e61, 32'h4157a4cb, 32'h42628f1b, 32'hc2bb057e, 32'h42aa01bb, 32'hc2597cf0};
test_output[912:919] = '{32'h40ad8079, 32'h0, 32'h405f7e61, 32'h4157a4cb, 32'h42628f1b, 32'h0, 32'h42aa01bb, 32'h0};
test_input[920:927] = '{32'hc2600f0f, 32'hc28cb12b, 32'hc2088be3, 32'h4189a2dc, 32'hc1d51fb5, 32'h429482d2, 32'h41049ab3, 32'hc09f86ab};
test_output[920:927] = '{32'h0, 32'h0, 32'h0, 32'h4189a2dc, 32'h0, 32'h429482d2, 32'h41049ab3, 32'h0};
test_input[928:935] = '{32'hc29490b4, 32'hc15858d8, 32'h42b6fd2e, 32'h3f0755b0, 32'hc27cf659, 32'hc27a0a88, 32'hc2c6f2b8, 32'hc2231e11};
test_output[928:935] = '{32'h0, 32'h0, 32'h42b6fd2e, 32'h3f0755b0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[936:943] = '{32'h3f17b8a1, 32'h413f0ec3, 32'hc295cf44, 32'hc259d361, 32'h4218d162, 32'h42bef436, 32'hc185a399, 32'h41ce6ecd};
test_output[936:943] = '{32'h3f17b8a1, 32'h413f0ec3, 32'h0, 32'h0, 32'h4218d162, 32'h42bef436, 32'h0, 32'h41ce6ecd};
test_input[944:951] = '{32'h41ddc0be, 32'hc29fb08c, 32'h4286a59a, 32'hc2ba88bc, 32'h41c9c0fd, 32'hc2c6d11e, 32'h4285247b, 32'hc29de6eb};
test_output[944:951] = '{32'h41ddc0be, 32'h0, 32'h4286a59a, 32'h0, 32'h41c9c0fd, 32'h0, 32'h4285247b, 32'h0};
test_input[952:959] = '{32'h4292a252, 32'h429a13bd, 32'h3fbca35c, 32'hc1354dd5, 32'h3f354792, 32'hc2a07d33, 32'hc284c06d, 32'h42c29a65};
test_output[952:959] = '{32'h4292a252, 32'h429a13bd, 32'h3fbca35c, 32'h0, 32'h3f354792, 32'h0, 32'h0, 32'h42c29a65};
test_input[960:967] = '{32'h422f43e7, 32'hc2c591cb, 32'hc0cee020, 32'hc2ae9638, 32'h40c25cc9, 32'h42bbf485, 32'hc2a0be00, 32'h42c097a8};
test_output[960:967] = '{32'h422f43e7, 32'h0, 32'h0, 32'h0, 32'h40c25cc9, 32'h42bbf485, 32'h0, 32'h42c097a8};
test_input[968:975] = '{32'h420778ea, 32'hc2c11b2c, 32'h42404284, 32'h4203705f, 32'hc1bdd958, 32'h42b06ab3, 32'h424f7609, 32'hc2479885};
test_output[968:975] = '{32'h420778ea, 32'h0, 32'h42404284, 32'h4203705f, 32'h0, 32'h42b06ab3, 32'h424f7609, 32'h0};
test_input[976:983] = '{32'h41f35fe4, 32'h41edd222, 32'h41373791, 32'h427b0b2b, 32'hc23e7304, 32'h42b2dd64, 32'hc1a57ebd, 32'hc2a07a38};
test_output[976:983] = '{32'h41f35fe4, 32'h41edd222, 32'h41373791, 32'h427b0b2b, 32'h0, 32'h42b2dd64, 32'h0, 32'h0};
test_input[984:991] = '{32'hc203015b, 32'h4211b33f, 32'h4277e98c, 32'h4254a09d, 32'hc01359b7, 32'h42376e3c, 32'hc2062b8b, 32'hc12a37b7};
test_output[984:991] = '{32'h0, 32'h4211b33f, 32'h4277e98c, 32'h4254a09d, 32'h0, 32'h42376e3c, 32'h0, 32'h0};
test_input[992:999] = '{32'hc2779ca4, 32'h41dcb723, 32'h40ffac97, 32'hc0d8d5eb, 32'hc1a30f70, 32'hc105e2e8, 32'hc2668e5d, 32'hc2a4b746};
test_output[992:999] = '{32'h0, 32'h41dcb723, 32'h40ffac97, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1000:1007] = '{32'hc2800ea6, 32'hc26f561f, 32'hc2107de2, 32'h4256746b, 32'hc209e565, 32'h42b5d83a, 32'hc13d97ad, 32'h42c0d81b};
test_output[1000:1007] = '{32'h0, 32'h0, 32'h0, 32'h4256746b, 32'h0, 32'h42b5d83a, 32'h0, 32'h42c0d81b};
test_input[1008:1015] = '{32'h42ae524d, 32'hc2356230, 32'h4282ddc2, 32'h42c304f7, 32'h41175da7, 32'hc2a16679, 32'h42c6558f, 32'hc1be49af};
test_output[1008:1015] = '{32'h42ae524d, 32'h0, 32'h4282ddc2, 32'h42c304f7, 32'h41175da7, 32'h0, 32'h42c6558f, 32'h0};
test_input[1016:1023] = '{32'hc2919ceb, 32'h42267740, 32'hc2b9d3f6, 32'h427358f0, 32'h419f71bd, 32'hc26455e7, 32'hc28ff452, 32'h42147d42};
test_output[1016:1023] = '{32'h0, 32'h42267740, 32'h0, 32'h427358f0, 32'h419f71bd, 32'h0, 32'h0, 32'h42147d42};
test_input[1024:1031] = '{32'h42902bbc, 32'hc2bfddc9, 32'hc2c04623, 32'hc20f5df1, 32'hc1b41018, 32'h421d8ca3, 32'hc29abc8c, 32'hc297789c};
test_output[1024:1031] = '{32'h42902bbc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h421d8ca3, 32'h0, 32'h0};
test_input[1032:1039] = '{32'hc2783c2f, 32'h4298d260, 32'hc20e5c1b, 32'hc278c02a, 32'h42220eb4, 32'hc2a68ebd, 32'h42785109, 32'hc23c92cb};
test_output[1032:1039] = '{32'h0, 32'h4298d260, 32'h0, 32'h0, 32'h42220eb4, 32'h0, 32'h42785109, 32'h0};
test_input[1040:1047] = '{32'h42165747, 32'h42bf7a38, 32'h427ee61c, 32'h4232b156, 32'h4268ebc4, 32'hc21ae3f2, 32'h427cca48, 32'hc2917179};
test_output[1040:1047] = '{32'h42165747, 32'h42bf7a38, 32'h427ee61c, 32'h4232b156, 32'h4268ebc4, 32'h0, 32'h427cca48, 32'h0};
test_input[1048:1055] = '{32'h42af831a, 32'h420a5e10, 32'h422db652, 32'hc166051a, 32'h42c54d3b, 32'h4281998e, 32'hc294b39d, 32'hc1581333};
test_output[1048:1055] = '{32'h42af831a, 32'h420a5e10, 32'h422db652, 32'h0, 32'h42c54d3b, 32'h4281998e, 32'h0, 32'h0};
test_input[1056:1063] = '{32'hc2c19817, 32'h418d4365, 32'hc0bb0cba, 32'h413d726d, 32'h4205b49d, 32'hc27dc0b9, 32'h41c64348, 32'hc1d7ffe6};
test_output[1056:1063] = '{32'h0, 32'h418d4365, 32'h0, 32'h413d726d, 32'h4205b49d, 32'h0, 32'h41c64348, 32'h0};
test_input[1064:1071] = '{32'hc1ec421b, 32'hc2839e4a, 32'hc284382d, 32'hbd959aee, 32'h428b2476, 32'hc28e1a99, 32'hc2a067cf, 32'hc11cef6b};
test_output[1064:1071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h428b2476, 32'h0, 32'h0, 32'h0};
test_input[1072:1079] = '{32'hc0b9c8ca, 32'hc13425cb, 32'h4261c450, 32'hc222a2e9, 32'h41b7b23c, 32'h42ae5b3e, 32'hc2668105, 32'h42c5d9c4};
test_output[1072:1079] = '{32'h0, 32'h0, 32'h4261c450, 32'h0, 32'h41b7b23c, 32'h42ae5b3e, 32'h0, 32'h42c5d9c4};
test_input[1080:1087] = '{32'hc0c599db, 32'hc101ada8, 32'h420b19f1, 32'h4094ccbb, 32'h41a428cf, 32'h3e3f1b62, 32'hc1cb8c07, 32'hc1aa3f1e};
test_output[1080:1087] = '{32'h0, 32'h0, 32'h420b19f1, 32'h4094ccbb, 32'h41a428cf, 32'h3e3f1b62, 32'h0, 32'h0};
test_input[1088:1095] = '{32'hc2351333, 32'h428475b7, 32'h429c8ccd, 32'h42b83896, 32'h40a57f4f, 32'hc237b0cc, 32'hc21f7a87, 32'hc2704070};
test_output[1088:1095] = '{32'h0, 32'h428475b7, 32'h429c8ccd, 32'h42b83896, 32'h40a57f4f, 32'h0, 32'h0, 32'h0};
test_input[1096:1103] = '{32'h422e4416, 32'hc18e986e, 32'hc2891c15, 32'hc28403b9, 32'hc19cb75f, 32'h420f6983, 32'hc1206ca6, 32'h41af7325};
test_output[1096:1103] = '{32'h422e4416, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420f6983, 32'h0, 32'h41af7325};
test_input[1104:1111] = '{32'hc23cddc8, 32'hc28dc23c, 32'h41f6a6bd, 32'h42925e5f, 32'h42bd29c3, 32'hc21db2a3, 32'h4229e929, 32'hc1aa9725};
test_output[1104:1111] = '{32'h0, 32'h0, 32'h41f6a6bd, 32'h42925e5f, 32'h42bd29c3, 32'h0, 32'h4229e929, 32'h0};
test_input[1112:1119] = '{32'hc2bc1981, 32'hc2616091, 32'h42874634, 32'h42a33896, 32'hc292aa9d, 32'hc213c7e2, 32'hc1773830, 32'hc00f39fd};
test_output[1112:1119] = '{32'h0, 32'h0, 32'h42874634, 32'h42a33896, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1120:1127] = '{32'hc2230976, 32'h4263a8cf, 32'hc2805143, 32'h42b7f6ba, 32'hc19432b8, 32'hc2b64591, 32'hc2a433a7, 32'h41ae34cc};
test_output[1120:1127] = '{32'h0, 32'h4263a8cf, 32'h0, 32'h42b7f6ba, 32'h0, 32'h0, 32'h0, 32'h41ae34cc};
test_input[1128:1135] = '{32'h423db3e8, 32'h42c3068d, 32'h4259af2e, 32'h429c2ba3, 32'h417669ef, 32'h42253e28, 32'h42b990af, 32'h42b46951};
test_output[1128:1135] = '{32'h423db3e8, 32'h42c3068d, 32'h4259af2e, 32'h429c2ba3, 32'h417669ef, 32'h42253e28, 32'h42b990af, 32'h42b46951};
test_input[1136:1143] = '{32'h423ccc7a, 32'h41ff1ef6, 32'h41b52c13, 32'h42905fdd, 32'h429c2963, 32'h418ff434, 32'hc1729c3b, 32'h406cd8c4};
test_output[1136:1143] = '{32'h423ccc7a, 32'h41ff1ef6, 32'h41b52c13, 32'h42905fdd, 32'h429c2963, 32'h418ff434, 32'h0, 32'h406cd8c4};
test_input[1144:1151] = '{32'hc2a8c9d0, 32'hc285da7d, 32'h41eba03d, 32'h428f78d4, 32'hc16891a5, 32'hc2a5f65e, 32'hc2b63c31, 32'hc28d315e};
test_output[1144:1151] = '{32'h0, 32'h0, 32'h41eba03d, 32'h428f78d4, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1152:1159] = '{32'h42303e19, 32'hc275c232, 32'hc2bef8f1, 32'hc0f68b3b, 32'hc2ba74dd, 32'hc171118e, 32'h42a3c0fc, 32'h42b02650};
test_output[1152:1159] = '{32'h42303e19, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a3c0fc, 32'h42b02650};
test_input[1160:1167] = '{32'hc156d4fe, 32'h41f21e1f, 32'h42b6eafd, 32'hc1b5e972, 32'h40d3bfc0, 32'hc2ad319d, 32'hc20bc5ee, 32'h4207e99c};
test_output[1160:1167] = '{32'h0, 32'h41f21e1f, 32'h42b6eafd, 32'h0, 32'h40d3bfc0, 32'h0, 32'h0, 32'h4207e99c};
test_input[1168:1175] = '{32'hc25892d2, 32'h42c52ebc, 32'h42a95d7c, 32'h4294bc91, 32'h4200e8b0, 32'h424ca9a2, 32'hc0e43678, 32'h42aaebec};
test_output[1168:1175] = '{32'h0, 32'h42c52ebc, 32'h42a95d7c, 32'h4294bc91, 32'h4200e8b0, 32'h424ca9a2, 32'h0, 32'h42aaebec};
test_input[1176:1183] = '{32'hc093f635, 32'h412872cc, 32'h4232a70a, 32'hc256846a, 32'h42ae4aee, 32'h4209f0c9, 32'h3fa9ca91, 32'hc23157bd};
test_output[1176:1183] = '{32'h0, 32'h412872cc, 32'h4232a70a, 32'h0, 32'h42ae4aee, 32'h4209f0c9, 32'h3fa9ca91, 32'h0};
test_input[1184:1191] = '{32'h42c6a4f5, 32'hc247e5aa, 32'hc1f03bac, 32'hc20af155, 32'h4273c344, 32'h42b853a3, 32'hc20c0559, 32'hc28b0a61};
test_output[1184:1191] = '{32'h42c6a4f5, 32'h0, 32'h0, 32'h0, 32'h4273c344, 32'h42b853a3, 32'h0, 32'h0};
test_input[1192:1199] = '{32'h42439b56, 32'hc2b60558, 32'hc2517f85, 32'h4196e904, 32'hc11b413e, 32'hc1bfff78, 32'h41cdf6bc, 32'hc265eade};
test_output[1192:1199] = '{32'h42439b56, 32'h0, 32'h0, 32'h4196e904, 32'h0, 32'h0, 32'h41cdf6bc, 32'h0};
test_input[1200:1207] = '{32'h425dab13, 32'h416e8ea3, 32'hc1b3bd82, 32'hc1820e89, 32'h42a16da8, 32'hc28f84d9, 32'hc29085fc, 32'h418acd07};
test_output[1200:1207] = '{32'h425dab13, 32'h416e8ea3, 32'h0, 32'h0, 32'h42a16da8, 32'h0, 32'h0, 32'h418acd07};
test_input[1208:1215] = '{32'h41e4c32c, 32'hc1a100b6, 32'h425ae33e, 32'hc18632df, 32'h42919e2e, 32'hc25d49fe, 32'hbeea1214, 32'hc28bc616};
test_output[1208:1215] = '{32'h41e4c32c, 32'h0, 32'h425ae33e, 32'h0, 32'h42919e2e, 32'h0, 32'h0, 32'h0};
test_input[1216:1223] = '{32'h426e0090, 32'h41157341, 32'h42c741ca, 32'hc26b7b8f, 32'h42202103, 32'h428171c2, 32'hc244c5c9, 32'h429c199c};
test_output[1216:1223] = '{32'h426e0090, 32'h41157341, 32'h42c741ca, 32'h0, 32'h42202103, 32'h428171c2, 32'h0, 32'h429c199c};
test_input[1224:1231] = '{32'hc0661606, 32'hc2a7658d, 32'hc229c6c6, 32'h4244c9c1, 32'hc26ab668, 32'h429cd326, 32'hc26f6f0b, 32'h429c6a32};
test_output[1224:1231] = '{32'h0, 32'h0, 32'h0, 32'h4244c9c1, 32'h0, 32'h429cd326, 32'h0, 32'h429c6a32};
test_input[1232:1239] = '{32'h423b9096, 32'hc1ba393d, 32'hc2443bae, 32'hc229bf11, 32'hc27cfd82, 32'h41d707dd, 32'hc2a9eef9, 32'hc116acd5};
test_output[1232:1239] = '{32'h423b9096, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41d707dd, 32'h0, 32'h0};
test_input[1240:1247] = '{32'h4200d62e, 32'h4297aae6, 32'h41d28def, 32'h4188bbab, 32'hc21cc4a3, 32'hc1d04915, 32'h418362fd, 32'h4143a785};
test_output[1240:1247] = '{32'h4200d62e, 32'h4297aae6, 32'h41d28def, 32'h4188bbab, 32'h0, 32'h0, 32'h418362fd, 32'h4143a785};
test_input[1248:1255] = '{32'hc2a55769, 32'h416e1d96, 32'hc0e03c61, 32'hc0c109f6, 32'hc28b7c81, 32'h42aff03d, 32'h41992e24, 32'h427aaead};
test_output[1248:1255] = '{32'h0, 32'h416e1d96, 32'h0, 32'h0, 32'h0, 32'h42aff03d, 32'h41992e24, 32'h427aaead};
test_input[1256:1263] = '{32'h4290b4e9, 32'h4211a81d, 32'hc1d73d57, 32'h42817f7a, 32'hc0079a69, 32'hc2804287, 32'hc2750a42, 32'hc28dca40};
test_output[1256:1263] = '{32'h4290b4e9, 32'h4211a81d, 32'h0, 32'h42817f7a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1264:1271] = '{32'hc238906f, 32'hc27d4f43, 32'hc2bd2890, 32'hc214e3d2, 32'hc2588167, 32'h4250ce53, 32'hc28a006f, 32'hc28f9880};
test_output[1264:1271] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4250ce53, 32'h0, 32'h0};
test_input[1272:1279] = '{32'h3fbaa381, 32'hc24e30bf, 32'h402d2b60, 32'h429f9bd2, 32'h421b776d, 32'h41e1aea2, 32'hc1c03a74, 32'hc222953c};
test_output[1272:1279] = '{32'h3fbaa381, 32'h0, 32'h402d2b60, 32'h429f9bd2, 32'h421b776d, 32'h41e1aea2, 32'h0, 32'h0};
test_input[1280:1287] = '{32'h41ddfcaf, 32'hc29bd043, 32'hc2357f89, 32'h425fc4bd, 32'hc240f2e3, 32'h42a887af, 32'h42adf466, 32'h428a55e1};
test_output[1280:1287] = '{32'h41ddfcaf, 32'h0, 32'h0, 32'h425fc4bd, 32'h0, 32'h42a887af, 32'h42adf466, 32'h428a55e1};
test_input[1288:1295] = '{32'hc1d6862a, 32'hc20850bf, 32'h42c589ba, 32'hc267a003, 32'hc2203612, 32'h42024a56, 32'hc28c3e21, 32'hc23687c4};
test_output[1288:1295] = '{32'h0, 32'h0, 32'h42c589ba, 32'h0, 32'h0, 32'h42024a56, 32'h0, 32'h0};
test_input[1296:1303] = '{32'hc255bf1c, 32'h41a7cfe4, 32'hc2c4414d, 32'h419caf5f, 32'h40b6b2fe, 32'hc20885a9, 32'hc1ef6cf0, 32'hc27b16e7};
test_output[1296:1303] = '{32'h0, 32'h41a7cfe4, 32'h0, 32'h419caf5f, 32'h40b6b2fe, 32'h0, 32'h0, 32'h0};
test_input[1304:1311] = '{32'hc108a6cc, 32'h429fd432, 32'hc2a6a5a6, 32'hc214f7f6, 32'h4239445b, 32'h4113c47a, 32'hc290a786, 32'h42baff85};
test_output[1304:1311] = '{32'h0, 32'h429fd432, 32'h0, 32'h0, 32'h4239445b, 32'h4113c47a, 32'h0, 32'h42baff85};
test_input[1312:1319] = '{32'hc23c7eac, 32'hc1a97702, 32'hc2a91846, 32'hc218d8fb, 32'h428a6bc5, 32'hc1fbb519, 32'h42365932, 32'hc2c04f8a};
test_output[1312:1319] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h428a6bc5, 32'h0, 32'h42365932, 32'h0};
test_input[1320:1327] = '{32'hc259775d, 32'h4258d468, 32'h42b09327, 32'h4299959a, 32'hc19b11fb, 32'hc1be745d, 32'h422547bf, 32'hc2818f45};
test_output[1320:1327] = '{32'h0, 32'h4258d468, 32'h42b09327, 32'h4299959a, 32'h0, 32'h0, 32'h422547bf, 32'h0};
test_input[1328:1335] = '{32'h426da1c3, 32'hc1dfa6bf, 32'h427012de, 32'h429100c0, 32'hc1e1b2ec, 32'hc1ec7796, 32'hc2158969, 32'h412c2d49};
test_output[1328:1335] = '{32'h426da1c3, 32'h0, 32'h427012de, 32'h429100c0, 32'h0, 32'h0, 32'h0, 32'h412c2d49};
test_input[1336:1343] = '{32'h41f0375a, 32'h42756b57, 32'hc2782675, 32'hc285fcfb, 32'hc2568835, 32'h42a359a2, 32'hc2220c8b, 32'hc261d467};
test_output[1336:1343] = '{32'h41f0375a, 32'h42756b57, 32'h0, 32'h0, 32'h0, 32'h42a359a2, 32'h0, 32'h0};
test_input[1344:1351] = '{32'h42b99574, 32'h42b69a80, 32'h42644e5f, 32'hc19dcdd6, 32'hc22a32bd, 32'hc1b80a9f, 32'hc25f6a6e, 32'hc22f0ec0};
test_output[1344:1351] = '{32'h42b99574, 32'h42b69a80, 32'h42644e5f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1352:1359] = '{32'h42b682a3, 32'h42a149d9, 32'hc19161c6, 32'hc19b9f11, 32'hc188654f, 32'h4177269b, 32'hbf1969bc, 32'h4247bbda};
test_output[1352:1359] = '{32'h42b682a3, 32'h42a149d9, 32'h0, 32'h0, 32'h0, 32'h4177269b, 32'h0, 32'h4247bbda};
test_input[1360:1367] = '{32'hc2024f05, 32'hc1ec5575, 32'hc2ad9acf, 32'h429a64c8, 32'hc225062b, 32'hc2a19c92, 32'h40e82b93, 32'h42b86fea};
test_output[1360:1367] = '{32'h0, 32'h0, 32'h0, 32'h429a64c8, 32'h0, 32'h0, 32'h40e82b93, 32'h42b86fea};
test_input[1368:1375] = '{32'hc1fa739f, 32'h419a5bfa, 32'hc2b04636, 32'hc23b8ecc, 32'hc2081c1b, 32'h4298efbb, 32'h42c71b44, 32'h42840374};
test_output[1368:1375] = '{32'h0, 32'h419a5bfa, 32'h0, 32'h0, 32'h0, 32'h4298efbb, 32'h42c71b44, 32'h42840374};
test_input[1376:1383] = '{32'hc2b0a568, 32'hc27aff3a, 32'hc25a53cf, 32'h428b0139, 32'hc164a1da, 32'hc2a8cf61, 32'h427ca15a, 32'h413210a2};
test_output[1376:1383] = '{32'h0, 32'h0, 32'h0, 32'h428b0139, 32'h0, 32'h0, 32'h427ca15a, 32'h413210a2};
test_input[1384:1391] = '{32'h42bd2ec6, 32'hc2550731, 32'hc216eed9, 32'h4100c8a0, 32'h42a910f9, 32'h40b00436, 32'hc1773363, 32'h418bc9f8};
test_output[1384:1391] = '{32'h42bd2ec6, 32'h0, 32'h0, 32'h4100c8a0, 32'h42a910f9, 32'h40b00436, 32'h0, 32'h418bc9f8};
test_input[1392:1399] = '{32'hc087f720, 32'h4264425c, 32'hc20ee731, 32'hc2a7916a, 32'h4122f582, 32'h40e8ef68, 32'hc1ad4d5a, 32'h4280b5b3};
test_output[1392:1399] = '{32'h0, 32'h4264425c, 32'h0, 32'h0, 32'h4122f582, 32'h40e8ef68, 32'h0, 32'h4280b5b3};
test_input[1400:1407] = '{32'hc1ac1c86, 32'hc2984d93, 32'h41b56a92, 32'hc29f1d00, 32'h41c9ed73, 32'h4109a174, 32'hc124c5d2, 32'h41a1a332};
test_output[1400:1407] = '{32'h0, 32'h0, 32'h41b56a92, 32'h0, 32'h41c9ed73, 32'h4109a174, 32'h0, 32'h41a1a332};
test_input[1408:1415] = '{32'h428ce97f, 32'hc16d5d5e, 32'h4027c60b, 32'hc20e21ca, 32'h41cc1f89, 32'h42b48010, 32'h42a800f1, 32'h42408a46};
test_output[1408:1415] = '{32'h428ce97f, 32'h0, 32'h4027c60b, 32'h0, 32'h41cc1f89, 32'h42b48010, 32'h42a800f1, 32'h42408a46};
test_input[1416:1423] = '{32'hc22e1e60, 32'h41c6fd29, 32'hc229c302, 32'h4198baa2, 32'h42a64008, 32'hc271505d, 32'h42bc9785, 32'h421c346f};
test_output[1416:1423] = '{32'h0, 32'h41c6fd29, 32'h0, 32'h4198baa2, 32'h42a64008, 32'h0, 32'h42bc9785, 32'h421c346f};
test_input[1424:1431] = '{32'h41c68d1b, 32'h42af7e9a, 32'h411889ca, 32'h423a8f33, 32'h42a60b40, 32'h424f1d97, 32'h428e88f2, 32'hc28e8074};
test_output[1424:1431] = '{32'h41c68d1b, 32'h42af7e9a, 32'h411889ca, 32'h423a8f33, 32'h42a60b40, 32'h424f1d97, 32'h428e88f2, 32'h0};
test_input[1432:1439] = '{32'h42b75fc3, 32'hc28b77a3, 32'hc22a33fa, 32'h428aa6de, 32'h42c520a4, 32'hc2bfcf55, 32'h429aa139, 32'h426b9870};
test_output[1432:1439] = '{32'h42b75fc3, 32'h0, 32'h0, 32'h428aa6de, 32'h42c520a4, 32'h0, 32'h429aa139, 32'h426b9870};
test_input[1440:1447] = '{32'hc24b6c51, 32'hc21535aa, 32'hc1a57e64, 32'hc29eb834, 32'h3fe46bf5, 32'h429192ca, 32'hc2675afb, 32'h42ac07f4};
test_output[1440:1447] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h3fe46bf5, 32'h429192ca, 32'h0, 32'h42ac07f4};
test_input[1448:1455] = '{32'h3efd08ea, 32'hc299fa2f, 32'hc27500fd, 32'hc29833a5, 32'h4287b2e9, 32'h417efdb0, 32'h424979e6, 32'hc1a58bda};
test_output[1448:1455] = '{32'h3efd08ea, 32'h0, 32'h0, 32'h0, 32'h4287b2e9, 32'h417efdb0, 32'h424979e6, 32'h0};
test_input[1456:1463] = '{32'h4285949f, 32'h428ca435, 32'hc24c0dad, 32'h42523df7, 32'h42014f1d, 32'hc148d026, 32'hc29877d3, 32'hc2a75558};
test_output[1456:1463] = '{32'h4285949f, 32'h428ca435, 32'h0, 32'h42523df7, 32'h42014f1d, 32'h0, 32'h0, 32'h0};
test_input[1464:1471] = '{32'h42c44bcb, 32'h42c72a51, 32'h41ebad80, 32'hbd97e084, 32'hc27224f9, 32'hc294fe67, 32'h41c1f26e, 32'h3fb24fc3};
test_output[1464:1471] = '{32'h42c44bcb, 32'h42c72a51, 32'h41ebad80, 32'h0, 32'h0, 32'h0, 32'h41c1f26e, 32'h3fb24fc3};
test_input[1472:1479] = '{32'h42780f44, 32'h42b3f3f0, 32'h41d9926a, 32'h428b1198, 32'hc2b8fb46, 32'hc1a7277d, 32'h401a07a7, 32'h428e91ab};
test_output[1472:1479] = '{32'h42780f44, 32'h42b3f3f0, 32'h41d9926a, 32'h428b1198, 32'h0, 32'h0, 32'h401a07a7, 32'h428e91ab};
test_input[1480:1487] = '{32'hc1773344, 32'h42c59f76, 32'h42ba645f, 32'h428ed027, 32'hc1954e59, 32'hc283eecb, 32'hc298368e, 32'hc2845b0b};
test_output[1480:1487] = '{32'h0, 32'h42c59f76, 32'h42ba645f, 32'h428ed027, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1488:1495] = '{32'h4130cebb, 32'h429bbeaa, 32'h41a81936, 32'h4165ee22, 32'h416bf99a, 32'h4177afab, 32'hc263067b, 32'hc23a67e6};
test_output[1488:1495] = '{32'h4130cebb, 32'h429bbeaa, 32'h41a81936, 32'h4165ee22, 32'h416bf99a, 32'h4177afab, 32'h0, 32'h0};
test_input[1496:1503] = '{32'hc11b0f23, 32'h41952a09, 32'hc20b516f, 32'h4283dd6b, 32'h423bd7a5, 32'hc229aa56, 32'h428a1452, 32'h4280fc07};
test_output[1496:1503] = '{32'h0, 32'h41952a09, 32'h0, 32'h4283dd6b, 32'h423bd7a5, 32'h0, 32'h428a1452, 32'h4280fc07};
test_input[1504:1511] = '{32'hc28a89f2, 32'h4223b96d, 32'hc24db17a, 32'h4296c05d, 32'hc18b454e, 32'hc26a7dcb, 32'hc29df961, 32'h42b145f1};
test_output[1504:1511] = '{32'h0, 32'h4223b96d, 32'h0, 32'h4296c05d, 32'h0, 32'h0, 32'h0, 32'h42b145f1};
test_input[1512:1519] = '{32'hc1eb7f33, 32'h41ef1229, 32'hc29a90e3, 32'h4277e14f, 32'hc1215cd4, 32'h4259275f, 32'h4186d1e5, 32'h3fa352b8};
test_output[1512:1519] = '{32'h0, 32'h41ef1229, 32'h0, 32'h4277e14f, 32'h0, 32'h4259275f, 32'h4186d1e5, 32'h3fa352b8};
test_input[1520:1527] = '{32'h42567cc0, 32'h42a5cbdf, 32'hc281e39b, 32'h41ed8b83, 32'h415063e5, 32'hc18b6b3a, 32'h42445504, 32'hc202935f};
test_output[1520:1527] = '{32'h42567cc0, 32'h42a5cbdf, 32'h0, 32'h41ed8b83, 32'h415063e5, 32'h0, 32'h42445504, 32'h0};
test_input[1528:1535] = '{32'h42191622, 32'h428497ed, 32'hc29a84d5, 32'h41ba3d7d, 32'hc2733c9a, 32'h41ef0157, 32'h42bf9133, 32'h4244e399};
test_output[1528:1535] = '{32'h42191622, 32'h428497ed, 32'h0, 32'h41ba3d7d, 32'h0, 32'h41ef0157, 32'h42bf9133, 32'h4244e399};
test_input[1536:1543] = '{32'h419ba963, 32'h42c0e260, 32'h4235efd5, 32'hc2bc0684, 32'h422b4989, 32'hc27ea07b, 32'hc2b5f822, 32'h41be0043};
test_output[1536:1543] = '{32'h419ba963, 32'h42c0e260, 32'h4235efd5, 32'h0, 32'h422b4989, 32'h0, 32'h0, 32'h41be0043};
test_input[1544:1551] = '{32'h42454220, 32'hc115a0df, 32'h42192cb3, 32'h424a95f9, 32'h42210c0d, 32'h40bed0d1, 32'h427c2793, 32'h428839c8};
test_output[1544:1551] = '{32'h42454220, 32'h0, 32'h42192cb3, 32'h424a95f9, 32'h42210c0d, 32'h40bed0d1, 32'h427c2793, 32'h428839c8};
test_input[1552:1559] = '{32'hc2a69b3a, 32'hc27f4e5f, 32'h41ed8006, 32'h41c665a0, 32'h41457277, 32'h42bb1e1f, 32'hc206786e, 32'hc23bffc7};
test_output[1552:1559] = '{32'h0, 32'h0, 32'h41ed8006, 32'h41c665a0, 32'h41457277, 32'h42bb1e1f, 32'h0, 32'h0};
test_input[1560:1567] = '{32'h419acf54, 32'hc2a35876, 32'h426e4299, 32'h424c8fc9, 32'h3f811f08, 32'h42970e30, 32'h42a77620, 32'h41b0e7d9};
test_output[1560:1567] = '{32'h419acf54, 32'h0, 32'h426e4299, 32'h424c8fc9, 32'h3f811f08, 32'h42970e30, 32'h42a77620, 32'h41b0e7d9};
test_input[1568:1575] = '{32'hc19babd2, 32'h4174edf1, 32'h419b024c, 32'hc284987c, 32'h42188c06, 32'h429691b7, 32'h428fbeca, 32'hc18a0ee8};
test_output[1568:1575] = '{32'h0, 32'h4174edf1, 32'h419b024c, 32'h0, 32'h42188c06, 32'h429691b7, 32'h428fbeca, 32'h0};
test_input[1576:1583] = '{32'h420610c7, 32'hc2b2e428, 32'h418c23a6, 32'hc2753883, 32'hc28e9b7d, 32'h42858970, 32'h4288f5b0, 32'hc2b3bdff};
test_output[1576:1583] = '{32'h420610c7, 32'h0, 32'h418c23a6, 32'h0, 32'h0, 32'h42858970, 32'h4288f5b0, 32'h0};
test_input[1584:1591] = '{32'hc2998cd0, 32'hc234a86a, 32'hc2b27914, 32'hc1ef4ae5, 32'hc0b57ab6, 32'h41ef3410, 32'hc22d4aa6, 32'h41e3dfdc};
test_output[1584:1591] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ef3410, 32'h0, 32'h41e3dfdc};
test_input[1592:1599] = '{32'hc14640b6, 32'h41a7c474, 32'h41ef766b, 32'hc291bd24, 32'hc211125d, 32'hc0917bc2, 32'hc1d9cbcd, 32'h3fa40caf};
test_output[1592:1599] = '{32'h0, 32'h41a7c474, 32'h41ef766b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3fa40caf};
test_input[1600:1607] = '{32'h427e300f, 32'hc2424061, 32'hc17c8803, 32'hc2a15951, 32'hc1237920, 32'hc1b45271, 32'h41f7df0d, 32'hbf4c97ca};
test_output[1600:1607] = '{32'h427e300f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f7df0d, 32'h0};
test_input[1608:1615] = '{32'h425c5c30, 32'h425edd72, 32'hc1fb5af7, 32'hc2b058fe, 32'hc0f43b80, 32'h42ba2ac9, 32'h42732c5d, 32'h429c8f44};
test_output[1608:1615] = '{32'h425c5c30, 32'h425edd72, 32'h0, 32'h0, 32'h0, 32'h42ba2ac9, 32'h42732c5d, 32'h429c8f44};
test_input[1616:1623] = '{32'h41aff2ef, 32'hc2ba33cf, 32'hc2b9c04e, 32'hc1f0b7d5, 32'h42229d60, 32'h420156bf, 32'hc2139e48, 32'h41645a02};
test_output[1616:1623] = '{32'h41aff2ef, 32'h0, 32'h0, 32'h0, 32'h42229d60, 32'h420156bf, 32'h0, 32'h41645a02};
test_input[1624:1631] = '{32'hc2bb1815, 32'hbf1c396f, 32'hc28b4406, 32'hc1452b0b, 32'hc2101aa1, 32'h415df693, 32'h42a78bc2, 32'h426c83bd};
test_output[1624:1631] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h415df693, 32'h42a78bc2, 32'h426c83bd};
test_input[1632:1639] = '{32'hc256ca84, 32'h42ab2bef, 32'h42c0c6ca, 32'h42b3d5c6, 32'h42c4e3e4, 32'h41ed8cdf, 32'h42c006b7, 32'hc20434bb};
test_output[1632:1639] = '{32'h0, 32'h42ab2bef, 32'h42c0c6ca, 32'h42b3d5c6, 32'h42c4e3e4, 32'h41ed8cdf, 32'h42c006b7, 32'h0};
test_input[1640:1647] = '{32'hc2bbf409, 32'hc0bb232c, 32'hc2b585cb, 32'h41b8b739, 32'hc2c42392, 32'h3f4dac99, 32'hc2beed19, 32'h42571065};
test_output[1640:1647] = '{32'h0, 32'h0, 32'h0, 32'h41b8b739, 32'h0, 32'h3f4dac99, 32'h0, 32'h42571065};
test_input[1648:1655] = '{32'h4286a7e1, 32'hc20da43b, 32'hc000eb27, 32'hc299fbed, 32'h42499ee5, 32'h42b5ea53, 32'h427979af, 32'h4221be9b};
test_output[1648:1655] = '{32'h4286a7e1, 32'h0, 32'h0, 32'h0, 32'h42499ee5, 32'h42b5ea53, 32'h427979af, 32'h4221be9b};
test_input[1656:1663] = '{32'h40c68c24, 32'h42a68d91, 32'hc2adaf43, 32'h41fc0939, 32'h42a6d963, 32'h41f77993, 32'h423c9525, 32'hc2c47a44};
test_output[1656:1663] = '{32'h40c68c24, 32'h42a68d91, 32'h0, 32'h41fc0939, 32'h42a6d963, 32'h41f77993, 32'h423c9525, 32'h0};
test_input[1664:1671] = '{32'h429769dd, 32'hc192121c, 32'hc120dddd, 32'hc189eaa8, 32'hc1be3c19, 32'hc23c218f, 32'hc18e40a2, 32'hc21a4346};
test_output[1664:1671] = '{32'h429769dd, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1672:1679] = '{32'h42426262, 32'h42af3e3b, 32'h428fd06a, 32'h42bee932, 32'h41dfaedf, 32'hc2a492f5, 32'h4209e695, 32'h42c2fb50};
test_output[1672:1679] = '{32'h42426262, 32'h42af3e3b, 32'h428fd06a, 32'h42bee932, 32'h41dfaedf, 32'h0, 32'h4209e695, 32'h42c2fb50};
test_input[1680:1687] = '{32'hc2a4c401, 32'hc1ac7b3d, 32'hc123abde, 32'hc2ae56f4, 32'h427f1cda, 32'h41f8c71c, 32'hc2412c1d, 32'h40e13b21};
test_output[1680:1687] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h427f1cda, 32'h41f8c71c, 32'h0, 32'h40e13b21};
test_input[1688:1695] = '{32'h42aec37f, 32'h42c2b057, 32'hc15efc09, 32'h41026425, 32'h3f2da239, 32'hc25eda2a, 32'hc2c70067, 32'h42732018};
test_output[1688:1695] = '{32'h42aec37f, 32'h42c2b057, 32'h0, 32'h41026425, 32'h3f2da239, 32'h0, 32'h0, 32'h42732018};
test_input[1696:1703] = '{32'h4299b55c, 32'hc25edd9d, 32'h41392b74, 32'h425dcaeb, 32'hc2636b11, 32'hc2bf7fb6, 32'h41abc198, 32'h426ff4b9};
test_output[1696:1703] = '{32'h4299b55c, 32'h0, 32'h41392b74, 32'h425dcaeb, 32'h0, 32'h0, 32'h41abc198, 32'h426ff4b9};
test_input[1704:1711] = '{32'h42be773e, 32'h411a67cc, 32'hc0108394, 32'h42588478, 32'hc1221d48, 32'h421acc25, 32'hc0b63522, 32'hc2371f04};
test_output[1704:1711] = '{32'h42be773e, 32'h411a67cc, 32'h0, 32'h42588478, 32'h0, 32'h421acc25, 32'h0, 32'h0};
test_input[1712:1719] = '{32'hc2792a38, 32'h41ce04f4, 32'h4212de03, 32'hc1ed768e, 32'h41224789, 32'h405459eb, 32'hc2c19aad, 32'hc181ae49};
test_output[1712:1719] = '{32'h0, 32'h41ce04f4, 32'h4212de03, 32'h0, 32'h41224789, 32'h405459eb, 32'h0, 32'h0};
test_input[1720:1727] = '{32'hc2939226, 32'h428474c6, 32'hc229b6dd, 32'h426e3dd2, 32'hc1a87cec, 32'hc286ee5e, 32'hc255c365, 32'h413b20a2};
test_output[1720:1727] = '{32'h0, 32'h428474c6, 32'h0, 32'h426e3dd2, 32'h0, 32'h0, 32'h0, 32'h413b20a2};
test_input[1728:1735] = '{32'hc2554613, 32'hc262b823, 32'h4188edad, 32'hc2b237a7, 32'h42ab6ed9, 32'hc2b546e7, 32'h42aaa1f4, 32'h4282e46f};
test_output[1728:1735] = '{32'h0, 32'h0, 32'h4188edad, 32'h0, 32'h42ab6ed9, 32'h0, 32'h42aaa1f4, 32'h4282e46f};
test_input[1736:1743] = '{32'h416f1a25, 32'h41ca0b0f, 32'hc2c7bd27, 32'h42048294, 32'hc2256176, 32'h40bb6675, 32'h4204fac4, 32'h41bad717};
test_output[1736:1743] = '{32'h416f1a25, 32'h41ca0b0f, 32'h0, 32'h42048294, 32'h0, 32'h40bb6675, 32'h4204fac4, 32'h41bad717};
test_input[1744:1751] = '{32'h42552b72, 32'hc235da98, 32'h4109ad87, 32'hc1b2327c, 32'hc228d98f, 32'h409030a0, 32'hc2478003, 32'h418e2ba7};
test_output[1744:1751] = '{32'h42552b72, 32'h0, 32'h4109ad87, 32'h0, 32'h0, 32'h409030a0, 32'h0, 32'h418e2ba7};
test_input[1752:1759] = '{32'h421b69de, 32'h428f4bd4, 32'hc215fb08, 32'h41cefca7, 32'h42b9332a, 32'hc243cca3, 32'hc2821beb, 32'h41bfb794};
test_output[1752:1759] = '{32'h421b69de, 32'h428f4bd4, 32'h0, 32'h41cefca7, 32'h42b9332a, 32'h0, 32'h0, 32'h41bfb794};
test_input[1760:1767] = '{32'h4203f0ee, 32'h42c11481, 32'h428210c1, 32'h41643991, 32'hc0b5758b, 32'h4280b430, 32'h42202d50, 32'h4180f3d9};
test_output[1760:1767] = '{32'h4203f0ee, 32'h42c11481, 32'h428210c1, 32'h41643991, 32'h0, 32'h4280b430, 32'h42202d50, 32'h4180f3d9};
test_input[1768:1775] = '{32'h42057d8d, 32'h421d9d86, 32'hc278109c, 32'hc0bab9a9, 32'hc2a12b75, 32'hc2759dd6, 32'h42a30591, 32'h42b53c1f};
test_output[1768:1775] = '{32'h42057d8d, 32'h421d9d86, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a30591, 32'h42b53c1f};
test_input[1776:1783] = '{32'h4270b6a3, 32'h41b18efe, 32'h41fdfa4f, 32'h42aedde8, 32'h41ee7db4, 32'h41aa7da0, 32'h4186cc25, 32'h410192a2};
test_output[1776:1783] = '{32'h4270b6a3, 32'h41b18efe, 32'h41fdfa4f, 32'h42aedde8, 32'h41ee7db4, 32'h41aa7da0, 32'h4186cc25, 32'h410192a2};
test_input[1784:1791] = '{32'h42290905, 32'h40300787, 32'h4107451a, 32'h429dfe47, 32'h42663ba1, 32'h40e70725, 32'h41810c2d, 32'h41577ede};
test_output[1784:1791] = '{32'h42290905, 32'h40300787, 32'h4107451a, 32'h429dfe47, 32'h42663ba1, 32'h40e70725, 32'h41810c2d, 32'h41577ede};
test_input[1792:1799] = '{32'h423121d2, 32'h422fb3e3, 32'hc2bd7c55, 32'h429cb03a, 32'h419dd1dc, 32'h41c732cd, 32'h42359d1d, 32'hc236c2e3};
test_output[1792:1799] = '{32'h423121d2, 32'h422fb3e3, 32'h0, 32'h429cb03a, 32'h419dd1dc, 32'h41c732cd, 32'h42359d1d, 32'h0};
test_input[1800:1807] = '{32'hc1aab248, 32'h415d9ab5, 32'h41c59f8f, 32'hc2a922b4, 32'h42c1e7f6, 32'h413e8330, 32'h423b10e1, 32'h3f806156};
test_output[1800:1807] = '{32'h0, 32'h415d9ab5, 32'h41c59f8f, 32'h0, 32'h42c1e7f6, 32'h413e8330, 32'h423b10e1, 32'h3f806156};
test_input[1808:1815] = '{32'h4278e9d1, 32'h424f8296, 32'hc2a5c135, 32'hc1f4d274, 32'h42173865, 32'hc23dfdb9, 32'hc27dd7e7, 32'hc1bd3c03};
test_output[1808:1815] = '{32'h4278e9d1, 32'h424f8296, 32'h0, 32'h0, 32'h42173865, 32'h0, 32'h0, 32'h0};
test_input[1816:1823] = '{32'hc2a00c16, 32'hc2c0ea29, 32'hc25db58a, 32'hc2bd19b3, 32'h428c5164, 32'hc05d451f, 32'h4232e747, 32'hc29cf369};
test_output[1816:1823] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h428c5164, 32'h0, 32'h4232e747, 32'h0};
test_input[1824:1831] = '{32'hc229e0f6, 32'hc12ec29f, 32'hc252e2fb, 32'hc269ec9e, 32'h41f27760, 32'hc1e5c652, 32'h42159413, 32'hc1a36ce6};
test_output[1824:1831] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41f27760, 32'h0, 32'h42159413, 32'h0};
test_input[1832:1839] = '{32'hc2b5a0b3, 32'h3fcdc473, 32'h4232a226, 32'h426610db, 32'h429ac33e, 32'hc296e24e, 32'h424a7143, 32'h41fe276f};
test_output[1832:1839] = '{32'h0, 32'h3fcdc473, 32'h4232a226, 32'h426610db, 32'h429ac33e, 32'h0, 32'h424a7143, 32'h41fe276f};
test_input[1840:1847] = '{32'h414b8973, 32'h40340c2f, 32'hc2958590, 32'h41fdc68c, 32'h42024910, 32'h42378b1f, 32'hc2826375, 32'h41f387c7};
test_output[1840:1847] = '{32'h414b8973, 32'h40340c2f, 32'h0, 32'h41fdc68c, 32'h42024910, 32'h42378b1f, 32'h0, 32'h41f387c7};
test_input[1848:1855] = '{32'h422260cc, 32'hc28e93b1, 32'h42bae2b8, 32'hc108f5a4, 32'hc283f780, 32'h41be904c, 32'hc2992d0b, 32'hc1f516c5};
test_output[1848:1855] = '{32'h422260cc, 32'h0, 32'h42bae2b8, 32'h0, 32'h0, 32'h41be904c, 32'h0, 32'h0};
test_input[1856:1863] = '{32'hc2924ba2, 32'h41f9382d, 32'h42c55c38, 32'hc216f113, 32'h414a3ed7, 32'h4095d444, 32'h42a12440, 32'hc193e2da};
test_output[1856:1863] = '{32'h0, 32'h41f9382d, 32'h42c55c38, 32'h0, 32'h414a3ed7, 32'h4095d444, 32'h42a12440, 32'h0};
test_input[1864:1871] = '{32'hc201648a, 32'hc2aecc87, 32'h4222772b, 32'hc1133d2d, 32'hc1a9aecb, 32'hc1c62edc, 32'h40eb96d9, 32'h4154762e};
test_output[1864:1871] = '{32'h0, 32'h0, 32'h4222772b, 32'h0, 32'h0, 32'h0, 32'h40eb96d9, 32'h4154762e};
test_input[1872:1879] = '{32'h416c9ee7, 32'hc29cd45e, 32'hc22dd74c, 32'h426f8736, 32'h42029558, 32'h42944b76, 32'h4214a776, 32'hc28a61b8};
test_output[1872:1879] = '{32'h416c9ee7, 32'h0, 32'h0, 32'h426f8736, 32'h42029558, 32'h42944b76, 32'h4214a776, 32'h0};
test_input[1880:1887] = '{32'h4180cbfa, 32'hc2bdd587, 32'h42562019, 32'hc10b0715, 32'hc2622e1c, 32'h4237ed24, 32'hc2409631, 32'hc24d610f};
test_output[1880:1887] = '{32'h4180cbfa, 32'h0, 32'h42562019, 32'h0, 32'h0, 32'h4237ed24, 32'h0, 32'h0};
test_input[1888:1895] = '{32'hc29d791c, 32'hc2be3358, 32'h41097dee, 32'hc21b0770, 32'hc26bb955, 32'hc2b23e02, 32'hc26786a6, 32'hc282f0ac};
test_output[1888:1895] = '{32'h0, 32'h0, 32'h41097dee, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1896:1903] = '{32'hbff93a54, 32'h420d9ed3, 32'hc1978dc1, 32'hc2c552dd, 32'h42861e56, 32'h42c6f14d, 32'h42a4e252, 32'h4278274a};
test_output[1896:1903] = '{32'h0, 32'h420d9ed3, 32'h0, 32'h0, 32'h42861e56, 32'h42c6f14d, 32'h42a4e252, 32'h4278274a};
test_input[1904:1911] = '{32'h42b28a73, 32'h41592f01, 32'hbd992243, 32'hc1aebeba, 32'h41fa474f, 32'hc223e2ee, 32'h42c79b99, 32'hc1a40865};
test_output[1904:1911] = '{32'h42b28a73, 32'h41592f01, 32'h0, 32'h0, 32'h41fa474f, 32'h0, 32'h42c79b99, 32'h0};
test_input[1912:1919] = '{32'h42b7683c, 32'h429e9754, 32'hc297d677, 32'hc2065562, 32'h427ddf8c, 32'h41f7caa1, 32'h42624742, 32'h40900a57};
test_output[1912:1919] = '{32'h42b7683c, 32'h429e9754, 32'h0, 32'h0, 32'h427ddf8c, 32'h41f7caa1, 32'h42624742, 32'h40900a57};
test_input[1920:1927] = '{32'hc0f78c7f, 32'h3f6b04dc, 32'hbe958f0e, 32'h42110fe0, 32'hc2ac1885, 32'h428d810c, 32'hc1318047, 32'h42bd02c5};
test_output[1920:1927] = '{32'h0, 32'h3f6b04dc, 32'h0, 32'h42110fe0, 32'h0, 32'h428d810c, 32'h0, 32'h42bd02c5};
test_input[1928:1935] = '{32'h402bc66b, 32'h41fcd877, 32'hc105783d, 32'hbf64afc6, 32'hc2a36283, 32'h42862064, 32'hc1f507fe, 32'h429c4f28};
test_output[1928:1935] = '{32'h402bc66b, 32'h41fcd877, 32'h0, 32'h0, 32'h0, 32'h42862064, 32'h0, 32'h429c4f28};
test_input[1936:1943] = '{32'h42888213, 32'h42ab9876, 32'hc28ee708, 32'h418b5ad0, 32'hc0892552, 32'hc2a63eef, 32'hc284f1bb, 32'hbfbae434};
test_output[1936:1943] = '{32'h42888213, 32'h42ab9876, 32'h0, 32'h418b5ad0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1944:1951] = '{32'hc284c795, 32'hc2603d85, 32'h4211eb4d, 32'h42764963, 32'h42c32df6, 32'h423f13fb, 32'h4201dff4, 32'h42ac9a53};
test_output[1944:1951] = '{32'h0, 32'h0, 32'h4211eb4d, 32'h42764963, 32'h42c32df6, 32'h423f13fb, 32'h4201dff4, 32'h42ac9a53};
test_input[1952:1959] = '{32'hc2b6ca95, 32'h422d91ed, 32'h42a9b93b, 32'h42b250bf, 32'hc2a47cca, 32'h4250a2b3, 32'h421514b5, 32'h42297ee0};
test_output[1952:1959] = '{32'h0, 32'h422d91ed, 32'h42a9b93b, 32'h42b250bf, 32'h0, 32'h4250a2b3, 32'h421514b5, 32'h42297ee0};
test_input[1960:1967] = '{32'h429a1fde, 32'hc15d191d, 32'hc186e960, 32'hc2c2f02f, 32'hc29042b8, 32'hc121eaf7, 32'hc134fdb4, 32'hc2428f02};
test_output[1960:1967] = '{32'h429a1fde, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1968:1975] = '{32'h4195592e, 32'hc0643ccb, 32'h421e4066, 32'h418dcda5, 32'h42c6b797, 32'h41d0f5ea, 32'hc0f1fbcb, 32'h421dae37};
test_output[1968:1975] = '{32'h4195592e, 32'h0, 32'h421e4066, 32'h418dcda5, 32'h42c6b797, 32'h41d0f5ea, 32'h0, 32'h421dae37};
test_input[1976:1983] = '{32'h42496352, 32'hc2a9f9b4, 32'h429aed42, 32'h4286c833, 32'hc28ead80, 32'h40ab1e82, 32'hc0679686, 32'hc2c21970};
test_output[1976:1983] = '{32'h42496352, 32'h0, 32'h429aed42, 32'h4286c833, 32'h0, 32'h40ab1e82, 32'h0, 32'h0};
test_input[1984:1991] = '{32'h413ba27d, 32'h41a40abb, 32'h4292fefb, 32'h42a58f46, 32'hc04f7885, 32'hc1f10d44, 32'h42adadc5, 32'hc23ca5cb};
test_output[1984:1991] = '{32'h413ba27d, 32'h41a40abb, 32'h4292fefb, 32'h42a58f46, 32'h0, 32'h0, 32'h42adadc5, 32'h0};
test_input[1992:1999] = '{32'h4192d189, 32'hc2ae9b86, 32'h42834c0c, 32'hc23d6bd9, 32'h42b0e02b, 32'h410f411f, 32'h41e58055, 32'hc2168c36};
test_output[1992:1999] = '{32'h4192d189, 32'h0, 32'h42834c0c, 32'h0, 32'h42b0e02b, 32'h410f411f, 32'h41e58055, 32'h0};
test_input[2000:2007] = '{32'hc27dd07c, 32'hc2195476, 32'hc28bdd72, 32'h42632bdc, 32'hc26b2dda, 32'h428146e3, 32'h4263ea34, 32'h42a514d9};
test_output[2000:2007] = '{32'h0, 32'h0, 32'h0, 32'h42632bdc, 32'h0, 32'h428146e3, 32'h4263ea34, 32'h42a514d9};
test_input[2008:2015] = '{32'h42bc0e7b, 32'hc22e280e, 32'hc23e26bd, 32'hc00a1db2, 32'hc20dbfdc, 32'hc28ac383, 32'h42a8f3e1, 32'hc2b0438f};
test_output[2008:2015] = '{32'h42bc0e7b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a8f3e1, 32'h0};
test_input[2016:2023] = '{32'h419bef61, 32'hc20aa218, 32'h427b8ed9, 32'hc2924ac1, 32'hc209bd44, 32'h423f368b, 32'h4207e5cf, 32'hc272d76a};
test_output[2016:2023] = '{32'h419bef61, 32'h0, 32'h427b8ed9, 32'h0, 32'h0, 32'h423f368b, 32'h4207e5cf, 32'h0};
test_input[2024:2031] = '{32'hc2c63828, 32'hc07690b7, 32'h42037351, 32'h40e692ac, 32'hc245c6b1, 32'h4153d5f1, 32'h42bbd01a, 32'hc2439ef0};
test_output[2024:2031] = '{32'h0, 32'h0, 32'h42037351, 32'h40e692ac, 32'h0, 32'h4153d5f1, 32'h42bbd01a, 32'h0};
test_input[2032:2039] = '{32'hc07e686c, 32'hc19ce695, 32'h41f95342, 32'h4203868e, 32'h4121a09f, 32'hc2b7f10a, 32'h41862081, 32'hc089bc81};
test_output[2032:2039] = '{32'h0, 32'h0, 32'h41f95342, 32'h4203868e, 32'h4121a09f, 32'h0, 32'h41862081, 32'h0};
test_input[2040:2047] = '{32'hc17ce42d, 32'h42a93487, 32'h401448ec, 32'hc248c494, 32'h422b6889, 32'hc24d830b, 32'hc2b6e80c, 32'hc12f5b07};
test_output[2040:2047] = '{32'h0, 32'h42a93487, 32'h401448ec, 32'h0, 32'h422b6889, 32'h0, 32'h0, 32'h0};
test_input[2048:2055] = '{32'hc1a67767, 32'hc295f554, 32'h418520cb, 32'h428cbb66, 32'hc2359b0c, 32'hc232367c, 32'h4177f1ed, 32'h42c23af5};
test_output[2048:2055] = '{32'h0, 32'h0, 32'h418520cb, 32'h428cbb66, 32'h0, 32'h0, 32'h4177f1ed, 32'h42c23af5};
test_input[2056:2063] = '{32'h416fe0fc, 32'hc239eb6b, 32'h423221d9, 32'h42c07e76, 32'hc28ba077, 32'h418386e3, 32'h428d5176, 32'h429aa096};
test_output[2056:2063] = '{32'h416fe0fc, 32'h0, 32'h423221d9, 32'h42c07e76, 32'h0, 32'h418386e3, 32'h428d5176, 32'h429aa096};
test_input[2064:2071] = '{32'h409f37da, 32'h415d4eac, 32'hc220eb2e, 32'h42c5f686, 32'hc2c3fa8e, 32'h429e5ed7, 32'h3f3ed710, 32'hc24e5e9f};
test_output[2064:2071] = '{32'h409f37da, 32'h415d4eac, 32'h0, 32'h42c5f686, 32'h0, 32'h429e5ed7, 32'h3f3ed710, 32'h0};
test_input[2072:2079] = '{32'hc2b1a20f, 32'hc29803d0, 32'h42a5a709, 32'h41f937eb, 32'h426676b0, 32'hc286e2b7, 32'h4230abe1, 32'hc2b088b6};
test_output[2072:2079] = '{32'h0, 32'h0, 32'h42a5a709, 32'h41f937eb, 32'h426676b0, 32'h0, 32'h4230abe1, 32'h0};
test_input[2080:2087] = '{32'hc2c53533, 32'h41d92f50, 32'h403ab145, 32'hc04eb815, 32'hc28264f9, 32'hbf713143, 32'h4255d9ed, 32'hc28978cd};
test_output[2080:2087] = '{32'h0, 32'h41d92f50, 32'h403ab145, 32'h0, 32'h0, 32'h0, 32'h4255d9ed, 32'h0};
test_input[2088:2095] = '{32'h426862b6, 32'hc2226ad1, 32'h42829e62, 32'hc1b4fad0, 32'h4204dd46, 32'hc137049e, 32'hc20a58de, 32'h42a41fe5};
test_output[2088:2095] = '{32'h426862b6, 32'h0, 32'h42829e62, 32'h0, 32'h4204dd46, 32'h0, 32'h0, 32'h42a41fe5};
test_input[2096:2103] = '{32'h423fd197, 32'hc2256d6d, 32'h42883e60, 32'hc12d0c78, 32'h42b8da3b, 32'hc22ecd2b, 32'h41e0f757, 32'hc2b44aeb};
test_output[2096:2103] = '{32'h423fd197, 32'h0, 32'h42883e60, 32'h0, 32'h42b8da3b, 32'h0, 32'h41e0f757, 32'h0};
test_input[2104:2111] = '{32'hc2b7d28c, 32'h41f84d3a, 32'hc255aefd, 32'hc258f108, 32'h42736d20, 32'hc2680345, 32'h4140330d, 32'h42553c47};
test_output[2104:2111] = '{32'h0, 32'h41f84d3a, 32'h0, 32'h0, 32'h42736d20, 32'h0, 32'h4140330d, 32'h42553c47};
test_input[2112:2119] = '{32'h42bcf310, 32'hc2769ca4, 32'hc2b08eee, 32'hc0ea30a3, 32'h42a5c464, 32'hc261ef56, 32'hc1ff1326, 32'hc2b0cfc8};
test_output[2112:2119] = '{32'h42bcf310, 32'h0, 32'h0, 32'h0, 32'h42a5c464, 32'h0, 32'h0, 32'h0};
test_input[2120:2127] = '{32'h423eaa5f, 32'h42be5767, 32'hc1c30a1e, 32'hc2331ee1, 32'hc1f98b5b, 32'h424dfd18, 32'h41201b4f, 32'h3ffe7f95};
test_output[2120:2127] = '{32'h423eaa5f, 32'h42be5767, 32'h0, 32'h0, 32'h0, 32'h424dfd18, 32'h41201b4f, 32'h3ffe7f95};
test_input[2128:2135] = '{32'h42b9b8b2, 32'hc08af457, 32'hc17bcaa6, 32'h412be57f, 32'hc1efe124, 32'hc214da11, 32'hc2467371, 32'hc1dc0169};
test_output[2128:2135] = '{32'h42b9b8b2, 32'h0, 32'h0, 32'h412be57f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2136:2143] = '{32'hc0d33752, 32'hc1b13c02, 32'h421d9bd8, 32'hc22d48a2, 32'h42968602, 32'h42a921d7, 32'hc2a78e94, 32'h40a1bd3b};
test_output[2136:2143] = '{32'h0, 32'h0, 32'h421d9bd8, 32'h0, 32'h42968602, 32'h42a921d7, 32'h0, 32'h40a1bd3b};
test_input[2144:2151] = '{32'h40fa8a6a, 32'h4192e34b, 32'hc278fa73, 32'hc255f658, 32'h428fcb7b, 32'h4291b084, 32'h42c1f6ae, 32'hc27ccd88};
test_output[2144:2151] = '{32'h40fa8a6a, 32'h4192e34b, 32'h0, 32'h0, 32'h428fcb7b, 32'h4291b084, 32'h42c1f6ae, 32'h0};
test_input[2152:2159] = '{32'hc2a9da8d, 32'h429b7890, 32'h42777adb, 32'hc1af12a0, 32'h42871200, 32'h42a7842f, 32'h42c71323, 32'h42105c41};
test_output[2152:2159] = '{32'h0, 32'h429b7890, 32'h42777adb, 32'h0, 32'h42871200, 32'h42a7842f, 32'h42c71323, 32'h42105c41};
test_input[2160:2167] = '{32'hc28feb1e, 32'hc09a503e, 32'h418914b4, 32'h413cf159, 32'h4212416e, 32'hc10a53d4, 32'h421a5dee, 32'h413e1796};
test_output[2160:2167] = '{32'h0, 32'h0, 32'h418914b4, 32'h413cf159, 32'h4212416e, 32'h0, 32'h421a5dee, 32'h413e1796};
test_input[2168:2175] = '{32'hc20cf3bd, 32'h429f9a54, 32'hc0e21c51, 32'h42b51f88, 32'h42c2550d, 32'h4219f59e, 32'h42a1b0c2, 32'hc2865fdf};
test_output[2168:2175] = '{32'h0, 32'h429f9a54, 32'h0, 32'h42b51f88, 32'h42c2550d, 32'h4219f59e, 32'h42a1b0c2, 32'h0};
test_input[2176:2183] = '{32'hc1f6568a, 32'hc17d6ea2, 32'h421f710f, 32'h429cd063, 32'hc24d4982, 32'h42c5020a, 32'h4149825e, 32'hc2be5403};
test_output[2176:2183] = '{32'h0, 32'h0, 32'h421f710f, 32'h429cd063, 32'h0, 32'h42c5020a, 32'h4149825e, 32'h0};
test_input[2184:2191] = '{32'h423db006, 32'h41ed0de1, 32'h427b7de3, 32'hc20c8384, 32'hc2acd9eb, 32'h42911bd7, 32'hc29ade0c, 32'h42983f23};
test_output[2184:2191] = '{32'h423db006, 32'h41ed0de1, 32'h427b7de3, 32'h0, 32'h0, 32'h42911bd7, 32'h0, 32'h42983f23};
test_input[2192:2199] = '{32'hc203d71b, 32'h401f10d4, 32'hc0964553, 32'h40ce5dbc, 32'hc26bd4b5, 32'h42082fe1, 32'hc28b979d, 32'h42b6d756};
test_output[2192:2199] = '{32'h0, 32'h401f10d4, 32'h0, 32'h40ce5dbc, 32'h0, 32'h42082fe1, 32'h0, 32'h42b6d756};
test_input[2200:2207] = '{32'hc16e2a15, 32'h417b21cf, 32'hc1e2a7f2, 32'h407a2bca, 32'h41fad26e, 32'h40e9a8ac, 32'hc0fca0d5, 32'h4242042c};
test_output[2200:2207] = '{32'h0, 32'h417b21cf, 32'h0, 32'h407a2bca, 32'h41fad26e, 32'h40e9a8ac, 32'h0, 32'h4242042c};
test_input[2208:2215] = '{32'h428bbc2d, 32'hc25173c8, 32'h4215376e, 32'hc24bf4f4, 32'h3fe842a7, 32'hc2a6eb79, 32'h3fd2cf31, 32'h42ba6e79};
test_output[2208:2215] = '{32'h428bbc2d, 32'h0, 32'h4215376e, 32'h0, 32'h3fe842a7, 32'h0, 32'h3fd2cf31, 32'h42ba6e79};
test_input[2216:2223] = '{32'h42b0865d, 32'hc049c66a, 32'h42514c01, 32'h42add7ff, 32'hc1e61b51, 32'h420c9711, 32'h41e47dc4, 32'h4295811d};
test_output[2216:2223] = '{32'h42b0865d, 32'h0, 32'h42514c01, 32'h42add7ff, 32'h0, 32'h420c9711, 32'h41e47dc4, 32'h4295811d};
test_input[2224:2231] = '{32'hc24abe3f, 32'h42604ad9, 32'hc1f1adf0, 32'h41d3d1fc, 32'hc29649d7, 32'hc2385556, 32'hc23bfa0c, 32'hc1b6ea38};
test_output[2224:2231] = '{32'h0, 32'h42604ad9, 32'h0, 32'h41d3d1fc, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2232:2239] = '{32'hc2b56503, 32'h40a511c8, 32'h42a29118, 32'hc0fdbbae, 32'hc18e4dcb, 32'hc270d221, 32'hc2804267, 32'hc25f8267};
test_output[2232:2239] = '{32'h0, 32'h40a511c8, 32'h42a29118, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2240:2247] = '{32'h40983efe, 32'hc25cf803, 32'h42837933, 32'hc1783e88, 32'h428520e3, 32'h4041354f, 32'hc21f4812, 32'hc22a5318};
test_output[2240:2247] = '{32'h40983efe, 32'h0, 32'h42837933, 32'h0, 32'h428520e3, 32'h4041354f, 32'h0, 32'h0};
test_input[2248:2255] = '{32'hc1a03760, 32'h422524b6, 32'hc11f787f, 32'h42c7f5bb, 32'h421fca4f, 32'h41739ded, 32'h4213eac4, 32'h419bf27d};
test_output[2248:2255] = '{32'h0, 32'h422524b6, 32'h0, 32'h42c7f5bb, 32'h421fca4f, 32'h41739ded, 32'h4213eac4, 32'h419bf27d};
test_input[2256:2263] = '{32'hc1b43022, 32'hc1b946f6, 32'h4249691d, 32'h416ae6e2, 32'h428c49fa, 32'hc1e56c1d, 32'hc2160625, 32'hc1d378b0};
test_output[2256:2263] = '{32'h0, 32'h0, 32'h4249691d, 32'h416ae6e2, 32'h428c49fa, 32'h0, 32'h0, 32'h0};
test_input[2264:2271] = '{32'h40b226c1, 32'h426ac450, 32'h42594ddd, 32'h429154b4, 32'h42a27769, 32'h428d7c6a, 32'h41b65f6f, 32'h421e1e5c};
test_output[2264:2271] = '{32'h40b226c1, 32'h426ac450, 32'h42594ddd, 32'h429154b4, 32'h42a27769, 32'h428d7c6a, 32'h41b65f6f, 32'h421e1e5c};
test_input[2272:2279] = '{32'hc248f8d9, 32'hc1d3654b, 32'h42606eb8, 32'h415c1260, 32'h425ea331, 32'hc20eefd3, 32'hc18ab0bb, 32'hc0af993f};
test_output[2272:2279] = '{32'h0, 32'h0, 32'h42606eb8, 32'h415c1260, 32'h425ea331, 32'h0, 32'h0, 32'h0};
test_input[2280:2287] = '{32'h428193b8, 32'h42b29ec0, 32'h42b22f8f, 32'hc1b13751, 32'h42b95091, 32'hc1be6492, 32'hc1ed19c7, 32'hc2318801};
test_output[2280:2287] = '{32'h428193b8, 32'h42b29ec0, 32'h42b22f8f, 32'h0, 32'h42b95091, 32'h0, 32'h0, 32'h0};
test_input[2288:2295] = '{32'hc28f3c9b, 32'h429e5f6b, 32'hc28db4a3, 32'h423d0cf6, 32'h423b4cb9, 32'hc1f26dbb, 32'h42569ab7, 32'h42b167ac};
test_output[2288:2295] = '{32'h0, 32'h429e5f6b, 32'h0, 32'h423d0cf6, 32'h423b4cb9, 32'h0, 32'h42569ab7, 32'h42b167ac};
test_input[2296:2303] = '{32'hc268cd37, 32'h418481c6, 32'hc2c04496, 32'hc28a7e25, 32'hc2685ef2, 32'h409c9c8b, 32'h418f2458, 32'h42b02c4c};
test_output[2296:2303] = '{32'h0, 32'h418481c6, 32'h0, 32'h0, 32'h0, 32'h409c9c8b, 32'h418f2458, 32'h42b02c4c};
test_input[2304:2311] = '{32'hc0b5ecd1, 32'h419e934f, 32'hc1897513, 32'hc246c5d0, 32'hc2c6006c, 32'hc262f913, 32'h4280cb76, 32'h428f4946};
test_output[2304:2311] = '{32'h0, 32'h419e934f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4280cb76, 32'h428f4946};
test_input[2312:2319] = '{32'h42bbdf6d, 32'hc2ae826c, 32'h42981970, 32'h42ad3146, 32'hc26b21e8, 32'h41f16170, 32'h40640a50, 32'hc217fefe};
test_output[2312:2319] = '{32'h42bbdf6d, 32'h0, 32'h42981970, 32'h42ad3146, 32'h0, 32'h41f16170, 32'h40640a50, 32'h0};
test_input[2320:2327] = '{32'hc2bc1286, 32'h4254bf07, 32'h42b2e784, 32'h4299551b, 32'hc281c707, 32'h42c6aaf4, 32'hc05b8169, 32'h4241d791};
test_output[2320:2327] = '{32'h0, 32'h4254bf07, 32'h42b2e784, 32'h4299551b, 32'h0, 32'h42c6aaf4, 32'h0, 32'h4241d791};
test_input[2328:2335] = '{32'h42936581, 32'hc2a05a8b, 32'h42440513, 32'hc21d4604, 32'hc0af3bb7, 32'hc27d5331, 32'hc2b8f76c, 32'h3fc12422};
test_output[2328:2335] = '{32'h42936581, 32'h0, 32'h42440513, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3fc12422};
test_input[2336:2343] = '{32'hc1099347, 32'hc0ce2666, 32'hc19f9f06, 32'h4263bd36, 32'h421e1df1, 32'hc2409573, 32'hc2ab58ff, 32'hc28b8a7b};
test_output[2336:2343] = '{32'h0, 32'h0, 32'h0, 32'h4263bd36, 32'h421e1df1, 32'h0, 32'h0, 32'h0};
test_input[2344:2351] = '{32'h42bd468a, 32'h42c61db8, 32'h428ee279, 32'h429ac50d, 32'hc295d10e, 32'h421958fa, 32'hc2a7238f, 32'hc269ac02};
test_output[2344:2351] = '{32'h42bd468a, 32'h42c61db8, 32'h428ee279, 32'h429ac50d, 32'h0, 32'h421958fa, 32'h0, 32'h0};
test_input[2352:2359] = '{32'h406aa3aa, 32'h42a0e4b5, 32'hc1001cb0, 32'h421a13a0, 32'hc2082dcc, 32'h4202959d, 32'hc12f7250, 32'hc0a6711e};
test_output[2352:2359] = '{32'h406aa3aa, 32'h42a0e4b5, 32'h0, 32'h421a13a0, 32'h0, 32'h4202959d, 32'h0, 32'h0};
test_input[2360:2367] = '{32'hc240c7b4, 32'h41a04361, 32'hc104427f, 32'h429daa39, 32'hc2979353, 32'h41e5505b, 32'hc25cb068, 32'h429723a7};
test_output[2360:2367] = '{32'h0, 32'h41a04361, 32'h0, 32'h429daa39, 32'h0, 32'h41e5505b, 32'h0, 32'h429723a7};
test_input[2368:2375] = '{32'h423d6294, 32'h42784a45, 32'hc27c68eb, 32'hc2024443, 32'hc2465142, 32'hc2c31eac, 32'hc2b3fb2d, 32'hc25f3d99};
test_output[2368:2375] = '{32'h423d6294, 32'h42784a45, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2376:2383] = '{32'hc1e449a7, 32'h428112bc, 32'hc17c7d83, 32'h42a4b695, 32'h4238ab13, 32'hc247c384, 32'hc1fdf4a9, 32'h42bcca14};
test_output[2376:2383] = '{32'h0, 32'h428112bc, 32'h0, 32'h42a4b695, 32'h4238ab13, 32'h0, 32'h0, 32'h42bcca14};
test_input[2384:2391] = '{32'hc22cf368, 32'hc2238a6b, 32'hc2a56a1c, 32'h422f84cb, 32'hc118bccc, 32'hc29b9ef3, 32'h4226742b, 32'hc29eb0f9};
test_output[2384:2391] = '{32'h0, 32'h0, 32'h0, 32'h422f84cb, 32'h0, 32'h0, 32'h4226742b, 32'h0};
test_input[2392:2399] = '{32'h41b625e7, 32'hc24691d1, 32'hc24af1af, 32'h41283248, 32'h41e348c1, 32'hc1a6e202, 32'h42c105d3, 32'h4257b1f1};
test_output[2392:2399] = '{32'h41b625e7, 32'h0, 32'h0, 32'h41283248, 32'h41e348c1, 32'h0, 32'h42c105d3, 32'h4257b1f1};
test_input[2400:2407] = '{32'h424cbdea, 32'h421749a2, 32'hc266b35d, 32'hc2944cc0, 32'h4294d351, 32'h40ec5feb, 32'h4260751c, 32'hc2adfddd};
test_output[2400:2407] = '{32'h424cbdea, 32'h421749a2, 32'h0, 32'h0, 32'h4294d351, 32'h40ec5feb, 32'h4260751c, 32'h0};
test_input[2408:2415] = '{32'h422ec316, 32'hc2bc2851, 32'hc2980917, 32'h42b2032f, 32'hc16e1d45, 32'h42547ed0, 32'h41c187bf, 32'hc2a0af95};
test_output[2408:2415] = '{32'h422ec316, 32'h0, 32'h0, 32'h42b2032f, 32'h0, 32'h42547ed0, 32'h41c187bf, 32'h0};
test_input[2416:2423] = '{32'hc0860751, 32'hc27fd169, 32'hc056a52e, 32'hc2979bc6, 32'hc2828844, 32'h42250da6, 32'hc1b4d855, 32'h415f09b6};
test_output[2416:2423] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42250da6, 32'h0, 32'h415f09b6};
test_input[2424:2431] = '{32'hc2b00d87, 32'h42c722bb, 32'hc2c24232, 32'h3f45fee1, 32'hc1a43bf4, 32'hc156dee3, 32'hc2a52c1d, 32'h42887798};
test_output[2424:2431] = '{32'h0, 32'h42c722bb, 32'h0, 32'h3f45fee1, 32'h0, 32'h0, 32'h0, 32'h42887798};
test_input[2432:2439] = '{32'h424ec307, 32'hc1d9fd0b, 32'hc0f925b7, 32'h4299e80b, 32'h42b61332, 32'hc2a414bb, 32'h421a1efd, 32'hc1639891};
test_output[2432:2439] = '{32'h424ec307, 32'h0, 32'h0, 32'h4299e80b, 32'h42b61332, 32'h0, 32'h421a1efd, 32'h0};
test_input[2440:2447] = '{32'h42a6929f, 32'hc0233dbe, 32'hc22ef853, 32'h429253a2, 32'h40edff6f, 32'h422a757b, 32'h428d3ba7, 32'hc2735c4e};
test_output[2440:2447] = '{32'h42a6929f, 32'h0, 32'h0, 32'h429253a2, 32'h40edff6f, 32'h422a757b, 32'h428d3ba7, 32'h0};
test_input[2448:2455] = '{32'hc29ac9e5, 32'h425f5bcf, 32'hc22ebf21, 32'hc21b49c8, 32'hc2be2df4, 32'hc28af242, 32'h42c5ea68, 32'h428e4a99};
test_output[2448:2455] = '{32'h0, 32'h425f5bcf, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c5ea68, 32'h428e4a99};
test_input[2456:2463] = '{32'h4237f628, 32'h423a3253, 32'hc2a956f5, 32'h420bb194, 32'hc2a74714, 32'h41f5dfa8, 32'hc285a20c, 32'h41b468f1};
test_output[2456:2463] = '{32'h4237f628, 32'h423a3253, 32'h0, 32'h420bb194, 32'h0, 32'h41f5dfa8, 32'h0, 32'h41b468f1};
test_input[2464:2471] = '{32'h429db47e, 32'h41001a30, 32'h40f80da7, 32'hc29e73c9, 32'h40e4068c, 32'h42bb8ca0, 32'h41256ee2, 32'hc20c3b6d};
test_output[2464:2471] = '{32'h429db47e, 32'h41001a30, 32'h40f80da7, 32'h0, 32'h40e4068c, 32'h42bb8ca0, 32'h41256ee2, 32'h0};
test_input[2472:2479] = '{32'hc292a1d8, 32'h42854216, 32'hc2bc5a2e, 32'h4285a745, 32'hc125ec46, 32'hc2bc5252, 32'h421b84fe, 32'hc293e3b8};
test_output[2472:2479] = '{32'h0, 32'h42854216, 32'h0, 32'h4285a745, 32'h0, 32'h0, 32'h421b84fe, 32'h0};
test_input[2480:2487] = '{32'h4267f2f2, 32'h42a85f10, 32'h425622bd, 32'hc2946a0f, 32'h42ba5269, 32'hc2bab949, 32'h40c0ca97, 32'h41e73b06};
test_output[2480:2487] = '{32'h4267f2f2, 32'h42a85f10, 32'h425622bd, 32'h0, 32'h42ba5269, 32'h0, 32'h40c0ca97, 32'h41e73b06};
test_input[2488:2495] = '{32'hc28715ba, 32'h4291ccf0, 32'h42338690, 32'hc2b1171e, 32'hc1aebc04, 32'hc29ed509, 32'h427a987a, 32'h41d4f1fc};
test_output[2488:2495] = '{32'h0, 32'h4291ccf0, 32'h42338690, 32'h0, 32'h0, 32'h0, 32'h427a987a, 32'h41d4f1fc};
test_input[2496:2503] = '{32'hc28527ac, 32'h418eea55, 32'hc260e8c5, 32'h4155b743, 32'hc2207f53, 32'h3ffd8092, 32'hc25aeedb, 32'hc17b1c94};
test_output[2496:2503] = '{32'h0, 32'h418eea55, 32'h0, 32'h4155b743, 32'h0, 32'h3ffd8092, 32'h0, 32'h0};
test_input[2504:2511] = '{32'hc29e492f, 32'h42770382, 32'h4103adb8, 32'hc1d15f4f, 32'h425f1972, 32'h3fb2ab7c, 32'h420f7063, 32'hc2b1a62d};
test_output[2504:2511] = '{32'h0, 32'h42770382, 32'h4103adb8, 32'h0, 32'h425f1972, 32'h3fb2ab7c, 32'h420f7063, 32'h0};
test_input[2512:2519] = '{32'h41d02345, 32'hc23eeb62, 32'h42183e8f, 32'hc2a6bea7, 32'h42a10b8b, 32'hc24dab9a, 32'hc08bf56f, 32'hc215123d};
test_output[2512:2519] = '{32'h41d02345, 32'h0, 32'h42183e8f, 32'h0, 32'h42a10b8b, 32'h0, 32'h0, 32'h0};
test_input[2520:2527] = '{32'hc19296b0, 32'h4251b843, 32'h42106757, 32'h42c2489f, 32'hc190917c, 32'hc0dc9b46, 32'h42aa1f46, 32'hc24250bb};
test_output[2520:2527] = '{32'h0, 32'h4251b843, 32'h42106757, 32'h42c2489f, 32'h0, 32'h0, 32'h42aa1f46, 32'h0};
test_input[2528:2535] = '{32'h428eedff, 32'hc2ad860d, 32'hbf563cdb, 32'h3e80cb78, 32'hc20c9298, 32'h4190c332, 32'h42024208, 32'hc2bdbdec};
test_output[2528:2535] = '{32'h428eedff, 32'h0, 32'h0, 32'h3e80cb78, 32'h0, 32'h4190c332, 32'h42024208, 32'h0};
test_input[2536:2543] = '{32'h42550ade, 32'h4112d491, 32'h42509e90, 32'hc2c55fe7, 32'hc05b8e09, 32'hc025a033, 32'h4253de42, 32'h412fbbdb};
test_output[2536:2543] = '{32'h42550ade, 32'h4112d491, 32'h42509e90, 32'h0, 32'h0, 32'h0, 32'h4253de42, 32'h412fbbdb};
test_input[2544:2551] = '{32'h41d685bc, 32'h42b9e44d, 32'h4234983b, 32'h42045e88, 32'h42ac274c, 32'h411ba787, 32'hc27112e0, 32'hc25e670a};
test_output[2544:2551] = '{32'h41d685bc, 32'h42b9e44d, 32'h4234983b, 32'h42045e88, 32'h42ac274c, 32'h411ba787, 32'h0, 32'h0};
test_input[2552:2559] = '{32'hc22b35d9, 32'h418d134c, 32'h42c6a14e, 32'hc28599d2, 32'hc2be306f, 32'h4285cffc, 32'hc28e7b33, 32'h421622e6};
test_output[2552:2559] = '{32'h0, 32'h418d134c, 32'h42c6a14e, 32'h0, 32'h0, 32'h4285cffc, 32'h0, 32'h421622e6};
test_input[2560:2567] = '{32'hc1222158, 32'h4206c665, 32'h429c8748, 32'hc21ab2e1, 32'h421a5eba, 32'h42990397, 32'hc2b29b39, 32'hc29ab705};
test_output[2560:2567] = '{32'h0, 32'h4206c665, 32'h429c8748, 32'h0, 32'h421a5eba, 32'h42990397, 32'h0, 32'h0};
test_input[2568:2575] = '{32'h426f59f7, 32'h40bbdd82, 32'h42be7462, 32'h3fca4c5b, 32'h42a597d5, 32'hc249ca7d, 32'hc1a90923, 32'hc22a89c9};
test_output[2568:2575] = '{32'h426f59f7, 32'h40bbdd82, 32'h42be7462, 32'h3fca4c5b, 32'h42a597d5, 32'h0, 32'h0, 32'h0};
test_input[2576:2583] = '{32'hc2b79e44, 32'h4256d4bc, 32'hc2bd3ff8, 32'h4206113c, 32'h410e5f70, 32'hc2b49640, 32'hc19d0ac7, 32'hc2225ee1};
test_output[2576:2583] = '{32'h0, 32'h4256d4bc, 32'h0, 32'h4206113c, 32'h410e5f70, 32'h0, 32'h0, 32'h0};
test_input[2584:2591] = '{32'hc2a09501, 32'h42c75484, 32'hc25497bf, 32'h407e0695, 32'hc25c7b35, 32'h423673bd, 32'h422ebbd7, 32'hc2114265};
test_output[2584:2591] = '{32'h0, 32'h42c75484, 32'h0, 32'h407e0695, 32'h0, 32'h423673bd, 32'h422ebbd7, 32'h0};
test_input[2592:2599] = '{32'h412caa88, 32'hc2c0525a, 32'hc1ac1a9d, 32'hc28e36cc, 32'h42928fde, 32'h4201ce54, 32'h4253c5b8, 32'h421d7980};
test_output[2592:2599] = '{32'h412caa88, 32'h0, 32'h0, 32'h0, 32'h42928fde, 32'h4201ce54, 32'h4253c5b8, 32'h421d7980};
test_input[2600:2607] = '{32'h425a4e9a, 32'hc21134e2, 32'hc2a2fd97, 32'hc0c4a225, 32'h40a175e4, 32'hc24398e0, 32'hc256c386, 32'hc20764dc};
test_output[2600:2607] = '{32'h425a4e9a, 32'h0, 32'h0, 32'h0, 32'h40a175e4, 32'h0, 32'h0, 32'h0};
test_input[2608:2615] = '{32'h422bbe38, 32'h42011522, 32'hc2807028, 32'h42a305c8, 32'hc2724e3b, 32'h411e0178, 32'hc209ac05, 32'h416fb439};
test_output[2608:2615] = '{32'h422bbe38, 32'h42011522, 32'h0, 32'h42a305c8, 32'h0, 32'h411e0178, 32'h0, 32'h416fb439};
test_input[2616:2623] = '{32'h421dcbca, 32'h42921319, 32'hc1f72800, 32'hc2077989, 32'h420d832f, 32'hc2555688, 32'h41d16471, 32'h41bdac11};
test_output[2616:2623] = '{32'h421dcbca, 32'h42921319, 32'h0, 32'h0, 32'h420d832f, 32'h0, 32'h41d16471, 32'h41bdac11};
test_input[2624:2631] = '{32'h4121cc34, 32'hc27f9d2c, 32'hc270f17e, 32'hc2a210e5, 32'h4272f5de, 32'h42bf2e57, 32'hc2b87096, 32'h422a8abc};
test_output[2624:2631] = '{32'h4121cc34, 32'h0, 32'h0, 32'h0, 32'h4272f5de, 32'h42bf2e57, 32'h0, 32'h422a8abc};
test_input[2632:2639] = '{32'hc20b0417, 32'hc281da74, 32'h428de2db, 32'hc2846ef5, 32'hc1f62b27, 32'h42aaf960, 32'hc28c2b14, 32'h421d9693};
test_output[2632:2639] = '{32'h0, 32'h0, 32'h428de2db, 32'h0, 32'h0, 32'h42aaf960, 32'h0, 32'h421d9693};
test_input[2640:2647] = '{32'hc26f3414, 32'h42a43c52, 32'hc207caf0, 32'h42140e0b, 32'h4282bd90, 32'h412655a6, 32'hc28b10d4, 32'hc2c0565c};
test_output[2640:2647] = '{32'h0, 32'h42a43c52, 32'h0, 32'h42140e0b, 32'h4282bd90, 32'h412655a6, 32'h0, 32'h0};
test_input[2648:2655] = '{32'h426fc956, 32'h3fbee2a2, 32'hbf5c938c, 32'hc149c1df, 32'hc2adf6b2, 32'h41997e65, 32'h4291b865, 32'h426d6aeb};
test_output[2648:2655] = '{32'h426fc956, 32'h3fbee2a2, 32'h0, 32'h0, 32'h0, 32'h41997e65, 32'h4291b865, 32'h426d6aeb};
test_input[2656:2663] = '{32'h424b971b, 32'h422d0878, 32'h41c0f0f8, 32'h41f196bf, 32'h42c46a28, 32'h4282ae45, 32'h414fcc5f, 32'h42560c79};
test_output[2656:2663] = '{32'h424b971b, 32'h422d0878, 32'h41c0f0f8, 32'h41f196bf, 32'h42c46a28, 32'h4282ae45, 32'h414fcc5f, 32'h42560c79};
test_input[2664:2671] = '{32'h4246c745, 32'h423ae563, 32'h41dfd0b5, 32'h4265df85, 32'h40c46bb0, 32'h4286ea3c, 32'h420d49a8, 32'hc14e7b10};
test_output[2664:2671] = '{32'h4246c745, 32'h423ae563, 32'h41dfd0b5, 32'h4265df85, 32'h40c46bb0, 32'h4286ea3c, 32'h420d49a8, 32'h0};
test_input[2672:2679] = '{32'h419ef47b, 32'hc0be14af, 32'hc12425d0, 32'hc1a6b484, 32'hc296b46c, 32'hc2a59e0f, 32'hc18d6f05, 32'h429a5b92};
test_output[2672:2679] = '{32'h419ef47b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429a5b92};
test_input[2680:2687] = '{32'h41b4a04e, 32'hc284d024, 32'hc293a882, 32'h419b12a2, 32'hc297315f, 32'h400676c3, 32'h423f1455, 32'hc2b81cdd};
test_output[2680:2687] = '{32'h41b4a04e, 32'h0, 32'h0, 32'h419b12a2, 32'h0, 32'h400676c3, 32'h423f1455, 32'h0};
test_input[2688:2695] = '{32'hc0cbf423, 32'hc1be4dc9, 32'hc1ede5bc, 32'hc2160b4a, 32'hc293ae4e, 32'h412624ac, 32'h4289834d, 32'hc13c83a6};
test_output[2688:2695] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h412624ac, 32'h4289834d, 32'h0};
test_input[2696:2703] = '{32'hc299a457, 32'hc03f7c5d, 32'h3e183a38, 32'hc164882a, 32'hc22b01a3, 32'h42a78e2a, 32'hc25042ce, 32'hc1dc28fd};
test_output[2696:2703] = '{32'h0, 32'h0, 32'h3e183a38, 32'h0, 32'h0, 32'h42a78e2a, 32'h0, 32'h0};
test_input[2704:2711] = '{32'h429c19ee, 32'hc0ac1a86, 32'h4264ce93, 32'hc291b787, 32'h42b7352c, 32'hc23338bf, 32'hc0a48f04, 32'hc2b987ac};
test_output[2704:2711] = '{32'h429c19ee, 32'h0, 32'h4264ce93, 32'h0, 32'h42b7352c, 32'h0, 32'h0, 32'h0};
test_input[2712:2719] = '{32'h420971c4, 32'hc21a281f, 32'h417154ab, 32'h414e504a, 32'h3f19c9fe, 32'h4291d105, 32'hc2abd23a, 32'h428db1c4};
test_output[2712:2719] = '{32'h420971c4, 32'h0, 32'h417154ab, 32'h414e504a, 32'h3f19c9fe, 32'h4291d105, 32'h0, 32'h428db1c4};
test_input[2720:2727] = '{32'h41fd1859, 32'h42a92486, 32'h425c5016, 32'h4293fad8, 32'h4039c347, 32'hc2c251f5, 32'hc23eb9f5, 32'h4298ed43};
test_output[2720:2727] = '{32'h41fd1859, 32'h42a92486, 32'h425c5016, 32'h4293fad8, 32'h4039c347, 32'h0, 32'h0, 32'h4298ed43};
test_input[2728:2735] = '{32'hc299d644, 32'hc2919955, 32'h41a97a46, 32'h42a371fb, 32'h423ca7fe, 32'hc1df0dff, 32'hc29dc0fd, 32'h42b656f8};
test_output[2728:2735] = '{32'h0, 32'h0, 32'h41a97a46, 32'h42a371fb, 32'h423ca7fe, 32'h0, 32'h0, 32'h42b656f8};
test_input[2736:2743] = '{32'hc2c51b21, 32'h4229d6bc, 32'hc1b03387, 32'hc2858b48, 32'hc28c7202, 32'hc2b36e71, 32'h4108bd96, 32'h404f73b9};
test_output[2736:2743] = '{32'h0, 32'h4229d6bc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4108bd96, 32'h404f73b9};
test_input[2744:2751] = '{32'hc1e21da9, 32'h41eb8a6d, 32'h42b3eba1, 32'hc2b7c461, 32'h4222d7d8, 32'hc2b1bd23, 32'hc27ed2c0, 32'hc2b5f402};
test_output[2744:2751] = '{32'h0, 32'h41eb8a6d, 32'h42b3eba1, 32'h0, 32'h4222d7d8, 32'h0, 32'h0, 32'h0};
test_input[2752:2759] = '{32'hbe2e8427, 32'hc22bf553, 32'h42317cee, 32'h4264159c, 32'h41e9733c, 32'h4274297f, 32'h4242efeb, 32'h42984e14};
test_output[2752:2759] = '{32'h0, 32'h0, 32'h42317cee, 32'h4264159c, 32'h41e9733c, 32'h4274297f, 32'h4242efeb, 32'h42984e14};
test_input[2760:2767] = '{32'h3e8c8ae9, 32'h42b127e2, 32'hc254162c, 32'hc1d50051, 32'h420cbe1b, 32'hc216c853, 32'hc204b7d8, 32'hc108d3b8};
test_output[2760:2767] = '{32'h3e8c8ae9, 32'h42b127e2, 32'h0, 32'h0, 32'h420cbe1b, 32'h0, 32'h0, 32'h0};
test_input[2768:2775] = '{32'h42a281d0, 32'h4228920e, 32'h405c85e4, 32'h4208da6a, 32'hc2098f70, 32'hc14480bd, 32'hc2547c94, 32'hc289f017};
test_output[2768:2775] = '{32'h42a281d0, 32'h4228920e, 32'h405c85e4, 32'h4208da6a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2776:2783] = '{32'h42b47290, 32'hc288170a, 32'h4252dea4, 32'hc227590c, 32'h425677fb, 32'hc2a69c00, 32'h41c74ef1, 32'h42ae6c22};
test_output[2776:2783] = '{32'h42b47290, 32'h0, 32'h4252dea4, 32'h0, 32'h425677fb, 32'h0, 32'h41c74ef1, 32'h42ae6c22};
test_input[2784:2791] = '{32'hc288ae9c, 32'hc266be80, 32'hc2c4d004, 32'h405f14cb, 32'hc233e466, 32'h425e7e91, 32'h42a36f0f, 32'h4222eecb};
test_output[2784:2791] = '{32'h0, 32'h0, 32'h0, 32'h405f14cb, 32'h0, 32'h425e7e91, 32'h42a36f0f, 32'h4222eecb};
test_input[2792:2799] = '{32'h42b4c70f, 32'h4268ddbc, 32'hc26bf237, 32'h41ca016b, 32'hc2361e99, 32'hc1dfc364, 32'hc135ac1a, 32'hc231faf4};
test_output[2792:2799] = '{32'h42b4c70f, 32'h4268ddbc, 32'h0, 32'h41ca016b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2800:2807] = '{32'h428089a3, 32'h42045a79, 32'h42b5863e, 32'hc2b37d6a, 32'hc19c1198, 32'h42518c8a, 32'hc19bbf29, 32'hc2b8c78c};
test_output[2800:2807] = '{32'h428089a3, 32'h42045a79, 32'h42b5863e, 32'h0, 32'h0, 32'h42518c8a, 32'h0, 32'h0};
test_input[2808:2815] = '{32'hc2c0f709, 32'hc2a279a6, 32'hc29f23d5, 32'h420e0e88, 32'h412d29a6, 32'hc2c3df54, 32'h41e203c9, 32'h41a345cd};
test_output[2808:2815] = '{32'h0, 32'h0, 32'h0, 32'h420e0e88, 32'h412d29a6, 32'h0, 32'h41e203c9, 32'h41a345cd};
test_input[2816:2823] = '{32'h408971f5, 32'h4265bc3f, 32'hc0849598, 32'hc2b3dafb, 32'h425918f6, 32'h422541ef, 32'h42c1817f, 32'hbf8e5a24};
test_output[2816:2823] = '{32'h408971f5, 32'h4265bc3f, 32'h0, 32'h0, 32'h425918f6, 32'h422541ef, 32'h42c1817f, 32'h0};
test_input[2824:2831] = '{32'hc217d499, 32'h41d3e523, 32'h411bc4ad, 32'h42b0cc4d, 32'hc07c23e4, 32'hc22f134f, 32'h427bfb9a, 32'hc24bbe2f};
test_output[2824:2831] = '{32'h0, 32'h41d3e523, 32'h411bc4ad, 32'h42b0cc4d, 32'h0, 32'h0, 32'h427bfb9a, 32'h0};
test_input[2832:2839] = '{32'hc18af98c, 32'hc090c0ad, 32'hc266f9b6, 32'hc28d3e61, 32'h422fe605, 32'h42a8f7cf, 32'h41d52d57, 32'h42248883};
test_output[2832:2839] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h422fe605, 32'h42a8f7cf, 32'h41d52d57, 32'h42248883};
test_input[2840:2847] = '{32'hc1bc1660, 32'hc2c1c486, 32'h42356cbe, 32'h40b1f01d, 32'h41dfe755, 32'hc1de8178, 32'hc2a3382e, 32'h3f4fc45f};
test_output[2840:2847] = '{32'h0, 32'h0, 32'h42356cbe, 32'h40b1f01d, 32'h41dfe755, 32'h0, 32'h0, 32'h3f4fc45f};
test_input[2848:2855] = '{32'hc2ad5e4f, 32'h40b97c50, 32'h42677114, 32'h42535ece, 32'h427082ef, 32'hc251166a, 32'h42aec070, 32'h407bc2c3};
test_output[2848:2855] = '{32'h0, 32'h40b97c50, 32'h42677114, 32'h42535ece, 32'h427082ef, 32'h0, 32'h42aec070, 32'h407bc2c3};
test_input[2856:2863] = '{32'h417928fd, 32'hc2b62e91, 32'h426649da, 32'hc2b2ad39, 32'hc2c4cbc1, 32'hc19822e9, 32'h4216fb73, 32'hc2b6402d};
test_output[2856:2863] = '{32'h417928fd, 32'h0, 32'h426649da, 32'h0, 32'h0, 32'h0, 32'h4216fb73, 32'h0};
test_input[2864:2871] = '{32'hc2aebd92, 32'hc23daa38, 32'hc2be164f, 32'hc298a92a, 32'h41b85eea, 32'hc24e48ec, 32'hc2429441, 32'hc2b37546};
test_output[2864:2871] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41b85eea, 32'h0, 32'h0, 32'h0};
test_input[2872:2879] = '{32'hc2c6f38b, 32'hc13e6ebf, 32'h4245d0af, 32'hc28fa5fb, 32'hc2407dd2, 32'h42bb5c27, 32'hc1282aaf, 32'h42924db9};
test_output[2872:2879] = '{32'h0, 32'h0, 32'h4245d0af, 32'h0, 32'h0, 32'h42bb5c27, 32'h0, 32'h42924db9};
test_input[2880:2887] = '{32'h4084bec6, 32'hc11c5e45, 32'h4278ba27, 32'h42938faf, 32'h42c28b1b, 32'hc1a0e2d7, 32'hc24f2003, 32'h41334d60};
test_output[2880:2887] = '{32'h4084bec6, 32'h0, 32'h4278ba27, 32'h42938faf, 32'h42c28b1b, 32'h0, 32'h0, 32'h41334d60};
test_input[2888:2895] = '{32'h4217314e, 32'hc2b1b3e0, 32'h42a79465, 32'h422fc998, 32'h42782ec1, 32'h415fe6cf, 32'hc26d654b, 32'hc0bf44f0};
test_output[2888:2895] = '{32'h4217314e, 32'h0, 32'h42a79465, 32'h422fc998, 32'h42782ec1, 32'h415fe6cf, 32'h0, 32'h0};
test_input[2896:2903] = '{32'hc28eabbe, 32'hc279074f, 32'h4297334d, 32'h422ef793, 32'hc092508f, 32'h4226ee06, 32'hc19b3993, 32'h410993d4};
test_output[2896:2903] = '{32'h0, 32'h0, 32'h4297334d, 32'h422ef793, 32'h0, 32'h4226ee06, 32'h0, 32'h410993d4};
test_input[2904:2911] = '{32'h41eae4da, 32'h41ddc813, 32'hc106bfcd, 32'hc28ef742, 32'h42667a42, 32'h420d8c4d, 32'h42c077be, 32'hc2afc2e7};
test_output[2904:2911] = '{32'h41eae4da, 32'h41ddc813, 32'h0, 32'h0, 32'h42667a42, 32'h420d8c4d, 32'h42c077be, 32'h0};
test_input[2912:2919] = '{32'hc2708efd, 32'hc29a5571, 32'hc1ff1ac5, 32'h41631cc4, 32'h417741e6, 32'hc2be17c7, 32'hbf919d3c, 32'h402f46ce};
test_output[2912:2919] = '{32'h0, 32'h0, 32'h0, 32'h41631cc4, 32'h417741e6, 32'h0, 32'h0, 32'h402f46ce};
test_input[2920:2927] = '{32'h423cc472, 32'h42a4da98, 32'hc298e778, 32'h41e9b877, 32'h4236ff21, 32'hc25aaf95, 32'hc29c5dba, 32'h425a8b3e};
test_output[2920:2927] = '{32'h423cc472, 32'h42a4da98, 32'h0, 32'h41e9b877, 32'h4236ff21, 32'h0, 32'h0, 32'h425a8b3e};
test_input[2928:2935] = '{32'h41c64802, 32'h425c1ef4, 32'hc210a4dc, 32'h41cb4038, 32'h41b71cac, 32'h42abfcde, 32'h421d3c86, 32'h41aa846a};
test_output[2928:2935] = '{32'h41c64802, 32'h425c1ef4, 32'h0, 32'h41cb4038, 32'h41b71cac, 32'h42abfcde, 32'h421d3c86, 32'h41aa846a};
test_input[2936:2943] = '{32'hc2980407, 32'hc25e05e6, 32'h41919090, 32'h428622db, 32'h42b2ca97, 32'hc2af0bbe, 32'h421dd722, 32'hc1977176};
test_output[2936:2943] = '{32'h0, 32'h0, 32'h41919090, 32'h428622db, 32'h42b2ca97, 32'h0, 32'h421dd722, 32'h0};
test_input[2944:2951] = '{32'hc13381d4, 32'h42bb9214, 32'hc20dc4fd, 32'h41b981ac, 32'h42242e3e, 32'hc1e61a80, 32'hc2233dc6, 32'h4273144d};
test_output[2944:2951] = '{32'h0, 32'h42bb9214, 32'h0, 32'h41b981ac, 32'h42242e3e, 32'h0, 32'h0, 32'h4273144d};
test_input[2952:2959] = '{32'hc2a8ef0d, 32'hc206ad17, 32'h42b633c4, 32'hc1ea7e50, 32'h423536dd, 32'hc2bf52b0, 32'hc2a00d27, 32'h42c19d9c};
test_output[2952:2959] = '{32'h0, 32'h0, 32'h42b633c4, 32'h0, 32'h423536dd, 32'h0, 32'h0, 32'h42c19d9c};
test_input[2960:2967] = '{32'hc29e197e, 32'h42aa4065, 32'hc27ef055, 32'h42714d12, 32'hc1ce3211, 32'h426bce2d, 32'hc2a5bcdb, 32'hc29a8685};
test_output[2960:2967] = '{32'h0, 32'h42aa4065, 32'h0, 32'h42714d12, 32'h0, 32'h426bce2d, 32'h0, 32'h0};
test_input[2968:2975] = '{32'hc1e6c331, 32'h42101c19, 32'hc2404cc7, 32'hc2829cfb, 32'h41ebca4d, 32'hc20cfc3c, 32'hc1fdb609, 32'hc21d5ca5};
test_output[2968:2975] = '{32'h0, 32'h42101c19, 32'h0, 32'h0, 32'h41ebca4d, 32'h0, 32'h0, 32'h0};
test_input[2976:2983] = '{32'h42bce599, 32'h424fa7a6, 32'hc2899aa9, 32'h42ac459f, 32'hbef8e118, 32'hc197751f, 32'h4239394a, 32'h42b7887c};
test_output[2976:2983] = '{32'h42bce599, 32'h424fa7a6, 32'h0, 32'h42ac459f, 32'h0, 32'h0, 32'h4239394a, 32'h42b7887c};
test_input[2984:2991] = '{32'h422e92ab, 32'h41c8d943, 32'h42952da1, 32'hc287b12b, 32'hc2858545, 32'hc2556a3a, 32'hc292661f, 32'h42baf6c3};
test_output[2984:2991] = '{32'h422e92ab, 32'h41c8d943, 32'h42952da1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42baf6c3};
test_input[2992:2999] = '{32'hc210dff3, 32'h42bb68ed, 32'hc28a14e0, 32'h42b79741, 32'h42b91023, 32'h41361d45, 32'h42420a80, 32'h41c04d72};
test_output[2992:2999] = '{32'h0, 32'h42bb68ed, 32'h0, 32'h42b79741, 32'h42b91023, 32'h41361d45, 32'h42420a80, 32'h41c04d72};
test_input[3000:3007] = '{32'h42adc9a8, 32'hc2c4fb23, 32'hc12694d4, 32'hc147fd3e, 32'h42bb453d, 32'h429f4e33, 32'h4208557c, 32'h4244deee};
test_output[3000:3007] = '{32'h42adc9a8, 32'h0, 32'h0, 32'h0, 32'h42bb453d, 32'h429f4e33, 32'h4208557c, 32'h4244deee};
test_input[3008:3015] = '{32'h4234436a, 32'h42809e2b, 32'hc247d2c8, 32'h422236bf, 32'h42c0258f, 32'hc141dde8, 32'hc292e8f1, 32'hc281271f};
test_output[3008:3015] = '{32'h4234436a, 32'h42809e2b, 32'h0, 32'h422236bf, 32'h42c0258f, 32'h0, 32'h0, 32'h0};
test_input[3016:3023] = '{32'hc24b0633, 32'hc0fb3912, 32'hc246bd9d, 32'hc257039a, 32'hc23cdf7c, 32'hc268b754, 32'h4191cd2b, 32'h419874e8};
test_output[3016:3023] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4191cd2b, 32'h419874e8};
test_input[3024:3031] = '{32'h42b3cf68, 32'h42abdece, 32'hc2c51ef7, 32'h4118c1bd, 32'h428a0d60, 32'hc2b99d55, 32'hc1683f5c, 32'h41f14212};
test_output[3024:3031] = '{32'h42b3cf68, 32'h42abdece, 32'h0, 32'h4118c1bd, 32'h428a0d60, 32'h0, 32'h0, 32'h41f14212};
test_input[3032:3039] = '{32'h40b93d0b, 32'h423821b9, 32'hc216bb60, 32'hc258c5b8, 32'hc2c32ae6, 32'hc2a8cef2, 32'hc2b7db4b, 32'hc29ec033};
test_output[3032:3039] = '{32'h40b93d0b, 32'h423821b9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3040:3047] = '{32'h41fba73e, 32'h4243b8be, 32'h426fa990, 32'h4277a5c8, 32'h41f56ba0, 32'h41b7dd19, 32'hc2b9853b, 32'h42bb0c8a};
test_output[3040:3047] = '{32'h41fba73e, 32'h4243b8be, 32'h426fa990, 32'h4277a5c8, 32'h41f56ba0, 32'h41b7dd19, 32'h0, 32'h42bb0c8a};
test_input[3048:3055] = '{32'hc2a283d4, 32'h42b28f6a, 32'hc2a5b9fb, 32'h429b855a, 32'h40d7dbca, 32'h428445f1, 32'hc28d0254, 32'hc2229479};
test_output[3048:3055] = '{32'h0, 32'h42b28f6a, 32'h0, 32'h429b855a, 32'h40d7dbca, 32'h428445f1, 32'h0, 32'h0};
test_input[3056:3063] = '{32'hc2940d7c, 32'hc15d8ff8, 32'hc223bef2, 32'hc2b61901, 32'h42440997, 32'h42b8768b, 32'h4245fc25, 32'hc2000d6e};
test_output[3056:3063] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42440997, 32'h42b8768b, 32'h4245fc25, 32'h0};
test_input[3064:3071] = '{32'hc09a13af, 32'hc1d5c2d1, 32'hc1aa1b20, 32'hc2369fa1, 32'h40d9f828, 32'h4230fee2, 32'hc2c02175, 32'hc210ecee};
test_output[3064:3071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40d9f828, 32'h4230fee2, 32'h0, 32'h0};
test_input[3072:3079] = '{32'hc21fa7ae, 32'h40f6335b, 32'hc0d3ed01, 32'h41aef386, 32'h42c7d5e7, 32'hc24d2b28, 32'hc2ac953d, 32'h41bde746};
test_output[3072:3079] = '{32'h0, 32'h40f6335b, 32'h0, 32'h41aef386, 32'h42c7d5e7, 32'h0, 32'h0, 32'h41bde746};
test_input[3080:3087] = '{32'hc0b8251e, 32'hc2979ab9, 32'h42245238, 32'hc285d308, 32'h41e2f2cd, 32'hc206dddd, 32'hc2bfdbb7, 32'hc23ba739};
test_output[3080:3087] = '{32'h0, 32'h0, 32'h42245238, 32'h0, 32'h41e2f2cd, 32'h0, 32'h0, 32'h0};
test_input[3088:3095] = '{32'h4261b127, 32'hc2925a5d, 32'h4157ea10, 32'hc2a7c0a7, 32'h42a0582a, 32'h41748d68, 32'h422a8c00, 32'h42b12444};
test_output[3088:3095] = '{32'h4261b127, 32'h0, 32'h4157ea10, 32'h0, 32'h42a0582a, 32'h41748d68, 32'h422a8c00, 32'h42b12444};
test_input[3096:3103] = '{32'hc2215d7f, 32'hc2af4f3c, 32'hc205b99f, 32'hc227f089, 32'hc2229e79, 32'hc285feea, 32'hc1535d2d, 32'h42a68411};
test_output[3096:3103] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a68411};
test_input[3104:3111] = '{32'hc2763636, 32'hc19699ef, 32'hc21806ce, 32'h423442dc, 32'hc10b3e0f, 32'hc2a90d95, 32'h423d9f9e, 32'h42b542e9};
test_output[3104:3111] = '{32'h0, 32'h0, 32'h0, 32'h423442dc, 32'h0, 32'h0, 32'h423d9f9e, 32'h42b542e9};
test_input[3112:3119] = '{32'h4239edc5, 32'hc09ee350, 32'hc1f186d9, 32'h424978b5, 32'hc1ad8865, 32'h42552e06, 32'h42a371d8, 32'h41f8ba7d};
test_output[3112:3119] = '{32'h4239edc5, 32'h0, 32'h0, 32'h424978b5, 32'h0, 32'h42552e06, 32'h42a371d8, 32'h41f8ba7d};
test_input[3120:3127] = '{32'h42c3199f, 32'hc28741c3, 32'h41deb785, 32'h426fed15, 32'h422c64fc, 32'hc22c2d51, 32'hc28e513b, 32'hc21f9f5e};
test_output[3120:3127] = '{32'h42c3199f, 32'h0, 32'h41deb785, 32'h426fed15, 32'h422c64fc, 32'h0, 32'h0, 32'h0};
test_input[3128:3135] = '{32'h41956689, 32'hc24f8cae, 32'hc27fbe7e, 32'h427f6e27, 32'h4180088b, 32'h4298fd5e, 32'hc20cf4d4, 32'h4247f5a5};
test_output[3128:3135] = '{32'h41956689, 32'h0, 32'h0, 32'h427f6e27, 32'h4180088b, 32'h4298fd5e, 32'h0, 32'h4247f5a5};
test_input[3136:3143] = '{32'hc2b6f254, 32'h411dca36, 32'hc206e0f9, 32'h42829dda, 32'h41f1dbce, 32'h427bc4c7, 32'h4286d167, 32'h428e0348};
test_output[3136:3143] = '{32'h0, 32'h411dca36, 32'h0, 32'h42829dda, 32'h41f1dbce, 32'h427bc4c7, 32'h4286d167, 32'h428e0348};
test_input[3144:3151] = '{32'hc2322f08, 32'hc2c52c69, 32'h41d797a6, 32'h420a2ff7, 32'hc1174eb8, 32'hc29ffc2a, 32'hc29a2c88, 32'h42644d12};
test_output[3144:3151] = '{32'h0, 32'h0, 32'h41d797a6, 32'h420a2ff7, 32'h0, 32'h0, 32'h0, 32'h42644d12};
test_input[3152:3159] = '{32'h428c7ef7, 32'hc29ac300, 32'h426e8b7c, 32'hc0acaecb, 32'h41166a83, 32'hc2895c8f, 32'h42c0609d, 32'hc06ceac5};
test_output[3152:3159] = '{32'h428c7ef7, 32'h0, 32'h426e8b7c, 32'h0, 32'h41166a83, 32'h0, 32'h42c0609d, 32'h0};
test_input[3160:3167] = '{32'h42ac036e, 32'h42a7a164, 32'hc13a58d8, 32'hc248529c, 32'hc298e25b, 32'hc2a55c7e, 32'hc295b1e2, 32'hc2b52a94};
test_output[3160:3167] = '{32'h42ac036e, 32'h42a7a164, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3168:3175] = '{32'hc10d60ae, 32'hbe358191, 32'h42a93bb0, 32'hc2b4618e, 32'hc2435633, 32'hc2034d90, 32'hc1a57254, 32'h420bd30d};
test_output[3168:3175] = '{32'h0, 32'h0, 32'h42a93bb0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420bd30d};
test_input[3176:3183] = '{32'hc29b9244, 32'hc1f882e6, 32'h4271b10d, 32'hc27072df, 32'h42afa0bd, 32'h42039ffe, 32'hc24740d3, 32'hc207fd14};
test_output[3176:3183] = '{32'h0, 32'h0, 32'h4271b10d, 32'h0, 32'h42afa0bd, 32'h42039ffe, 32'h0, 32'h0};
test_input[3184:3191] = '{32'hc2008ad6, 32'h42ab9045, 32'hc29d0321, 32'hc2acacef, 32'h429e55f0, 32'hc29444be, 32'hc20e1b29, 32'hc227d618};
test_output[3184:3191] = '{32'h0, 32'h42ab9045, 32'h0, 32'h0, 32'h429e55f0, 32'h0, 32'h0, 32'h0};
test_input[3192:3199] = '{32'hc10c81e7, 32'h42af1cd7, 32'h42becbd2, 32'hc276e877, 32'hc1d4f033, 32'hc137cfb8, 32'h42a267f0, 32'hc1a75100};
test_output[3192:3199] = '{32'h0, 32'h42af1cd7, 32'h42becbd2, 32'h0, 32'h0, 32'h0, 32'h42a267f0, 32'h0};
test_input[3200:3207] = '{32'h4215f330, 32'h42812382, 32'h4297cd9d, 32'h416370d3, 32'h42094153, 32'h422b5801, 32'h40eb647e, 32'hc22da964};
test_output[3200:3207] = '{32'h4215f330, 32'h42812382, 32'h4297cd9d, 32'h416370d3, 32'h42094153, 32'h422b5801, 32'h40eb647e, 32'h0};
test_input[3208:3215] = '{32'hc2ac1c5a, 32'h42b7e066, 32'h428d69e7, 32'hc29d1360, 32'hc2272081, 32'hc2aa93ab, 32'hc209f17f, 32'h41ebc950};
test_output[3208:3215] = '{32'h0, 32'h42b7e066, 32'h428d69e7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ebc950};
test_input[3216:3223] = '{32'hc2202fc1, 32'h4297abd7, 32'h3f3e7242, 32'h413c8743, 32'hc207eea2, 32'h4259bbdb, 32'hc28af922, 32'hc22fcfde};
test_output[3216:3223] = '{32'h0, 32'h4297abd7, 32'h3f3e7242, 32'h413c8743, 32'h0, 32'h4259bbdb, 32'h0, 32'h0};
test_input[3224:3231] = '{32'hc2bbdc98, 32'h42bb5a77, 32'h420400de, 32'hc286a254, 32'h41726e7d, 32'h426a7d82, 32'hc2101b42, 32'h427c6907};
test_output[3224:3231] = '{32'h0, 32'h42bb5a77, 32'h420400de, 32'h0, 32'h41726e7d, 32'h426a7d82, 32'h0, 32'h427c6907};
test_input[3232:3239] = '{32'hc2b47e4b, 32'hc2150ec4, 32'hc27113fc, 32'h419b3a67, 32'hc21a27a2, 32'h42b7057f, 32'hc2779f02, 32'h42813d09};
test_output[3232:3239] = '{32'h0, 32'h0, 32'h0, 32'h419b3a67, 32'h0, 32'h42b7057f, 32'h0, 32'h42813d09};
test_input[3240:3247] = '{32'hc1acc650, 32'h427d582b, 32'hc0498836, 32'hc2849f49, 32'h41f7f6b5, 32'hc2142d5f, 32'hc1a9296e, 32'h42a02be9};
test_output[3240:3247] = '{32'h0, 32'h427d582b, 32'h0, 32'h0, 32'h41f7f6b5, 32'h0, 32'h0, 32'h42a02be9};
test_input[3248:3255] = '{32'h41fede11, 32'hc2c11f54, 32'h413eac2c, 32'hc2b3a46c, 32'hc1e63163, 32'h402ee87d, 32'h42041f85, 32'hbfe154a3};
test_output[3248:3255] = '{32'h41fede11, 32'h0, 32'h413eac2c, 32'h0, 32'h0, 32'h402ee87d, 32'h42041f85, 32'h0};
test_input[3256:3263] = '{32'h40d7f564, 32'hc1bfc35d, 32'h421e5df8, 32'hc2351ff0, 32'hc1ee804f, 32'hc2146916, 32'hc1a493b0, 32'h41bce2ea};
test_output[3256:3263] = '{32'h40d7f564, 32'h0, 32'h421e5df8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41bce2ea};
test_input[3264:3271] = '{32'hc1faa419, 32'hc1584ea9, 32'h42c6a02a, 32'h41efca73, 32'h4211c66e, 32'hc29b6257, 32'h40f9b69a, 32'h4050de65};
test_output[3264:3271] = '{32'h0, 32'h0, 32'h42c6a02a, 32'h41efca73, 32'h4211c66e, 32'h0, 32'h40f9b69a, 32'h4050de65};
test_input[3272:3279] = '{32'h42a1abe4, 32'hc1a309fb, 32'hbfd49ee0, 32'hc2ad7c33, 32'hc2936b2e, 32'h427c1f4a, 32'h4280f612, 32'h42817c54};
test_output[3272:3279] = '{32'h42a1abe4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427c1f4a, 32'h4280f612, 32'h42817c54};
test_input[3280:3287] = '{32'hc22b664a, 32'h41145546, 32'hc24eef3c, 32'hc26dc8c8, 32'h42a5e200, 32'h4224f89f, 32'hc24cc902, 32'h428da7ba};
test_output[3280:3287] = '{32'h0, 32'h41145546, 32'h0, 32'h0, 32'h42a5e200, 32'h4224f89f, 32'h0, 32'h428da7ba};
test_input[3288:3295] = '{32'hc1f5ecb7, 32'h42b4c600, 32'h403bc1be, 32'hc2a437d1, 32'h41cb856a, 32'hc1efd0e7, 32'hc2b53895, 32'h412b3327};
test_output[3288:3295] = '{32'h0, 32'h42b4c600, 32'h403bc1be, 32'h0, 32'h41cb856a, 32'h0, 32'h0, 32'h412b3327};
test_input[3296:3303] = '{32'hc1923dad, 32'hc28caa60, 32'h3f624a33, 32'h41135b65, 32'h41802b58, 32'hc281dce1, 32'h42821391, 32'h42a050ba};
test_output[3296:3303] = '{32'h0, 32'h0, 32'h3f624a33, 32'h41135b65, 32'h41802b58, 32'h0, 32'h42821391, 32'h42a050ba};
test_input[3304:3311] = '{32'h424034b2, 32'h4283a0f7, 32'h40e284e3, 32'hc2ba166e, 32'hc287c44a, 32'h421eb89c, 32'hc18ca421, 32'h4261d684};
test_output[3304:3311] = '{32'h424034b2, 32'h4283a0f7, 32'h40e284e3, 32'h0, 32'h0, 32'h421eb89c, 32'h0, 32'h4261d684};
test_input[3312:3319] = '{32'hc1a933c1, 32'hc11e359a, 32'h42410241, 32'h422901d3, 32'h403fb749, 32'hc1065f75, 32'h42b82d42, 32'hc2ac51d7};
test_output[3312:3319] = '{32'h0, 32'h0, 32'h42410241, 32'h422901d3, 32'h403fb749, 32'h0, 32'h42b82d42, 32'h0};
test_input[3320:3327] = '{32'h42b5e9a7, 32'h41a76a0e, 32'h42ae95f1, 32'hc2145cba, 32'h428a440b, 32'hc2ad6e74, 32'h412dfdda, 32'h41beb416};
test_output[3320:3327] = '{32'h42b5e9a7, 32'h41a76a0e, 32'h42ae95f1, 32'h0, 32'h428a440b, 32'h0, 32'h412dfdda, 32'h41beb416};
test_input[3328:3335] = '{32'h4143723a, 32'h4245e385, 32'hc271702f, 32'hc2351302, 32'hc27f3c98, 32'hc0bd85ca, 32'hc2819a21, 32'hc2229edf};
test_output[3328:3335] = '{32'h4143723a, 32'h4245e385, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3336:3343] = '{32'h41d7af7b, 32'hc290d2f1, 32'h41d888f6, 32'h42b03d10, 32'hc21ecd19, 32'hc22d381a, 32'hc2bb1bbb, 32'h423205b5};
test_output[3336:3343] = '{32'h41d7af7b, 32'h0, 32'h41d888f6, 32'h42b03d10, 32'h0, 32'h0, 32'h0, 32'h423205b5};
test_input[3344:3351] = '{32'hc2372527, 32'hc19f56a7, 32'hc27c10d0, 32'h42b32105, 32'hc2030ca2, 32'h422241d5, 32'hc2b1bf50, 32'hc288f0ca};
test_output[3344:3351] = '{32'h0, 32'h0, 32'h0, 32'h42b32105, 32'h0, 32'h422241d5, 32'h0, 32'h0};
test_input[3352:3359] = '{32'h42a06c4e, 32'h42470a80, 32'hc2a97bbc, 32'hc2846527, 32'h42bc94b6, 32'h42aabfb2, 32'h428cee12, 32'h4203cd0f};
test_output[3352:3359] = '{32'h42a06c4e, 32'h42470a80, 32'h0, 32'h0, 32'h42bc94b6, 32'h42aabfb2, 32'h428cee12, 32'h4203cd0f};
test_input[3360:3367] = '{32'h425bdb25, 32'hc20d8a94, 32'hc0fb1d52, 32'hc178bdd8, 32'h4042209f, 32'h41e8ac75, 32'hc24e1a78, 32'h42bb4bd8};
test_output[3360:3367] = '{32'h425bdb25, 32'h0, 32'h0, 32'h0, 32'h4042209f, 32'h41e8ac75, 32'h0, 32'h42bb4bd8};
test_input[3368:3375] = '{32'hc2b5b9e4, 32'h4246f2a5, 32'hc1c50f3f, 32'h42bdf88a, 32'h425a148e, 32'h41c3d67f, 32'hc26469e6, 32'hc2743d53};
test_output[3368:3375] = '{32'h0, 32'h4246f2a5, 32'h0, 32'h42bdf88a, 32'h425a148e, 32'h41c3d67f, 32'h0, 32'h0};
test_input[3376:3383] = '{32'h428f13ba, 32'h410a46d0, 32'hc0aec1a9, 32'hc2857a72, 32'h403d39ba, 32'hc01c283b, 32'h424aa09f, 32'hbf6fc717};
test_output[3376:3383] = '{32'h428f13ba, 32'h410a46d0, 32'h0, 32'h0, 32'h403d39ba, 32'h0, 32'h424aa09f, 32'h0};
test_input[3384:3391] = '{32'h42a10b72, 32'h4244326c, 32'hc238e2a7, 32'h42393e12, 32'hbf92f55f, 32'hc2a2745a, 32'hc1b6cd61, 32'hc21c68a4};
test_output[3384:3391] = '{32'h42a10b72, 32'h4244326c, 32'h0, 32'h42393e12, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3392:3399] = '{32'hc2748b26, 32'h41c4e035, 32'h4260aa40, 32'hc28a551c, 32'h42aaa3f3, 32'hc2b3bb8f, 32'h41e2f1e8, 32'hc2c78449};
test_output[3392:3399] = '{32'h0, 32'h41c4e035, 32'h4260aa40, 32'h0, 32'h42aaa3f3, 32'h0, 32'h41e2f1e8, 32'h0};
test_input[3400:3407] = '{32'hc29e9cde, 32'h42a44114, 32'hc233e48f, 32'h41420b49, 32'hc2a43f12, 32'h423f6770, 32'h415c2471, 32'h42686e77};
test_output[3400:3407] = '{32'h0, 32'h42a44114, 32'h0, 32'h41420b49, 32'h0, 32'h423f6770, 32'h415c2471, 32'h42686e77};
test_input[3408:3415] = '{32'hc26ed21a, 32'hc255f4d0, 32'h41cdeb79, 32'hc2bd4702, 32'hc2ade681, 32'h420ae52e, 32'hc12bcf5a, 32'h41b4388e};
test_output[3408:3415] = '{32'h0, 32'h0, 32'h41cdeb79, 32'h0, 32'h0, 32'h420ae52e, 32'h0, 32'h41b4388e};
test_input[3416:3423] = '{32'hc2c61c6a, 32'h40e4608a, 32'hc2132915, 32'hc29f0d04, 32'h428e677e, 32'hc22e7124, 32'h42bcf333, 32'hc1196514};
test_output[3416:3423] = '{32'h0, 32'h40e4608a, 32'h0, 32'h0, 32'h428e677e, 32'h0, 32'h42bcf333, 32'h0};
test_input[3424:3431] = '{32'h4250cb38, 32'hc170c868, 32'hc210a509, 32'h42342423, 32'h3ff1286f, 32'hc1b95ee3, 32'hc23694e7, 32'hc242b17a};
test_output[3424:3431] = '{32'h4250cb38, 32'h0, 32'h0, 32'h42342423, 32'h3ff1286f, 32'h0, 32'h0, 32'h0};
test_input[3432:3439] = '{32'h42335384, 32'hc2bb4da0, 32'hc1d974c3, 32'hc2b94ddb, 32'hc1f1813e, 32'hc2935eb1, 32'hc246bab1, 32'h42b65b55};
test_output[3432:3439] = '{32'h42335384, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b65b55};
test_input[3440:3447] = '{32'hc2af5aec, 32'hc2b2b68a, 32'hc22460c1, 32'hbf6c2fc7, 32'h4285aa4a, 32'hc2b455e0, 32'hc28622a4, 32'h423969bf};
test_output[3440:3447] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4285aa4a, 32'h0, 32'h0, 32'h423969bf};
test_input[3448:3455] = '{32'h4198b49d, 32'h4243eea9, 32'hc167807d, 32'hc2915855, 32'hc2a78730, 32'h4240924a, 32'hc1c73ab1, 32'hc23d86ca};
test_output[3448:3455] = '{32'h4198b49d, 32'h4243eea9, 32'h0, 32'h0, 32'h0, 32'h4240924a, 32'h0, 32'h0};
test_input[3456:3463] = '{32'h40f9a2c3, 32'hc2c64492, 32'h3f576e73, 32'hc143752d, 32'h42669660, 32'hc24de6d1, 32'hc2c00b00, 32'hc118be76};
test_output[3456:3463] = '{32'h40f9a2c3, 32'h0, 32'h3f576e73, 32'h0, 32'h42669660, 32'h0, 32'h0, 32'h0};
test_input[3464:3471] = '{32'hc2bac218, 32'h419b0ff1, 32'h4180ada7, 32'h425f1d37, 32'hc28dccfe, 32'hc137a1e1, 32'h427eb165, 32'hc2843d52};
test_output[3464:3471] = '{32'h0, 32'h419b0ff1, 32'h4180ada7, 32'h425f1d37, 32'h0, 32'h0, 32'h427eb165, 32'h0};
test_input[3472:3479] = '{32'hc2a639e1, 32'h42913d12, 32'hc2378ad5, 32'h4289493f, 32'hc18d3989, 32'h42285ec5, 32'h4244e96a, 32'hc21f5307};
test_output[3472:3479] = '{32'h0, 32'h42913d12, 32'h0, 32'h4289493f, 32'h0, 32'h42285ec5, 32'h4244e96a, 32'h0};
test_input[3480:3487] = '{32'h4217c9de, 32'h4238df60, 32'hc0da8559, 32'hc2c4e65a, 32'hc1f805f6, 32'hc1d8058e, 32'hc1baa1b7, 32'hc2ae9667};
test_output[3480:3487] = '{32'h4217c9de, 32'h4238df60, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3488:3495] = '{32'h426c8769, 32'h429c1195, 32'hc21d94a1, 32'h3fd54100, 32'hc2566415, 32'h42302abc, 32'h42905968, 32'hc192ab2b};
test_output[3488:3495] = '{32'h426c8769, 32'h429c1195, 32'h0, 32'h3fd54100, 32'h0, 32'h42302abc, 32'h42905968, 32'h0};
test_input[3496:3503] = '{32'h41c243a5, 32'h3e2e5f3d, 32'hbfba9f45, 32'h42898253, 32'hc21711c6, 32'h42ac4a73, 32'hc2512e59, 32'h42c764ab};
test_output[3496:3503] = '{32'h41c243a5, 32'h3e2e5f3d, 32'h0, 32'h42898253, 32'h0, 32'h42ac4a73, 32'h0, 32'h42c764ab};
test_input[3504:3511] = '{32'hc294ba81, 32'h426fd261, 32'h40de9b49, 32'h42052131, 32'hc203a903, 32'hc292a5e4, 32'h42bcd1af, 32'h42550e8a};
test_output[3504:3511] = '{32'h0, 32'h426fd261, 32'h40de9b49, 32'h42052131, 32'h0, 32'h0, 32'h42bcd1af, 32'h42550e8a};
test_input[3512:3519] = '{32'h427229a2, 32'hc2962db4, 32'h3f81db0d, 32'h427a56f5, 32'hc17c5c74, 32'h4261ddc3, 32'h4280e64e, 32'h423e8d90};
test_output[3512:3519] = '{32'h427229a2, 32'h0, 32'h3f81db0d, 32'h427a56f5, 32'h0, 32'h4261ddc3, 32'h4280e64e, 32'h423e8d90};
test_input[3520:3527] = '{32'hbe995c43, 32'h428e8368, 32'h3f119cae, 32'hc25e7774, 32'hc14d2126, 32'hc0b1f0f8, 32'hc26a093a, 32'hc23e0984};
test_output[3520:3527] = '{32'h0, 32'h428e8368, 32'h3f119cae, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3528:3535] = '{32'h42605d35, 32'h42bfbbec, 32'hc2c60693, 32'h428434df, 32'h40fc9bdd, 32'hc27a292e, 32'hc2af1aab, 32'h42a733ed};
test_output[3528:3535] = '{32'h42605d35, 32'h42bfbbec, 32'h0, 32'h428434df, 32'h40fc9bdd, 32'h0, 32'h0, 32'h42a733ed};
test_input[3536:3543] = '{32'h42be64b4, 32'h428a62fc, 32'h420ac4ab, 32'h40f2555e, 32'hc286829c, 32'h426d031f, 32'hc198b608, 32'h4116e618};
test_output[3536:3543] = '{32'h42be64b4, 32'h428a62fc, 32'h420ac4ab, 32'h40f2555e, 32'h0, 32'h426d031f, 32'h0, 32'h4116e618};
test_input[3544:3551] = '{32'h428b7a5a, 32'hc2b08b0f, 32'hc2c21e3c, 32'h4183c6ae, 32'hc159f5db, 32'hc27f83a2, 32'hc121f4ae, 32'h4198eb25};
test_output[3544:3551] = '{32'h428b7a5a, 32'h0, 32'h0, 32'h4183c6ae, 32'h0, 32'h0, 32'h0, 32'h4198eb25};
test_input[3552:3559] = '{32'hc0ca331a, 32'h428c848b, 32'h41d0a59d, 32'h42b7b928, 32'hc2519927, 32'hc2480617, 32'h4194beaf, 32'h4154e51c};
test_output[3552:3559] = '{32'h0, 32'h428c848b, 32'h41d0a59d, 32'h42b7b928, 32'h0, 32'h0, 32'h4194beaf, 32'h4154e51c};
test_input[3560:3567] = '{32'h41253a34, 32'h41b1b2f8, 32'hc2c5d8e4, 32'hc0fead2c, 32'hc28c4228, 32'h4120f44c, 32'hc2694bc5, 32'h420cd48e};
test_output[3560:3567] = '{32'h41253a34, 32'h41b1b2f8, 32'h0, 32'h0, 32'h0, 32'h4120f44c, 32'h0, 32'h420cd48e};
test_input[3568:3575] = '{32'h41befc20, 32'hc1ea4a21, 32'hc262dff8, 32'hc2736592, 32'hc1551b68, 32'hc110f501, 32'hc2aaaad3, 32'hc0aac5b7};
test_output[3568:3575] = '{32'h41befc20, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3576:3583] = '{32'h41efff9d, 32'h42302fec, 32'hc2a0369e, 32'h4216fab1, 32'hc2a8eb0f, 32'h423343f3, 32'hc29592f6, 32'hc2235f5d};
test_output[3576:3583] = '{32'h41efff9d, 32'h42302fec, 32'h0, 32'h4216fab1, 32'h0, 32'h423343f3, 32'h0, 32'h0};
test_input[3584:3591] = '{32'hc20cf50c, 32'hc231ecda, 32'h42abb73f, 32'h4259e4ac, 32'hc286f310, 32'h42b3d0d6, 32'hc18d6fd2, 32'hc1145514};
test_output[3584:3591] = '{32'h0, 32'h0, 32'h42abb73f, 32'h4259e4ac, 32'h0, 32'h42b3d0d6, 32'h0, 32'h0};
test_input[3592:3599] = '{32'h42532173, 32'hc148db93, 32'h410f1555, 32'hc2b2b5f1, 32'hc0885cb5, 32'h429ae174, 32'hc2c3afa3, 32'hbf138473};
test_output[3592:3599] = '{32'h42532173, 32'h0, 32'h410f1555, 32'h0, 32'h0, 32'h429ae174, 32'h0, 32'h0};
test_input[3600:3607] = '{32'h41185884, 32'h418eeed6, 32'hc0bf7576, 32'hc28c0c5b, 32'hc24c0ca4, 32'h42a03dc1, 32'h42b9e381, 32'hc1f766bd};
test_output[3600:3607] = '{32'h41185884, 32'h418eeed6, 32'h0, 32'h0, 32'h0, 32'h42a03dc1, 32'h42b9e381, 32'h0};
test_input[3608:3615] = '{32'h4268428b, 32'h42098704, 32'h42a75ebb, 32'hc18e9055, 32'h42a7b5d0, 32'hc2bf5f33, 32'h41dc6c7f, 32'hc1eb9901};
test_output[3608:3615] = '{32'h4268428b, 32'h42098704, 32'h42a75ebb, 32'h0, 32'h42a7b5d0, 32'h0, 32'h41dc6c7f, 32'h0};
test_input[3616:3623] = '{32'h418b6997, 32'h42b4faae, 32'h42bdb848, 32'hc1ef610a, 32'hc296944c, 32'hc2b8905d, 32'hc2a79caa, 32'h423ec3e3};
test_output[3616:3623] = '{32'h418b6997, 32'h42b4faae, 32'h42bdb848, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423ec3e3};
test_input[3624:3631] = '{32'hc2a265ed, 32'hc1f4f52c, 32'h42c3b8d7, 32'hc1636227, 32'hc1c986d9, 32'hc1fbab22, 32'hc281bbf4, 32'h42ba1a71};
test_output[3624:3631] = '{32'h0, 32'h0, 32'h42c3b8d7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ba1a71};
test_input[3632:3639] = '{32'h42039698, 32'hc1cc8a85, 32'h40d37d53, 32'h41bb7302, 32'hc24beac8, 32'h4293fe35, 32'hc2902233, 32'hc2a437e2};
test_output[3632:3639] = '{32'h42039698, 32'h0, 32'h40d37d53, 32'h41bb7302, 32'h0, 32'h4293fe35, 32'h0, 32'h0};
test_input[3640:3647] = '{32'h429f16ad, 32'h420eccb0, 32'hc234e4a7, 32'h41b27b9a, 32'hc092fc28, 32'h4211fae8, 32'h3f7c26b9, 32'h42b7d6b1};
test_output[3640:3647] = '{32'h429f16ad, 32'h420eccb0, 32'h0, 32'h41b27b9a, 32'h0, 32'h4211fae8, 32'h3f7c26b9, 32'h42b7d6b1};
test_input[3648:3655] = '{32'h40a8daf2, 32'h42257c7c, 32'h41ae5632, 32'hc2aa8388, 32'hc1539fbf, 32'h429a9696, 32'h4283746f, 32'h427347ab};
test_output[3648:3655] = '{32'h40a8daf2, 32'h42257c7c, 32'h41ae5632, 32'h0, 32'h0, 32'h429a9696, 32'h4283746f, 32'h427347ab};
test_input[3656:3663] = '{32'h42c2df4d, 32'hc27116e6, 32'hc2665b67, 32'h4184a7c2, 32'h409b7243, 32'h41ca78a3, 32'hc16bab37, 32'h42ab5924};
test_output[3656:3663] = '{32'h42c2df4d, 32'h0, 32'h0, 32'h4184a7c2, 32'h409b7243, 32'h41ca78a3, 32'h0, 32'h42ab5924};
test_input[3664:3671] = '{32'h42443179, 32'h426f60ea, 32'hc29bda2d, 32'hc2ae5f53, 32'h42825e9d, 32'h427ee31c, 32'hc2c655e0, 32'hc107a624};
test_output[3664:3671] = '{32'h42443179, 32'h426f60ea, 32'h0, 32'h0, 32'h42825e9d, 32'h427ee31c, 32'h0, 32'h0};
test_input[3672:3679] = '{32'h4282c862, 32'hc1911a8b, 32'h428cdeb9, 32'hc2b7fa9b, 32'hc2beeb39, 32'h42035cad, 32'hc203b7eb, 32'h4271f7fc};
test_output[3672:3679] = '{32'h4282c862, 32'h0, 32'h428cdeb9, 32'h0, 32'h0, 32'h42035cad, 32'h0, 32'h4271f7fc};
test_input[3680:3687] = '{32'hc28a86d7, 32'h41d9daa5, 32'hc0739e11, 32'h421b03a0, 32'hc206a485, 32'h42949fe9, 32'hc19a1269, 32'hc1ea68b0};
test_output[3680:3687] = '{32'h0, 32'h41d9daa5, 32'h0, 32'h421b03a0, 32'h0, 32'h42949fe9, 32'h0, 32'h0};
test_input[3688:3695] = '{32'hc2835760, 32'hc22da0c2, 32'hc26c32f2, 32'h428de8e0, 32'h42477a00, 32'hc0de0386, 32'hc18cb6cf, 32'h428b469c};
test_output[3688:3695] = '{32'h0, 32'h0, 32'h0, 32'h428de8e0, 32'h42477a00, 32'h0, 32'h0, 32'h428b469c};
test_input[3696:3703] = '{32'hc11700b0, 32'h42974ff1, 32'hc1667240, 32'hc290731b, 32'hc2379dd3, 32'hc26286a6, 32'hc29fedbd, 32'hc1500b64};
test_output[3696:3703] = '{32'h0, 32'h42974ff1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3704:3711] = '{32'hc2452c46, 32'h419a66df, 32'h41e51bd9, 32'h40bff14a, 32'h41cfc94a, 32'hc1bb73c0, 32'hc26dfb80, 32'h422fc269};
test_output[3704:3711] = '{32'h0, 32'h419a66df, 32'h41e51bd9, 32'h40bff14a, 32'h41cfc94a, 32'h0, 32'h0, 32'h422fc269};
test_input[3712:3719] = '{32'hc12d3be2, 32'hc2b8a156, 32'h42a848b2, 32'h42991c19, 32'h42ad0068, 32'hc2931406, 32'hc1987772, 32'hc2577db1};
test_output[3712:3719] = '{32'h0, 32'h0, 32'h42a848b2, 32'h42991c19, 32'h42ad0068, 32'h0, 32'h0, 32'h0};
test_input[3720:3727] = '{32'h4084ab76, 32'hc25db28e, 32'h422520e7, 32'h425378fb, 32'h4202c028, 32'hc1d1aed1, 32'hc28de5ea, 32'hc2a5ede7};
test_output[3720:3727] = '{32'h4084ab76, 32'h0, 32'h422520e7, 32'h425378fb, 32'h4202c028, 32'h0, 32'h0, 32'h0};
test_input[3728:3735] = '{32'hc1abc7e0, 32'h425004e1, 32'hc2a01fc8, 32'h424ac540, 32'hc262d309, 32'hc2c4acf5, 32'hc2938998, 32'hc2abab72};
test_output[3728:3735] = '{32'h0, 32'h425004e1, 32'h0, 32'h424ac540, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3736:3743] = '{32'hc2b7c27c, 32'hc2946b04, 32'h41234aa9, 32'hc1118168, 32'hc2a668c8, 32'h42977dc3, 32'hc09604a3, 32'h4255b8cf};
test_output[3736:3743] = '{32'h0, 32'h0, 32'h41234aa9, 32'h0, 32'h0, 32'h42977dc3, 32'h0, 32'h4255b8cf};
test_input[3744:3751] = '{32'hc2216ac0, 32'h42364b25, 32'h42a1c8ad, 32'h3f854d9e, 32'hc2791629, 32'h426351d7, 32'hc29662ea, 32'hc276c702};
test_output[3744:3751] = '{32'h0, 32'h42364b25, 32'h42a1c8ad, 32'h3f854d9e, 32'h0, 32'h426351d7, 32'h0, 32'h0};
test_input[3752:3759] = '{32'hc2b9c4da, 32'hc22be3b0, 32'hc295a10a, 32'h416e1df7, 32'hc0f0d3e2, 32'h425e5751, 32'h4285a7b8, 32'hc239c81b};
test_output[3752:3759] = '{32'h0, 32'h0, 32'h0, 32'h416e1df7, 32'h0, 32'h425e5751, 32'h4285a7b8, 32'h0};
test_input[3760:3767] = '{32'h41369e79, 32'hc2c58e6f, 32'hc19a171d, 32'hc1e960f3, 32'h42873020, 32'hbe86e0b1, 32'hc293f78f, 32'hc209846c};
test_output[3760:3767] = '{32'h41369e79, 32'h0, 32'h0, 32'h0, 32'h42873020, 32'h0, 32'h0, 32'h0};
test_input[3768:3775] = '{32'h401243be, 32'hc04f405b, 32'h42c2c27c, 32'hc2401e4f, 32'hc19d3732, 32'h41a6d16c, 32'hc260ee57, 32'h4237e84c};
test_output[3768:3775] = '{32'h401243be, 32'h0, 32'h42c2c27c, 32'h0, 32'h0, 32'h41a6d16c, 32'h0, 32'h4237e84c};
test_input[3776:3783] = '{32'h42c1b34d, 32'hc2b15efa, 32'h4273c778, 32'hc257608c, 32'hc20e0c55, 32'h41c03728, 32'hc1be9251, 32'h4254a6de};
test_output[3776:3783] = '{32'h42c1b34d, 32'h0, 32'h4273c778, 32'h0, 32'h0, 32'h41c03728, 32'h0, 32'h4254a6de};
test_input[3784:3791] = '{32'hc0f6e8ff, 32'hc1022ef8, 32'hc2336955, 32'h42889df1, 32'h42878052, 32'hc28f10e9, 32'hc21bad24, 32'hc2af4152};
test_output[3784:3791] = '{32'h0, 32'h0, 32'h0, 32'h42889df1, 32'h42878052, 32'h0, 32'h0, 32'h0};
test_input[3792:3799] = '{32'h41714ba2, 32'hc234b04a, 32'hc29308b4, 32'hc29e6387, 32'h429c5ed7, 32'h41d9d7cf, 32'hc2b8ca0b, 32'h42a257a3};
test_output[3792:3799] = '{32'h41714ba2, 32'h0, 32'h0, 32'h0, 32'h429c5ed7, 32'h41d9d7cf, 32'h0, 32'h42a257a3};
test_input[3800:3807] = '{32'h420bcd4a, 32'hc25a2433, 32'hc137ad1f, 32'hc2ba7652, 32'hc2162d11, 32'h402f346f, 32'h423dea55, 32'h42a499b6};
test_output[3800:3807] = '{32'h420bcd4a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h402f346f, 32'h423dea55, 32'h42a499b6};
test_input[3808:3815] = '{32'hc20b8a35, 32'h428ccec8, 32'h42879a16, 32'h42bfabb5, 32'h424bee84, 32'hc256cd18, 32'hc1e4c041, 32'h3fd94a72};
test_output[3808:3815] = '{32'h0, 32'h428ccec8, 32'h42879a16, 32'h42bfabb5, 32'h424bee84, 32'h0, 32'h0, 32'h3fd94a72};
test_input[3816:3823] = '{32'h41b41f58, 32'h42373f23, 32'hc27ea847, 32'h41d6361e, 32'hc1bb3afc, 32'hc1100cf9, 32'h4193d2e2, 32'hc2bc6667};
test_output[3816:3823] = '{32'h41b41f58, 32'h42373f23, 32'h0, 32'h41d6361e, 32'h0, 32'h0, 32'h4193d2e2, 32'h0};
test_input[3824:3831] = '{32'h42c6e56f, 32'h4221b0ca, 32'h4294b0b1, 32'h42212d8b, 32'hc2a3f77c, 32'hc28c644f, 32'hc29d5d0b, 32'hc28fdc5e};
test_output[3824:3831] = '{32'h42c6e56f, 32'h4221b0ca, 32'h4294b0b1, 32'h42212d8b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3832:3839] = '{32'hc29b33e1, 32'hc2950997, 32'hc1951e86, 32'h4296dc5e, 32'hc1cbbe12, 32'hc2992e3e, 32'h423b9560, 32'hc2c23dc9};
test_output[3832:3839] = '{32'h0, 32'h0, 32'h0, 32'h4296dc5e, 32'h0, 32'h0, 32'h423b9560, 32'h0};
test_input[3840:3847] = '{32'hc0e4a2c2, 32'hc1f40dd7, 32'hc244e738, 32'hc24b88bd, 32'hc02e9295, 32'h428bc232, 32'hc24d78a3, 32'h42a38a12};
test_output[3840:3847] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428bc232, 32'h0, 32'h42a38a12};
test_input[3848:3855] = '{32'hc1c7367c, 32'h4260c538, 32'h428acd34, 32'h421ab787, 32'h41781da5, 32'hc2c4e6ed, 32'hc271f11c, 32'h425cf568};
test_output[3848:3855] = '{32'h0, 32'h4260c538, 32'h428acd34, 32'h421ab787, 32'h41781da5, 32'h0, 32'h0, 32'h425cf568};
test_input[3856:3863] = '{32'h41951443, 32'hc28985e5, 32'h429a479a, 32'h422427c9, 32'hc22f5d50, 32'h4241c8ab, 32'h42b4aa62, 32'h42545bf9};
test_output[3856:3863] = '{32'h41951443, 32'h0, 32'h429a479a, 32'h422427c9, 32'h0, 32'h4241c8ab, 32'h42b4aa62, 32'h42545bf9};
test_input[3864:3871] = '{32'h4271033c, 32'h4283045e, 32'h4210b887, 32'hc200c865, 32'hc279e519, 32'h42ae3742, 32'h42a7eae1, 32'h42947510};
test_output[3864:3871] = '{32'h4271033c, 32'h4283045e, 32'h4210b887, 32'h0, 32'h0, 32'h42ae3742, 32'h42a7eae1, 32'h42947510};
test_input[3872:3879] = '{32'h4113ce1f, 32'h417580e2, 32'hc27d4a59, 32'hc29fcb38, 32'hc2c130c5, 32'hc2a4fcfe, 32'hc256fc6c, 32'hc00aea87};
test_output[3872:3879] = '{32'h4113ce1f, 32'h417580e2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3880:3887] = '{32'h41628937, 32'h4243691d, 32'h420e8417, 32'h42516844, 32'h42ba7102, 32'hc08c7897, 32'hc262377c, 32'hc26ae61e};
test_output[3880:3887] = '{32'h41628937, 32'h4243691d, 32'h420e8417, 32'h42516844, 32'h42ba7102, 32'h0, 32'h0, 32'h0};
test_input[3888:3895] = '{32'hc2a07ac2, 32'hc2210c49, 32'h41365a04, 32'hc187797c, 32'hc21f6057, 32'h42932293, 32'h423b5299, 32'h42c61827};
test_output[3888:3895] = '{32'h0, 32'h0, 32'h41365a04, 32'h0, 32'h0, 32'h42932293, 32'h423b5299, 32'h42c61827};
test_input[3896:3903] = '{32'hc1464065, 32'h42a953f5, 32'h42c0b246, 32'h416a7a3d, 32'hc19e2df1, 32'hc25fbdc5, 32'h4091f791, 32'hc251f3b6};
test_output[3896:3903] = '{32'h0, 32'h42a953f5, 32'h42c0b246, 32'h416a7a3d, 32'h0, 32'h0, 32'h4091f791, 32'h0};
test_input[3904:3911] = '{32'h41b6ede2, 32'h42837d37, 32'h4299bc75, 32'h42391212, 32'h40b6b8cf, 32'h41d70b8a, 32'h41a5b0e8, 32'hc156a448};
test_output[3904:3911] = '{32'h41b6ede2, 32'h42837d37, 32'h4299bc75, 32'h42391212, 32'h40b6b8cf, 32'h41d70b8a, 32'h41a5b0e8, 32'h0};
test_input[3912:3919] = '{32'h4226c559, 32'hc1a29e46, 32'hc2747712, 32'hc2bae3b7, 32'hc28a3f8b, 32'hc2162ce2, 32'hc2376b53, 32'h4113209a};
test_output[3912:3919] = '{32'h4226c559, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4113209a};
test_input[3920:3927] = '{32'hc2adc208, 32'hc185b2f5, 32'hc1888495, 32'h4203f103, 32'h42a7f04a, 32'h418846d3, 32'hc28395f0, 32'hc2b35cac};
test_output[3920:3927] = '{32'h0, 32'h0, 32'h0, 32'h4203f103, 32'h42a7f04a, 32'h418846d3, 32'h0, 32'h0};
test_input[3928:3935] = '{32'h4289d72c, 32'hc27be6d2, 32'h4263946c, 32'h42c51e9c, 32'hc150e0bf, 32'h419d6ac3, 32'hc252396b, 32'hc289ff92};
test_output[3928:3935] = '{32'h4289d72c, 32'h0, 32'h4263946c, 32'h42c51e9c, 32'h0, 32'h419d6ac3, 32'h0, 32'h0};
test_input[3936:3943] = '{32'hc25b088f, 32'h422b9e86, 32'hc2231fd0, 32'h4220a1ca, 32'h424030da, 32'h420f2344, 32'hc1752147, 32'hc0527a23};
test_output[3936:3943] = '{32'h0, 32'h422b9e86, 32'h0, 32'h4220a1ca, 32'h424030da, 32'h420f2344, 32'h0, 32'h0};
test_input[3944:3951] = '{32'hc14fa151, 32'h4003a54f, 32'h40d5058f, 32'h428f1ed7, 32'hc2252a13, 32'h4285c816, 32'h42958cea, 32'h41c8d92a};
test_output[3944:3951] = '{32'h0, 32'h4003a54f, 32'h40d5058f, 32'h428f1ed7, 32'h0, 32'h4285c816, 32'h42958cea, 32'h41c8d92a};
test_input[3952:3959] = '{32'hc2938314, 32'h42a5e86a, 32'h42554c11, 32'hc2b75a9a, 32'hc0e0e05b, 32'hc1b35bbb, 32'h412b62f5, 32'h401ffed2};
test_output[3952:3959] = '{32'h0, 32'h42a5e86a, 32'h42554c11, 32'h0, 32'h0, 32'h0, 32'h412b62f5, 32'h401ffed2};
test_input[3960:3967] = '{32'h429102d5, 32'h42275668, 32'h411e51f9, 32'hc0f7860c, 32'hc298f490, 32'hc2bb9e08, 32'h42a3ab40, 32'h419057a1};
test_output[3960:3967] = '{32'h429102d5, 32'h42275668, 32'h411e51f9, 32'h0, 32'h0, 32'h0, 32'h42a3ab40, 32'h419057a1};
test_input[3968:3975] = '{32'hc29b5c53, 32'hc1faf45f, 32'h40850ae0, 32'h41c02b8e, 32'h421e930c, 32'h428dba32, 32'hc11d9344, 32'h425a4e12};
test_output[3968:3975] = '{32'h0, 32'h0, 32'h40850ae0, 32'h41c02b8e, 32'h421e930c, 32'h428dba32, 32'h0, 32'h425a4e12};
test_input[3976:3983] = '{32'hc2c678a4, 32'h403915eb, 32'hbff551f3, 32'h41a90737, 32'h4278136f, 32'h41ee426b, 32'h41e96d5e, 32'h4217e1e7};
test_output[3976:3983] = '{32'h0, 32'h403915eb, 32'h0, 32'h41a90737, 32'h4278136f, 32'h41ee426b, 32'h41e96d5e, 32'h4217e1e7};
test_input[3984:3991] = '{32'hc21f04da, 32'h418bc849, 32'h42375cf2, 32'h41b21e1f, 32'h4054a215, 32'h4268a913, 32'hc2609de3, 32'h42835647};
test_output[3984:3991] = '{32'h0, 32'h418bc849, 32'h42375cf2, 32'h41b21e1f, 32'h4054a215, 32'h4268a913, 32'h0, 32'h42835647};
test_input[3992:3999] = '{32'h42950194, 32'h4294a629, 32'hc1bdaf9e, 32'h427583cd, 32'h428858e0, 32'h421b9fa7, 32'h413a4d30, 32'hc2269fed};
test_output[3992:3999] = '{32'h42950194, 32'h4294a629, 32'h0, 32'h427583cd, 32'h428858e0, 32'h421b9fa7, 32'h413a4d30, 32'h0};
test_input[4000:4007] = '{32'hc28ad4e1, 32'hc25441c0, 32'hc24352b8, 32'hc2920aa1, 32'h3db67356, 32'h427e9f45, 32'hc2c29c37, 32'hc27104a0};
test_output[4000:4007] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h3db67356, 32'h427e9f45, 32'h0, 32'h0};
test_input[4008:4015] = '{32'h42692c03, 32'hc2aad471, 32'h4128ea5e, 32'hc236016d, 32'hc08b859a, 32'hc29489a8, 32'h422ad6f7, 32'hc2c531e7};
test_output[4008:4015] = '{32'h42692c03, 32'h0, 32'h4128ea5e, 32'h0, 32'h0, 32'h0, 32'h422ad6f7, 32'h0};
test_input[4016:4023] = '{32'h427687b0, 32'hc255a57c, 32'hc2583c10, 32'h414945c6, 32'h42c6904f, 32'h41ab6be3, 32'h425c258a, 32'h427b0445};
test_output[4016:4023] = '{32'h427687b0, 32'h0, 32'h0, 32'h414945c6, 32'h42c6904f, 32'h41ab6be3, 32'h425c258a, 32'h427b0445};
test_input[4024:4031] = '{32'h41852b31, 32'h4193360f, 32'h41532a1d, 32'hc29ce278, 32'hc2251f79, 32'hc21b39c0, 32'h42b0b1a3, 32'h41d12882};
test_output[4024:4031] = '{32'h41852b31, 32'h4193360f, 32'h41532a1d, 32'h0, 32'h0, 32'h0, 32'h42b0b1a3, 32'h41d12882};
test_input[4032:4039] = '{32'hc2680f8a, 32'h427266bc, 32'hc042aec3, 32'h42c76cd7, 32'hc183bcd7, 32'hc2a0e659, 32'hc1686783, 32'hc28579aa};
test_output[4032:4039] = '{32'h0, 32'h427266bc, 32'h0, 32'h42c76cd7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4040:4047] = '{32'h42934c98, 32'hc191e383, 32'hc212d498, 32'hc2025557, 32'h426af430, 32'hc2834c51, 32'h415c21d7, 32'h42308caf};
test_output[4040:4047] = '{32'h42934c98, 32'h0, 32'h0, 32'h0, 32'h426af430, 32'h0, 32'h415c21d7, 32'h42308caf};
test_input[4048:4055] = '{32'h429b829a, 32'hc2106f6f, 32'hc2c587e6, 32'h4285e98c, 32'h42af3b3b, 32'h42a8caab, 32'hc2beab63, 32'hc2819968};
test_output[4048:4055] = '{32'h429b829a, 32'h0, 32'h0, 32'h4285e98c, 32'h42af3b3b, 32'h42a8caab, 32'h0, 32'h0};
test_input[4056:4063] = '{32'h42051031, 32'hc16be0a0, 32'hc24cd01c, 32'h42b2131f, 32'h42c5d861, 32'h4243d550, 32'h420921c9, 32'h42757d1c};
test_output[4056:4063] = '{32'h42051031, 32'h0, 32'h0, 32'h42b2131f, 32'h42c5d861, 32'h4243d550, 32'h420921c9, 32'h42757d1c};
test_input[4064:4071] = '{32'hc299eb13, 32'hc1d5d024, 32'hc222c919, 32'h405324df, 32'hc2a16cba, 32'hc11db7e6, 32'h42a29529, 32'hc2227e46};
test_output[4064:4071] = '{32'h0, 32'h0, 32'h0, 32'h405324df, 32'h0, 32'h0, 32'h42a29529, 32'h0};
test_input[4072:4079] = '{32'hc23d9727, 32'hc2c0fdaa, 32'h42a9eb8a, 32'hc25f9ee5, 32'hc2b52931, 32'h426a12a5, 32'hc2960f47, 32'hc1e30ac5};
test_output[4072:4079] = '{32'h0, 32'h0, 32'h42a9eb8a, 32'h0, 32'h0, 32'h426a12a5, 32'h0, 32'h0};
test_input[4080:4087] = '{32'hc2073a5a, 32'h42a3245a, 32'h4231f59a, 32'hc20ab9df, 32'hc29dd29a, 32'h42a16e46, 32'h427c3d3e, 32'h408d54f0};
test_output[4080:4087] = '{32'h0, 32'h42a3245a, 32'h4231f59a, 32'h0, 32'h0, 32'h42a16e46, 32'h427c3d3e, 32'h408d54f0};
test_input[4088:4095] = '{32'h428b2732, 32'hc236c231, 32'hc2a4ded4, 32'h41e0e5c1, 32'h41aae64f, 32'h42ae3c14, 32'hc2123a92, 32'hc00b1098};
test_output[4088:4095] = '{32'h428b2732, 32'h0, 32'h0, 32'h41e0e5c1, 32'h41aae64f, 32'h42ae3c14, 32'h0, 32'h0};
test_input[4096:4103] = '{32'h427605af, 32'h42b1304f, 32'hc21d3d61, 32'hc20d78b3, 32'hc20494f5, 32'h411de982, 32'h42a9aacd, 32'hc26caab3};
test_output[4096:4103] = '{32'h427605af, 32'h42b1304f, 32'h0, 32'h0, 32'h0, 32'h411de982, 32'h42a9aacd, 32'h0};
test_input[4104:4111] = '{32'h42871f19, 32'hc2bfa3a8, 32'h414a5422, 32'h42689cc6, 32'hc1c78c2d, 32'h4242532b, 32'hc2b47d3e, 32'hc2a172ee};
test_output[4104:4111] = '{32'h42871f19, 32'h0, 32'h414a5422, 32'h42689cc6, 32'h0, 32'h4242532b, 32'h0, 32'h0};
test_input[4112:4119] = '{32'hc28b2d26, 32'h426a873c, 32'h412192f8, 32'hc11a4aea, 32'hc0a1b014, 32'h41d56dce, 32'h409bd217, 32'hc180fcc3};
test_output[4112:4119] = '{32'h0, 32'h426a873c, 32'h412192f8, 32'h0, 32'h0, 32'h41d56dce, 32'h409bd217, 32'h0};
test_input[4120:4127] = '{32'h425aaadd, 32'h4287ee6e, 32'h41ad04d6, 32'h428c06cf, 32'h4152aa0c, 32'h41232432, 32'hc28e43d3, 32'hc0691347};
test_output[4120:4127] = '{32'h425aaadd, 32'h4287ee6e, 32'h41ad04d6, 32'h428c06cf, 32'h4152aa0c, 32'h41232432, 32'h0, 32'h0};
test_input[4128:4135] = '{32'hc150c25c, 32'hc25edd8d, 32'hc166fe4f, 32'h42a380d0, 32'h42171b8a, 32'h4058356b, 32'hc2c3a5b4, 32'hbe10efa4};
test_output[4128:4135] = '{32'h0, 32'h0, 32'h0, 32'h42a380d0, 32'h42171b8a, 32'h4058356b, 32'h0, 32'h0};
test_input[4136:4143] = '{32'h4200b623, 32'h4122e37f, 32'h427ecb3d, 32'hc28c03a8, 32'hc2a1464b, 32'h421c4bb3, 32'hc2b0f841, 32'hc0c848c4};
test_output[4136:4143] = '{32'h4200b623, 32'h4122e37f, 32'h427ecb3d, 32'h0, 32'h0, 32'h421c4bb3, 32'h0, 32'h0};
test_input[4144:4151] = '{32'hc299bd87, 32'h42ba5a89, 32'hc1d0ae6c, 32'h4290f890, 32'h41e8a82d, 32'hc2c17ea8, 32'hc266554a, 32'h42031257};
test_output[4144:4151] = '{32'h0, 32'h42ba5a89, 32'h0, 32'h4290f890, 32'h41e8a82d, 32'h0, 32'h0, 32'h42031257};
test_input[4152:4159] = '{32'h428b1527, 32'h4209e94b, 32'hc1ff368a, 32'hc2b86d84, 32'h41aeb305, 32'hc2b26aef, 32'hc273493f, 32'hc19b1fb5};
test_output[4152:4159] = '{32'h428b1527, 32'h4209e94b, 32'h0, 32'h0, 32'h41aeb305, 32'h0, 32'h0, 32'h0};
test_input[4160:4167] = '{32'hc287a8b0, 32'h42a381cc, 32'hc0628a8e, 32'hc2a08ff4, 32'hc2b734e6, 32'hc1cce593, 32'hc28acf6b, 32'hc27648c8};
test_output[4160:4167] = '{32'h0, 32'h42a381cc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4168:4175] = '{32'h423ff952, 32'h42bedf16, 32'hc233be39, 32'hc2a15431, 32'hc23998a9, 32'hc2ba073c, 32'h418a9149, 32'hc2274637};
test_output[4168:4175] = '{32'h423ff952, 32'h42bedf16, 32'h0, 32'h0, 32'h0, 32'h0, 32'h418a9149, 32'h0};
test_input[4176:4183] = '{32'hc1f1d151, 32'hc24124de, 32'h42b94460, 32'h418eff19, 32'hc18f4056, 32'hc012ab25, 32'h4234fb38, 32'hc231a3ed};
test_output[4176:4183] = '{32'h0, 32'h0, 32'h42b94460, 32'h418eff19, 32'h0, 32'h0, 32'h4234fb38, 32'h0};
test_input[4184:4191] = '{32'h42b2c571, 32'hc20afd6d, 32'hc299ff62, 32'hc29343ab, 32'hc2939886, 32'hc265f49b, 32'hc27d9f89, 32'hc10de5a5};
test_output[4184:4191] = '{32'h42b2c571, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4192:4199] = '{32'hc2aca4b8, 32'h419f6646, 32'hc2bf5af5, 32'hc295509c, 32'h41506d4e, 32'hc2acf154, 32'hc11fa8ff, 32'h41da427f};
test_output[4192:4199] = '{32'h0, 32'h419f6646, 32'h0, 32'h0, 32'h41506d4e, 32'h0, 32'h0, 32'h41da427f};
test_input[4200:4207] = '{32'hc28809cb, 32'hc2346722, 32'hc136cdbe, 32'h42956ad1, 32'hc26a9809, 32'hc28aa99b, 32'hc25cefb2, 32'h421e9455};
test_output[4200:4207] = '{32'h0, 32'h0, 32'h0, 32'h42956ad1, 32'h0, 32'h0, 32'h0, 32'h421e9455};
test_input[4208:4215] = '{32'h426a236a, 32'hc27b47b6, 32'h4236f1d8, 32'hc2a34e36, 32'h423008c3, 32'hc2a188a3, 32'h424aa90f, 32'h42771ebd};
test_output[4208:4215] = '{32'h426a236a, 32'h0, 32'h4236f1d8, 32'h0, 32'h423008c3, 32'h0, 32'h424aa90f, 32'h42771ebd};
test_input[4216:4223] = '{32'h41cec846, 32'h4206a8c2, 32'hc290d3ee, 32'h41ca13df, 32'h4230885b, 32'h40f5f8b4, 32'hc2c1d0d7, 32'h4285affe};
test_output[4216:4223] = '{32'h41cec846, 32'h4206a8c2, 32'h0, 32'h41ca13df, 32'h4230885b, 32'h40f5f8b4, 32'h0, 32'h4285affe};
test_input[4224:4231] = '{32'hc2a7ad66, 32'h41c7024b, 32'hc2ac6f4d, 32'h425e8bdd, 32'h423ac11e, 32'h4270e273, 32'h4282f346, 32'hc29038d0};
test_output[4224:4231] = '{32'h0, 32'h41c7024b, 32'h0, 32'h425e8bdd, 32'h423ac11e, 32'h4270e273, 32'h4282f346, 32'h0};
test_input[4232:4239] = '{32'hc2606825, 32'h417d2cfd, 32'hc1d0b786, 32'hc1e25cd0, 32'h41cf5be8, 32'hc1bdb2e2, 32'h41fc03d8, 32'hc20cb89d};
test_output[4232:4239] = '{32'h0, 32'h417d2cfd, 32'h0, 32'h0, 32'h41cf5be8, 32'h0, 32'h41fc03d8, 32'h0};
test_input[4240:4247] = '{32'hc2bf4cb9, 32'hc29c9661, 32'hc280c44e, 32'hc1628c65, 32'h4294e180, 32'hc2afc46c, 32'h42659fe5, 32'hc287d50d};
test_output[4240:4247] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4294e180, 32'h0, 32'h42659fe5, 32'h0};
test_input[4248:4255] = '{32'h42931d0d, 32'h42800058, 32'hc23c2669, 32'h420960c9, 32'h4188e96a, 32'h4281cf32, 32'h429c9f4f, 32'h42908406};
test_output[4248:4255] = '{32'h42931d0d, 32'h42800058, 32'h0, 32'h420960c9, 32'h4188e96a, 32'h4281cf32, 32'h429c9f4f, 32'h42908406};
test_input[4256:4263] = '{32'h40d79f85, 32'h423f0c5d, 32'h42395754, 32'hc2754a54, 32'h42b770fe, 32'h42a8f78f, 32'h4269ab91, 32'h413aca77};
test_output[4256:4263] = '{32'h40d79f85, 32'h423f0c5d, 32'h42395754, 32'h0, 32'h42b770fe, 32'h42a8f78f, 32'h4269ab91, 32'h413aca77};
test_input[4264:4271] = '{32'h4280eb3c, 32'hc2a95e84, 32'h42439cf6, 32'h423fab81, 32'h4276bf29, 32'h425560ed, 32'hc24d08f7, 32'h422e8f28};
test_output[4264:4271] = '{32'h4280eb3c, 32'h0, 32'h42439cf6, 32'h423fab81, 32'h4276bf29, 32'h425560ed, 32'h0, 32'h422e8f28};
test_input[4272:4279] = '{32'hc1605bc1, 32'hc28e11cf, 32'h422fb1cc, 32'h428cae70, 32'h41824500, 32'hc23ebf58, 32'h42392a25, 32'hc1fdfc99};
test_output[4272:4279] = '{32'h0, 32'h0, 32'h422fb1cc, 32'h428cae70, 32'h41824500, 32'h0, 32'h42392a25, 32'h0};
test_input[4280:4287] = '{32'h4090e592, 32'h42841dfa, 32'hc1914b40, 32'h42b6ab22, 32'h3f9746f1, 32'h42a3846a, 32'hc2a409fc, 32'h423f0971};
test_output[4280:4287] = '{32'h4090e592, 32'h42841dfa, 32'h0, 32'h42b6ab22, 32'h3f9746f1, 32'h42a3846a, 32'h0, 32'h423f0971};
test_input[4288:4295] = '{32'hc12dd80d, 32'hc25d11fc, 32'hc2a07ee9, 32'hc29c206b, 32'hc1902758, 32'h42bd7a42, 32'h4188cda5, 32'hc2bb24b5};
test_output[4288:4295] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bd7a42, 32'h4188cda5, 32'h0};
test_input[4296:4303] = '{32'hc2a1b7f3, 32'h418f7d03, 32'hc292eb86, 32'h42bb9337, 32'hc2b32cde, 32'hc290e450, 32'h428aa00b, 32'hc197f937};
test_output[4296:4303] = '{32'h0, 32'h418f7d03, 32'h0, 32'h42bb9337, 32'h0, 32'h0, 32'h428aa00b, 32'h0};
test_input[4304:4311] = '{32'h40f9d897, 32'hc2596804, 32'hc24feed7, 32'hc0ae4cca, 32'hc239a066, 32'h429f21e2, 32'hc2735ce4, 32'h40c4a56f};
test_output[4304:4311] = '{32'h40f9d897, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429f21e2, 32'h0, 32'h40c4a56f};
test_input[4312:4319] = '{32'hc1b6083e, 32'h42aa8070, 32'h421fec6e, 32'h4253c1bc, 32'hc28871a4, 32'h424d180a, 32'h42231f04, 32'hc25db14b};
test_output[4312:4319] = '{32'h0, 32'h42aa8070, 32'h421fec6e, 32'h4253c1bc, 32'h0, 32'h424d180a, 32'h42231f04, 32'h0};
test_input[4320:4327] = '{32'h428958a8, 32'h42aec522, 32'h423d74d0, 32'hc2555676, 32'h428f0af4, 32'hc25bcab2, 32'h40973467, 32'hc267483d};
test_output[4320:4327] = '{32'h428958a8, 32'h42aec522, 32'h423d74d0, 32'h0, 32'h428f0af4, 32'h0, 32'h40973467, 32'h0};
test_input[4328:4335] = '{32'hc21650ab, 32'hc0b7924d, 32'h42985b57, 32'hc1f7a8cb, 32'hc28fee97, 32'h41987ff0, 32'h42c4dcec, 32'hc1be3e62};
test_output[4328:4335] = '{32'h0, 32'h0, 32'h42985b57, 32'h0, 32'h0, 32'h41987ff0, 32'h42c4dcec, 32'h0};
test_input[4336:4343] = '{32'h42a513e0, 32'h42b401f5, 32'h429c1e40, 32'h428c1e77, 32'h4193d93c, 32'h42a8ea2a, 32'hc29cffd0, 32'h42b9d7e9};
test_output[4336:4343] = '{32'h42a513e0, 32'h42b401f5, 32'h429c1e40, 32'h428c1e77, 32'h4193d93c, 32'h42a8ea2a, 32'h0, 32'h42b9d7e9};
test_input[4344:4351] = '{32'h4277614e, 32'hc245fc93, 32'hc2174f1b, 32'hc2391c12, 32'hc27580ee, 32'h4250c963, 32'h426d5b2e, 32'h41f4c22c};
test_output[4344:4351] = '{32'h4277614e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4250c963, 32'h426d5b2e, 32'h41f4c22c};
test_input[4352:4359] = '{32'hc11047b2, 32'h42c6b383, 32'h42379024, 32'h42bc7124, 32'h418d4f67, 32'h417d6a29, 32'hc252ec13, 32'hc16a1f19};
test_output[4352:4359] = '{32'h0, 32'h42c6b383, 32'h42379024, 32'h42bc7124, 32'h418d4f67, 32'h417d6a29, 32'h0, 32'h0};
test_input[4360:4367] = '{32'h41a65e6e, 32'h42671771, 32'h42541676, 32'h42bd0b30, 32'h42a401e4, 32'h420caff3, 32'hc28eb4b3, 32'hc23b21d8};
test_output[4360:4367] = '{32'h41a65e6e, 32'h42671771, 32'h42541676, 32'h42bd0b30, 32'h42a401e4, 32'h420caff3, 32'h0, 32'h0};
test_input[4368:4375] = '{32'h42bfa7a1, 32'h42271685, 32'hc293dd7e, 32'h42711a83, 32'hc2c3d20d, 32'hc286a2a6, 32'hc2a5bf73, 32'hc20b7f0b};
test_output[4368:4375] = '{32'h42bfa7a1, 32'h42271685, 32'h0, 32'h42711a83, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4376:4383] = '{32'hc2c0ef0e, 32'hc179b834, 32'h3f1f36a6, 32'hc27723df, 32'hc249ed60, 32'h42b25e28, 32'h4123f50b, 32'hc2279ad5};
test_output[4376:4383] = '{32'h0, 32'h0, 32'h3f1f36a6, 32'h0, 32'h0, 32'h42b25e28, 32'h4123f50b, 32'h0};
test_input[4384:4391] = '{32'h4283b71f, 32'h4299d060, 32'hc27c8217, 32'h42c70864, 32'h4266b46c, 32'hc20859f2, 32'hc2a9450a, 32'h4172de94};
test_output[4384:4391] = '{32'h4283b71f, 32'h4299d060, 32'h0, 32'h42c70864, 32'h4266b46c, 32'h0, 32'h0, 32'h4172de94};
test_input[4392:4399] = '{32'h418fa1dd, 32'h42915cde, 32'h429ff4ba, 32'hc2a6f017, 32'h42617fb6, 32'hc27422d4, 32'h421f4c19, 32'hc2a49073};
test_output[4392:4399] = '{32'h418fa1dd, 32'h42915cde, 32'h429ff4ba, 32'h0, 32'h42617fb6, 32'h0, 32'h421f4c19, 32'h0};
test_input[4400:4407] = '{32'hc0ac0262, 32'h41bf0c99, 32'hc2295724, 32'h41699976, 32'h427fd2ee, 32'h429ea331, 32'hc17a08df, 32'h429bc975};
test_output[4400:4407] = '{32'h0, 32'h41bf0c99, 32'h0, 32'h41699976, 32'h427fd2ee, 32'h429ea331, 32'h0, 32'h429bc975};
test_input[4408:4415] = '{32'hc2b691ed, 32'h41a1c51b, 32'h424e4a68, 32'h4273f480, 32'hc18e9bde, 32'hc2286cb5, 32'h41e1dace, 32'h42c52db0};
test_output[4408:4415] = '{32'h0, 32'h41a1c51b, 32'h424e4a68, 32'h4273f480, 32'h0, 32'h0, 32'h41e1dace, 32'h42c52db0};
test_input[4416:4423] = '{32'hc2a123a2, 32'hc025b45d, 32'hc173f4ec, 32'hc13b93a1, 32'h42505a18, 32'hc26bd173, 32'h42b041c0, 32'h42392e38};
test_output[4416:4423] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42505a18, 32'h0, 32'h42b041c0, 32'h42392e38};
test_input[4424:4431] = '{32'h42850fc1, 32'h420bb356, 32'hc29d0976, 32'hc20998d3, 32'hc1c8e7c5, 32'hc1ab79c7, 32'hc23e1542, 32'hc2c78896};
test_output[4424:4431] = '{32'h42850fc1, 32'h420bb356, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4432:4439] = '{32'hc2be5c1d, 32'hc2743a2a, 32'hc28b6c61, 32'h42687652, 32'hc17cfdf2, 32'h4201cc26, 32'hc29a7ac6, 32'h41fcbf32};
test_output[4432:4439] = '{32'h0, 32'h0, 32'h0, 32'h42687652, 32'h0, 32'h4201cc26, 32'h0, 32'h41fcbf32};
test_input[4440:4447] = '{32'h41d207ce, 32'hc10ac124, 32'hc2a474e8, 32'hc042bf4d, 32'h4255a28a, 32'h3fa64e40, 32'h42b39f8e, 32'h4281d018};
test_output[4440:4447] = '{32'h41d207ce, 32'h0, 32'h0, 32'h0, 32'h4255a28a, 32'h3fa64e40, 32'h42b39f8e, 32'h4281d018};
test_input[4448:4455] = '{32'hc1c741d6, 32'h40661801, 32'h426d4621, 32'h4212c52c, 32'h42010030, 32'h414e4dd6, 32'hc1851259, 32'h41db7f52};
test_output[4448:4455] = '{32'h0, 32'h40661801, 32'h426d4621, 32'h4212c52c, 32'h42010030, 32'h414e4dd6, 32'h0, 32'h41db7f52};
test_input[4456:4463] = '{32'hc1db79c9, 32'hc2b74eea, 32'hc28fdd7b, 32'h42ba5b8c, 32'hc2873cab, 32'hc23ab882, 32'hc22971a5, 32'hc2c5db55};
test_output[4456:4463] = '{32'h0, 32'h0, 32'h0, 32'h42ba5b8c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4464:4471] = '{32'hc1c65041, 32'hc28d8e99, 32'h428a3527, 32'hc2478fdb, 32'hc1fbb5ff, 32'h42af91c0, 32'h42a666b9, 32'hc28bf660};
test_output[4464:4471] = '{32'h0, 32'h0, 32'h428a3527, 32'h0, 32'h0, 32'h42af91c0, 32'h42a666b9, 32'h0};
test_input[4472:4479] = '{32'h4245d868, 32'hc1bc102e, 32'h42a14983, 32'h42c2cae6, 32'h42ad6525, 32'h40fa45ab, 32'hc235f821, 32'h420bc366};
test_output[4472:4479] = '{32'h4245d868, 32'h0, 32'h42a14983, 32'h42c2cae6, 32'h42ad6525, 32'h40fa45ab, 32'h0, 32'h420bc366};
test_input[4480:4487] = '{32'h4234abff, 32'h422e3bab, 32'h3f238362, 32'hbfb09df5, 32'hc0aa44de, 32'h41777589, 32'h42988b64, 32'h41300355};
test_output[4480:4487] = '{32'h4234abff, 32'h422e3bab, 32'h3f238362, 32'h0, 32'h0, 32'h41777589, 32'h42988b64, 32'h41300355};
test_input[4488:4495] = '{32'h41eeaf0d, 32'h415e5271, 32'hc13ad00c, 32'h42b8ad52, 32'h3fd7abbb, 32'h42783662, 32'hc101aceb, 32'hc22d19bb};
test_output[4488:4495] = '{32'h41eeaf0d, 32'h415e5271, 32'h0, 32'h42b8ad52, 32'h3fd7abbb, 32'h42783662, 32'h0, 32'h0};
test_input[4496:4503] = '{32'h42bba806, 32'hc2313fb4, 32'h4298ab92, 32'h422b0b53, 32'hc2c6de67, 32'hc2534bfc, 32'hc2c721ce, 32'h4160c53d};
test_output[4496:4503] = '{32'h42bba806, 32'h0, 32'h4298ab92, 32'h422b0b53, 32'h0, 32'h0, 32'h0, 32'h4160c53d};
test_input[4504:4511] = '{32'hc2b19759, 32'h426a3177, 32'hc0e7c937, 32'hc2890e67, 32'hc232886b, 32'hc24a25b2, 32'h42c459f7, 32'h42563bc1};
test_output[4504:4511] = '{32'h0, 32'h426a3177, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c459f7, 32'h42563bc1};
test_input[4512:4519] = '{32'h41a0575e, 32'h411b7e52, 32'hc10f5371, 32'h4293efd5, 32'hc2884d37, 32'hc200cda1, 32'hc2bdb58c, 32'h42ba6b5c};
test_output[4512:4519] = '{32'h41a0575e, 32'h411b7e52, 32'h0, 32'h4293efd5, 32'h0, 32'h0, 32'h0, 32'h42ba6b5c};
test_input[4520:4527] = '{32'hc2c279df, 32'h4209302b, 32'hc2812ecb, 32'h4236b25b, 32'hc06f3b94, 32'h41de804e, 32'h42b198a9, 32'hc036771f};
test_output[4520:4527] = '{32'h0, 32'h4209302b, 32'h0, 32'h4236b25b, 32'h0, 32'h41de804e, 32'h42b198a9, 32'h0};
test_input[4528:4535] = '{32'hc1e2219f, 32'h41a1cff8, 32'h42acb60e, 32'h415979aa, 32'hbfd9bf2b, 32'h424bae13, 32'hc2863c78, 32'hc21b1c87};
test_output[4528:4535] = '{32'h0, 32'h41a1cff8, 32'h42acb60e, 32'h415979aa, 32'h0, 32'h424bae13, 32'h0, 32'h0};
test_input[4536:4543] = '{32'h41842690, 32'hc0f3a989, 32'hc27aa7cc, 32'h41a30d12, 32'hc24eac46, 32'h403e2c4a, 32'h41e77904, 32'hc1a28038};
test_output[4536:4543] = '{32'h41842690, 32'h0, 32'h0, 32'h41a30d12, 32'h0, 32'h403e2c4a, 32'h41e77904, 32'h0};
test_input[4544:4551] = '{32'hc1910e04, 32'h429c1ae0, 32'h42464116, 32'h42405cc9, 32'h42b3f1dd, 32'hc2c23f12, 32'hc25f7daf, 32'hc29dfd6d};
test_output[4544:4551] = '{32'h0, 32'h429c1ae0, 32'h42464116, 32'h42405cc9, 32'h42b3f1dd, 32'h0, 32'h0, 32'h0};
test_input[4552:4559] = '{32'hc293a4f9, 32'h422cb01c, 32'hc2ac9fb1, 32'h4238509c, 32'hc295cf67, 32'h41f229b4, 32'hc2142f04, 32'h42368f0f};
test_output[4552:4559] = '{32'h0, 32'h422cb01c, 32'h0, 32'h4238509c, 32'h0, 32'h41f229b4, 32'h0, 32'h42368f0f};
test_input[4560:4567] = '{32'hc2071a65, 32'h4187f942, 32'h42ac8c4f, 32'h3ed93838, 32'h41aeaddd, 32'h42a1b184, 32'h40a3bf46, 32'h420ea157};
test_output[4560:4567] = '{32'h0, 32'h4187f942, 32'h42ac8c4f, 32'h3ed93838, 32'h41aeaddd, 32'h42a1b184, 32'h40a3bf46, 32'h420ea157};
test_input[4568:4575] = '{32'h42bc9dd8, 32'hc2683270, 32'hc2c55c95, 32'h41cc5735, 32'h4105d842, 32'hc2aaa7d5, 32'hc0f18e9c, 32'hc27af673};
test_output[4568:4575] = '{32'h42bc9dd8, 32'h0, 32'h0, 32'h41cc5735, 32'h4105d842, 32'h0, 32'h0, 32'h0};
test_input[4576:4583] = '{32'h417c5c59, 32'hc2a4a33a, 32'h42b908c9, 32'hc2ad9ab7, 32'hc2c0836a, 32'h41d0cf4b, 32'h402f7efe, 32'h42630755};
test_output[4576:4583] = '{32'h417c5c59, 32'h0, 32'h42b908c9, 32'h0, 32'h0, 32'h41d0cf4b, 32'h402f7efe, 32'h42630755};
test_input[4584:4591] = '{32'h42c32627, 32'h428bea95, 32'hc2708b21, 32'hc29828e0, 32'hc24beef7, 32'hc2bb005d, 32'hc26a3fb4, 32'h41f95dc2};
test_output[4584:4591] = '{32'h42c32627, 32'h428bea95, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f95dc2};
test_input[4592:4599] = '{32'h419f75ce, 32'h4273b5ca, 32'h42acb552, 32'h41205fc3, 32'h4254d80c, 32'h42b7fc30, 32'hc26a85cb, 32'h42a167da};
test_output[4592:4599] = '{32'h419f75ce, 32'h4273b5ca, 32'h42acb552, 32'h41205fc3, 32'h4254d80c, 32'h42b7fc30, 32'h0, 32'h42a167da};
test_input[4600:4607] = '{32'hc280e949, 32'hc27fad65, 32'h42a7d75d, 32'h42b64432, 32'h4210873c, 32'hc268e094, 32'h412dbaa3, 32'hc21ef3dd};
test_output[4600:4607] = '{32'h0, 32'h0, 32'h42a7d75d, 32'h42b64432, 32'h4210873c, 32'h0, 32'h412dbaa3, 32'h0};
test_input[4608:4615] = '{32'h423a31ce, 32'hc28dd052, 32'h418d7ac7, 32'h41517a04, 32'hc26f2c39, 32'h42abc6f2, 32'hc0c7ee34, 32'hc207789b};
test_output[4608:4615] = '{32'h423a31ce, 32'h0, 32'h418d7ac7, 32'h41517a04, 32'h0, 32'h42abc6f2, 32'h0, 32'h0};
test_input[4616:4623] = '{32'h41eb95bb, 32'h42430408, 32'hc2a2212b, 32'hc2bf42cc, 32'h41b1d53a, 32'h429cfaae, 32'hc2bacdfe, 32'hc209be2a};
test_output[4616:4623] = '{32'h41eb95bb, 32'h42430408, 32'h0, 32'h0, 32'h41b1d53a, 32'h429cfaae, 32'h0, 32'h0};
test_input[4624:4631] = '{32'hc24aabd7, 32'h41afeb57, 32'h41bf9f20, 32'h421b8156, 32'h42c66fa9, 32'h4264b0ae, 32'h42077132, 32'h428d0e2f};
test_output[4624:4631] = '{32'h0, 32'h41afeb57, 32'h41bf9f20, 32'h421b8156, 32'h42c66fa9, 32'h4264b0ae, 32'h42077132, 32'h428d0e2f};
test_input[4632:4639] = '{32'hc2bb2b70, 32'h42247eb7, 32'h41213a31, 32'h41908a47, 32'h421a0bb5, 32'h42a2100d, 32'hc210e74d, 32'hc27131e1};
test_output[4632:4639] = '{32'h0, 32'h42247eb7, 32'h41213a31, 32'h41908a47, 32'h421a0bb5, 32'h42a2100d, 32'h0, 32'h0};
test_input[4640:4647] = '{32'hc24e122d, 32'h42afbd78, 32'h42959ac1, 32'h425d5ee9, 32'h40bb4d38, 32'h42aa473d, 32'h424af912, 32'hbea3054b};
test_output[4640:4647] = '{32'h0, 32'h42afbd78, 32'h42959ac1, 32'h425d5ee9, 32'h40bb4d38, 32'h42aa473d, 32'h424af912, 32'h0};
test_input[4648:4655] = '{32'hc258690c, 32'h41ee9025, 32'h4282a016, 32'hc28f21ed, 32'hc263413e, 32'hc1af485a, 32'hc1c24c4c, 32'hc1c14583};
test_output[4648:4655] = '{32'h0, 32'h41ee9025, 32'h4282a016, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4656:4663] = '{32'hc2bdee74, 32'h42abc5e2, 32'h42bf377c, 32'h416cc5f7, 32'h42b7291b, 32'h4040bc23, 32'h4257034e, 32'h4214a0b1};
test_output[4656:4663] = '{32'h0, 32'h42abc5e2, 32'h42bf377c, 32'h416cc5f7, 32'h42b7291b, 32'h4040bc23, 32'h4257034e, 32'h4214a0b1};
test_input[4664:4671] = '{32'hc06e0c2b, 32'hc2074125, 32'h40ace0dc, 32'h42c25689, 32'hc2864c5e, 32'h42a9d25b, 32'h42b344f2, 32'hc23923a5};
test_output[4664:4671] = '{32'h0, 32'h0, 32'h40ace0dc, 32'h42c25689, 32'h0, 32'h42a9d25b, 32'h42b344f2, 32'h0};
test_input[4672:4679] = '{32'h428a014d, 32'h428971f7, 32'h42934940, 32'h420265c2, 32'hc1a7baff, 32'hc1b8c2fb, 32'hc22e28e1, 32'h42808ef8};
test_output[4672:4679] = '{32'h428a014d, 32'h428971f7, 32'h42934940, 32'h420265c2, 32'h0, 32'h0, 32'h0, 32'h42808ef8};
test_input[4680:4687] = '{32'hc20b920b, 32'h42435add, 32'hc2b93d09, 32'h4145bb5b, 32'hc224f6d1, 32'hc219bc0a, 32'hc1ba87df, 32'hc1507586};
test_output[4680:4687] = '{32'h0, 32'h42435add, 32'h0, 32'h4145bb5b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4688:4695] = '{32'hc2925740, 32'hc2a1e00c, 32'hc2bea093, 32'hc2a09494, 32'hc285e87c, 32'h424a2b96, 32'hc09ce5c7, 32'hc10fe796};
test_output[4688:4695] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h424a2b96, 32'h0, 32'h0};
test_input[4696:4703] = '{32'h4284c8fb, 32'hc0b0ab5e, 32'h422a329a, 32'hc272fa78, 32'h421ddff4, 32'hc2b3a2d8, 32'hc2336070, 32'h42860714};
test_output[4696:4703] = '{32'h4284c8fb, 32'h0, 32'h422a329a, 32'h0, 32'h421ddff4, 32'h0, 32'h0, 32'h42860714};
test_input[4704:4711] = '{32'h3f51ce0c, 32'hc2c4bd76, 32'hc27fa182, 32'h4182d51e, 32'h42b5352a, 32'h40ab530b, 32'hc12e8e39, 32'hc29cba89};
test_output[4704:4711] = '{32'h3f51ce0c, 32'h0, 32'h0, 32'h4182d51e, 32'h42b5352a, 32'h40ab530b, 32'h0, 32'h0};
test_input[4712:4719] = '{32'h42222055, 32'hc0ca9783, 32'hc2b2e762, 32'h4268984b, 32'hc1959cae, 32'h40f00a30, 32'h40bfc843, 32'hc2a5c851};
test_output[4712:4719] = '{32'h42222055, 32'h0, 32'h0, 32'h4268984b, 32'h0, 32'h40f00a30, 32'h40bfc843, 32'h0};
test_input[4720:4727] = '{32'hbfc0a98e, 32'hc0a3b107, 32'hc2652082, 32'h42ab79e8, 32'hc1ca7367, 32'h4244d122, 32'hc28052b8, 32'hc0ce88ec};
test_output[4720:4727] = '{32'h0, 32'h0, 32'h0, 32'h42ab79e8, 32'h0, 32'h4244d122, 32'h0, 32'h0};
test_input[4728:4735] = '{32'h4214e57d, 32'hc25f8009, 32'h42a07a60, 32'hc1ada4a6, 32'h41b0b617, 32'h427f11d7, 32'hc21fbd1f, 32'hc26b640a};
test_output[4728:4735] = '{32'h4214e57d, 32'h0, 32'h42a07a60, 32'h0, 32'h41b0b617, 32'h427f11d7, 32'h0, 32'h0};
test_input[4736:4743] = '{32'hc2720db2, 32'h42b0b824, 32'h424aeed0, 32'hc2910c91, 32'h41ab31a8, 32'h42b8d567, 32'hc2241fe0, 32'hc2b4cefe};
test_output[4736:4743] = '{32'h0, 32'h42b0b824, 32'h424aeed0, 32'h0, 32'h41ab31a8, 32'h42b8d567, 32'h0, 32'h0};
test_input[4744:4751] = '{32'h42c2ebec, 32'hc2c6e0f8, 32'hc2b1d26c, 32'h426eff70, 32'hc222c78e, 32'hc27db920, 32'h4182ecae, 32'hc2632140};
test_output[4744:4751] = '{32'h42c2ebec, 32'h0, 32'h0, 32'h426eff70, 32'h0, 32'h0, 32'h4182ecae, 32'h0};
test_input[4752:4759] = '{32'hc1b77de6, 32'h41e65e86, 32'h421e1888, 32'hc26cdc79, 32'hc2341adc, 32'h42c6d76e, 32'hc2b1e136, 32'hc1c37e2e};
test_output[4752:4759] = '{32'h0, 32'h41e65e86, 32'h421e1888, 32'h0, 32'h0, 32'h42c6d76e, 32'h0, 32'h0};
test_input[4760:4767] = '{32'h3c96b341, 32'hc222f132, 32'h4234eab3, 32'hc2963ca4, 32'h428b824e, 32'h42b501c3, 32'hc2813329, 32'hc2859f6b};
test_output[4760:4767] = '{32'h3c96b341, 32'h0, 32'h4234eab3, 32'h0, 32'h428b824e, 32'h42b501c3, 32'h0, 32'h0};
test_input[4768:4775] = '{32'hc2a7a824, 32'h42bfc4fd, 32'h429f1ee9, 32'h4216f003, 32'hc248753b, 32'h42897b45, 32'h41417fe4, 32'hc29cee78};
test_output[4768:4775] = '{32'h0, 32'h42bfc4fd, 32'h429f1ee9, 32'h4216f003, 32'h0, 32'h42897b45, 32'h41417fe4, 32'h0};
test_input[4776:4783] = '{32'h41bb0a93, 32'h41c8f93f, 32'hc281010c, 32'hc2aa0744, 32'hc12cdaa7, 32'hc27446d3, 32'h4166f27f, 32'hc29e3593};
test_output[4776:4783] = '{32'h41bb0a93, 32'h41c8f93f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4166f27f, 32'h0};
test_input[4784:4791] = '{32'hc2c52f4f, 32'hc2843fb1, 32'h41e6f76d, 32'h4293418c, 32'hc1a61163, 32'h420afd8a, 32'h4221ea1e, 32'h417df6f8};
test_output[4784:4791] = '{32'h0, 32'h0, 32'h41e6f76d, 32'h4293418c, 32'h0, 32'h420afd8a, 32'h4221ea1e, 32'h417df6f8};
test_input[4792:4799] = '{32'hc10146c8, 32'hc20e6bae, 32'h4281197f, 32'h4206c346, 32'h4292188c, 32'hc21b039e, 32'h42c6d705, 32'h41807d2c};
test_output[4792:4799] = '{32'h0, 32'h0, 32'h4281197f, 32'h4206c346, 32'h4292188c, 32'h0, 32'h42c6d705, 32'h41807d2c};
test_input[4800:4807] = '{32'hc2856df9, 32'hc22948be, 32'h4232642d, 32'h40436c0e, 32'h42871c95, 32'hbf5b3fe6, 32'hc20e03e0, 32'hc140c35a};
test_output[4800:4807] = '{32'h0, 32'h0, 32'h4232642d, 32'h40436c0e, 32'h42871c95, 32'h0, 32'h0, 32'h0};
test_input[4808:4815] = '{32'h424dfec5, 32'hc2a42f50, 32'hc27cc14a, 32'hc288301b, 32'h402f6b2c, 32'hc0716ab3, 32'hc071fbc5, 32'h429862e7};
test_output[4808:4815] = '{32'h424dfec5, 32'h0, 32'h0, 32'h0, 32'h402f6b2c, 32'h0, 32'h0, 32'h429862e7};
test_input[4816:4823] = '{32'h42a9d633, 32'h41ce656f, 32'hc2bf6ad3, 32'h42958121, 32'h41d3199d, 32'hc26526ca, 32'h42110169, 32'hc27c66b9};
test_output[4816:4823] = '{32'h42a9d633, 32'h41ce656f, 32'h0, 32'h42958121, 32'h41d3199d, 32'h0, 32'h42110169, 32'h0};
test_input[4824:4831] = '{32'hc0d154a6, 32'hbfa7961d, 32'h410a584b, 32'hc0fd458b, 32'hc1878101, 32'hc1a636de, 32'h40c43734, 32'hc2a74a62};
test_output[4824:4831] = '{32'h0, 32'h0, 32'h410a584b, 32'h0, 32'h0, 32'h0, 32'h40c43734, 32'h0};
test_input[4832:4839] = '{32'h42830f50, 32'hc2be0295, 32'hc2aab50c, 32'h41a539aa, 32'h42b36e81, 32'hc201ed78, 32'h407a9b03, 32'hc2a7f6b7};
test_output[4832:4839] = '{32'h42830f50, 32'h0, 32'h0, 32'h41a539aa, 32'h42b36e81, 32'h0, 32'h407a9b03, 32'h0};
test_input[4840:4847] = '{32'hc2a9b266, 32'hc2360542, 32'hc2a0435d, 32'hc2817e37, 32'hc26d3066, 32'h42966bf0, 32'hc1b281cd, 32'hc2c7ff34};
test_output[4840:4847] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42966bf0, 32'h0, 32'h0};
test_input[4848:4855] = '{32'hc29eec5c, 32'h42b3be8b, 32'h40b265e1, 32'h429af1d4, 32'h41c5cbb8, 32'hc25141fa, 32'hc150c534, 32'hc1e7eb21};
test_output[4848:4855] = '{32'h0, 32'h42b3be8b, 32'h40b265e1, 32'h429af1d4, 32'h41c5cbb8, 32'h0, 32'h0, 32'h0};
test_input[4856:4863] = '{32'hc2aa97a7, 32'hc2199249, 32'hc210a458, 32'h42aaee16, 32'hc272b0f9, 32'hc26842d8, 32'h42ab6ad2, 32'h4258cfd9};
test_output[4856:4863] = '{32'h0, 32'h0, 32'h0, 32'h42aaee16, 32'h0, 32'h0, 32'h42ab6ad2, 32'h4258cfd9};
test_input[4864:4871] = '{32'h42c33305, 32'hc18a1e01, 32'hc1a24a22, 32'hc2ace0fe, 32'h41e4dee3, 32'h4294ca54, 32'h41c33513, 32'hc244e3e6};
test_output[4864:4871] = '{32'h42c33305, 32'h0, 32'h0, 32'h0, 32'h41e4dee3, 32'h4294ca54, 32'h41c33513, 32'h0};
test_input[4872:4879] = '{32'hc2357e9a, 32'h4263815b, 32'h427e2a7c, 32'hc1b8cb49, 32'h42308698, 32'h4186bc52, 32'hc175f95b, 32'hc25d9789};
test_output[4872:4879] = '{32'h0, 32'h4263815b, 32'h427e2a7c, 32'h0, 32'h42308698, 32'h4186bc52, 32'h0, 32'h0};
test_input[4880:4887] = '{32'hc28a77fc, 32'h424444ef, 32'hc1c70321, 32'h4261b572, 32'hc2c7ea01, 32'h42b5f080, 32'h42a289c9, 32'h3fa94442};
test_output[4880:4887] = '{32'h0, 32'h424444ef, 32'h0, 32'h4261b572, 32'h0, 32'h42b5f080, 32'h42a289c9, 32'h3fa94442};
test_input[4888:4895] = '{32'h423b3d73, 32'h42a11681, 32'h4286a0b0, 32'h4282b1e0, 32'h426cc460, 32'hc27901f3, 32'hc1c6f452, 32'h4204bcfa};
test_output[4888:4895] = '{32'h423b3d73, 32'h42a11681, 32'h4286a0b0, 32'h4282b1e0, 32'h426cc460, 32'h0, 32'h0, 32'h4204bcfa};
test_input[4896:4903] = '{32'h40682ffe, 32'hc049083f, 32'h429fa2f0, 32'hc22c4948, 32'h42c77719, 32'hc25c73db, 32'h42c62b62, 32'h40963f78};
test_output[4896:4903] = '{32'h40682ffe, 32'h0, 32'h429fa2f0, 32'h0, 32'h42c77719, 32'h0, 32'h42c62b62, 32'h40963f78};
test_input[4904:4911] = '{32'hc23b3de8, 32'hc1ff3257, 32'hc28f9d6b, 32'h42a6dafb, 32'h428a67ab, 32'hc25e4bf9, 32'h42c3863e, 32'hc2bdbc89};
test_output[4904:4911] = '{32'h0, 32'h0, 32'h0, 32'h42a6dafb, 32'h428a67ab, 32'h0, 32'h42c3863e, 32'h0};
test_input[4912:4919] = '{32'h42b5833a, 32'hc22deddc, 32'hc2c6ca15, 32'h42778e11, 32'hc178e26f, 32'h424b0505, 32'h422c03a1, 32'h42528a93};
test_output[4912:4919] = '{32'h42b5833a, 32'h0, 32'h0, 32'h42778e11, 32'h0, 32'h424b0505, 32'h422c03a1, 32'h42528a93};
test_input[4920:4927] = '{32'hc1db36db, 32'hc1ed4313, 32'hc10ac079, 32'hc21c9ce6, 32'hc24e4c3f, 32'h41dc0b85, 32'hc23c1b04, 32'hc2a8b2d7};
test_output[4920:4927] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41dc0b85, 32'h0, 32'h0};
test_input[4928:4935] = '{32'h418b4bc9, 32'h42a82319, 32'h3fa9bb19, 32'h4295f6a3, 32'hc1f00cce, 32'h418a44c5, 32'hc28b9676, 32'h428926d5};
test_output[4928:4935] = '{32'h418b4bc9, 32'h42a82319, 32'h3fa9bb19, 32'h4295f6a3, 32'h0, 32'h418a44c5, 32'h0, 32'h428926d5};
test_input[4936:4943] = '{32'h42144f33, 32'hc1c13bf3, 32'hc21536e0, 32'h4234ffe0, 32'hc2580779, 32'hc2152518, 32'h415fe714, 32'hc13c0e85};
test_output[4936:4943] = '{32'h42144f33, 32'h0, 32'h0, 32'h4234ffe0, 32'h0, 32'h0, 32'h415fe714, 32'h0};
test_input[4944:4951] = '{32'hbf888ae9, 32'hc2977b0a, 32'h418932a2, 32'h40ac6713, 32'hc22d0abb, 32'h42a8bb77, 32'h41e635ab, 32'h42b1f5c7};
test_output[4944:4951] = '{32'h0, 32'h0, 32'h418932a2, 32'h40ac6713, 32'h0, 32'h42a8bb77, 32'h41e635ab, 32'h42b1f5c7};
test_input[4952:4959] = '{32'h42184a7d, 32'hc208561e, 32'hc23f7d62, 32'hc1c90ecc, 32'h42b1f491, 32'h427678da, 32'hc29b21c9, 32'h42a8b5e1};
test_output[4952:4959] = '{32'h42184a7d, 32'h0, 32'h0, 32'h0, 32'h42b1f491, 32'h427678da, 32'h0, 32'h42a8b5e1};
test_input[4960:4967] = '{32'hc235755c, 32'h4293c88d, 32'hc289b10a, 32'hc2a197e0, 32'hc1747681, 32'h41dd9a0f, 32'h42c393de, 32'h41efbaa7};
test_output[4960:4967] = '{32'h0, 32'h4293c88d, 32'h0, 32'h0, 32'h0, 32'h41dd9a0f, 32'h42c393de, 32'h41efbaa7};
test_input[4968:4975] = '{32'h41be7503, 32'hc241a499, 32'h42a6e44e, 32'hc1ee15ee, 32'h419131af, 32'h42a40715, 32'h412f2816, 32'h41a97025};
test_output[4968:4975] = '{32'h41be7503, 32'h0, 32'h42a6e44e, 32'h0, 32'h419131af, 32'h42a40715, 32'h412f2816, 32'h41a97025};
test_input[4976:4983] = '{32'hc2c736e4, 32'hc2464a47, 32'hc2ab9ddc, 32'hc254ef01, 32'hc1cc7cb4, 32'h42382f51, 32'h41b5bf5c, 32'h4238dd77};
test_output[4976:4983] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42382f51, 32'h41b5bf5c, 32'h4238dd77};
test_input[4984:4991] = '{32'hc13f3bd0, 32'h418c458f, 32'hc2bf022c, 32'h42918d26, 32'hc29a0287, 32'hc25f7490, 32'h42895ecf, 32'hc016d5c8};
test_output[4984:4991] = '{32'h0, 32'h418c458f, 32'h0, 32'h42918d26, 32'h0, 32'h0, 32'h42895ecf, 32'h0};
test_input[4992:4999] = '{32'h429a2c29, 32'h42c49fe1, 32'h42a4c07a, 32'hc1855b36, 32'h418642fb, 32'h41fbed70, 32'hc21d816a, 32'h420d59d9};
test_output[4992:4999] = '{32'h429a2c29, 32'h42c49fe1, 32'h42a4c07a, 32'h0, 32'h418642fb, 32'h41fbed70, 32'h0, 32'h420d59d9};
test_input[5000:5007] = '{32'hc22d86c4, 32'hc0e6cd18, 32'hc20f1d59, 32'hc1845c05, 32'h42a60b6f, 32'hc207ac7e, 32'h42024982, 32'hc2a4f4fe};
test_output[5000:5007] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a60b6f, 32'h0, 32'h42024982, 32'h0};
test_input[5008:5015] = '{32'hc219b3f2, 32'hc22a672b, 32'hc216ba86, 32'hc10a4b5a, 32'hc2b99a57, 32'h41acd2b6, 32'hc2575835, 32'hc2bf984c};
test_output[5008:5015] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41acd2b6, 32'h0, 32'h0};
test_input[5016:5023] = '{32'h4203956f, 32'hc2ab6642, 32'hc242b344, 32'h4280f008, 32'hc24bd18a, 32'h429ecfdd, 32'hbdfe10f4, 32'h42882568};
test_output[5016:5023] = '{32'h4203956f, 32'h0, 32'h0, 32'h4280f008, 32'h0, 32'h429ecfdd, 32'h0, 32'h42882568};
test_input[5024:5031] = '{32'hc24ef596, 32'hc2c008f6, 32'hc194a62f, 32'h422422fc, 32'h422c77b3, 32'h42060fb9, 32'hbf94c71b, 32'hc2868843};
test_output[5024:5031] = '{32'h0, 32'h0, 32'h0, 32'h422422fc, 32'h422c77b3, 32'h42060fb9, 32'h0, 32'h0};
test_input[5032:5039] = '{32'hc271e330, 32'hc2b1601a, 32'hbe7e4e01, 32'hc270513d, 32'hc2140358, 32'h4162219a, 32'h4299b33e, 32'hbff31997};
test_output[5032:5039] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4162219a, 32'h4299b33e, 32'h0};
test_input[5040:5047] = '{32'h428089cf, 32'hc27586c8, 32'hc2984f3c, 32'h4167dfb6, 32'hc2abeabd, 32'hc09455b3, 32'h40046ac2, 32'h42c765d9};
test_output[5040:5047] = '{32'h428089cf, 32'h0, 32'h0, 32'h4167dfb6, 32'h0, 32'h0, 32'h40046ac2, 32'h42c765d9};
test_input[5048:5055] = '{32'hc2abbc41, 32'hc291ba68, 32'h428287d8, 32'h428e93d2, 32'hc2b07897, 32'h4285d0c2, 32'hc1720f29, 32'h42a5033a};
test_output[5048:5055] = '{32'h0, 32'h0, 32'h428287d8, 32'h428e93d2, 32'h0, 32'h4285d0c2, 32'h0, 32'h42a5033a};
test_input[5056:5063] = '{32'h4196e957, 32'hc0742564, 32'hc2a91f28, 32'hc2a012c6, 32'h4298d89c, 32'h41ed48aa, 32'h42bdc8cc, 32'h4162c1e2};
test_output[5056:5063] = '{32'h4196e957, 32'h0, 32'h0, 32'h0, 32'h4298d89c, 32'h41ed48aa, 32'h42bdc8cc, 32'h4162c1e2};
test_input[5064:5071] = '{32'hc129619f, 32'hc12eaece, 32'h3f474109, 32'h429395bf, 32'hc0627635, 32'hc29fd7ba, 32'h42bd083f, 32'hc29e3ea6};
test_output[5064:5071] = '{32'h0, 32'h0, 32'h3f474109, 32'h429395bf, 32'h0, 32'h0, 32'h42bd083f, 32'h0};
test_input[5072:5079] = '{32'hc29a851d, 32'hc28460f9, 32'h421e7d26, 32'hc19f10c2, 32'hc21fd97b, 32'hc0a7fa78, 32'hc228351e, 32'h3f792518};
test_output[5072:5079] = '{32'h0, 32'h0, 32'h421e7d26, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3f792518};
test_input[5080:5087] = '{32'h41d363a5, 32'hc10635b1, 32'h42c3cdf0, 32'hc02a003d, 32'h4108bff3, 32'hc1894ce4, 32'h40653c7d, 32'h4260cd51};
test_output[5080:5087] = '{32'h41d363a5, 32'h0, 32'h42c3cdf0, 32'h0, 32'h4108bff3, 32'h0, 32'h40653c7d, 32'h4260cd51};
test_input[5088:5095] = '{32'hc1d11ed2, 32'h42995814, 32'hc21d2a69, 32'hc27dd59d, 32'hc2c2553e, 32'hc2590b04, 32'h42c7edc3, 32'hc2bdd117};
test_output[5088:5095] = '{32'h0, 32'h42995814, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c7edc3, 32'h0};
test_input[5096:5103] = '{32'h426cccf9, 32'h42c04743, 32'hc28a68fc, 32'hc2a35f17, 32'hc250f53c, 32'h42b30fde, 32'hc14c21dd, 32'hc0e56e41};
test_output[5096:5103] = '{32'h426cccf9, 32'h42c04743, 32'h0, 32'h0, 32'h0, 32'h42b30fde, 32'h0, 32'h0};
test_input[5104:5111] = '{32'hc2b5a22b, 32'hc2ba565c, 32'hc21ce3ad, 32'hc25b6bd5, 32'hc2399241, 32'h42c73ee6, 32'hc17d930f, 32'h40774dad};
test_output[5104:5111] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c73ee6, 32'h0, 32'h40774dad};
test_input[5112:5119] = '{32'hc2b15320, 32'hc2b8670f, 32'h41b8c767, 32'hc20caa1f, 32'hc26ebc95, 32'h41a462ce, 32'hc26fc5cd, 32'h421fc51f};
test_output[5112:5119] = '{32'h0, 32'h0, 32'h41b8c767, 32'h0, 32'h0, 32'h41a462ce, 32'h0, 32'h421fc51f};
test_input[5120:5127] = '{32'h421e23b4, 32'hc2a28bb2, 32'hc2c076cf, 32'hc223cea9, 32'hc273c078, 32'hc1220640, 32'hc1e9080d, 32'hc1babc9f};
test_output[5120:5127] = '{32'h421e23b4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5128:5135] = '{32'h4238b44b, 32'h41511dc3, 32'h418b9911, 32'h41f06bc9, 32'h428ea3c7, 32'hc1b43b65, 32'h41d3ac31, 32'h4235fd8e};
test_output[5128:5135] = '{32'h4238b44b, 32'h41511dc3, 32'h418b9911, 32'h41f06bc9, 32'h428ea3c7, 32'h0, 32'h41d3ac31, 32'h4235fd8e};
test_input[5136:5143] = '{32'h4235ea2c, 32'h42c6c805, 32'hc28d788c, 32'h424445a5, 32'hc23c242e, 32'hc25c6720, 32'h42a1df2b, 32'hc199b3e3};
test_output[5136:5143] = '{32'h4235ea2c, 32'h42c6c805, 32'h0, 32'h424445a5, 32'h0, 32'h0, 32'h42a1df2b, 32'h0};
test_input[5144:5151] = '{32'h42c72b4c, 32'h42ac760c, 32'hc227bde3, 32'h425481c9, 32'hc024d59b, 32'hc2c2cc9a, 32'h426f7376, 32'hc1ba62c3};
test_output[5144:5151] = '{32'h42c72b4c, 32'h42ac760c, 32'h0, 32'h425481c9, 32'h0, 32'h0, 32'h426f7376, 32'h0};
test_input[5152:5159] = '{32'h42b5f40b, 32'hc25a4927, 32'h4246a9b7, 32'h42909c9a, 32'h42a4d3cf, 32'h42c56c14, 32'hc1b78797, 32'hc29ed177};
test_output[5152:5159] = '{32'h42b5f40b, 32'h0, 32'h4246a9b7, 32'h42909c9a, 32'h42a4d3cf, 32'h42c56c14, 32'h0, 32'h0};
test_input[5160:5167] = '{32'h42b672c1, 32'h42a3dee7, 32'hc1460d46, 32'h42a7cff5, 32'hc29a38d5, 32'hc2bb8111, 32'hc1041f31, 32'hc2990d9f};
test_output[5160:5167] = '{32'h42b672c1, 32'h42a3dee7, 32'h0, 32'h42a7cff5, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5168:5175] = '{32'hc20c5bb6, 32'hc204f78b, 32'h40e9faf1, 32'h42582ce1, 32'h42571be0, 32'hc1047e93, 32'hc252f4d8, 32'hc2917766};
test_output[5168:5175] = '{32'h0, 32'h0, 32'h40e9faf1, 32'h42582ce1, 32'h42571be0, 32'h0, 32'h0, 32'h0};
test_input[5176:5183] = '{32'h41e0e0ae, 32'h41e34984, 32'h41970f9b, 32'hc2555f3b, 32'h423be1ca, 32'hc297ec28, 32'h421c8987, 32'h4295c2e4};
test_output[5176:5183] = '{32'h41e0e0ae, 32'h41e34984, 32'h41970f9b, 32'h0, 32'h423be1ca, 32'h0, 32'h421c8987, 32'h4295c2e4};
test_input[5184:5191] = '{32'h42a5285c, 32'hc00d10e3, 32'hc228167e, 32'hc29af7af, 32'h4231170e, 32'hc208ad4b, 32'h42584184, 32'hc28a4e96};
test_output[5184:5191] = '{32'h42a5285c, 32'h0, 32'h0, 32'h0, 32'h4231170e, 32'h0, 32'h42584184, 32'h0};
test_input[5192:5199] = '{32'hc240eeb0, 32'h425ef140, 32'hc2c46348, 32'hc2936f5d, 32'h41e2b270, 32'h42640ff0, 32'h42b643bc, 32'hc0fe55d2};
test_output[5192:5199] = '{32'h0, 32'h425ef140, 32'h0, 32'h0, 32'h41e2b270, 32'h42640ff0, 32'h42b643bc, 32'h0};
test_input[5200:5207] = '{32'hc2058436, 32'hc253d5aa, 32'hc2151e99, 32'hc0f9f996, 32'hc299b1e1, 32'h42bf26cc, 32'h425703c1, 32'h4278b276};
test_output[5200:5207] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bf26cc, 32'h425703c1, 32'h4278b276};
test_input[5208:5215] = '{32'h41e11451, 32'h421b6ac4, 32'h41a38da6, 32'hc27a1cfe, 32'h42ae18a5, 32'h42931b08, 32'hc25f16cf, 32'hc28d7466};
test_output[5208:5215] = '{32'h41e11451, 32'h421b6ac4, 32'h41a38da6, 32'h0, 32'h42ae18a5, 32'h42931b08, 32'h0, 32'h0};
test_input[5216:5223] = '{32'h42a591f7, 32'h4269993d, 32'hc2a9d45a, 32'h42701a9e, 32'h423a60e6, 32'h42355f98, 32'hc067b6fd, 32'hc1ee8736};
test_output[5216:5223] = '{32'h42a591f7, 32'h4269993d, 32'h0, 32'h42701a9e, 32'h423a60e6, 32'h42355f98, 32'h0, 32'h0};
test_input[5224:5231] = '{32'h422d1a51, 32'h41a5ca45, 32'hbf0bb461, 32'hc2bcb60a, 32'hc2861a86, 32'hc24cec5e, 32'h42302690, 32'hc2a3c9cf};
test_output[5224:5231] = '{32'h422d1a51, 32'h41a5ca45, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42302690, 32'h0};
test_input[5232:5239] = '{32'hc2767747, 32'h426d4e50, 32'h42c46374, 32'hc2ad2280, 32'hc1c93d53, 32'h4256e8bc, 32'h41fc4921, 32'h42552422};
test_output[5232:5239] = '{32'h0, 32'h426d4e50, 32'h42c46374, 32'h0, 32'h0, 32'h4256e8bc, 32'h41fc4921, 32'h42552422};
test_input[5240:5247] = '{32'h41f7b0d7, 32'hbf214fb0, 32'h42996a01, 32'h425e678b, 32'h406653ce, 32'hc2865239, 32'h423d499a, 32'hc13b3280};
test_output[5240:5247] = '{32'h41f7b0d7, 32'h0, 32'h42996a01, 32'h425e678b, 32'h406653ce, 32'h0, 32'h423d499a, 32'h0};
test_input[5248:5255] = '{32'h42a981a4, 32'hc2529024, 32'h41e3e66a, 32'hc27c1947, 32'hc1260b93, 32'h3d89744e, 32'hc24addfe, 32'h42558eb2};
test_output[5248:5255] = '{32'h42a981a4, 32'h0, 32'h41e3e66a, 32'h0, 32'h0, 32'h3d89744e, 32'h0, 32'h42558eb2};
test_input[5256:5263] = '{32'hc24a0975, 32'h4109ed17, 32'hc25ab486, 32'h409d957c, 32'h428c4599, 32'h42925496, 32'hc29c18a1, 32'hc219c75c};
test_output[5256:5263] = '{32'h0, 32'h4109ed17, 32'h0, 32'h409d957c, 32'h428c4599, 32'h42925496, 32'h0, 32'h0};
test_input[5264:5271] = '{32'h4247ea9f, 32'h41e65999, 32'hc2707191, 32'h42a685d8, 32'hc1cbddc9, 32'hc11cdaa9, 32'hc256b3c4, 32'h415e3d09};
test_output[5264:5271] = '{32'h4247ea9f, 32'h41e65999, 32'h0, 32'h42a685d8, 32'h0, 32'h0, 32'h0, 32'h415e3d09};
test_input[5272:5279] = '{32'h4216c350, 32'hc2b8ff01, 32'h422ff1bf, 32'hc26c91eb, 32'hc245765d, 32'h42a390d0, 32'hc2381cdc, 32'hc291e8ff};
test_output[5272:5279] = '{32'h4216c350, 32'h0, 32'h422ff1bf, 32'h0, 32'h0, 32'h42a390d0, 32'h0, 32'h0};
test_input[5280:5287] = '{32'hc2b271b3, 32'hc2b105e8, 32'hc2be5d06, 32'h42befe8b, 32'h4270319a, 32'hc2ad3d55, 32'hc231efae, 32'h422293a9};
test_output[5280:5287] = '{32'h0, 32'h0, 32'h0, 32'h42befe8b, 32'h4270319a, 32'h0, 32'h0, 32'h422293a9};
test_input[5288:5295] = '{32'hc0b3c92f, 32'hc2a10542, 32'h416832a2, 32'hc287d57b, 32'hc2c3b7b8, 32'hc1a1933a, 32'hc14cb182, 32'hc1c58c6f};
test_output[5288:5295] = '{32'h0, 32'h0, 32'h416832a2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5296:5303] = '{32'hc2a12eee, 32'h423593e4, 32'h42631050, 32'h42816aad, 32'h41fe7d42, 32'h42a61856, 32'hc1dca6a1, 32'hc2a94a5f};
test_output[5296:5303] = '{32'h0, 32'h423593e4, 32'h42631050, 32'h42816aad, 32'h41fe7d42, 32'h42a61856, 32'h0, 32'h0};
test_input[5304:5311] = '{32'h42bc95ec, 32'h426b9c1d, 32'hc2a7307c, 32'h42661ce2, 32'h4262c840, 32'hc2b4095e, 32'h41ebea5f, 32'hc29c59dd};
test_output[5304:5311] = '{32'h42bc95ec, 32'h426b9c1d, 32'h0, 32'h42661ce2, 32'h4262c840, 32'h0, 32'h41ebea5f, 32'h0};
test_input[5312:5319] = '{32'hc2a41150, 32'h4289be1e, 32'hc28ebdbf, 32'hc293f376, 32'hc294331f, 32'h428dd56b, 32'h42a50265, 32'h413b39ff};
test_output[5312:5319] = '{32'h0, 32'h4289be1e, 32'h0, 32'h0, 32'h0, 32'h428dd56b, 32'h42a50265, 32'h413b39ff};
test_input[5320:5327] = '{32'h427febc2, 32'h4201538d, 32'h42c4bd46, 32'h42b385b6, 32'h42a77768, 32'h41e1d07c, 32'hc1e3cd58, 32'hc24dcf36};
test_output[5320:5327] = '{32'h427febc2, 32'h4201538d, 32'h42c4bd46, 32'h42b385b6, 32'h42a77768, 32'h41e1d07c, 32'h0, 32'h0};
test_input[5328:5335] = '{32'hc16ef21e, 32'h420b599a, 32'hc1311629, 32'h4220fb48, 32'hc19fc41a, 32'h4231402d, 32'h42b92099, 32'h42838220};
test_output[5328:5335] = '{32'h0, 32'h420b599a, 32'h0, 32'h4220fb48, 32'h0, 32'h4231402d, 32'h42b92099, 32'h42838220};
test_input[5336:5343] = '{32'h407a0b21, 32'hc1a3fe91, 32'h42ba19b5, 32'hc1a55a77, 32'h429d7e7b, 32'hc28ac864, 32'h4249e599, 32'hc18203f9};
test_output[5336:5343] = '{32'h407a0b21, 32'h0, 32'h42ba19b5, 32'h0, 32'h429d7e7b, 32'h0, 32'h4249e599, 32'h0};
test_input[5344:5351] = '{32'hc28767d1, 32'h42ad4278, 32'h42821372, 32'h40aeb4c3, 32'h429f0799, 32'hc2639bcc, 32'h421ef9ae, 32'h4115abad};
test_output[5344:5351] = '{32'h0, 32'h42ad4278, 32'h42821372, 32'h40aeb4c3, 32'h429f0799, 32'h0, 32'h421ef9ae, 32'h4115abad};
test_input[5352:5359] = '{32'hc0be7a1b, 32'hc0b9fd12, 32'hc24adc18, 32'hc28f23a5, 32'hc253eb70, 32'hc2be3fc8, 32'h429113a3, 32'h3f6696c8};
test_output[5352:5359] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429113a3, 32'h3f6696c8};
test_input[5360:5367] = '{32'hc28d378d, 32'hc2927fb1, 32'hbe95ef31, 32'h42a5f38f, 32'hc2918b8c, 32'hc0b3cedd, 32'h4217c936, 32'hc1b4983a};
test_output[5360:5367] = '{32'h0, 32'h0, 32'h0, 32'h42a5f38f, 32'h0, 32'h0, 32'h4217c936, 32'h0};
test_input[5368:5375] = '{32'hc102b722, 32'hc1405b51, 32'h42a78bf1, 32'h423c9ca6, 32'h42b520a8, 32'hc1ec179d, 32'h429df37b, 32'hc2b47793};
test_output[5368:5375] = '{32'h0, 32'h0, 32'h42a78bf1, 32'h423c9ca6, 32'h42b520a8, 32'h0, 32'h429df37b, 32'h0};
test_input[5376:5383] = '{32'hc2057dbd, 32'hc29fc2f0, 32'h423caf6f, 32'hc24c3fcc, 32'hc288869e, 32'hc02b0af5, 32'h42c1ec99, 32'hc2bdd29a};
test_output[5376:5383] = '{32'h0, 32'h0, 32'h423caf6f, 32'h0, 32'h0, 32'h0, 32'h42c1ec99, 32'h0};
test_input[5384:5391] = '{32'hc23524b3, 32'hc259cf4e, 32'hbf20cd29, 32'hc2a55f37, 32'h4162fdcc, 32'hc205490d, 32'h413afa5f, 32'hc2c2cb26};
test_output[5384:5391] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4162fdcc, 32'h0, 32'h413afa5f, 32'h0};
test_input[5392:5399] = '{32'h429f9cbb, 32'h41ab5a60, 32'hc2baf248, 32'h42446939, 32'hc293c067, 32'h41dd2fc9, 32'h4206922c, 32'hc2129714};
test_output[5392:5399] = '{32'h429f9cbb, 32'h41ab5a60, 32'h0, 32'h42446939, 32'h0, 32'h41dd2fc9, 32'h4206922c, 32'h0};
test_input[5400:5407] = '{32'hc0395e9d, 32'hc29e944f, 32'h41ff768f, 32'h41841319, 32'hc28896e9, 32'hc1f76cf5, 32'hc2a52902, 32'hc0a8f2e4};
test_output[5400:5407] = '{32'h0, 32'h0, 32'h41ff768f, 32'h41841319, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5408:5415] = '{32'hc199c9fe, 32'h42c0b5a8, 32'h420fa55c, 32'hc2c60f24, 32'hc110d07f, 32'h4270ca57, 32'h4207cefd, 32'hc2a3401d};
test_output[5408:5415] = '{32'h0, 32'h42c0b5a8, 32'h420fa55c, 32'h0, 32'h0, 32'h4270ca57, 32'h4207cefd, 32'h0};
test_input[5416:5423] = '{32'h42570518, 32'h4225d2c9, 32'h4287631c, 32'hc22b44e0, 32'hc230351f, 32'hc273ee47, 32'hc2835875, 32'h425ab008};
test_output[5416:5423] = '{32'h42570518, 32'h4225d2c9, 32'h4287631c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425ab008};
test_input[5424:5431] = '{32'hc1cd0ab7, 32'hc092267f, 32'hc0e4546e, 32'h4229ef5f, 32'h428aaf1d, 32'hc2ac3d1d, 32'h409f39f9, 32'h42743b81};
test_output[5424:5431] = '{32'h0, 32'h0, 32'h0, 32'h4229ef5f, 32'h428aaf1d, 32'h0, 32'h409f39f9, 32'h42743b81};
test_input[5432:5439] = '{32'h41c8f48f, 32'h41b7f90c, 32'hc2c67638, 32'hc186a556, 32'h4261c3d1, 32'hc29fcb03, 32'h4171d100, 32'hc20e8822};
test_output[5432:5439] = '{32'h41c8f48f, 32'h41b7f90c, 32'h0, 32'h0, 32'h4261c3d1, 32'h0, 32'h4171d100, 32'h0};
test_input[5440:5447] = '{32'h42ba5563, 32'h42876271, 32'hc28dfe0a, 32'hc170355e, 32'hc258d250, 32'hc080129b, 32'h3eead0ca, 32'h42a694dd};
test_output[5440:5447] = '{32'h42ba5563, 32'h42876271, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3eead0ca, 32'h42a694dd};
test_input[5448:5455] = '{32'hc159c56c, 32'hc15193e9, 32'hc2201f92, 32'hc08b3468, 32'hc226767b, 32'hc1e7d34b, 32'h41fe2918, 32'hc228b4e1};
test_output[5448:5455] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41fe2918, 32'h0};
test_input[5456:5463] = '{32'hc146a6de, 32'h4213e77b, 32'h4084a834, 32'h411199bc, 32'h427dad6b, 32'hc2ae0307, 32'hc259816b, 32'h420b2513};
test_output[5456:5463] = '{32'h0, 32'h4213e77b, 32'h4084a834, 32'h411199bc, 32'h427dad6b, 32'h0, 32'h0, 32'h420b2513};
test_input[5464:5471] = '{32'h42c56407, 32'hc225cb5c, 32'h428f4aa2, 32'h420472a8, 32'h42864808, 32'hc2c326a0, 32'hc29d7d23, 32'hc1a14b3d};
test_output[5464:5471] = '{32'h42c56407, 32'h0, 32'h428f4aa2, 32'h420472a8, 32'h42864808, 32'h0, 32'h0, 32'h0};
test_input[5472:5479] = '{32'hc0e6cf1e, 32'h422a700d, 32'hc114e156, 32'hc2c47a2d, 32'h409afe8d, 32'h42773d20, 32'hc10b0e36, 32'h42aa2e87};
test_output[5472:5479] = '{32'h0, 32'h422a700d, 32'h0, 32'h0, 32'h409afe8d, 32'h42773d20, 32'h0, 32'h42aa2e87};
test_input[5480:5487] = '{32'h41945805, 32'h427cbc00, 32'hc20bc7e6, 32'h426556ae, 32'hc294923e, 32'h42aa6e7d, 32'h42556a3f, 32'hc16df275};
test_output[5480:5487] = '{32'h41945805, 32'h427cbc00, 32'h0, 32'h426556ae, 32'h0, 32'h42aa6e7d, 32'h42556a3f, 32'h0};
test_input[5488:5495] = '{32'hc13cb4d8, 32'hc28917ad, 32'h426ad033, 32'h428072e6, 32'h428ca140, 32'hc27c1399, 32'h42a197ef, 32'hc2111cf0};
test_output[5488:5495] = '{32'h0, 32'h0, 32'h426ad033, 32'h428072e6, 32'h428ca140, 32'h0, 32'h42a197ef, 32'h0};
test_input[5496:5503] = '{32'h41cbaa05, 32'h421e6a83, 32'h42c71eb2, 32'h426c8d7a, 32'h42879ebe, 32'h429d1a7e, 32'hc1a07199, 32'h400f21a1};
test_output[5496:5503] = '{32'h41cbaa05, 32'h421e6a83, 32'h42c71eb2, 32'h426c8d7a, 32'h42879ebe, 32'h429d1a7e, 32'h0, 32'h400f21a1};
test_input[5504:5511] = '{32'h4215f7bc, 32'hc2c6c47e, 32'h40daf572, 32'hc267adb4, 32'hc243bfe0, 32'h418fbf7f, 32'h404f1515, 32'hc1a045d7};
test_output[5504:5511] = '{32'h4215f7bc, 32'h0, 32'h40daf572, 32'h0, 32'h0, 32'h418fbf7f, 32'h404f1515, 32'h0};
test_input[5512:5519] = '{32'h4251f8cb, 32'h42043bde, 32'h41ecf696, 32'hc1192590, 32'hc2c4b781, 32'hc29374de, 32'h42ba5324, 32'h4298ab42};
test_output[5512:5519] = '{32'h4251f8cb, 32'h42043bde, 32'h41ecf696, 32'h0, 32'h0, 32'h0, 32'h42ba5324, 32'h4298ab42};
test_input[5520:5527] = '{32'h421781a7, 32'h4222bf2f, 32'hc25ba141, 32'hc1fa04c8, 32'h41f2acea, 32'h42a50758, 32'hc28bb3bb, 32'hc2bc14c8};
test_output[5520:5527] = '{32'h421781a7, 32'h4222bf2f, 32'h0, 32'h0, 32'h41f2acea, 32'h42a50758, 32'h0, 32'h0};
test_input[5528:5535] = '{32'h428880ae, 32'h428f2a71, 32'hc236f93b, 32'hc2af7675, 32'hc273b40e, 32'h4259314f, 32'hc2b1dd30, 32'hc0958a50};
test_output[5528:5535] = '{32'h428880ae, 32'h428f2a71, 32'h0, 32'h0, 32'h0, 32'h4259314f, 32'h0, 32'h0};
test_input[5536:5543] = '{32'h419dfee8, 32'h42b3105d, 32'hc2aacb63, 32'hc15de4d6, 32'hc22602c1, 32'h42335942, 32'hc2a58bf4, 32'h428667b8};
test_output[5536:5543] = '{32'h419dfee8, 32'h42b3105d, 32'h0, 32'h0, 32'h0, 32'h42335942, 32'h0, 32'h428667b8};
test_input[5544:5551] = '{32'h41fe06b2, 32'hc27eeb38, 32'hc20c302f, 32'h429b42f6, 32'hc2c0ba17, 32'h42b8edef, 32'hc29ffc79, 32'h428b1092};
test_output[5544:5551] = '{32'h41fe06b2, 32'h0, 32'h0, 32'h429b42f6, 32'h0, 32'h42b8edef, 32'h0, 32'h428b1092};
test_input[5552:5559] = '{32'h4239599c, 32'h42694a4e, 32'hc2a77682, 32'hc2ab4e97, 32'h42a7206e, 32'hc2c7663f, 32'h424c6294, 32'hc19d18ec};
test_output[5552:5559] = '{32'h4239599c, 32'h42694a4e, 32'h0, 32'h0, 32'h42a7206e, 32'h0, 32'h424c6294, 32'h0};
test_input[5560:5567] = '{32'h4213cadf, 32'hc20fd9fd, 32'hc285602d, 32'hc206ed88, 32'hc2b73f2e, 32'hc21e778a, 32'h42349deb, 32'hc1f9d4d5};
test_output[5560:5567] = '{32'h4213cadf, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42349deb, 32'h0};
test_input[5568:5575] = '{32'h4299c648, 32'h4221889d, 32'h41e14c87, 32'h4286aa53, 32'hc2b57466, 32'hc1a70434, 32'hc263314a, 32'h424e12e6};
test_output[5568:5575] = '{32'h4299c648, 32'h4221889d, 32'h41e14c87, 32'h4286aa53, 32'h0, 32'h0, 32'h0, 32'h424e12e6};
test_input[5576:5583] = '{32'h4290d659, 32'hc1b27f9a, 32'h42a6f5b2, 32'h423ab225, 32'h403ea6d4, 32'h4113f47a, 32'h41acd7a1, 32'hc2c4194a};
test_output[5576:5583] = '{32'h4290d659, 32'h0, 32'h42a6f5b2, 32'h423ab225, 32'h403ea6d4, 32'h4113f47a, 32'h41acd7a1, 32'h0};
test_input[5584:5591] = '{32'h41e183b7, 32'hc21163fa, 32'h4283e239, 32'hc28ced2b, 32'h422b4448, 32'h41c19ead, 32'hc2aaf656, 32'hc0c6ee45};
test_output[5584:5591] = '{32'h41e183b7, 32'h0, 32'h4283e239, 32'h0, 32'h422b4448, 32'h41c19ead, 32'h0, 32'h0};
test_input[5592:5599] = '{32'h42924bfc, 32'h42708780, 32'hc247b433, 32'h42b10a4b, 32'h42bdd6c4, 32'h423342f8, 32'hc23dd742, 32'h42b00c6e};
test_output[5592:5599] = '{32'h42924bfc, 32'h42708780, 32'h0, 32'h42b10a4b, 32'h42bdd6c4, 32'h423342f8, 32'h0, 32'h42b00c6e};
test_input[5600:5607] = '{32'hc2c0e04c, 32'hc28ed457, 32'h4035b92e, 32'h4299c1e2, 32'hc09a54c0, 32'h42984675, 32'h41dc51e3, 32'hbf10fe01};
test_output[5600:5607] = '{32'h0, 32'h0, 32'h4035b92e, 32'h4299c1e2, 32'h0, 32'h42984675, 32'h41dc51e3, 32'h0};
test_input[5608:5615] = '{32'hc23c3548, 32'h4126c71f, 32'h416a985f, 32'hc04eef09, 32'h427fe7ec, 32'h4231a533, 32'hc2be7ecc, 32'h42971cac};
test_output[5608:5615] = '{32'h0, 32'h4126c71f, 32'h416a985f, 32'h0, 32'h427fe7ec, 32'h4231a533, 32'h0, 32'h42971cac};
test_input[5616:5623] = '{32'hc27408d1, 32'hc2a31c18, 32'hc2ab9e00, 32'h42a36168, 32'h3fe2a61d, 32'hc294050a, 32'hc23de83a, 32'hc251a79d};
test_output[5616:5623] = '{32'h0, 32'h0, 32'h0, 32'h42a36168, 32'h3fe2a61d, 32'h0, 32'h0, 32'h0};
test_input[5624:5631] = '{32'h429aa82f, 32'h40435f93, 32'hc29337f4, 32'h42a7f143, 32'hc2925acd, 32'hc2c5ada8, 32'hc24c0d0a, 32'h411ea6db};
test_output[5624:5631] = '{32'h429aa82f, 32'h40435f93, 32'h0, 32'h42a7f143, 32'h0, 32'h0, 32'h0, 32'h411ea6db};
test_input[5632:5639] = '{32'hc2282b85, 32'h423b6a57, 32'h42896fd0, 32'h42930b70, 32'hc280ce33, 32'hc1198408, 32'hc2744d9f, 32'h42526f60};
test_output[5632:5639] = '{32'h0, 32'h423b6a57, 32'h42896fd0, 32'h42930b70, 32'h0, 32'h0, 32'h0, 32'h42526f60};
test_input[5640:5647] = '{32'h41e3fd6b, 32'hc15cbf19, 32'h4291737e, 32'h4283f397, 32'h42af4442, 32'hc295092f, 32'hc2370e8b, 32'hc1f357a1};
test_output[5640:5647] = '{32'h41e3fd6b, 32'h0, 32'h4291737e, 32'h4283f397, 32'h42af4442, 32'h0, 32'h0, 32'h0};
test_input[5648:5655] = '{32'h42b3d76e, 32'h425795d6, 32'hc23e1805, 32'h4189ff9d, 32'h409c9163, 32'hc2b6d457, 32'h42acba61, 32'h42a369bf};
test_output[5648:5655] = '{32'h42b3d76e, 32'h425795d6, 32'h0, 32'h4189ff9d, 32'h409c9163, 32'h0, 32'h42acba61, 32'h42a369bf};
test_input[5656:5663] = '{32'hc291adf7, 32'hc27ecec3, 32'hc0d94416, 32'h42942e6a, 32'h41dd0f1b, 32'hc235dfd6, 32'hc1f5df8b, 32'hc2798f9d};
test_output[5656:5663] = '{32'h0, 32'h0, 32'h0, 32'h42942e6a, 32'h41dd0f1b, 32'h0, 32'h0, 32'h0};
test_input[5664:5671] = '{32'hc28ff48e, 32'h41555e03, 32'h42673a1d, 32'hc236a5b9, 32'h42a9f272, 32'hc2ada368, 32'hc1cd053e, 32'h41e5de39};
test_output[5664:5671] = '{32'h0, 32'h41555e03, 32'h42673a1d, 32'h0, 32'h42a9f272, 32'h0, 32'h0, 32'h41e5de39};
test_input[5672:5679] = '{32'h4277e45b, 32'hc2bb39cc, 32'hc2340ed2, 32'hc2c33960, 32'h420ff362, 32'h4104aff5, 32'h429fc41c, 32'h421a00ac};
test_output[5672:5679] = '{32'h4277e45b, 32'h0, 32'h0, 32'h0, 32'h420ff362, 32'h4104aff5, 32'h429fc41c, 32'h421a00ac};
test_input[5680:5687] = '{32'hc200e62d, 32'hc21f2f4a, 32'hc2836cb3, 32'hc1a0a806, 32'h41b580ca, 32'h41af0f4d, 32'h42ad1a93, 32'h4285c82f};
test_output[5680:5687] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41b580ca, 32'h41af0f4d, 32'h42ad1a93, 32'h4285c82f};
test_input[5688:5695] = '{32'h42009951, 32'h428a1f24, 32'h429b09ce, 32'hc2891247, 32'hc2933a5a, 32'hc2c28cad, 32'hc2bdb668, 32'hc24cf5fe};
test_output[5688:5695] = '{32'h42009951, 32'h428a1f24, 32'h429b09ce, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5696:5703] = '{32'h4292cbd2, 32'hc2a5522f, 32'hc237242f, 32'hc2b778ae, 32'h42528bc2, 32'h41d384c1, 32'h40f316c8, 32'h42812b55};
test_output[5696:5703] = '{32'h4292cbd2, 32'h0, 32'h0, 32'h0, 32'h42528bc2, 32'h41d384c1, 32'h40f316c8, 32'h42812b55};
test_input[5704:5711] = '{32'hc215a04a, 32'hc2af5751, 32'h429561ab, 32'hc24aa7c3, 32'h422a99b3, 32'hc2aa1114, 32'h42b1dc0c, 32'h41b08c62};
test_output[5704:5711] = '{32'h0, 32'h0, 32'h429561ab, 32'h0, 32'h422a99b3, 32'h0, 32'h42b1dc0c, 32'h41b08c62};
test_input[5712:5719] = '{32'h4268337f, 32'hc2760afb, 32'hc2887036, 32'h426260c3, 32'hc124d81c, 32'h42059669, 32'hc297b8cc, 32'h411b4f0d};
test_output[5712:5719] = '{32'h4268337f, 32'h0, 32'h0, 32'h426260c3, 32'h0, 32'h42059669, 32'h0, 32'h411b4f0d};
test_input[5720:5727] = '{32'hc00e16b8, 32'hc2655e2e, 32'hc205fef2, 32'h408da062, 32'h428b0348, 32'h3f9a976f, 32'hc2270124, 32'hc23aab49};
test_output[5720:5727] = '{32'h0, 32'h0, 32'h0, 32'h408da062, 32'h428b0348, 32'h3f9a976f, 32'h0, 32'h0};
test_input[5728:5735] = '{32'h42befe26, 32'hc286223d, 32'h4295230b, 32'h415397e6, 32'h42b338a9, 32'hbf1614b7, 32'hc1b86e4f, 32'hc1d9ac1e};
test_output[5728:5735] = '{32'h42befe26, 32'h0, 32'h4295230b, 32'h415397e6, 32'h42b338a9, 32'h0, 32'h0, 32'h0};
test_input[5736:5743] = '{32'hc2b40fa8, 32'hc2bf006e, 32'h42909929, 32'hc2920546, 32'h420567cb, 32'h42129fd8, 32'h42255013, 32'h420f3a10};
test_output[5736:5743] = '{32'h0, 32'h0, 32'h42909929, 32'h0, 32'h420567cb, 32'h42129fd8, 32'h42255013, 32'h420f3a10};
test_input[5744:5751] = '{32'h42b60b15, 32'hc2c19d40, 32'h42191b3a, 32'hc2af71d0, 32'hc243e7c8, 32'hc275a307, 32'hc272cd5a, 32'h41f01cfc};
test_output[5744:5751] = '{32'h42b60b15, 32'h0, 32'h42191b3a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f01cfc};
test_input[5752:5759] = '{32'h428fbe6b, 32'hc241e3de, 32'h42c3f927, 32'h42b20f5d, 32'h41ea7b8b, 32'h42001683, 32'hc07d67e8, 32'hc22145a8};
test_output[5752:5759] = '{32'h428fbe6b, 32'h0, 32'h42c3f927, 32'h42b20f5d, 32'h41ea7b8b, 32'h42001683, 32'h0, 32'h0};
test_input[5760:5767] = '{32'hc286bd42, 32'h426c4a53, 32'h42847ab3, 32'hc0a1250c, 32'h4236cbc0, 32'h417d6dc0, 32'hc27e44e9, 32'hc265a32a};
test_output[5760:5767] = '{32'h0, 32'h426c4a53, 32'h42847ab3, 32'h0, 32'h4236cbc0, 32'h417d6dc0, 32'h0, 32'h0};
test_input[5768:5775] = '{32'h4210d45e, 32'hc2bf2d6c, 32'h428b67fc, 32'h42a85b15, 32'h40f4810e, 32'h40fc6795, 32'h42a36792, 32'hc2bea045};
test_output[5768:5775] = '{32'h4210d45e, 32'h0, 32'h428b67fc, 32'h42a85b15, 32'h40f4810e, 32'h40fc6795, 32'h42a36792, 32'h0};
test_input[5776:5783] = '{32'hc203272f, 32'hc2532970, 32'hc2c7128c, 32'h41e21c0c, 32'hc1bc1941, 32'h41aabaf9, 32'h4234e50d, 32'h41c9665d};
test_output[5776:5783] = '{32'h0, 32'h0, 32'h0, 32'h41e21c0c, 32'h0, 32'h41aabaf9, 32'h4234e50d, 32'h41c9665d};
test_input[5784:5791] = '{32'h42b7ed00, 32'h42b62822, 32'hc22158ad, 32'h41f5f3d0, 32'hc000637f, 32'hc1e37478, 32'hc2a83c95, 32'h41ad6ce7};
test_output[5784:5791] = '{32'h42b7ed00, 32'h42b62822, 32'h0, 32'h41f5f3d0, 32'h0, 32'h0, 32'h0, 32'h41ad6ce7};
test_input[5792:5799] = '{32'h411493b7, 32'h42034afe, 32'h4205b829, 32'hc18fe8fd, 32'h41ec0c04, 32'h42962953, 32'hc225e4ac, 32'hc225e6bf};
test_output[5792:5799] = '{32'h411493b7, 32'h42034afe, 32'h4205b829, 32'h0, 32'h41ec0c04, 32'h42962953, 32'h0, 32'h0};
test_input[5800:5807] = '{32'h41372ddb, 32'h419e5b32, 32'h422b8766, 32'h41686762, 32'h4184934f, 32'hc0db4513, 32'hc1c2ec6b, 32'hc20e638f};
test_output[5800:5807] = '{32'h41372ddb, 32'h419e5b32, 32'h422b8766, 32'h41686762, 32'h4184934f, 32'h0, 32'h0, 32'h0};
test_input[5808:5815] = '{32'h42afbcf7, 32'h42905f19, 32'h42c746f9, 32'hc2be319f, 32'hc2af1d44, 32'h42b4463b, 32'h425bc147, 32'hc2548b39};
test_output[5808:5815] = '{32'h42afbcf7, 32'h42905f19, 32'h42c746f9, 32'h0, 32'h0, 32'h42b4463b, 32'h425bc147, 32'h0};
test_input[5816:5823] = '{32'h428577d5, 32'hc2c64075, 32'hc2193838, 32'h41812353, 32'h427ace81, 32'hc1178b9b, 32'h41f91233, 32'hc29e6fa8};
test_output[5816:5823] = '{32'h428577d5, 32'h0, 32'h0, 32'h41812353, 32'h427ace81, 32'h0, 32'h41f91233, 32'h0};
test_input[5824:5831] = '{32'hc202e52e, 32'h4212d07f, 32'hc20ea476, 32'h42569722, 32'h418dae0f, 32'h41bf32d7, 32'h41c3bc6f, 32'h42bea587};
test_output[5824:5831] = '{32'h0, 32'h4212d07f, 32'h0, 32'h42569722, 32'h418dae0f, 32'h41bf32d7, 32'h41c3bc6f, 32'h42bea587};
test_input[5832:5839] = '{32'hc202675f, 32'h424ac288, 32'hc2b702a0, 32'hc22589c7, 32'hc2af01f0, 32'hc229780e, 32'hc0856e0d, 32'h41de8918};
test_output[5832:5839] = '{32'h0, 32'h424ac288, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41de8918};
test_input[5840:5847] = '{32'h42b5e667, 32'hc2be1ab1, 32'h42b9532f, 32'hc1344ff3, 32'hc2b7d679, 32'hc1166eff, 32'h41d4bfde, 32'h41bb0fa2};
test_output[5840:5847] = '{32'h42b5e667, 32'h0, 32'h42b9532f, 32'h0, 32'h0, 32'h0, 32'h41d4bfde, 32'h41bb0fa2};
test_input[5848:5855] = '{32'h41a88ab3, 32'hc28575f1, 32'h42943f3c, 32'h4108ca4e, 32'hc29d214d, 32'hc2b46693, 32'h409a5fb2, 32'h4170a861};
test_output[5848:5855] = '{32'h41a88ab3, 32'h0, 32'h42943f3c, 32'h4108ca4e, 32'h0, 32'h0, 32'h409a5fb2, 32'h4170a861};
test_input[5856:5863] = '{32'hc2a07b45, 32'h425b748a, 32'h427ba2eb, 32'hc0979993, 32'h415b63a7, 32'hc22429f5, 32'hc1859d93, 32'hc287e9b1};
test_output[5856:5863] = '{32'h0, 32'h425b748a, 32'h427ba2eb, 32'h0, 32'h415b63a7, 32'h0, 32'h0, 32'h0};
test_input[5864:5871] = '{32'h42bfbb6b, 32'h42a4012c, 32'hc2a37cea, 32'hc17e38fc, 32'h42c71e60, 32'hc2bc2725, 32'hc2bd3002, 32'hc1abefb2};
test_output[5864:5871] = '{32'h42bfbb6b, 32'h42a4012c, 32'h0, 32'h0, 32'h42c71e60, 32'h0, 32'h0, 32'h0};
test_input[5872:5879] = '{32'h42acd0fc, 32'hc21f574b, 32'hc1ad733f, 32'h42c34c73, 32'hc286b0a1, 32'h400cd046, 32'hc291efcc, 32'h42455b02};
test_output[5872:5879] = '{32'h42acd0fc, 32'h0, 32'h0, 32'h42c34c73, 32'h0, 32'h400cd046, 32'h0, 32'h42455b02};
test_input[5880:5887] = '{32'hc14b2249, 32'h425ad02f, 32'h41cd7acb, 32'h42a2ae67, 32'h4257637b, 32'h419f45b5, 32'hc1842f20, 32'h42a0be69};
test_output[5880:5887] = '{32'h0, 32'h425ad02f, 32'h41cd7acb, 32'h42a2ae67, 32'h4257637b, 32'h419f45b5, 32'h0, 32'h42a0be69};
test_input[5888:5895] = '{32'hc217c661, 32'hc2a6555e, 32'hc2b8aefd, 32'h42af8153, 32'hc2ba3775, 32'h428329f8, 32'hc20ee810, 32'h42633f31};
test_output[5888:5895] = '{32'h0, 32'h0, 32'h0, 32'h42af8153, 32'h0, 32'h428329f8, 32'h0, 32'h42633f31};
test_input[5896:5903] = '{32'hc163b4d6, 32'h41e3e16e, 32'hc2805179, 32'h422d264f, 32'h42186682, 32'hc1c1b5c5, 32'h41a351e6, 32'h4211f68b};
test_output[5896:5903] = '{32'h0, 32'h41e3e16e, 32'h0, 32'h422d264f, 32'h42186682, 32'h0, 32'h41a351e6, 32'h4211f68b};
test_input[5904:5911] = '{32'h42bac823, 32'hc2a3f92d, 32'hc2b37d62, 32'h42bfbfe8, 32'hc1827471, 32'h400faa09, 32'hc2bb0c51, 32'hc28510bb};
test_output[5904:5911] = '{32'h42bac823, 32'h0, 32'h0, 32'h42bfbfe8, 32'h0, 32'h400faa09, 32'h0, 32'h0};
test_input[5912:5919] = '{32'h42799fb7, 32'hc2362e8f, 32'h42446a7f, 32'h41387e11, 32'h42bb5309, 32'hc2a8f017, 32'h42a33a11, 32'h424090d9};
test_output[5912:5919] = '{32'h42799fb7, 32'h0, 32'h42446a7f, 32'h41387e11, 32'h42bb5309, 32'h0, 32'h42a33a11, 32'h424090d9};
test_input[5920:5927] = '{32'h41fbf7b6, 32'h42afbd61, 32'h4287b381, 32'h42893ac6, 32'h4185e55d, 32'h421f247a, 32'h429d8044, 32'h42ab676a};
test_output[5920:5927] = '{32'h41fbf7b6, 32'h42afbd61, 32'h4287b381, 32'h42893ac6, 32'h4185e55d, 32'h421f247a, 32'h429d8044, 32'h42ab676a};
test_input[5928:5935] = '{32'hc2aa1e65, 32'h41d196ef, 32'hc25ace92, 32'h41800946, 32'hc281d546, 32'hc1bfc89f, 32'h428ea4e9, 32'h42c3cb91};
test_output[5928:5935] = '{32'h0, 32'h41d196ef, 32'h0, 32'h41800946, 32'h0, 32'h0, 32'h428ea4e9, 32'h42c3cb91};
test_input[5936:5943] = '{32'hbfc0500f, 32'h42be9fb9, 32'h42291579, 32'hc1d3f6d8, 32'hc1df07d9, 32'h429141a5, 32'h421fdc22, 32'hc2b89528};
test_output[5936:5943] = '{32'h0, 32'h42be9fb9, 32'h42291579, 32'h0, 32'h0, 32'h429141a5, 32'h421fdc22, 32'h0};
test_input[5944:5951] = '{32'h429f556e, 32'hc2340e7f, 32'h42bf9646, 32'hc288fafc, 32'h429d44a6, 32'h423d2741, 32'h410fe6f8, 32'h40f840b8};
test_output[5944:5951] = '{32'h429f556e, 32'h0, 32'h42bf9646, 32'h0, 32'h429d44a6, 32'h423d2741, 32'h410fe6f8, 32'h40f840b8};
test_input[5952:5959] = '{32'hc1ea06b1, 32'hc21de2e7, 32'h405e2f20, 32'h41c428ff, 32'h426e8349, 32'hc2624552, 32'h42b8c4fb, 32'hc213557e};
test_output[5952:5959] = '{32'h0, 32'h0, 32'h405e2f20, 32'h41c428ff, 32'h426e8349, 32'h0, 32'h42b8c4fb, 32'h0};
test_input[5960:5967] = '{32'h41c2140a, 32'hc2946d78, 32'h41c3f140, 32'hc187f6c8, 32'hc298e6a6, 32'hc1c1c90f, 32'hc2c36052, 32'hc2a7635d};
test_output[5960:5967] = '{32'h41c2140a, 32'h0, 32'h41c3f140, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5968:5975] = '{32'h41cfd6ed, 32'hc1836d5a, 32'h425c7d98, 32'h424d6be7, 32'h4180ecf8, 32'h41253db1, 32'h421bea4c, 32'hc2c3838c};
test_output[5968:5975] = '{32'h41cfd6ed, 32'h0, 32'h425c7d98, 32'h424d6be7, 32'h4180ecf8, 32'h41253db1, 32'h421bea4c, 32'h0};
test_input[5976:5983] = '{32'hc24e1793, 32'hc246edbe, 32'h42a044f1, 32'h4186e556, 32'h420559d5, 32'hc25fc314, 32'h429f51bc, 32'h420220f8};
test_output[5976:5983] = '{32'h0, 32'h0, 32'h42a044f1, 32'h4186e556, 32'h420559d5, 32'h0, 32'h429f51bc, 32'h420220f8};
test_input[5984:5991] = '{32'hc2178b52, 32'hc239873d, 32'hc23ceb0e, 32'hc2bd4141, 32'h429dfe41, 32'hc2c2cfae, 32'h42c2e8b6, 32'hc29a3ced};
test_output[5984:5991] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429dfe41, 32'h0, 32'h42c2e8b6, 32'h0};
test_input[5992:5999] = '{32'hc1d5f30d, 32'hc0f370f0, 32'hc1d4f520, 32'h42a4bbe6, 32'h4260b356, 32'hc135e846, 32'hc27fec0e, 32'hc2ade11d};
test_output[5992:5999] = '{32'h0, 32'h0, 32'h0, 32'h42a4bbe6, 32'h4260b356, 32'h0, 32'h0, 32'h0};
test_input[6000:6007] = '{32'h428dba5b, 32'hc20548c7, 32'h42058eab, 32'h4110528a, 32'hc2728340, 32'h4149a85d, 32'h4169011e, 32'hc26d7e61};
test_output[6000:6007] = '{32'h428dba5b, 32'h0, 32'h42058eab, 32'h4110528a, 32'h0, 32'h4149a85d, 32'h4169011e, 32'h0};
test_input[6008:6015] = '{32'hc2a38514, 32'h42af70de, 32'hc0b15e68, 32'h408973a9, 32'hc205b81e, 32'h42be5681, 32'hc26258f3, 32'hc2ad6c4c};
test_output[6008:6015] = '{32'h0, 32'h42af70de, 32'h0, 32'h408973a9, 32'h0, 32'h42be5681, 32'h0, 32'h0};
test_input[6016:6023] = '{32'hc295f88f, 32'h429b0b31, 32'hc29d6419, 32'hc2038684, 32'h42a4a05c, 32'h4214d1ae, 32'h425e6d86, 32'hc0d2433b};
test_output[6016:6023] = '{32'h0, 32'h429b0b31, 32'h0, 32'h0, 32'h42a4a05c, 32'h4214d1ae, 32'h425e6d86, 32'h0};
test_input[6024:6031] = '{32'hc2b9d8da, 32'hc09413c0, 32'h4292b976, 32'hc02bcc9e, 32'h42c27feb, 32'h428df73e, 32'h41713c57, 32'hc042c0b2};
test_output[6024:6031] = '{32'h0, 32'h0, 32'h4292b976, 32'h0, 32'h42c27feb, 32'h428df73e, 32'h41713c57, 32'h0};
test_input[6032:6039] = '{32'h424211da, 32'hc1b3b4ee, 32'h4016a374, 32'hc1e1deb6, 32'hc1405db2, 32'hc14a2787, 32'h4212cd6d, 32'h40fd94c0};
test_output[6032:6039] = '{32'h424211da, 32'h0, 32'h4016a374, 32'h0, 32'h0, 32'h0, 32'h4212cd6d, 32'h40fd94c0};
test_input[6040:6047] = '{32'h42807a35, 32'h42a0ba17, 32'h41ee748c, 32'h428b9b6f, 32'h4048363f, 32'h42c0da1b, 32'hc28aa843, 32'hc240170a};
test_output[6040:6047] = '{32'h42807a35, 32'h42a0ba17, 32'h41ee748c, 32'h428b9b6f, 32'h4048363f, 32'h42c0da1b, 32'h0, 32'h0};
test_input[6048:6055] = '{32'h40abc629, 32'hc2339a83, 32'h42324076, 32'h42b33f28, 32'h4282af37, 32'h42b2a1c3, 32'hc216716e, 32'hc2842909};
test_output[6048:6055] = '{32'h40abc629, 32'h0, 32'h42324076, 32'h42b33f28, 32'h4282af37, 32'h42b2a1c3, 32'h0, 32'h0};
test_input[6056:6063] = '{32'hc297d33b, 32'hc2222bbb, 32'h42af7845, 32'h4252fefc, 32'hc21ba501, 32'h42223d50, 32'hc2a5e411, 32'h428c752d};
test_output[6056:6063] = '{32'h0, 32'h0, 32'h42af7845, 32'h4252fefc, 32'h0, 32'h42223d50, 32'h0, 32'h428c752d};
test_input[6064:6071] = '{32'hc28bb6a4, 32'hc1c40b30, 32'hc2a2585b, 32'hc233d8ae, 32'hc0f2df35, 32'h42450079, 32'h42c6f58d, 32'h4232fcb5};
test_output[6064:6071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42450079, 32'h42c6f58d, 32'h4232fcb5};
test_input[6072:6079] = '{32'hc1568135, 32'hc1c7fd95, 32'hc19695d9, 32'hc27795c6, 32'h424e0b68, 32'hc1cc2a16, 32'hc2a7e87b, 32'hc27d50a9};
test_output[6072:6079] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h424e0b68, 32'h0, 32'h0, 32'h0};
test_input[6080:6087] = '{32'hc2040753, 32'hc2589010, 32'hc28a6c5b, 32'hc239967b, 32'hc186c9b5, 32'h42b82683, 32'h422f9bd5, 32'h4179c518};
test_output[6080:6087] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b82683, 32'h422f9bd5, 32'h4179c518};
test_input[6088:6095] = '{32'h4274e173, 32'h4236ca14, 32'h42728cf5, 32'h4231ef0e, 32'h42b06200, 32'h4094d5be, 32'hc2938f47, 32'hc27a7dac};
test_output[6088:6095] = '{32'h4274e173, 32'h4236ca14, 32'h42728cf5, 32'h4231ef0e, 32'h42b06200, 32'h4094d5be, 32'h0, 32'h0};
test_input[6096:6103] = '{32'hc0748335, 32'h414f5756, 32'hc2b75be4, 32'h415cdf9f, 32'hc29ad13b, 32'h42a1fbfa, 32'hc1eed066, 32'hbfad143d};
test_output[6096:6103] = '{32'h0, 32'h414f5756, 32'h0, 32'h415cdf9f, 32'h0, 32'h42a1fbfa, 32'h0, 32'h0};
test_input[6104:6111] = '{32'h42a6a6b2, 32'h3f8346ba, 32'hc26fea4f, 32'h42309d0a, 32'hc227e3bf, 32'h42828b40, 32'hc27ea1f5, 32'h42a3ea7b};
test_output[6104:6111] = '{32'h42a6a6b2, 32'h3f8346ba, 32'h0, 32'h42309d0a, 32'h0, 32'h42828b40, 32'h0, 32'h42a3ea7b};
test_input[6112:6119] = '{32'hc203ac82, 32'h41097356, 32'h40960670, 32'hc168605b, 32'h424a52f6, 32'h425e5548, 32'hc23609c8, 32'h425b5b14};
test_output[6112:6119] = '{32'h0, 32'h41097356, 32'h40960670, 32'h0, 32'h424a52f6, 32'h425e5548, 32'h0, 32'h425b5b14};
test_input[6120:6127] = '{32'h41f19948, 32'hc26d3de8, 32'hc2889c0d, 32'h42449506, 32'h4222fd00, 32'h426e8001, 32'hc24bf02d, 32'hc1861370};
test_output[6120:6127] = '{32'h41f19948, 32'h0, 32'h0, 32'h42449506, 32'h4222fd00, 32'h426e8001, 32'h0, 32'h0};
test_input[6128:6135] = '{32'h4247f25e, 32'hc21908c3, 32'h42884df8, 32'hc25f1fb0, 32'h422823c8, 32'hc277b96f, 32'h42021734, 32'hc2b3d775};
test_output[6128:6135] = '{32'h4247f25e, 32'h0, 32'h42884df8, 32'h0, 32'h422823c8, 32'h0, 32'h42021734, 32'h0};
test_input[6136:6143] = '{32'hc2a981b9, 32'hc2778d26, 32'h4290f891, 32'h41bafe7a, 32'hc1b089b9, 32'h42bad6bc, 32'hc27f1916, 32'h42a0528d};
test_output[6136:6143] = '{32'h0, 32'h0, 32'h4290f891, 32'h41bafe7a, 32'h0, 32'h42bad6bc, 32'h0, 32'h42a0528d};
test_input[6144:6151] = '{32'h40ee5d2d, 32'hc2068079, 32'h414e6e1b, 32'h412a589c, 32'hc2ad6cc1, 32'h4148906d, 32'hc2642bce, 32'h4292957d};
test_output[6144:6151] = '{32'h40ee5d2d, 32'h0, 32'h414e6e1b, 32'h412a589c, 32'h0, 32'h4148906d, 32'h0, 32'h4292957d};
test_input[6152:6159] = '{32'hc29abc4f, 32'h42bff393, 32'hc297c7f5, 32'h427a3054, 32'h428e7be9, 32'h428e83a0, 32'h41d7b29c, 32'h41f78a11};
test_output[6152:6159] = '{32'h0, 32'h42bff393, 32'h0, 32'h427a3054, 32'h428e7be9, 32'h428e83a0, 32'h41d7b29c, 32'h41f78a11};
test_input[6160:6167] = '{32'h42c439c2, 32'h42c5573c, 32'h4296d8b9, 32'hc250b542, 32'hc1b570f2, 32'hc241eadf, 32'h42bc7140, 32'hc24fcd64};
test_output[6160:6167] = '{32'h42c439c2, 32'h42c5573c, 32'h4296d8b9, 32'h0, 32'h0, 32'h0, 32'h42bc7140, 32'h0};
test_input[6168:6175] = '{32'h41544f10, 32'h4249487d, 32'h41fbdfea, 32'hc24c21e6, 32'h41dfe103, 32'hc1d59f32, 32'h42c433bc, 32'hc1d0463b};
test_output[6168:6175] = '{32'h41544f10, 32'h4249487d, 32'h41fbdfea, 32'h0, 32'h41dfe103, 32'h0, 32'h42c433bc, 32'h0};
test_input[6176:6183] = '{32'hc1ba45dc, 32'h41735254, 32'hc179e189, 32'hc1ea6f77, 32'h428728cc, 32'h3eb436ef, 32'hc2bb1f04, 32'h41e3562c};
test_output[6176:6183] = '{32'h0, 32'h41735254, 32'h0, 32'h0, 32'h428728cc, 32'h3eb436ef, 32'h0, 32'h41e3562c};
test_input[6184:6191] = '{32'h42c362f4, 32'h42142ea0, 32'hc2bd25ba, 32'hc2a48687, 32'hc1bc2cbf, 32'h4201cae4, 32'h420b53ed, 32'hc18efba5};
test_output[6184:6191] = '{32'h42c362f4, 32'h42142ea0, 32'h0, 32'h0, 32'h0, 32'h4201cae4, 32'h420b53ed, 32'h0};
test_input[6192:6199] = '{32'hc253e598, 32'hc16fa5b5, 32'hc2a17395, 32'hc29490d4, 32'hc2a32dfb, 32'hc15bc9ca, 32'hc2852090, 32'hc2bf8ecd};
test_output[6192:6199] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6200:6207] = '{32'h42c26090, 32'hc254598a, 32'h41ffea08, 32'hc28cd9e6, 32'hc20938b0, 32'h4255a180, 32'h42c7382c, 32'h3e9ea0a5};
test_output[6200:6207] = '{32'h42c26090, 32'h0, 32'h41ffea08, 32'h0, 32'h0, 32'h4255a180, 32'h42c7382c, 32'h3e9ea0a5};
test_input[6208:6215] = '{32'h42073784, 32'h4047e271, 32'hc2a6209f, 32'hc1e6b5b7, 32'h42586811, 32'h428a0547, 32'hc292c092, 32'h42997c5f};
test_output[6208:6215] = '{32'h42073784, 32'h4047e271, 32'h0, 32'h0, 32'h42586811, 32'h428a0547, 32'h0, 32'h42997c5f};
test_input[6216:6223] = '{32'hc22894cd, 32'h4282e749, 32'h41e4573f, 32'hc26b8a03, 32'h42a3b76a, 32'hc23756e2, 32'h42626b0f, 32'hc2614197};
test_output[6216:6223] = '{32'h0, 32'h4282e749, 32'h41e4573f, 32'h0, 32'h42a3b76a, 32'h0, 32'h42626b0f, 32'h0};
test_input[6224:6231] = '{32'h429a89e2, 32'hc28895fe, 32'hc1044d71, 32'h4140ccdd, 32'hc22b8edd, 32'hc2a41594, 32'hc1fa8194, 32'h4287c064};
test_output[6224:6231] = '{32'h429a89e2, 32'h0, 32'h0, 32'h4140ccdd, 32'h0, 32'h0, 32'h0, 32'h4287c064};
test_input[6232:6239] = '{32'hc2be243a, 32'hc22deaf7, 32'h41ed344b, 32'h42a00fbb, 32'h4284c725, 32'hc097a337, 32'hc2b73660, 32'hc23fa7b8};
test_output[6232:6239] = '{32'h0, 32'h0, 32'h41ed344b, 32'h42a00fbb, 32'h4284c725, 32'h0, 32'h0, 32'h0};
test_input[6240:6247] = '{32'hc214d177, 32'h42aedc49, 32'hc21b5553, 32'h42b42698, 32'hc26a52c6, 32'hc2c3cbed, 32'h40ab187d, 32'hc2bd15f1};
test_output[6240:6247] = '{32'h0, 32'h42aedc49, 32'h0, 32'h42b42698, 32'h0, 32'h0, 32'h40ab187d, 32'h0};
test_input[6248:6255] = '{32'h42910e18, 32'h4280aba9, 32'hc1a3ea69, 32'h41a49aef, 32'h4248779c, 32'hc2c5d49b, 32'h41dafda2, 32'hc214066d};
test_output[6248:6255] = '{32'h42910e18, 32'h4280aba9, 32'h0, 32'h41a49aef, 32'h4248779c, 32'h0, 32'h41dafda2, 32'h0};
test_input[6256:6263] = '{32'h41bef6fb, 32'hc0e2c69e, 32'hc1fd0a2d, 32'hc1feb08e, 32'hc1bf3bb3, 32'h420eaf0a, 32'h42083cb9, 32'hc0709bc7};
test_output[6256:6263] = '{32'h41bef6fb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420eaf0a, 32'h42083cb9, 32'h0};
test_input[6264:6271] = '{32'h4207558a, 32'h4280c711, 32'h427f4af1, 32'h40ffa4af, 32'hc2665d08, 32'h4172c71b, 32'hc2809cbe, 32'hc21e31d8};
test_output[6264:6271] = '{32'h4207558a, 32'h4280c711, 32'h427f4af1, 32'h40ffa4af, 32'h0, 32'h4172c71b, 32'h0, 32'h0};
test_input[6272:6279] = '{32'hc241d9a9, 32'h404fbe78, 32'hc2828f26, 32'hc2a14bc2, 32'hc25cd72d, 32'h41236be1, 32'hc041e580, 32'hc2b9746a};
test_output[6272:6279] = '{32'h0, 32'h404fbe78, 32'h0, 32'h0, 32'h0, 32'h41236be1, 32'h0, 32'h0};
test_input[6280:6287] = '{32'hc26fc3dd, 32'hc2bd158c, 32'h41a4540d, 32'h429aa69c, 32'hc2bf5328, 32'hc29d0bb9, 32'hc286c140, 32'hc2441af8};
test_output[6280:6287] = '{32'h0, 32'h0, 32'h41a4540d, 32'h429aa69c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6288:6295] = '{32'hc2aa15de, 32'hc295a38b, 32'h3eb8fde8, 32'hc2255ef2, 32'hc251ca24, 32'hc04421c0, 32'h420a3165, 32'h40d3b3b4};
test_output[6288:6295] = '{32'h0, 32'h0, 32'h3eb8fde8, 32'h0, 32'h0, 32'h0, 32'h420a3165, 32'h40d3b3b4};
test_input[6296:6303] = '{32'hc2b24280, 32'h42040084, 32'h4291f153, 32'h4225efc1, 32'h3f1670e0, 32'h42b3ad1f, 32'hc17e5241, 32'hc285a1c9};
test_output[6296:6303] = '{32'h0, 32'h42040084, 32'h4291f153, 32'h4225efc1, 32'h3f1670e0, 32'h42b3ad1f, 32'h0, 32'h0};
test_input[6304:6311] = '{32'h42b4e47f, 32'hc23cd9a9, 32'h422e70e4, 32'h429d5245, 32'h4244177c, 32'hc294a8af, 32'h42c48471, 32'h42741d1f};
test_output[6304:6311] = '{32'h42b4e47f, 32'h0, 32'h422e70e4, 32'h429d5245, 32'h4244177c, 32'h0, 32'h42c48471, 32'h42741d1f};
test_input[6312:6319] = '{32'hc241087b, 32'h4287130c, 32'hc239c852, 32'hc2882079, 32'h4259b73f, 32'h421fd921, 32'h42a3ed88, 32'h427d4438};
test_output[6312:6319] = '{32'h0, 32'h4287130c, 32'h0, 32'h0, 32'h4259b73f, 32'h421fd921, 32'h42a3ed88, 32'h427d4438};
test_input[6320:6327] = '{32'h42572b4a, 32'h426b1849, 32'h4182ac9b, 32'hc1f6fe5d, 32'h41e2df88, 32'h42b0e4da, 32'h428df80b, 32'h420f65eb};
test_output[6320:6327] = '{32'h42572b4a, 32'h426b1849, 32'h4182ac9b, 32'h0, 32'h41e2df88, 32'h42b0e4da, 32'h428df80b, 32'h420f65eb};
test_input[6328:6335] = '{32'h42c056c4, 32'hc013cd38, 32'h426724fa, 32'h418a7ede, 32'h42987767, 32'hc2aaae68, 32'h42b0dff5, 32'hc2911f8f};
test_output[6328:6335] = '{32'h42c056c4, 32'h0, 32'h426724fa, 32'h418a7ede, 32'h42987767, 32'h0, 32'h42b0dff5, 32'h0};
test_input[6336:6343] = '{32'hc2b30c85, 32'hc1c6329a, 32'hc28db204, 32'hc26b5b1f, 32'hc2c393e8, 32'h42b74b6b, 32'hc1fa417f, 32'h4227b68c};
test_output[6336:6343] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b74b6b, 32'h0, 32'h4227b68c};
test_input[6344:6351] = '{32'hc1183fe3, 32'hc2b785d1, 32'h426e0896, 32'hc23a3f07, 32'hc24b1bdb, 32'hc1e37813, 32'h4145869e, 32'h4284c1bb};
test_output[6344:6351] = '{32'h0, 32'h0, 32'h426e0896, 32'h0, 32'h0, 32'h0, 32'h4145869e, 32'h4284c1bb};
test_input[6352:6359] = '{32'hc2b97ba5, 32'hc10f5b39, 32'hc1cd6520, 32'h421852c3, 32'hc2b1f98f, 32'hc2460464, 32'hc1cf0fdf, 32'h4200d998};
test_output[6352:6359] = '{32'h0, 32'h0, 32'h0, 32'h421852c3, 32'h0, 32'h0, 32'h0, 32'h4200d998};
test_input[6360:6367] = '{32'hc27d059a, 32'h4298a78c, 32'hc20c7196, 32'h400df41b, 32'hc2c5e618, 32'hc10db400, 32'hc1ec0385, 32'hc1b3b81f};
test_output[6360:6367] = '{32'h0, 32'h4298a78c, 32'h0, 32'h400df41b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6368:6375] = '{32'h41f50819, 32'h42a3813f, 32'h42c1c508, 32'h4216a048, 32'h425cc744, 32'hc284b85a, 32'hc0d04c2e, 32'hc1d0f900};
test_output[6368:6375] = '{32'h41f50819, 32'h42a3813f, 32'h42c1c508, 32'h4216a048, 32'h425cc744, 32'h0, 32'h0, 32'h0};
test_input[6376:6383] = '{32'h42bb5d80, 32'hc263912f, 32'hc1bf975c, 32'h42075518, 32'h412104f7, 32'h429a0e19, 32'h42c72fd5, 32'h4119c05b};
test_output[6376:6383] = '{32'h42bb5d80, 32'h0, 32'h0, 32'h42075518, 32'h412104f7, 32'h429a0e19, 32'h42c72fd5, 32'h4119c05b};
test_input[6384:6391] = '{32'h42b2904f, 32'h3e511ed6, 32'h42180bb0, 32'hc0c67c2e, 32'h4230a6f3, 32'h42b7851b, 32'h42c0a4cd, 32'hc291ff7c};
test_output[6384:6391] = '{32'h42b2904f, 32'h3e511ed6, 32'h42180bb0, 32'h0, 32'h4230a6f3, 32'h42b7851b, 32'h42c0a4cd, 32'h0};
test_input[6392:6399] = '{32'h429fadf5, 32'hc1dc7830, 32'hc2a2a80c, 32'h40f0e1f1, 32'hc2c7942a, 32'h425876f9, 32'hc28a7ddd, 32'h42b270ad};
test_output[6392:6399] = '{32'h429fadf5, 32'h0, 32'h0, 32'h40f0e1f1, 32'h0, 32'h425876f9, 32'h0, 32'h42b270ad};
test_input[6400:6407] = '{32'h40d85095, 32'hc1288f95, 32'hc274d3a2, 32'hc26a5c12, 32'h42111172, 32'hc24593a6, 32'h429120ee, 32'h41ea2cd8};
test_output[6400:6407] = '{32'h40d85095, 32'h0, 32'h0, 32'h0, 32'h42111172, 32'h0, 32'h429120ee, 32'h41ea2cd8};
test_input[6408:6415] = '{32'hc203f919, 32'hc2c251bb, 32'hc2bc370a, 32'h42a6cb4a, 32'hc1e337be, 32'h42b3dd99, 32'hc27f484d, 32'h4286a026};
test_output[6408:6415] = '{32'h0, 32'h0, 32'h0, 32'h42a6cb4a, 32'h0, 32'h42b3dd99, 32'h0, 32'h4286a026};
test_input[6416:6423] = '{32'hc0874a6f, 32'h429ee655, 32'h42be4e70, 32'hc1bf7ff3, 32'h429d9473, 32'h4235b6b7, 32'hc2288349, 32'h42a9bb14};
test_output[6416:6423] = '{32'h0, 32'h429ee655, 32'h42be4e70, 32'h0, 32'h429d9473, 32'h4235b6b7, 32'h0, 32'h42a9bb14};
test_input[6424:6431] = '{32'hc2369643, 32'hc213a61a, 32'h4256e127, 32'h42b14c6d, 32'h42c5cba6, 32'h421b7687, 32'h4082c92a, 32'h420b679e};
test_output[6424:6431] = '{32'h0, 32'h0, 32'h4256e127, 32'h42b14c6d, 32'h42c5cba6, 32'h421b7687, 32'h4082c92a, 32'h420b679e};
test_input[6432:6439] = '{32'h42bfad3d, 32'hc278b7d0, 32'hc28e5ac9, 32'hc1b0147c, 32'hc2c3a513, 32'h42a30309, 32'h421541bc, 32'h4279f398};
test_output[6432:6439] = '{32'h42bfad3d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a30309, 32'h421541bc, 32'h4279f398};
test_input[6440:6447] = '{32'h4241504b, 32'hc0fe2b60, 32'hc297276b, 32'hc2552e27, 32'h419d44b8, 32'hc2316d14, 32'hc1c27498, 32'h42a236a5};
test_output[6440:6447] = '{32'h4241504b, 32'h0, 32'h0, 32'h0, 32'h419d44b8, 32'h0, 32'h0, 32'h42a236a5};
test_input[6448:6455] = '{32'hc1379d6e, 32'hc16b2337, 32'h40578d52, 32'hc28668a2, 32'hc2b4eef4, 32'h413937de, 32'h421ab174, 32'hc282b16d};
test_output[6448:6455] = '{32'h0, 32'h0, 32'h40578d52, 32'h0, 32'h0, 32'h413937de, 32'h421ab174, 32'h0};
test_input[6456:6463] = '{32'h4283c302, 32'h41983da2, 32'h41613e92, 32'h41bf12ed, 32'h4289a281, 32'hc27ba3ab, 32'hc1126922, 32'h424d784f};
test_output[6456:6463] = '{32'h4283c302, 32'h41983da2, 32'h41613e92, 32'h41bf12ed, 32'h4289a281, 32'h0, 32'h0, 32'h424d784f};
test_input[6464:6471] = '{32'hc2935b19, 32'hc2969518, 32'hc2b8e911, 32'hc267766d, 32'h422c4608, 32'hc226f2b2, 32'hc26fbd39, 32'h40efde90};
test_output[6464:6471] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h422c4608, 32'h0, 32'h0, 32'h40efde90};
test_input[6472:6479] = '{32'h423e1944, 32'hc2934647, 32'h41e73d86, 32'h421b86ba, 32'h429621d4, 32'hc2249076, 32'h4286c549, 32'hc2a6c4e9};
test_output[6472:6479] = '{32'h423e1944, 32'h0, 32'h41e73d86, 32'h421b86ba, 32'h429621d4, 32'h0, 32'h4286c549, 32'h0};
test_input[6480:6487] = '{32'h42c3a206, 32'hc295fdd3, 32'hc2c4e90f, 32'hc265bd1f, 32'h42406b6d, 32'h422717fe, 32'h41255556, 32'hc2845eae};
test_output[6480:6487] = '{32'h42c3a206, 32'h0, 32'h0, 32'h0, 32'h42406b6d, 32'h422717fe, 32'h41255556, 32'h0};
test_input[6488:6495] = '{32'h42b6e5ae, 32'h421b93a5, 32'h419d3d92, 32'h424c52ab, 32'h4271a7ef, 32'h41b87122, 32'hbfd4070f, 32'h4121233f};
test_output[6488:6495] = '{32'h42b6e5ae, 32'h421b93a5, 32'h419d3d92, 32'h424c52ab, 32'h4271a7ef, 32'h41b87122, 32'h0, 32'h4121233f};
test_input[6496:6503] = '{32'hc180648c, 32'hc287b312, 32'hc28031da, 32'hc2a77e73, 32'hc22cc37b, 32'h429fea25, 32'hc2be3783, 32'hc19361ac};
test_output[6496:6503] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429fea25, 32'h0, 32'h0};
test_input[6504:6511] = '{32'hc1f564ca, 32'hc2ab93ac, 32'hc2c6c74a, 32'hc28f7f5f, 32'h4153ca61, 32'h4286a036, 32'h42ac5dfd, 32'hbfefa714};
test_output[6504:6511] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4153ca61, 32'h4286a036, 32'h42ac5dfd, 32'h0};
test_input[6512:6519] = '{32'h405d99ad, 32'hc2819e5c, 32'h4284af95, 32'h418815ed, 32'hc2bb7c4d, 32'hc2643645, 32'hc1fcc339, 32'h42a45286};
test_output[6512:6519] = '{32'h405d99ad, 32'h0, 32'h4284af95, 32'h418815ed, 32'h0, 32'h0, 32'h0, 32'h42a45286};
test_input[6520:6527] = '{32'hc28626b2, 32'h42abe85a, 32'hc247b85a, 32'h41773a5d, 32'h4266ffe3, 32'h42b9eb7b, 32'h3f971a4e, 32'h416eb8a2};
test_output[6520:6527] = '{32'h0, 32'h42abe85a, 32'h0, 32'h41773a5d, 32'h4266ffe3, 32'h42b9eb7b, 32'h3f971a4e, 32'h416eb8a2};
test_input[6528:6535] = '{32'hc19ea801, 32'hc1886a64, 32'h427dd4b6, 32'h40e87a9f, 32'hbff9dacd, 32'hc28f10e5, 32'hc1a81ec2, 32'hc2895261};
test_output[6528:6535] = '{32'h0, 32'h0, 32'h427dd4b6, 32'h40e87a9f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6536:6543] = '{32'hc2ab5466, 32'hc204a4b0, 32'h42686211, 32'h422d771a, 32'hc2814767, 32'hc091c10c, 32'h42b9a4e6, 32'hc2140e16};
test_output[6536:6543] = '{32'h0, 32'h0, 32'h42686211, 32'h422d771a, 32'h0, 32'h0, 32'h42b9a4e6, 32'h0};
test_input[6544:6551] = '{32'hc29fb9ec, 32'h42490e29, 32'hc26a5e24, 32'hc214322b, 32'hc08b1f9c, 32'h413876d7, 32'h41e3c21f, 32'hc284e216};
test_output[6544:6551] = '{32'h0, 32'h42490e29, 32'h0, 32'h0, 32'h0, 32'h413876d7, 32'h41e3c21f, 32'h0};
test_input[6552:6559] = '{32'h41b5b64c, 32'h41469dbb, 32'h40ab6c85, 32'hc12ae703, 32'h4247337b, 32'h428b381b, 32'h42c51352, 32'hc168def9};
test_output[6552:6559] = '{32'h41b5b64c, 32'h41469dbb, 32'h40ab6c85, 32'h0, 32'h4247337b, 32'h428b381b, 32'h42c51352, 32'h0};
test_input[6560:6567] = '{32'h4103d038, 32'hc29b2438, 32'hc2bde7b6, 32'hc2b026c5, 32'h4126ef2d, 32'hc289ce76, 32'h42a782c8, 32'h4283751c};
test_output[6560:6567] = '{32'h4103d038, 32'h0, 32'h0, 32'h0, 32'h4126ef2d, 32'h0, 32'h42a782c8, 32'h4283751c};
test_input[6568:6575] = '{32'h42ba97a0, 32'hc28de9b5, 32'h3f787899, 32'hc22b8083, 32'hc26dc4f5, 32'h416a4c5b, 32'hc25c728a, 32'h417e86ce};
test_output[6568:6575] = '{32'h42ba97a0, 32'h0, 32'h3f787899, 32'h0, 32'h0, 32'h416a4c5b, 32'h0, 32'h417e86ce};
test_input[6576:6583] = '{32'hc1a6d14b, 32'h4205c2f1, 32'hc22d0b05, 32'hc0221bf7, 32'h41a75c13, 32'hc285a50a, 32'h4285c833, 32'h4267d830};
test_output[6576:6583] = '{32'h0, 32'h4205c2f1, 32'h0, 32'h0, 32'h41a75c13, 32'h0, 32'h4285c833, 32'h4267d830};
test_input[6584:6591] = '{32'h4285fa5e, 32'h420e10a1, 32'hc1faf752, 32'h41732bdb, 32'h41cfd357, 32'h42105a01, 32'h420cc690, 32'h419f2767};
test_output[6584:6591] = '{32'h4285fa5e, 32'h420e10a1, 32'h0, 32'h41732bdb, 32'h41cfd357, 32'h42105a01, 32'h420cc690, 32'h419f2767};
test_input[6592:6599] = '{32'h420b9b9b, 32'hc295e994, 32'h416873a2, 32'hc2c2ccdc, 32'hc10d1b72, 32'h42b48809, 32'hc2849906, 32'h41d8ea60};
test_output[6592:6599] = '{32'h420b9b9b, 32'h0, 32'h416873a2, 32'h0, 32'h0, 32'h42b48809, 32'h0, 32'h41d8ea60};
test_input[6600:6607] = '{32'h4140c87b, 32'h42988297, 32'hc12d2025, 32'h413ea5af, 32'h42245415, 32'hc21010f7, 32'hc2307775, 32'hc2c4c302};
test_output[6600:6607] = '{32'h4140c87b, 32'h42988297, 32'h0, 32'h413ea5af, 32'h42245415, 32'h0, 32'h0, 32'h0};
test_input[6608:6615] = '{32'h42bb958f, 32'hc277f203, 32'hc266f910, 32'hc28f393c, 32'hc2963312, 32'hc266fb15, 32'h413a104a, 32'hc2240e0e};
test_output[6608:6615] = '{32'h42bb958f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h413a104a, 32'h0};
test_input[6616:6623] = '{32'hc2c787eb, 32'hc22da9e3, 32'h416e81a4, 32'h4112ec15, 32'hc047d24d, 32'h42c0a100, 32'h42b23be3, 32'h4217929f};
test_output[6616:6623] = '{32'h0, 32'h0, 32'h416e81a4, 32'h4112ec15, 32'h0, 32'h42c0a100, 32'h42b23be3, 32'h4217929f};
test_input[6624:6631] = '{32'hc2268544, 32'hc299c652, 32'hc22dc876, 32'hbf6ad300, 32'hc2105702, 32'h428d924f, 32'hc27d7942, 32'h4292baad};
test_output[6624:6631] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428d924f, 32'h0, 32'h4292baad};
test_input[6632:6639] = '{32'hc18ba5bc, 32'h42ae0567, 32'h4264f140, 32'hc1814355, 32'hc1bfa4d4, 32'hc2b2df69, 32'hc241a98a, 32'hc0f2b790};
test_output[6632:6639] = '{32'h0, 32'h42ae0567, 32'h4264f140, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6640:6647] = '{32'hc1fb3b5e, 32'hc220888f, 32'h429d8133, 32'h4280a019, 32'h4290e22a, 32'hc16d4ef8, 32'h4193b0d5, 32'hc06c7c21};
test_output[6640:6647] = '{32'h0, 32'h0, 32'h429d8133, 32'h4280a019, 32'h4290e22a, 32'h0, 32'h4193b0d5, 32'h0};
test_input[6648:6655] = '{32'hc2a2d6b8, 32'h418c2675, 32'hc23b0cc6, 32'h4120ef3f, 32'hc287f1fa, 32'h420c1d9b, 32'h42a826c6, 32'h42c0391f};
test_output[6648:6655] = '{32'h0, 32'h418c2675, 32'h0, 32'h4120ef3f, 32'h0, 32'h420c1d9b, 32'h42a826c6, 32'h42c0391f};
test_input[6656:6663] = '{32'hc2516b50, 32'h42558d67, 32'h421208a9, 32'h42124e4b, 32'hc210a68a, 32'h421f4456, 32'h42c6b798, 32'hc2a00048};
test_output[6656:6663] = '{32'h0, 32'h42558d67, 32'h421208a9, 32'h42124e4b, 32'h0, 32'h421f4456, 32'h42c6b798, 32'h0};
test_input[6664:6671] = '{32'h4206637a, 32'hc22a63cf, 32'h41aaf79c, 32'h4102d9eb, 32'h42528ead, 32'hc27a019d, 32'hc26af0cc, 32'h41a6b855};
test_output[6664:6671] = '{32'h4206637a, 32'h0, 32'h41aaf79c, 32'h4102d9eb, 32'h42528ead, 32'h0, 32'h0, 32'h41a6b855};
test_input[6672:6679] = '{32'h420943e5, 32'hc294ebb5, 32'hc2a49c16, 32'hc1f8aac5, 32'hc207a2e1, 32'hc28a9b44, 32'hc15f0887, 32'hc0ef5c74};
test_output[6672:6679] = '{32'h420943e5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6680:6687] = '{32'h421bfa77, 32'h4291bb34, 32'h424c6dfc, 32'hc0bb78bd, 32'hc293dfca, 32'hc2c36c93, 32'h425e56fe, 32'h425f59bc};
test_output[6680:6687] = '{32'h421bfa77, 32'h4291bb34, 32'h424c6dfc, 32'h0, 32'h0, 32'h0, 32'h425e56fe, 32'h425f59bc};
test_input[6688:6695] = '{32'hc27beed2, 32'hc29526d0, 32'hc2179202, 32'h41c3d5fa, 32'h42293ca1, 32'h42237858, 32'h41b7e01d, 32'h422f1d08};
test_output[6688:6695] = '{32'h0, 32'h0, 32'h0, 32'h41c3d5fa, 32'h42293ca1, 32'h42237858, 32'h41b7e01d, 32'h422f1d08};
test_input[6696:6703] = '{32'h40598ede, 32'hc283d396, 32'hc2443f75, 32'h418d6afe, 32'hc273cd26, 32'hc1f20ce4, 32'h42984087, 32'hc2b4977f};
test_output[6696:6703] = '{32'h40598ede, 32'h0, 32'h0, 32'h418d6afe, 32'h0, 32'h0, 32'h42984087, 32'h0};
test_input[6704:6711] = '{32'h4259f357, 32'h42147834, 32'h42a5c3f4, 32'h42a14f86, 32'hc1ee2f48, 32'h4246a996, 32'h429b9793, 32'h413943aa};
test_output[6704:6711] = '{32'h4259f357, 32'h42147834, 32'h42a5c3f4, 32'h42a14f86, 32'h0, 32'h4246a996, 32'h429b9793, 32'h413943aa};
test_input[6712:6719] = '{32'h42127ab2, 32'hc010c615, 32'hc169724c, 32'h413aa6f9, 32'hc2414027, 32'h425f31fb, 32'hc217e079, 32'h42849ac8};
test_output[6712:6719] = '{32'h42127ab2, 32'h0, 32'h0, 32'h413aa6f9, 32'h0, 32'h425f31fb, 32'h0, 32'h42849ac8};
test_input[6720:6727] = '{32'hc28b8bbe, 32'hc2c3eddd, 32'hc2aaf5a6, 32'hc2c595a6, 32'hc28d8669, 32'h41258bb8, 32'h42c28a5d, 32'hc1495f82};
test_output[6720:6727] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41258bb8, 32'h42c28a5d, 32'h0};
test_input[6728:6735] = '{32'h42bd5876, 32'h4258c0c1, 32'hc288257c, 32'h4295605b, 32'h42bed555, 32'hc253a58e, 32'h41c4e86a, 32'hc247651f};
test_output[6728:6735] = '{32'h42bd5876, 32'h4258c0c1, 32'h0, 32'h4295605b, 32'h42bed555, 32'h0, 32'h41c4e86a, 32'h0};
test_input[6736:6743] = '{32'hc1ab95fa, 32'hc2090ff7, 32'h417fa611, 32'hc1fc2fa6, 32'hc2a8f3b7, 32'hc28fef4b, 32'h41122fd9, 32'h426cfdbf};
test_output[6736:6743] = '{32'h0, 32'h0, 32'h417fa611, 32'h0, 32'h0, 32'h0, 32'h41122fd9, 32'h426cfdbf};
test_input[6744:6751] = '{32'h42b36288, 32'h42862774, 32'hc23aa26e, 32'h420f514d, 32'h4275ca55, 32'hc2392773, 32'h42b0e3ea, 32'hc2c729a2};
test_output[6744:6751] = '{32'h42b36288, 32'h42862774, 32'h0, 32'h420f514d, 32'h4275ca55, 32'h0, 32'h42b0e3ea, 32'h0};
test_input[6752:6759] = '{32'hbf9e0a99, 32'h420a7e01, 32'h428420eb, 32'h427f3077, 32'hc2007316, 32'hc2840a1d, 32'hc28a5fb6, 32'hc081ffa4};
test_output[6752:6759] = '{32'h0, 32'h420a7e01, 32'h428420eb, 32'h427f3077, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6760:6767] = '{32'h40af4ca8, 32'h42ab559e, 32'hc27e5c95, 32'hc1010fc5, 32'h428a1ad5, 32'hc19b12b7, 32'h40a56a86, 32'h425b871f};
test_output[6760:6767] = '{32'h40af4ca8, 32'h42ab559e, 32'h0, 32'h0, 32'h428a1ad5, 32'h0, 32'h40a56a86, 32'h425b871f};
test_input[6768:6775] = '{32'hc20ebc47, 32'h42a58c18, 32'hc23d3a69, 32'h4291eba8, 32'h422e784c, 32'h427c4398, 32'hc225eae8, 32'h40980329};
test_output[6768:6775] = '{32'h0, 32'h42a58c18, 32'h0, 32'h4291eba8, 32'h422e784c, 32'h427c4398, 32'h0, 32'h40980329};
test_input[6776:6783] = '{32'hc29cdd79, 32'h422f1cc5, 32'h422b7ff3, 32'hc2c7fe17, 32'h427170e8, 32'hc2338129, 32'hc12e739c, 32'h4297598e};
test_output[6776:6783] = '{32'h0, 32'h422f1cc5, 32'h422b7ff3, 32'h0, 32'h427170e8, 32'h0, 32'h0, 32'h4297598e};
test_input[6784:6791] = '{32'h42aea61e, 32'hc2c0838b, 32'h427cad41, 32'hc2b554d4, 32'h4275a4d7, 32'hc1b216ad, 32'h42832269, 32'h42a6f2b7};
test_output[6784:6791] = '{32'h42aea61e, 32'h0, 32'h427cad41, 32'h0, 32'h4275a4d7, 32'h0, 32'h42832269, 32'h42a6f2b7};
test_input[6792:6799] = '{32'h41b050c5, 32'hc20cc8fc, 32'hc0b3d50d, 32'hc1a044d9, 32'h4130592d, 32'hc201f628, 32'hc233a4e7, 32'hc15c1943};
test_output[6792:6799] = '{32'h41b050c5, 32'h0, 32'h0, 32'h0, 32'h4130592d, 32'h0, 32'h0, 32'h0};
test_input[6800:6807] = '{32'hc0f7410a, 32'h410a3038, 32'h42998233, 32'h42204f8e, 32'h429480b9, 32'hc2a7a1e7, 32'h41806d04, 32'hc24d87da};
test_output[6800:6807] = '{32'h0, 32'h410a3038, 32'h42998233, 32'h42204f8e, 32'h429480b9, 32'h0, 32'h41806d04, 32'h0};
test_input[6808:6815] = '{32'h42ac467d, 32'hc08b24a4, 32'h42b9069f, 32'hc225589e, 32'hc1870603, 32'h425bae25, 32'h429bb746, 32'hc213b6f8};
test_output[6808:6815] = '{32'h42ac467d, 32'h0, 32'h42b9069f, 32'h0, 32'h0, 32'h425bae25, 32'h429bb746, 32'h0};
test_input[6816:6823] = '{32'hc1cfa4cc, 32'hc2c641e4, 32'h428743d8, 32'h4252c5e3, 32'h40ce5b0a, 32'h42a5290c, 32'h41290eec, 32'h42ac0dbc};
test_output[6816:6823] = '{32'h0, 32'h0, 32'h428743d8, 32'h4252c5e3, 32'h40ce5b0a, 32'h42a5290c, 32'h41290eec, 32'h42ac0dbc};
test_input[6824:6831] = '{32'hbf8813dd, 32'hc2032eeb, 32'h4110ce8f, 32'h4243758a, 32'h423c1533, 32'h424e20d7, 32'h428492d9, 32'h4241a866};
test_output[6824:6831] = '{32'h0, 32'h0, 32'h4110ce8f, 32'h4243758a, 32'h423c1533, 32'h424e20d7, 32'h428492d9, 32'h4241a866};
test_input[6832:6839] = '{32'h4142cbb0, 32'h429866fb, 32'hc2c19fd4, 32'hc244aa4c, 32'h421dd887, 32'h41e450b6, 32'h42895192, 32'hc2be34b8};
test_output[6832:6839] = '{32'h4142cbb0, 32'h429866fb, 32'h0, 32'h0, 32'h421dd887, 32'h41e450b6, 32'h42895192, 32'h0};
test_input[6840:6847] = '{32'h42c64e3e, 32'hc2391d8e, 32'hc2446e07, 32'h429fb9ad, 32'hc125c0fd, 32'hc12a6322, 32'h4282825d, 32'h41fc355d};
test_output[6840:6847] = '{32'h42c64e3e, 32'h0, 32'h0, 32'h429fb9ad, 32'h0, 32'h0, 32'h4282825d, 32'h41fc355d};
test_input[6848:6855] = '{32'h4149dd31, 32'hc1029496, 32'h41a6d51b, 32'h41e0940b, 32'hc1b448e3, 32'hc2ae12fb, 32'h42a0cdff, 32'hc2b1392b};
test_output[6848:6855] = '{32'h4149dd31, 32'h0, 32'h41a6d51b, 32'h41e0940b, 32'h0, 32'h0, 32'h42a0cdff, 32'h0};
test_input[6856:6863] = '{32'h429e032b, 32'hc2b44ee0, 32'hc2162439, 32'h425dc9be, 32'h423fccd3, 32'hc29f87a6, 32'hc1172a73, 32'h415a0533};
test_output[6856:6863] = '{32'h429e032b, 32'h0, 32'h0, 32'h425dc9be, 32'h423fccd3, 32'h0, 32'h0, 32'h415a0533};
test_input[6864:6871] = '{32'h3e10b8d6, 32'hc162b9db, 32'hc192be07, 32'hc20b9650, 32'h40b3d214, 32'h426bef57, 32'h41524915, 32'h420c8e46};
test_output[6864:6871] = '{32'h3e10b8d6, 32'h0, 32'h0, 32'h0, 32'h40b3d214, 32'h426bef57, 32'h41524915, 32'h420c8e46};
test_input[6872:6879] = '{32'hc23e6bce, 32'hc1d08073, 32'h421d53d7, 32'h429ab417, 32'hc25d1db4, 32'hc2c3ee5a, 32'h42ad2bb6, 32'hc29f146a};
test_output[6872:6879] = '{32'h0, 32'h0, 32'h421d53d7, 32'h429ab417, 32'h0, 32'h0, 32'h42ad2bb6, 32'h0};
test_input[6880:6887] = '{32'hc2b53c0e, 32'hc1520b19, 32'hc108690e, 32'hc23a7fc6, 32'h422cc69a, 32'hc2c5b863, 32'h42a10ca5, 32'hc13b3420};
test_output[6880:6887] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h422cc69a, 32'h0, 32'h42a10ca5, 32'h0};
test_input[6888:6895] = '{32'h42a63ff2, 32'h42972046, 32'hc1d57d17, 32'h42aa9d98, 32'hc28eb1b5, 32'h4115171f, 32'hc2c3a6aa, 32'hc233f91c};
test_output[6888:6895] = '{32'h42a63ff2, 32'h42972046, 32'h0, 32'h42aa9d98, 32'h0, 32'h4115171f, 32'h0, 32'h0};
test_input[6896:6903] = '{32'h427590ca, 32'hc206bdd6, 32'hc2978ca5, 32'h428192a2, 32'hc2ba7794, 32'h41ea0393, 32'hc0ec6af3, 32'hc1a9fab0};
test_output[6896:6903] = '{32'h427590ca, 32'h0, 32'h0, 32'h428192a2, 32'h0, 32'h41ea0393, 32'h0, 32'h0};
test_input[6904:6911] = '{32'h4264c362, 32'h417175fc, 32'hc205612c, 32'h42541f0b, 32'h42b3ffea, 32'h42a6b0d4, 32'h419620aa, 32'h4195024a};
test_output[6904:6911] = '{32'h4264c362, 32'h417175fc, 32'h0, 32'h42541f0b, 32'h42b3ffea, 32'h42a6b0d4, 32'h419620aa, 32'h4195024a};
test_input[6912:6919] = '{32'h42b8898d, 32'hc19b531c, 32'h424ca003, 32'h429109d8, 32'hc2918cba, 32'hc28bdda4, 32'hc1b82345, 32'hc1d59fa8};
test_output[6912:6919] = '{32'h42b8898d, 32'h0, 32'h424ca003, 32'h429109d8, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6920:6927] = '{32'h42896855, 32'h42918d0f, 32'h42a78c1e, 32'h416b2b28, 32'h42bf9277, 32'hc29ea920, 32'h41f5dd3f, 32'hc2bc0f5a};
test_output[6920:6927] = '{32'h42896855, 32'h42918d0f, 32'h42a78c1e, 32'h416b2b28, 32'h42bf9277, 32'h0, 32'h41f5dd3f, 32'h0};
test_input[6928:6935] = '{32'h426d3fa0, 32'h42a7f5a5, 32'h424200db, 32'h422ec7a4, 32'h41efe1fe, 32'h42010b36, 32'h418deb4c, 32'hc15d42eb};
test_output[6928:6935] = '{32'h426d3fa0, 32'h42a7f5a5, 32'h424200db, 32'h422ec7a4, 32'h41efe1fe, 32'h42010b36, 32'h418deb4c, 32'h0};
test_input[6936:6943] = '{32'h41d96a65, 32'h42259cf2, 32'h426315ed, 32'hc14cb05a, 32'hc0928324, 32'hc0cb6637, 32'h429725c7, 32'h424532cb};
test_output[6936:6943] = '{32'h41d96a65, 32'h42259cf2, 32'h426315ed, 32'h0, 32'h0, 32'h0, 32'h429725c7, 32'h424532cb};
test_input[6944:6951] = '{32'h42a1c03a, 32'hc2ae186a, 32'h412a7a98, 32'h4236c9ed, 32'h423f5667, 32'hc18bb5ea, 32'hc1bb0c65, 32'hc2744822};
test_output[6944:6951] = '{32'h42a1c03a, 32'h0, 32'h412a7a98, 32'h4236c9ed, 32'h423f5667, 32'h0, 32'h0, 32'h0};
test_input[6952:6959] = '{32'hc2656edb, 32'h4207fb46, 32'h42a51792, 32'hc299c571, 32'hc2b3437e, 32'h42b24692, 32'h419ac056, 32'h42a0b0e2};
test_output[6952:6959] = '{32'h0, 32'h4207fb46, 32'h42a51792, 32'h0, 32'h0, 32'h42b24692, 32'h419ac056, 32'h42a0b0e2};
test_input[6960:6967] = '{32'hc285763a, 32'hc1283e6e, 32'hc2bcf7f9, 32'hc1eda144, 32'hc21713dc, 32'hc25ddb8d, 32'h42c22a06, 32'hc2798139};
test_output[6960:6967] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c22a06, 32'h0};
test_input[6968:6975] = '{32'h4257b680, 32'hc2ab0c4e, 32'hc213e89a, 32'hc11303f9, 32'h42632522, 32'hc23e9186, 32'h42c3adac, 32'h421b58b4};
test_output[6968:6975] = '{32'h4257b680, 32'h0, 32'h0, 32'h0, 32'h42632522, 32'h0, 32'h42c3adac, 32'h421b58b4};
test_input[6976:6983] = '{32'h42bfdff9, 32'hc2a7d2b7, 32'hc2b4d847, 32'hc26833a1, 32'h41b37c83, 32'h42710288, 32'hc24d7292, 32'hc2826629};
test_output[6976:6983] = '{32'h42bfdff9, 32'h0, 32'h0, 32'h0, 32'h41b37c83, 32'h42710288, 32'h0, 32'h0};
test_input[6984:6991] = '{32'hc2bb9366, 32'h42142e6b, 32'h418d2682, 32'hbf169f87, 32'h42b0f545, 32'h4240ecc0, 32'hc1b01f86, 32'h428b6733};
test_output[6984:6991] = '{32'h0, 32'h42142e6b, 32'h418d2682, 32'h0, 32'h42b0f545, 32'h4240ecc0, 32'h0, 32'h428b6733};
test_input[6992:6999] = '{32'hc0d425ed, 32'h41269e9b, 32'h42873803, 32'hc2783460, 32'h429aa4c6, 32'h4168e943, 32'hc2b94177, 32'h42917f86};
test_output[6992:6999] = '{32'h0, 32'h41269e9b, 32'h42873803, 32'h0, 32'h429aa4c6, 32'h4168e943, 32'h0, 32'h42917f86};
test_input[7000:7007] = '{32'h412d5a35, 32'h42a1f4ca, 32'h42026fba, 32'h40fcb972, 32'hc1f4eba4, 32'h421f4637, 32'hc2a8b23b, 32'hc16c10e0};
test_output[7000:7007] = '{32'h412d5a35, 32'h42a1f4ca, 32'h42026fba, 32'h40fcb972, 32'h0, 32'h421f4637, 32'h0, 32'h0};
test_input[7008:7015] = '{32'h4110b5ad, 32'h4258b072, 32'hc2583235, 32'h41ff539b, 32'hc24b57c1, 32'h41e14fa9, 32'hc240346c, 32'hc23d9840};
test_output[7008:7015] = '{32'h4110b5ad, 32'h4258b072, 32'h0, 32'h41ff539b, 32'h0, 32'h41e14fa9, 32'h0, 32'h0};
test_input[7016:7023] = '{32'hc29e79e9, 32'h41ad5733, 32'h41b90707, 32'h420bac0d, 32'h4206f5f0, 32'h429968ae, 32'h423fb781, 32'h424f9980};
test_output[7016:7023] = '{32'h0, 32'h41ad5733, 32'h41b90707, 32'h420bac0d, 32'h4206f5f0, 32'h429968ae, 32'h423fb781, 32'h424f9980};
test_input[7024:7031] = '{32'h4060a960, 32'hc21c3516, 32'hc2b0f670, 32'hc2803455, 32'hc2bde861, 32'hc2731631, 32'hc232914d, 32'h429471fd};
test_output[7024:7031] = '{32'h4060a960, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429471fd};
test_input[7032:7039] = '{32'hc26e042e, 32'h4293300a, 32'hc2bb6d18, 32'h427b5f0f, 32'h41e2e6b0, 32'hc2c2be25, 32'h42c6f6a8, 32'hc26d5034};
test_output[7032:7039] = '{32'h0, 32'h4293300a, 32'h0, 32'h427b5f0f, 32'h41e2e6b0, 32'h0, 32'h42c6f6a8, 32'h0};
test_input[7040:7047] = '{32'h428d418c, 32'hc2a23500, 32'h42b4ab3c, 32'h4115798c, 32'hc25f9bde, 32'h40eb3ceb, 32'h4296796c, 32'hc1db279a};
test_output[7040:7047] = '{32'h428d418c, 32'h0, 32'h42b4ab3c, 32'h4115798c, 32'h0, 32'h40eb3ceb, 32'h4296796c, 32'h0};
test_input[7048:7055] = '{32'h426414f3, 32'h425ddd4a, 32'hc2154867, 32'h41e5f429, 32'hc2b989f0, 32'h42b9076f, 32'h427cbffc, 32'h41dca2cf};
test_output[7048:7055] = '{32'h426414f3, 32'h425ddd4a, 32'h0, 32'h41e5f429, 32'h0, 32'h42b9076f, 32'h427cbffc, 32'h41dca2cf};
test_input[7056:7063] = '{32'hc27ffaa9, 32'h425a6e6b, 32'hc0f0d31e, 32'hc288cd8a, 32'h4127afa3, 32'h42bebacc, 32'h42a34c04, 32'h429e846c};
test_output[7056:7063] = '{32'h0, 32'h425a6e6b, 32'h0, 32'h0, 32'h4127afa3, 32'h42bebacc, 32'h42a34c04, 32'h429e846c};
test_input[7064:7071] = '{32'h42b4c630, 32'hc1eda217, 32'h42c0d358, 32'hc28d38cc, 32'hc2c05ed8, 32'h42ab84ab, 32'h424607f1, 32'h4245393f};
test_output[7064:7071] = '{32'h42b4c630, 32'h0, 32'h42c0d358, 32'h0, 32'h0, 32'h42ab84ab, 32'h424607f1, 32'h4245393f};
test_input[7072:7079] = '{32'h428b8eb6, 32'hc2c4fc29, 32'h41ff055d, 32'h40177aac, 32'h423c1b0b, 32'h40e46fda, 32'h4250cc24, 32'hc2401337};
test_output[7072:7079] = '{32'h428b8eb6, 32'h0, 32'h41ff055d, 32'h40177aac, 32'h423c1b0b, 32'h40e46fda, 32'h4250cc24, 32'h0};
test_input[7080:7087] = '{32'hc2ac5a26, 32'h429e3d57, 32'h42867524, 32'h42522e18, 32'h42bb3f4a, 32'hc2937765, 32'hc1d20eaa, 32'h4248d878};
test_output[7080:7087] = '{32'h0, 32'h429e3d57, 32'h42867524, 32'h42522e18, 32'h42bb3f4a, 32'h0, 32'h0, 32'h4248d878};
test_input[7088:7095] = '{32'h428589bb, 32'hc168d2b7, 32'hc2ae5dc8, 32'h41abf44f, 32'h42702b7e, 32'hc2aab11b, 32'hc18b0fd7, 32'hc049d72c};
test_output[7088:7095] = '{32'h428589bb, 32'h0, 32'h0, 32'h41abf44f, 32'h42702b7e, 32'h0, 32'h0, 32'h0};
test_input[7096:7103] = '{32'hc26d8144, 32'h42684e60, 32'h42724353, 32'h4172e7cd, 32'hc28e78c9, 32'hc2adb3cf, 32'hc2020509, 32'h4293bb33};
test_output[7096:7103] = '{32'h0, 32'h42684e60, 32'h42724353, 32'h4172e7cd, 32'h0, 32'h0, 32'h0, 32'h4293bb33};
test_input[7104:7111] = '{32'hc1128c86, 32'hc2b92e6b, 32'h425737a3, 32'hc2c7ee4c, 32'hc0e59ab3, 32'hc2b4a3b4, 32'hc1e7706c, 32'hc28742ee};
test_output[7104:7111] = '{32'h0, 32'h0, 32'h425737a3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7112:7119] = '{32'hc271ac03, 32'h4227803b, 32'h42825074, 32'hc22cdd46, 32'h4160b258, 32'h4261ecab, 32'h42c72aad, 32'hc260d05a};
test_output[7112:7119] = '{32'h0, 32'h4227803b, 32'h42825074, 32'h0, 32'h4160b258, 32'h4261ecab, 32'h42c72aad, 32'h0};
test_input[7120:7127] = '{32'hc29a91bc, 32'hc28a7b2d, 32'hc2697811, 32'h425bed48, 32'h40a47a95, 32'h418188df, 32'h4280b26f, 32'h42ac1360};
test_output[7120:7127] = '{32'h0, 32'h0, 32'h0, 32'h425bed48, 32'h40a47a95, 32'h418188df, 32'h4280b26f, 32'h42ac1360};
test_input[7128:7135] = '{32'hc285210d, 32'h41ed8db0, 32'h4287e51f, 32'hc2a3937b, 32'hc289131f, 32'h420d469d, 32'hc103aa1c, 32'h428c8270};
test_output[7128:7135] = '{32'h0, 32'h41ed8db0, 32'h4287e51f, 32'h0, 32'h0, 32'h420d469d, 32'h0, 32'h428c8270};
test_input[7136:7143] = '{32'hc29a2ffb, 32'hc2b3da90, 32'h42782500, 32'h42b1de63, 32'hc2448061, 32'hc20b1124, 32'h41da9eb3, 32'hc1da3f51};
test_output[7136:7143] = '{32'h0, 32'h0, 32'h42782500, 32'h42b1de63, 32'h0, 32'h0, 32'h41da9eb3, 32'h0};
test_input[7144:7151] = '{32'h42453df8, 32'hc27bbf80, 32'hc24ae979, 32'h42c67025, 32'hc27221f1, 32'hc2a1bd7f, 32'hc2ae16e3, 32'hc2b9b5bb};
test_output[7144:7151] = '{32'h42453df8, 32'h0, 32'h0, 32'h42c67025, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7152:7159] = '{32'h41c10a10, 32'hc291568c, 32'hc1e8d36b, 32'h41e2d2b6, 32'h416a019e, 32'h428d3f96, 32'h42a41a86, 32'h42aa4a90};
test_output[7152:7159] = '{32'h41c10a10, 32'h0, 32'h0, 32'h41e2d2b6, 32'h416a019e, 32'h428d3f96, 32'h42a41a86, 32'h42aa4a90};
test_input[7160:7167] = '{32'hc2b2d4d3, 32'h40eed641, 32'hc289222a, 32'h41e0e7e5, 32'h422f3545, 32'h4215d63e, 32'h4299eb8b, 32'h42b635ce};
test_output[7160:7167] = '{32'h0, 32'h40eed641, 32'h0, 32'h41e0e7e5, 32'h422f3545, 32'h4215d63e, 32'h4299eb8b, 32'h42b635ce};
test_input[7168:7175] = '{32'h42768b29, 32'h42a39421, 32'h429b1bef, 32'hc22feaaf, 32'hc2975485, 32'h42333955, 32'h4194ffec, 32'h3fc055ce};
test_output[7168:7175] = '{32'h42768b29, 32'h42a39421, 32'h429b1bef, 32'h0, 32'h0, 32'h42333955, 32'h4194ffec, 32'h3fc055ce};
test_input[7176:7183] = '{32'h416a2a23, 32'h42b79498, 32'h42adfcfb, 32'hc0819de2, 32'hc1e0b7c1, 32'hc1ecfce3, 32'h40396691, 32'hc246179f};
test_output[7176:7183] = '{32'h416a2a23, 32'h42b79498, 32'h42adfcfb, 32'h0, 32'h0, 32'h0, 32'h40396691, 32'h0};
test_input[7184:7191] = '{32'hc267b16d, 32'h42a11ad1, 32'h429d55d4, 32'h42c221ad, 32'h429472c7, 32'hc21a3697, 32'hc27acfa6, 32'hc1c6dc8f};
test_output[7184:7191] = '{32'h0, 32'h42a11ad1, 32'h429d55d4, 32'h42c221ad, 32'h429472c7, 32'h0, 32'h0, 32'h0};
test_input[7192:7199] = '{32'h4299982e, 32'h413bace4, 32'hc2a7f5ce, 32'hc1f2e5b2, 32'hc21ad738, 32'h42b948de, 32'h41a77987, 32'h423eeb86};
test_output[7192:7199] = '{32'h4299982e, 32'h413bace4, 32'h0, 32'h0, 32'h0, 32'h42b948de, 32'h41a77987, 32'h423eeb86};
test_input[7200:7207] = '{32'hc2788e2d, 32'hc1d405e6, 32'hc2be61c0, 32'h42918273, 32'h4285d455, 32'h42316e4e, 32'h421dc460, 32'h41e20468};
test_output[7200:7207] = '{32'h0, 32'h0, 32'h0, 32'h42918273, 32'h4285d455, 32'h42316e4e, 32'h421dc460, 32'h41e20468};
test_input[7208:7215] = '{32'hc1707c5f, 32'h42b751be, 32'hc10a00df, 32'hbfbbe6ad, 32'h429e3e33, 32'hc29a584d, 32'h424959c8, 32'hc25f0334};
test_output[7208:7215] = '{32'h0, 32'h42b751be, 32'h0, 32'h0, 32'h429e3e33, 32'h0, 32'h424959c8, 32'h0};
test_input[7216:7223] = '{32'h40daf1be, 32'h41929660, 32'hc284d1d7, 32'hc139f30b, 32'hc1f9a593, 32'h429c6a28, 32'h42889a09, 32'h424effa5};
test_output[7216:7223] = '{32'h40daf1be, 32'h41929660, 32'h0, 32'h0, 32'h0, 32'h429c6a28, 32'h42889a09, 32'h424effa5};
test_input[7224:7231] = '{32'hc1a443a1, 32'hc272cad1, 32'hc27b36a3, 32'h42417429, 32'h42c0f640, 32'hc0d99959, 32'h426d5620, 32'h4270b3d9};
test_output[7224:7231] = '{32'h0, 32'h0, 32'h0, 32'h42417429, 32'h42c0f640, 32'h0, 32'h426d5620, 32'h4270b3d9};
test_input[7232:7239] = '{32'h425c70b0, 32'h42c2f05f, 32'hc25ea3dc, 32'h419fcec2, 32'hc2b808db, 32'h40b60126, 32'h42bcfaa8, 32'hc2961ba7};
test_output[7232:7239] = '{32'h425c70b0, 32'h42c2f05f, 32'h0, 32'h419fcec2, 32'h0, 32'h40b60126, 32'h42bcfaa8, 32'h0};
test_input[7240:7247] = '{32'hc03d6dd7, 32'h41dffe7d, 32'hc1119fcc, 32'h42bce6c5, 32'hc29d3707, 32'hc2a7138b, 32'h4122c605, 32'h4297b14f};
test_output[7240:7247] = '{32'h0, 32'h41dffe7d, 32'h0, 32'h42bce6c5, 32'h0, 32'h0, 32'h4122c605, 32'h4297b14f};
test_input[7248:7255] = '{32'hc2a557b1, 32'hc22fa205, 32'h418b9815, 32'hc20f734b, 32'hc29cc11a, 32'h42c4ec23, 32'hc2bff3f9, 32'h41c546c7};
test_output[7248:7255] = '{32'h0, 32'h0, 32'h418b9815, 32'h0, 32'h0, 32'h42c4ec23, 32'h0, 32'h41c546c7};
test_input[7256:7263] = '{32'hc2799aba, 32'hc274b51d, 32'hc190a805, 32'h42ba228c, 32'hc228de6f, 32'h422db0a5, 32'h41520590, 32'h42b2c0e9};
test_output[7256:7263] = '{32'h0, 32'h0, 32'h0, 32'h42ba228c, 32'h0, 32'h422db0a5, 32'h41520590, 32'h42b2c0e9};
test_input[7264:7271] = '{32'h42227feb, 32'hc21a7f0f, 32'h4277797a, 32'hc2c770d0, 32'h42c1df2f, 32'h40c004f2, 32'h419a0e8f, 32'hc24a1a53};
test_output[7264:7271] = '{32'h42227feb, 32'h0, 32'h4277797a, 32'h0, 32'h42c1df2f, 32'h40c004f2, 32'h419a0e8f, 32'h0};
test_input[7272:7279] = '{32'h4225fbeb, 32'hbe652355, 32'h42811407, 32'hc26885cd, 32'hc0b31da7, 32'hc27f2b70, 32'hc223f70a, 32'hc1a0a771};
test_output[7272:7279] = '{32'h4225fbeb, 32'h0, 32'h42811407, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7280:7287] = '{32'h40cfd47d, 32'h41a532f6, 32'h411fa7be, 32'hc1ff5dbc, 32'h4233c5a4, 32'h428ee38b, 32'hc243a17e, 32'hc23ed67d};
test_output[7280:7287] = '{32'h40cfd47d, 32'h41a532f6, 32'h411fa7be, 32'h0, 32'h4233c5a4, 32'h428ee38b, 32'h0, 32'h0};
test_input[7288:7295] = '{32'hc19fe69c, 32'h42830995, 32'hc1cddfb6, 32'h42a02399, 32'hc2b2483a, 32'h41679ff2, 32'hc1575b1d, 32'h4285c644};
test_output[7288:7295] = '{32'h0, 32'h42830995, 32'h0, 32'h42a02399, 32'h0, 32'h41679ff2, 32'h0, 32'h4285c644};
test_input[7296:7303] = '{32'hc1a08d72, 32'hc287f8e8, 32'hc280f66b, 32'hc2c4df11, 32'hc1119a29, 32'h3fbfe26b, 32'hc2b756a7, 32'h42c6e2d7};
test_output[7296:7303] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3fbfe26b, 32'h0, 32'h42c6e2d7};
test_input[7304:7311] = '{32'hc2b53aa3, 32'hc278f9a9, 32'hc166b0e2, 32'h410f29d3, 32'h42a9102d, 32'hc1dca1f7, 32'hc18a9d27, 32'h41f3f51a};
test_output[7304:7311] = '{32'h0, 32'h0, 32'h0, 32'h410f29d3, 32'h42a9102d, 32'h0, 32'h0, 32'h41f3f51a};
test_input[7312:7319] = '{32'h419aa629, 32'h41b9f171, 32'h4120554c, 32'h42ab63bd, 32'h41b6fb0c, 32'h4299c8ed, 32'hc136af51, 32'hbf4d8aae};
test_output[7312:7319] = '{32'h419aa629, 32'h41b9f171, 32'h4120554c, 32'h42ab63bd, 32'h41b6fb0c, 32'h4299c8ed, 32'h0, 32'h0};
test_input[7320:7327] = '{32'hc2a93935, 32'hc29f8d48, 32'h41c01878, 32'hc2be8c9a, 32'hc24d1ea6, 32'h418aaab3, 32'h41aee115, 32'hc00dd2cd};
test_output[7320:7327] = '{32'h0, 32'h0, 32'h41c01878, 32'h0, 32'h0, 32'h418aaab3, 32'h41aee115, 32'h0};
test_input[7328:7335] = '{32'h425c773d, 32'hc21bbec9, 32'h4251ca51, 32'hc25b907c, 32'h4234ec74, 32'h411a3ac9, 32'h422bac4a, 32'hc24520f5};
test_output[7328:7335] = '{32'h425c773d, 32'h0, 32'h4251ca51, 32'h0, 32'h4234ec74, 32'h411a3ac9, 32'h422bac4a, 32'h0};
test_input[7336:7343] = '{32'h4269f6ce, 32'h3f3c66ea, 32'hc2ad747d, 32'hc21270cd, 32'hc29510db, 32'hc2a94312, 32'hc2695e15, 32'h41dc7516};
test_output[7336:7343] = '{32'h4269f6ce, 32'h3f3c66ea, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41dc7516};
test_input[7344:7351] = '{32'h42c7dd55, 32'h4209664c, 32'hc2ad4fd2, 32'h420c6b01, 32'hc1cefbdf, 32'hc265c4ce, 32'hc24fbefe, 32'h41eea627};
test_output[7344:7351] = '{32'h42c7dd55, 32'h4209664c, 32'h0, 32'h420c6b01, 32'h0, 32'h0, 32'h0, 32'h41eea627};
test_input[7352:7359] = '{32'h40eef693, 32'h425cc149, 32'h429b0fb8, 32'hc2c41743, 32'hc0ee432c, 32'hc2b68d52, 32'hc21f1a77, 32'h4012c5a5};
test_output[7352:7359] = '{32'h40eef693, 32'h425cc149, 32'h429b0fb8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4012c5a5};
test_input[7360:7367] = '{32'h425f9adc, 32'h4138776c, 32'hc20f023a, 32'hc17ebf0c, 32'h4141ad4d, 32'hc2912aff, 32'hc22c85ba, 32'h42b6e3bb};
test_output[7360:7367] = '{32'h425f9adc, 32'h4138776c, 32'h0, 32'h0, 32'h4141ad4d, 32'h0, 32'h0, 32'h42b6e3bb};
test_input[7368:7375] = '{32'h42b23ffe, 32'h4195e592, 32'hc2317b73, 32'hc2192f2b, 32'h428db684, 32'hc2c4572f, 32'hc17e6c7b, 32'hc2c1094d};
test_output[7368:7375] = '{32'h42b23ffe, 32'h4195e592, 32'h0, 32'h0, 32'h428db684, 32'h0, 32'h0, 32'h0};
test_input[7376:7383] = '{32'hc2291f6d, 32'hc2c4258e, 32'hc2adac83, 32'hc296e64b, 32'hc244cfc0, 32'hc24571b8, 32'hc1e6df45, 32'hc1f82041};
test_output[7376:7383] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7384:7391] = '{32'hc19cc91e, 32'h4244deb2, 32'h42049139, 32'h40bdb0d9, 32'h428ac9e7, 32'h42294692, 32'hc28d381a, 32'h42046ab5};
test_output[7384:7391] = '{32'h0, 32'h4244deb2, 32'h42049139, 32'h40bdb0d9, 32'h428ac9e7, 32'h42294692, 32'h0, 32'h42046ab5};
test_input[7392:7399] = '{32'hc2b0228a, 32'hc2b41c00, 32'hbfdb511b, 32'hc2452170, 32'hc26989b7, 32'hc23f4f48, 32'h41f1e13a, 32'hc18a448c};
test_output[7392:7399] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f1e13a, 32'h0};
test_input[7400:7407] = '{32'h42c5b87a, 32'hc204cc26, 32'hc264cf85, 32'h429aa3e4, 32'hc12494fb, 32'hc27870a6, 32'hc2b30195, 32'h40f9765f};
test_output[7400:7407] = '{32'h42c5b87a, 32'h0, 32'h0, 32'h429aa3e4, 32'h0, 32'h0, 32'h0, 32'h40f9765f};
test_input[7408:7415] = '{32'hc100006e, 32'hc0f5254a, 32'h4260f519, 32'hc20d1c8f, 32'h423784ff, 32'h41b31bbf, 32'hc2b5034e, 32'hc254b4e0};
test_output[7408:7415] = '{32'h0, 32'h0, 32'h4260f519, 32'h0, 32'h423784ff, 32'h41b31bbf, 32'h0, 32'h0};
test_input[7416:7423] = '{32'hc2a73a4a, 32'hc27d5257, 32'hc27a3ad5, 32'hc293cce9, 32'h426f3c68, 32'h42a502f5, 32'hc2c4a52e, 32'hc18d5f55};
test_output[7416:7423] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h426f3c68, 32'h42a502f5, 32'h0, 32'h0};
test_input[7424:7431] = '{32'h42a6135d, 32'h4284453c, 32'h41d1490d, 32'hc20f705e, 32'hc1f9471d, 32'h4151c287, 32'hc17719fc, 32'hc2a2ec6a};
test_output[7424:7431] = '{32'h42a6135d, 32'h4284453c, 32'h41d1490d, 32'h0, 32'h0, 32'h4151c287, 32'h0, 32'h0};
test_input[7432:7439] = '{32'h418455cc, 32'h41cb33cf, 32'hc153860d, 32'h41949fd5, 32'hc2417d19, 32'h42901d15, 32'hc29d817e, 32'h41e22a62};
test_output[7432:7439] = '{32'h418455cc, 32'h41cb33cf, 32'h0, 32'h41949fd5, 32'h0, 32'h42901d15, 32'h0, 32'h41e22a62};
test_input[7440:7447] = '{32'h40ff71a5, 32'h422cbfc2, 32'hc2bfa8dc, 32'hc22643c0, 32'h41a65549, 32'hc18b5bcf, 32'hc25747b1, 32'h429373de};
test_output[7440:7447] = '{32'h40ff71a5, 32'h422cbfc2, 32'h0, 32'h0, 32'h41a65549, 32'h0, 32'h0, 32'h429373de};
test_input[7448:7455] = '{32'h42a10ccc, 32'h42a87a0e, 32'hc27789d9, 32'h429af775, 32'h42889747, 32'hc20a7c83, 32'h42747fde, 32'hc282e6e0};
test_output[7448:7455] = '{32'h42a10ccc, 32'h42a87a0e, 32'h0, 32'h429af775, 32'h42889747, 32'h0, 32'h42747fde, 32'h0};
test_input[7456:7463] = '{32'hc1494b6c, 32'h42a1235f, 32'hc11366c4, 32'h42ad1500, 32'h4212c476, 32'h4297860b, 32'h42aa4084, 32'h408c8587};
test_output[7456:7463] = '{32'h0, 32'h42a1235f, 32'h0, 32'h42ad1500, 32'h4212c476, 32'h4297860b, 32'h42aa4084, 32'h408c8587};
test_input[7464:7471] = '{32'h41a09c70, 32'hc255bbc7, 32'hc219f42c, 32'hc2bf07dc, 32'h41f7c649, 32'h41847603, 32'h4201e964, 32'hc27063f5};
test_output[7464:7471] = '{32'h41a09c70, 32'h0, 32'h0, 32'h0, 32'h41f7c649, 32'h41847603, 32'h4201e964, 32'h0};
test_input[7472:7479] = '{32'hc2a82073, 32'hc25eecd8, 32'h418e7429, 32'hc268d3f2, 32'hc27fa9e7, 32'hc2500193, 32'hc1935764, 32'h4249c060};
test_output[7472:7479] = '{32'h0, 32'h0, 32'h418e7429, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4249c060};
test_input[7480:7487] = '{32'hc24e81c1, 32'hc25e5589, 32'hc2834794, 32'h42bf75d6, 32'hc0bd6f02, 32'h40338d0b, 32'h3fe64fb6, 32'h4279dd7e};
test_output[7480:7487] = '{32'h0, 32'h0, 32'h0, 32'h42bf75d6, 32'h0, 32'h40338d0b, 32'h3fe64fb6, 32'h4279dd7e};
test_input[7488:7495] = '{32'h41bc2a99, 32'h4215c2d8, 32'h422668a5, 32'h41ada149, 32'hc27a3cc9, 32'h42bdfaa1, 32'hc29ac5e9, 32'h42a87dff};
test_output[7488:7495] = '{32'h41bc2a99, 32'h4215c2d8, 32'h422668a5, 32'h41ada149, 32'h0, 32'h42bdfaa1, 32'h0, 32'h42a87dff};
test_input[7496:7503] = '{32'h4292fd9a, 32'hbf16bfc8, 32'hc2beafe0, 32'hc2b18f50, 32'hc2a8d9b8, 32'h424d927d, 32'hc2c7a77a, 32'hc209d877};
test_output[7496:7503] = '{32'h4292fd9a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h424d927d, 32'h0, 32'h0};
test_input[7504:7511] = '{32'hc2b3970d, 32'h40e9ab56, 32'hc1a7de07, 32'hc0d24109, 32'hc2854f9d, 32'hc2996251, 32'hc2a35106, 32'h41c59f84};
test_output[7504:7511] = '{32'h0, 32'h40e9ab56, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41c59f84};
test_input[7512:7519] = '{32'hc1ede585, 32'h42327a62, 32'hc2880e20, 32'h412d7809, 32'h42b42f3e, 32'h4119489b, 32'hc2bfd697, 32'h3fdb8d63};
test_output[7512:7519] = '{32'h0, 32'h42327a62, 32'h0, 32'h412d7809, 32'h42b42f3e, 32'h4119489b, 32'h0, 32'h3fdb8d63};
test_input[7520:7527] = '{32'h426d7494, 32'h420f6f2b, 32'hc2053fc3, 32'h4234499d, 32'hc29f2756, 32'h410d38c9, 32'hc039c2e6, 32'h4296e338};
test_output[7520:7527] = '{32'h426d7494, 32'h420f6f2b, 32'h0, 32'h4234499d, 32'h0, 32'h410d38c9, 32'h0, 32'h4296e338};
test_input[7528:7535] = '{32'h409fd4fb, 32'hc26fe564, 32'h428de2b2, 32'h41fcc5dd, 32'hbe4e0567, 32'hc125aa80, 32'hc20594db, 32'hc25010cb};
test_output[7528:7535] = '{32'h409fd4fb, 32'h0, 32'h428de2b2, 32'h41fcc5dd, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7536:7543] = '{32'hc25c2750, 32'hc1bb202a, 32'hc2a1eb78, 32'hc21282b2, 32'h41bccb12, 32'hbe320d12, 32'h41b02fde, 32'hc195a5bf};
test_output[7536:7543] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41bccb12, 32'h0, 32'h41b02fde, 32'h0};
test_input[7544:7551] = '{32'hc24e01ba, 32'h41f20624, 32'hc2447484, 32'h42afcde6, 32'hc2040bc2, 32'h42424115, 32'hc2939caf, 32'hc25e5c2e};
test_output[7544:7551] = '{32'h0, 32'h41f20624, 32'h0, 32'h42afcde6, 32'h0, 32'h42424115, 32'h0, 32'h0};
test_input[7552:7559] = '{32'hc2b5c8ba, 32'hc27e43de, 32'h426b8063, 32'hc2c515b7, 32'h42a5666f, 32'hc2199334, 32'h42a8d535, 32'hc2bc65b3};
test_output[7552:7559] = '{32'h0, 32'h0, 32'h426b8063, 32'h0, 32'h42a5666f, 32'h0, 32'h42a8d535, 32'h0};
test_input[7560:7567] = '{32'hc117f820, 32'h42857d8d, 32'h42877f56, 32'h428ede80, 32'h42a7b647, 32'hc1e80cbe, 32'hc2c0a4b7, 32'hc113dff5};
test_output[7560:7567] = '{32'h0, 32'h42857d8d, 32'h42877f56, 32'h428ede80, 32'h42a7b647, 32'h0, 32'h0, 32'h0};
test_input[7568:7575] = '{32'h42840d0e, 32'hc2b53484, 32'h4206249c, 32'h41db1b38, 32'h4295da3c, 32'h42b9bec0, 32'h42c081cd, 32'hbfbffd2b};
test_output[7568:7575] = '{32'h42840d0e, 32'h0, 32'h4206249c, 32'h41db1b38, 32'h4295da3c, 32'h42b9bec0, 32'h42c081cd, 32'h0};
test_input[7576:7583] = '{32'hbfbe5648, 32'h4288d081, 32'h4296fa74, 32'h427fcdec, 32'hc1821d5d, 32'hc28c4486, 32'hc24c2a4e, 32'h4234c911};
test_output[7576:7583] = '{32'h0, 32'h4288d081, 32'h4296fa74, 32'h427fcdec, 32'h0, 32'h0, 32'h0, 32'h4234c911};
test_input[7584:7591] = '{32'h422c7573, 32'hc2ad3992, 32'h427c7dae, 32'h411141a2, 32'hc1224833, 32'h42701a63, 32'h421b4f8d, 32'h42c70181};
test_output[7584:7591] = '{32'h422c7573, 32'h0, 32'h427c7dae, 32'h411141a2, 32'h0, 32'h42701a63, 32'h421b4f8d, 32'h42c70181};
test_input[7592:7599] = '{32'hc232f4c5, 32'h4269488a, 32'hc2acda40, 32'hc21830fd, 32'hc1e257b3, 32'h42255587, 32'h42940c58, 32'h3f3daf66};
test_output[7592:7599] = '{32'h0, 32'h4269488a, 32'h0, 32'h0, 32'h0, 32'h42255587, 32'h42940c58, 32'h3f3daf66};
test_input[7600:7607] = '{32'h429eec6b, 32'h4283627a, 32'h422cb549, 32'h428919a5, 32'hc2086538, 32'hc20e0e78, 32'h419e7696, 32'hc17a2203};
test_output[7600:7607] = '{32'h429eec6b, 32'h4283627a, 32'h422cb549, 32'h428919a5, 32'h0, 32'h0, 32'h419e7696, 32'h0};
test_input[7608:7615] = '{32'hc2319bb6, 32'h413c153c, 32'h408aee68, 32'h42c6b029, 32'hc2a4e3d1, 32'h3f8bf14c, 32'hc1edf8a2, 32'h41b0c0a3};
test_output[7608:7615] = '{32'h0, 32'h413c153c, 32'h408aee68, 32'h42c6b029, 32'h0, 32'h3f8bf14c, 32'h0, 32'h41b0c0a3};
test_input[7616:7623] = '{32'h4276c1c8, 32'h42b46483, 32'h42050085, 32'h42242779, 32'h41e76ac8, 32'hc2429734, 32'h42359feb, 32'h424c5d10};
test_output[7616:7623] = '{32'h4276c1c8, 32'h42b46483, 32'h42050085, 32'h42242779, 32'h41e76ac8, 32'h0, 32'h42359feb, 32'h424c5d10};
test_input[7624:7631] = '{32'hc2c6ba36, 32'hc1aa1ac4, 32'h4280ad33, 32'hc2969032, 32'h41d7976a, 32'hc26d7479, 32'hc29232be, 32'h41423e30};
test_output[7624:7631] = '{32'h0, 32'h0, 32'h4280ad33, 32'h0, 32'h41d7976a, 32'h0, 32'h0, 32'h41423e30};
test_input[7632:7639] = '{32'h426e015a, 32'h3fcc7f8c, 32'h42206678, 32'hc2a47a28, 32'h4272e9c7, 32'hc28aaca5, 32'hc2c71e57, 32'hc2902072};
test_output[7632:7639] = '{32'h426e015a, 32'h3fcc7f8c, 32'h42206678, 32'h0, 32'h4272e9c7, 32'h0, 32'h0, 32'h0};
test_input[7640:7647] = '{32'h3f5b5d4d, 32'hc28820f2, 32'h4258da3a, 32'hc2773a4a, 32'hc167c552, 32'hc2bb5ae6, 32'h40ff6339, 32'hc21e32e7};
test_output[7640:7647] = '{32'h3f5b5d4d, 32'h0, 32'h4258da3a, 32'h0, 32'h0, 32'h0, 32'h40ff6339, 32'h0};
test_input[7648:7655] = '{32'h42a1c6af, 32'h41b9a6d8, 32'hc2ae059b, 32'hc237adc9, 32'hc23865f8, 32'h42a151fa, 32'hbe873344, 32'h4213b730};
test_output[7648:7655] = '{32'h42a1c6af, 32'h41b9a6d8, 32'h0, 32'h0, 32'h0, 32'h42a151fa, 32'h0, 32'h4213b730};
test_input[7656:7663] = '{32'hc2b223e2, 32'h42aaa0cc, 32'hc1c8783a, 32'h42a219af, 32'hc2006ab4, 32'h41b49f82, 32'hbeeaaba8, 32'h42b87b61};
test_output[7656:7663] = '{32'h0, 32'h42aaa0cc, 32'h0, 32'h42a219af, 32'h0, 32'h41b49f82, 32'h0, 32'h42b87b61};
test_input[7664:7671] = '{32'hc2889bb3, 32'h42862be0, 32'hc2a68f52, 32'h4248fc6c, 32'hc2894ec4, 32'h41d88a39, 32'hc28a8f62, 32'hc0813aaa};
test_output[7664:7671] = '{32'h0, 32'h42862be0, 32'h0, 32'h4248fc6c, 32'h0, 32'h41d88a39, 32'h0, 32'h0};
test_input[7672:7679] = '{32'hc23fa0d2, 32'hc1f629a7, 32'hc2b50838, 32'h4286174b, 32'hc275c0f7, 32'h40a63257, 32'h422d4fb4, 32'h42418cb3};
test_output[7672:7679] = '{32'h0, 32'h0, 32'h0, 32'h4286174b, 32'h0, 32'h40a63257, 32'h422d4fb4, 32'h42418cb3};
test_input[7680:7687] = '{32'hc1175cfa, 32'h42c36016, 32'h42984659, 32'hc1160765, 32'hc195b2fb, 32'hc0c9c539, 32'hc27206bf, 32'hc125ca7d};
test_output[7680:7687] = '{32'h0, 32'h42c36016, 32'h42984659, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7688:7695] = '{32'h41cbd279, 32'h425fc5ac, 32'hc21e3715, 32'h4232704f, 32'h42388150, 32'h418c3dc3, 32'h42778a73, 32'hc2bf89a6};
test_output[7688:7695] = '{32'h41cbd279, 32'h425fc5ac, 32'h0, 32'h4232704f, 32'h42388150, 32'h418c3dc3, 32'h42778a73, 32'h0};
test_input[7696:7703] = '{32'h42a5d7be, 32'hc2a19fbc, 32'h41b1ad52, 32'hc22e314b, 32'hc23c62f3, 32'h42059423, 32'hc1b70a09, 32'hc29c7efb};
test_output[7696:7703] = '{32'h42a5d7be, 32'h0, 32'h41b1ad52, 32'h0, 32'h0, 32'h42059423, 32'h0, 32'h0};
test_input[7704:7711] = '{32'hc29ebef8, 32'hbf285bfe, 32'hc1846790, 32'h42adfd46, 32'hc281d07a, 32'hc10935f1, 32'hc0f43d3c, 32'h41afd92c};
test_output[7704:7711] = '{32'h0, 32'h0, 32'h0, 32'h42adfd46, 32'h0, 32'h0, 32'h0, 32'h41afd92c};
test_input[7712:7719] = '{32'hc287f868, 32'h428a2f55, 32'hc2bb016f, 32'h426aa2df, 32'hc215c41d, 32'h405417a9, 32'h42c5a035, 32'h42bf2c5b};
test_output[7712:7719] = '{32'h0, 32'h428a2f55, 32'h0, 32'h426aa2df, 32'h0, 32'h405417a9, 32'h42c5a035, 32'h42bf2c5b};
test_input[7720:7727] = '{32'hc2619abf, 32'hbfa8985f, 32'h428d4f4d, 32'h42207c10, 32'h42076a8e, 32'hc26e0e8b, 32'h42b3629a, 32'hc294b41e};
test_output[7720:7727] = '{32'h0, 32'h0, 32'h428d4f4d, 32'h42207c10, 32'h42076a8e, 32'h0, 32'h42b3629a, 32'h0};
test_input[7728:7735] = '{32'h41126cb3, 32'h4277c7bc, 32'h42983287, 32'hc1f4bcf0, 32'h4274d8ba, 32'h421eabc0, 32'h41a245f4, 32'hc1cda9d3};
test_output[7728:7735] = '{32'h41126cb3, 32'h4277c7bc, 32'h42983287, 32'h0, 32'h4274d8ba, 32'h421eabc0, 32'h41a245f4, 32'h0};
test_input[7736:7743] = '{32'h4233cd02, 32'hc2b4a02d, 32'hc2b76d86, 32'h415f5ea8, 32'h415c538c, 32'hc27c59e2, 32'hc2b99dcb, 32'hc279c5d3};
test_output[7736:7743] = '{32'h4233cd02, 32'h0, 32'h0, 32'h415f5ea8, 32'h415c538c, 32'h0, 32'h0, 32'h0};
test_input[7744:7751] = '{32'h419d07e6, 32'h410aeda4, 32'h41404f40, 32'h427d2bc5, 32'hc285ef20, 32'h427cf34d, 32'hc2bf9ff2, 32'h426e866d};
test_output[7744:7751] = '{32'h419d07e6, 32'h410aeda4, 32'h41404f40, 32'h427d2bc5, 32'h0, 32'h427cf34d, 32'h0, 32'h426e866d};
test_input[7752:7759] = '{32'h420cf830, 32'hc1211cc4, 32'h4226bfa0, 32'h41b968ab, 32'h42bccb65, 32'hc2963a2d, 32'h42071d6f, 32'hc0707ea9};
test_output[7752:7759] = '{32'h420cf830, 32'h0, 32'h4226bfa0, 32'h41b968ab, 32'h42bccb65, 32'h0, 32'h42071d6f, 32'h0};
test_input[7760:7767] = '{32'hc2c5ea3b, 32'h4244df52, 32'hc1ce5414, 32'hc11175c2, 32'h412d1057, 32'hc163ee29, 32'h422da6d8, 32'h418b978b};
test_output[7760:7767] = '{32'h0, 32'h4244df52, 32'h0, 32'h0, 32'h412d1057, 32'h0, 32'h422da6d8, 32'h418b978b};
test_input[7768:7775] = '{32'hc1c9bef3, 32'h4256b5e2, 32'hc0d0cca8, 32'hc11ac124, 32'h404df81d, 32'h41e05453, 32'h428c8eec, 32'h428e6975};
test_output[7768:7775] = '{32'h0, 32'h4256b5e2, 32'h0, 32'h0, 32'h404df81d, 32'h41e05453, 32'h428c8eec, 32'h428e6975};
test_input[7776:7783] = '{32'h41d419bf, 32'hc2a98545, 32'hc216a053, 32'hc2c6a598, 32'hc1088b5c, 32'h429feed9, 32'h4226e178, 32'hc2653e8c};
test_output[7776:7783] = '{32'h41d419bf, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429feed9, 32'h4226e178, 32'h0};
test_input[7784:7791] = '{32'hc24a0ff5, 32'h41f29134, 32'hc27fbe63, 32'h41f98cb8, 32'hc28bd990, 32'hc262724c, 32'hc16676a8, 32'hc224eeeb};
test_output[7784:7791] = '{32'h0, 32'h41f29134, 32'h0, 32'h41f98cb8, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7792:7799] = '{32'h4275d260, 32'h42bf031a, 32'hc2aadf89, 32'hbfb2b020, 32'hc2c6f71b, 32'hc1d9e1d6, 32'hc2672334, 32'hc29b9ddf};
test_output[7792:7799] = '{32'h4275d260, 32'h42bf031a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7800:7807] = '{32'h4238e1c7, 32'hc18dcc8a, 32'hc28da062, 32'hc1f945d9, 32'hc2c092e3, 32'hc29de597, 32'h41858b17, 32'hc29fd041};
test_output[7800:7807] = '{32'h4238e1c7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41858b17, 32'h0};
test_input[7808:7815] = '{32'h4132e9a1, 32'hc12b4e48, 32'hc2282d57, 32'h424a6a7d, 32'h41974d0c, 32'hc2035729, 32'h42b9e107, 32'h422e236d};
test_output[7808:7815] = '{32'h4132e9a1, 32'h0, 32'h0, 32'h424a6a7d, 32'h41974d0c, 32'h0, 32'h42b9e107, 32'h422e236d};
test_input[7816:7823] = '{32'hc287f901, 32'hc2bedbf6, 32'hc29e7c85, 32'h42736429, 32'h42243e23, 32'hc134626a, 32'hc28ee55e, 32'hc2344dba};
test_output[7816:7823] = '{32'h0, 32'h0, 32'h0, 32'h42736429, 32'h42243e23, 32'h0, 32'h0, 32'h0};
test_input[7824:7831] = '{32'hc29022da, 32'h4291b9dd, 32'hc20b1b40, 32'hc20d6d37, 32'h42b9d086, 32'h4259f42b, 32'h429303f7, 32'h4283aec2};
test_output[7824:7831] = '{32'h0, 32'h4291b9dd, 32'h0, 32'h0, 32'h42b9d086, 32'h4259f42b, 32'h429303f7, 32'h4283aec2};
test_input[7832:7839] = '{32'h41df29d9, 32'hc264eaa6, 32'hc27bdfe9, 32'hc291b7b2, 32'hc238093a, 32'h419326c4, 32'h41b5efcd, 32'h41fe06d6};
test_output[7832:7839] = '{32'h41df29d9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h419326c4, 32'h41b5efcd, 32'h41fe06d6};
test_input[7840:7847] = '{32'h4165c739, 32'h428af9ba, 32'hc26805a0, 32'hc25499cc, 32'hc28f177b, 32'h42a9ee26, 32'hc12b2bbe, 32'h424bc16d};
test_output[7840:7847] = '{32'h4165c739, 32'h428af9ba, 32'h0, 32'h0, 32'h0, 32'h42a9ee26, 32'h0, 32'h424bc16d};
test_input[7848:7855] = '{32'hc2ad9405, 32'h423f251c, 32'hc2bc84f8, 32'h428a9ebb, 32'h42a35d89, 32'h4088bc54, 32'h41ab58be, 32'hc2512ebc};
test_output[7848:7855] = '{32'h0, 32'h423f251c, 32'h0, 32'h428a9ebb, 32'h42a35d89, 32'h4088bc54, 32'h41ab58be, 32'h0};
test_input[7856:7863] = '{32'h421ef719, 32'hc1d14ed4, 32'hc0ae99c0, 32'h41fb1995, 32'h42425d8b, 32'hc1c71bbb, 32'h41c1da12, 32'hc2c2c153};
test_output[7856:7863] = '{32'h421ef719, 32'h0, 32'h0, 32'h41fb1995, 32'h42425d8b, 32'h0, 32'h41c1da12, 32'h0};
test_input[7864:7871] = '{32'hc167da6d, 32'hc2b1383c, 32'hc2601daf, 32'h425dd050, 32'hc2c6d6e5, 32'hc2c2b9e6, 32'hbef91d5b, 32'hc25a8a88};
test_output[7864:7871] = '{32'h0, 32'h0, 32'h0, 32'h425dd050, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7872:7879] = '{32'hc237f879, 32'h414e4447, 32'h41ec7857, 32'h42333a91, 32'h42b5fefd, 32'h4275edc0, 32'h42687b98, 32'h418dc0a5};
test_output[7872:7879] = '{32'h0, 32'h414e4447, 32'h41ec7857, 32'h42333a91, 32'h42b5fefd, 32'h4275edc0, 32'h42687b98, 32'h418dc0a5};
test_input[7880:7887] = '{32'hc2b2f184, 32'h42a78fad, 32'hc24bfebf, 32'hc2b2ca9b, 32'h3fdcd5af, 32'hc20609eb, 32'h42a97214, 32'h41fbb465};
test_output[7880:7887] = '{32'h0, 32'h42a78fad, 32'h0, 32'h0, 32'h3fdcd5af, 32'h0, 32'h42a97214, 32'h41fbb465};
test_input[7888:7895] = '{32'h423ea17b, 32'hc245c09c, 32'h42aea6ea, 32'hc25e1eb1, 32'hc200b370, 32'hc2b44635, 32'hc18c38dc, 32'h41512cf9};
test_output[7888:7895] = '{32'h423ea17b, 32'h0, 32'h42aea6ea, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41512cf9};
test_input[7896:7903] = '{32'hc2826957, 32'hc147253e, 32'h42c13e90, 32'hc294dfd6, 32'hc2506649, 32'h424d1314, 32'h4281bb57, 32'hc292e3b7};
test_output[7896:7903] = '{32'h0, 32'h0, 32'h42c13e90, 32'h0, 32'h0, 32'h424d1314, 32'h4281bb57, 32'h0};
test_input[7904:7911] = '{32'h4280fe2b, 32'h428a24fb, 32'h41fcb020, 32'h42afc2b7, 32'hc2608cde, 32'h421e831e, 32'hc1b64c5d, 32'hc28d990d};
test_output[7904:7911] = '{32'h4280fe2b, 32'h428a24fb, 32'h41fcb020, 32'h42afc2b7, 32'h0, 32'h421e831e, 32'h0, 32'h0};
test_input[7912:7919] = '{32'hc2039682, 32'hc1c48acc, 32'h428b3566, 32'h40d2c4a3, 32'h40bd4ab2, 32'h42b5c478, 32'hc29eca87, 32'hc113cbe5};
test_output[7912:7919] = '{32'h0, 32'h0, 32'h428b3566, 32'h40d2c4a3, 32'h40bd4ab2, 32'h42b5c478, 32'h0, 32'h0};
test_input[7920:7927] = '{32'hc19b26cc, 32'hc201ba91, 32'h42b2c701, 32'hc2a2273a, 32'h42a77a7a, 32'hc21ed38d, 32'h42872e4e, 32'hc13ba90a};
test_output[7920:7927] = '{32'h0, 32'h0, 32'h42b2c701, 32'h0, 32'h42a77a7a, 32'h0, 32'h42872e4e, 32'h0};
test_input[7928:7935] = '{32'hc2b1aeb7, 32'h416a8708, 32'h42ae8f77, 32'hc26aaf66, 32'hc28201ce, 32'hc211d061, 32'hc17d1519, 32'hc2b7214a};
test_output[7928:7935] = '{32'h0, 32'h416a8708, 32'h42ae8f77, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7936:7943] = '{32'hc2a5c9f6, 32'hc22eef5e, 32'h42a3c797, 32'hc2b42804, 32'hc26d1fd6, 32'hc0ae4d2c, 32'h41b32376, 32'hc2394047};
test_output[7936:7943] = '{32'h0, 32'h0, 32'h42a3c797, 32'h0, 32'h0, 32'h0, 32'h41b32376, 32'h0};
test_input[7944:7951] = '{32'hc2aa9375, 32'hc2aa1375, 32'h42353153, 32'h41b273aa, 32'h428e83e1, 32'hc0e6e6e4, 32'hc19feff3, 32'h419a6129};
test_output[7944:7951] = '{32'h0, 32'h0, 32'h42353153, 32'h41b273aa, 32'h428e83e1, 32'h0, 32'h0, 32'h419a6129};
test_input[7952:7959] = '{32'h42a2ca42, 32'hc20bb717, 32'hc17d2104, 32'hc293e3d3, 32'hc2ba7ddc, 32'h42858122, 32'hc1d4a81f, 32'hc207c16e};
test_output[7952:7959] = '{32'h42a2ca42, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42858122, 32'h0, 32'h0};
test_input[7960:7967] = '{32'h4217491f, 32'hc2c2d876, 32'hc213130c, 32'hc2952c15, 32'hc24cea52, 32'hc1a8187c, 32'h425c7d1d, 32'hc2c4ee4b};
test_output[7960:7967] = '{32'h4217491f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425c7d1d, 32'h0};
test_input[7968:7975] = '{32'hc2900329, 32'h42ab71fd, 32'h4281e49f, 32'hc202b38f, 32'h42730732, 32'hc213db0f, 32'hc2bea732, 32'hc204938d};
test_output[7968:7975] = '{32'h0, 32'h42ab71fd, 32'h4281e49f, 32'h0, 32'h42730732, 32'h0, 32'h0, 32'h0};
test_input[7976:7983] = '{32'h418ac925, 32'h420daa87, 32'h4290e2d2, 32'h422c18ec, 32'hc2bf1a3c, 32'hc2835ef8, 32'hc28fd409, 32'h3fbc8cfb};
test_output[7976:7983] = '{32'h418ac925, 32'h420daa87, 32'h4290e2d2, 32'h422c18ec, 32'h0, 32'h0, 32'h0, 32'h3fbc8cfb};
test_input[7984:7991] = '{32'hc275e6f3, 32'h429d4e25, 32'hc228fb4d, 32'hc2a894bd, 32'h4259cbef, 32'h41b43ed0, 32'h41d343ff, 32'h40a4567a};
test_output[7984:7991] = '{32'h0, 32'h429d4e25, 32'h0, 32'h0, 32'h4259cbef, 32'h41b43ed0, 32'h41d343ff, 32'h40a4567a};
test_input[7992:7999] = '{32'h428456c0, 32'hc22e787c, 32'hc1a5cfff, 32'h422411b2, 32'hc287b6ef, 32'h40a23cfc, 32'hc29d9618, 32'hc2925b31};
test_output[7992:7999] = '{32'h428456c0, 32'h0, 32'h0, 32'h422411b2, 32'h0, 32'h40a23cfc, 32'h0, 32'h0};
test_input[8000:8007] = '{32'hc10ad292, 32'h41cfec62, 32'hc2054206, 32'h406a1b4b, 32'h42288819, 32'h42b04cfc, 32'h42165cf6, 32'hc10752bb};
test_output[8000:8007] = '{32'h0, 32'h41cfec62, 32'h0, 32'h406a1b4b, 32'h42288819, 32'h42b04cfc, 32'h42165cf6, 32'h0};
test_input[8008:8015] = '{32'h411dc7c9, 32'hc29dc4e3, 32'h42867695, 32'h41e05ea3, 32'hc2ae17bb, 32'h42738e9e, 32'h42898c06, 32'hc169f548};
test_output[8008:8015] = '{32'h411dc7c9, 32'h0, 32'h42867695, 32'h41e05ea3, 32'h0, 32'h42738e9e, 32'h42898c06, 32'h0};
test_input[8016:8023] = '{32'h424da31d, 32'h40ab638d, 32'hc288f38d, 32'h42236786, 32'h429173ae, 32'hc2bee9f1, 32'hc2bd80b0, 32'h42ab5d41};
test_output[8016:8023] = '{32'h424da31d, 32'h40ab638d, 32'h0, 32'h42236786, 32'h429173ae, 32'h0, 32'h0, 32'h42ab5d41};
test_input[8024:8031] = '{32'hc2be6fca, 32'h42990f8c, 32'hc20f3253, 32'h42318aee, 32'h42891f06, 32'h42a2127c, 32'h41949019, 32'h41fd374a};
test_output[8024:8031] = '{32'h0, 32'h42990f8c, 32'h0, 32'h42318aee, 32'h42891f06, 32'h42a2127c, 32'h41949019, 32'h41fd374a};
test_input[8032:8039] = '{32'h4231dbe9, 32'hc295a39b, 32'hc2441149, 32'h42c7d19b, 32'h40c9ab0f, 32'h429d0584, 32'hc2bfaa56, 32'h42671781};
test_output[8032:8039] = '{32'h4231dbe9, 32'h0, 32'h0, 32'h42c7d19b, 32'h40c9ab0f, 32'h429d0584, 32'h0, 32'h42671781};
test_input[8040:8047] = '{32'hc2090749, 32'hc19cc944, 32'h4295c1d0, 32'h4292df4b, 32'hc2a90b94, 32'hc2180b9e, 32'h418d8ac0, 32'hc21303c7};
test_output[8040:8047] = '{32'h0, 32'h0, 32'h4295c1d0, 32'h4292df4b, 32'h0, 32'h0, 32'h418d8ac0, 32'h0};
test_input[8048:8055] = '{32'hc2b9bb6c, 32'hc2309a54, 32'hc22cd9eb, 32'hc276d727, 32'hc1fc8c5a, 32'hc203121d, 32'h4279661b, 32'h42076ab6};
test_output[8048:8055] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4279661b, 32'h42076ab6};
test_input[8056:8063] = '{32'hc20bad27, 32'hc014d3df, 32'hc2a71f48, 32'hc2a616de, 32'h414bed1b, 32'hc29b6c15, 32'hc20a46e2, 32'h41115cb6};
test_output[8056:8063] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h414bed1b, 32'h0, 32'h0, 32'h41115cb6};
test_input[8064:8071] = '{32'hc1e8a3ee, 32'hc2976fca, 32'hc1b97624, 32'hc298ef45, 32'h422c3e11, 32'h4269c9ed, 32'hc205ce7f, 32'h41f86e37};
test_output[8064:8071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h422c3e11, 32'h4269c9ed, 32'h0, 32'h41f86e37};
test_input[8072:8079] = '{32'h424341da, 32'hc1fbc95c, 32'hc28a61e7, 32'hc23529a8, 32'hc212e688, 32'hc191214a, 32'hc28e0fbc, 32'hc127ff2b};
test_output[8072:8079] = '{32'h424341da, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8080:8087] = '{32'hc284e38e, 32'h42813188, 32'hc24a12c3, 32'h41b68c42, 32'hc2939efd, 32'hc02367f2, 32'hc26d883a, 32'h42863ce1};
test_output[8080:8087] = '{32'h0, 32'h42813188, 32'h0, 32'h41b68c42, 32'h0, 32'h0, 32'h0, 32'h42863ce1};
test_input[8088:8095] = '{32'hc2519879, 32'h42ab7cc0, 32'h42aa6669, 32'h4283c83a, 32'hc118a6e1, 32'hc214654b, 32'hc1901755, 32'hc2b729e6};
test_output[8088:8095] = '{32'h0, 32'h42ab7cc0, 32'h42aa6669, 32'h4283c83a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8096:8103] = '{32'h42bb7965, 32'h42b531b4, 32'h4187af08, 32'h42b444d6, 32'h4128eeff, 32'hc28d23dc, 32'hc26be3fa, 32'h42ba2421};
test_output[8096:8103] = '{32'h42bb7965, 32'h42b531b4, 32'h4187af08, 32'h42b444d6, 32'h4128eeff, 32'h0, 32'h0, 32'h42ba2421};
test_input[8104:8111] = '{32'h426a2120, 32'h4288ca3a, 32'hc2adb53f, 32'h413a2971, 32'h41ccd06d, 32'hc2bd39cc, 32'h40b55a39, 32'hc2903661};
test_output[8104:8111] = '{32'h426a2120, 32'h4288ca3a, 32'h0, 32'h413a2971, 32'h41ccd06d, 32'h0, 32'h40b55a39, 32'h0};
test_input[8112:8119] = '{32'hc29904fd, 32'hc2b55cd7, 32'h429a1859, 32'h42bc1119, 32'hc13fce0c, 32'hc215abb6, 32'h425884a5, 32'hc2661d71};
test_output[8112:8119] = '{32'h0, 32'h0, 32'h429a1859, 32'h42bc1119, 32'h0, 32'h0, 32'h425884a5, 32'h0};
test_input[8120:8127] = '{32'h4065ed62, 32'hc294f9f8, 32'h42a54ed1, 32'hc28d37ef, 32'h41ed7ff2, 32'h42c28d19, 32'h41ab7516, 32'h427e1bf8};
test_output[8120:8127] = '{32'h4065ed62, 32'h0, 32'h42a54ed1, 32'h0, 32'h41ed7ff2, 32'h42c28d19, 32'h41ab7516, 32'h427e1bf8};
test_input[8128:8135] = '{32'hc2564e08, 32'h42539a84, 32'h428df39a, 32'h429d9d88, 32'h42b2e465, 32'h42123ce0, 32'h411986e5, 32'hc1d3596a};
test_output[8128:8135] = '{32'h0, 32'h42539a84, 32'h428df39a, 32'h429d9d88, 32'h42b2e465, 32'h42123ce0, 32'h411986e5, 32'h0};
test_input[8136:8143] = '{32'h420830cd, 32'hc1e9c933, 32'h412b3de2, 32'h428e3384, 32'h428bfa68, 32'h429920ae, 32'h42c16a33, 32'hc299a484};
test_output[8136:8143] = '{32'h420830cd, 32'h0, 32'h412b3de2, 32'h428e3384, 32'h428bfa68, 32'h429920ae, 32'h42c16a33, 32'h0};
test_input[8144:8151] = '{32'h42020b80, 32'h4217ab95, 32'h422409e4, 32'hc21e4c42, 32'h42953e85, 32'h41703637, 32'hc21a40f3, 32'h42030021};
test_output[8144:8151] = '{32'h42020b80, 32'h4217ab95, 32'h422409e4, 32'h0, 32'h42953e85, 32'h41703637, 32'h0, 32'h42030021};
test_input[8152:8159] = '{32'hc216206c, 32'h41be8fae, 32'hc28dfddb, 32'h42b44e6d, 32'h423d7ef3, 32'h41e5c5b8, 32'h41db7380, 32'hc25160e2};
test_output[8152:8159] = '{32'h0, 32'h41be8fae, 32'h0, 32'h42b44e6d, 32'h423d7ef3, 32'h41e5c5b8, 32'h41db7380, 32'h0};
test_input[8160:8167] = '{32'hc2b82e0a, 32'hc2b8bda4, 32'h42675fd3, 32'h42a84975, 32'h42b2373f, 32'h41fe990e, 32'hc1aa82ae, 32'h41a8b6a4};
test_output[8160:8167] = '{32'h0, 32'h0, 32'h42675fd3, 32'h42a84975, 32'h42b2373f, 32'h41fe990e, 32'h0, 32'h41a8b6a4};
test_input[8168:8175] = '{32'hc21b8a39, 32'h42906ccb, 32'hc1f0e7d4, 32'h410097af, 32'hc2959c22, 32'hc1e3d092, 32'hc2be2428, 32'h420bc5e9};
test_output[8168:8175] = '{32'h0, 32'h42906ccb, 32'h0, 32'h410097af, 32'h0, 32'h0, 32'h0, 32'h420bc5e9};
test_input[8176:8183] = '{32'hc1e3cf48, 32'h408139ec, 32'hc2c47526, 32'hc0f5b561, 32'hc2c2b14a, 32'hc2532d74, 32'hc1c043aa, 32'hc2af6a9f};
test_output[8176:8183] = '{32'h0, 32'h408139ec, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8184:8191] = '{32'hc2bc5d8b, 32'hc231fffe, 32'hc271b5d0, 32'h4058bc9d, 32'h3fbdf09e, 32'hc2692d19, 32'h4244f670, 32'hc2200a37};
test_output[8184:8191] = '{32'h0, 32'h0, 32'h0, 32'h4058bc9d, 32'h3fbdf09e, 32'h0, 32'h4244f670, 32'h0};
test_input[8192:8199] = '{32'hc2b696f4, 32'h4294859a, 32'hc2740346, 32'h41749f58, 32'h40404cb8, 32'h429162b9, 32'h425bd078, 32'h41867422};
test_output[8192:8199] = '{32'h0, 32'h4294859a, 32'h0, 32'h41749f58, 32'h40404cb8, 32'h429162b9, 32'h425bd078, 32'h41867422};
test_input[8200:8207] = '{32'hc2773c06, 32'h42b842bb, 32'hc26111eb, 32'h427c60ae, 32'hc22075c7, 32'hc0fb406d, 32'h42536333, 32'h42658f50};
test_output[8200:8207] = '{32'h0, 32'h42b842bb, 32'h0, 32'h427c60ae, 32'h0, 32'h0, 32'h42536333, 32'h42658f50};
test_input[8208:8215] = '{32'h428988e6, 32'h402be3e5, 32'h427d9ee2, 32'h40d8905b, 32'hbfe30348, 32'hc2aaae1e, 32'hc25a6310, 32'hc2a63d14};
test_output[8208:8215] = '{32'h428988e6, 32'h402be3e5, 32'h427d9ee2, 32'h40d8905b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8216:8223] = '{32'h42b0016c, 32'h42b3e3ab, 32'hc2a11912, 32'h42ba1693, 32'h41ef6ef3, 32'h4280e540, 32'h428eebc0, 32'hc24e689a};
test_output[8216:8223] = '{32'h42b0016c, 32'h42b3e3ab, 32'h0, 32'h42ba1693, 32'h41ef6ef3, 32'h4280e540, 32'h428eebc0, 32'h0};
test_input[8224:8231] = '{32'h3d8ed8df, 32'h42a25cc1, 32'hc2c35536, 32'h428b621e, 32'hc2ae5fc1, 32'hc1b71996, 32'hc23d2e5c, 32'h42001215};
test_output[8224:8231] = '{32'h3d8ed8df, 32'h42a25cc1, 32'h0, 32'h428b621e, 32'h0, 32'h0, 32'h0, 32'h42001215};
test_input[8232:8239] = '{32'hc24a9fd7, 32'h4260f7ae, 32'hc2b5964c, 32'hc1f3563a, 32'h424305ae, 32'h42c72de3, 32'h428063c0, 32'h425a506b};
test_output[8232:8239] = '{32'h0, 32'h4260f7ae, 32'h0, 32'h0, 32'h424305ae, 32'h42c72de3, 32'h428063c0, 32'h425a506b};
test_input[8240:8247] = '{32'h4217e312, 32'hc22d98cc, 32'h41dc90ce, 32'hc2810213, 32'h428f9f4c, 32'h429df62b, 32'hc219956c, 32'h409c4340};
test_output[8240:8247] = '{32'h4217e312, 32'h0, 32'h41dc90ce, 32'h0, 32'h428f9f4c, 32'h429df62b, 32'h0, 32'h409c4340};
test_input[8248:8255] = '{32'h4093428d, 32'h42205b93, 32'h41b265e2, 32'h41dd3cb1, 32'h42a2fea5, 32'hc2b820bf, 32'h426456d1, 32'h42784be5};
test_output[8248:8255] = '{32'h4093428d, 32'h42205b93, 32'h41b265e2, 32'h41dd3cb1, 32'h42a2fea5, 32'h0, 32'h426456d1, 32'h42784be5};
test_input[8256:8263] = '{32'h4252204d, 32'h425b5ad9, 32'h42703efe, 32'h41c8841d, 32'hc199b3ec, 32'h42a94c00, 32'h42b61b95, 32'h42790c38};
test_output[8256:8263] = '{32'h4252204d, 32'h425b5ad9, 32'h42703efe, 32'h41c8841d, 32'h0, 32'h42a94c00, 32'h42b61b95, 32'h42790c38};
test_input[8264:8271] = '{32'hc2186899, 32'hbe7f9d44, 32'h42c7d714, 32'h421eed84, 32'h41ecfa42, 32'h423bde86, 32'h42058162, 32'hc24bdde0};
test_output[8264:8271] = '{32'h0, 32'h0, 32'h42c7d714, 32'h421eed84, 32'h41ecfa42, 32'h423bde86, 32'h42058162, 32'h0};
test_input[8272:8279] = '{32'h42809b2c, 32'hc2c499dd, 32'h428a4f03, 32'h42bdb0ac, 32'h42314775, 32'hc0e87781, 32'h424906d1, 32'h42b81527};
test_output[8272:8279] = '{32'h42809b2c, 32'h0, 32'h428a4f03, 32'h42bdb0ac, 32'h42314775, 32'h0, 32'h424906d1, 32'h42b81527};
test_input[8280:8287] = '{32'h42a514e0, 32'h41af4944, 32'hc24aba12, 32'hbfd6af2a, 32'h428852b6, 32'hc21e1e0d, 32'hc242e253, 32'hc1b11efd};
test_output[8280:8287] = '{32'h42a514e0, 32'h41af4944, 32'h0, 32'h0, 32'h428852b6, 32'h0, 32'h0, 32'h0};
test_input[8288:8295] = '{32'h42bb7ac6, 32'hc28a6639, 32'hc1ac1b59, 32'h42b7021f, 32'hc2867c69, 32'h417a8d54, 32'hc28d13da, 32'hc1c6b7a9};
test_output[8288:8295] = '{32'h42bb7ac6, 32'h0, 32'h0, 32'h42b7021f, 32'h0, 32'h417a8d54, 32'h0, 32'h0};
test_input[8296:8303] = '{32'h42c392b9, 32'hc2312b04, 32'h42b23a90, 32'hc2093dcd, 32'h42912cdb, 32'hc2ab82ec, 32'h4237b936, 32'hc204c6e9};
test_output[8296:8303] = '{32'h42c392b9, 32'h0, 32'h42b23a90, 32'h0, 32'h42912cdb, 32'h0, 32'h4237b936, 32'h0};
test_input[8304:8311] = '{32'h425a5ff1, 32'h429012be, 32'h4285fba1, 32'h409b4dd3, 32'hc1211780, 32'hc2ba85af, 32'h42a99ed3, 32'hc10b4ee6};
test_output[8304:8311] = '{32'h425a5ff1, 32'h429012be, 32'h4285fba1, 32'h409b4dd3, 32'h0, 32'h0, 32'h42a99ed3, 32'h0};
test_input[8312:8319] = '{32'hc22f33ff, 32'h4285f411, 32'hc079647b, 32'hc1da2182, 32'hc1a39a7f, 32'hc2360c96, 32'hc29fb014, 32'hc24566d5};
test_output[8312:8319] = '{32'h0, 32'h4285f411, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8320:8327] = '{32'h4182ac8b, 32'hc2ad897f, 32'hc2962157, 32'h4291c735, 32'h418117fd, 32'h42b065a8, 32'hc10b57bf, 32'h42a53d3f};
test_output[8320:8327] = '{32'h4182ac8b, 32'h0, 32'h0, 32'h4291c735, 32'h418117fd, 32'h42b065a8, 32'h0, 32'h42a53d3f};
test_input[8328:8335] = '{32'hc11b376d, 32'h42141b2e, 32'h41dabc06, 32'h424cd60c, 32'hc19947d4, 32'hc2c7619e, 32'hc03b624e, 32'hc283384b};
test_output[8328:8335] = '{32'h0, 32'h42141b2e, 32'h41dabc06, 32'h424cd60c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8336:8343] = '{32'h40df9af0, 32'h419684ec, 32'h408e953d, 32'h413e929d, 32'h42865c3a, 32'h428e51d9, 32'h41749cdf, 32'h42623493};
test_output[8336:8343] = '{32'h40df9af0, 32'h419684ec, 32'h408e953d, 32'h413e929d, 32'h42865c3a, 32'h428e51d9, 32'h41749cdf, 32'h42623493};
test_input[8344:8351] = '{32'h420b4703, 32'h42a9eb6f, 32'h422ba6a5, 32'hc1fdb148, 32'h4281d2e7, 32'h4281bd0f, 32'hc28631c2, 32'hc23b262c};
test_output[8344:8351] = '{32'h420b4703, 32'h42a9eb6f, 32'h422ba6a5, 32'h0, 32'h4281d2e7, 32'h4281bd0f, 32'h0, 32'h0};
test_input[8352:8359] = '{32'hc24fb051, 32'h426cae9d, 32'h42674bde, 32'h42981fbd, 32'h41d93824, 32'hc18cd80f, 32'hc2c42b23, 32'h4287d1da};
test_output[8352:8359] = '{32'h0, 32'h426cae9d, 32'h42674bde, 32'h42981fbd, 32'h41d93824, 32'h0, 32'h0, 32'h4287d1da};
test_input[8360:8367] = '{32'hc2705e9e, 32'hc1bd36d6, 32'h425d5f16, 32'hc288d082, 32'h426484ed, 32'hc21a67be, 32'h3fd714cb, 32'h42857195};
test_output[8360:8367] = '{32'h0, 32'h0, 32'h425d5f16, 32'h0, 32'h426484ed, 32'h0, 32'h3fd714cb, 32'h42857195};
test_input[8368:8375] = '{32'hc2b60dc6, 32'h4253f80a, 32'hc292b41f, 32'hc280e3da, 32'h42692a64, 32'h40cbe4b4, 32'hc2069d86, 32'hc19dbc7d};
test_output[8368:8375] = '{32'h0, 32'h4253f80a, 32'h0, 32'h0, 32'h42692a64, 32'h40cbe4b4, 32'h0, 32'h0};
test_input[8376:8383] = '{32'hc21b35bd, 32'h42c271ad, 32'h428c7b71, 32'hc1701594, 32'hc1af8b88, 32'hc26b474a, 32'hc29eeaf4, 32'hc2ac88fa};
test_output[8376:8383] = '{32'h0, 32'h42c271ad, 32'h428c7b71, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8384:8391] = '{32'hc2a0b64a, 32'hc1d2078a, 32'h409f2b3e, 32'hc2b09325, 32'hc28a47a8, 32'hc2138e4b, 32'hc27d86ad, 32'h423144f3};
test_output[8384:8391] = '{32'h0, 32'h0, 32'h409f2b3e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423144f3};
test_input[8392:8399] = '{32'hc27e099c, 32'hc26f57d9, 32'hc1cde84a, 32'h42767a38, 32'hc2b5469d, 32'hc1947d4a, 32'hc2a73c73, 32'h41b3988b};
test_output[8392:8399] = '{32'h0, 32'h0, 32'h0, 32'h42767a38, 32'h0, 32'h0, 32'h0, 32'h41b3988b};
test_input[8400:8407] = '{32'h42a1d785, 32'hc1d2fcd4, 32'hc2b8d0ea, 32'hc1cc49aa, 32'h42a83564, 32'h4111ba1c, 32'h420ea793, 32'h40b40b69};
test_output[8400:8407] = '{32'h42a1d785, 32'h0, 32'h0, 32'h0, 32'h42a83564, 32'h4111ba1c, 32'h420ea793, 32'h40b40b69};
test_input[8408:8415] = '{32'h42b16a7f, 32'h42199b65, 32'hc0d4d2e6, 32'hc2a231f6, 32'hc25f0278, 32'hc21c8c6b, 32'h41197bff, 32'h41096a84};
test_output[8408:8415] = '{32'h42b16a7f, 32'h42199b65, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41197bff, 32'h41096a84};
test_input[8416:8423] = '{32'h42a2908a, 32'hc2c7745f, 32'h4271565a, 32'hc27efd99, 32'hc285891f, 32'h422b0610, 32'h42a50e9d, 32'h4298f1dd};
test_output[8416:8423] = '{32'h42a2908a, 32'h0, 32'h4271565a, 32'h0, 32'h0, 32'h422b0610, 32'h42a50e9d, 32'h4298f1dd};
test_input[8424:8431] = '{32'hc0b32722, 32'hc2967225, 32'hc1dd283f, 32'hc118cedc, 32'h42c04c48, 32'hc2a282d3, 32'h41ea8430, 32'hc19118ec};
test_output[8424:8431] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42c04c48, 32'h0, 32'h41ea8430, 32'h0};
test_input[8432:8439] = '{32'h41df758c, 32'hc2bb2abb, 32'h428c5c9e, 32'h41cd61dd, 32'hc2565a15, 32'hc2993985, 32'hc2406ed3, 32'h41f75330};
test_output[8432:8439] = '{32'h41df758c, 32'h0, 32'h428c5c9e, 32'h41cd61dd, 32'h0, 32'h0, 32'h0, 32'h41f75330};
test_input[8440:8447] = '{32'hc1271e89, 32'h4296487b, 32'h423ac5fd, 32'hc2c1c4c1, 32'hc26fed86, 32'h420f3b9d, 32'hc2a96bed, 32'h4276e762};
test_output[8440:8447] = '{32'h0, 32'h4296487b, 32'h423ac5fd, 32'h0, 32'h0, 32'h420f3b9d, 32'h0, 32'h4276e762};
test_input[8448:8455] = '{32'h429f52cb, 32'h42ba576e, 32'h42938f50, 32'h41ac5184, 32'hc294cf7a, 32'h427bc3ea, 32'hc2888b6e, 32'h422b06e2};
test_output[8448:8455] = '{32'h429f52cb, 32'h42ba576e, 32'h42938f50, 32'h41ac5184, 32'h0, 32'h427bc3ea, 32'h0, 32'h422b06e2};
test_input[8456:8463] = '{32'hc161972b, 32'hc297a6ed, 32'h41f38580, 32'h428ed563, 32'hc2bd1861, 32'h420b789a, 32'h423d3c60, 32'hc0d2c734};
test_output[8456:8463] = '{32'h0, 32'h0, 32'h41f38580, 32'h428ed563, 32'h0, 32'h420b789a, 32'h423d3c60, 32'h0};
test_input[8464:8471] = '{32'hbfe5c254, 32'h4040115c, 32'hc239e2ab, 32'hc13cda4d, 32'h41c399db, 32'hc2a21a9c, 32'hc17650bf, 32'h41c6d0cf};
test_output[8464:8471] = '{32'h0, 32'h4040115c, 32'h0, 32'h0, 32'h41c399db, 32'h0, 32'h0, 32'h41c6d0cf};
test_input[8472:8479] = '{32'h42af064d, 32'h42395e55, 32'hc207ef5b, 32'hc2bad556, 32'hc1902da9, 32'hc25bd529, 32'hc21af5fb, 32'h42b9e089};
test_output[8472:8479] = '{32'h42af064d, 32'h42395e55, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b9e089};
test_input[8480:8487] = '{32'h427b85d2, 32'h42c48baf, 32'hc2bd43e8, 32'h413b1333, 32'h4266d1d5, 32'h42b5f6b4, 32'h41ce39ae, 32'h42532eb4};
test_output[8480:8487] = '{32'h427b85d2, 32'h42c48baf, 32'h0, 32'h413b1333, 32'h4266d1d5, 32'h42b5f6b4, 32'h41ce39ae, 32'h42532eb4};
test_input[8488:8495] = '{32'hc1a9ff3d, 32'h414aff10, 32'h400575cb, 32'h42936295, 32'hc24b0afb, 32'h42273c2a, 32'hc18cae38, 32'hc2ad6387};
test_output[8488:8495] = '{32'h0, 32'h414aff10, 32'h400575cb, 32'h42936295, 32'h0, 32'h42273c2a, 32'h0, 32'h0};
test_input[8496:8503] = '{32'h42a858d4, 32'h4299aeec, 32'h4250aa18, 32'hc257f32f, 32'h427e0f42, 32'hc1ba082e, 32'hc1b79fde, 32'hc0815ac1};
test_output[8496:8503] = '{32'h42a858d4, 32'h4299aeec, 32'h4250aa18, 32'h0, 32'h427e0f42, 32'h0, 32'h0, 32'h0};
test_input[8504:8511] = '{32'h42960d7e, 32'hc260a3b3, 32'hc1e7e0a6, 32'h428c7b8b, 32'h40de904a, 32'hc27cc589, 32'h42be75a4, 32'hc2530b4c};
test_output[8504:8511] = '{32'h42960d7e, 32'h0, 32'h0, 32'h428c7b8b, 32'h40de904a, 32'h0, 32'h42be75a4, 32'h0};
test_input[8512:8519] = '{32'hc1fd2adb, 32'hc214de8a, 32'h41a52b0c, 32'hc26e6147, 32'h42007356, 32'h427e0a7c, 32'hc1ec19f3, 32'hc1d0a296};
test_output[8512:8519] = '{32'h0, 32'h0, 32'h41a52b0c, 32'h0, 32'h42007356, 32'h427e0a7c, 32'h0, 32'h0};
test_input[8520:8527] = '{32'h3f568fc2, 32'h422d7a18, 32'hc2b48669, 32'h42b3e3a3, 32'h42ac0510, 32'h41635ccc, 32'h419c1a0c, 32'h42129f64};
test_output[8520:8527] = '{32'h3f568fc2, 32'h422d7a18, 32'h0, 32'h42b3e3a3, 32'h42ac0510, 32'h41635ccc, 32'h419c1a0c, 32'h42129f64};
test_input[8528:8535] = '{32'h42515518, 32'h41c858ba, 32'h4261efa6, 32'h41d92345, 32'h41ccab26, 32'hc2338ae0, 32'h428214bc, 32'hc1a691e4};
test_output[8528:8535] = '{32'h42515518, 32'h41c858ba, 32'h4261efa6, 32'h41d92345, 32'h41ccab26, 32'h0, 32'h428214bc, 32'h0};
test_input[8536:8543] = '{32'h42b3bc0a, 32'h3fdd15ff, 32'hc234e185, 32'h4198517d, 32'hc1eb783b, 32'hc12ca5b4, 32'h425e372a, 32'hc2a62b94};
test_output[8536:8543] = '{32'h42b3bc0a, 32'h3fdd15ff, 32'h0, 32'h4198517d, 32'h0, 32'h0, 32'h425e372a, 32'h0};
test_input[8544:8551] = '{32'hc293154b, 32'h41880e38, 32'h41b00046, 32'h42aafd9f, 32'hc2c0e7cf, 32'hc2807b6d, 32'hc221074b, 32'hc2a59cf9};
test_output[8544:8551] = '{32'h0, 32'h41880e38, 32'h41b00046, 32'h42aafd9f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8552:8559] = '{32'h42ad91f2, 32'hc2046a7d, 32'h42c5972b, 32'h41488f67, 32'hc27567e6, 32'h422162d6, 32'hc1a58d75, 32'hc28b1d7a};
test_output[8552:8559] = '{32'h42ad91f2, 32'h0, 32'h42c5972b, 32'h41488f67, 32'h0, 32'h422162d6, 32'h0, 32'h0};
test_input[8560:8567] = '{32'hc2930316, 32'h41237d44, 32'hc28cb098, 32'hc24bd62e, 32'hc2021be4, 32'hc2852c6f, 32'h40d6525c, 32'h41219550};
test_output[8560:8567] = '{32'h0, 32'h41237d44, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40d6525c, 32'h41219550};
test_input[8568:8575] = '{32'hc25a02fc, 32'h41e142d2, 32'hc29fc3ea, 32'hc2745fdb, 32'h41c5330d, 32'hc18b9997, 32'hc2046676, 32'hc20640bc};
test_output[8568:8575] = '{32'h0, 32'h41e142d2, 32'h0, 32'h0, 32'h41c5330d, 32'h0, 32'h0, 32'h0};
test_input[8576:8583] = '{32'hc201f3e0, 32'hc2117d89, 32'hc2b9a288, 32'h4169d6dc, 32'h42c445f8, 32'hc2b20b42, 32'hc27943d4, 32'hc24e39e5};
test_output[8576:8583] = '{32'h0, 32'h0, 32'h0, 32'h4169d6dc, 32'h42c445f8, 32'h0, 32'h0, 32'h0};
test_input[8584:8591] = '{32'hc121d191, 32'h407f6bb7, 32'hc171aafc, 32'hc28187c6, 32'hc2107158, 32'hc29fbc11, 32'h4298c77d, 32'h4265a314};
test_output[8584:8591] = '{32'h0, 32'h407f6bb7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4298c77d, 32'h4265a314};
test_input[8592:8599] = '{32'hc2559010, 32'h42c537b8, 32'hc1e5b4be, 32'h422244c8, 32'h41f9c344, 32'hbf925b21, 32'hc19620db, 32'h42bc0ca2};
test_output[8592:8599] = '{32'h0, 32'h42c537b8, 32'h0, 32'h422244c8, 32'h41f9c344, 32'h0, 32'h0, 32'h42bc0ca2};
test_input[8600:8607] = '{32'h4295952a, 32'h41cf1ee4, 32'h423361a8, 32'h42af6a29, 32'h402e116e, 32'hc29d6d99, 32'hc21d5adb, 32'h421db857};
test_output[8600:8607] = '{32'h4295952a, 32'h41cf1ee4, 32'h423361a8, 32'h42af6a29, 32'h402e116e, 32'h0, 32'h0, 32'h421db857};
test_input[8608:8615] = '{32'h41f495eb, 32'h4275572e, 32'hc2abbc1d, 32'hc0392513, 32'h424a2743, 32'h41933bdd, 32'hc2b51ec8, 32'hc21385ce};
test_output[8608:8615] = '{32'h41f495eb, 32'h4275572e, 32'h0, 32'h0, 32'h424a2743, 32'h41933bdd, 32'h0, 32'h0};
test_input[8616:8623] = '{32'hc2aae311, 32'h418d60c6, 32'hc282a31c, 32'hc193a782, 32'hc1ee6bc6, 32'h3fa9e156, 32'hc2bedf4e, 32'hc206f590};
test_output[8616:8623] = '{32'h0, 32'h418d60c6, 32'h0, 32'h0, 32'h0, 32'h3fa9e156, 32'h0, 32'h0};
test_input[8624:8631] = '{32'h417cf185, 32'hc297f2f1, 32'hc1fa73c6, 32'h421a6e51, 32'h40aadfc0, 32'hc2c358d6, 32'h4227f063, 32'h40e18fde};
test_output[8624:8631] = '{32'h417cf185, 32'h0, 32'h0, 32'h421a6e51, 32'h40aadfc0, 32'h0, 32'h4227f063, 32'h40e18fde};
test_input[8632:8639] = '{32'hc2ae1c9c, 32'hc231848b, 32'hc0dfb2bb, 32'hc1e298e2, 32'hc22b1fcd, 32'h426f80ee, 32'h42baae1f, 32'h42c420fe};
test_output[8632:8639] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426f80ee, 32'h42baae1f, 32'h42c420fe};
test_input[8640:8647] = '{32'hc2b49ea1, 32'hc229b524, 32'h424cf8d9, 32'h41ec58ac, 32'hc29f79f3, 32'hc17d8ce4, 32'hc299fac4, 32'h42abf7f4};
test_output[8640:8647] = '{32'h0, 32'h0, 32'h424cf8d9, 32'h41ec58ac, 32'h0, 32'h0, 32'h0, 32'h42abf7f4};
test_input[8648:8655] = '{32'hc1b9df52, 32'hc26ad677, 32'hc2b7852c, 32'hc27346af, 32'h42acadc3, 32'h415b6c81, 32'hc2941bf0, 32'h42b97a1a};
test_output[8648:8655] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42acadc3, 32'h415b6c81, 32'h0, 32'h42b97a1a};
test_input[8656:8663] = '{32'hc0acfc45, 32'h42bbcb74, 32'h40e0fd5f, 32'hc2b25e65, 32'hc197f0bd, 32'h42c245a3, 32'h42485ef2, 32'hc1ba309c};
test_output[8656:8663] = '{32'h0, 32'h42bbcb74, 32'h40e0fd5f, 32'h0, 32'h0, 32'h42c245a3, 32'h42485ef2, 32'h0};
test_input[8664:8671] = '{32'h4004861d, 32'hc0beb942, 32'h4223850b, 32'hc24a0073, 32'h417a79af, 32'hc22d0239, 32'h4125cdb5, 32'hc29345b3};
test_output[8664:8671] = '{32'h4004861d, 32'h0, 32'h4223850b, 32'h0, 32'h417a79af, 32'h0, 32'h4125cdb5, 32'h0};
test_input[8672:8679] = '{32'h423d0c22, 32'h42447f75, 32'h406daeba, 32'h42291660, 32'h408ae02d, 32'hc278be3d, 32'h3fdf4def, 32'h41e3b6d7};
test_output[8672:8679] = '{32'h423d0c22, 32'h42447f75, 32'h406daeba, 32'h42291660, 32'h408ae02d, 32'h0, 32'h3fdf4def, 32'h41e3b6d7};
test_input[8680:8687] = '{32'hc22ebb67, 32'h42be2f8b, 32'hc1606046, 32'h42b54597, 32'hc29f0958, 32'hc24d4e67, 32'h41ea21e4, 32'hc2154336};
test_output[8680:8687] = '{32'h0, 32'h42be2f8b, 32'h0, 32'h42b54597, 32'h0, 32'h0, 32'h41ea21e4, 32'h0};
test_input[8688:8695] = '{32'hc20535a9, 32'hc2634391, 32'h4150c1dd, 32'h4180c234, 32'h42b9af2b, 32'h418f3bd0, 32'h42094637, 32'h42856f87};
test_output[8688:8695] = '{32'h0, 32'h0, 32'h4150c1dd, 32'h4180c234, 32'h42b9af2b, 32'h418f3bd0, 32'h42094637, 32'h42856f87};
test_input[8696:8703] = '{32'hc2977f17, 32'h42a45fc5, 32'hc2a9bd04, 32'hc2a1012d, 32'h4272a671, 32'h41a9ab7e, 32'hc19a720e, 32'h42a81c60};
test_output[8696:8703] = '{32'h0, 32'h42a45fc5, 32'h0, 32'h0, 32'h4272a671, 32'h41a9ab7e, 32'h0, 32'h42a81c60};
test_input[8704:8711] = '{32'hc2b34930, 32'hc204c585, 32'h4124a051, 32'hc203f6f1, 32'h4293ca8d, 32'hc19849d0, 32'h42c7f699, 32'h40bacc3a};
test_output[8704:8711] = '{32'h0, 32'h0, 32'h4124a051, 32'h0, 32'h4293ca8d, 32'h0, 32'h42c7f699, 32'h40bacc3a};
test_input[8712:8719] = '{32'hc2b73780, 32'hc272f494, 32'hc17cd27c, 32'h4217c430, 32'hc1c5c8d6, 32'hc2b0e601, 32'hc2bd3b0b, 32'hc2b909df};
test_output[8712:8719] = '{32'h0, 32'h0, 32'h0, 32'h4217c430, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8720:8727] = '{32'h41c8997c, 32'hc2729091, 32'hc1a39821, 32'hc01ca926, 32'hc28c5f37, 32'h42175f55, 32'h428829d4, 32'hc171122a};
test_output[8720:8727] = '{32'h41c8997c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42175f55, 32'h428829d4, 32'h0};
test_input[8728:8735] = '{32'h421bce69, 32'hc1a90f52, 32'h4262c4da, 32'hc206ec86, 32'h4254447a, 32'hc2bbc700, 32'hc25f36dc, 32'h424306ea};
test_output[8728:8735] = '{32'h421bce69, 32'h0, 32'h4262c4da, 32'h0, 32'h4254447a, 32'h0, 32'h0, 32'h424306ea};
test_input[8736:8743] = '{32'hc2c31871, 32'hc1a4cdbf, 32'h411002cc, 32'h42158730, 32'h422f769f, 32'h42566d3e, 32'hc1dc5d7c, 32'hc18356b5};
test_output[8736:8743] = '{32'h0, 32'h0, 32'h411002cc, 32'h42158730, 32'h422f769f, 32'h42566d3e, 32'h0, 32'h0};
test_input[8744:8751] = '{32'h4265deca, 32'h420fc794, 32'h41603bde, 32'hc2840e66, 32'h42a17e6d, 32'hc0e9cc39, 32'hc21c6459, 32'h41c4eabe};
test_output[8744:8751] = '{32'h4265deca, 32'h420fc794, 32'h41603bde, 32'h0, 32'h42a17e6d, 32'h0, 32'h0, 32'h41c4eabe};
test_input[8752:8759] = '{32'h42496b5c, 32'h42920387, 32'h429c573e, 32'h429bb35e, 32'hc281a9ec, 32'hc1b92a61, 32'h41fd2a3e, 32'h3f8299de};
test_output[8752:8759] = '{32'h42496b5c, 32'h42920387, 32'h429c573e, 32'h429bb35e, 32'h0, 32'h0, 32'h41fd2a3e, 32'h3f8299de};
test_input[8760:8767] = '{32'hc2332461, 32'hc1843c63, 32'h41f1cd7c, 32'h40c60bbe, 32'h40fefa00, 32'h4282b83b, 32'h41e9a87e, 32'h41a9dad4};
test_output[8760:8767] = '{32'h0, 32'h0, 32'h41f1cd7c, 32'h40c60bbe, 32'h40fefa00, 32'h4282b83b, 32'h41e9a87e, 32'h41a9dad4};
test_input[8768:8775] = '{32'h42c27771, 32'h4247956b, 32'h4157c27b, 32'hc292e1ae, 32'h42739961, 32'h41b8b0c1, 32'hc2aaac87, 32'hc28a661c};
test_output[8768:8775] = '{32'h42c27771, 32'h4247956b, 32'h4157c27b, 32'h0, 32'h42739961, 32'h41b8b0c1, 32'h0, 32'h0};
test_input[8776:8783] = '{32'h420e3b38, 32'hc0ce6fa9, 32'hc28bb3cb, 32'h429e2e9a, 32'hc286e28d, 32'hc2b24741, 32'h42be758c, 32'hc27f6642};
test_output[8776:8783] = '{32'h420e3b38, 32'h0, 32'h0, 32'h429e2e9a, 32'h0, 32'h0, 32'h42be758c, 32'h0};
test_input[8784:8791] = '{32'hc1550834, 32'h41410820, 32'h4234c410, 32'hc0e8b72f, 32'hc2134b37, 32'h426c4cac, 32'h41682f89, 32'hc2a77027};
test_output[8784:8791] = '{32'h0, 32'h41410820, 32'h4234c410, 32'h0, 32'h0, 32'h426c4cac, 32'h41682f89, 32'h0};
test_input[8792:8799] = '{32'hc206e98e, 32'h42be60c1, 32'hc0fab58c, 32'h4298b023, 32'hc214a6f6, 32'hc1fd78fd, 32'hc0b7af01, 32'h4293e0f2};
test_output[8792:8799] = '{32'h0, 32'h42be60c1, 32'h0, 32'h4298b023, 32'h0, 32'h0, 32'h0, 32'h4293e0f2};
test_input[8800:8807] = '{32'hc2a61474, 32'hc2be6a4a, 32'hc2c4bfc1, 32'h426f6091, 32'hc29e10ef, 32'h4268ed15, 32'h428caf3a, 32'hc1f4b53b};
test_output[8800:8807] = '{32'h0, 32'h0, 32'h0, 32'h426f6091, 32'h0, 32'h4268ed15, 32'h428caf3a, 32'h0};
test_input[8808:8815] = '{32'h41ebcd19, 32'h429107c9, 32'hc23a1ad0, 32'h42930a5a, 32'hc1c6140d, 32'hc0975350, 32'h42363de3, 32'hc13fd106};
test_output[8808:8815] = '{32'h41ebcd19, 32'h429107c9, 32'h0, 32'h42930a5a, 32'h0, 32'h0, 32'h42363de3, 32'h0};
test_input[8816:8823] = '{32'hc202e81a, 32'hc29a7447, 32'hc2340454, 32'hc2716973, 32'hc289cfc3, 32'hc2b58740, 32'hc1c6fb5c, 32'hc266d658};
test_output[8816:8823] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8824:8831] = '{32'h428a9e44, 32'hc1926b05, 32'h426b6f93, 32'h41a3ba1c, 32'hc1abf090, 32'h42694d64, 32'h42c444f7, 32'hc2c22b88};
test_output[8824:8831] = '{32'h428a9e44, 32'h0, 32'h426b6f93, 32'h41a3ba1c, 32'h0, 32'h42694d64, 32'h42c444f7, 32'h0};
test_input[8832:8839] = '{32'h428eaf13, 32'h42b34929, 32'hc2934bd6, 32'h425bbae8, 32'hc28778ca, 32'hc2a981fd, 32'hc2944816, 32'h41e6db31};
test_output[8832:8839] = '{32'h428eaf13, 32'h42b34929, 32'h0, 32'h425bbae8, 32'h0, 32'h0, 32'h0, 32'h41e6db31};
test_input[8840:8847] = '{32'hc26fecfb, 32'h427c11f4, 32'h4299d72f, 32'hc1d36eff, 32'hc2b81a9f, 32'hc1ff97dc, 32'hc2095755, 32'h41d0f958};
test_output[8840:8847] = '{32'h0, 32'h427c11f4, 32'h4299d72f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41d0f958};
test_input[8848:8855] = '{32'hc223dc34, 32'hc1db446a, 32'hc2694102, 32'hc2016bc1, 32'hc257beda, 32'h42b071b5, 32'h4192b023, 32'hc299fa62};
test_output[8848:8855] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b071b5, 32'h4192b023, 32'h0};
test_input[8856:8863] = '{32'h42b6862b, 32'hc19ddbf6, 32'hc21cdd9f, 32'hc17432c5, 32'h42802b9b, 32'hc1304089, 32'hc1462d2d, 32'h4187ebd6};
test_output[8856:8863] = '{32'h42b6862b, 32'h0, 32'h0, 32'h0, 32'h42802b9b, 32'h0, 32'h0, 32'h4187ebd6};
test_input[8864:8871] = '{32'hc1cbad33, 32'h42398679, 32'h40d0b76f, 32'h42b9b489, 32'hc2ab8e45, 32'hc28a7c59, 32'hc06ca58b, 32'h42163eeb};
test_output[8864:8871] = '{32'h0, 32'h42398679, 32'h40d0b76f, 32'h42b9b489, 32'h0, 32'h0, 32'h0, 32'h42163eeb};
test_input[8872:8879] = '{32'hc19ef499, 32'hc084789e, 32'hc1a57a63, 32'h41f44b98, 32'h403eb89e, 32'h429a69b1, 32'h4286cbc4, 32'hc2b0b1a9};
test_output[8872:8879] = '{32'h0, 32'h0, 32'h0, 32'h41f44b98, 32'h403eb89e, 32'h429a69b1, 32'h4286cbc4, 32'h0};
test_input[8880:8887] = '{32'h41bf2953, 32'h424db20a, 32'h42bafa36, 32'h42c5f2cc, 32'h4278a126, 32'hc2977ab4, 32'h42910971, 32'h42442341};
test_output[8880:8887] = '{32'h41bf2953, 32'h424db20a, 32'h42bafa36, 32'h42c5f2cc, 32'h4278a126, 32'h0, 32'h42910971, 32'h42442341};
test_input[8888:8895] = '{32'hc2b17a1c, 32'h42593fc3, 32'h3f1bb46c, 32'hc2b0ae5d, 32'h41f11440, 32'hc2c18307, 32'hc17987d2, 32'h403e661a};
test_output[8888:8895] = '{32'h0, 32'h42593fc3, 32'h3f1bb46c, 32'h0, 32'h41f11440, 32'h0, 32'h0, 32'h403e661a};
test_input[8896:8903] = '{32'h426f3a18, 32'h41da61ea, 32'hc1f32094, 32'h42898b4f, 32'h424e5756, 32'hc2313a20, 32'h426856d5, 32'hc29d88e2};
test_output[8896:8903] = '{32'h426f3a18, 32'h41da61ea, 32'h0, 32'h42898b4f, 32'h424e5756, 32'h0, 32'h426856d5, 32'h0};
test_input[8904:8911] = '{32'hc1adfc2e, 32'hc1dcac56, 32'hc23cb0a3, 32'h413cde41, 32'hc20bd056, 32'h40bd47e6, 32'hc2c524d2, 32'hc288aed5};
test_output[8904:8911] = '{32'h0, 32'h0, 32'h0, 32'h413cde41, 32'h0, 32'h40bd47e6, 32'h0, 32'h0};
test_input[8912:8919] = '{32'h420f9b90, 32'hc1a16943, 32'h3f988fbc, 32'hc245a09e, 32'h4291ad33, 32'hc22f63fb, 32'hc2b34cc9, 32'hc21e5939};
test_output[8912:8919] = '{32'h420f9b90, 32'h0, 32'h3f988fbc, 32'h0, 32'h4291ad33, 32'h0, 32'h0, 32'h0};
test_input[8920:8927] = '{32'hc29bb383, 32'hc2a681c1, 32'h4236c9eb, 32'h427506f3, 32'hc28100df, 32'h422814ef, 32'hc2aec249, 32'hc040849d};
test_output[8920:8927] = '{32'h0, 32'h0, 32'h4236c9eb, 32'h427506f3, 32'h0, 32'h422814ef, 32'h0, 32'h0};
test_input[8928:8935] = '{32'h42304d1b, 32'h42a61e00, 32'h42ae8c11, 32'h42580518, 32'h429cba8a, 32'hc2554f8f, 32'h41421612, 32'hc28bc2a4};
test_output[8928:8935] = '{32'h42304d1b, 32'h42a61e00, 32'h42ae8c11, 32'h42580518, 32'h429cba8a, 32'h0, 32'h41421612, 32'h0};
test_input[8936:8943] = '{32'h428eade5, 32'h4190849d, 32'h42c4ebbc, 32'h428c1e7a, 32'hc2860bad, 32'hbf3e0101, 32'h41b49670, 32'hc2bb09b6};
test_output[8936:8943] = '{32'h428eade5, 32'h4190849d, 32'h42c4ebbc, 32'h428c1e7a, 32'h0, 32'h0, 32'h41b49670, 32'h0};
test_input[8944:8951] = '{32'hc2b68687, 32'hc0efefd0, 32'hc2084bee, 32'h42aae63c, 32'hc2b85a53, 32'h3f9b8064, 32'hc15c326d, 32'h411ff66b};
test_output[8944:8951] = '{32'h0, 32'h0, 32'h0, 32'h42aae63c, 32'h0, 32'h3f9b8064, 32'h0, 32'h411ff66b};
test_input[8952:8959] = '{32'h41f71891, 32'h42bc8d3d, 32'hc23918f4, 32'hc02fa461, 32'hc2bdb397, 32'hc1a41996, 32'hc2aa1b0f, 32'h42628d34};
test_output[8952:8959] = '{32'h41f71891, 32'h42bc8d3d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42628d34};
test_input[8960:8967] = '{32'hc25bd469, 32'h40ce2a33, 32'hc223e1c3, 32'h424e4825, 32'h420530cb, 32'h427b19eb, 32'hc1c62b21, 32'hc2715fa6};
test_output[8960:8967] = '{32'h0, 32'h40ce2a33, 32'h0, 32'h424e4825, 32'h420530cb, 32'h427b19eb, 32'h0, 32'h0};
test_input[8968:8975] = '{32'hc289d497, 32'h42b6c731, 32'h42071015, 32'hc18a39d1, 32'hc22fee19, 32'h42c62605, 32'h415ac4c5, 32'hbfeddd13};
test_output[8968:8975] = '{32'h0, 32'h42b6c731, 32'h42071015, 32'h0, 32'h0, 32'h42c62605, 32'h415ac4c5, 32'h0};
test_input[8976:8983] = '{32'h40bcafa0, 32'h42c1e41c, 32'h41f8b690, 32'hc22ea24c, 32'hc27abcd5, 32'h406f2a22, 32'hc2b09ab6, 32'h41c6e660};
test_output[8976:8983] = '{32'h40bcafa0, 32'h42c1e41c, 32'h41f8b690, 32'h0, 32'h0, 32'h406f2a22, 32'h0, 32'h41c6e660};
test_input[8984:8991] = '{32'hc2a8dddf, 32'hc295d589, 32'hc0e24c7e, 32'h41694a6d, 32'hc29bbdc9, 32'hc2409da0, 32'hc261a592, 32'h4279d740};
test_output[8984:8991] = '{32'h0, 32'h0, 32'h0, 32'h41694a6d, 32'h0, 32'h0, 32'h0, 32'h4279d740};
test_input[8992:8999] = '{32'hc222af3d, 32'hc2059965, 32'hc292ca04, 32'hc287f3ee, 32'h4281c07b, 32'hc26347d5, 32'hc2652d8f, 32'hc26ede6e};
test_output[8992:8999] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4281c07b, 32'h0, 32'h0, 32'h0};
test_input[9000:9007] = '{32'hbf1d9e2a, 32'h41fde55d, 32'h4034f64a, 32'hc1dbce34, 32'hc297c611, 32'hc1e97fd7, 32'hc21d4add, 32'hc10a24d6};
test_output[9000:9007] = '{32'h0, 32'h41fde55d, 32'h4034f64a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9008:9015] = '{32'hc19353ad, 32'hc292899a, 32'hc271049a, 32'h42149d4b, 32'h41b1f162, 32'hc24045fa, 32'hc2b10a32, 32'h4240d5b9};
test_output[9008:9015] = '{32'h0, 32'h0, 32'h0, 32'h42149d4b, 32'h41b1f162, 32'h0, 32'h0, 32'h4240d5b9};
test_input[9016:9023] = '{32'h41d77f19, 32'h41459715, 32'hc246eaf0, 32'h42689d9c, 32'hc0ce94e5, 32'hc1d11a29, 32'hc21476b6, 32'hc299d236};
test_output[9016:9023] = '{32'h41d77f19, 32'h41459715, 32'h0, 32'h42689d9c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9024:9031] = '{32'hc03a79ea, 32'h42903090, 32'hc28b15ac, 32'hc2b2bd88, 32'hc22c0849, 32'hc17bb008, 32'hc2a03d5f, 32'hc2a268c5};
test_output[9024:9031] = '{32'h0, 32'h42903090, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9032:9039] = '{32'hc28000c7, 32'h42b719d6, 32'hc22a7c9d, 32'hc0dc65f1, 32'hc21862b6, 32'h42498649, 32'hc20259ea, 32'hc22e7e44};
test_output[9032:9039] = '{32'h0, 32'h42b719d6, 32'h0, 32'h0, 32'h0, 32'h42498649, 32'h0, 32'h0};
test_input[9040:9047] = '{32'h41cb58e5, 32'h42c08516, 32'hc29ccce6, 32'hc222211d, 32'h421eafa4, 32'hc1a803a8, 32'h41edc0f7, 32'hc2950ccf};
test_output[9040:9047] = '{32'h41cb58e5, 32'h42c08516, 32'h0, 32'h0, 32'h421eafa4, 32'h0, 32'h41edc0f7, 32'h0};
test_input[9048:9055] = '{32'h41ecf996, 32'hc2bd9414, 32'h419d37f0, 32'hc19b0b80, 32'hc1d0ecd7, 32'h42883de6, 32'hc283ef41, 32'h422fa5fc};
test_output[9048:9055] = '{32'h41ecf996, 32'h0, 32'h419d37f0, 32'h0, 32'h0, 32'h42883de6, 32'h0, 32'h422fa5fc};
test_input[9056:9063] = '{32'h420b85d9, 32'h42bf239e, 32'hc1e48295, 32'hbf947acd, 32'hc2c10256, 32'hc2be3ef0, 32'hc28f5976, 32'h42065326};
test_output[9056:9063] = '{32'h420b85d9, 32'h42bf239e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42065326};
test_input[9064:9071] = '{32'h41e3f3fd, 32'hc1e54079, 32'h40d75ec5, 32'hc2c4aa63, 32'h42819f8c, 32'h423eb941, 32'h41b6f27c, 32'hc20a4655};
test_output[9064:9071] = '{32'h41e3f3fd, 32'h0, 32'h40d75ec5, 32'h0, 32'h42819f8c, 32'h423eb941, 32'h41b6f27c, 32'h0};
test_input[9072:9079] = '{32'hc28f4ec8, 32'hc1b1cb91, 32'h41a4ca58, 32'h41e40ad5, 32'h42c4b662, 32'hc208f90a, 32'hc1d9fed8, 32'hc23a0bf6};
test_output[9072:9079] = '{32'h0, 32'h0, 32'h41a4ca58, 32'h41e40ad5, 32'h42c4b662, 32'h0, 32'h0, 32'h0};
test_input[9080:9087] = '{32'hc2638d5e, 32'h42800443, 32'h42013a06, 32'h42b945c5, 32'hc2a0c563, 32'h4174356d, 32'h422ee4c3, 32'hc18013d8};
test_output[9080:9087] = '{32'h0, 32'h42800443, 32'h42013a06, 32'h42b945c5, 32'h0, 32'h4174356d, 32'h422ee4c3, 32'h0};
test_input[9088:9095] = '{32'hc20f450b, 32'h3e9718f1, 32'hc264707e, 32'hc2a9f7aa, 32'hc2917bd4, 32'hc2a41a8e, 32'h423ab9f7, 32'h42a8a82b};
test_output[9088:9095] = '{32'h0, 32'h3e9718f1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423ab9f7, 32'h42a8a82b};
test_input[9096:9103] = '{32'hc09a8b6a, 32'h42c1f57c, 32'h42928403, 32'hc29555dc, 32'hc277050a, 32'h424136de, 32'h424e6d83, 32'hc2b0bab7};
test_output[9096:9103] = '{32'h0, 32'h42c1f57c, 32'h42928403, 32'h0, 32'h0, 32'h424136de, 32'h424e6d83, 32'h0};
test_input[9104:9111] = '{32'h424d1731, 32'h4204a445, 32'hc20de55b, 32'h413ae86e, 32'h417254c7, 32'h429eb34b, 32'h424fb1c9, 32'hc213f8b3};
test_output[9104:9111] = '{32'h424d1731, 32'h4204a445, 32'h0, 32'h413ae86e, 32'h417254c7, 32'h429eb34b, 32'h424fb1c9, 32'h0};
test_input[9112:9119] = '{32'hc2725656, 32'h4263a8aa, 32'h425fb612, 32'hc285d619, 32'h427c9dff, 32'hc28ffad1, 32'h422ff261, 32'hc2a98471};
test_output[9112:9119] = '{32'h0, 32'h4263a8aa, 32'h425fb612, 32'h0, 32'h427c9dff, 32'h0, 32'h422ff261, 32'h0};
test_input[9120:9127] = '{32'hc1be23f3, 32'h402d35ea, 32'hc0586cdc, 32'h41c9fc16, 32'hc2bb2e44, 32'hc2a4df37, 32'h42517b28, 32'h427826ae};
test_output[9120:9127] = '{32'h0, 32'h402d35ea, 32'h0, 32'h41c9fc16, 32'h0, 32'h0, 32'h42517b28, 32'h427826ae};
test_input[9128:9135] = '{32'hc277c746, 32'hc0ff8aae, 32'h426b8cd7, 32'h42a75574, 32'hc2b1b2fc, 32'h412b323c, 32'h4299d041, 32'hc2963f75};
test_output[9128:9135] = '{32'h0, 32'h0, 32'h426b8cd7, 32'h42a75574, 32'h0, 32'h412b323c, 32'h4299d041, 32'h0};
test_input[9136:9143] = '{32'hc1ac331f, 32'hc1c6b03d, 32'hc1ebfb21, 32'hc1d843d0, 32'hc21cc254, 32'h42bf027d, 32'h424eb1bf, 32'hc20067e9};
test_output[9136:9143] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bf027d, 32'h424eb1bf, 32'h0};
test_input[9144:9151] = '{32'hc2081557, 32'hc2b02dcd, 32'h409e50c4, 32'hc1ffd243, 32'h41d3509f, 32'h42a06154, 32'hc2ae2cc8, 32'hc280c044};
test_output[9144:9151] = '{32'h0, 32'h0, 32'h409e50c4, 32'h0, 32'h41d3509f, 32'h42a06154, 32'h0, 32'h0};
test_input[9152:9159] = '{32'hc23d2600, 32'hc243fe29, 32'hc2a29b24, 32'h41172600, 32'hc2622b65, 32'h42c17a7d, 32'h41dce7ea, 32'h42938ad5};
test_output[9152:9159] = '{32'h0, 32'h0, 32'h0, 32'h41172600, 32'h0, 32'h42c17a7d, 32'h41dce7ea, 32'h42938ad5};
test_input[9160:9167] = '{32'h42a59076, 32'h42a1d90a, 32'hc218727b, 32'hc2224b14, 32'h42139805, 32'h41cd5cb9, 32'hc21aa05e, 32'h42c15f75};
test_output[9160:9167] = '{32'h42a59076, 32'h42a1d90a, 32'h0, 32'h0, 32'h42139805, 32'h41cd5cb9, 32'h0, 32'h42c15f75};
test_input[9168:9175] = '{32'h4257114c, 32'hc25bbd65, 32'h422c5311, 32'h41bb0b9b, 32'h42c61174, 32'hc269d211, 32'hc2341dba, 32'h423081df};
test_output[9168:9175] = '{32'h4257114c, 32'h0, 32'h422c5311, 32'h41bb0b9b, 32'h42c61174, 32'h0, 32'h0, 32'h423081df};
test_input[9176:9183] = '{32'hc16db8c2, 32'h4299911e, 32'hc254cb57, 32'hc2bf3cbd, 32'hc1fb4e06, 32'h412f4f43, 32'h42a99257, 32'h424472f3};
test_output[9176:9183] = '{32'h0, 32'h4299911e, 32'h0, 32'h0, 32'h0, 32'h412f4f43, 32'h42a99257, 32'h424472f3};
test_input[9184:9191] = '{32'hc1b8b1f9, 32'hc2c069f7, 32'h411087d9, 32'h41970f8d, 32'h4298d6f8, 32'hc26383fb, 32'h4227a645, 32'h42ac2183};
test_output[9184:9191] = '{32'h0, 32'h0, 32'h411087d9, 32'h41970f8d, 32'h4298d6f8, 32'h0, 32'h4227a645, 32'h42ac2183};
test_input[9192:9199] = '{32'hc26b2120, 32'hbf31d8fe, 32'hc235aae5, 32'hc26a3b42, 32'h427ed208, 32'hc189b349, 32'h40c7d251, 32'h4297ae74};
test_output[9192:9199] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h427ed208, 32'h0, 32'h40c7d251, 32'h4297ae74};
test_input[9200:9207] = '{32'h423ca640, 32'hc2595c9c, 32'hc21d737f, 32'hc20864f9, 32'hc2929fb2, 32'h42444338, 32'hc1854972, 32'h42a5ce1c};
test_output[9200:9207] = '{32'h423ca640, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42444338, 32'h0, 32'h42a5ce1c};
test_input[9208:9215] = '{32'hc20b443b, 32'hc247c308, 32'hc28ce6de, 32'hc2bd6d17, 32'h429219b7, 32'h4281b40e, 32'hc2bd6961, 32'hc2b53413};
test_output[9208:9215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429219b7, 32'h4281b40e, 32'h0, 32'h0};
test_input[9216:9223] = '{32'hc1ebf9c0, 32'h42b9c284, 32'h41ea1322, 32'hc06b8d2d, 32'hc29f718e, 32'h428232f7, 32'hc1fd20b6, 32'hc2bc953f};
test_output[9216:9223] = '{32'h0, 32'h42b9c284, 32'h41ea1322, 32'h0, 32'h0, 32'h428232f7, 32'h0, 32'h0};
test_input[9224:9231] = '{32'h40dbf11e, 32'hc235aece, 32'hc2c36844, 32'h412fe504, 32'hc2a61f8c, 32'h41970276, 32'hc2231dab, 32'h42ad1378};
test_output[9224:9231] = '{32'h40dbf11e, 32'h0, 32'h0, 32'h412fe504, 32'h0, 32'h41970276, 32'h0, 32'h42ad1378};
test_input[9232:9239] = '{32'h425518d4, 32'hc13b8db4, 32'h429ea455, 32'h42c0cde7, 32'hc2b3cb07, 32'hc1b70194, 32'hbfd1f6b2, 32'hc25d274f};
test_output[9232:9239] = '{32'h425518d4, 32'h0, 32'h429ea455, 32'h42c0cde7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9240:9247] = '{32'hc2591dfd, 32'hc141e46b, 32'hc215aeed, 32'hc2c1d6e2, 32'h424d0fb0, 32'hc2bb6cf2, 32'hc26298fe, 32'hbfc45a0f};
test_output[9240:9247] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h424d0fb0, 32'h0, 32'h0, 32'h0};
test_input[9248:9255] = '{32'h40c6c4e1, 32'h429293cd, 32'h4251e60c, 32'h41511a20, 32'h4284c908, 32'h42302b7a, 32'h427a687b, 32'h42828a8e};
test_output[9248:9255] = '{32'h40c6c4e1, 32'h429293cd, 32'h4251e60c, 32'h41511a20, 32'h4284c908, 32'h42302b7a, 32'h427a687b, 32'h42828a8e};
test_input[9256:9263] = '{32'h40a9ab5c, 32'h417c7f31, 32'h42c0cc5b, 32'hc2bc690f, 32'h421ccfe9, 32'hc1ddd974, 32'h42611178, 32'h42be9d8b};
test_output[9256:9263] = '{32'h40a9ab5c, 32'h417c7f31, 32'h42c0cc5b, 32'h0, 32'h421ccfe9, 32'h0, 32'h42611178, 32'h42be9d8b};
test_input[9264:9271] = '{32'hc281a068, 32'h40f99d21, 32'hc131d200, 32'h42b3e7f0, 32'hc231defa, 32'hc1498482, 32'hc1579604, 32'hc21497a4};
test_output[9264:9271] = '{32'h0, 32'h40f99d21, 32'h0, 32'h42b3e7f0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9272:9279] = '{32'hc20dac40, 32'h41898c75, 32'h42174ef0, 32'hc25790ae, 32'hc2045c60, 32'h4207821d, 32'h4226f053, 32'h41b026b4};
test_output[9272:9279] = '{32'h0, 32'h41898c75, 32'h42174ef0, 32'h0, 32'h0, 32'h4207821d, 32'h4226f053, 32'h41b026b4};
test_input[9280:9287] = '{32'h42b54835, 32'hc18d12c9, 32'h41e5444a, 32'h426f538f, 32'hc2bee4f0, 32'h416e3f75, 32'h425a0f1e, 32'hc27fd261};
test_output[9280:9287] = '{32'h42b54835, 32'h0, 32'h41e5444a, 32'h426f538f, 32'h0, 32'h416e3f75, 32'h425a0f1e, 32'h0};
test_input[9288:9295] = '{32'h40ea48ed, 32'h4103a8c7, 32'h42a92ff4, 32'h408e38d1, 32'h427a67af, 32'h429fcf20, 32'hc1592d2e, 32'hc2353773};
test_output[9288:9295] = '{32'h40ea48ed, 32'h4103a8c7, 32'h42a92ff4, 32'h408e38d1, 32'h427a67af, 32'h429fcf20, 32'h0, 32'h0};
test_input[9296:9303] = '{32'h4292ab69, 32'h4285b676, 32'h42aaf226, 32'h41c4b4ef, 32'hc2bf1b30, 32'h41649691, 32'h42bc4107, 32'hc2c03938};
test_output[9296:9303] = '{32'h4292ab69, 32'h4285b676, 32'h42aaf226, 32'h41c4b4ef, 32'h0, 32'h41649691, 32'h42bc4107, 32'h0};
test_input[9304:9311] = '{32'hc285c2a7, 32'h424aac08, 32'hc2595efc, 32'hc2542182, 32'h40f4fd17, 32'h4292c15f, 32'hc1b86ba7, 32'h42ba5f92};
test_output[9304:9311] = '{32'h0, 32'h424aac08, 32'h0, 32'h0, 32'h40f4fd17, 32'h4292c15f, 32'h0, 32'h42ba5f92};
test_input[9312:9319] = '{32'hc1a45204, 32'hc152e148, 32'h42497eb2, 32'hc25b6f24, 32'h42b9d604, 32'h41bae862, 32'h4209e5f9, 32'h42964183};
test_output[9312:9319] = '{32'h0, 32'h0, 32'h42497eb2, 32'h0, 32'h42b9d604, 32'h41bae862, 32'h4209e5f9, 32'h42964183};
test_input[9320:9327] = '{32'hc25562a2, 32'hc2c514a0, 32'h414d164a, 32'h42a46448, 32'hc2437c23, 32'h4107d745, 32'h42a01162, 32'hc2894048};
test_output[9320:9327] = '{32'h0, 32'h0, 32'h414d164a, 32'h42a46448, 32'h0, 32'h4107d745, 32'h42a01162, 32'h0};
test_input[9328:9335] = '{32'hc2b3b9f3, 32'hc291817b, 32'hc2c1c462, 32'h427f209a, 32'h413ec0c1, 32'h4292ca7f, 32'hc2c4d692, 32'h42ba5e8d};
test_output[9328:9335] = '{32'h0, 32'h0, 32'h0, 32'h427f209a, 32'h413ec0c1, 32'h4292ca7f, 32'h0, 32'h42ba5e8d};
test_input[9336:9343] = '{32'hc2a40762, 32'h42840ea9, 32'hc2178c98, 32'h42c0e71b, 32'h417261db, 32'h42bb829b, 32'hc0674b70, 32'hc2c374e8};
test_output[9336:9343] = '{32'h0, 32'h42840ea9, 32'h0, 32'h42c0e71b, 32'h417261db, 32'h42bb829b, 32'h0, 32'h0};
test_input[9344:9351] = '{32'h41a3416a, 32'h421d7bf7, 32'hc2855c58, 32'h415b23b4, 32'hc102b3a7, 32'h41cc892a, 32'h427d489e, 32'hc1f2254e};
test_output[9344:9351] = '{32'h41a3416a, 32'h421d7bf7, 32'h0, 32'h415b23b4, 32'h0, 32'h41cc892a, 32'h427d489e, 32'h0};
test_input[9352:9359] = '{32'h410a8b21, 32'hc2a721b2, 32'hc2af2215, 32'hc290970a, 32'hc2811fe5, 32'hc251148c, 32'hc21e84c4, 32'hc1a91365};
test_output[9352:9359] = '{32'h410a8b21, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9360:9367] = '{32'hc0c6c5b9, 32'h428a2a7c, 32'h41f3b0a4, 32'h42511a3d, 32'hc29fee11, 32'hc09a18ce, 32'hc26280ff, 32'h42882424};
test_output[9360:9367] = '{32'h0, 32'h428a2a7c, 32'h41f3b0a4, 32'h42511a3d, 32'h0, 32'h0, 32'h0, 32'h42882424};
test_input[9368:9375] = '{32'h41c542f2, 32'h42714efd, 32'hc194f286, 32'hc116ce1a, 32'h42483ed3, 32'h42591527, 32'hc20b7ce7, 32'h428d5db9};
test_output[9368:9375] = '{32'h41c542f2, 32'h42714efd, 32'h0, 32'h0, 32'h42483ed3, 32'h42591527, 32'h0, 32'h428d5db9};
test_input[9376:9383] = '{32'hc1e051ac, 32'h428810a9, 32'h4275d6e4, 32'h42626ef4, 32'hc2a025aa, 32'hbf2cfb61, 32'h42b8cde1, 32'hc00a2e52};
test_output[9376:9383] = '{32'h0, 32'h428810a9, 32'h4275d6e4, 32'h42626ef4, 32'h0, 32'h0, 32'h42b8cde1, 32'h0};
test_input[9384:9391] = '{32'h42bbf777, 32'hc2815575, 32'hc255ea76, 32'hc11dafed, 32'hc2c739f2, 32'h42803c4a, 32'h4132075e, 32'h424c9fff};
test_output[9384:9391] = '{32'h42bbf777, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42803c4a, 32'h4132075e, 32'h424c9fff};
test_input[9392:9399] = '{32'hc224e614, 32'h419415e1, 32'hc2b76c45, 32'hc26fd87b, 32'h421e0f3b, 32'h428184dc, 32'h429a92e6, 32'h420bc617};
test_output[9392:9399] = '{32'h0, 32'h419415e1, 32'h0, 32'h0, 32'h421e0f3b, 32'h428184dc, 32'h429a92e6, 32'h420bc617};
test_input[9400:9407] = '{32'hc1ec8cc4, 32'h41cc20ae, 32'h421f5f82, 32'hc1bd1d19, 32'h42b1093f, 32'h40e68eef, 32'hc20ecbfc, 32'h41986bc5};
test_output[9400:9407] = '{32'h0, 32'h41cc20ae, 32'h421f5f82, 32'h0, 32'h42b1093f, 32'h40e68eef, 32'h0, 32'h41986bc5};
test_input[9408:9415] = '{32'h41d0392b, 32'h4180fd0e, 32'h425e9f3a, 32'h42a89b46, 32'h41a466f3, 32'hc20ac108, 32'h4280aadc, 32'hc12af121};
test_output[9408:9415] = '{32'h41d0392b, 32'h4180fd0e, 32'h425e9f3a, 32'h42a89b46, 32'h41a466f3, 32'h0, 32'h4280aadc, 32'h0};
test_input[9416:9423] = '{32'hc298a096, 32'hc1ae98ad, 32'h418db730, 32'h428380f9, 32'h429d47c5, 32'h413b4c7b, 32'hc0d33e99, 32'h42593941};
test_output[9416:9423] = '{32'h0, 32'h0, 32'h418db730, 32'h428380f9, 32'h429d47c5, 32'h413b4c7b, 32'h0, 32'h42593941};
test_input[9424:9431] = '{32'h41610893, 32'h42887eff, 32'hc2bedeb1, 32'hc1b9ac3a, 32'h40c2c0dd, 32'h41843aa0, 32'hc09ab825, 32'h42896e9d};
test_output[9424:9431] = '{32'h41610893, 32'h42887eff, 32'h0, 32'h0, 32'h40c2c0dd, 32'h41843aa0, 32'h0, 32'h42896e9d};
test_input[9432:9439] = '{32'h42c684ec, 32'h422aeaab, 32'hc219a20d, 32'hc176c86b, 32'h417d34e0, 32'hc2a3dc7a, 32'hc2b14bc0, 32'h4235c9ab};
test_output[9432:9439] = '{32'h42c684ec, 32'h422aeaab, 32'h0, 32'h0, 32'h417d34e0, 32'h0, 32'h0, 32'h4235c9ab};
test_input[9440:9447] = '{32'h4275b282, 32'h41d278f7, 32'hbeaaa7b7, 32'h41d3b115, 32'h425d357f, 32'hc2b0f490, 32'hc1487f6d, 32'hc1eb5852};
test_output[9440:9447] = '{32'h4275b282, 32'h41d278f7, 32'h0, 32'h41d3b115, 32'h425d357f, 32'h0, 32'h0, 32'h0};
test_input[9448:9455] = '{32'h428e9115, 32'h42bc258c, 32'hc20e6fad, 32'hc2babd5a, 32'h42a8c5d8, 32'h42900d94, 32'h4130459f, 32'hc240ca53};
test_output[9448:9455] = '{32'h428e9115, 32'h42bc258c, 32'h0, 32'h0, 32'h42a8c5d8, 32'h42900d94, 32'h4130459f, 32'h0};
test_input[9456:9463] = '{32'hc2aaa019, 32'hc1e47e59, 32'h42b2ae4c, 32'hc29340b8, 32'h426fa1cc, 32'hc155af3f, 32'hc25ad35f, 32'h42c5d943};
test_output[9456:9463] = '{32'h0, 32'h0, 32'h42b2ae4c, 32'h0, 32'h426fa1cc, 32'h0, 32'h0, 32'h42c5d943};
test_input[9464:9471] = '{32'hc224085e, 32'hc275f298, 32'hc2bc6427, 32'h42bddafd, 32'hc2bdb6dd, 32'hc08e82b6, 32'h42c2408d, 32'h422d5792};
test_output[9464:9471] = '{32'h0, 32'h0, 32'h0, 32'h42bddafd, 32'h0, 32'h0, 32'h42c2408d, 32'h422d5792};
test_input[9472:9479] = '{32'h42521cc8, 32'hc2c27ec2, 32'h429973bb, 32'hc21d338c, 32'h42c14636, 32'hc249bde0, 32'h4228f5d1, 32'h4290e856};
test_output[9472:9479] = '{32'h42521cc8, 32'h0, 32'h429973bb, 32'h0, 32'h42c14636, 32'h0, 32'h4228f5d1, 32'h4290e856};
test_input[9480:9487] = '{32'hc26d44fc, 32'hc0967ddf, 32'hc26e0c57, 32'h42b18a4a, 32'hc23ab099, 32'h41368cbb, 32'hc2b7a7d7, 32'hc2a10715};
test_output[9480:9487] = '{32'h0, 32'h0, 32'h0, 32'h42b18a4a, 32'h0, 32'h41368cbb, 32'h0, 32'h0};
test_input[9488:9495] = '{32'hc28cec7a, 32'h41f08607, 32'hc2aca816, 32'hc2a3861f, 32'hc213ab42, 32'h41dc3251, 32'h42514290, 32'h4255774d};
test_output[9488:9495] = '{32'h0, 32'h41f08607, 32'h0, 32'h0, 32'h0, 32'h41dc3251, 32'h42514290, 32'h4255774d};
test_input[9496:9503] = '{32'h42c3cd8d, 32'hc1e42580, 32'hc1c25bb8, 32'hc29893d0, 32'h414a85c1, 32'h41c0ab74, 32'h426ff228, 32'hc1a6cc26};
test_output[9496:9503] = '{32'h42c3cd8d, 32'h0, 32'h0, 32'h0, 32'h414a85c1, 32'h41c0ab74, 32'h426ff228, 32'h0};
test_input[9504:9511] = '{32'h4226200b, 32'h42a0e98b, 32'h4239e85d, 32'hc29dd422, 32'h42a96898, 32'hc2b039e7, 32'h426f9aba, 32'hc189323f};
test_output[9504:9511] = '{32'h4226200b, 32'h42a0e98b, 32'h4239e85d, 32'h0, 32'h42a96898, 32'h0, 32'h426f9aba, 32'h0};
test_input[9512:9519] = '{32'hc21d89b2, 32'hc20e6cca, 32'hc26f75ec, 32'hc1af4304, 32'hc2c13c9f, 32'h42333042, 32'hc25ea7c7, 32'h42bca3c6};
test_output[9512:9519] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42333042, 32'h0, 32'h42bca3c6};
test_input[9520:9527] = '{32'h4265bf89, 32'hc1292f38, 32'h41dcaad3, 32'h42c4d728, 32'hc111fcfd, 32'h41d694d1, 32'hc292cd79, 32'h42c344fe};
test_output[9520:9527] = '{32'h4265bf89, 32'h0, 32'h41dcaad3, 32'h42c4d728, 32'h0, 32'h41d694d1, 32'h0, 32'h42c344fe};
test_input[9528:9535] = '{32'h423b5e14, 32'h41af9d09, 32'h417651d8, 32'hc240bb3e, 32'h4283cc2f, 32'h41f7fab7, 32'h413c28ad, 32'h4231aff2};
test_output[9528:9535] = '{32'h423b5e14, 32'h41af9d09, 32'h417651d8, 32'h0, 32'h4283cc2f, 32'h41f7fab7, 32'h413c28ad, 32'h4231aff2};
test_input[9536:9543] = '{32'hc29b2be5, 32'h42b6f3e8, 32'hc21cab8a, 32'hc2a93184, 32'hc23e5880, 32'hc28f0ca2, 32'h41db8405, 32'hc1f96190};
test_output[9536:9543] = '{32'h0, 32'h42b6f3e8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41db8405, 32'h0};
test_input[9544:9551] = '{32'h42a14994, 32'h423511cf, 32'h413310fa, 32'hc29754ad, 32'h40936db0, 32'hc281546a, 32'h42283563, 32'h42822644};
test_output[9544:9551] = '{32'h42a14994, 32'h423511cf, 32'h413310fa, 32'h0, 32'h40936db0, 32'h0, 32'h42283563, 32'h42822644};
test_input[9552:9559] = '{32'h42381592, 32'h41e20fc8, 32'hc260e310, 32'h4252e099, 32'h41005b64, 32'h418932c7, 32'hc130d3dd, 32'hc2c45467};
test_output[9552:9559] = '{32'h42381592, 32'h41e20fc8, 32'h0, 32'h4252e099, 32'h41005b64, 32'h418932c7, 32'h0, 32'h0};
test_input[9560:9567] = '{32'hc20062f6, 32'hc1541d18, 32'h4252558a, 32'hc2c10363, 32'hc2934716, 32'h41dc21d6, 32'h41bce4c2, 32'h3d2d9395};
test_output[9560:9567] = '{32'h0, 32'h0, 32'h4252558a, 32'h0, 32'h0, 32'h41dc21d6, 32'h41bce4c2, 32'h3d2d9395};
test_input[9568:9575] = '{32'h421ab24e, 32'hc270e1d2, 32'h4259eecd, 32'hc02fee5a, 32'h42709180, 32'hc292a650, 32'hc2b51a1a, 32'h428d3f1d};
test_output[9568:9575] = '{32'h421ab24e, 32'h0, 32'h4259eecd, 32'h0, 32'h42709180, 32'h0, 32'h0, 32'h428d3f1d};
test_input[9576:9583] = '{32'h42654436, 32'h4208ff2d, 32'h421dd91c, 32'hc1304625, 32'h406b8e8e, 32'h42b01eec, 32'hc22c7745, 32'h42c28c41};
test_output[9576:9583] = '{32'h42654436, 32'h4208ff2d, 32'h421dd91c, 32'h0, 32'h406b8e8e, 32'h42b01eec, 32'h0, 32'h42c28c41};
test_input[9584:9591] = '{32'h41368ec3, 32'h42182eff, 32'hc2c3e842, 32'h4220a16c, 32'h42861903, 32'h41e2b166, 32'hc26ac9b1, 32'hc173fcd4};
test_output[9584:9591] = '{32'h41368ec3, 32'h42182eff, 32'h0, 32'h4220a16c, 32'h42861903, 32'h41e2b166, 32'h0, 32'h0};
test_input[9592:9599] = '{32'hc25bdf5c, 32'h41a45f85, 32'h42c300b6, 32'h424ca02b, 32'hc26a08d1, 32'hc239f307, 32'h421e6c11, 32'hc1b559a6};
test_output[9592:9599] = '{32'h0, 32'h41a45f85, 32'h42c300b6, 32'h424ca02b, 32'h0, 32'h0, 32'h421e6c11, 32'h0};
test_input[9600:9607] = '{32'h4212158f, 32'h4294ce53, 32'h41c25f7e, 32'h42a5aba8, 32'hc12c6abd, 32'hc1961574, 32'h42b2001d, 32'hc1e6775a};
test_output[9600:9607] = '{32'h4212158f, 32'h4294ce53, 32'h41c25f7e, 32'h42a5aba8, 32'h0, 32'h0, 32'h42b2001d, 32'h0};
test_input[9608:9615] = '{32'hc221605d, 32'hc26f77db, 32'hc2c6ed06, 32'h41166d5a, 32'hc2939fa0, 32'hc2708e82, 32'hc13b54b5, 32'hc26d3b6e};
test_output[9608:9615] = '{32'h0, 32'h0, 32'h0, 32'h41166d5a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9616:9623] = '{32'hc29089d3, 32'h42b30194, 32'h427baa38, 32'hc2c3087e, 32'h41eff618, 32'hc1987a1b, 32'h42c53c5d, 32'h421323d4};
test_output[9616:9623] = '{32'h0, 32'h42b30194, 32'h427baa38, 32'h0, 32'h41eff618, 32'h0, 32'h42c53c5d, 32'h421323d4};
test_input[9624:9631] = '{32'h41e59725, 32'h4298fa61, 32'h40da7ac8, 32'h423d13f6, 32'h403e2aef, 32'h42b04ec2, 32'hc292ca58, 32'h423ae26d};
test_output[9624:9631] = '{32'h41e59725, 32'h4298fa61, 32'h40da7ac8, 32'h423d13f6, 32'h403e2aef, 32'h42b04ec2, 32'h0, 32'h423ae26d};
test_input[9632:9639] = '{32'h4229e653, 32'hc1577134, 32'h425485ed, 32'hc1e992d7, 32'h42a6f945, 32'hc25ef730, 32'hc23aa11c, 32'hc1e5dc15};
test_output[9632:9639] = '{32'h4229e653, 32'h0, 32'h425485ed, 32'h0, 32'h42a6f945, 32'h0, 32'h0, 32'h0};
test_input[9640:9647] = '{32'hc2928af6, 32'hc2129e22, 32'hc1089f99, 32'hc2b1a94b, 32'hc2a35a96, 32'h41de3923, 32'hc1bab5b4, 32'hc1d108ca};
test_output[9640:9647] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41de3923, 32'h0, 32'h0};
test_input[9648:9655] = '{32'h42bff1ba, 32'hc27689b4, 32'hc2937466, 32'h42bd9654, 32'hc19780dd, 32'hbf23f0f9, 32'h42a6c574, 32'h40f73c0d};
test_output[9648:9655] = '{32'h42bff1ba, 32'h0, 32'h0, 32'h42bd9654, 32'h0, 32'h0, 32'h42a6c574, 32'h40f73c0d};
test_input[9656:9663] = '{32'h4288e872, 32'h4259c8f0, 32'hc2418ed8, 32'h42865ab9, 32'hc2bcf0e3, 32'hc162ab35, 32'h42a45adb, 32'h42b410c9};
test_output[9656:9663] = '{32'h4288e872, 32'h4259c8f0, 32'h0, 32'h42865ab9, 32'h0, 32'h0, 32'h42a45adb, 32'h42b410c9};
test_input[9664:9671] = '{32'h40a44a4b, 32'h4143c7c3, 32'hc12f9fb1, 32'h42a6cfba, 32'h428aee45, 32'h41b7e14c, 32'hc2a5f8ba, 32'h429c3fef};
test_output[9664:9671] = '{32'h40a44a4b, 32'h4143c7c3, 32'h0, 32'h42a6cfba, 32'h428aee45, 32'h41b7e14c, 32'h0, 32'h429c3fef};
test_input[9672:9679] = '{32'hc2764f91, 32'h424a2548, 32'h423d3c50, 32'hc2b284c0, 32'hc13f0100, 32'hc21af8b8, 32'h414dbf95, 32'h412e5b8a};
test_output[9672:9679] = '{32'h0, 32'h424a2548, 32'h423d3c50, 32'h0, 32'h0, 32'h0, 32'h414dbf95, 32'h412e5b8a};
test_input[9680:9687] = '{32'h3fc3640b, 32'hc1a7b6ac, 32'h41acb2f9, 32'hbea17448, 32'hc2b8ccb2, 32'h42b9a10e, 32'h42c31e31, 32'hc248274e};
test_output[9680:9687] = '{32'h3fc3640b, 32'h0, 32'h41acb2f9, 32'h0, 32'h0, 32'h42b9a10e, 32'h42c31e31, 32'h0};
test_input[9688:9695] = '{32'hc27e2d73, 32'h422d9dee, 32'hc2b1705c, 32'hc1a75f42, 32'h42c42621, 32'hc126be23, 32'hbd81d2ba, 32'h422fba14};
test_output[9688:9695] = '{32'h0, 32'h422d9dee, 32'h0, 32'h0, 32'h42c42621, 32'h0, 32'h0, 32'h422fba14};
test_input[9696:9703] = '{32'hc2ada0d3, 32'hc29c5363, 32'hc08685d8, 32'h42b89d95, 32'h42980039, 32'hc13730b8, 32'hc16ae26b, 32'h4294ab36};
test_output[9696:9703] = '{32'h0, 32'h0, 32'h0, 32'h42b89d95, 32'h42980039, 32'h0, 32'h0, 32'h4294ab36};
test_input[9704:9711] = '{32'hc27dad3e, 32'hc2678950, 32'hc1910c98, 32'h41296727, 32'h420fbde4, 32'hc2243bac, 32'h428cb8ca, 32'h4155148c};
test_output[9704:9711] = '{32'h0, 32'h0, 32'h0, 32'h41296727, 32'h420fbde4, 32'h0, 32'h428cb8ca, 32'h4155148c};
test_input[9712:9719] = '{32'h42138253, 32'h3ff86a45, 32'h4206341d, 32'hc2513ddc, 32'hc2aa30db, 32'hc2281f03, 32'h3f7f9d30, 32'hc1ee6dba};
test_output[9712:9719] = '{32'h42138253, 32'h3ff86a45, 32'h4206341d, 32'h0, 32'h0, 32'h0, 32'h3f7f9d30, 32'h0};
test_input[9720:9727] = '{32'hc244b6a5, 32'h4140e914, 32'hc13c10b7, 32'hc0cb2db5, 32'hc238c608, 32'hc266bb3c, 32'h4234c1dc, 32'h41faf692};
test_output[9720:9727] = '{32'h0, 32'h4140e914, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4234c1dc, 32'h41faf692};
test_input[9728:9735] = '{32'hc2a7033b, 32'hc28edeed, 32'hc221ba18, 32'hc275ade1, 32'hc1cdad87, 32'h42548a62, 32'h42242749, 32'hc10a4e8f};
test_output[9728:9735] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42548a62, 32'h42242749, 32'h0};
test_input[9736:9743] = '{32'hc27d2c9a, 32'h42736e6f, 32'hc29e9991, 32'h429cdcbd, 32'hc01b67b7, 32'h428c0089, 32'hc20fe48c, 32'h42137627};
test_output[9736:9743] = '{32'h0, 32'h42736e6f, 32'h0, 32'h429cdcbd, 32'h0, 32'h428c0089, 32'h0, 32'h42137627};
test_input[9744:9751] = '{32'hc250bee0, 32'hc2453706, 32'h40fa939a, 32'h3fe7ebca, 32'h41df2e40, 32'h41f945b2, 32'hc20afc5b, 32'h42a25e53};
test_output[9744:9751] = '{32'h0, 32'h0, 32'h40fa939a, 32'h3fe7ebca, 32'h41df2e40, 32'h41f945b2, 32'h0, 32'h42a25e53};
test_input[9752:9759] = '{32'h41ccd61f, 32'h41b4e820, 32'hc1d69ffc, 32'h427352bf, 32'hc1613d86, 32'hc286772c, 32'hc11b2818, 32'hc1908bc7};
test_output[9752:9759] = '{32'h41ccd61f, 32'h41b4e820, 32'h0, 32'h427352bf, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9760:9767] = '{32'h41a5fae5, 32'hc11b03d7, 32'h41a2290f, 32'h42327ac1, 32'h42c5c2eb, 32'hc2b294b0, 32'h423cc510, 32'h42925f41};
test_output[9760:9767] = '{32'h41a5fae5, 32'h0, 32'h41a2290f, 32'h42327ac1, 32'h42c5c2eb, 32'h0, 32'h423cc510, 32'h42925f41};
test_input[9768:9775] = '{32'hc2491e0f, 32'h41babce5, 32'h410f1e73, 32'h42152df7, 32'hc156e891, 32'h409fe4bf, 32'h42b672ca, 32'h406f8de4};
test_output[9768:9775] = '{32'h0, 32'h41babce5, 32'h410f1e73, 32'h42152df7, 32'h0, 32'h409fe4bf, 32'h42b672ca, 32'h406f8de4};
test_input[9776:9783] = '{32'h40c1dd86, 32'h42c2340e, 32'hc290e7b6, 32'h4268afa7, 32'h426d9dca, 32'hc12a3305, 32'hc2a386fb, 32'h4186791a};
test_output[9776:9783] = '{32'h40c1dd86, 32'h42c2340e, 32'h0, 32'h4268afa7, 32'h426d9dca, 32'h0, 32'h0, 32'h4186791a};
test_input[9784:9791] = '{32'hc288016c, 32'h42937bf7, 32'hc1436114, 32'hc23b3144, 32'hc1bcd5f4, 32'h42b1d17e, 32'h427cc0d6, 32'h41aff9ed};
test_output[9784:9791] = '{32'h0, 32'h42937bf7, 32'h0, 32'h0, 32'h0, 32'h42b1d17e, 32'h427cc0d6, 32'h41aff9ed};
test_input[9792:9799] = '{32'hc2ab6781, 32'h4078ce27, 32'h414607b5, 32'h4243b95d, 32'h42c00346, 32'h42906c77, 32'hc21915fd, 32'hc29662d6};
test_output[9792:9799] = '{32'h0, 32'h4078ce27, 32'h414607b5, 32'h4243b95d, 32'h42c00346, 32'h42906c77, 32'h0, 32'h0};
test_input[9800:9807] = '{32'h4226ffda, 32'h425415e0, 32'hc2b49e88, 32'h426594a2, 32'hc295f133, 32'h428b23ae, 32'hc231df2e, 32'h42a6619b};
test_output[9800:9807] = '{32'h4226ffda, 32'h425415e0, 32'h0, 32'h426594a2, 32'h0, 32'h428b23ae, 32'h0, 32'h42a6619b};
test_input[9808:9815] = '{32'hc0140129, 32'h421152a0, 32'hc2aa8e69, 32'hc26da0e4, 32'hc2be6db6, 32'hc2866aa8, 32'hc228b43b, 32'h42482bca};
test_output[9808:9815] = '{32'h0, 32'h421152a0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42482bca};
test_input[9816:9823] = '{32'h42a9ca2c, 32'hc14f5833, 32'h41d99b8f, 32'h4206cd91, 32'h4237679e, 32'h41ace821, 32'h426048e3, 32'hc228cef0};
test_output[9816:9823] = '{32'h42a9ca2c, 32'h0, 32'h41d99b8f, 32'h4206cd91, 32'h4237679e, 32'h41ace821, 32'h426048e3, 32'h0};
test_input[9824:9831] = '{32'h42943d3a, 32'hc2a7a09d, 32'hc1c39f85, 32'hc1654dc7, 32'hc2292147, 32'hc2836c7e, 32'h42180c88, 32'hc17099f4};
test_output[9824:9831] = '{32'h42943d3a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42180c88, 32'h0};
test_input[9832:9839] = '{32'h4082fd5f, 32'hc1232b9c, 32'h4254e2f5, 32'hc207ed70, 32'hc1d1554d, 32'hc10e0fe6, 32'hc2224fd9, 32'h4147dc53};
test_output[9832:9839] = '{32'h4082fd5f, 32'h0, 32'h4254e2f5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4147dc53};
test_input[9840:9847] = '{32'h429d8964, 32'h41d5401e, 32'hc0976ec8, 32'hc200b4cd, 32'hc1d0853f, 32'h426b5d6e, 32'hc28a128d, 32'hc0bc1675};
test_output[9840:9847] = '{32'h429d8964, 32'h41d5401e, 32'h0, 32'h0, 32'h0, 32'h426b5d6e, 32'h0, 32'h0};
test_input[9848:9855] = '{32'hc295482e, 32'h421ebd92, 32'hc2702d00, 32'hc26f1059, 32'h428418a7, 32'h4260a280, 32'h42158c13, 32'h41792fba};
test_output[9848:9855] = '{32'h0, 32'h421ebd92, 32'h0, 32'h0, 32'h428418a7, 32'h4260a280, 32'h42158c13, 32'h41792fba};
test_input[9856:9863] = '{32'hc2ba987e, 32'hc182255b, 32'h421df9a5, 32'h41588e6f, 32'h42bbd141, 32'h42aae97c, 32'h42adff90, 32'hc25c9ef2};
test_output[9856:9863] = '{32'h0, 32'h0, 32'h421df9a5, 32'h41588e6f, 32'h42bbd141, 32'h42aae97c, 32'h42adff90, 32'h0};
test_input[9864:9871] = '{32'hc22503fd, 32'hc2bf54f9, 32'h41e39bc7, 32'hc1b57f63, 32'h42833f76, 32'h41e5fcee, 32'h4243a306, 32'hc24e34e8};
test_output[9864:9871] = '{32'h0, 32'h0, 32'h41e39bc7, 32'h0, 32'h42833f76, 32'h41e5fcee, 32'h4243a306, 32'h0};
test_input[9872:9879] = '{32'hc28e5528, 32'h41be441f, 32'hc070ba59, 32'hc2b804ca, 32'h4278c15d, 32'h4296056f, 32'h4198c46e, 32'h4096c4d2};
test_output[9872:9879] = '{32'h0, 32'h41be441f, 32'h0, 32'h0, 32'h4278c15d, 32'h4296056f, 32'h4198c46e, 32'h4096c4d2};
test_input[9880:9887] = '{32'hc1abf514, 32'h4238e2da, 32'h426b9d8d, 32'h42c44054, 32'h42b33eee, 32'hc280eb10, 32'hc2c6c8d6, 32'hc1e2b082};
test_output[9880:9887] = '{32'h0, 32'h4238e2da, 32'h426b9d8d, 32'h42c44054, 32'h42b33eee, 32'h0, 32'h0, 32'h0};
test_input[9888:9895] = '{32'hc2026924, 32'h40365c5c, 32'hc1eb60ee, 32'h415d93d1, 32'hc210ebee, 32'hc1eb6bfd, 32'h428a848b, 32'hc1ee45bb};
test_output[9888:9895] = '{32'h0, 32'h40365c5c, 32'h0, 32'h415d93d1, 32'h0, 32'h0, 32'h428a848b, 32'h0};
test_input[9896:9903] = '{32'h4279c275, 32'hc2b1466d, 32'h41a55f20, 32'hc236bb42, 32'h42a238e3, 32'h42c5109d, 32'h42ad00e5, 32'hc2255ba3};
test_output[9896:9903] = '{32'h4279c275, 32'h0, 32'h41a55f20, 32'h0, 32'h42a238e3, 32'h42c5109d, 32'h42ad00e5, 32'h0};
test_input[9904:9911] = '{32'h40f8f97c, 32'h4201f5c7, 32'h42ba5c87, 32'h42849203, 32'h425d3057, 32'h41c5206b, 32'hc2a34eaf, 32'hc09a2f38};
test_output[9904:9911] = '{32'h40f8f97c, 32'h4201f5c7, 32'h42ba5c87, 32'h42849203, 32'h425d3057, 32'h41c5206b, 32'h0, 32'h0};
test_input[9912:9919] = '{32'hc2afaeff, 32'h4205f733, 32'h41b4edd4, 32'hc24f0583, 32'h41cbaa92, 32'hc235cf20, 32'h425ef9b3, 32'h4232f7ee};
test_output[9912:9919] = '{32'h0, 32'h4205f733, 32'h41b4edd4, 32'h0, 32'h41cbaa92, 32'h0, 32'h425ef9b3, 32'h4232f7ee};
test_input[9920:9927] = '{32'h4207e8b5, 32'hc2c17b16, 32'hc2859c03, 32'h4242197b, 32'hbf8069d6, 32'h4142714a, 32'h41a71550, 32'h41a15078};
test_output[9920:9927] = '{32'h4207e8b5, 32'h0, 32'h0, 32'h4242197b, 32'h0, 32'h4142714a, 32'h41a71550, 32'h41a15078};
test_input[9928:9935] = '{32'hc2030574, 32'hc2bd21c0, 32'hc212028a, 32'hc262123d, 32'hc21f2776, 32'h424d259c, 32'hc2af9b9e, 32'hc216fed5};
test_output[9928:9935] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h424d259c, 32'h0, 32'h0};
test_input[9936:9943] = '{32'hc045d897, 32'h4249c47b, 32'h42a3849f, 32'h42c03c1b, 32'hc1a2bbc9, 32'hc1a0462e, 32'h42420c5c, 32'hc2be97dc};
test_output[9936:9943] = '{32'h0, 32'h4249c47b, 32'h42a3849f, 32'h42c03c1b, 32'h0, 32'h0, 32'h42420c5c, 32'h0};
test_input[9944:9951] = '{32'hc21011e1, 32'h4258328e, 32'hc2311181, 32'h41365eab, 32'h425ee1f9, 32'h42261b21, 32'h423016a3, 32'h428dddf9};
test_output[9944:9951] = '{32'h0, 32'h4258328e, 32'h0, 32'h41365eab, 32'h425ee1f9, 32'h42261b21, 32'h423016a3, 32'h428dddf9};
test_input[9952:9959] = '{32'h3f90a806, 32'hc18202ba, 32'h42a28f1e, 32'hc08865bd, 32'hc20367b5, 32'h4280cc19, 32'hc1e25479, 32'hc267f291};
test_output[9952:9959] = '{32'h3f90a806, 32'h0, 32'h42a28f1e, 32'h0, 32'h0, 32'h4280cc19, 32'h0, 32'h0};
test_input[9960:9967] = '{32'hc00bc088, 32'hc2913df2, 32'h410d20cc, 32'hc2af07c0, 32'hc1095dff, 32'h41b56034, 32'h4258158b, 32'h41c7496e};
test_output[9960:9967] = '{32'h0, 32'h0, 32'h410d20cc, 32'h0, 32'h0, 32'h41b56034, 32'h4258158b, 32'h41c7496e};
test_input[9968:9975] = '{32'hc2a3ed75, 32'h400fd487, 32'h420cdf15, 32'h4296c137, 32'hc1c9364a, 32'hbfb9632a, 32'h418c53cc, 32'h42bdaefa};
test_output[9968:9975] = '{32'h0, 32'h400fd487, 32'h420cdf15, 32'h4296c137, 32'h0, 32'h0, 32'h418c53cc, 32'h42bdaefa};
test_input[9976:9983] = '{32'hc2b79bd5, 32'h427ec7e8, 32'h4189470c, 32'h42507e8f, 32'hc27d038d, 32'h41832f88, 32'hc108685c, 32'h41a02ee0};
test_output[9976:9983] = '{32'h0, 32'h427ec7e8, 32'h4189470c, 32'h42507e8f, 32'h0, 32'h41832f88, 32'h0, 32'h41a02ee0};
test_input[9984:9991] = '{32'hc286a7f1, 32'h3c811107, 32'hc20ed0ec, 32'h426878ae, 32'h42abcb48, 32'h42424330, 32'hc1ef4a1d, 32'h4282ac1b};
test_output[9984:9991] = '{32'h0, 32'h3c811107, 32'h0, 32'h426878ae, 32'h42abcb48, 32'h42424330, 32'h0, 32'h4282ac1b};
test_input[9992:9999] = '{32'h4181f581, 32'hc24bb223, 32'h426b76aa, 32'hc1cd4658, 32'hbf55f23d, 32'h42a72a31, 32'h42956810, 32'hc296bb6d};
test_output[9992:9999] = '{32'h4181f581, 32'h0, 32'h426b76aa, 32'h0, 32'h0, 32'h42a72a31, 32'h42956810, 32'h0};
test_input[10000:10007] = '{32'h420720ec, 32'hc14ff3e0, 32'hc20777fe, 32'h425369a4, 32'h3f8e45a1, 32'h42136d78, 32'h42be81ae, 32'hc21e46fb};
test_output[10000:10007] = '{32'h420720ec, 32'h0, 32'h0, 32'h425369a4, 32'h3f8e45a1, 32'h42136d78, 32'h42be81ae, 32'h0};
test_input[10008:10015] = '{32'hc23950bf, 32'hc212040c, 32'hc28430fc, 32'h425179fb, 32'hc2b3adba, 32'h42191e72, 32'hc0ae79b6, 32'h42773a7d};
test_output[10008:10015] = '{32'h0, 32'h0, 32'h0, 32'h425179fb, 32'h0, 32'h42191e72, 32'h0, 32'h42773a7d};
test_input[10016:10023] = '{32'hc09c6963, 32'h42260ac0, 32'h402a9f1a, 32'h40bab673, 32'h4234f42a, 32'h408f213b, 32'h3dd1169c, 32'hc2508777};
test_output[10016:10023] = '{32'h0, 32'h42260ac0, 32'h402a9f1a, 32'h40bab673, 32'h4234f42a, 32'h408f213b, 32'h3dd1169c, 32'h0};
test_input[10024:10031] = '{32'hc23f3fcf, 32'h40a91063, 32'hc2aee73e, 32'h42c7c59b, 32'hc2c6acc0, 32'h41a780a2, 32'h429f39ea, 32'h4277078c};
test_output[10024:10031] = '{32'h0, 32'h40a91063, 32'h0, 32'h42c7c59b, 32'h0, 32'h41a780a2, 32'h429f39ea, 32'h4277078c};
test_input[10032:10039] = '{32'hc28c5008, 32'hc29a713c, 32'hc1c96c02, 32'h420cd1ac, 32'hc2ac1e8f, 32'h428e3aff, 32'hc2632704, 32'h41a6f8f0};
test_output[10032:10039] = '{32'h0, 32'h0, 32'h0, 32'h420cd1ac, 32'h0, 32'h428e3aff, 32'h0, 32'h41a6f8f0};
test_input[10040:10047] = '{32'hc27106f0, 32'hc2ac8091, 32'h4246b4a8, 32'h41d2fbf4, 32'h426e614b, 32'h42031ea5, 32'hc2abe508, 32'h41c9c1b7};
test_output[10040:10047] = '{32'h0, 32'h0, 32'h4246b4a8, 32'h41d2fbf4, 32'h426e614b, 32'h42031ea5, 32'h0, 32'h41c9c1b7};
test_input[10048:10055] = '{32'hc2bfdde6, 32'h42096800, 32'h42a1e5a3, 32'h41ccd904, 32'h428b7ca6, 32'h42bf50a6, 32'h4258aac4, 32'hc1728350};
test_output[10048:10055] = '{32'h0, 32'h42096800, 32'h42a1e5a3, 32'h41ccd904, 32'h428b7ca6, 32'h42bf50a6, 32'h4258aac4, 32'h0};
test_input[10056:10063] = '{32'hc1fd0fbd, 32'hc1c6f51c, 32'hc0e02503, 32'h41510aa1, 32'h4291f47d, 32'hc2b27f82, 32'h42a6d5a8, 32'h420793ce};
test_output[10056:10063] = '{32'h0, 32'h0, 32'h0, 32'h41510aa1, 32'h4291f47d, 32'h0, 32'h42a6d5a8, 32'h420793ce};
test_input[10064:10071] = '{32'h429a0e6d, 32'hc2ad57ad, 32'hc29d26dc, 32'h42130e18, 32'hc292f2f1, 32'h42277816, 32'h42757b2f, 32'hc246f0a3};
test_output[10064:10071] = '{32'h429a0e6d, 32'h0, 32'h0, 32'h42130e18, 32'h0, 32'h42277816, 32'h42757b2f, 32'h0};
test_input[10072:10079] = '{32'hc2c4f6e6, 32'hc24542e9, 32'h42b1bf1d, 32'hc2a0fc15, 32'h42180753, 32'h41a23f35, 32'hc27d0c62, 32'h428c8f3e};
test_output[10072:10079] = '{32'h0, 32'h0, 32'h42b1bf1d, 32'h0, 32'h42180753, 32'h41a23f35, 32'h0, 32'h428c8f3e};
test_input[10080:10087] = '{32'hc237e7a0, 32'h416a367e, 32'h41a5da18, 32'hc20019bf, 32'hc0a63ace, 32'h41b7db2f, 32'h41dfd266, 32'hc1dde0a9};
test_output[10080:10087] = '{32'h0, 32'h416a367e, 32'h41a5da18, 32'h0, 32'h0, 32'h41b7db2f, 32'h41dfd266, 32'h0};
test_input[10088:10095] = '{32'h41f2684e, 32'hc2464c23, 32'h41e213d3, 32'hc268014c, 32'hc259e8ee, 32'h4228bc24, 32'h4284df2d, 32'hc0712661};
test_output[10088:10095] = '{32'h41f2684e, 32'h0, 32'h41e213d3, 32'h0, 32'h0, 32'h4228bc24, 32'h4284df2d, 32'h0};
test_input[10096:10103] = '{32'h421c4206, 32'h42c392a7, 32'hc291f84f, 32'hc1ec8ce1, 32'h4294a9ef, 32'h429e1807, 32'h42bf945a, 32'h42002164};
test_output[10096:10103] = '{32'h421c4206, 32'h42c392a7, 32'h0, 32'h0, 32'h4294a9ef, 32'h429e1807, 32'h42bf945a, 32'h42002164};
test_input[10104:10111] = '{32'h3e36d533, 32'h4116aca4, 32'h4246774f, 32'h424b62ba, 32'hc231099b, 32'hc2a44f17, 32'h41c715f1, 32'hc2b67980};
test_output[10104:10111] = '{32'h3e36d533, 32'h4116aca4, 32'h4246774f, 32'h424b62ba, 32'h0, 32'h0, 32'h41c715f1, 32'h0};
test_input[10112:10119] = '{32'hc2a1da7c, 32'hc089efcc, 32'hc21ec046, 32'h41443a74, 32'hc29e82e1, 32'hc2a3d3ca, 32'h4275d46e, 32'h4275bbb4};
test_output[10112:10119] = '{32'h0, 32'h0, 32'h0, 32'h41443a74, 32'h0, 32'h0, 32'h4275d46e, 32'h4275bbb4};
test_input[10120:10127] = '{32'h4290df5c, 32'h429868b4, 32'h42bdb17b, 32'hc12a7801, 32'hc2214397, 32'hc288909f, 32'hc2a2c00f, 32'h424718ce};
test_output[10120:10127] = '{32'h4290df5c, 32'h429868b4, 32'h42bdb17b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h424718ce};
test_input[10128:10135] = '{32'hc275d6fb, 32'h42a9329b, 32'h422350ac, 32'hc1c065c3, 32'hc2a63306, 32'hc2949ff7, 32'h42a72be3, 32'hc1d59328};
test_output[10128:10135] = '{32'h0, 32'h42a9329b, 32'h422350ac, 32'h0, 32'h0, 32'h0, 32'h42a72be3, 32'h0};
test_input[10136:10143] = '{32'hbf91933d, 32'hc20506f2, 32'h423ec41b, 32'hc01e4cfa, 32'h424c21b5, 32'h42232aa6, 32'hc004dd60, 32'hbee824c9};
test_output[10136:10143] = '{32'h0, 32'h0, 32'h423ec41b, 32'h0, 32'h424c21b5, 32'h42232aa6, 32'h0, 32'h0};
test_input[10144:10151] = '{32'h41ad5a3c, 32'h42499506, 32'h41e29fc5, 32'hc1b4b8f9, 32'h4228b3ee, 32'h42695924, 32'hc1e1b8bc, 32'hc2807392};
test_output[10144:10151] = '{32'h41ad5a3c, 32'h42499506, 32'h41e29fc5, 32'h0, 32'h4228b3ee, 32'h42695924, 32'h0, 32'h0};
test_input[10152:10159] = '{32'hc1ca566b, 32'hc2604a3b, 32'hc25a503b, 32'h4225f459, 32'hc1c0b0a6, 32'h42ad385e, 32'hc251a426, 32'h410afea9};
test_output[10152:10159] = '{32'h0, 32'h0, 32'h0, 32'h4225f459, 32'h0, 32'h42ad385e, 32'h0, 32'h410afea9};
test_input[10160:10167] = '{32'h422da930, 32'hc291dcef, 32'h3fa9722d, 32'h429f7bc4, 32'h42c62554, 32'hc24da02d, 32'h42b53565, 32'hc1f984ca};
test_output[10160:10167] = '{32'h422da930, 32'h0, 32'h3fa9722d, 32'h429f7bc4, 32'h42c62554, 32'h0, 32'h42b53565, 32'h0};
test_input[10168:10175] = '{32'h42ac710f, 32'hc1add68c, 32'hc274dde2, 32'hbf642b21, 32'h40457751, 32'h425ec041, 32'h42c49d62, 32'hc115be99};
test_output[10168:10175] = '{32'h42ac710f, 32'h0, 32'h0, 32'h0, 32'h40457751, 32'h425ec041, 32'h42c49d62, 32'h0};
test_input[10176:10183] = '{32'hc1fa48bf, 32'h42449fdf, 32'h42832e9a, 32'hc18aecdf, 32'hc22f4cdf, 32'hbfa2e8e7, 32'h4255f07b, 32'h41dc1958};
test_output[10176:10183] = '{32'h0, 32'h42449fdf, 32'h42832e9a, 32'h0, 32'h0, 32'h0, 32'h4255f07b, 32'h41dc1958};
test_input[10184:10191] = '{32'hbfe85b87, 32'h42b988ac, 32'hc200755d, 32'hc2c2c904, 32'h3f78aa79, 32'hc1bdfad3, 32'hc27226bb, 32'h42239c47};
test_output[10184:10191] = '{32'h0, 32'h42b988ac, 32'h0, 32'h0, 32'h3f78aa79, 32'h0, 32'h0, 32'h42239c47};
test_input[10192:10199] = '{32'hc2b41817, 32'h42b9f542, 32'hc2bd62f8, 32'hc2a73bfb, 32'h42842a7b, 32'hc0ca0c47, 32'hc287da3f, 32'hc27e3584};
test_output[10192:10199] = '{32'h0, 32'h42b9f542, 32'h0, 32'h0, 32'h42842a7b, 32'h0, 32'h0, 32'h0};
test_input[10200:10207] = '{32'hc1eaa962, 32'h418daf42, 32'hc2958bb4, 32'hc19f0382, 32'hc28080f3, 32'hc2b5bf80, 32'h422f4dd5, 32'hc101e246};
test_output[10200:10207] = '{32'h0, 32'h418daf42, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422f4dd5, 32'h0};
test_input[10208:10215] = '{32'h427db35d, 32'h42c00b76, 32'hc20f4f7e, 32'hc26ea702, 32'hc215442f, 32'hc2a4dc9a, 32'h426c885e, 32'hc2af9081};
test_output[10208:10215] = '{32'h427db35d, 32'h42c00b76, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426c885e, 32'h0};
test_input[10216:10223] = '{32'h42c1f98c, 32'h425be9c9, 32'h42a3db7c, 32'hc2c200b1, 32'hc0dd56ac, 32'hc1a2bd7e, 32'hc27e5232, 32'h428a9e22};
test_output[10216:10223] = '{32'h42c1f98c, 32'h425be9c9, 32'h42a3db7c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428a9e22};
test_input[10224:10231] = '{32'hc0a90b78, 32'h42482eca, 32'h42c3469c, 32'hc2bea46f, 32'h42b58b39, 32'h41372d4d, 32'h4219fff5, 32'h4233aa7f};
test_output[10224:10231] = '{32'h0, 32'h42482eca, 32'h42c3469c, 32'h0, 32'h42b58b39, 32'h41372d4d, 32'h4219fff5, 32'h4233aa7f};
test_input[10232:10239] = '{32'hc285def1, 32'h42a184b6, 32'h42b252c5, 32'h41e81627, 32'hc12afbca, 32'hc24cc2bd, 32'hc29b3e08, 32'hc24866f1};
test_output[10232:10239] = '{32'h0, 32'h42a184b6, 32'h42b252c5, 32'h41e81627, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10240:10247] = '{32'h3f179129, 32'hc258b770, 32'hc2ac38d2, 32'h42a04ff9, 32'hc2424d6c, 32'hc2128cb8, 32'hc2772b37, 32'h426b6ee4};
test_output[10240:10247] = '{32'h3f179129, 32'h0, 32'h0, 32'h42a04ff9, 32'h0, 32'h0, 32'h0, 32'h426b6ee4};
test_input[10248:10255] = '{32'hc1317de6, 32'hc2c12797, 32'hc1186346, 32'h414b40be, 32'h420b9c97, 32'hc2944767, 32'hc24d6319, 32'h42a64fc6};
test_output[10248:10255] = '{32'h0, 32'h0, 32'h0, 32'h414b40be, 32'h420b9c97, 32'h0, 32'h0, 32'h42a64fc6};
test_input[10256:10263] = '{32'hc2863973, 32'hc2391b89, 32'hc239f28e, 32'h42752fa7, 32'h4295f16a, 32'h42a2682a, 32'hc296ecbe, 32'hc1a7e541};
test_output[10256:10263] = '{32'h0, 32'h0, 32'h0, 32'h42752fa7, 32'h4295f16a, 32'h42a2682a, 32'h0, 32'h0};
test_input[10264:10271] = '{32'h422447ab, 32'h4208e3bd, 32'hc2baef38, 32'h421909f6, 32'hc2af0e92, 32'h42b17e2e, 32'h421a021c, 32'h4121c858};
test_output[10264:10271] = '{32'h422447ab, 32'h4208e3bd, 32'h0, 32'h421909f6, 32'h0, 32'h42b17e2e, 32'h421a021c, 32'h4121c858};
test_input[10272:10279] = '{32'h429adf40, 32'hc22c6bba, 32'hc0f15574, 32'hc260014b, 32'hc1426389, 32'hc240283d, 32'hc29929a5, 32'hc2635853};
test_output[10272:10279] = '{32'h429adf40, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10280:10287] = '{32'hc154ca38, 32'h428ea4c7, 32'hc2a49fec, 32'h3f620c61, 32'h40d56685, 32'hc1ba3d33, 32'hc1d6e397, 32'h429d6754};
test_output[10280:10287] = '{32'h0, 32'h428ea4c7, 32'h0, 32'h3f620c61, 32'h40d56685, 32'h0, 32'h0, 32'h429d6754};
test_input[10288:10295] = '{32'hc2423e5d, 32'h410f3874, 32'h422de4d8, 32'h42a11f67, 32'hc04865f2, 32'hc29f4afc, 32'h42c0af37, 32'hc2614272};
test_output[10288:10295] = '{32'h0, 32'h410f3874, 32'h422de4d8, 32'h42a11f67, 32'h0, 32'h0, 32'h42c0af37, 32'h0};
test_input[10296:10303] = '{32'h420042e5, 32'hc1bd93f0, 32'h429663a3, 32'h42bfc85e, 32'hc2bf3297, 32'hc2a92174, 32'hc290e0da, 32'h42426acf};
test_output[10296:10303] = '{32'h420042e5, 32'h0, 32'h429663a3, 32'h42bfc85e, 32'h0, 32'h0, 32'h0, 32'h42426acf};
test_input[10304:10311] = '{32'h42b24a79, 32'hc2b0b7a4, 32'h418ad13d, 32'hc1a7cbb4, 32'hc18e4234, 32'h418918e3, 32'h4294eba2, 32'hc231663e};
test_output[10304:10311] = '{32'h42b24a79, 32'h0, 32'h418ad13d, 32'h0, 32'h0, 32'h418918e3, 32'h4294eba2, 32'h0};
test_input[10312:10319] = '{32'h4293d3c8, 32'hc0235acf, 32'hc2a54441, 32'hc125b980, 32'h41d514c2, 32'hbf2c3eb2, 32'hc23f144f, 32'hc1a524af};
test_output[10312:10319] = '{32'h4293d3c8, 32'h0, 32'h0, 32'h0, 32'h41d514c2, 32'h0, 32'h0, 32'h0};
test_input[10320:10327] = '{32'hc25a4213, 32'hc21c2a0c, 32'h41852423, 32'h41cb9a70, 32'hc23afdf1, 32'h42046919, 32'hc2200a29, 32'h41ad46d0};
test_output[10320:10327] = '{32'h0, 32'h0, 32'h41852423, 32'h41cb9a70, 32'h0, 32'h42046919, 32'h0, 32'h41ad46d0};
test_input[10328:10335] = '{32'h4228534e, 32'hc2977a4f, 32'h4257eb70, 32'hc142991c, 32'h40333915, 32'hc28de15e, 32'hc2abe610, 32'h41e9f79e};
test_output[10328:10335] = '{32'h4228534e, 32'h0, 32'h4257eb70, 32'h0, 32'h40333915, 32'h0, 32'h0, 32'h41e9f79e};
test_input[10336:10343] = '{32'hc2795367, 32'h42c1a248, 32'hc20ab103, 32'h4210fc09, 32'hc2b32c81, 32'hc2a12826, 32'h428d6783, 32'h420c5270};
test_output[10336:10343] = '{32'h0, 32'h42c1a248, 32'h0, 32'h4210fc09, 32'h0, 32'h0, 32'h428d6783, 32'h420c5270};
test_input[10344:10351] = '{32'hc27b2f65, 32'h4281515f, 32'hc120a3ea, 32'hc1d002f9, 32'h42855d60, 32'h4205177d, 32'hc2c66ff9, 32'hc29dbca3};
test_output[10344:10351] = '{32'h0, 32'h4281515f, 32'h0, 32'h0, 32'h42855d60, 32'h4205177d, 32'h0, 32'h0};
test_input[10352:10359] = '{32'h42546be7, 32'hc166f0a2, 32'h42a8f8fe, 32'hc209eed9, 32'h42aa87a0, 32'h421f4a81, 32'hc2866080, 32'hc2aed698};
test_output[10352:10359] = '{32'h42546be7, 32'h0, 32'h42a8f8fe, 32'h0, 32'h42aa87a0, 32'h421f4a81, 32'h0, 32'h0};
test_input[10360:10367] = '{32'h426b7882, 32'h42140341, 32'hc1c5b696, 32'hc25e7067, 32'hc28512ad, 32'h4221fe51, 32'hc12e0f15, 32'hc2406d48};
test_output[10360:10367] = '{32'h426b7882, 32'h42140341, 32'h0, 32'h0, 32'h0, 32'h4221fe51, 32'h0, 32'h0};
test_input[10368:10375] = '{32'h41951604, 32'hc16daed2, 32'hc2b0543a, 32'h42950816, 32'hc2964f4d, 32'h41de1220, 32'h4288bbc1, 32'hc2b0642b};
test_output[10368:10375] = '{32'h41951604, 32'h0, 32'h0, 32'h42950816, 32'h0, 32'h41de1220, 32'h4288bbc1, 32'h0};
test_input[10376:10383] = '{32'hc2944d47, 32'hc299e4db, 32'hc284c7c8, 32'hc2a4bf55, 32'hc2749491, 32'hc291a25f, 32'hc29e7725, 32'hc1f023e2};
test_output[10376:10383] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10384:10391] = '{32'h41e892e9, 32'hc1fe10ff, 32'h421c1aac, 32'h41d7b4b5, 32'h424e7015, 32'h429c214a, 32'hc2596429, 32'h41f9a50c};
test_output[10384:10391] = '{32'h41e892e9, 32'h0, 32'h421c1aac, 32'h41d7b4b5, 32'h424e7015, 32'h429c214a, 32'h0, 32'h41f9a50c};
test_input[10392:10399] = '{32'hc16abd2e, 32'hc1f46ecf, 32'h4187bf7f, 32'h411aeb13, 32'h41cff887, 32'hc29db9f9, 32'h427cd29e, 32'hc25ee795};
test_output[10392:10399] = '{32'h0, 32'h0, 32'h4187bf7f, 32'h411aeb13, 32'h41cff887, 32'h0, 32'h427cd29e, 32'h0};
test_input[10400:10407] = '{32'hc0891c11, 32'hc2723f7a, 32'h42a663fa, 32'hbf93f72c, 32'h422a6efc, 32'h4248381d, 32'h420b3dcd, 32'hc28fa1e5};
test_output[10400:10407] = '{32'h0, 32'h0, 32'h42a663fa, 32'h0, 32'h422a6efc, 32'h4248381d, 32'h420b3dcd, 32'h0};
test_input[10408:10415] = '{32'h403c52fb, 32'hc0c5b0e7, 32'h42beac38, 32'h428e910b, 32'hc2a8e5e0, 32'hc2193372, 32'h422e82b7, 32'h41e19df6};
test_output[10408:10415] = '{32'h403c52fb, 32'h0, 32'h42beac38, 32'h428e910b, 32'h0, 32'h0, 32'h422e82b7, 32'h41e19df6};
test_input[10416:10423] = '{32'hc2375c4c, 32'hc2bc39f0, 32'h419019a6, 32'h41d435af, 32'hc2058eaf, 32'h422cc2d9, 32'h42b5bea4, 32'hc1503012};
test_output[10416:10423] = '{32'h0, 32'h0, 32'h419019a6, 32'h41d435af, 32'h0, 32'h422cc2d9, 32'h42b5bea4, 32'h0};
test_input[10424:10431] = '{32'hc2161814, 32'hc1b97037, 32'h42269caa, 32'hc1f3be04, 32'hc29a1c69, 32'hc243353d, 32'h4276e8b6, 32'hc2466e8d};
test_output[10424:10431] = '{32'h0, 32'h0, 32'h42269caa, 32'h0, 32'h0, 32'h0, 32'h4276e8b6, 32'h0};
test_input[10432:10439] = '{32'hc2b934e0, 32'h42856a29, 32'h4282b88d, 32'h402ff88b, 32'h420fa987, 32'hc2c21086, 32'hc18c39e1, 32'hc1e508ce};
test_output[10432:10439] = '{32'h0, 32'h42856a29, 32'h4282b88d, 32'h402ff88b, 32'h420fa987, 32'h0, 32'h0, 32'h0};
test_input[10440:10447] = '{32'h40c00aea, 32'h42295966, 32'hc2b03600, 32'h3fd7b1a1, 32'h42a607a3, 32'h422adc6b, 32'hc215439f, 32'hc0aff999};
test_output[10440:10447] = '{32'h40c00aea, 32'h42295966, 32'h0, 32'h3fd7b1a1, 32'h42a607a3, 32'h422adc6b, 32'h0, 32'h0};
test_input[10448:10455] = '{32'h4143d886, 32'hc2824140, 32'h420370f2, 32'hc1446e20, 32'h419d3d32, 32'hc2830267, 32'hc17efc21, 32'hc2c62361};
test_output[10448:10455] = '{32'h4143d886, 32'h0, 32'h420370f2, 32'h0, 32'h419d3d32, 32'h0, 32'h0, 32'h0};
test_input[10456:10463] = '{32'hc2afffc4, 32'h41014900, 32'h41a33be9, 32'hc1e2966e, 32'hc24cc143, 32'hc025094e, 32'h427b2d27, 32'hc2581d62};
test_output[10456:10463] = '{32'h0, 32'h41014900, 32'h41a33be9, 32'h0, 32'h0, 32'h0, 32'h427b2d27, 32'h0};
test_input[10464:10471] = '{32'h41df6a0f, 32'hbfd9dba9, 32'h4194744a, 32'h41bdcc1b, 32'h41baf7e6, 32'h429410d5, 32'hc1fcfbf8, 32'hc19a4cd9};
test_output[10464:10471] = '{32'h41df6a0f, 32'h0, 32'h4194744a, 32'h41bdcc1b, 32'h41baf7e6, 32'h429410d5, 32'h0, 32'h0};
test_input[10472:10479] = '{32'h4131c988, 32'hc18bcccb, 32'h42887c46, 32'h42698b5a, 32'hc2b00282, 32'hc293ec73, 32'h42b96bb7, 32'h425fce7a};
test_output[10472:10479] = '{32'h4131c988, 32'h0, 32'h42887c46, 32'h42698b5a, 32'h0, 32'h0, 32'h42b96bb7, 32'h425fce7a};
test_input[10480:10487] = '{32'hc29b823d, 32'hc2b257fa, 32'h4207d7a5, 32'hc2820dce, 32'h41102204, 32'h422b82c8, 32'h4280126a, 32'h4172ed06};
test_output[10480:10487] = '{32'h0, 32'h0, 32'h4207d7a5, 32'h0, 32'h41102204, 32'h422b82c8, 32'h4280126a, 32'h4172ed06};
test_input[10488:10495] = '{32'h4265ca46, 32'h42c66f07, 32'h42924c3a, 32'hc25652ed, 32'hc1980c9d, 32'h42098d25, 32'hc1e5461b, 32'h42ac787e};
test_output[10488:10495] = '{32'h4265ca46, 32'h42c66f07, 32'h42924c3a, 32'h0, 32'h0, 32'h42098d25, 32'h0, 32'h42ac787e};
test_input[10496:10503] = '{32'h41671c19, 32'hc21ef9d8, 32'hc2372320, 32'hc15d4675, 32'hc2ad4cb6, 32'hc2ae45bb, 32'h42c0b088, 32'h41581efa};
test_output[10496:10503] = '{32'h41671c19, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c0b088, 32'h41581efa};
test_input[10504:10511] = '{32'hc2c642f3, 32'h428ba53f, 32'h421951e5, 32'h429c3c44, 32'hc213f2de, 32'hc28dbf97, 32'h40c267a7, 32'h41fc685e};
test_output[10504:10511] = '{32'h0, 32'h428ba53f, 32'h421951e5, 32'h429c3c44, 32'h0, 32'h0, 32'h40c267a7, 32'h41fc685e};
test_input[10512:10519] = '{32'hc18e2176, 32'h42a1c2c2, 32'hc24a2c28, 32'hc23bebcd, 32'hc17a2179, 32'h40fec53e, 32'h4292eb5c, 32'hc20195a7};
test_output[10512:10519] = '{32'h0, 32'h42a1c2c2, 32'h0, 32'h0, 32'h0, 32'h40fec53e, 32'h4292eb5c, 32'h0};
test_input[10520:10527] = '{32'h41d35795, 32'hc0bf8958, 32'hc1b5c28d, 32'h429793e5, 32'hc272b36a, 32'h42c56978, 32'hc2a9b566, 32'h42562ab5};
test_output[10520:10527] = '{32'h41d35795, 32'h0, 32'h0, 32'h429793e5, 32'h0, 32'h42c56978, 32'h0, 32'h42562ab5};
test_input[10528:10535] = '{32'h420fc27c, 32'hbda4b540, 32'h4289e1f8, 32'h41101838, 32'hc2b8b3c6, 32'h42461681, 32'h42705022, 32'hc1a7ced3};
test_output[10528:10535] = '{32'h420fc27c, 32'h0, 32'h4289e1f8, 32'h41101838, 32'h0, 32'h42461681, 32'h42705022, 32'h0};
test_input[10536:10543] = '{32'hc2367814, 32'h41af59be, 32'hc2b26440, 32'h42a2087f, 32'h422a01de, 32'hc291f113, 32'h41dec437, 32'h4294effc};
test_output[10536:10543] = '{32'h0, 32'h41af59be, 32'h0, 32'h42a2087f, 32'h422a01de, 32'h0, 32'h41dec437, 32'h4294effc};
test_input[10544:10551] = '{32'hc2be0b60, 32'h42857e1b, 32'h42c0575e, 32'hc2bd048e, 32'hc288455c, 32'hc2684a01, 32'h426a1a13, 32'h42976b65};
test_output[10544:10551] = '{32'h0, 32'h42857e1b, 32'h42c0575e, 32'h0, 32'h0, 32'h0, 32'h426a1a13, 32'h42976b65};
test_input[10552:10559] = '{32'hc2c65d96, 32'hc299df1b, 32'h42aab9cd, 32'hc21cd76e, 32'hc0144899, 32'hc2ae06a5, 32'hc2753feb, 32'h41f0d2ba};
test_output[10552:10559] = '{32'h0, 32'h0, 32'h42aab9cd, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f0d2ba};
test_input[10560:10567] = '{32'h41efd56e, 32'h421ab9c2, 32'hc20ea123, 32'h418b4ed1, 32'h42a42ff0, 32'hc0d01742, 32'hc206e1a2, 32'hc2908287};
test_output[10560:10567] = '{32'h41efd56e, 32'h421ab9c2, 32'h0, 32'h418b4ed1, 32'h42a42ff0, 32'h0, 32'h0, 32'h0};
test_input[10568:10575] = '{32'h4207242a, 32'h4292d263, 32'hc2a17228, 32'hc22b7df8, 32'h41f9e549, 32'hc276ac4f, 32'hc2952a05, 32'h419ecad4};
test_output[10568:10575] = '{32'h4207242a, 32'h4292d263, 32'h0, 32'h0, 32'h41f9e549, 32'h0, 32'h0, 32'h419ecad4};
test_input[10576:10583] = '{32'h4236395d, 32'h3fdac143, 32'hc230e3dc, 32'h4288e758, 32'hc0fe04ad, 32'h42c19149, 32'hbf8a5459, 32'h42499fc0};
test_output[10576:10583] = '{32'h4236395d, 32'h3fdac143, 32'h0, 32'h4288e758, 32'h0, 32'h42c19149, 32'h0, 32'h42499fc0};
test_input[10584:10591] = '{32'hc2910fef, 32'hc0efd255, 32'hc2be82a5, 32'hc2200c92, 32'hc27ec89f, 32'hc232f9e5, 32'h42809a5e, 32'hbf972648};
test_output[10584:10591] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42809a5e, 32'h0};
test_input[10592:10599] = '{32'hc1699ef4, 32'hc2b9ca05, 32'h41ed7aa6, 32'hc2a963bd, 32'hc29fbc7f, 32'h42c54dd6, 32'h42b0a001, 32'h41fd4806};
test_output[10592:10599] = '{32'h0, 32'h0, 32'h41ed7aa6, 32'h0, 32'h0, 32'h42c54dd6, 32'h42b0a001, 32'h41fd4806};
test_input[10600:10607] = '{32'hc27224f7, 32'hc2a2245f, 32'h42b45ae3, 32'h420a2c1c, 32'hc24126a8, 32'hc20971c6, 32'hc2905186, 32'hc1e81446};
test_output[10600:10607] = '{32'h0, 32'h0, 32'h42b45ae3, 32'h420a2c1c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10608:10615] = '{32'h41ca688f, 32'h42aebda1, 32'hc29bc025, 32'hc2301b07, 32'h428fbcc8, 32'h41d5c96a, 32'h42517b8e, 32'hc2a07277};
test_output[10608:10615] = '{32'h41ca688f, 32'h42aebda1, 32'h0, 32'h0, 32'h428fbcc8, 32'h41d5c96a, 32'h42517b8e, 32'h0};
test_input[10616:10623] = '{32'h4299e4f5, 32'hc2ae17d5, 32'hc2c5eb61, 32'hc16b3397, 32'h410f7372, 32'h429168ac, 32'h41d5be73, 32'hc20fc11a};
test_output[10616:10623] = '{32'h4299e4f5, 32'h0, 32'h0, 32'h0, 32'h410f7372, 32'h429168ac, 32'h41d5be73, 32'h0};
test_input[10624:10631] = '{32'hc23c46e6, 32'hc2aef0a6, 32'hc1951675, 32'h42a20396, 32'h427bb2ee, 32'hc2ae8177, 32'h421115da, 32'h411a655b};
test_output[10624:10631] = '{32'h0, 32'h0, 32'h0, 32'h42a20396, 32'h427bb2ee, 32'h0, 32'h421115da, 32'h411a655b};
test_input[10632:10639] = '{32'hc2171482, 32'hc1f4d636, 32'h429a192e, 32'h423f4d40, 32'h42731338, 32'hc203fc8b, 32'hc212034e, 32'h429cc656};
test_output[10632:10639] = '{32'h0, 32'h0, 32'h429a192e, 32'h423f4d40, 32'h42731338, 32'h0, 32'h0, 32'h429cc656};
test_input[10640:10647] = '{32'h41ce1a33, 32'hc214ffe6, 32'hc2a17c83, 32'h41eb71e6, 32'hc2077322, 32'h418d7b1b, 32'h41e86349, 32'h4255539b};
test_output[10640:10647] = '{32'h41ce1a33, 32'h0, 32'h0, 32'h41eb71e6, 32'h0, 32'h418d7b1b, 32'h41e86349, 32'h4255539b};
test_input[10648:10655] = '{32'h41a0e72f, 32'h41d1ede8, 32'h4277a9ea, 32'h42530c8b, 32'hc28842c1, 32'hc2ad9a10, 32'hc1c1c034, 32'h418a3a18};
test_output[10648:10655] = '{32'h41a0e72f, 32'h41d1ede8, 32'h4277a9ea, 32'h42530c8b, 32'h0, 32'h0, 32'h0, 32'h418a3a18};
test_input[10656:10663] = '{32'hc22310f9, 32'h4264fd94, 32'hc24356d6, 32'hc23dcad9, 32'hc0899799, 32'h418c3ee6, 32'h4202cb3d, 32'hc25fc3ed};
test_output[10656:10663] = '{32'h0, 32'h4264fd94, 32'h0, 32'h0, 32'h0, 32'h418c3ee6, 32'h4202cb3d, 32'h0};
test_input[10664:10671] = '{32'hc096386a, 32'hc1d902f0, 32'hc24f481a, 32'hc193d8bb, 32'h4246b66e, 32'h423dceb4, 32'h411b181c, 32'h41b86749};
test_output[10664:10671] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4246b66e, 32'h423dceb4, 32'h411b181c, 32'h41b86749};
test_input[10672:10679] = '{32'hc145309b, 32'hc2660429, 32'hc28aad40, 32'hc28650f0, 32'hc21cb523, 32'h42b7be44, 32'hc26aec43, 32'h42252f59};
test_output[10672:10679] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b7be44, 32'h0, 32'h42252f59};
test_input[10680:10687] = '{32'hc292acc6, 32'h429f19fe, 32'h42aedd19, 32'hc2a1ba35, 32'h42aefad2, 32'h42a79d6b, 32'hc28f356d, 32'hc27e2fd8};
test_output[10680:10687] = '{32'h0, 32'h429f19fe, 32'h42aedd19, 32'h0, 32'h42aefad2, 32'h42a79d6b, 32'h0, 32'h0};
test_input[10688:10695] = '{32'h422f4360, 32'hc223bd53, 32'h424e7670, 32'hc29f41c9, 32'hc23f0896, 32'hc242d890, 32'hc211a394, 32'h4251ab65};
test_output[10688:10695] = '{32'h422f4360, 32'h0, 32'h424e7670, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4251ab65};
test_input[10696:10703] = '{32'h403ea34d, 32'hc234f45d, 32'hc236577e, 32'h42c781f2, 32'h4294dbe1, 32'h4287f98b, 32'h42542465, 32'hc275a890};
test_output[10696:10703] = '{32'h403ea34d, 32'h0, 32'h0, 32'h42c781f2, 32'h4294dbe1, 32'h4287f98b, 32'h42542465, 32'h0};
test_input[10704:10711] = '{32'h42aa8a7a, 32'h423e28d9, 32'hc286174f, 32'h42b21de6, 32'h424d957d, 32'hc22ff593, 32'hc290f29d, 32'hc28c958e};
test_output[10704:10711] = '{32'h42aa8a7a, 32'h423e28d9, 32'h0, 32'h42b21de6, 32'h424d957d, 32'h0, 32'h0, 32'h0};
test_input[10712:10719] = '{32'h415841b5, 32'hc286145e, 32'h42bda600, 32'h429ed003, 32'h42a86444, 32'h428ea7f1, 32'hc154ce06, 32'hc2abf83d};
test_output[10712:10719] = '{32'h415841b5, 32'h0, 32'h42bda600, 32'h429ed003, 32'h42a86444, 32'h428ea7f1, 32'h0, 32'h0};
test_input[10720:10727] = '{32'h4202b54a, 32'hc16b89c1, 32'h41aa8b2d, 32'hbf95041b, 32'h40e69905, 32'h416a3b0a, 32'h425ac565, 32'hc1cc6e94};
test_output[10720:10727] = '{32'h4202b54a, 32'h0, 32'h41aa8b2d, 32'h0, 32'h40e69905, 32'h416a3b0a, 32'h425ac565, 32'h0};
test_input[10728:10735] = '{32'h4189537e, 32'hc20353c5, 32'h41b6971a, 32'h41c4ed7a, 32'hc29335e0, 32'hc221101b, 32'h4268d8a0, 32'h4144bbec};
test_output[10728:10735] = '{32'h4189537e, 32'h0, 32'h41b6971a, 32'h41c4ed7a, 32'h0, 32'h0, 32'h4268d8a0, 32'h4144bbec};
test_input[10736:10743] = '{32'hc23e5572, 32'h421a16a7, 32'h421f49ee, 32'hc2a709c2, 32'hc2986957, 32'hc18d1480, 32'hc27de15d, 32'hc29239b2};
test_output[10736:10743] = '{32'h0, 32'h421a16a7, 32'h421f49ee, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10744:10751] = '{32'h40f84343, 32'hc23e0ed5, 32'h4183d24c, 32'h4135504a, 32'h41f79f59, 32'h406f6f2c, 32'hc2c13dd8, 32'h428cee73};
test_output[10744:10751] = '{32'h40f84343, 32'h0, 32'h4183d24c, 32'h4135504a, 32'h41f79f59, 32'h406f6f2c, 32'h0, 32'h428cee73};
test_input[10752:10759] = '{32'hc2694114, 32'h40f7b1b0, 32'h429158a1, 32'h42324844, 32'hc26266e7, 32'hc212e306, 32'hc2428e26, 32'h4299c10d};
test_output[10752:10759] = '{32'h0, 32'h40f7b1b0, 32'h429158a1, 32'h42324844, 32'h0, 32'h0, 32'h0, 32'h4299c10d};
test_input[10760:10767] = '{32'hc294a78e, 32'hc1e4f491, 32'h408f25a9, 32'h42ae1437, 32'hc2b63dc9, 32'h4244fbab, 32'hc2127786, 32'h423b6410};
test_output[10760:10767] = '{32'h0, 32'h0, 32'h408f25a9, 32'h42ae1437, 32'h0, 32'h4244fbab, 32'h0, 32'h423b6410};
test_input[10768:10775] = '{32'h42304e31, 32'hc1abf405, 32'hc2b0e667, 32'h427ad45a, 32'h428b5e9c, 32'hc21eaf15, 32'hc20eb133, 32'hc088832d};
test_output[10768:10775] = '{32'h42304e31, 32'h0, 32'h0, 32'h427ad45a, 32'h428b5e9c, 32'h0, 32'h0, 32'h0};
test_input[10776:10783] = '{32'h4274b988, 32'h42a26614, 32'hc1940ee1, 32'h4151339f, 32'h41384823, 32'h41e825a3, 32'h42a0279c, 32'h4287cbe2};
test_output[10776:10783] = '{32'h4274b988, 32'h42a26614, 32'h0, 32'h4151339f, 32'h41384823, 32'h41e825a3, 32'h42a0279c, 32'h4287cbe2};
test_input[10784:10791] = '{32'h42baf1df, 32'hc2a463dc, 32'hc24a3584, 32'hc1d19263, 32'hc200e861, 32'h41deaaff, 32'hc1bf17f5, 32'hc2849523};
test_output[10784:10791] = '{32'h42baf1df, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41deaaff, 32'h0, 32'h0};
test_input[10792:10799] = '{32'h42817d7e, 32'hc28ac5e4, 32'h421ff79f, 32'h4110c3db, 32'h428e8c02, 32'hc22507ec, 32'hc223fdba, 32'hc2263fd0};
test_output[10792:10799] = '{32'h42817d7e, 32'h0, 32'h421ff79f, 32'h4110c3db, 32'h428e8c02, 32'h0, 32'h0, 32'h0};
test_input[10800:10807] = '{32'h4256edac, 32'hc240202b, 32'h42c2e05f, 32'hc29fb924, 32'h4215f5b0, 32'hc2949eb3, 32'hc2963efb, 32'hc1844007};
test_output[10800:10807] = '{32'h4256edac, 32'h0, 32'h42c2e05f, 32'h0, 32'h4215f5b0, 32'h0, 32'h0, 32'h0};
test_input[10808:10815] = '{32'h4191b234, 32'hc2a2a88d, 32'h428a9e18, 32'h42b4e33e, 32'h3f931b93, 32'hc2b89eaf, 32'hc209bf7b, 32'h42a942d2};
test_output[10808:10815] = '{32'h4191b234, 32'h0, 32'h428a9e18, 32'h42b4e33e, 32'h3f931b93, 32'h0, 32'h0, 32'h42a942d2};
test_input[10816:10823] = '{32'hc2969cf9, 32'h4131d3a7, 32'h424de397, 32'h42b74de3, 32'h4247c6b6, 32'hc1aad588, 32'h42885c61, 32'hc2b49b1e};
test_output[10816:10823] = '{32'h0, 32'h4131d3a7, 32'h424de397, 32'h42b74de3, 32'h4247c6b6, 32'h0, 32'h42885c61, 32'h0};
test_input[10824:10831] = '{32'h428d4a6c, 32'h426d4c1e, 32'hbf1c82ee, 32'h419d5b1a, 32'hc292099f, 32'hc22a2018, 32'hc1dfd9a4, 32'hc0e1c1ac};
test_output[10824:10831] = '{32'h428d4a6c, 32'h426d4c1e, 32'h0, 32'h419d5b1a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10832:10839] = '{32'hc24553c5, 32'hc0f2a498, 32'hc26e4a94, 32'h421c4dfa, 32'hc2a0c1f4, 32'hc29bbf34, 32'hc19a7f20, 32'h42b50397};
test_output[10832:10839] = '{32'h0, 32'h0, 32'h0, 32'h421c4dfa, 32'h0, 32'h0, 32'h0, 32'h42b50397};
test_input[10840:10847] = '{32'h42a51e45, 32'hc2475d02, 32'h422e5f1a, 32'h425f3435, 32'h42653a6e, 32'hc18b4c18, 32'h42a79c16, 32'h40d88982};
test_output[10840:10847] = '{32'h42a51e45, 32'h0, 32'h422e5f1a, 32'h425f3435, 32'h42653a6e, 32'h0, 32'h42a79c16, 32'h40d88982};
test_input[10848:10855] = '{32'h42b2aca0, 32'h42960d10, 32'hc13c2f9b, 32'h424231f1, 32'h42628972, 32'hc139521a, 32'hc2720b85, 32'h406425dc};
test_output[10848:10855] = '{32'h42b2aca0, 32'h42960d10, 32'h0, 32'h424231f1, 32'h42628972, 32'h0, 32'h0, 32'h406425dc};
test_input[10856:10863] = '{32'hc21d93df, 32'h424fe1c3, 32'hc18dfeab, 32'hc21cad26, 32'hc1821ef9, 32'hc1e01ebb, 32'hc0770ef1, 32'h42bffec8};
test_output[10856:10863] = '{32'h0, 32'h424fe1c3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bffec8};
test_input[10864:10871] = '{32'hc1ab1f72, 32'h4186afa6, 32'h413b54bf, 32'hc272c21f, 32'h42644f74, 32'hc19802c0, 32'hc27bb20d, 32'hc199f42a};
test_output[10864:10871] = '{32'h0, 32'h4186afa6, 32'h413b54bf, 32'h0, 32'h42644f74, 32'h0, 32'h0, 32'h0};
test_input[10872:10879] = '{32'hc1696dde, 32'hc0c37c89, 32'hc188414b, 32'hc26e6ed7, 32'h4253e583, 32'hc2563dc9, 32'hc276ec33, 32'h42c47704};
test_output[10872:10879] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4253e583, 32'h0, 32'h0, 32'h42c47704};
test_input[10880:10887] = '{32'hc1712a29, 32'h423f1ee2, 32'h422fd3b8, 32'h42af7986, 32'h42aeea40, 32'h416b5ff7, 32'h40a1c811, 32'h41cbcbfd};
test_output[10880:10887] = '{32'h0, 32'h423f1ee2, 32'h422fd3b8, 32'h42af7986, 32'h42aeea40, 32'h416b5ff7, 32'h40a1c811, 32'h41cbcbfd};
test_input[10888:10895] = '{32'h414b8b8f, 32'h423d087b, 32'hc1fccb58, 32'hc29052ca, 32'h409a982f, 32'h42b7d95a, 32'h42719d83, 32'hc284cd75};
test_output[10888:10895] = '{32'h414b8b8f, 32'h423d087b, 32'h0, 32'h0, 32'h409a982f, 32'h42b7d95a, 32'h42719d83, 32'h0};
test_input[10896:10903] = '{32'h42a3932c, 32'h417d6a70, 32'h42841e08, 32'hc1ce6284, 32'hc23d0805, 32'h41b24661, 32'hc24191be, 32'hc2826ca9};
test_output[10896:10903] = '{32'h42a3932c, 32'h417d6a70, 32'h42841e08, 32'h0, 32'h0, 32'h41b24661, 32'h0, 32'h0};
test_input[10904:10911] = '{32'h3f9c622b, 32'hc218b1f3, 32'h4261c897, 32'hc24e58df, 32'h428d6233, 32'h421afc3a, 32'h42140ee4, 32'hc1307e6a};
test_output[10904:10911] = '{32'h3f9c622b, 32'h0, 32'h4261c897, 32'h0, 32'h428d6233, 32'h421afc3a, 32'h42140ee4, 32'h0};
test_input[10912:10919] = '{32'hc216b309, 32'hc03be741, 32'h42bb5e9f, 32'hc235ca2e, 32'hc27fe28f, 32'h4281c3ba, 32'h4143ae12, 32'h42ba9847};
test_output[10912:10919] = '{32'h0, 32'h0, 32'h42bb5e9f, 32'h0, 32'h0, 32'h4281c3ba, 32'h4143ae12, 32'h42ba9847};
test_input[10920:10927] = '{32'h429414e1, 32'h42bed7f4, 32'h41ce6a6b, 32'h4213642a, 32'hc247407a, 32'h41c69d26, 32'hc20c35b9, 32'hc257418a};
test_output[10920:10927] = '{32'h429414e1, 32'h42bed7f4, 32'h41ce6a6b, 32'h4213642a, 32'h0, 32'h41c69d26, 32'h0, 32'h0};
test_input[10928:10935] = '{32'h42853829, 32'h41dfbb82, 32'hc19ace40, 32'hc11255f0, 32'hc175bc22, 32'hc28722c4, 32'h418332fa, 32'h42ab39e8};
test_output[10928:10935] = '{32'h42853829, 32'h41dfbb82, 32'h0, 32'h0, 32'h0, 32'h0, 32'h418332fa, 32'h42ab39e8};
test_input[10936:10943] = '{32'hc20da8a8, 32'h426d40c6, 32'hc21e6e55, 32'h426df23f, 32'hc20fdaf6, 32'h41fb2716, 32'hc23eb9c7, 32'hc269cb04};
test_output[10936:10943] = '{32'h0, 32'h426d40c6, 32'h0, 32'h426df23f, 32'h0, 32'h41fb2716, 32'h0, 32'h0};
test_input[10944:10951] = '{32'h421b04bf, 32'h412b7edb, 32'h42a65f5b, 32'h42c4cb9a, 32'hc1bd7d8c, 32'hc1b72abe, 32'h427b67fa, 32'h420f7072};
test_output[10944:10951] = '{32'h421b04bf, 32'h412b7edb, 32'h42a65f5b, 32'h42c4cb9a, 32'h0, 32'h0, 32'h427b67fa, 32'h420f7072};
test_input[10952:10959] = '{32'hc29c6c5c, 32'h42a16884, 32'hc23e13c4, 32'h42b56ee2, 32'h42c0bb22, 32'h41844c45, 32'h4251e58d, 32'h41d396e4};
test_output[10952:10959] = '{32'h0, 32'h42a16884, 32'h0, 32'h42b56ee2, 32'h42c0bb22, 32'h41844c45, 32'h4251e58d, 32'h41d396e4};
test_input[10960:10967] = '{32'hc292f482, 32'hc23ea5a9, 32'h40dc33ce, 32'hc2c524a8, 32'hc1a7b0f8, 32'h4138743c, 32'h41776689, 32'h42b1244d};
test_output[10960:10967] = '{32'h0, 32'h0, 32'h40dc33ce, 32'h0, 32'h0, 32'h4138743c, 32'h41776689, 32'h42b1244d};
test_input[10968:10975] = '{32'hc109c6c9, 32'hc2c04d22, 32'hc18439af, 32'hc2159fd8, 32'h429bd936, 32'hc180cfe5, 32'hc2aa3087, 32'h40de43b9};
test_output[10968:10975] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429bd936, 32'h0, 32'h0, 32'h40de43b9};
test_input[10976:10983] = '{32'hc2088126, 32'hc16b244e, 32'h4292d271, 32'h422ec8df, 32'hc2551289, 32'hc24b2f94, 32'hc284fcf0, 32'hc1d49402};
test_output[10976:10983] = '{32'h0, 32'h0, 32'h4292d271, 32'h422ec8df, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10984:10991] = '{32'hc0b8ef08, 32'hbfe44323, 32'h4136d90e, 32'h42c7c728, 32'hc26a1ee6, 32'h42143e30, 32'hc251b462, 32'hc25f18ac};
test_output[10984:10991] = '{32'h0, 32'h0, 32'h4136d90e, 32'h42c7c728, 32'h0, 32'h42143e30, 32'h0, 32'h0};
test_input[10992:10999] = '{32'hc28ee054, 32'hc29f2e13, 32'h42c5cecb, 32'h4002a609, 32'h40627e8b, 32'h425cf776, 32'h41e075c1, 32'h4082c309};
test_output[10992:10999] = '{32'h0, 32'h0, 32'h42c5cecb, 32'h4002a609, 32'h40627e8b, 32'h425cf776, 32'h41e075c1, 32'h4082c309};
test_input[11000:11007] = '{32'hc2c5a51e, 32'h40bbb858, 32'hc1feb970, 32'hc1e202d5, 32'h42c61bd8, 32'h3f914b01, 32'h428bac4e, 32'h426d9567};
test_output[11000:11007] = '{32'h0, 32'h40bbb858, 32'h0, 32'h0, 32'h42c61bd8, 32'h3f914b01, 32'h428bac4e, 32'h426d9567};
test_input[11008:11015] = '{32'hc1075cbd, 32'hc137c48f, 32'hc03fd818, 32'h424f93fd, 32'hc296e1b5, 32'h4258849a, 32'h42a1465a, 32'hc0ca8f03};
test_output[11008:11015] = '{32'h0, 32'h0, 32'h0, 32'h424f93fd, 32'h0, 32'h4258849a, 32'h42a1465a, 32'h0};
test_input[11016:11023] = '{32'h4283b527, 32'hc2ab9bf3, 32'hc0b122f1, 32'h42bb25af, 32'hc1b143eb, 32'h40dc186c, 32'hc2af4ed0, 32'h42bb9277};
test_output[11016:11023] = '{32'h4283b527, 32'h0, 32'h0, 32'h42bb25af, 32'h0, 32'h40dc186c, 32'h0, 32'h42bb9277};
test_input[11024:11031] = '{32'h428f6971, 32'h42952581, 32'hc2011b2f, 32'hc274a9f3, 32'hc22bad50, 32'hc28ce9bb, 32'hc2bdc9b2, 32'h42c5a21c};
test_output[11024:11031] = '{32'h428f6971, 32'h42952581, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c5a21c};
test_input[11032:11039] = '{32'hbf74c62c, 32'h41bad52e, 32'hc1daefc9, 32'hc28f52a6, 32'h424c0923, 32'hc212a760, 32'hc22bb978, 32'hc29bc37c};
test_output[11032:11039] = '{32'h0, 32'h41bad52e, 32'h0, 32'h0, 32'h424c0923, 32'h0, 32'h0, 32'h0};
test_input[11040:11047] = '{32'h41c8de12, 32'hc13992a7, 32'hc29d5f63, 32'hc2ba5bd8, 32'h426f7bf6, 32'h410994c9, 32'h425e5d4b, 32'hc29d2a4a};
test_output[11040:11047] = '{32'h41c8de12, 32'h0, 32'h0, 32'h0, 32'h426f7bf6, 32'h410994c9, 32'h425e5d4b, 32'h0};
test_input[11048:11055] = '{32'hc2bf36e3, 32'hc285971b, 32'h415bbbec, 32'hc0c9606b, 32'h42c7a186, 32'h41b84509, 32'h42768fa5, 32'h429cd8f9};
test_output[11048:11055] = '{32'h0, 32'h0, 32'h415bbbec, 32'h0, 32'h42c7a186, 32'h41b84509, 32'h42768fa5, 32'h429cd8f9};
test_input[11056:11063] = '{32'h428f0162, 32'h41fcb825, 32'hc1fbae5d, 32'h4299bedc, 32'hc2ab6345, 32'h42b8fe54, 32'hc273a1c5, 32'hc296fa59};
test_output[11056:11063] = '{32'h428f0162, 32'h41fcb825, 32'h0, 32'h4299bedc, 32'h0, 32'h42b8fe54, 32'h0, 32'h0};
test_input[11064:11071] = '{32'hc2a5def2, 32'h405c48bc, 32'h4186253a, 32'h42821c85, 32'h41aa4909, 32'hc1c7174f, 32'hc2997bd8, 32'h42187b2d};
test_output[11064:11071] = '{32'h0, 32'h405c48bc, 32'h4186253a, 32'h42821c85, 32'h41aa4909, 32'h0, 32'h0, 32'h42187b2d};
test_input[11072:11079] = '{32'hc2513baa, 32'h42c78948, 32'h42a24ff9, 32'hc2ab21f1, 32'h429477e0, 32'h420c17af, 32'h4271293d, 32'hc20fbee0};
test_output[11072:11079] = '{32'h0, 32'h42c78948, 32'h42a24ff9, 32'h0, 32'h429477e0, 32'h420c17af, 32'h4271293d, 32'h0};
test_input[11080:11087] = '{32'hc20e7845, 32'h427161f7, 32'h426bae08, 32'hc193846e, 32'h41d5dd7b, 32'h427e4143, 32'hc282fe82, 32'hc27dfd48};
test_output[11080:11087] = '{32'h0, 32'h427161f7, 32'h426bae08, 32'h0, 32'h41d5dd7b, 32'h427e4143, 32'h0, 32'h0};
test_input[11088:11095] = '{32'hc29e388a, 32'hc175083d, 32'hc24efcd0, 32'h41cfc94b, 32'h423b016c, 32'hc1d0d163, 32'hc23b682d, 32'h42bfd14c};
test_output[11088:11095] = '{32'h0, 32'h0, 32'h0, 32'h41cfc94b, 32'h423b016c, 32'h0, 32'h0, 32'h42bfd14c};
test_input[11096:11103] = '{32'h42b40589, 32'hc13fa413, 32'hc1de512c, 32'h421403bb, 32'hc224f51e, 32'h42579f3b, 32'hc216577d, 32'h418c38e6};
test_output[11096:11103] = '{32'h42b40589, 32'h0, 32'h0, 32'h421403bb, 32'h0, 32'h42579f3b, 32'h0, 32'h418c38e6};
test_input[11104:11111] = '{32'h428e8950, 32'hc2a5f640, 32'h42c7d61f, 32'hc2b48ee3, 32'h428d67b3, 32'hc282ccab, 32'h41ccc505, 32'h4194c307};
test_output[11104:11111] = '{32'h428e8950, 32'h0, 32'h42c7d61f, 32'h0, 32'h428d67b3, 32'h0, 32'h41ccc505, 32'h4194c307};
test_input[11112:11119] = '{32'h4230e5ab, 32'h40aac41d, 32'h42282122, 32'h41f699e1, 32'h42b656fc, 32'hc2a12472, 32'h423c0349, 32'h42ba2e4e};
test_output[11112:11119] = '{32'h4230e5ab, 32'h40aac41d, 32'h42282122, 32'h41f699e1, 32'h42b656fc, 32'h0, 32'h423c0349, 32'h42ba2e4e};
test_input[11120:11127] = '{32'h42859db3, 32'hc1ed160d, 32'h420e20a8, 32'hc290125e, 32'hc1cd8415, 32'h4173be14, 32'hc29e9cd4, 32'h42562c28};
test_output[11120:11127] = '{32'h42859db3, 32'h0, 32'h420e20a8, 32'h0, 32'h0, 32'h4173be14, 32'h0, 32'h42562c28};
test_input[11128:11135] = '{32'hc2316338, 32'h421783a1, 32'h40d048e4, 32'h42b78f89, 32'h3f524add, 32'hc2257eca, 32'hc28460b4, 32'hc1864df9};
test_output[11128:11135] = '{32'h0, 32'h421783a1, 32'h40d048e4, 32'h42b78f89, 32'h3f524add, 32'h0, 32'h0, 32'h0};
test_input[11136:11143] = '{32'hc2838870, 32'hc1788bc9, 32'h42138fbb, 32'h42bd05de, 32'h42914d12, 32'h4229291b, 32'h4112f217, 32'hc292e3da};
test_output[11136:11143] = '{32'h0, 32'h0, 32'h42138fbb, 32'h42bd05de, 32'h42914d12, 32'h4229291b, 32'h4112f217, 32'h0};
test_input[11144:11151] = '{32'hc24ca081, 32'hc18823a4, 32'hc13d1f02, 32'hc1ac8410, 32'h427b3e68, 32'h40ed47a8, 32'hc19469b5, 32'h41ec02e1};
test_output[11144:11151] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h427b3e68, 32'h40ed47a8, 32'h0, 32'h41ec02e1};
test_input[11152:11159] = '{32'hc21c56bc, 32'hc2a0be8d, 32'h421e60e2, 32'h421b9c61, 32'h4156d987, 32'h42a3be86, 32'h41c98a85, 32'h42aad695};
test_output[11152:11159] = '{32'h0, 32'h0, 32'h421e60e2, 32'h421b9c61, 32'h4156d987, 32'h42a3be86, 32'h41c98a85, 32'h42aad695};
test_input[11160:11167] = '{32'h419c84ae, 32'h41e1a092, 32'hc2092ba5, 32'hc160fdaf, 32'hc2168881, 32'h415df64d, 32'hc15aa893, 32'hc2c3fe18};
test_output[11160:11167] = '{32'h419c84ae, 32'h41e1a092, 32'h0, 32'h0, 32'h0, 32'h415df64d, 32'h0, 32'h0};
test_input[11168:11175] = '{32'hc17d165c, 32'h42ae53a7, 32'h429c51b5, 32'h42b03129, 32'hc291011b, 32'h41c652ad, 32'h42374c48, 32'h425c6d8c};
test_output[11168:11175] = '{32'h0, 32'h42ae53a7, 32'h429c51b5, 32'h42b03129, 32'h0, 32'h41c652ad, 32'h42374c48, 32'h425c6d8c};
test_input[11176:11183] = '{32'hc1ab1f7f, 32'hc2c2af37, 32'hc2afbdce, 32'hc1db1c62, 32'h4086f677, 32'hc1b93d19, 32'h4202c498, 32'hc29b65da};
test_output[11176:11183] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4086f677, 32'h0, 32'h4202c498, 32'h0};
test_input[11184:11191] = '{32'h41f04960, 32'hc0bca83c, 32'hc28d4574, 32'h4223cfae, 32'h4286d4f4, 32'h425fc5a8, 32'hc116f3e2, 32'h420d8e8b};
test_output[11184:11191] = '{32'h41f04960, 32'h0, 32'h0, 32'h4223cfae, 32'h4286d4f4, 32'h425fc5a8, 32'h0, 32'h420d8e8b};
test_input[11192:11199] = '{32'hc2ac1535, 32'h3f190dd9, 32'h40dec4dc, 32'hc2ba92ac, 32'h41216120, 32'h4224aa1f, 32'h41b32439, 32'h42c66d0f};
test_output[11192:11199] = '{32'h0, 32'h3f190dd9, 32'h40dec4dc, 32'h0, 32'h41216120, 32'h4224aa1f, 32'h41b32439, 32'h42c66d0f};
test_input[11200:11207] = '{32'h427628f4, 32'h42a4bb42, 32'hc1e8b6af, 32'h42a43c30, 32'h42a24b12, 32'hc1d5f514, 32'h42b22f6c, 32'h41199fe8};
test_output[11200:11207] = '{32'h427628f4, 32'h42a4bb42, 32'h0, 32'h42a43c30, 32'h42a24b12, 32'h0, 32'h42b22f6c, 32'h41199fe8};
test_input[11208:11215] = '{32'hc2ab827a, 32'hc2184f12, 32'hc299ca50, 32'hc2878abc, 32'h41969c6d, 32'h41eb1172, 32'h428dd519, 32'hc210bb8a};
test_output[11208:11215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41969c6d, 32'h41eb1172, 32'h428dd519, 32'h0};
test_input[11216:11223] = '{32'h427d9002, 32'h422947fe, 32'h42a9502f, 32'hc1d19e0a, 32'h42c4f1a0, 32'hc250168b, 32'h42821cf6, 32'hc2bb92d3};
test_output[11216:11223] = '{32'h427d9002, 32'h422947fe, 32'h42a9502f, 32'h0, 32'h42c4f1a0, 32'h0, 32'h42821cf6, 32'h0};
test_input[11224:11231] = '{32'hc18df8a3, 32'h41b0a297, 32'h4288eae8, 32'h423aa205, 32'h42267927, 32'h42118a5e, 32'hc206f847, 32'hc2ac0f57};
test_output[11224:11231] = '{32'h0, 32'h41b0a297, 32'h4288eae8, 32'h423aa205, 32'h42267927, 32'h42118a5e, 32'h0, 32'h0};
test_input[11232:11239] = '{32'h42af13ae, 32'hc2bad727, 32'hc2278a0a, 32'h4287f595, 32'h4213d86c, 32'hc29cfeb0, 32'h428eb04b, 32'h42b0ca69};
test_output[11232:11239] = '{32'h42af13ae, 32'h0, 32'h0, 32'h4287f595, 32'h4213d86c, 32'h0, 32'h428eb04b, 32'h42b0ca69};
test_input[11240:11247] = '{32'h423fb590, 32'h415bebae, 32'hc27ac307, 32'hc2c5911a, 32'h419f5099, 32'h41fdb638, 32'hc2133de1, 32'h4291a46a};
test_output[11240:11247] = '{32'h423fb590, 32'h415bebae, 32'h0, 32'h0, 32'h419f5099, 32'h41fdb638, 32'h0, 32'h4291a46a};
test_input[11248:11255] = '{32'h42636a66, 32'h42b8788f, 32'h4286fd08, 32'hc27b6cef, 32'hc28fe739, 32'hc2abbbf3, 32'h41ee33c2, 32'hc1f806cc};
test_output[11248:11255] = '{32'h42636a66, 32'h42b8788f, 32'h4286fd08, 32'h0, 32'h0, 32'h0, 32'h41ee33c2, 32'h0};
test_input[11256:11263] = '{32'hc2b24f3a, 32'hc28a261b, 32'h4208d09e, 32'h41194b58, 32'hc28b7b2e, 32'h4255c44d, 32'hc283c455, 32'hc294d653};
test_output[11256:11263] = '{32'h0, 32'h0, 32'h4208d09e, 32'h41194b58, 32'h0, 32'h4255c44d, 32'h0, 32'h0};
test_input[11264:11271] = '{32'hc2a07f4c, 32'h422d4408, 32'hc2701008, 32'h426a3371, 32'hc1de13fd, 32'hc2340eb9, 32'h429b4bcb, 32'h41c1eb0e};
test_output[11264:11271] = '{32'h0, 32'h422d4408, 32'h0, 32'h426a3371, 32'h0, 32'h0, 32'h429b4bcb, 32'h41c1eb0e};
test_input[11272:11279] = '{32'h42c05e48, 32'hc1b909c6, 32'hc2206a4c, 32'h4251d720, 32'h42807573, 32'hc28fb381, 32'h409868fe, 32'h421cf212};
test_output[11272:11279] = '{32'h42c05e48, 32'h0, 32'h0, 32'h4251d720, 32'h42807573, 32'h0, 32'h409868fe, 32'h421cf212};
test_input[11280:11287] = '{32'h42090027, 32'h42c00fee, 32'hc2a30f2f, 32'hc2a21c2d, 32'hc220c0d0, 32'hc29c811a, 32'h411ae09d, 32'hc25bc8d9};
test_output[11280:11287] = '{32'h42090027, 32'h42c00fee, 32'h0, 32'h0, 32'h0, 32'h0, 32'h411ae09d, 32'h0};
test_input[11288:11295] = '{32'h42c0b032, 32'hc2282a16, 32'h420fc775, 32'h42a84eab, 32'hc2b4c9bc, 32'h42af5544, 32'hc2ae263b, 32'hc1c757f0};
test_output[11288:11295] = '{32'h42c0b032, 32'h0, 32'h420fc775, 32'h42a84eab, 32'h0, 32'h42af5544, 32'h0, 32'h0};
test_input[11296:11303] = '{32'hc24d63ba, 32'h424acfc7, 32'hc2c13e97, 32'h428011c5, 32'hc25dda0c, 32'hc0a59642, 32'h40a91770, 32'hc25b8fa4};
test_output[11296:11303] = '{32'h0, 32'h424acfc7, 32'h0, 32'h428011c5, 32'h0, 32'h0, 32'h40a91770, 32'h0};
test_input[11304:11311] = '{32'hbf1400ff, 32'hc24a8325, 32'h40fbaa64, 32'h4240a490, 32'h41b0d89b, 32'hc0ce3ac0, 32'h42ac00e9, 32'hc216d558};
test_output[11304:11311] = '{32'h0, 32'h0, 32'h40fbaa64, 32'h4240a490, 32'h41b0d89b, 32'h0, 32'h42ac00e9, 32'h0};
test_input[11312:11319] = '{32'hc15292dd, 32'hc285f6b2, 32'h423cfb12, 32'h40cdf557, 32'h42aaeb27, 32'hc2147897, 32'hc29c6448, 32'hc29eaef8};
test_output[11312:11319] = '{32'h0, 32'h0, 32'h423cfb12, 32'h40cdf557, 32'h42aaeb27, 32'h0, 32'h0, 32'h0};
test_input[11320:11327] = '{32'h42765bce, 32'hc2c69c37, 32'h428b3ae0, 32'h405a5873, 32'hc22a527c, 32'h4134768e, 32'hc18bc7ce, 32'h426f1647};
test_output[11320:11327] = '{32'h42765bce, 32'h0, 32'h428b3ae0, 32'h405a5873, 32'h0, 32'h4134768e, 32'h0, 32'h426f1647};
test_input[11328:11335] = '{32'h429936de, 32'hc2561a53, 32'hc2ae1da3, 32'hc21018db, 32'hc2b808c2, 32'h4235fd71, 32'h423f2e8f, 32'h4256115a};
test_output[11328:11335] = '{32'h429936de, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4235fd71, 32'h423f2e8f, 32'h4256115a};
test_input[11336:11343] = '{32'hc268afb0, 32'hc2ab7cef, 32'h41638f84, 32'h41686beb, 32'hc27e31be, 32'hc2bbb844, 32'h41137fc0, 32'h3fd9275c};
test_output[11336:11343] = '{32'h0, 32'h0, 32'h41638f84, 32'h41686beb, 32'h0, 32'h0, 32'h41137fc0, 32'h3fd9275c};
test_input[11344:11351] = '{32'hc1853e03, 32'h40a7d4d8, 32'h42335c22, 32'h42afa71d, 32'h42849e2c, 32'hc2aa3b39, 32'h42bc415c, 32'h42a9b691};
test_output[11344:11351] = '{32'h0, 32'h40a7d4d8, 32'h42335c22, 32'h42afa71d, 32'h42849e2c, 32'h0, 32'h42bc415c, 32'h42a9b691};
test_input[11352:11359] = '{32'h42a20e2a, 32'hc155159f, 32'hc15820da, 32'h40f6dbf5, 32'hc12302e6, 32'hc239d45f, 32'h42a41c27, 32'hc2824a15};
test_output[11352:11359] = '{32'h42a20e2a, 32'h0, 32'h0, 32'h40f6dbf5, 32'h0, 32'h0, 32'h42a41c27, 32'h0};
test_input[11360:11367] = '{32'h42536122, 32'h429a93d3, 32'hc2735f2c, 32'hc290db31, 32'hc242b464, 32'hc25d0685, 32'h428ca57a, 32'h42973151};
test_output[11360:11367] = '{32'h42536122, 32'h429a93d3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428ca57a, 32'h42973151};
test_input[11368:11375] = '{32'hc20574ae, 32'h42bc5d15, 32'hc2227117, 32'hc2779924, 32'h41ee9dda, 32'hc19e1fa5, 32'hc272244c, 32'hc2469f2e};
test_output[11368:11375] = '{32'h0, 32'h42bc5d15, 32'h0, 32'h0, 32'h41ee9dda, 32'h0, 32'h0, 32'h0};
test_input[11376:11383] = '{32'hc28a9aa2, 32'hc1f29a83, 32'hc2a4da57, 32'h42c0dd27, 32'h422241b5, 32'hc2ad97f8, 32'hc173a3b8, 32'hc29744ca};
test_output[11376:11383] = '{32'h0, 32'h0, 32'h0, 32'h42c0dd27, 32'h422241b5, 32'h0, 32'h0, 32'h0};
test_input[11384:11391] = '{32'h424e7c24, 32'h41801352, 32'h42a83a54, 32'hc2164778, 32'h42b03d54, 32'h42a95f13, 32'hc1b21512, 32'hc2102c2f};
test_output[11384:11391] = '{32'h424e7c24, 32'h41801352, 32'h42a83a54, 32'h0, 32'h42b03d54, 32'h42a95f13, 32'h0, 32'h0};
test_input[11392:11399] = '{32'h4291027b, 32'h428d7e5e, 32'hc2218c99, 32'h4214ebf3, 32'hc26a53b2, 32'h428bd59f, 32'h4298a9d3, 32'h4265d007};
test_output[11392:11399] = '{32'h4291027b, 32'h428d7e5e, 32'h0, 32'h4214ebf3, 32'h0, 32'h428bd59f, 32'h4298a9d3, 32'h4265d007};
test_input[11400:11407] = '{32'hc14c972c, 32'hc1f73c28, 32'hc2580a20, 32'hc24fb478, 32'hc2b23df0, 32'h42b1ca7c, 32'h41121d58, 32'h4179f7e9};
test_output[11400:11407] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b1ca7c, 32'h41121d58, 32'h4179f7e9};
test_input[11408:11415] = '{32'h42a242ef, 32'hc28fd73a, 32'h41fcb184, 32'h3f9dc01c, 32'h41cd6eba, 32'hc20b4b62, 32'hc1a1c7d8, 32'hc22c479d};
test_output[11408:11415] = '{32'h42a242ef, 32'h0, 32'h41fcb184, 32'h3f9dc01c, 32'h41cd6eba, 32'h0, 32'h0, 32'h0};
test_input[11416:11423] = '{32'h413b5f51, 32'h4165a516, 32'h423ddad8, 32'hc219620a, 32'h418ccc4b, 32'h423c70c6, 32'hc25a24f6, 32'hc14c6db1};
test_output[11416:11423] = '{32'h413b5f51, 32'h4165a516, 32'h423ddad8, 32'h0, 32'h418ccc4b, 32'h423c70c6, 32'h0, 32'h0};
test_input[11424:11431] = '{32'hc2ba4140, 32'h428b6eb8, 32'hc246c5c5, 32'hc19b30e3, 32'h4229fbfe, 32'h42225cdf, 32'hc0fe847c, 32'h42c30268};
test_output[11424:11431] = '{32'h0, 32'h428b6eb8, 32'h0, 32'h0, 32'h4229fbfe, 32'h42225cdf, 32'h0, 32'h42c30268};
test_input[11432:11439] = '{32'hc29a7431, 32'hc27595ae, 32'h42523de4, 32'h42957c76, 32'hc2c36859, 32'hc2785d3e, 32'h42a365bc, 32'hc2b6a22b};
test_output[11432:11439] = '{32'h0, 32'h0, 32'h42523de4, 32'h42957c76, 32'h0, 32'h0, 32'h42a365bc, 32'h0};
test_input[11440:11447] = '{32'h422ca479, 32'hc2a60d06, 32'hc287b850, 32'hc2909e2a, 32'h421cead2, 32'hc25a0bd4, 32'h42c4156f, 32'h42835e1c};
test_output[11440:11447] = '{32'h422ca479, 32'h0, 32'h0, 32'h0, 32'h421cead2, 32'h0, 32'h42c4156f, 32'h42835e1c};
test_input[11448:11455] = '{32'hc1df3662, 32'h42997d5f, 32'hc232a35b, 32'h428dcbe7, 32'h41d364d1, 32'hc2359639, 32'hc2008ea5, 32'hc2b12e4d};
test_output[11448:11455] = '{32'h0, 32'h42997d5f, 32'h0, 32'h428dcbe7, 32'h41d364d1, 32'h0, 32'h0, 32'h0};
test_input[11456:11463] = '{32'hc1b012ae, 32'h42b1d744, 32'h42908fe8, 32'hc0bc37d6, 32'h42b685b9, 32'hc2a8b890, 32'h42bc54e6, 32'hc19d7bf3};
test_output[11456:11463] = '{32'h0, 32'h42b1d744, 32'h42908fe8, 32'h0, 32'h42b685b9, 32'h0, 32'h42bc54e6, 32'h0};
test_input[11464:11471] = '{32'hc2b9595e, 32'hc22ee13d, 32'hc29be781, 32'h422a6615, 32'hc2b0a3c8, 32'hbfa49f85, 32'hc22fb3d9, 32'hc21a226c};
test_output[11464:11471] = '{32'h0, 32'h0, 32'h0, 32'h422a6615, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11472:11479] = '{32'h426af488, 32'hc1aa5907, 32'h413ba5e1, 32'hc20489d8, 32'h4014ede6, 32'h42b31419, 32'h4109938a, 32'hc1463889};
test_output[11472:11479] = '{32'h426af488, 32'h0, 32'h413ba5e1, 32'h0, 32'h4014ede6, 32'h42b31419, 32'h4109938a, 32'h0};
test_input[11480:11487] = '{32'h3ef644cd, 32'h4176ef8e, 32'hc2b28c96, 32'hc2b9d0bb, 32'h4278f66c, 32'hc2c0ba26, 32'hbf5095df, 32'hc254fcb3};
test_output[11480:11487] = '{32'h3ef644cd, 32'h4176ef8e, 32'h0, 32'h0, 32'h4278f66c, 32'h0, 32'h0, 32'h0};
test_input[11488:11495] = '{32'hc2ac081d, 32'h429346bd, 32'hc22c0647, 32'h4238de11, 32'h4215d76e, 32'h40b4ee52, 32'hc2c2c5ad, 32'hc14c14ff};
test_output[11488:11495] = '{32'h0, 32'h429346bd, 32'h0, 32'h4238de11, 32'h4215d76e, 32'h40b4ee52, 32'h0, 32'h0};
test_input[11496:11503] = '{32'hc2c0cbfc, 32'h4197dd4a, 32'h419835cb, 32'hc278a4e5, 32'hc1e26865, 32'hc191547a, 32'hc1ad7485, 32'h4245f95c};
test_output[11496:11503] = '{32'h0, 32'h4197dd4a, 32'h419835cb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4245f95c};
test_input[11504:11511] = '{32'h42197068, 32'hc2b8f686, 32'h42a3fca9, 32'hc2bad684, 32'h40cec1f2, 32'h425d28c4, 32'hc1e73ccc, 32'hc1afeadf};
test_output[11504:11511] = '{32'h42197068, 32'h0, 32'h42a3fca9, 32'h0, 32'h40cec1f2, 32'h425d28c4, 32'h0, 32'h0};
test_input[11512:11519] = '{32'hc1f39e47, 32'hc1dccd57, 32'hc2b579d2, 32'h409a0e3a, 32'hc21f2601, 32'h424a5234, 32'h4183b3b1, 32'h428d9488};
test_output[11512:11519] = '{32'h0, 32'h0, 32'h0, 32'h409a0e3a, 32'h0, 32'h424a5234, 32'h4183b3b1, 32'h428d9488};
test_input[11520:11527] = '{32'hc268fea0, 32'hc2517fac, 32'hc1860c1b, 32'h41c9f503, 32'hc25e6393, 32'hc1986b15, 32'h423e16e6, 32'h4292e837};
test_output[11520:11527] = '{32'h0, 32'h0, 32'h0, 32'h41c9f503, 32'h0, 32'h0, 32'h423e16e6, 32'h4292e837};
test_input[11528:11535] = '{32'hc25023b9, 32'hc1b06ba7, 32'h427e993a, 32'h425a8e87, 32'hc20ef9ab, 32'hc20217d4, 32'h428b909d, 32'h4132478d};
test_output[11528:11535] = '{32'h0, 32'h0, 32'h427e993a, 32'h425a8e87, 32'h0, 32'h0, 32'h428b909d, 32'h4132478d};
test_input[11536:11543] = '{32'hc25864d6, 32'hc20e458a, 32'h41ccd9fa, 32'hc1b15187, 32'h424ef28d, 32'h4268a3e7, 32'hc141e0ed, 32'hc00f4f57};
test_output[11536:11543] = '{32'h0, 32'h0, 32'h41ccd9fa, 32'h0, 32'h424ef28d, 32'h4268a3e7, 32'h0, 32'h0};
test_input[11544:11551] = '{32'hc1f0c15f, 32'h4286d73d, 32'h406d627c, 32'hc2c60474, 32'h42708fe2, 32'h3f3953f4, 32'h42c6ef99, 32'hc22bfa58};
test_output[11544:11551] = '{32'h0, 32'h4286d73d, 32'h406d627c, 32'h0, 32'h42708fe2, 32'h3f3953f4, 32'h42c6ef99, 32'h0};
test_input[11552:11559] = '{32'hc23aef3b, 32'hc1f8924c, 32'hc27e11af, 32'hc2b94db8, 32'hc21bb515, 32'h42bd5336, 32'h420fc051, 32'hc2299a68};
test_output[11552:11559] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bd5336, 32'h420fc051, 32'h0};
test_input[11560:11567] = '{32'hc172db27, 32'hc1d795d4, 32'hc2c2d69b, 32'hc156576d, 32'h42af699f, 32'h4091e262, 32'h40dce6aa, 32'h42c2b173};
test_output[11560:11567] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42af699f, 32'h4091e262, 32'h40dce6aa, 32'h42c2b173};
test_input[11568:11575] = '{32'hc2c2be56, 32'h41b69b00, 32'h41bd3af4, 32'hc2873619, 32'h42af7432, 32'hc2887954, 32'hc2b02a0f, 32'hc0cdf9c0};
test_output[11568:11575] = '{32'h0, 32'h41b69b00, 32'h41bd3af4, 32'h0, 32'h42af7432, 32'h0, 32'h0, 32'h0};
test_input[11576:11583] = '{32'hc1512a1b, 32'hc126baa9, 32'h4261f5ab, 32'h42bc6134, 32'h42860dac, 32'h414bbab2, 32'hc26124a5, 32'h422036fe};
test_output[11576:11583] = '{32'h0, 32'h0, 32'h4261f5ab, 32'h42bc6134, 32'h42860dac, 32'h414bbab2, 32'h0, 32'h422036fe};
test_input[11584:11591] = '{32'hc2414430, 32'h4270c39c, 32'h41f997f0, 32'h424c833c, 32'hc0fb9293, 32'h42bd160f, 32'h41eec052, 32'hc16ca702};
test_output[11584:11591] = '{32'h0, 32'h4270c39c, 32'h41f997f0, 32'h424c833c, 32'h0, 32'h42bd160f, 32'h41eec052, 32'h0};
test_input[11592:11599] = '{32'h428cdb59, 32'h41cdb54a, 32'h422a5e71, 32'hc28c221d, 32'h419da4e4, 32'hc1d4e888, 32'h42afd10e, 32'hc2879145};
test_output[11592:11599] = '{32'h428cdb59, 32'h41cdb54a, 32'h422a5e71, 32'h0, 32'h419da4e4, 32'h0, 32'h42afd10e, 32'h0};
test_input[11600:11607] = '{32'hc18e475d, 32'hc10441aa, 32'hc2144a88, 32'hc1d69c2b, 32'hc1190abd, 32'hc27c8526, 32'h42441bb0, 32'hc2add4d4};
test_output[11600:11607] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42441bb0, 32'h0};
test_input[11608:11615] = '{32'hc2a17954, 32'hc292bb64, 32'h42bf157f, 32'hc1a098b3, 32'hc2bd6b3e, 32'hc288cc77, 32'h42353686, 32'h41e0f119};
test_output[11608:11615] = '{32'h0, 32'h0, 32'h42bf157f, 32'h0, 32'h0, 32'h0, 32'h42353686, 32'h41e0f119};
test_input[11616:11623] = '{32'h427d826a, 32'h41beea4b, 32'hc2a0b5b8, 32'hc2c4f71c, 32'hc2b8253d, 32'hc28612df, 32'hc25fb95b, 32'h4283755b};
test_output[11616:11623] = '{32'h427d826a, 32'h41beea4b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4283755b};
test_input[11624:11631] = '{32'hc2517014, 32'hc258ace6, 32'hc0075195, 32'hc280001f, 32'hc2673b69, 32'h42831dec, 32'hc2c64bc9, 32'h421cc989};
test_output[11624:11631] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42831dec, 32'h0, 32'h421cc989};
test_input[11632:11639] = '{32'h41808637, 32'h413b874f, 32'h4216a6d8, 32'hc1c9856c, 32'h41b091aa, 32'hc2843a10, 32'h42372720, 32'hc241da49};
test_output[11632:11639] = '{32'h41808637, 32'h413b874f, 32'h4216a6d8, 32'h0, 32'h41b091aa, 32'h0, 32'h42372720, 32'h0};
test_input[11640:11647] = '{32'hc22a064b, 32'hc2a87f3e, 32'hc28b5820, 32'h42bcbacc, 32'h42b6393a, 32'h41a769d4, 32'h414b42e6, 32'h42c0e397};
test_output[11640:11647] = '{32'h0, 32'h0, 32'h0, 32'h42bcbacc, 32'h42b6393a, 32'h41a769d4, 32'h414b42e6, 32'h42c0e397};
test_input[11648:11655] = '{32'hc1aa7ad0, 32'hc1b77f88, 32'h428a9efa, 32'h41e0ec16, 32'h422ce983, 32'hc215d0cd, 32'hc29003a9, 32'h41babfcb};
test_output[11648:11655] = '{32'h0, 32'h0, 32'h428a9efa, 32'h41e0ec16, 32'h422ce983, 32'h0, 32'h0, 32'h41babfcb};
test_input[11656:11663] = '{32'hc24106a1, 32'hc2c04470, 32'hc25bff32, 32'h425db5f6, 32'h42a5ba58, 32'hc23facc6, 32'hc240a741, 32'h42c0b277};
test_output[11656:11663] = '{32'h0, 32'h0, 32'h0, 32'h425db5f6, 32'h42a5ba58, 32'h0, 32'h0, 32'h42c0b277};
test_input[11664:11671] = '{32'hc2a70e4f, 32'hc219af3c, 32'hc2c438f0, 32'hc2047073, 32'h42b42f51, 32'hc1d08569, 32'hc24ca32d, 32'hc2a1a384};
test_output[11664:11671] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42b42f51, 32'h0, 32'h0, 32'h0};
test_input[11672:11679] = '{32'h4132b293, 32'h42bed0d7, 32'h421b997b, 32'hbe977e6f, 32'h42bfaf13, 32'h423557bf, 32'hc1c03345, 32'hc2b31719};
test_output[11672:11679] = '{32'h4132b293, 32'h42bed0d7, 32'h421b997b, 32'h0, 32'h42bfaf13, 32'h423557bf, 32'h0, 32'h0};
test_input[11680:11687] = '{32'hc29a791e, 32'hc22c790a, 32'h42abbbe2, 32'hc217ea1c, 32'hc2a0c7a9, 32'h42a90d38, 32'h42b93387, 32'hc29afbe2};
test_output[11680:11687] = '{32'h0, 32'h0, 32'h42abbbe2, 32'h0, 32'h0, 32'h42a90d38, 32'h42b93387, 32'h0};
test_input[11688:11695] = '{32'h42a7e682, 32'h423877e8, 32'hc2b8a8b5, 32'hc292246f, 32'hc29ce712, 32'h42c01cf5, 32'hc229dcbd, 32'h42030a5a};
test_output[11688:11695] = '{32'h42a7e682, 32'h423877e8, 32'h0, 32'h0, 32'h0, 32'h42c01cf5, 32'h0, 32'h42030a5a};
test_input[11696:11703] = '{32'hc1c538b3, 32'h42a5e360, 32'hc2b24aa7, 32'h42551620, 32'hc11882be, 32'h4216a48c, 32'h42738a7b, 32'hc2951dc2};
test_output[11696:11703] = '{32'h0, 32'h42a5e360, 32'h0, 32'h42551620, 32'h0, 32'h4216a48c, 32'h42738a7b, 32'h0};
test_input[11704:11711] = '{32'h42a80dd1, 32'hc13ec44c, 32'h41c6ace1, 32'h429d13ae, 32'h428bc7c7, 32'hc27a441e, 32'hc1e6f14b, 32'h420117db};
test_output[11704:11711] = '{32'h42a80dd1, 32'h0, 32'h41c6ace1, 32'h429d13ae, 32'h428bc7c7, 32'h0, 32'h0, 32'h420117db};
test_input[11712:11719] = '{32'h4217c2de, 32'h41a84376, 32'hc17cad22, 32'h41a4ed98, 32'h41f3b94e, 32'h42c75ce1, 32'h4281f610, 32'h42a3bb21};
test_output[11712:11719] = '{32'h4217c2de, 32'h41a84376, 32'h0, 32'h41a4ed98, 32'h41f3b94e, 32'h42c75ce1, 32'h4281f610, 32'h42a3bb21};
test_input[11720:11727] = '{32'h416c8850, 32'h42bd4a00, 32'h41c15c2e, 32'h4053217a, 32'hc248631b, 32'h424a7c47, 32'hbfc8b817, 32'hc17b8856};
test_output[11720:11727] = '{32'h416c8850, 32'h42bd4a00, 32'h41c15c2e, 32'h4053217a, 32'h0, 32'h424a7c47, 32'h0, 32'h0};
test_input[11728:11735] = '{32'hc1de08e6, 32'h42a5993c, 32'hc21085d3, 32'h4230a254, 32'hc28551ff, 32'h421a4846, 32'h42968f85, 32'h41957ae4};
test_output[11728:11735] = '{32'h0, 32'h42a5993c, 32'h0, 32'h4230a254, 32'h0, 32'h421a4846, 32'h42968f85, 32'h41957ae4};
test_input[11736:11743] = '{32'hc1e6db72, 32'h424ff5f5, 32'h42056b43, 32'hc0751d51, 32'hc2263663, 32'h41d6b2fa, 32'hc26757d9, 32'hc2187ab7};
test_output[11736:11743] = '{32'h0, 32'h424ff5f5, 32'h42056b43, 32'h0, 32'h0, 32'h41d6b2fa, 32'h0, 32'h0};
test_input[11744:11751] = '{32'h415f3b6c, 32'h4288942e, 32'hc1069f13, 32'h42623e7f, 32'hc0310088, 32'hc1104948, 32'h4232b288, 32'hc1a0aa1b};
test_output[11744:11751] = '{32'h415f3b6c, 32'h4288942e, 32'h0, 32'h42623e7f, 32'h0, 32'h0, 32'h4232b288, 32'h0};
test_input[11752:11759] = '{32'hc1190b2d, 32'h425f0dd0, 32'h42911caf, 32'h4160bea5, 32'hc237ea46, 32'h40cd7b61, 32'h42b51760, 32'hc29f6898};
test_output[11752:11759] = '{32'h0, 32'h425f0dd0, 32'h42911caf, 32'h4160bea5, 32'h0, 32'h40cd7b61, 32'h42b51760, 32'h0};
test_input[11760:11767] = '{32'hc0b8fe05, 32'hc150b816, 32'hc24715fa, 32'h41b3db97, 32'hc26e1ac3, 32'hc22a6729, 32'hc2b4d711, 32'hc254ae4b};
test_output[11760:11767] = '{32'h0, 32'h0, 32'h0, 32'h41b3db97, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11768:11775] = '{32'hc2bdab83, 32'h42b5e030, 32'hc10b0419, 32'h41fd1139, 32'hc24cd3cd, 32'hc18531e8, 32'h427c4771, 32'h419e4312};
test_output[11768:11775] = '{32'h0, 32'h42b5e030, 32'h0, 32'h41fd1139, 32'h0, 32'h0, 32'h427c4771, 32'h419e4312};
test_input[11776:11783] = '{32'hc2ab135a, 32'h429a01a5, 32'h41748874, 32'hc2aaa132, 32'hc23ec0da, 32'h4155cc1e, 32'hc2241cf0, 32'h412bfe88};
test_output[11776:11783] = '{32'h0, 32'h429a01a5, 32'h41748874, 32'h0, 32'h0, 32'h4155cc1e, 32'h0, 32'h412bfe88};
test_input[11784:11791] = '{32'hc2c2d851, 32'h42bc5849, 32'hc29622b8, 32'h41c33216, 32'h42c25bb8, 32'h42c3bbcb, 32'h417931f4, 32'h429e87d1};
test_output[11784:11791] = '{32'h0, 32'h42bc5849, 32'h0, 32'h41c33216, 32'h42c25bb8, 32'h42c3bbcb, 32'h417931f4, 32'h429e87d1};
test_input[11792:11799] = '{32'h4080963c, 32'h42b2a16c, 32'hc241ea49, 32'hc0179dd5, 32'h41d585a0, 32'hc0ddb9ab, 32'hc1f599db, 32'hc0d2aa64};
test_output[11792:11799] = '{32'h4080963c, 32'h42b2a16c, 32'h0, 32'h0, 32'h41d585a0, 32'h0, 32'h0, 32'h0};
test_input[11800:11807] = '{32'h42838dea, 32'hc2153ae3, 32'hc1562deb, 32'hc24c4582, 32'hc1a5e72b, 32'hc1aabcac, 32'h4282f44c, 32'hc200b18e};
test_output[11800:11807] = '{32'h42838dea, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4282f44c, 32'h0};
test_input[11808:11815] = '{32'h4288a9d8, 32'hc1c3c665, 32'hc2648457, 32'hc2a8b44a, 32'hc1c43079, 32'hc0953393, 32'h413fc583, 32'h41ecbe10};
test_output[11808:11815] = '{32'h4288a9d8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h413fc583, 32'h41ecbe10};
test_input[11816:11823] = '{32'h42a0dfc2, 32'hc088a1ce, 32'h4207860c, 32'h42a1dc32, 32'hc2a9035b, 32'hc1930b7d, 32'h42376a5e, 32'h422f348c};
test_output[11816:11823] = '{32'h42a0dfc2, 32'h0, 32'h4207860c, 32'h42a1dc32, 32'h0, 32'h0, 32'h42376a5e, 32'h422f348c};
test_input[11824:11831] = '{32'hc2b51a9d, 32'h42544816, 32'hc2a293f2, 32'h42003123, 32'h4251e77c, 32'hc1d90e79, 32'h4298e8da, 32'h4297cb93};
test_output[11824:11831] = '{32'h0, 32'h42544816, 32'h0, 32'h42003123, 32'h4251e77c, 32'h0, 32'h4298e8da, 32'h4297cb93};
test_input[11832:11839] = '{32'h42a4d492, 32'h42b33fe6, 32'h42c08f2d, 32'h42a48cec, 32'hc2814c2b, 32'hc1d43853, 32'hc21672d2, 32'hc1e60fb6};
test_output[11832:11839] = '{32'h42a4d492, 32'h42b33fe6, 32'h42c08f2d, 32'h42a48cec, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11840:11847] = '{32'hc22144df, 32'hc13bf695, 32'h4150de27, 32'h400c064e, 32'hc28a641f, 32'h428d0867, 32'hc228b69a, 32'hc1043acd};
test_output[11840:11847] = '{32'h0, 32'h0, 32'h4150de27, 32'h400c064e, 32'h0, 32'h428d0867, 32'h0, 32'h0};
test_input[11848:11855] = '{32'h42a7853f, 32'h42ac1727, 32'h428e0702, 32'h425b7605, 32'h42a5880a, 32'hc136fef7, 32'hc28f57ab, 32'h4293778c};
test_output[11848:11855] = '{32'h42a7853f, 32'h42ac1727, 32'h428e0702, 32'h425b7605, 32'h42a5880a, 32'h0, 32'h0, 32'h4293778c};
test_input[11856:11863] = '{32'h428a2fb7, 32'hc270ccc7, 32'hc2070c4d, 32'h401ef368, 32'hc29a1604, 32'hc2a2142a, 32'h42904dd9, 32'hc1e39d8e};
test_output[11856:11863] = '{32'h428a2fb7, 32'h0, 32'h0, 32'h401ef368, 32'h0, 32'h0, 32'h42904dd9, 32'h0};
test_input[11864:11871] = '{32'h41f7cecb, 32'h410847be, 32'hc22fd973, 32'h429c43a6, 32'h42386bce, 32'hc130b2e8, 32'h42347a51, 32'h3f5d6824};
test_output[11864:11871] = '{32'h41f7cecb, 32'h410847be, 32'h0, 32'h429c43a6, 32'h42386bce, 32'h0, 32'h42347a51, 32'h3f5d6824};
test_input[11872:11879] = '{32'hc16ae8f0, 32'hc24d8813, 32'h42680d26, 32'h4154b1c8, 32'h421fd6ff, 32'hc2618f3c, 32'h41c39905, 32'h42489e22};
test_output[11872:11879] = '{32'h0, 32'h0, 32'h42680d26, 32'h4154b1c8, 32'h421fd6ff, 32'h0, 32'h41c39905, 32'h42489e22};
test_input[11880:11887] = '{32'h41164f24, 32'hc1ca9000, 32'hc1bbd9fa, 32'h4299863a, 32'hc26a2dfa, 32'hc2600f07, 32'hc2bc0bca, 32'hc136c757};
test_output[11880:11887] = '{32'h41164f24, 32'h0, 32'h0, 32'h4299863a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11888:11895] = '{32'hc264fe9a, 32'h4239111c, 32'hc21f04a1, 32'h429d91e9, 32'h42391812, 32'hc1a105a4, 32'h42925a7f, 32'h4240c7b9};
test_output[11888:11895] = '{32'h0, 32'h4239111c, 32'h0, 32'h429d91e9, 32'h42391812, 32'h0, 32'h42925a7f, 32'h4240c7b9};
test_input[11896:11903] = '{32'h42b8a8da, 32'hc261e750, 32'h42a8c303, 32'hc24c49bd, 32'hc1edf6b6, 32'h42c724e4, 32'h4218fc3c, 32'h42a5bf24};
test_output[11896:11903] = '{32'h42b8a8da, 32'h0, 32'h42a8c303, 32'h0, 32'h0, 32'h42c724e4, 32'h4218fc3c, 32'h42a5bf24};
test_input[11904:11911] = '{32'h4193d447, 32'hc23c701a, 32'h42817cff, 32'h418a03e1, 32'hc22aac12, 32'h407fd5b4, 32'h42b51aed, 32'h428befc4};
test_output[11904:11911] = '{32'h4193d447, 32'h0, 32'h42817cff, 32'h418a03e1, 32'h0, 32'h407fd5b4, 32'h42b51aed, 32'h428befc4};
test_input[11912:11919] = '{32'h410f7c2a, 32'h4263db3c, 32'h4236a1ee, 32'hc20dba80, 32'hc2292f37, 32'h418e71db, 32'hc21a0c4c, 32'hc1246323};
test_output[11912:11919] = '{32'h410f7c2a, 32'h4263db3c, 32'h4236a1ee, 32'h0, 32'h0, 32'h418e71db, 32'h0, 32'h0};
test_input[11920:11927] = '{32'h4286d625, 32'hc29c3b2c, 32'hc094933b, 32'h41df8380, 32'hc24a233c, 32'h42342d2b, 32'h428833ec, 32'h417514ee};
test_output[11920:11927] = '{32'h4286d625, 32'h0, 32'h0, 32'h41df8380, 32'h0, 32'h42342d2b, 32'h428833ec, 32'h417514ee};
test_input[11928:11935] = '{32'h403bba17, 32'hc246d4e8, 32'h41dc9f30, 32'hc28aaccd, 32'h4275b165, 32'h3e5f1b1e, 32'hc07c0629, 32'h427e478a};
test_output[11928:11935] = '{32'h403bba17, 32'h0, 32'h41dc9f30, 32'h0, 32'h4275b165, 32'h3e5f1b1e, 32'h0, 32'h427e478a};
test_input[11936:11943] = '{32'hc2b6e7e3, 32'h42abd30c, 32'hc2928ae8, 32'h42a3d5f6, 32'hc2934415, 32'h426b2bdd, 32'hc20e4bf8, 32'hc27491b4};
test_output[11936:11943] = '{32'h0, 32'h42abd30c, 32'h0, 32'h42a3d5f6, 32'h0, 32'h426b2bdd, 32'h0, 32'h0};
test_input[11944:11951] = '{32'hc0d76cad, 32'h425160d3, 32'hc24244dd, 32'hc0fbd95e, 32'hc28f94e7, 32'h4274f9bd, 32'h42a9cf12, 32'h41cc1612};
test_output[11944:11951] = '{32'h0, 32'h425160d3, 32'h0, 32'h0, 32'h0, 32'h4274f9bd, 32'h42a9cf12, 32'h41cc1612};
test_input[11952:11959] = '{32'h4260e3d3, 32'h42adc586, 32'h41d82076, 32'hc01e242f, 32'h42a9ce7d, 32'hc2c67d3c, 32'hbf94453d, 32'hc2151e14};
test_output[11952:11959] = '{32'h4260e3d3, 32'h42adc586, 32'h41d82076, 32'h0, 32'h42a9ce7d, 32'h0, 32'h0, 32'h0};
test_input[11960:11967] = '{32'hc2756208, 32'h42c26abc, 32'hc233f445, 32'h428845e6, 32'hc280b7c1, 32'h421690be, 32'hbc26fd42, 32'hc284e858};
test_output[11960:11967] = '{32'h0, 32'h42c26abc, 32'h0, 32'h428845e6, 32'h0, 32'h421690be, 32'h0, 32'h0};
test_input[11968:11975] = '{32'h41d82c1f, 32'h4275b197, 32'hc280a916, 32'h426ae7f4, 32'hc295983a, 32'h428924e3, 32'hc28bc2b0, 32'h41cee294};
test_output[11968:11975] = '{32'h41d82c1f, 32'h4275b197, 32'h0, 32'h426ae7f4, 32'h0, 32'h428924e3, 32'h0, 32'h41cee294};
test_input[11976:11983] = '{32'hc146688b, 32'h42b4b375, 32'h42408116, 32'hc25c9c2f, 32'h42892851, 32'hc2a21250, 32'hc2a3a0c4, 32'h413c5bad};
test_output[11976:11983] = '{32'h0, 32'h42b4b375, 32'h42408116, 32'h0, 32'h42892851, 32'h0, 32'h0, 32'h413c5bad};
test_input[11984:11991] = '{32'h42a53d3d, 32'h42bf4b57, 32'hc29dc7cc, 32'hc29daf09, 32'h41a1b791, 32'h429d18b9, 32'h41615603, 32'hc2b6e034};
test_output[11984:11991] = '{32'h42a53d3d, 32'h42bf4b57, 32'h0, 32'h0, 32'h41a1b791, 32'h429d18b9, 32'h41615603, 32'h0};
test_input[11992:11999] = '{32'hc1e98ae8, 32'h428a1769, 32'hc26c6b39, 32'h41f49d6e, 32'h428d6cb5, 32'h42bc8f14, 32'hc1321aec, 32'h41184dac};
test_output[11992:11999] = '{32'h0, 32'h428a1769, 32'h0, 32'h41f49d6e, 32'h428d6cb5, 32'h42bc8f14, 32'h0, 32'h41184dac};
test_input[12000:12007] = '{32'hc02a60fe, 32'hc193845f, 32'hc1a1eee2, 32'hc28aed0a, 32'hc24fb532, 32'h428ad13c, 32'h429b1b43, 32'hc20931f0};
test_output[12000:12007] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428ad13c, 32'h429b1b43, 32'h0};
test_input[12008:12015] = '{32'hc195296b, 32'hc29bf5a1, 32'hc2b5be86, 32'h42a747b1, 32'h428fed04, 32'h41fd9d82, 32'h421c66f3, 32'hc20289ce};
test_output[12008:12015] = '{32'h0, 32'h0, 32'h0, 32'h42a747b1, 32'h428fed04, 32'h41fd9d82, 32'h421c66f3, 32'h0};
test_input[12016:12023] = '{32'hc195f005, 32'hc2aec8ec, 32'h422cd1a5, 32'h4270a346, 32'h42284176, 32'hc20913ba, 32'hc1f4e757, 32'hc2964c60};
test_output[12016:12023] = '{32'h0, 32'h0, 32'h422cd1a5, 32'h4270a346, 32'h42284176, 32'h0, 32'h0, 32'h0};
test_input[12024:12031] = '{32'hc08394a8, 32'h429d5646, 32'hc19f362d, 32'hc060cd82, 32'h41ef54b1, 32'h42c471aa, 32'h42830ad6, 32'h401e2b20};
test_output[12024:12031] = '{32'h0, 32'h429d5646, 32'h0, 32'h0, 32'h41ef54b1, 32'h42c471aa, 32'h42830ad6, 32'h401e2b20};
test_input[12032:12039] = '{32'h42a3b8da, 32'hc22f7975, 32'hc24919ab, 32'h42778b4d, 32'hc151cdc1, 32'hc2c50404, 32'h421d7d03, 32'h41fc7bb0};
test_output[12032:12039] = '{32'h42a3b8da, 32'h0, 32'h0, 32'h42778b4d, 32'h0, 32'h0, 32'h421d7d03, 32'h41fc7bb0};
test_input[12040:12047] = '{32'h40fad754, 32'h42a2b4da, 32'hc23011a0, 32'h415ee80a, 32'h4178b623, 32'h41facf4f, 32'hc206a09e, 32'hc29440a4};
test_output[12040:12047] = '{32'h40fad754, 32'h42a2b4da, 32'h0, 32'h415ee80a, 32'h4178b623, 32'h41facf4f, 32'h0, 32'h0};
test_input[12048:12055] = '{32'hc28e214d, 32'hc2a7820c, 32'h4133b3ce, 32'hc2b7e62e, 32'h4262a0d2, 32'h42889334, 32'h426b655c, 32'h42453eda};
test_output[12048:12055] = '{32'h0, 32'h0, 32'h4133b3ce, 32'h0, 32'h4262a0d2, 32'h42889334, 32'h426b655c, 32'h42453eda};
test_input[12056:12063] = '{32'h415c8fbf, 32'h41a38dc1, 32'hc2c3ce9c, 32'hc0da319f, 32'hc197fd75, 32'hc27dc88c, 32'hc20690fb, 32'hc1f85cda};
test_output[12056:12063] = '{32'h415c8fbf, 32'h41a38dc1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12064:12071] = '{32'h4297257c, 32'hc2711590, 32'hc20e5ab6, 32'hc1b8d767, 32'h4230e214, 32'hc296a174, 32'hc2a8b7b6, 32'hc10295bc};
test_output[12064:12071] = '{32'h4297257c, 32'h0, 32'h0, 32'h0, 32'h4230e214, 32'h0, 32'h0, 32'h0};
test_input[12072:12079] = '{32'h40af7c0a, 32'hc1d9d63e, 32'h42758e20, 32'hc2938bb6, 32'hc28da05d, 32'h3f2a1252, 32'h425926b4, 32'hc2a3e7b6};
test_output[12072:12079] = '{32'h40af7c0a, 32'h0, 32'h42758e20, 32'h0, 32'h0, 32'h3f2a1252, 32'h425926b4, 32'h0};
test_input[12080:12087] = '{32'h41dea898, 32'h428c5729, 32'hc232cccb, 32'hc1885555, 32'h42c0d524, 32'h42130d4d, 32'hc2880ca0, 32'hc27839fa};
test_output[12080:12087] = '{32'h41dea898, 32'h428c5729, 32'h0, 32'h0, 32'h42c0d524, 32'h42130d4d, 32'h0, 32'h0};
test_input[12088:12095] = '{32'hc238e44b, 32'h418a7e9b, 32'h42b402c4, 32'h421b9b00, 32'hc2953646, 32'h42c00e30, 32'hc0810762, 32'h42aa93d1};
test_output[12088:12095] = '{32'h0, 32'h418a7e9b, 32'h42b402c4, 32'h421b9b00, 32'h0, 32'h42c00e30, 32'h0, 32'h42aa93d1};
test_input[12096:12103] = '{32'hbe4c94e1, 32'hc1ed2fc7, 32'h41dd0015, 32'h42a154ca, 32'h4285e5b4, 32'h414f822e, 32'hc1355458, 32'hc0a94ed2};
test_output[12096:12103] = '{32'h0, 32'h0, 32'h41dd0015, 32'h42a154ca, 32'h4285e5b4, 32'h414f822e, 32'h0, 32'h0};
test_input[12104:12111] = '{32'h42756937, 32'hc28ecf1b, 32'h42b59927, 32'h420fc4ec, 32'hc2bb22b3, 32'hc0fefe89, 32'hc2737427, 32'hc18c4faf};
test_output[12104:12111] = '{32'h42756937, 32'h0, 32'h42b59927, 32'h420fc4ec, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12112:12119] = '{32'h42afe299, 32'h41a8821d, 32'hc2909129, 32'h42bb5f0a, 32'hc2817ed9, 32'h417a01c7, 32'h42a96f1c, 32'hc2c5104a};
test_output[12112:12119] = '{32'h42afe299, 32'h41a8821d, 32'h0, 32'h42bb5f0a, 32'h0, 32'h417a01c7, 32'h42a96f1c, 32'h0};
test_input[12120:12127] = '{32'hc2b81ad9, 32'hc2829bc8, 32'h42b653cd, 32'h42b63c35, 32'hc263913c, 32'h41400f4e, 32'hc21a0376, 32'h4285a11a};
test_output[12120:12127] = '{32'h0, 32'h0, 32'h42b653cd, 32'h42b63c35, 32'h0, 32'h41400f4e, 32'h0, 32'h4285a11a};
test_input[12128:12135] = '{32'h40dd5c85, 32'hc180f905, 32'hc256dafc, 32'h426b0818, 32'h425ced3b, 32'hc2a42233, 32'h3f19e8c8, 32'hc26cd93f};
test_output[12128:12135] = '{32'h40dd5c85, 32'h0, 32'h0, 32'h426b0818, 32'h425ced3b, 32'h0, 32'h3f19e8c8, 32'h0};
test_input[12136:12143] = '{32'h40a7469b, 32'hc1bc077a, 32'h424e29a6, 32'h428389c5, 32'hc2950e21, 32'h42198e00, 32'h426c342e, 32'h41640a2f};
test_output[12136:12143] = '{32'h40a7469b, 32'h0, 32'h424e29a6, 32'h428389c5, 32'h0, 32'h42198e00, 32'h426c342e, 32'h41640a2f};
test_input[12144:12151] = '{32'h42016c04, 32'h41943561, 32'hc1a7db19, 32'hc25faa79, 32'h41eb3b24, 32'hc190aee4, 32'h42699506, 32'hc252cb6d};
test_output[12144:12151] = '{32'h42016c04, 32'h41943561, 32'h0, 32'h0, 32'h41eb3b24, 32'h0, 32'h42699506, 32'h0};
test_input[12152:12159] = '{32'h4190d55a, 32'hc233a859, 32'hc230af9c, 32'h42892e46, 32'hc270d00c, 32'hbf366779, 32'hc28016b8, 32'h42c65620};
test_output[12152:12159] = '{32'h4190d55a, 32'h0, 32'h0, 32'h42892e46, 32'h0, 32'h0, 32'h0, 32'h42c65620};
test_input[12160:12167] = '{32'hc2a5d0be, 32'h426b8e18, 32'hc1be8305, 32'h424e4e51, 32'hc2840958, 32'hc2aa7522, 32'hc2244e0d, 32'hc25e98d9};
test_output[12160:12167] = '{32'h0, 32'h426b8e18, 32'h0, 32'h424e4e51, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12168:12175] = '{32'hc1fed00d, 32'hc1af3aa3, 32'hc2877860, 32'h42bc3696, 32'h41c9b5ca, 32'hc28129d4, 32'h4281b856, 32'h4143f440};
test_output[12168:12175] = '{32'h0, 32'h0, 32'h0, 32'h42bc3696, 32'h41c9b5ca, 32'h0, 32'h4281b856, 32'h4143f440};
test_input[12176:12183] = '{32'hc25a9129, 32'hc2b3505d, 32'hbed7332c, 32'h41fd6df2, 32'hc26f1e8d, 32'hc21ff22b, 32'h42bc07cf, 32'h41b84aa0};
test_output[12176:12183] = '{32'h0, 32'h0, 32'h0, 32'h41fd6df2, 32'h0, 32'h0, 32'h42bc07cf, 32'h41b84aa0};
test_input[12184:12191] = '{32'h42a6d451, 32'h41c98cc2, 32'h425c9ba6, 32'hc299c5dc, 32'h41603a3f, 32'hc2221da7, 32'h42ab40c5, 32'hc16dbc26};
test_output[12184:12191] = '{32'h42a6d451, 32'h41c98cc2, 32'h425c9ba6, 32'h0, 32'h41603a3f, 32'h0, 32'h42ab40c5, 32'h0};
test_input[12192:12199] = '{32'hc2581441, 32'h4282b980, 32'h4258adf3, 32'h42be9d31, 32'hc122ebf9, 32'h42bbbd42, 32'hc263f359, 32'hc2abc330};
test_output[12192:12199] = '{32'h0, 32'h4282b980, 32'h4258adf3, 32'h42be9d31, 32'h0, 32'h42bbbd42, 32'h0, 32'h0};
test_input[12200:12207] = '{32'h42a18147, 32'h42c5d916, 32'hc253c6f0, 32'h4036fec7, 32'h41cf2668, 32'h428291bc, 32'h429c58ae, 32'h42b4b3d3};
test_output[12200:12207] = '{32'h42a18147, 32'h42c5d916, 32'h0, 32'h4036fec7, 32'h41cf2668, 32'h428291bc, 32'h429c58ae, 32'h42b4b3d3};
test_input[12208:12215] = '{32'hc14d82c0, 32'hc240a6d6, 32'hc2a2debb, 32'h427bac12, 32'h420582ff, 32'h42b485bc, 32'h40d2e6c6, 32'h4181f04a};
test_output[12208:12215] = '{32'h0, 32'h0, 32'h0, 32'h427bac12, 32'h420582ff, 32'h42b485bc, 32'h40d2e6c6, 32'h4181f04a};
test_input[12216:12223] = '{32'h41eb12b7, 32'hc2b91054, 32'h4205c747, 32'hc2963041, 32'h42918777, 32'h428c5c82, 32'hc1e6142f, 32'hc124df7a};
test_output[12216:12223] = '{32'h41eb12b7, 32'h0, 32'h4205c747, 32'h0, 32'h42918777, 32'h428c5c82, 32'h0, 32'h0};
test_input[12224:12231] = '{32'h42aa7878, 32'hc2247dc5, 32'h41ef0f22, 32'hc275be04, 32'hc1b21814, 32'hc22e5bf3, 32'h42b78fe9, 32'hc205c9ad};
test_output[12224:12231] = '{32'h42aa7878, 32'h0, 32'h41ef0f22, 32'h0, 32'h0, 32'h0, 32'h42b78fe9, 32'h0};
test_input[12232:12239] = '{32'hbfd0d235, 32'hc26ce2c6, 32'h4283dae5, 32'hc14fa76f, 32'h419681c2, 32'h4175e3fe, 32'h419c35b3, 32'h41483b8c};
test_output[12232:12239] = '{32'h0, 32'h0, 32'h4283dae5, 32'h0, 32'h419681c2, 32'h4175e3fe, 32'h419c35b3, 32'h41483b8c};
test_input[12240:12247] = '{32'h4234b405, 32'h41b4349a, 32'hc2245314, 32'h413be1c4, 32'hc24d5885, 32'h42649384, 32'h42a82b44, 32'hc112d85c};
test_output[12240:12247] = '{32'h4234b405, 32'h41b4349a, 32'h0, 32'h413be1c4, 32'h0, 32'h42649384, 32'h42a82b44, 32'h0};
test_input[12248:12255] = '{32'h42699be0, 32'hc21219e5, 32'hc2959915, 32'hc280d1b7, 32'h41c6abc8, 32'h42901f63, 32'hc22cd784, 32'h42aaaf91};
test_output[12248:12255] = '{32'h42699be0, 32'h0, 32'h0, 32'h0, 32'h41c6abc8, 32'h42901f63, 32'h0, 32'h42aaaf91};
test_input[12256:12263] = '{32'h420842d1, 32'h3fc00d4f, 32'hc145f2aa, 32'hc18e0bba, 32'h42bc6522, 32'h42afa6e9, 32'hc254251a, 32'h408db85b};
test_output[12256:12263] = '{32'h420842d1, 32'h3fc00d4f, 32'h0, 32'h0, 32'h42bc6522, 32'h42afa6e9, 32'h0, 32'h408db85b};
test_input[12264:12271] = '{32'hc0fbdc6a, 32'h41b643b0, 32'hc2ae01e8, 32'hc26990a0, 32'hc272b845, 32'hc2828732, 32'hc1ef5309, 32'h428684dd};
test_output[12264:12271] = '{32'h0, 32'h41b643b0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428684dd};
test_input[12272:12279] = '{32'h404390b9, 32'h41a33bc3, 32'hc13688e7, 32'hc0a26029, 32'hc175c723, 32'h40ccd4ef, 32'h4224ab85, 32'h414384de};
test_output[12272:12279] = '{32'h404390b9, 32'h41a33bc3, 32'h0, 32'h0, 32'h0, 32'h40ccd4ef, 32'h4224ab85, 32'h414384de};
test_input[12280:12287] = '{32'h3fd80abb, 32'hc26444f8, 32'hc28aa5b9, 32'hc20873e8, 32'h42898bcf, 32'hc2619ccc, 32'hc22a2c22, 32'h4245fb38};
test_output[12280:12287] = '{32'h3fd80abb, 32'h0, 32'h0, 32'h0, 32'h42898bcf, 32'h0, 32'h0, 32'h4245fb38};
test_input[12288:12295] = '{32'h3fc2e96b, 32'hc2ad0c2c, 32'hc2674ed8, 32'hc17f3fdd, 32'hc2bfd604, 32'hc27cc235, 32'hc288cc73, 32'hc28a7420};
test_output[12288:12295] = '{32'h3fc2e96b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12296:12303] = '{32'h42a92b9c, 32'hc254576f, 32'h420859e5, 32'hc16728c1, 32'hc1ea6153, 32'hc26c73a5, 32'h42738c71, 32'hc18c7825};
test_output[12296:12303] = '{32'h42a92b9c, 32'h0, 32'h420859e5, 32'h0, 32'h0, 32'h0, 32'h42738c71, 32'h0};
test_input[12304:12311] = '{32'hc29fbd55, 32'h42ac02fb, 32'hc10b5015, 32'h428acc67, 32'h41a2a816, 32'h41752b31, 32'h42190779, 32'h42a587f6};
test_output[12304:12311] = '{32'h0, 32'h42ac02fb, 32'h0, 32'h428acc67, 32'h41a2a816, 32'h41752b31, 32'h42190779, 32'h42a587f6};
test_input[12312:12319] = '{32'hc196916d, 32'hc200a996, 32'h42ae54bd, 32'h422e0f6e, 32'hc0e1f6c5, 32'hc1e95594, 32'hc292f711, 32'h42a7d6fc};
test_output[12312:12319] = '{32'h0, 32'h0, 32'h42ae54bd, 32'h422e0f6e, 32'h0, 32'h0, 32'h0, 32'h42a7d6fc};
test_input[12320:12327] = '{32'h41a7aa78, 32'h4259b225, 32'h4214f158, 32'h42b63009, 32'hc03d4ec7, 32'hc276f3b1, 32'hc2b66590, 32'h42a21cf4};
test_output[12320:12327] = '{32'h41a7aa78, 32'h4259b225, 32'h4214f158, 32'h42b63009, 32'h0, 32'h0, 32'h0, 32'h42a21cf4};
test_input[12328:12335] = '{32'h41ffe0ce, 32'hc2934dcb, 32'h4234f715, 32'hc28d09c6, 32'h426ee91d, 32'hc1b86435, 32'hc200e672, 32'hc23b8ee1};
test_output[12328:12335] = '{32'h41ffe0ce, 32'h0, 32'h4234f715, 32'h0, 32'h426ee91d, 32'h0, 32'h0, 32'h0};
test_input[12336:12343] = '{32'h42ac68fc, 32'hc2be027d, 32'h424fb83d, 32'hc0caf887, 32'hc1a77e13, 32'hc2929476, 32'hc2197711, 32'hc2a3abbb};
test_output[12336:12343] = '{32'h42ac68fc, 32'h0, 32'h424fb83d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12344:12351] = '{32'h42342e5f, 32'h41f7a9b9, 32'h4280f54b, 32'hc214b080, 32'h421d4812, 32'h42bb20b6, 32'hc2916221, 32'hc288f9a3};
test_output[12344:12351] = '{32'h42342e5f, 32'h41f7a9b9, 32'h4280f54b, 32'h0, 32'h421d4812, 32'h42bb20b6, 32'h0, 32'h0};
test_input[12352:12359] = '{32'hc1862094, 32'h42702e77, 32'hc2783069, 32'hc1a5ee4e, 32'h42104bda, 32'hc28b8539, 32'hc29c1f7c, 32'h422bcb11};
test_output[12352:12359] = '{32'h0, 32'h42702e77, 32'h0, 32'h0, 32'h42104bda, 32'h0, 32'h0, 32'h422bcb11};
test_input[12360:12367] = '{32'hc26ac791, 32'h42016ef7, 32'hc1b10c66, 32'h42b59d04, 32'h4248b2db, 32'h42287ce5, 32'hc22954ac, 32'hc1e636e8};
test_output[12360:12367] = '{32'h0, 32'h42016ef7, 32'h0, 32'h42b59d04, 32'h4248b2db, 32'h42287ce5, 32'h0, 32'h0};
test_input[12368:12375] = '{32'hc1b144a9, 32'h42801ad2, 32'hc2b3d2a8, 32'hc28ee745, 32'hc27f279a, 32'h41ef9eef, 32'h41b20820, 32'hc2a748ec};
test_output[12368:12375] = '{32'h0, 32'h42801ad2, 32'h0, 32'h0, 32'h0, 32'h41ef9eef, 32'h41b20820, 32'h0};
test_input[12376:12383] = '{32'hc2138741, 32'hc221e0f5, 32'h4206de69, 32'h3fe120b3, 32'hc2b193f3, 32'h42b641e7, 32'h3f380b77, 32'h420edb6e};
test_output[12376:12383] = '{32'h0, 32'h0, 32'h4206de69, 32'h3fe120b3, 32'h0, 32'h42b641e7, 32'h3f380b77, 32'h420edb6e};
test_input[12384:12391] = '{32'h42be4238, 32'h42832a6c, 32'h42270aab, 32'h42763a18, 32'h4158bd3c, 32'hc1aadd48, 32'hc1d9b9fc, 32'hc277f41c};
test_output[12384:12391] = '{32'h42be4238, 32'h42832a6c, 32'h42270aab, 32'h42763a18, 32'h4158bd3c, 32'h0, 32'h0, 32'h0};
test_input[12392:12399] = '{32'hc22ed100, 32'hc221da23, 32'h41ea6cb1, 32'h42044158, 32'h42c1b80f, 32'h42925c8d, 32'hc08dfe33, 32'hc1125fd9};
test_output[12392:12399] = '{32'h0, 32'h0, 32'h41ea6cb1, 32'h42044158, 32'h42c1b80f, 32'h42925c8d, 32'h0, 32'h0};
test_input[12400:12407] = '{32'h41687a69, 32'h4197377e, 32'hc1592ea4, 32'hc228bb84, 32'hc03da3b0, 32'hc1e466e6, 32'hc26df045, 32'hc1ffccec};
test_output[12400:12407] = '{32'h41687a69, 32'h4197377e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12408:12415] = '{32'h425d1769, 32'h42ba085e, 32'hc2ba974f, 32'hc0e71766, 32'hc28e560f, 32'hc1f6ded4, 32'h422f20d8, 32'h41ba18df};
test_output[12408:12415] = '{32'h425d1769, 32'h42ba085e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422f20d8, 32'h41ba18df};
test_input[12416:12423] = '{32'hc28b1895, 32'h3e013e15, 32'h4251fa63, 32'h4223a622, 32'hc2a60618, 32'hc18bce78, 32'h42ab2431, 32'h4111862a};
test_output[12416:12423] = '{32'h0, 32'h3e013e15, 32'h4251fa63, 32'h4223a622, 32'h0, 32'h0, 32'h42ab2431, 32'h4111862a};
test_input[12424:12431] = '{32'h42b39cce, 32'h4154774b, 32'hc2b519d9, 32'hc250616f, 32'h4236f5cc, 32'hc19836cf, 32'hc15342f9, 32'h42aa9f99};
test_output[12424:12431] = '{32'h42b39cce, 32'h4154774b, 32'h0, 32'h0, 32'h4236f5cc, 32'h0, 32'h0, 32'h42aa9f99};
test_input[12432:12439] = '{32'hc288ff5d, 32'hc1ca0148, 32'hc2a7c158, 32'h42be92e5, 32'hc1e20b3e, 32'hc2641c8d, 32'hbec36820, 32'h42782c75};
test_output[12432:12439] = '{32'h0, 32'h0, 32'h0, 32'h42be92e5, 32'h0, 32'h0, 32'h0, 32'h42782c75};
test_input[12440:12447] = '{32'h42a82ac2, 32'h42398bcc, 32'h40a51231, 32'h42514308, 32'hc27a85e8, 32'hc1f71926, 32'hc27f423b, 32'hc18f9332};
test_output[12440:12447] = '{32'h42a82ac2, 32'h42398bcc, 32'h40a51231, 32'h42514308, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12448:12455] = '{32'hbf81ee59, 32'hc1aff8df, 32'hc254d624, 32'hc2a00579, 32'h4215e066, 32'h42b54e55, 32'hc2b3b7aa, 32'hc296b75c};
test_output[12448:12455] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4215e066, 32'h42b54e55, 32'h0, 32'h0};
test_input[12456:12463] = '{32'hc2c192b0, 32'hc29e9cf7, 32'h41cffa38, 32'h41f0aa68, 32'hc25b8096, 32'h42599871, 32'hc2bfae1f, 32'h41fa6b44};
test_output[12456:12463] = '{32'h0, 32'h0, 32'h41cffa38, 32'h41f0aa68, 32'h0, 32'h42599871, 32'h0, 32'h41fa6b44};
test_input[12464:12471] = '{32'h426937ba, 32'hc20c94b8, 32'h429665d7, 32'h420f6468, 32'hc1841e5e, 32'h41887193, 32'hc0af8f25, 32'h42b28b1e};
test_output[12464:12471] = '{32'h426937ba, 32'h0, 32'h429665d7, 32'h420f6468, 32'h0, 32'h41887193, 32'h0, 32'h42b28b1e};
test_input[12472:12479] = '{32'hc101abec, 32'hc2a140ba, 32'h42b73ae7, 32'h41a89943, 32'hc23077f7, 32'h4015d03d, 32'hc2799c5c, 32'h42803fb4};
test_output[12472:12479] = '{32'h0, 32'h0, 32'h42b73ae7, 32'h41a89943, 32'h0, 32'h4015d03d, 32'h0, 32'h42803fb4};
test_input[12480:12487] = '{32'hc2ad4f91, 32'hc214a703, 32'hc1932363, 32'h40da1b61, 32'hc2735282, 32'hc1cf1394, 32'hc2362203, 32'hc106f1aa};
test_output[12480:12487] = '{32'h0, 32'h0, 32'h0, 32'h40da1b61, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12488:12495] = '{32'hc27e02ce, 32'h4208f70e, 32'hc2a84029, 32'hc2b409ad, 32'hc14b662b, 32'h4206e065, 32'h42457693, 32'h419d77ac};
test_output[12488:12495] = '{32'h0, 32'h4208f70e, 32'h0, 32'h0, 32'h0, 32'h4206e065, 32'h42457693, 32'h419d77ac};
test_input[12496:12503] = '{32'hc233bc85, 32'h41b6758a, 32'h3ef38f0d, 32'h41df0c4d, 32'h4211da4e, 32'hc2c66e6f, 32'hc1c2b6f4, 32'h42b2bb14};
test_output[12496:12503] = '{32'h0, 32'h41b6758a, 32'h3ef38f0d, 32'h41df0c4d, 32'h4211da4e, 32'h0, 32'h0, 32'h42b2bb14};
test_input[12504:12511] = '{32'hc21b90f9, 32'h427b4580, 32'h41cfdf3e, 32'h424184b3, 32'h427f1f19, 32'h40f9ce33, 32'hc0625ead, 32'hc2c27dc8};
test_output[12504:12511] = '{32'h0, 32'h427b4580, 32'h41cfdf3e, 32'h424184b3, 32'h427f1f19, 32'h40f9ce33, 32'h0, 32'h0};
test_input[12512:12519] = '{32'hc2094959, 32'hc2603759, 32'hc29fad44, 32'h41afba86, 32'hc246a2b2, 32'hc24ab7e5, 32'h42a04852, 32'hc1078316};
test_output[12512:12519] = '{32'h0, 32'h0, 32'h0, 32'h41afba86, 32'h0, 32'h0, 32'h42a04852, 32'h0};
test_input[12520:12527] = '{32'h427e9709, 32'h4291203e, 32'hc2c557f0, 32'h42bfa7de, 32'hc22246a4, 32'h40e37db3, 32'h42818587, 32'hc275f3d2};
test_output[12520:12527] = '{32'h427e9709, 32'h4291203e, 32'h0, 32'h42bfa7de, 32'h0, 32'h40e37db3, 32'h42818587, 32'h0};
test_input[12528:12535] = '{32'h42b59ce5, 32'h42a9f567, 32'h42a67379, 32'hc13c0415, 32'h410aac6a, 32'h42c6066f, 32'hc0b35600, 32'hc19abed6};
test_output[12528:12535] = '{32'h42b59ce5, 32'h42a9f567, 32'h42a67379, 32'h0, 32'h410aac6a, 32'h42c6066f, 32'h0, 32'h0};
test_input[12536:12543] = '{32'h41a8fc69, 32'h42452303, 32'h4281bde6, 32'h4241f6cd, 32'h422af0a8, 32'h40f5bf9c, 32'hc2a4384f, 32'h413badf2};
test_output[12536:12543] = '{32'h41a8fc69, 32'h42452303, 32'h4281bde6, 32'h4241f6cd, 32'h422af0a8, 32'h40f5bf9c, 32'h0, 32'h413badf2};
test_input[12544:12551] = '{32'h41c107b7, 32'hc20d3b74, 32'h41ce8512, 32'hc298a917, 32'hc28bbcf5, 32'hc21b524a, 32'h417b2974, 32'h42c3d49d};
test_output[12544:12551] = '{32'h41c107b7, 32'h0, 32'h41ce8512, 32'h0, 32'h0, 32'h0, 32'h417b2974, 32'h42c3d49d};
test_input[12552:12559] = '{32'h40195afa, 32'hc2c31d3c, 32'hc28aad2e, 32'h4283b4fe, 32'hc2c60f29, 32'h41361f68, 32'h4199586e, 32'hc2619e73};
test_output[12552:12559] = '{32'h40195afa, 32'h0, 32'h0, 32'h4283b4fe, 32'h0, 32'h41361f68, 32'h4199586e, 32'h0};
test_input[12560:12567] = '{32'hc1ce4658, 32'h428d3a71, 32'hc1d184e6, 32'h4171b144, 32'hc2a889fd, 32'h428a58a2, 32'hc2ac8931, 32'h4219a3d7};
test_output[12560:12567] = '{32'h0, 32'h428d3a71, 32'h0, 32'h4171b144, 32'h0, 32'h428a58a2, 32'h0, 32'h4219a3d7};
test_input[12568:12575] = '{32'hc2072d39, 32'hc0b82345, 32'h42ac159f, 32'h41bb6130, 32'h41443b14, 32'h40eafcaa, 32'h423eaf89, 32'hc2a34ef2};
test_output[12568:12575] = '{32'h0, 32'h0, 32'h42ac159f, 32'h41bb6130, 32'h41443b14, 32'h40eafcaa, 32'h423eaf89, 32'h0};
test_input[12576:12583] = '{32'hc246e5a6, 32'hc011c052, 32'hc2799e9d, 32'h42a036da, 32'h4243e646, 32'hc2a46055, 32'h4092c930, 32'h41cc2d22};
test_output[12576:12583] = '{32'h0, 32'h0, 32'h0, 32'h42a036da, 32'h4243e646, 32'h0, 32'h4092c930, 32'h41cc2d22};
test_input[12584:12591] = '{32'hc2b8aa46, 32'h42b5123b, 32'hc2b5beed, 32'h41cb7c56, 32'h42b0c4f0, 32'hc239bcb6, 32'hc24199be, 32'hc19d033f};
test_output[12584:12591] = '{32'h0, 32'h42b5123b, 32'h0, 32'h41cb7c56, 32'h42b0c4f0, 32'h0, 32'h0, 32'h0};
test_input[12592:12599] = '{32'h41953e52, 32'h41bc6f4f, 32'hc29847d6, 32'h41b7e408, 32'h421b5436, 32'h429e6bde, 32'hc2c68095, 32'hc2afbb03};
test_output[12592:12599] = '{32'h41953e52, 32'h41bc6f4f, 32'h0, 32'h41b7e408, 32'h421b5436, 32'h429e6bde, 32'h0, 32'h0};
test_input[12600:12607] = '{32'hc1c6df59, 32'h425962f4, 32'h42acf50b, 32'hc2076016, 32'h426e3ead, 32'h420d3107, 32'h41b6ce29, 32'h42625b89};
test_output[12600:12607] = '{32'h0, 32'h425962f4, 32'h42acf50b, 32'h0, 32'h426e3ead, 32'h420d3107, 32'h41b6ce29, 32'h42625b89};
test_input[12608:12615] = '{32'h42934881, 32'h420f4b1c, 32'h422629d3, 32'h410512e8, 32'h402fbc56, 32'hc2abf75d, 32'hc1183622, 32'hc1d0ff45};
test_output[12608:12615] = '{32'h42934881, 32'h420f4b1c, 32'h422629d3, 32'h410512e8, 32'h402fbc56, 32'h0, 32'h0, 32'h0};
test_input[12616:12623] = '{32'hc2c52f1d, 32'h41b6b81c, 32'h41b56e15, 32'h426434d3, 32'hc2a4b711, 32'h40bb639a, 32'h42995bd0, 32'hc1ab19d5};
test_output[12616:12623] = '{32'h0, 32'h41b6b81c, 32'h41b56e15, 32'h426434d3, 32'h0, 32'h40bb639a, 32'h42995bd0, 32'h0};
test_input[12624:12631] = '{32'hc27ad5f2, 32'hc24e1de5, 32'hc1babc8c, 32'h417f6ba1, 32'hc2574863, 32'hc24a87d0, 32'h4184b7de, 32'h422ef286};
test_output[12624:12631] = '{32'h0, 32'h0, 32'h0, 32'h417f6ba1, 32'h0, 32'h0, 32'h4184b7de, 32'h422ef286};
test_input[12632:12639] = '{32'hc0ff50cb, 32'h40957a56, 32'hc290b8d9, 32'hc28bde2f, 32'h4231d154, 32'h429d8a15, 32'hc2aadd39, 32'hc25d7972};
test_output[12632:12639] = '{32'h0, 32'h40957a56, 32'h0, 32'h0, 32'h4231d154, 32'h429d8a15, 32'h0, 32'h0};
test_input[12640:12647] = '{32'hc2bdef12, 32'hc154ddce, 32'h4236e156, 32'h40ec4144, 32'hc1932c2f, 32'hc20c59f7, 32'hc1e2406f, 32'hc2a780bf};
test_output[12640:12647] = '{32'h0, 32'h0, 32'h4236e156, 32'h40ec4144, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12648:12655] = '{32'hc22056a4, 32'hc2a1c8a3, 32'h41e99ee1, 32'hc230126b, 32'hc2972c74, 32'h41a15860, 32'h42a8e298, 32'h42599a99};
test_output[12648:12655] = '{32'h0, 32'h0, 32'h41e99ee1, 32'h0, 32'h0, 32'h41a15860, 32'h42a8e298, 32'h42599a99};
test_input[12656:12663] = '{32'hc21c09bb, 32'hc1c222c7, 32'hc1981bbd, 32'hc11f726e, 32'hc1d9f389, 32'h42c74639, 32'hc18e2305, 32'h4281b09c};
test_output[12656:12663] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c74639, 32'h0, 32'h4281b09c};
test_input[12664:12671] = '{32'hc2b9dc92, 32'h42774529, 32'hc1e248ff, 32'h427e1bc6, 32'h424549e8, 32'h4263e199, 32'h41f7c8c3, 32'h42b36767};
test_output[12664:12671] = '{32'h0, 32'h42774529, 32'h0, 32'h427e1bc6, 32'h424549e8, 32'h4263e199, 32'h41f7c8c3, 32'h42b36767};
test_input[12672:12679] = '{32'h41c6e371, 32'h41d02fa6, 32'h42a89f16, 32'h4083986a, 32'h422d534d, 32'hc0eaa21a, 32'h42ab8ef6, 32'h42ad33d6};
test_output[12672:12679] = '{32'h41c6e371, 32'h41d02fa6, 32'h42a89f16, 32'h4083986a, 32'h422d534d, 32'h0, 32'h42ab8ef6, 32'h42ad33d6};
test_input[12680:12687] = '{32'h41449735, 32'hc1fe8caf, 32'hc23659e2, 32'h4292d96a, 32'hc26d3a67, 32'h41d4993c, 32'hc2bc78b4, 32'hc2a15b98};
test_output[12680:12687] = '{32'h41449735, 32'h0, 32'h0, 32'h4292d96a, 32'h0, 32'h41d4993c, 32'h0, 32'h0};
test_input[12688:12695] = '{32'hc143fafb, 32'hc196ffe6, 32'hc2238cd8, 32'hc2125179, 32'h420c7ba1, 32'hc2a88b81, 32'h41114494, 32'hc292378e};
test_output[12688:12695] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h420c7ba1, 32'h0, 32'h41114494, 32'h0};
test_input[12696:12703] = '{32'hc2474997, 32'h3f063a4a, 32'h41d9cf94, 32'hc29bd64d, 32'h41f82a60, 32'h3e52b877, 32'hc1a9fd1e, 32'hc16d0349};
test_output[12696:12703] = '{32'h0, 32'h3f063a4a, 32'h41d9cf94, 32'h0, 32'h41f82a60, 32'h3e52b877, 32'h0, 32'h0};
test_input[12704:12711] = '{32'h41fcb1aa, 32'hc0ae54d7, 32'h41e4338b, 32'hc18cd0fe, 32'h42b8e40e, 32'hc2036d3b, 32'h42b02537, 32'h42a780a5};
test_output[12704:12711] = '{32'h41fcb1aa, 32'h0, 32'h41e4338b, 32'h0, 32'h42b8e40e, 32'h0, 32'h42b02537, 32'h42a780a5};
test_input[12712:12719] = '{32'h428d1f4e, 32'hc028c6ed, 32'hc18348d4, 32'h42c10f7a, 32'h41d1485a, 32'hc1a7e2c1, 32'h42aad1a5, 32'h424170c3};
test_output[12712:12719] = '{32'h428d1f4e, 32'h0, 32'h0, 32'h42c10f7a, 32'h41d1485a, 32'h0, 32'h42aad1a5, 32'h424170c3};
test_input[12720:12727] = '{32'hc232b513, 32'hc276806d, 32'h426875fb, 32'hc219d059, 32'h406a11ae, 32'hc19b64fd, 32'hc03d930e, 32'h42b52c31};
test_output[12720:12727] = '{32'h0, 32'h0, 32'h426875fb, 32'h0, 32'h406a11ae, 32'h0, 32'h0, 32'h42b52c31};
test_input[12728:12735] = '{32'h410d31c2, 32'h429be2be, 32'h4246f4a0, 32'hc2432a8d, 32'h4264ed11, 32'h4085e09d, 32'hc2359c96, 32'h42c2f6bc};
test_output[12728:12735] = '{32'h410d31c2, 32'h429be2be, 32'h4246f4a0, 32'h0, 32'h4264ed11, 32'h4085e09d, 32'h0, 32'h42c2f6bc};
test_input[12736:12743] = '{32'h422048ff, 32'hc297b2f5, 32'h426383c9, 32'hc1e052ad, 32'hc202e110, 32'hc1ccd1c3, 32'hc23b787b, 32'hc222494f};
test_output[12736:12743] = '{32'h422048ff, 32'h0, 32'h426383c9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12744:12751] = '{32'hc215f5a8, 32'hc28c0576, 32'hc2be54bd, 32'hc28e2040, 32'h4270a134, 32'h423ba5d6, 32'h42755ac0, 32'hc0a317fc};
test_output[12744:12751] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4270a134, 32'h423ba5d6, 32'h42755ac0, 32'h0};
test_input[12752:12759] = '{32'hc2601d01, 32'hc00f8523, 32'h41b8daa3, 32'hc2b66b26, 32'h425e1a20, 32'hc2361875, 32'hc27deb55, 32'hc1c331a8};
test_output[12752:12759] = '{32'h0, 32'h0, 32'h41b8daa3, 32'h0, 32'h425e1a20, 32'h0, 32'h0, 32'h0};
test_input[12760:12767] = '{32'h4200fd17, 32'hc2a2a548, 32'hc0ab132b, 32'hc2aef0f2, 32'h41f11035, 32'h4295ffcd, 32'h41c9b12f, 32'hc2bbdb52};
test_output[12760:12767] = '{32'h4200fd17, 32'h0, 32'h0, 32'h0, 32'h41f11035, 32'h4295ffcd, 32'h41c9b12f, 32'h0};
test_input[12768:12775] = '{32'h423aaecd, 32'hc18c4a10, 32'hc26990bb, 32'h4206c2d3, 32'hc20e3bd3, 32'hc2b89289, 32'h429668ce, 32'h428cb448};
test_output[12768:12775] = '{32'h423aaecd, 32'h0, 32'h0, 32'h4206c2d3, 32'h0, 32'h0, 32'h429668ce, 32'h428cb448};
test_input[12776:12783] = '{32'hc1a74d4d, 32'h42865a67, 32'h42c6266e, 32'h42aef222, 32'hc2ad199f, 32'hc29e4a19, 32'h420355fd, 32'hc236944e};
test_output[12776:12783] = '{32'h0, 32'h42865a67, 32'h42c6266e, 32'h42aef222, 32'h0, 32'h0, 32'h420355fd, 32'h0};
test_input[12784:12791] = '{32'hc225a2c4, 32'hc18359f6, 32'hc26e1e2b, 32'h42813c0f, 32'hc2116dd2, 32'h42befba9, 32'h429ea087, 32'hc2bff068};
test_output[12784:12791] = '{32'h0, 32'h0, 32'h0, 32'h42813c0f, 32'h0, 32'h42befba9, 32'h429ea087, 32'h0};
test_input[12792:12799] = '{32'hc251e2a7, 32'h427075b7, 32'hbfea48e7, 32'hc22d1442, 32'h413b0262, 32'hc2b08594, 32'hc226ce62, 32'h419440f0};
test_output[12792:12799] = '{32'h0, 32'h427075b7, 32'h0, 32'h0, 32'h413b0262, 32'h0, 32'h0, 32'h419440f0};
test_input[12800:12807] = '{32'hc220067b, 32'h42ab9fe4, 32'hc24bac88, 32'hc18a98d7, 32'hc0c30fa6, 32'hc1dba401, 32'h42bc948d, 32'h422f12ff};
test_output[12800:12807] = '{32'h0, 32'h42ab9fe4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bc948d, 32'h422f12ff};
test_input[12808:12815] = '{32'h42b462d8, 32'hc2862185, 32'h42b45726, 32'hc2b126d5, 32'h41a8b978, 32'hc284b695, 32'h42aee00a, 32'h424107ab};
test_output[12808:12815] = '{32'h42b462d8, 32'h0, 32'h42b45726, 32'h0, 32'h41a8b978, 32'h0, 32'h42aee00a, 32'h424107ab};
test_input[12816:12823] = '{32'h421c75b1, 32'hc2878f39, 32'h429d9c52, 32'hc2ace5da, 32'hc28797ba, 32'hc264143e, 32'h3ef4239a, 32'hc2287819};
test_output[12816:12823] = '{32'h421c75b1, 32'h0, 32'h429d9c52, 32'h0, 32'h0, 32'h0, 32'h3ef4239a, 32'h0};
test_input[12824:12831] = '{32'hc1541d7c, 32'hc29bf071, 32'h4095dbd8, 32'hc2b8b76f, 32'hc10d6302, 32'h41f78fcd, 32'hc21fbcb0, 32'hc29afb7a};
test_output[12824:12831] = '{32'h0, 32'h0, 32'h4095dbd8, 32'h0, 32'h0, 32'h41f78fcd, 32'h0, 32'h0};
test_input[12832:12839] = '{32'h41f365aa, 32'hc26dd0dd, 32'h427058fb, 32'hc2963ec9, 32'hc2583746, 32'h420a46f5, 32'hc288a9f1, 32'hc2334fbf};
test_output[12832:12839] = '{32'h41f365aa, 32'h0, 32'h427058fb, 32'h0, 32'h0, 32'h420a46f5, 32'h0, 32'h0};
test_input[12840:12847] = '{32'h41f4397d, 32'hc2bbe1cf, 32'h424dae3a, 32'h42c15990, 32'h423c9301, 32'hc20d2570, 32'hc2b28626, 32'hc29ae401};
test_output[12840:12847] = '{32'h41f4397d, 32'h0, 32'h424dae3a, 32'h42c15990, 32'h423c9301, 32'h0, 32'h0, 32'h0};
test_input[12848:12855] = '{32'hc28ea32e, 32'hbec20a8c, 32'h40ff9737, 32'h42835a13, 32'h4245c1e5, 32'h42791ca9, 32'hc27218cf, 32'hc238d9a3};
test_output[12848:12855] = '{32'h0, 32'h0, 32'h40ff9737, 32'h42835a13, 32'h4245c1e5, 32'h42791ca9, 32'h0, 32'h0};
test_input[12856:12863] = '{32'hc1ae8354, 32'h42342b3a, 32'h42844a9b, 32'hc2822045, 32'h4081f779, 32'h428dc180, 32'h41f9ce3d, 32'hc1e5eb83};
test_output[12856:12863] = '{32'h0, 32'h42342b3a, 32'h42844a9b, 32'h0, 32'h4081f779, 32'h428dc180, 32'h41f9ce3d, 32'h0};
test_input[12864:12871] = '{32'h4299ddea, 32'h42c247b6, 32'hc2643f75, 32'h42ac9b35, 32'hc28b2d97, 32'hc23d451e, 32'hc2bd4434, 32'h429e0dec};
test_output[12864:12871] = '{32'h4299ddea, 32'h42c247b6, 32'h0, 32'h42ac9b35, 32'h0, 32'h0, 32'h0, 32'h429e0dec};
test_input[12872:12879] = '{32'h4286c2d7, 32'hc1874e7a, 32'hc2ae396c, 32'hc2a49b89, 32'h419c1d6d, 32'h4293f7eb, 32'h424bc355, 32'hc238662c};
test_output[12872:12879] = '{32'h4286c2d7, 32'h0, 32'h0, 32'h0, 32'h419c1d6d, 32'h4293f7eb, 32'h424bc355, 32'h0};
test_input[12880:12887] = '{32'h41c40928, 32'hc24181ec, 32'h4237bbb6, 32'hc1b3ed6e, 32'h428f7ab8, 32'h42c54ad1, 32'h41a5a79f, 32'hbfa7d831};
test_output[12880:12887] = '{32'h41c40928, 32'h0, 32'h4237bbb6, 32'h0, 32'h428f7ab8, 32'h42c54ad1, 32'h41a5a79f, 32'h0};
test_input[12888:12895] = '{32'h42245782, 32'h41f80dd1, 32'hc0198d9a, 32'h417f3ae6, 32'h42673db2, 32'hc1e88c91, 32'hc281e053, 32'hc1a8caf0};
test_output[12888:12895] = '{32'h42245782, 32'h41f80dd1, 32'h0, 32'h417f3ae6, 32'h42673db2, 32'h0, 32'h0, 32'h0};
test_input[12896:12903] = '{32'h412c05dc, 32'hc29b115f, 32'hc19c06a5, 32'h41c5fd38, 32'hbf5163bd, 32'hc130462b, 32'h4096d5f6, 32'hc109ddf3};
test_output[12896:12903] = '{32'h412c05dc, 32'h0, 32'h0, 32'h41c5fd38, 32'h0, 32'h0, 32'h4096d5f6, 32'h0};
test_input[12904:12911] = '{32'hc1bfe185, 32'hc26aa542, 32'h4274756f, 32'hc24784d4, 32'hc1e409bb, 32'hc0436499, 32'hc2c0aa15, 32'hc20438c2};
test_output[12904:12911] = '{32'h0, 32'h0, 32'h4274756f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12912:12919] = '{32'hc2a3c993, 32'h42a1a65d, 32'h4060ae30, 32'h4046bcfb, 32'hc2b5a70b, 32'h42844bd4, 32'hc13bf1ff, 32'hc2b3ac55};
test_output[12912:12919] = '{32'h0, 32'h42a1a65d, 32'h4060ae30, 32'h4046bcfb, 32'h0, 32'h42844bd4, 32'h0, 32'h0};
test_input[12920:12927] = '{32'hc274439e, 32'h40bd5f49, 32'h421e670b, 32'h40a2685d, 32'hbf58e582, 32'h420b7d0c, 32'h41a2fb85, 32'h419dec2e};
test_output[12920:12927] = '{32'h0, 32'h40bd5f49, 32'h421e670b, 32'h40a2685d, 32'h0, 32'h420b7d0c, 32'h41a2fb85, 32'h419dec2e};
test_input[12928:12935] = '{32'h420423ce, 32'hbf93ae9c, 32'hc2546dc0, 32'hc04d70e0, 32'hc28b43e8, 32'hc2571282, 32'h420a575c, 32'hc2ac0769};
test_output[12928:12935] = '{32'h420423ce, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420a575c, 32'h0};
test_input[12936:12943] = '{32'h42560a00, 32'h428f76e9, 32'hc22c21eb, 32'h4212a7b7, 32'h4139452a, 32'hc10d1239, 32'hc1b85196, 32'h424d0d47};
test_output[12936:12943] = '{32'h42560a00, 32'h428f76e9, 32'h0, 32'h4212a7b7, 32'h4139452a, 32'h0, 32'h0, 32'h424d0d47};
test_input[12944:12951] = '{32'hc2b79e90, 32'hc16d7b6e, 32'h428b00c6, 32'hc18bf4c3, 32'h42c5d498, 32'hc28e957c, 32'hc25c5cc9, 32'h42215367};
test_output[12944:12951] = '{32'h0, 32'h0, 32'h428b00c6, 32'h0, 32'h42c5d498, 32'h0, 32'h0, 32'h42215367};
test_input[12952:12959] = '{32'hc26c1116, 32'hc2a45753, 32'hc290aede, 32'hc2813ba2, 32'hbeb364a6, 32'h42c654de, 32'hc20da8f3, 32'hc21d136d};
test_output[12952:12959] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c654de, 32'h0, 32'h0};
test_input[12960:12967] = '{32'hc2a9ff4c, 32'h42aecd08, 32'hc22877c2, 32'hc117b7df, 32'hc27eb1cc, 32'hc218536d, 32'h40f597a2, 32'h42882391};
test_output[12960:12967] = '{32'h0, 32'h42aecd08, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40f597a2, 32'h42882391};
test_input[12968:12975] = '{32'hc22907ab, 32'h42a038b2, 32'hc2a7ebb7, 32'h40b1920f, 32'hc23de898, 32'h4245fd5c, 32'h42212ae7, 32'hc2ab77f0};
test_output[12968:12975] = '{32'h0, 32'h42a038b2, 32'h0, 32'h40b1920f, 32'h0, 32'h4245fd5c, 32'h42212ae7, 32'h0};
test_input[12976:12983] = '{32'hc2449e59, 32'h424a0147, 32'h42655e16, 32'h4201e428, 32'hc21813ef, 32'h40d9f696, 32'h41369041, 32'h420ee777};
test_output[12976:12983] = '{32'h0, 32'h424a0147, 32'h42655e16, 32'h4201e428, 32'h0, 32'h40d9f696, 32'h41369041, 32'h420ee777};
test_input[12984:12991] = '{32'h41afc0e2, 32'hc25394d8, 32'hc283c430, 32'h40a7664e, 32'hc210ae1a, 32'h425dbd09, 32'h417bee93, 32'hc0a5b737};
test_output[12984:12991] = '{32'h41afc0e2, 32'h0, 32'h0, 32'h40a7664e, 32'h0, 32'h425dbd09, 32'h417bee93, 32'h0};
test_input[12992:12999] = '{32'hc2400d6a, 32'hc2c36f31, 32'h42829a83, 32'h4287b2e0, 32'hc292dee2, 32'hc20e1a11, 32'h41029753, 32'h416419ff};
test_output[12992:12999] = '{32'h0, 32'h0, 32'h42829a83, 32'h4287b2e0, 32'h0, 32'h0, 32'h41029753, 32'h416419ff};
test_input[13000:13007] = '{32'hc27a0877, 32'h4280478f, 32'h4038e71b, 32'hc0b77957, 32'hc1cc1663, 32'hc2133605, 32'hc2908b74, 32'h42620b7f};
test_output[13000:13007] = '{32'h0, 32'h4280478f, 32'h4038e71b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42620b7f};
test_input[13008:13015] = '{32'h4275ef08, 32'hc1e9e839, 32'h4150f6cb, 32'hc126d9e3, 32'h4289baf6, 32'h42551393, 32'hc187f8f6, 32'h41b16992};
test_output[13008:13015] = '{32'h4275ef08, 32'h0, 32'h4150f6cb, 32'h0, 32'h4289baf6, 32'h42551393, 32'h0, 32'h41b16992};
test_input[13016:13023] = '{32'hc27fe8e9, 32'hc211d642, 32'h4208609a, 32'hc20b3ada, 32'h428d561a, 32'hc2203db9, 32'h42956eac, 32'hc24e0863};
test_output[13016:13023] = '{32'h0, 32'h0, 32'h4208609a, 32'h0, 32'h428d561a, 32'h0, 32'h42956eac, 32'h0};
test_input[13024:13031] = '{32'hc1fa2bbb, 32'hc1cc9a6b, 32'hc2bc7e35, 32'h42a02a80, 32'h42a8baed, 32'h415ba61c, 32'hc1e5ede6, 32'h42b03f89};
test_output[13024:13031] = '{32'h0, 32'h0, 32'h0, 32'h42a02a80, 32'h42a8baed, 32'h415ba61c, 32'h0, 32'h42b03f89};
test_input[13032:13039] = '{32'h42ba4472, 32'hc1dc94fa, 32'h4172421c, 32'h428b710b, 32'h42140e6a, 32'h42c5ed92, 32'h42a88de9, 32'h41b966e1};
test_output[13032:13039] = '{32'h42ba4472, 32'h0, 32'h4172421c, 32'h428b710b, 32'h42140e6a, 32'h42c5ed92, 32'h42a88de9, 32'h41b966e1};
test_input[13040:13047] = '{32'hc2217556, 32'h429e20a4, 32'hc28cc15c, 32'h42a2caa9, 32'h42644844, 32'hc06e7d77, 32'h42c10c66, 32'h42beb692};
test_output[13040:13047] = '{32'h0, 32'h429e20a4, 32'h0, 32'h42a2caa9, 32'h42644844, 32'h0, 32'h42c10c66, 32'h42beb692};
test_input[13048:13055] = '{32'hc2840e94, 32'h41a1204c, 32'h41e93864, 32'hc1a22173, 32'hc1b95750, 32'h42878ec3, 32'hc16c0743, 32'hc27ba162};
test_output[13048:13055] = '{32'h0, 32'h41a1204c, 32'h41e93864, 32'h0, 32'h0, 32'h42878ec3, 32'h0, 32'h0};
test_input[13056:13063] = '{32'hc215b91c, 32'hc1098792, 32'h4294330d, 32'hc24c42a0, 32'h4158871c, 32'hc1af9890, 32'h42a6c34b, 32'hc25c15d8};
test_output[13056:13063] = '{32'h0, 32'h0, 32'h4294330d, 32'h0, 32'h4158871c, 32'h0, 32'h42a6c34b, 32'h0};
test_input[13064:13071] = '{32'h428e6dd2, 32'h41ae4b1d, 32'h41f08bc8, 32'hc17f4b4a, 32'h4237fa10, 32'hc2acc3c5, 32'hc10b3546, 32'h4195118a};
test_output[13064:13071] = '{32'h428e6dd2, 32'h41ae4b1d, 32'h41f08bc8, 32'h0, 32'h4237fa10, 32'h0, 32'h0, 32'h4195118a};
test_input[13072:13079] = '{32'h425aeab3, 32'hc2a17bb6, 32'hc1abc0f3, 32'hc2b22aa5, 32'h42af41d7, 32'hc2c3de2e, 32'hc1f08da0, 32'hbfa9fdc2};
test_output[13072:13079] = '{32'h425aeab3, 32'h0, 32'h0, 32'h0, 32'h42af41d7, 32'h0, 32'h0, 32'h0};
test_input[13080:13087] = '{32'hc1fdd7e7, 32'hc20d0c65, 32'hc2089a8e, 32'hc25eb7a8, 32'h4208c778, 32'h41bce0b8, 32'hbfd038e6, 32'h423b2332};
test_output[13080:13087] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4208c778, 32'h41bce0b8, 32'h0, 32'h423b2332};
test_input[13088:13095] = '{32'h42ab06a9, 32'h4250aaed, 32'hc29e5f34, 32'hc288ee6f, 32'hc26521a8, 32'h42806037, 32'hc235a9df, 32'h425e98ce};
test_output[13088:13095] = '{32'h42ab06a9, 32'h4250aaed, 32'h0, 32'h0, 32'h0, 32'h42806037, 32'h0, 32'h425e98ce};
test_input[13096:13103] = '{32'h42c7f300, 32'h421254c7, 32'hc2862ec8, 32'hc283c897, 32'h42293f28, 32'h41b8f82e, 32'h4184263f, 32'h42a5325d};
test_output[13096:13103] = '{32'h42c7f300, 32'h421254c7, 32'h0, 32'h0, 32'h42293f28, 32'h41b8f82e, 32'h4184263f, 32'h42a5325d};
test_input[13104:13111] = '{32'h41c91ef2, 32'h422ea578, 32'h42178b06, 32'h425f6c4c, 32'h4279b59e, 32'hc2874292, 32'hc1d2803e, 32'h4298b8bc};
test_output[13104:13111] = '{32'h41c91ef2, 32'h422ea578, 32'h42178b06, 32'h425f6c4c, 32'h4279b59e, 32'h0, 32'h0, 32'h4298b8bc};
test_input[13112:13119] = '{32'h4267188a, 32'hc2c76ec7, 32'hc2af9d2e, 32'hc2a3ce9a, 32'h41c3327b, 32'hc24f835c, 32'h42c59bd4, 32'hc2940803};
test_output[13112:13119] = '{32'h4267188a, 32'h0, 32'h0, 32'h0, 32'h41c3327b, 32'h0, 32'h42c59bd4, 32'h0};
test_input[13120:13127] = '{32'hc21cf30e, 32'hc0a4f40f, 32'h42aacdc4, 32'h4221e3db, 32'h421a9d53, 32'hc16f0402, 32'hc02f3c5c, 32'h428021b3};
test_output[13120:13127] = '{32'h0, 32'h0, 32'h42aacdc4, 32'h4221e3db, 32'h421a9d53, 32'h0, 32'h0, 32'h428021b3};
test_input[13128:13135] = '{32'h428dc3eb, 32'hc251afc0, 32'h42a6f901, 32'hc23a8882, 32'h428162f9, 32'h427aad1d, 32'h42b45a2f, 32'hc22bdb10};
test_output[13128:13135] = '{32'h428dc3eb, 32'h0, 32'h42a6f901, 32'h0, 32'h428162f9, 32'h427aad1d, 32'h42b45a2f, 32'h0};
test_input[13136:13143] = '{32'h4285c2f3, 32'h41dd986e, 32'h41fd7eb2, 32'hc121fcd7, 32'hc14112a9, 32'h41e295aa, 32'hc2224acc, 32'hc23c85a4};
test_output[13136:13143] = '{32'h4285c2f3, 32'h41dd986e, 32'h41fd7eb2, 32'h0, 32'h0, 32'h41e295aa, 32'h0, 32'h0};
test_input[13144:13151] = '{32'h42c5a4d3, 32'h42b8bb8c, 32'hc291b2f7, 32'h423ba27a, 32'h412299ac, 32'hc28cd514, 32'h414e7096, 32'hc208f4e2};
test_output[13144:13151] = '{32'h42c5a4d3, 32'h42b8bb8c, 32'h0, 32'h423ba27a, 32'h412299ac, 32'h0, 32'h414e7096, 32'h0};
test_input[13152:13159] = '{32'hc123c377, 32'hc0895c49, 32'hc12856f3, 32'h41f2233e, 32'h418cb68e, 32'hc204445b, 32'h40e29471, 32'h42bbf861};
test_output[13152:13159] = '{32'h0, 32'h0, 32'h0, 32'h41f2233e, 32'h418cb68e, 32'h0, 32'h40e29471, 32'h42bbf861};
test_input[13160:13167] = '{32'hc29e7c81, 32'hc2bb7cef, 32'hc295819d, 32'h4203e73e, 32'h42677cc6, 32'hc2796583, 32'hc2ba5229, 32'h424a690e};
test_output[13160:13167] = '{32'h0, 32'h0, 32'h0, 32'h4203e73e, 32'h42677cc6, 32'h0, 32'h0, 32'h424a690e};
test_input[13168:13175] = '{32'h41d03b34, 32'hc2991741, 32'hc279a3ed, 32'h42962f1a, 32'h424c7f79, 32'h41f32d17, 32'hc28cea88, 32'h42b9c4b0};
test_output[13168:13175] = '{32'h41d03b34, 32'h0, 32'h0, 32'h42962f1a, 32'h424c7f79, 32'h41f32d17, 32'h0, 32'h42b9c4b0};
test_input[13176:13183] = '{32'h41d6d127, 32'h429bd9c3, 32'hc1162d65, 32'h42310388, 32'hc1c11627, 32'h41cff107, 32'h41a00a7c, 32'h4242f75e};
test_output[13176:13183] = '{32'h41d6d127, 32'h429bd9c3, 32'h0, 32'h42310388, 32'h0, 32'h41cff107, 32'h41a00a7c, 32'h4242f75e};
test_input[13184:13191] = '{32'h42b30d30, 32'hc28cc351, 32'h3f8da3a5, 32'hc2341c69, 32'h420fa406, 32'hc2849f56, 32'h41ac8d1a, 32'h425d2f8a};
test_output[13184:13191] = '{32'h42b30d30, 32'h0, 32'h3f8da3a5, 32'h0, 32'h420fa406, 32'h0, 32'h41ac8d1a, 32'h425d2f8a};
test_input[13192:13199] = '{32'hc09d210d, 32'h42bfd076, 32'h4231abea, 32'h4216b007, 32'hc266642e, 32'h42a38748, 32'h428caccf, 32'hc2601b66};
test_output[13192:13199] = '{32'h0, 32'h42bfd076, 32'h4231abea, 32'h4216b007, 32'h0, 32'h42a38748, 32'h428caccf, 32'h0};
test_input[13200:13207] = '{32'hc2b75643, 32'hc1a19c31, 32'h42c5e1e7, 32'hc293f980, 32'h42a13403, 32'hc1dcd223, 32'h4265bec1, 32'hc2c0c2af};
test_output[13200:13207] = '{32'h0, 32'h0, 32'h42c5e1e7, 32'h0, 32'h42a13403, 32'h0, 32'h4265bec1, 32'h0};
test_input[13208:13215] = '{32'h4250f9e8, 32'h41a92e16, 32'hc28daa86, 32'h41af45fc, 32'h41fc82a5, 32'hc202218e, 32'hc1973ee3, 32'h42c4541a};
test_output[13208:13215] = '{32'h4250f9e8, 32'h41a92e16, 32'h0, 32'h41af45fc, 32'h41fc82a5, 32'h0, 32'h0, 32'h42c4541a};
test_input[13216:13223] = '{32'h42a176d2, 32'hc2c59b35, 32'h409f9052, 32'hc288b6dd, 32'h425f52af, 32'hc2538a1b, 32'hc1d9a7f6, 32'hc15b8f6c};
test_output[13216:13223] = '{32'h42a176d2, 32'h0, 32'h409f9052, 32'h0, 32'h425f52af, 32'h0, 32'h0, 32'h0};
test_input[13224:13231] = '{32'hc2958744, 32'hc08c42d4, 32'h42220320, 32'hc27f797d, 32'hc2c148f5, 32'h4219d17f, 32'hc24db219, 32'h42146d21};
test_output[13224:13231] = '{32'h0, 32'h0, 32'h42220320, 32'h0, 32'h0, 32'h4219d17f, 32'h0, 32'h42146d21};
test_input[13232:13239] = '{32'h428f91bb, 32'hc221d708, 32'h42a9468a, 32'hc28a9b3b, 32'h42c060f8, 32'h42889a32, 32'h42a4f70d, 32'h41cb9e1a};
test_output[13232:13239] = '{32'h428f91bb, 32'h0, 32'h42a9468a, 32'h0, 32'h42c060f8, 32'h42889a32, 32'h42a4f70d, 32'h41cb9e1a};
test_input[13240:13247] = '{32'hc1c28602, 32'hc262dac1, 32'h4198818c, 32'h42bf2310, 32'hc240b10e, 32'h40107070, 32'h422281e5, 32'h426110d2};
test_output[13240:13247] = '{32'h0, 32'h0, 32'h4198818c, 32'h42bf2310, 32'h0, 32'h40107070, 32'h422281e5, 32'h426110d2};
test_input[13248:13255] = '{32'hc2a513d0, 32'h417efde0, 32'h42279deb, 32'hc2c1dc70, 32'hc21b8788, 32'hc1c5407f, 32'hc2bd1750, 32'h424754ae};
test_output[13248:13255] = '{32'h0, 32'h417efde0, 32'h42279deb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h424754ae};
test_input[13256:13263] = '{32'h3f86485e, 32'h41083b30, 32'h428af40e, 32'h423ab0cc, 32'hc2547304, 32'h425817c9, 32'h4262f479, 32'hc1f2aa2a};
test_output[13256:13263] = '{32'h3f86485e, 32'h41083b30, 32'h428af40e, 32'h423ab0cc, 32'h0, 32'h425817c9, 32'h4262f479, 32'h0};
test_input[13264:13271] = '{32'h42aca24c, 32'hc18d0c93, 32'h4204325a, 32'hc17fbcd0, 32'h42b79237, 32'hc23ca0cd, 32'hc2664332, 32'hc18f972a};
test_output[13264:13271] = '{32'h42aca24c, 32'h0, 32'h4204325a, 32'h0, 32'h42b79237, 32'h0, 32'h0, 32'h0};
test_input[13272:13279] = '{32'hc262e6df, 32'h42b2fa85, 32'hc29d2738, 32'hc2c7bc9d, 32'hbe16f0c4, 32'h422d2642, 32'hc2438552, 32'h4119d8cc};
test_output[13272:13279] = '{32'h0, 32'h42b2fa85, 32'h0, 32'h0, 32'h0, 32'h422d2642, 32'h0, 32'h4119d8cc};
test_input[13280:13287] = '{32'h4140ef67, 32'h4195b2c2, 32'h41ed77e5, 32'h4285f548, 32'hc295bee0, 32'h42acb351, 32'h42996b2d, 32'h424ef6a0};
test_output[13280:13287] = '{32'h4140ef67, 32'h4195b2c2, 32'h41ed77e5, 32'h4285f548, 32'h0, 32'h42acb351, 32'h42996b2d, 32'h424ef6a0};
test_input[13288:13295] = '{32'h4290b099, 32'hc287ff89, 32'h42a0a334, 32'hc29592d7, 32'h4261cc12, 32'hc28ee04f, 32'hc29ee381, 32'hc1bd7541};
test_output[13288:13295] = '{32'h4290b099, 32'h0, 32'h42a0a334, 32'h0, 32'h4261cc12, 32'h0, 32'h0, 32'h0};
test_input[13296:13303] = '{32'hc286b984, 32'h41cbf965, 32'hc2b75832, 32'hc28ba60c, 32'hc297393f, 32'h40eab1e0, 32'h4284318b, 32'h40d9ef22};
test_output[13296:13303] = '{32'h0, 32'h41cbf965, 32'h0, 32'h0, 32'h0, 32'h40eab1e0, 32'h4284318b, 32'h40d9ef22};
test_input[13304:13311] = '{32'h41c3486f, 32'h429b382e, 32'hc2538707, 32'h42bcb807, 32'hc226ebf2, 32'hc25ebd18, 32'h410c97b9, 32'hc23d6cb3};
test_output[13304:13311] = '{32'h41c3486f, 32'h429b382e, 32'h0, 32'h42bcb807, 32'h0, 32'h0, 32'h410c97b9, 32'h0};
test_input[13312:13319] = '{32'h41c930b0, 32'h428b59c2, 32'hbfd4628e, 32'hc297b1de, 32'h420e6c25, 32'hc23d1895, 32'h421a2d32, 32'hc2aa77d5};
test_output[13312:13319] = '{32'h41c930b0, 32'h428b59c2, 32'h0, 32'h0, 32'h420e6c25, 32'h0, 32'h421a2d32, 32'h0};
test_input[13320:13327] = '{32'hc2ad3346, 32'hc2b00901, 32'h4280084d, 32'h41ffcaff, 32'h42524b8f, 32'hc28973a8, 32'h422563fa, 32'hc1ee2cee};
test_output[13320:13327] = '{32'h0, 32'h0, 32'h4280084d, 32'h41ffcaff, 32'h42524b8f, 32'h0, 32'h422563fa, 32'h0};
test_input[13328:13335] = '{32'h42944608, 32'hc276e504, 32'hc2a4a67d, 32'hc2993c87, 32'hc2ac99e2, 32'h42c2eae5, 32'h41843494, 32'hc184767b};
test_output[13328:13335] = '{32'h42944608, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c2eae5, 32'h41843494, 32'h0};
test_input[13336:13343] = '{32'h40ef7dec, 32'h423eb5bd, 32'h41f630ca, 32'hc2bf3921, 32'h42b90569, 32'hc1fc58e9, 32'hc21e66e9, 32'h421507ce};
test_output[13336:13343] = '{32'h40ef7dec, 32'h423eb5bd, 32'h41f630ca, 32'h0, 32'h42b90569, 32'h0, 32'h0, 32'h421507ce};
test_input[13344:13351] = '{32'hc18c9b7e, 32'hc13f79a1, 32'h4261b0e5, 32'h4291c36c, 32'h42690e90, 32'hc2809d57, 32'h42689ae9, 32'h411b1a18};
test_output[13344:13351] = '{32'h0, 32'h0, 32'h4261b0e5, 32'h4291c36c, 32'h42690e90, 32'h0, 32'h42689ae9, 32'h411b1a18};
test_input[13352:13359] = '{32'hc1629a50, 32'hc191c666, 32'hc1ad3901, 32'h42988c45, 32'h413b8f98, 32'h425f2541, 32'h41a1f628, 32'h42bd4b8f};
test_output[13352:13359] = '{32'h0, 32'h0, 32'h0, 32'h42988c45, 32'h413b8f98, 32'h425f2541, 32'h41a1f628, 32'h42bd4b8f};
test_input[13360:13367] = '{32'hc13a6454, 32'hc21148c8, 32'hc0e1d0cb, 32'hc2862750, 32'h4276476e, 32'hc22381a3, 32'hc25b4b77, 32'h42b7a587};
test_output[13360:13367] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4276476e, 32'h0, 32'h0, 32'h42b7a587};
test_input[13368:13375] = '{32'hc28ab12d, 32'h42a255d0, 32'hc1e48e35, 32'h417d936a, 32'hc0bf7dae, 32'h4211fe64, 32'h424784fd, 32'h41f6e2db};
test_output[13368:13375] = '{32'h0, 32'h42a255d0, 32'h0, 32'h417d936a, 32'h0, 32'h4211fe64, 32'h424784fd, 32'h41f6e2db};
test_input[13376:13383] = '{32'hc1d19313, 32'h42b15822, 32'h412b7a66, 32'h41553c7f, 32'hc236e4f9, 32'hc18a2ea9, 32'h428f4a6f, 32'h428c52fe};
test_output[13376:13383] = '{32'h0, 32'h42b15822, 32'h412b7a66, 32'h41553c7f, 32'h0, 32'h0, 32'h428f4a6f, 32'h428c52fe};
test_input[13384:13391] = '{32'h4281e2d5, 32'h4230316d, 32'h42b4f932, 32'h4228bd39, 32'h40145109, 32'hc2ad2f45, 32'hc1bd8175, 32'hc246fa1e};
test_output[13384:13391] = '{32'h4281e2d5, 32'h4230316d, 32'h42b4f932, 32'h4228bd39, 32'h40145109, 32'h0, 32'h0, 32'h0};
test_input[13392:13399] = '{32'h42aec1d2, 32'h42481c43, 32'hc282d4c1, 32'h4231610f, 32'h4295181e, 32'hc2285f3e, 32'h42c6b66e, 32'h42ba5ba2};
test_output[13392:13399] = '{32'h42aec1d2, 32'h42481c43, 32'h0, 32'h4231610f, 32'h4295181e, 32'h0, 32'h42c6b66e, 32'h42ba5ba2};
test_input[13400:13407] = '{32'hc2853c08, 32'h42a2d28a, 32'h420d2817, 32'h42965f25, 32'h41a6c37a, 32'h41e5387a, 32'hc189651d, 32'hc226a12f};
test_output[13400:13407] = '{32'h0, 32'h42a2d28a, 32'h420d2817, 32'h42965f25, 32'h41a6c37a, 32'h41e5387a, 32'h0, 32'h0};
test_input[13408:13415] = '{32'h4279cd01, 32'hc2823b31, 32'h42376551, 32'hc2c4baab, 32'h42a6ad20, 32'hc281d6db, 32'hc1895df1, 32'hc1dab9d5};
test_output[13408:13415] = '{32'h4279cd01, 32'h0, 32'h42376551, 32'h0, 32'h42a6ad20, 32'h0, 32'h0, 32'h0};
test_input[13416:13423] = '{32'h4148ad04, 32'hc15d947a, 32'hc2c5d9a1, 32'h41df8270, 32'h42200313, 32'hc0affaab, 32'h4248fc90, 32'hc2c0e3d0};
test_output[13416:13423] = '{32'h4148ad04, 32'h0, 32'h0, 32'h41df8270, 32'h42200313, 32'h0, 32'h4248fc90, 32'h0};
test_input[13424:13431] = '{32'hc193c891, 32'h4285a13a, 32'hc274cf21, 32'hc1881f71, 32'hbf01445f, 32'hc2c0b0c7, 32'hc206ca02, 32'hc2bf9a1e};
test_output[13424:13431] = '{32'h0, 32'h4285a13a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13432:13439] = '{32'hc29bf09f, 32'h41f19892, 32'h428c5f70, 32'hc28aef90, 32'hc2c6a4bf, 32'h42bffa6e, 32'h4216871f, 32'hc2248705};
test_output[13432:13439] = '{32'h0, 32'h41f19892, 32'h428c5f70, 32'h0, 32'h0, 32'h42bffa6e, 32'h4216871f, 32'h0};
test_input[13440:13447] = '{32'h42b01089, 32'h42015510, 32'h428cb709, 32'hc2340af0, 32'h42af852a, 32'hc22a5dc2, 32'h42080f73, 32'hc22cd81c};
test_output[13440:13447] = '{32'h42b01089, 32'h42015510, 32'h428cb709, 32'h0, 32'h42af852a, 32'h0, 32'h42080f73, 32'h0};
test_input[13448:13455] = '{32'h42a70495, 32'hc1cd1efc, 32'hc1eaf330, 32'h424cfecc, 32'h415318a9, 32'h41d9cb25, 32'hc2b5195f, 32'h42c4b87a};
test_output[13448:13455] = '{32'h42a70495, 32'h0, 32'h0, 32'h424cfecc, 32'h415318a9, 32'h41d9cb25, 32'h0, 32'h42c4b87a};
test_input[13456:13463] = '{32'h4134dcd4, 32'hc2557e00, 32'h42125fc9, 32'h420bab7f, 32'hc08b88de, 32'h428e0044, 32'h41def922, 32'h420f0bcf};
test_output[13456:13463] = '{32'h4134dcd4, 32'h0, 32'h42125fc9, 32'h420bab7f, 32'h0, 32'h428e0044, 32'h41def922, 32'h420f0bcf};
test_input[13464:13471] = '{32'h3f7ea9a2, 32'h42517c4c, 32'h42729335, 32'hc279c53e, 32'hc1b770e8, 32'hc13ba0b2, 32'h42c69f01, 32'hc2306e9f};
test_output[13464:13471] = '{32'h3f7ea9a2, 32'h42517c4c, 32'h42729335, 32'h0, 32'h0, 32'h0, 32'h42c69f01, 32'h0};
test_input[13472:13479] = '{32'hc292ea85, 32'hc2434a1a, 32'hc09c20e7, 32'h429148a2, 32'h420268f8, 32'h41a21b60, 32'hc1617f12, 32'h41afe2da};
test_output[13472:13479] = '{32'h0, 32'h0, 32'h0, 32'h429148a2, 32'h420268f8, 32'h41a21b60, 32'h0, 32'h41afe2da};
test_input[13480:13487] = '{32'h42621f6a, 32'hc1831607, 32'h42b66d86, 32'h41eba1be, 32'hc21fa51c, 32'h42ac2e89, 32'h40b39ab7, 32'h4274024b};
test_output[13480:13487] = '{32'h42621f6a, 32'h0, 32'h42b66d86, 32'h41eba1be, 32'h0, 32'h42ac2e89, 32'h40b39ab7, 32'h4274024b};
test_input[13488:13495] = '{32'hc234e8f9, 32'h424207e5, 32'hc291198d, 32'hc2c41f0b, 32'hc14569df, 32'hc2a87022, 32'h420837b8, 32'h41bba91e};
test_output[13488:13495] = '{32'h0, 32'h424207e5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420837b8, 32'h41bba91e};
test_input[13496:13503] = '{32'h4283c5bb, 32'h42ae1476, 32'h41ee17a8, 32'h42b3c724, 32'hc2847265, 32'h42aaef35, 32'hc297023b, 32'hc19ec6d1};
test_output[13496:13503] = '{32'h4283c5bb, 32'h42ae1476, 32'h41ee17a8, 32'h42b3c724, 32'h0, 32'h42aaef35, 32'h0, 32'h0};
test_input[13504:13511] = '{32'hc2033312, 32'h427645b1, 32'h42510beb, 32'hc2b4ca62, 32'h427930a2, 32'h4066a7ef, 32'hc2ba2699, 32'hc1ef8b0d};
test_output[13504:13511] = '{32'h0, 32'h427645b1, 32'h42510beb, 32'h0, 32'h427930a2, 32'h4066a7ef, 32'h0, 32'h0};
test_input[13512:13519] = '{32'hc2b8c908, 32'hc2879a0a, 32'hc21e882c, 32'hc256d8a9, 32'h428d5d3c, 32'h42b8ecc2, 32'hc26519bd, 32'hc117d2a2};
test_output[13512:13519] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h428d5d3c, 32'h42b8ecc2, 32'h0, 32'h0};
test_input[13520:13527] = '{32'h41e4f8f0, 32'hc182cb7a, 32'h42828cb8, 32'h41835b64, 32'hc206ea11, 32'hc2239c7e, 32'h40d3f130, 32'h41fa28af};
test_output[13520:13527] = '{32'h41e4f8f0, 32'h0, 32'h42828cb8, 32'h41835b64, 32'h0, 32'h0, 32'h40d3f130, 32'h41fa28af};
test_input[13528:13535] = '{32'hc29139a9, 32'hc20bec72, 32'h41980208, 32'hc1ec24cb, 32'h4189980b, 32'hc21d4e2a, 32'hc22bcd12, 32'hc1a640cf};
test_output[13528:13535] = '{32'h0, 32'h0, 32'h41980208, 32'h0, 32'h4189980b, 32'h0, 32'h0, 32'h0};
test_input[13536:13543] = '{32'h425f6dbb, 32'hbecc7a8a, 32'h424459c6, 32'h41c2dd45, 32'hc297b03c, 32'hc1e6b8b7, 32'hc1c97ba7, 32'hc1229ff3};
test_output[13536:13543] = '{32'h425f6dbb, 32'h0, 32'h424459c6, 32'h41c2dd45, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13544:13551] = '{32'hc1056b39, 32'hc0d701d5, 32'hc29b8339, 32'hbeebdbfc, 32'hc1e7b956, 32'h41b4cf73, 32'h420f893c, 32'hc1c2ab27};
test_output[13544:13551] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b4cf73, 32'h420f893c, 32'h0};
test_input[13552:13559] = '{32'h3f4f56f4, 32'h427bd0b2, 32'hc2a5673f, 32'hc2c46f97, 32'hc1e9b629, 32'hc2140a32, 32'hc2905bb9, 32'h4236bc35};
test_output[13552:13559] = '{32'h3f4f56f4, 32'h427bd0b2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4236bc35};
test_input[13560:13567] = '{32'hc21d2745, 32'h4287fb12, 32'h42c1826b, 32'h41a2656b, 32'hc2c11127, 32'h4196061c, 32'hc2324088, 32'hc224e74d};
test_output[13560:13567] = '{32'h0, 32'h4287fb12, 32'h42c1826b, 32'h41a2656b, 32'h0, 32'h4196061c, 32'h0, 32'h0};
test_input[13568:13575] = '{32'hc28f7808, 32'h41428266, 32'h41bfc7fc, 32'h42b8f91f, 32'h4183bdd5, 32'hc19e1dfc, 32'hc20464c5, 32'h42098ce2};
test_output[13568:13575] = '{32'h0, 32'h41428266, 32'h41bfc7fc, 32'h42b8f91f, 32'h4183bdd5, 32'h0, 32'h0, 32'h42098ce2};
test_input[13576:13583] = '{32'hc1809033, 32'h428b904b, 32'hc0c02e26, 32'hc2592234, 32'h4133306d, 32'hc2c441be, 32'h41109a2a, 32'h419f6b39};
test_output[13576:13583] = '{32'h0, 32'h428b904b, 32'h0, 32'h0, 32'h4133306d, 32'h0, 32'h41109a2a, 32'h419f6b39};
test_input[13584:13591] = '{32'hc29adb29, 32'hc1a6a7b9, 32'h42aae123, 32'hc2c6338f, 32'h429e4b53, 32'h429ad237, 32'h42a5e196, 32'h42282f2f};
test_output[13584:13591] = '{32'h0, 32'h0, 32'h42aae123, 32'h0, 32'h429e4b53, 32'h429ad237, 32'h42a5e196, 32'h42282f2f};
test_input[13592:13599] = '{32'h4243fb45, 32'hc1bc0cb0, 32'hc28c346c, 32'h42961e64, 32'h42890d72, 32'hc2005799, 32'h400a0d90, 32'h42af3fc6};
test_output[13592:13599] = '{32'h4243fb45, 32'h0, 32'h0, 32'h42961e64, 32'h42890d72, 32'h0, 32'h400a0d90, 32'h42af3fc6};
test_input[13600:13607] = '{32'h40f64491, 32'h4194732f, 32'h41f8dc19, 32'h426269d8, 32'h4209b8ca, 32'hc26be0da, 32'hc21112c1, 32'hc1ea1285};
test_output[13600:13607] = '{32'h40f64491, 32'h4194732f, 32'h41f8dc19, 32'h426269d8, 32'h4209b8ca, 32'h0, 32'h0, 32'h0};
test_input[13608:13615] = '{32'hc231fb2a, 32'hc23a02c2, 32'hc1720fc5, 32'hc287fe6f, 32'h40c7c391, 32'h42bfddf8, 32'h41d198e6, 32'hc1ecacb4};
test_output[13608:13615] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40c7c391, 32'h42bfddf8, 32'h41d198e6, 32'h0};
test_input[13616:13623] = '{32'h429178a7, 32'h42b57fa4, 32'h3eb57081, 32'h412dde23, 32'h425955a6, 32'hc2553b7a, 32'hc20a4ce7, 32'hc1d323ee};
test_output[13616:13623] = '{32'h429178a7, 32'h42b57fa4, 32'h3eb57081, 32'h412dde23, 32'h425955a6, 32'h0, 32'h0, 32'h0};
test_input[13624:13631] = '{32'hc23913ed, 32'h41669d49, 32'h4066bf5d, 32'hc0b22eee, 32'h42aec3e3, 32'h422e3a47, 32'h42bcae0d, 32'h41830b8f};
test_output[13624:13631] = '{32'h0, 32'h41669d49, 32'h4066bf5d, 32'h0, 32'h42aec3e3, 32'h422e3a47, 32'h42bcae0d, 32'h41830b8f};
test_input[13632:13639] = '{32'hc272da39, 32'hc2a10e19, 32'hc2c220d8, 32'hc116233b, 32'hc24f4a8b, 32'hc18d83b1, 32'h4226ae2a, 32'hc212d7a9};
test_output[13632:13639] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4226ae2a, 32'h0};
test_input[13640:13647] = '{32'h41ba1be2, 32'hc28c68ef, 32'h41fd380d, 32'hc2960fef, 32'hc195ad1b, 32'h425a0821, 32'hc255ecdd, 32'hc22ca6f7};
test_output[13640:13647] = '{32'h41ba1be2, 32'h0, 32'h41fd380d, 32'h0, 32'h0, 32'h425a0821, 32'h0, 32'h0};
test_input[13648:13655] = '{32'hc24c5be3, 32'hc1acff96, 32'hc25020ff, 32'hc2a17878, 32'hc285464e, 32'h41a938f0, 32'h428716b9, 32'hc21dbeae};
test_output[13648:13655] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41a938f0, 32'h428716b9, 32'h0};
test_input[13656:13663] = '{32'hc2b897eb, 32'h42bb80b6, 32'hc174f257, 32'hc1573cb8, 32'h42b4a153, 32'h420422b7, 32'hc21c3a25, 32'h42c3bdd1};
test_output[13656:13663] = '{32'h0, 32'h42bb80b6, 32'h0, 32'h0, 32'h42b4a153, 32'h420422b7, 32'h0, 32'h42c3bdd1};
test_input[13664:13671] = '{32'hc1e8accd, 32'hc2c10a66, 32'h42944fd1, 32'h4257bf98, 32'h42831522, 32'h4296ad07, 32'hc2a66bb2, 32'hc21c5f95};
test_output[13664:13671] = '{32'h0, 32'h0, 32'h42944fd1, 32'h4257bf98, 32'h42831522, 32'h4296ad07, 32'h0, 32'h0};
test_input[13672:13679] = '{32'hc29ac4b7, 32'h42aeca66, 32'h40714202, 32'h41601847, 32'hc2959f69, 32'h42b7a3e1, 32'h403bd5eb, 32'h424ead03};
test_output[13672:13679] = '{32'h0, 32'h42aeca66, 32'h40714202, 32'h41601847, 32'h0, 32'h42b7a3e1, 32'h403bd5eb, 32'h424ead03};
test_input[13680:13687] = '{32'hc2c2a882, 32'h4285d35a, 32'h42b258c1, 32'h42af72ff, 32'h418dc859, 32'h42981ce0, 32'h424b52c5, 32'h4291355d};
test_output[13680:13687] = '{32'h0, 32'h4285d35a, 32'h42b258c1, 32'h42af72ff, 32'h418dc859, 32'h42981ce0, 32'h424b52c5, 32'h4291355d};
test_input[13688:13695] = '{32'h424a566b, 32'h42ade819, 32'h4297a191, 32'h426f788f, 32'hc27a050d, 32'h426e75f8, 32'hc15d6f88, 32'h4251c50f};
test_output[13688:13695] = '{32'h424a566b, 32'h42ade819, 32'h4297a191, 32'h426f788f, 32'h0, 32'h426e75f8, 32'h0, 32'h4251c50f};
test_input[13696:13703] = '{32'h427c2dc0, 32'h422473d1, 32'h415686c4, 32'hc1775f98, 32'h4246be53, 32'hc28b7574, 32'h42122bfa, 32'hc2b32a94};
test_output[13696:13703] = '{32'h427c2dc0, 32'h422473d1, 32'h415686c4, 32'h0, 32'h4246be53, 32'h0, 32'h42122bfa, 32'h0};
test_input[13704:13711] = '{32'h4242b68d, 32'hc2477293, 32'h4296ff54, 32'hc2003abf, 32'h423cc170, 32'h40ae5a00, 32'h42b04046, 32'h420a8e35};
test_output[13704:13711] = '{32'h4242b68d, 32'h0, 32'h4296ff54, 32'h0, 32'h423cc170, 32'h40ae5a00, 32'h42b04046, 32'h420a8e35};
test_input[13712:13719] = '{32'hc28516b8, 32'h42932f35, 32'hc2ab301e, 32'h41e81051, 32'h41235b9a, 32'h42812f5a, 32'h42c1cfaa, 32'hc2917381};
test_output[13712:13719] = '{32'h0, 32'h42932f35, 32'h0, 32'h41e81051, 32'h41235b9a, 32'h42812f5a, 32'h42c1cfaa, 32'h0};
test_input[13720:13727] = '{32'hc2b65149, 32'h4287ab8e, 32'h40c9f968, 32'h41dbb847, 32'hc2937609, 32'h42128942, 32'hc257e896, 32'h429c2f77};
test_output[13720:13727] = '{32'h0, 32'h4287ab8e, 32'h40c9f968, 32'h41dbb847, 32'h0, 32'h42128942, 32'h0, 32'h429c2f77};
test_input[13728:13735] = '{32'hc25d4503, 32'h409b07e1, 32'hc276a96f, 32'h420b707b, 32'hc2510c10, 32'hc27a768e, 32'h42575f4f, 32'hc2891f77};
test_output[13728:13735] = '{32'h0, 32'h409b07e1, 32'h0, 32'h420b707b, 32'h0, 32'h0, 32'h42575f4f, 32'h0};
test_input[13736:13743] = '{32'h42b2131f, 32'h424e5f17, 32'h4291eb3e, 32'hc2a07237, 32'hc2af4b8b, 32'hc1f0beea, 32'hc1e93f79, 32'hc20bbe31};
test_output[13736:13743] = '{32'h42b2131f, 32'h424e5f17, 32'h4291eb3e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13744:13751] = '{32'hc29119fe, 32'h428bc7da, 32'hc23146ed, 32'h419644ad, 32'h4111e85d, 32'hc225e232, 32'hc2a9ae7e, 32'h42afe485};
test_output[13744:13751] = '{32'h0, 32'h428bc7da, 32'h0, 32'h419644ad, 32'h4111e85d, 32'h0, 32'h0, 32'h42afe485};
test_input[13752:13759] = '{32'hc29e14d5, 32'hc2485817, 32'hc1c8786a, 32'hc2b0607e, 32'hc21a9109, 32'h42997f13, 32'hc1991b9a, 32'h41fce65d};
test_output[13752:13759] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42997f13, 32'h0, 32'h41fce65d};
test_input[13760:13767] = '{32'h420c139e, 32'h408a460c, 32'hc26ae6ee, 32'h425def80, 32'hc1b3f75e, 32'h429e17fe, 32'hc22ca7c6, 32'hc282efa2};
test_output[13760:13767] = '{32'h420c139e, 32'h408a460c, 32'h0, 32'h425def80, 32'h0, 32'h429e17fe, 32'h0, 32'h0};
test_input[13768:13775] = '{32'hc25e2492, 32'h41f976df, 32'hc21ec6fe, 32'h42c585db, 32'hc2964f1e, 32'hc28259a5, 32'h429a66a7, 32'h4291db68};
test_output[13768:13775] = '{32'h0, 32'h41f976df, 32'h0, 32'h42c585db, 32'h0, 32'h0, 32'h429a66a7, 32'h4291db68};
test_input[13776:13783] = '{32'h41a00889, 32'hc0975c1d, 32'h4223ba9e, 32'h4296ab28, 32'h412144c5, 32'h424f3752, 32'hc2bcc3f5, 32'h41d5494e};
test_output[13776:13783] = '{32'h41a00889, 32'h0, 32'h4223ba9e, 32'h4296ab28, 32'h412144c5, 32'h424f3752, 32'h0, 32'h41d5494e};
test_input[13784:13791] = '{32'hc28c04a8, 32'hc256283b, 32'h42b7c2ff, 32'hc1b5f753, 32'h41cc7350, 32'h41b6c52f, 32'hc1a3382b, 32'h416b51e3};
test_output[13784:13791] = '{32'h0, 32'h0, 32'h42b7c2ff, 32'h0, 32'h41cc7350, 32'h41b6c52f, 32'h0, 32'h416b51e3};
test_input[13792:13799] = '{32'h425bbe1c, 32'h3f20b7dd, 32'hc290958d, 32'hc2203a86, 32'hc2ac3c55, 32'h4285a73f, 32'h426e5c39, 32'h42b9c57d};
test_output[13792:13799] = '{32'h425bbe1c, 32'h3f20b7dd, 32'h0, 32'h0, 32'h0, 32'h4285a73f, 32'h426e5c39, 32'h42b9c57d};
test_input[13800:13807] = '{32'h42c0b21f, 32'hc24560ae, 32'hc1f4095f, 32'hc09a83c3, 32'h42b052cb, 32'hc2bd08ce, 32'h4294f211, 32'h421557c1};
test_output[13800:13807] = '{32'h42c0b21f, 32'h0, 32'h0, 32'h0, 32'h42b052cb, 32'h0, 32'h4294f211, 32'h421557c1};
test_input[13808:13815] = '{32'h41d45560, 32'h42433b08, 32'h42ad8221, 32'hc2c4a3a6, 32'h4274c28a, 32'hc29dde86, 32'h42986f04, 32'h412bfcd2};
test_output[13808:13815] = '{32'h41d45560, 32'h42433b08, 32'h42ad8221, 32'h0, 32'h4274c28a, 32'h0, 32'h42986f04, 32'h412bfcd2};
test_input[13816:13823] = '{32'hc285a35e, 32'hc27cdc22, 32'h408ffcd4, 32'h424e3f72, 32'hc28f5d19, 32'h428c2a03, 32'h42a2a6f6, 32'h424e1f12};
test_output[13816:13823] = '{32'h0, 32'h0, 32'h408ffcd4, 32'h424e3f72, 32'h0, 32'h428c2a03, 32'h42a2a6f6, 32'h424e1f12};
test_input[13824:13831] = '{32'hc2c70a05, 32'hc250eaeb, 32'h42034c74, 32'h4143c27d, 32'hc28c3bac, 32'hc0ad9b24, 32'h42bd9aaf, 32'h42af7717};
test_output[13824:13831] = '{32'h0, 32'h0, 32'h42034c74, 32'h4143c27d, 32'h0, 32'h0, 32'h42bd9aaf, 32'h42af7717};
test_input[13832:13839] = '{32'h42a108bc, 32'h4119058c, 32'h42c16c31, 32'hc0bb09ae, 32'hc2abec0f, 32'h42477789, 32'h41cb04c3, 32'h41ac575d};
test_output[13832:13839] = '{32'h42a108bc, 32'h4119058c, 32'h42c16c31, 32'h0, 32'h0, 32'h42477789, 32'h41cb04c3, 32'h41ac575d};
test_input[13840:13847] = '{32'hc2b27c62, 32'h4272e9a7, 32'h422351af, 32'h4285a1fa, 32'hc183e12d, 32'hc1753269, 32'hc29f6be8, 32'h4229c9c9};
test_output[13840:13847] = '{32'h0, 32'h4272e9a7, 32'h422351af, 32'h4285a1fa, 32'h0, 32'h0, 32'h0, 32'h4229c9c9};
test_input[13848:13855] = '{32'h4227416d, 32'hc2032027, 32'hc1e27cfa, 32'hc28cf3fd, 32'hc23b18ff, 32'hc2357506, 32'hc2a9fc05, 32'hc29012e3};
test_output[13848:13855] = '{32'h4227416d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13856:13863] = '{32'hc26c4d7a, 32'h426ee219, 32'h4161a54f, 32'hc2aaba90, 32'h41e897a8, 32'h4283d4df, 32'h42c2dda3, 32'h407b54a5};
test_output[13856:13863] = '{32'h0, 32'h426ee219, 32'h4161a54f, 32'h0, 32'h41e897a8, 32'h4283d4df, 32'h42c2dda3, 32'h407b54a5};
test_input[13864:13871] = '{32'hc27ee994, 32'hc2885278, 32'hc2435bb7, 32'hc28b7aa4, 32'h4266bb1c, 32'hc216f6de, 32'hc2b83e4b, 32'hc210ab5a};
test_output[13864:13871] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4266bb1c, 32'h0, 32'h0, 32'h0};
test_input[13872:13879] = '{32'hc279d8cd, 32'hc2892e76, 32'h42c64c7e, 32'h4276b794, 32'hc2024ce0, 32'h4299d0e5, 32'h425e6aac, 32'h42b939a6};
test_output[13872:13879] = '{32'h0, 32'h0, 32'h42c64c7e, 32'h4276b794, 32'h0, 32'h4299d0e5, 32'h425e6aac, 32'h42b939a6};
test_input[13880:13887] = '{32'hc269d22c, 32'hc1214c55, 32'h420c6fc0, 32'hc2a7cf17, 32'h4141c617, 32'hc0ad7ed2, 32'hc260f450, 32'h42a02e88};
test_output[13880:13887] = '{32'h0, 32'h0, 32'h420c6fc0, 32'h0, 32'h4141c617, 32'h0, 32'h0, 32'h42a02e88};
test_input[13888:13895] = '{32'hc28fb8f6, 32'hc24e03db, 32'h422d9cdb, 32'h41cdc52d, 32'h42435f44, 32'h420e9387, 32'hc29b459b, 32'h427328b5};
test_output[13888:13895] = '{32'h0, 32'h0, 32'h422d9cdb, 32'h41cdc52d, 32'h42435f44, 32'h420e9387, 32'h0, 32'h427328b5};
test_input[13896:13903] = '{32'hc18181b1, 32'hc1ab53b8, 32'hc1cd8ad0, 32'h41d044be, 32'hc24e2543, 32'h42b7ee1d, 32'h426e1649, 32'hc278383b};
test_output[13896:13903] = '{32'h0, 32'h0, 32'h0, 32'h41d044be, 32'h0, 32'h42b7ee1d, 32'h426e1649, 32'h0};
test_input[13904:13911] = '{32'hc1edc948, 32'h41854d8a, 32'hc2ae62a5, 32'h424c32f5, 32'hc1f21e9d, 32'h418f839f, 32'h42bc0ff0, 32'h41b52755};
test_output[13904:13911] = '{32'h0, 32'h41854d8a, 32'h0, 32'h424c32f5, 32'h0, 32'h418f839f, 32'h42bc0ff0, 32'h41b52755};
test_input[13912:13919] = '{32'hc2b6a280, 32'hc1f18765, 32'hc22d3369, 32'h41dc01bf, 32'h40577363, 32'hc24f7321, 32'hc25e690e, 32'h42abef8c};
test_output[13912:13919] = '{32'h0, 32'h0, 32'h0, 32'h41dc01bf, 32'h40577363, 32'h0, 32'h0, 32'h42abef8c};
test_input[13920:13927] = '{32'h42c0c35d, 32'h424e8a15, 32'hc22fd53b, 32'hc1d21d4c, 32'hbd7be5f7, 32'h42b89e05, 32'hc023ad9a, 32'h42818e51};
test_output[13920:13927] = '{32'h42c0c35d, 32'h424e8a15, 32'h0, 32'h0, 32'h0, 32'h42b89e05, 32'h0, 32'h42818e51};
test_input[13928:13935] = '{32'hc2c07e17, 32'h42ac0bdf, 32'hbee28737, 32'hc2a67a6e, 32'h4253fa5d, 32'h418fdc1d, 32'hc2c26b97, 32'h42bf539a};
test_output[13928:13935] = '{32'h0, 32'h42ac0bdf, 32'h0, 32'h0, 32'h4253fa5d, 32'h418fdc1d, 32'h0, 32'h42bf539a};
test_input[13936:13943] = '{32'hc2bbcabd, 32'hc0dbf10a, 32'h41e8418d, 32'hc18acce8, 32'h425a8d25, 32'hc28a01a2, 32'hc1c9b0aa, 32'hc244b66d};
test_output[13936:13943] = '{32'h0, 32'h0, 32'h41e8418d, 32'h0, 32'h425a8d25, 32'h0, 32'h0, 32'h0};
test_input[13944:13951] = '{32'h41ab98f2, 32'h421a8752, 32'h421e7d50, 32'h418e6c96, 32'hc0d4752e, 32'hc184b4a0, 32'hbf8113b3, 32'h42ad1769};
test_output[13944:13951] = '{32'h41ab98f2, 32'h421a8752, 32'h421e7d50, 32'h418e6c96, 32'h0, 32'h0, 32'h0, 32'h42ad1769};
test_input[13952:13959] = '{32'h4288243b, 32'hc29d66fd, 32'h42bf7432, 32'hc07bbc75, 32'hc112d463, 32'h42916411, 32'h41542fea, 32'hc144b2da};
test_output[13952:13959] = '{32'h4288243b, 32'h0, 32'h42bf7432, 32'h0, 32'h0, 32'h42916411, 32'h41542fea, 32'h0};
test_input[13960:13967] = '{32'h422b76b1, 32'h423c5112, 32'h42c46771, 32'h42434e69, 32'hc1c40f1f, 32'h4265db5f, 32'hc2035452, 32'h41d48f20};
test_output[13960:13967] = '{32'h422b76b1, 32'h423c5112, 32'h42c46771, 32'h42434e69, 32'h0, 32'h4265db5f, 32'h0, 32'h41d48f20};
test_input[13968:13975] = '{32'hc22e6af7, 32'h42ace286, 32'hc06fe4ea, 32'h42bfc27d, 32'h4291333d, 32'hc1f7c648, 32'hc2a836d8, 32'hc125452f};
test_output[13968:13975] = '{32'h0, 32'h42ace286, 32'h0, 32'h42bfc27d, 32'h4291333d, 32'h0, 32'h0, 32'h0};
test_input[13976:13983] = '{32'h4259b18f, 32'h4135aaf7, 32'hc2c28616, 32'h414e6f87, 32'h420c69e3, 32'hc2a486a1, 32'h4206635b, 32'h42bc9b7d};
test_output[13976:13983] = '{32'h4259b18f, 32'h4135aaf7, 32'h0, 32'h414e6f87, 32'h420c69e3, 32'h0, 32'h4206635b, 32'h42bc9b7d};
test_input[13984:13991] = '{32'h42a41edc, 32'h426bae5c, 32'h40d180e5, 32'hc274eb39, 32'hc2439748, 32'h40fcace3, 32'h42a79b95, 32'hc2371506};
test_output[13984:13991] = '{32'h42a41edc, 32'h426bae5c, 32'h40d180e5, 32'h0, 32'h0, 32'h40fcace3, 32'h42a79b95, 32'h0};
test_input[13992:13999] = '{32'h42795cb2, 32'h424f48c9, 32'h428160b5, 32'h427208a0, 32'h413dbbcd, 32'h4299aa33, 32'hc16c9774, 32'h4284c2d7};
test_output[13992:13999] = '{32'h42795cb2, 32'h424f48c9, 32'h428160b5, 32'h427208a0, 32'h413dbbcd, 32'h4299aa33, 32'h0, 32'h4284c2d7};
test_input[14000:14007] = '{32'hc10d11ab, 32'h423cc008, 32'hc1d6dc62, 32'h41874ba8, 32'hc2a1526e, 32'h42847db0, 32'h41919c50, 32'h4241c45f};
test_output[14000:14007] = '{32'h0, 32'h423cc008, 32'h0, 32'h41874ba8, 32'h0, 32'h42847db0, 32'h41919c50, 32'h4241c45f};
test_input[14008:14015] = '{32'hc2540941, 32'hc229ac5f, 32'h422aa1c8, 32'hc1c641a1, 32'h4210d8cf, 32'h407b6613, 32'hc251616b, 32'h425bfe0b};
test_output[14008:14015] = '{32'h0, 32'h0, 32'h422aa1c8, 32'h0, 32'h4210d8cf, 32'h407b6613, 32'h0, 32'h425bfe0b};
test_input[14016:14023] = '{32'hc2505352, 32'hc171f52f, 32'h4206966e, 32'hc114947b, 32'hc2939fee, 32'h42b03b81, 32'hc04190af, 32'hc2ac1900};
test_output[14016:14023] = '{32'h0, 32'h0, 32'h4206966e, 32'h0, 32'h0, 32'h42b03b81, 32'h0, 32'h0};
test_input[14024:14031] = '{32'hc1920002, 32'h42a22846, 32'h42a0d745, 32'h42c346db, 32'hc2518fff, 32'h42c6ba72, 32'h41d00f10, 32'h422aa078};
test_output[14024:14031] = '{32'h0, 32'h42a22846, 32'h42a0d745, 32'h42c346db, 32'h0, 32'h42c6ba72, 32'h41d00f10, 32'h422aa078};
test_input[14032:14039] = '{32'hc2296db0, 32'hc1f611c9, 32'h4222bd1a, 32'h41fd1817, 32'hc2981f5d, 32'hc270ebdf, 32'hc0acf29b, 32'h413e301f};
test_output[14032:14039] = '{32'h0, 32'h0, 32'h4222bd1a, 32'h41fd1817, 32'h0, 32'h0, 32'h0, 32'h413e301f};
test_input[14040:14047] = '{32'hc250d874, 32'h424d4351, 32'h421022e8, 32'h425f6b78, 32'hc20366fe, 32'h42ba686e, 32'hc1e3e40a, 32'h42942574};
test_output[14040:14047] = '{32'h0, 32'h424d4351, 32'h421022e8, 32'h425f6b78, 32'h0, 32'h42ba686e, 32'h0, 32'h42942574};
test_input[14048:14055] = '{32'h428e526a, 32'h42c5e2e9, 32'hc24f1e67, 32'h425822de, 32'h42959df1, 32'h4281c9ad, 32'hc109eace, 32'hc24d987d};
test_output[14048:14055] = '{32'h428e526a, 32'h42c5e2e9, 32'h0, 32'h425822de, 32'h42959df1, 32'h4281c9ad, 32'h0, 32'h0};
test_input[14056:14063] = '{32'h423c8519, 32'hc2992121, 32'hc20c5139, 32'h423ee370, 32'h419c83f6, 32'hc0047c58, 32'hc0596c5a, 32'hc2c158db};
test_output[14056:14063] = '{32'h423c8519, 32'h0, 32'h0, 32'h423ee370, 32'h419c83f6, 32'h0, 32'h0, 32'h0};
test_input[14064:14071] = '{32'h411e9101, 32'hc2a8073f, 32'hc2a66728, 32'h429ab9f0, 32'hc20c9c2e, 32'h42a1de0b, 32'hc281b6a9, 32'hc1e78050};
test_output[14064:14071] = '{32'h411e9101, 32'h0, 32'h0, 32'h429ab9f0, 32'h0, 32'h42a1de0b, 32'h0, 32'h0};
test_input[14072:14079] = '{32'h423cb6b5, 32'hc1be64f1, 32'h41bfb82a, 32'h41aae9a0, 32'hc2140edb, 32'hc2832b5e, 32'hc130a786, 32'h41dc72ec};
test_output[14072:14079] = '{32'h423cb6b5, 32'h0, 32'h41bfb82a, 32'h41aae9a0, 32'h0, 32'h0, 32'h0, 32'h41dc72ec};
test_input[14080:14087] = '{32'hc1f53bf0, 32'hc198dc7b, 32'hc29e514c, 32'h42b7204f, 32'hc2554f1f, 32'hbfd41e71, 32'h429f647e, 32'h41a8d62a};
test_output[14080:14087] = '{32'h0, 32'h0, 32'h0, 32'h42b7204f, 32'h0, 32'h0, 32'h429f647e, 32'h41a8d62a};
test_input[14088:14095] = '{32'h41ffd32c, 32'hc282f346, 32'h42ad8103, 32'hc24baac3, 32'hc2253e5c, 32'h42a77dae, 32'hc2b65819, 32'h42a28630};
test_output[14088:14095] = '{32'h41ffd32c, 32'h0, 32'h42ad8103, 32'h0, 32'h0, 32'h42a77dae, 32'h0, 32'h42a28630};
test_input[14096:14103] = '{32'h411244c5, 32'hc20ef98d, 32'h424d76a2, 32'hc2c52390, 32'hc2c314df, 32'hc2992a64, 32'hc1cc4803, 32'h42b47cc6};
test_output[14096:14103] = '{32'h411244c5, 32'h0, 32'h424d76a2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b47cc6};
test_input[14104:14111] = '{32'h41044db0, 32'hc2c5f28e, 32'hc14a74b0, 32'hc178eeb8, 32'h41b7915c, 32'hc2b04322, 32'hc2adb093, 32'h41bc8420};
test_output[14104:14111] = '{32'h41044db0, 32'h0, 32'h0, 32'h0, 32'h41b7915c, 32'h0, 32'h0, 32'h41bc8420};
test_input[14112:14119] = '{32'h42175a4d, 32'h4235333f, 32'h3f833b29, 32'hc1107079, 32'hc1813d1c, 32'h423f7dd0, 32'h4283e579, 32'h4129082f};
test_output[14112:14119] = '{32'h42175a4d, 32'h4235333f, 32'h3f833b29, 32'h0, 32'h0, 32'h423f7dd0, 32'h4283e579, 32'h4129082f};
test_input[14120:14127] = '{32'hc264f0fc, 32'hc203165b, 32'hc1d6fe85, 32'h41e99955, 32'hc167a6b2, 32'hc206c085, 32'hc09c4788, 32'hc1f38d9e};
test_output[14120:14127] = '{32'h0, 32'h0, 32'h0, 32'h41e99955, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14128:14135] = '{32'h41ce1d6c, 32'hc213eeb3, 32'h426d2cf8, 32'hc26a48a1, 32'hc264b4fc, 32'h423385e7, 32'hc2beaeb4, 32'hc29841bc};
test_output[14128:14135] = '{32'h41ce1d6c, 32'h0, 32'h426d2cf8, 32'h0, 32'h0, 32'h423385e7, 32'h0, 32'h0};
test_input[14136:14143] = '{32'h419b6c26, 32'hc1c90cfc, 32'h4189781e, 32'hc2c660ff, 32'hc27bf0fb, 32'h41cfba68, 32'h4271b33f, 32'h41a67d65};
test_output[14136:14143] = '{32'h419b6c26, 32'h0, 32'h4189781e, 32'h0, 32'h0, 32'h41cfba68, 32'h4271b33f, 32'h41a67d65};
test_input[14144:14151] = '{32'hc1452a2d, 32'h427ada02, 32'h423e6c58, 32'hc18c2581, 32'hc2b7ea80, 32'h40f7e9ae, 32'h4254a9d6, 32'h429839e6};
test_output[14144:14151] = '{32'h0, 32'h427ada02, 32'h423e6c58, 32'h0, 32'h0, 32'h40f7e9ae, 32'h4254a9d6, 32'h429839e6};
test_input[14152:14159] = '{32'hc1f8c76a, 32'h42c40431, 32'hc24f10a7, 32'hc1ae9cc2, 32'h42aad89a, 32'h41a91742, 32'hc2c6c782, 32'h429c3891};
test_output[14152:14159] = '{32'h0, 32'h42c40431, 32'h0, 32'h0, 32'h42aad89a, 32'h41a91742, 32'h0, 32'h429c3891};
test_input[14160:14167] = '{32'hc24b63ed, 32'h41859ec9, 32'hc1f4bdd9, 32'hc0cbd6f7, 32'hc21115be, 32'hc26b5c23, 32'hc2942d00, 32'hc1b0a34b};
test_output[14160:14167] = '{32'h0, 32'h41859ec9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14168:14175] = '{32'hc270cb5f, 32'h423208ef, 32'h4240bd54, 32'h418bd84d, 32'hc171e5ca, 32'h40f6b8e6, 32'hc10b8607, 32'hc2340317};
test_output[14168:14175] = '{32'h0, 32'h423208ef, 32'h4240bd54, 32'h418bd84d, 32'h0, 32'h40f6b8e6, 32'h0, 32'h0};
test_input[14176:14183] = '{32'hc28f6de5, 32'h41b3a015, 32'h413aade7, 32'h42bab8b2, 32'h4261f2dd, 32'h428d349c, 32'h41d9a251, 32'h42af3f9c};
test_output[14176:14183] = '{32'h0, 32'h41b3a015, 32'h413aade7, 32'h42bab8b2, 32'h4261f2dd, 32'h428d349c, 32'h41d9a251, 32'h42af3f9c};
test_input[14184:14191] = '{32'h42226a59, 32'h40d7353f, 32'hc281262b, 32'hc2836a11, 32'h4286476c, 32'h421b2d9d, 32'hc0fc57bf, 32'h422ab04a};
test_output[14184:14191] = '{32'h42226a59, 32'h40d7353f, 32'h0, 32'h0, 32'h4286476c, 32'h421b2d9d, 32'h0, 32'h422ab04a};
test_input[14192:14199] = '{32'h422ff7b2, 32'h42903355, 32'hc25afd36, 32'h42469f0b, 32'h4145ffdd, 32'h42ae2e4e, 32'hc27a6197, 32'hc2913ede};
test_output[14192:14199] = '{32'h422ff7b2, 32'h42903355, 32'h0, 32'h42469f0b, 32'h4145ffdd, 32'h42ae2e4e, 32'h0, 32'h0};
test_input[14200:14207] = '{32'hc112ba96, 32'h41fcc05c, 32'hbe90d4b9, 32'h42133083, 32'h42a19f08, 32'hc19686a4, 32'hc1395f07, 32'hc114b3fc};
test_output[14200:14207] = '{32'h0, 32'h41fcc05c, 32'h0, 32'h42133083, 32'h42a19f08, 32'h0, 32'h0, 32'h0};
test_input[14208:14215] = '{32'h41dae7d1, 32'hc21b16c4, 32'h425a7903, 32'hc2888aa5, 32'hc2a881e8, 32'hc20ae4df, 32'hc1848fbd, 32'h4224080c};
test_output[14208:14215] = '{32'h41dae7d1, 32'h0, 32'h425a7903, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4224080c};
test_input[14216:14223] = '{32'hc1cd604b, 32'hc1ccba4d, 32'hc2ac1cba, 32'hc18857c4, 32'hc2a6a2ec, 32'h41e1156f, 32'h42b9dfa0, 32'hc197071d};
test_output[14216:14223] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41e1156f, 32'h42b9dfa0, 32'h0};
test_input[14224:14231] = '{32'h42296ce9, 32'hc29e976a, 32'hc1f1f44b, 32'h426f50ea, 32'hc2b97130, 32'hc29e711a, 32'h40438aa3, 32'hc224b128};
test_output[14224:14231] = '{32'h42296ce9, 32'h0, 32'h0, 32'h426f50ea, 32'h0, 32'h0, 32'h40438aa3, 32'h0};
test_input[14232:14239] = '{32'hc2365e66, 32'hc1f42d72, 32'hc20587ae, 32'h4255968a, 32'h41fc9d7b, 32'hc290145f, 32'hc1ba935b, 32'h40102a14};
test_output[14232:14239] = '{32'h0, 32'h0, 32'h0, 32'h4255968a, 32'h41fc9d7b, 32'h0, 32'h0, 32'h40102a14};
test_input[14240:14247] = '{32'hc1137ccc, 32'h40b388f5, 32'hc1c188ce, 32'hc18a9222, 32'hc1092bb0, 32'h42c14b88, 32'hc1ce03c7, 32'hc1f260c8};
test_output[14240:14247] = '{32'h0, 32'h40b388f5, 32'h0, 32'h0, 32'h0, 32'h42c14b88, 32'h0, 32'h0};
test_input[14248:14255] = '{32'h424715c3, 32'h413a1a22, 32'h3f39bbc7, 32'hc2166ca3, 32'h404bcc9b, 32'hc28eec18, 32'hc294d285, 32'hc2745346};
test_output[14248:14255] = '{32'h424715c3, 32'h413a1a22, 32'h3f39bbc7, 32'h0, 32'h404bcc9b, 32'h0, 32'h0, 32'h0};
test_input[14256:14263] = '{32'h40bb11e1, 32'hc2c346b6, 32'hc1b3950a, 32'h41aecd78, 32'hc24d45e2, 32'hc242d021, 32'h423467b9, 32'h41cedab1};
test_output[14256:14263] = '{32'h40bb11e1, 32'h0, 32'h0, 32'h41aecd78, 32'h0, 32'h0, 32'h423467b9, 32'h41cedab1};
test_input[14264:14271] = '{32'h424e2d52, 32'h429aadd6, 32'hc19dae75, 32'hc20dbeef, 32'hc12570f6, 32'hc17aec7d, 32'h41a46830, 32'h42b8d8dc};
test_output[14264:14271] = '{32'h424e2d52, 32'h429aadd6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41a46830, 32'h42b8d8dc};
test_input[14272:14279] = '{32'hc248a701, 32'hc259547a, 32'hc26b66f4, 32'hc297575d, 32'hc228932b, 32'h428fb091, 32'h426c92e3, 32'h423048e3};
test_output[14272:14279] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428fb091, 32'h426c92e3, 32'h423048e3};
test_input[14280:14287] = '{32'hc258fb70, 32'h4263fc50, 32'hc23b267f, 32'hc16d26ba, 32'hc28fcc4b, 32'hc2836e65, 32'h4072643b, 32'h41260d2b};
test_output[14280:14287] = '{32'h0, 32'h4263fc50, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4072643b, 32'h41260d2b};
test_input[14288:14295] = '{32'hc297c3fb, 32'h40ab0fe3, 32'h41cc0fef, 32'h421b711e, 32'h4259c2b4, 32'h40ca9846, 32'hbfffa0ad, 32'hc0cd83f4};
test_output[14288:14295] = '{32'h0, 32'h40ab0fe3, 32'h41cc0fef, 32'h421b711e, 32'h4259c2b4, 32'h40ca9846, 32'h0, 32'h0};
test_input[14296:14303] = '{32'h411d1a41, 32'hc2b3faa2, 32'h424f11c4, 32'hc16acdb2, 32'hc0f722d3, 32'hc01571a8, 32'h4228e9e7, 32'h416b347a};
test_output[14296:14303] = '{32'h411d1a41, 32'h0, 32'h424f11c4, 32'h0, 32'h0, 32'h0, 32'h4228e9e7, 32'h416b347a};
test_input[14304:14311] = '{32'hc2b957f4, 32'hc2aad4b1, 32'hc2655e71, 32'h4278173a, 32'h4290fca3, 32'hc2c19b1b, 32'hc2514412, 32'hc2241ffd};
test_output[14304:14311] = '{32'h0, 32'h0, 32'h0, 32'h4278173a, 32'h4290fca3, 32'h0, 32'h0, 32'h0};
test_input[14312:14319] = '{32'hc271551c, 32'hc293ba52, 32'h4290c4aa, 32'hc1ad4809, 32'h41094bc0, 32'hc2958770, 32'h40fcec10, 32'h42447a08};
test_output[14312:14319] = '{32'h0, 32'h0, 32'h4290c4aa, 32'h0, 32'h41094bc0, 32'h0, 32'h40fcec10, 32'h42447a08};
test_input[14320:14327] = '{32'h42c1c8a1, 32'h42c686f4, 32'h41b049dd, 32'h4224b844, 32'hc1551be5, 32'h4207767c, 32'h4081f407, 32'h42c3bdc4};
test_output[14320:14327] = '{32'h42c1c8a1, 32'h42c686f4, 32'h41b049dd, 32'h4224b844, 32'h0, 32'h4207767c, 32'h4081f407, 32'h42c3bdc4};
test_input[14328:14335] = '{32'hc2a5fa19, 32'h41dda4d3, 32'h416abaa4, 32'hc2208a18, 32'h41d80e56, 32'h429b58be, 32'h42b9547f, 32'hc16ebce9};
test_output[14328:14335] = '{32'h0, 32'h41dda4d3, 32'h416abaa4, 32'h0, 32'h41d80e56, 32'h429b58be, 32'h42b9547f, 32'h0};
test_input[14336:14343] = '{32'h428d2e0a, 32'h4223f14f, 32'h410dbaaf, 32'hc1a6f147, 32'h41e5cc8d, 32'h4187d50a, 32'hc1d7aec8, 32'hc24d8a41};
test_output[14336:14343] = '{32'h428d2e0a, 32'h4223f14f, 32'h410dbaaf, 32'h0, 32'h41e5cc8d, 32'h4187d50a, 32'h0, 32'h0};
test_input[14344:14351] = '{32'h42861a6b, 32'hc2967758, 32'h42819311, 32'hc0c1fd1c, 32'h425fbd0a, 32'h4283c102, 32'h42485a63, 32'h42a02418};
test_output[14344:14351] = '{32'h42861a6b, 32'h0, 32'h42819311, 32'h0, 32'h425fbd0a, 32'h4283c102, 32'h42485a63, 32'h42a02418};
test_input[14352:14359] = '{32'h4252451b, 32'h42a90aa8, 32'h42bc02e1, 32'h42709c23, 32'h41de63cf, 32'hc1cc5c9e, 32'h42b3108f, 32'hc1c0e2d2};
test_output[14352:14359] = '{32'h4252451b, 32'h42a90aa8, 32'h42bc02e1, 32'h42709c23, 32'h41de63cf, 32'h0, 32'h42b3108f, 32'h0};
test_input[14360:14367] = '{32'hc1b43abe, 32'hc2c73d11, 32'h429ba7df, 32'h419c0ee5, 32'h3f7c024b, 32'hc295b0fe, 32'h41890120, 32'hc162f686};
test_output[14360:14367] = '{32'h0, 32'h0, 32'h429ba7df, 32'h419c0ee5, 32'h3f7c024b, 32'h0, 32'h41890120, 32'h0};
test_input[14368:14375] = '{32'h40e58a6e, 32'hc2372b8a, 32'hc1cead62, 32'h4210aeb5, 32'h4169787b, 32'hc29422fa, 32'hc2b701d3, 32'hc1392367};
test_output[14368:14375] = '{32'h40e58a6e, 32'h0, 32'h0, 32'h4210aeb5, 32'h4169787b, 32'h0, 32'h0, 32'h0};
test_input[14376:14383] = '{32'hc2834710, 32'hc24a7b41, 32'h42bf6339, 32'hc2961655, 32'h42a6e28a, 32'hc2a14589, 32'hc2c15fe2, 32'hc27d6b66};
test_output[14376:14383] = '{32'h0, 32'h0, 32'h42bf6339, 32'h0, 32'h42a6e28a, 32'h0, 32'h0, 32'h0};
test_input[14384:14391] = '{32'h428711d2, 32'hc2a39223, 32'hc2be54ab, 32'h413828f9, 32'hc2887933, 32'hc29e40f9, 32'h421ddce4, 32'h40fbb658};
test_output[14384:14391] = '{32'h428711d2, 32'h0, 32'h0, 32'h413828f9, 32'h0, 32'h0, 32'h421ddce4, 32'h40fbb658};
test_input[14392:14399] = '{32'hc266fd67, 32'hc24e60be, 32'h41829dfd, 32'h4297e7e0, 32'hc22920ed, 32'h428df8de, 32'hc261a66b, 32'h429b4016};
test_output[14392:14399] = '{32'h0, 32'h0, 32'h41829dfd, 32'h4297e7e0, 32'h0, 32'h428df8de, 32'h0, 32'h429b4016};
test_input[14400:14407] = '{32'hc0ba6b2f, 32'h42b44606, 32'h423e67a6, 32'h4294a601, 32'hc25628cc, 32'h415badb9, 32'hc291c977, 32'h422dff6a};
test_output[14400:14407] = '{32'h0, 32'h42b44606, 32'h423e67a6, 32'h4294a601, 32'h0, 32'h415badb9, 32'h0, 32'h422dff6a};
test_input[14408:14415] = '{32'hc28fd2df, 32'hc18a7b32, 32'h4250d2e5, 32'hc2a29b10, 32'hc280c20b, 32'h4241edbc, 32'hc242aee2, 32'h42386e6a};
test_output[14408:14415] = '{32'h0, 32'h0, 32'h4250d2e5, 32'h0, 32'h0, 32'h4241edbc, 32'h0, 32'h42386e6a};
test_input[14416:14423] = '{32'h3fd51c0e, 32'h423f87c9, 32'h41b96711, 32'h42185342, 32'h4247a511, 32'hc2c6845c, 32'hc0c2ab5f, 32'hc25d04da};
test_output[14416:14423] = '{32'h3fd51c0e, 32'h423f87c9, 32'h41b96711, 32'h42185342, 32'h4247a511, 32'h0, 32'h0, 32'h0};
test_input[14424:14431] = '{32'h402a6569, 32'hc22713bd, 32'hc2bee173, 32'hc23735f4, 32'h4288c191, 32'hc1d6aa6f, 32'hc279b9ba, 32'h42b6dd0a};
test_output[14424:14431] = '{32'h402a6569, 32'h0, 32'h0, 32'h0, 32'h4288c191, 32'h0, 32'h0, 32'h42b6dd0a};
test_input[14432:14439] = '{32'hc2975968, 32'h41b624d6, 32'h428712ee, 32'hc28547e1, 32'hc2ae60b3, 32'h42a61906, 32'hc0bbb790, 32'hc2ad1488};
test_output[14432:14439] = '{32'h0, 32'h41b624d6, 32'h428712ee, 32'h0, 32'h0, 32'h42a61906, 32'h0, 32'h0};
test_input[14440:14447] = '{32'hc111f09f, 32'hc1510d66, 32'hc27aa9b7, 32'h428fbfe1, 32'hc20311cc, 32'hc2a3fcb2, 32'h41cf6f3e, 32'h428f3974};
test_output[14440:14447] = '{32'h0, 32'h0, 32'h0, 32'h428fbfe1, 32'h0, 32'h0, 32'h41cf6f3e, 32'h428f3974};
test_input[14448:14455] = '{32'hc20439ac, 32'h4294643b, 32'h42bfe131, 32'h41610ce9, 32'h3f03ceb9, 32'h429f35fc, 32'h420cc4ca, 32'h42b0eb59};
test_output[14448:14455] = '{32'h0, 32'h4294643b, 32'h42bfe131, 32'h41610ce9, 32'h3f03ceb9, 32'h429f35fc, 32'h420cc4ca, 32'h42b0eb59};
test_input[14456:14463] = '{32'h429671a7, 32'h4239ff6d, 32'h41758505, 32'h4287f10e, 32'h4289e0e3, 32'hc29aa635, 32'h42214a9f, 32'hc21fad34};
test_output[14456:14463] = '{32'h429671a7, 32'h4239ff6d, 32'h41758505, 32'h4287f10e, 32'h4289e0e3, 32'h0, 32'h42214a9f, 32'h0};
test_input[14464:14471] = '{32'h429c7c78, 32'h4234f718, 32'h4050c2fd, 32'hc24e0736, 32'h4289c579, 32'hc2b909c9, 32'hc28b1262, 32'hc219b836};
test_output[14464:14471] = '{32'h429c7c78, 32'h4234f718, 32'h4050c2fd, 32'h0, 32'h4289c579, 32'h0, 32'h0, 32'h0};
test_input[14472:14479] = '{32'hc2982f58, 32'h4195cfa6, 32'hc1ced7ed, 32'hc10f2f41, 32'hc282756c, 32'h42bdd764, 32'h4289bc73, 32'hc1b5ff84};
test_output[14472:14479] = '{32'h0, 32'h4195cfa6, 32'h0, 32'h0, 32'h0, 32'h42bdd764, 32'h4289bc73, 32'h0};
test_input[14480:14487] = '{32'hc2a75888, 32'h41bb3ff2, 32'h42bb162a, 32'h4118abe4, 32'hc23b582b, 32'hc1afdfd9, 32'h42bec7f0, 32'hc29e8500};
test_output[14480:14487] = '{32'h0, 32'h41bb3ff2, 32'h42bb162a, 32'h4118abe4, 32'h0, 32'h0, 32'h42bec7f0, 32'h0};
test_input[14488:14495] = '{32'h4215bcaf, 32'hc28febcc, 32'h42824967, 32'h427c4624, 32'h422a9fe2, 32'hc0e39d0c, 32'hc2a00145, 32'hc2c09614};
test_output[14488:14495] = '{32'h4215bcaf, 32'h0, 32'h42824967, 32'h427c4624, 32'h422a9fe2, 32'h0, 32'h0, 32'h0};
test_input[14496:14503] = '{32'hc162ea39, 32'hc12833c4, 32'h42b07066, 32'h41d9de31, 32'h429dbc11, 32'h408e08bd, 32'hc2377b29, 32'h3f99ab5e};
test_output[14496:14503] = '{32'h0, 32'h0, 32'h42b07066, 32'h41d9de31, 32'h429dbc11, 32'h408e08bd, 32'h0, 32'h3f99ab5e};
test_input[14504:14511] = '{32'hc282a5f1, 32'hc2ae9fd4, 32'h42ad10e6, 32'h41b3984d, 32'hc18eb6c4, 32'hc211fc52, 32'hc28bf86c, 32'h42c590e4};
test_output[14504:14511] = '{32'h0, 32'h0, 32'h42ad10e6, 32'h41b3984d, 32'h0, 32'h0, 32'h0, 32'h42c590e4};
test_input[14512:14519] = '{32'hc2b0341b, 32'h41c2fc5a, 32'hc26f450e, 32'h422e3188, 32'h427e7c8c, 32'hc25e4921, 32'hc2423690, 32'h4162577c};
test_output[14512:14519] = '{32'h0, 32'h41c2fc5a, 32'h0, 32'h422e3188, 32'h427e7c8c, 32'h0, 32'h0, 32'h4162577c};
test_input[14520:14527] = '{32'hc2836d1b, 32'h426cf520, 32'h41b3dd75, 32'hc25f413f, 32'h42558763, 32'hc2aab0ab, 32'hc23f866a, 32'hc28f09ed};
test_output[14520:14527] = '{32'h0, 32'h426cf520, 32'h41b3dd75, 32'h0, 32'h42558763, 32'h0, 32'h0, 32'h0};
test_input[14528:14535] = '{32'hc01a3f4b, 32'hc05c1522, 32'h426b45f0, 32'h41f5138a, 32'h425de87e, 32'hc005f7e9, 32'h4297f35f, 32'hc2a0ef2a};
test_output[14528:14535] = '{32'h0, 32'h0, 32'h426b45f0, 32'h41f5138a, 32'h425de87e, 32'h0, 32'h4297f35f, 32'h0};
test_input[14536:14543] = '{32'hc2b40aca, 32'hc2941710, 32'hc28d3e51, 32'h4200ba92, 32'h4298f406, 32'hc28e903e, 32'hc0bb5dc7, 32'h40fad5d7};
test_output[14536:14543] = '{32'h0, 32'h0, 32'h0, 32'h4200ba92, 32'h4298f406, 32'h0, 32'h0, 32'h40fad5d7};
test_input[14544:14551] = '{32'h404482d7, 32'hc256289a, 32'h42a3d1b3, 32'hc2bd362d, 32'h40675172, 32'h40f6ebdc, 32'h42431054, 32'hc1c71559};
test_output[14544:14551] = '{32'h404482d7, 32'h0, 32'h42a3d1b3, 32'h0, 32'h40675172, 32'h40f6ebdc, 32'h42431054, 32'h0};
test_input[14552:14559] = '{32'hc2ab8dc3, 32'h422a635f, 32'hc2521ae8, 32'hc2659fff, 32'h4289b6d1, 32'h41c2805c, 32'h41b2a0c6, 32'hc1934d42};
test_output[14552:14559] = '{32'h0, 32'h422a635f, 32'h0, 32'h0, 32'h4289b6d1, 32'h41c2805c, 32'h41b2a0c6, 32'h0};
test_input[14560:14567] = '{32'h4206ca72, 32'h42458569, 32'h423af1c3, 32'hc182d64a, 32'hc1b1d7d3, 32'hc29247e1, 32'h42aab11b, 32'hc2ba8e93};
test_output[14560:14567] = '{32'h4206ca72, 32'h42458569, 32'h423af1c3, 32'h0, 32'h0, 32'h0, 32'h42aab11b, 32'h0};
test_input[14568:14575] = '{32'h4282b50c, 32'hc117f728, 32'hc2b8d2b8, 32'h42b4df74, 32'hc1c20a4e, 32'hc16e6dcf, 32'hc24b583f, 32'h4245d2d6};
test_output[14568:14575] = '{32'h4282b50c, 32'h0, 32'h0, 32'h42b4df74, 32'h0, 32'h0, 32'h0, 32'h4245d2d6};
test_input[14576:14583] = '{32'h42428c46, 32'h420a3621, 32'h420822e1, 32'hc13dd0b0, 32'h4251fce4, 32'h427f85cf, 32'h405efb1b, 32'h41df0980};
test_output[14576:14583] = '{32'h42428c46, 32'h420a3621, 32'h420822e1, 32'h0, 32'h4251fce4, 32'h427f85cf, 32'h405efb1b, 32'h41df0980};
test_input[14584:14591] = '{32'hc2b48d3d, 32'h4233fd8a, 32'h41a9d00d, 32'hc261832d, 32'h41d2b1bf, 32'h42669009, 32'h4297f1f6, 32'h42082987};
test_output[14584:14591] = '{32'h0, 32'h4233fd8a, 32'h41a9d00d, 32'h0, 32'h41d2b1bf, 32'h42669009, 32'h4297f1f6, 32'h42082987};
test_input[14592:14599] = '{32'h3fa4e727, 32'h4262bd95, 32'hc1fc5fec, 32'hc273262c, 32'hc1ce6930, 32'h42bb1b14, 32'h4243ef31, 32'h42481a63};
test_output[14592:14599] = '{32'h3fa4e727, 32'h4262bd95, 32'h0, 32'h0, 32'h0, 32'h42bb1b14, 32'h4243ef31, 32'h42481a63};
test_input[14600:14607] = '{32'h4288a7c8, 32'hc25e9a95, 32'h4053ea8b, 32'hc2b05629, 32'h41fdce04, 32'hc2b78328, 32'hc2868b68, 32'h42a8ec4d};
test_output[14600:14607] = '{32'h4288a7c8, 32'h0, 32'h4053ea8b, 32'h0, 32'h41fdce04, 32'h0, 32'h0, 32'h42a8ec4d};
test_input[14608:14615] = '{32'h41700db5, 32'hc2bd448c, 32'h415e5c69, 32'hc2a63ba8, 32'h40fb187d, 32'hc0fbda0c, 32'hc2161103, 32'hc2788a39};
test_output[14608:14615] = '{32'h41700db5, 32'h0, 32'h415e5c69, 32'h0, 32'h40fb187d, 32'h0, 32'h0, 32'h0};
test_input[14616:14623] = '{32'h428099d1, 32'hc24cb659, 32'hc19aa5ae, 32'h426886df, 32'h4219c53d, 32'hc24c1da1, 32'h426ec2cd, 32'hc25c0bc6};
test_output[14616:14623] = '{32'h428099d1, 32'h0, 32'h0, 32'h426886df, 32'h4219c53d, 32'h0, 32'h426ec2cd, 32'h0};
test_input[14624:14631] = '{32'h41cb0b94, 32'hc19f367d, 32'hc27044a0, 32'hc165811a, 32'hc2b8fd29, 32'h417e05cf, 32'hc21c48a7, 32'h418d2b84};
test_output[14624:14631] = '{32'h41cb0b94, 32'h0, 32'h0, 32'h0, 32'h0, 32'h417e05cf, 32'h0, 32'h418d2b84};
test_input[14632:14639] = '{32'h413775f3, 32'h418668f2, 32'h4221507e, 32'hc0e9c713, 32'h422c4acf, 32'hc2b64864, 32'hc2bd92b8, 32'h4220102a};
test_output[14632:14639] = '{32'h413775f3, 32'h418668f2, 32'h4221507e, 32'h0, 32'h422c4acf, 32'h0, 32'h0, 32'h4220102a};
test_input[14640:14647] = '{32'h40a8ed52, 32'hc214c1ba, 32'hc2bd940c, 32'h429ef827, 32'hc1616e01, 32'h425b9dd3, 32'h42142e73, 32'h411c31a6};
test_output[14640:14647] = '{32'h40a8ed52, 32'h0, 32'h0, 32'h429ef827, 32'h0, 32'h425b9dd3, 32'h42142e73, 32'h411c31a6};
test_input[14648:14655] = '{32'h42472bee, 32'hc1df0cff, 32'h42b5520c, 32'hc2b50904, 32'h420bae18, 32'h42b54d38, 32'h42a661cd, 32'hc24b402b};
test_output[14648:14655] = '{32'h42472bee, 32'h0, 32'h42b5520c, 32'h0, 32'h420bae18, 32'h42b54d38, 32'h42a661cd, 32'h0};
test_input[14656:14663] = '{32'hc13b966f, 32'h427e667a, 32'hc2a1a4ad, 32'h42b310bb, 32'hc25b465d, 32'h4204479a, 32'h41ecd71c, 32'h4278df51};
test_output[14656:14663] = '{32'h0, 32'h427e667a, 32'h0, 32'h42b310bb, 32'h0, 32'h4204479a, 32'h41ecd71c, 32'h4278df51};
test_input[14664:14671] = '{32'h4267aaa5, 32'hc1a1d944, 32'h42259a8e, 32'h425021cc, 32'hc14d3edb, 32'hc16097d4, 32'h4273f35d, 32'h42273b74};
test_output[14664:14671] = '{32'h4267aaa5, 32'h0, 32'h42259a8e, 32'h425021cc, 32'h0, 32'h0, 32'h4273f35d, 32'h42273b74};
test_input[14672:14679] = '{32'h421e1d67, 32'h41065299, 32'hc2c48b09, 32'hc1d41f0b, 32'h425873ad, 32'h407096fe, 32'h41c22079, 32'hc2b17178};
test_output[14672:14679] = '{32'h421e1d67, 32'h41065299, 32'h0, 32'h0, 32'h425873ad, 32'h407096fe, 32'h41c22079, 32'h0};
test_input[14680:14687] = '{32'h41e11378, 32'hc2b605d3, 32'h419cdb50, 32'h4186a07c, 32'h42a5bab3, 32'h41831c50, 32'hc2a19d52, 32'hc26ddabc};
test_output[14680:14687] = '{32'h41e11378, 32'h0, 32'h419cdb50, 32'h4186a07c, 32'h42a5bab3, 32'h41831c50, 32'h0, 32'h0};
test_input[14688:14695] = '{32'h425efc14, 32'h41a9ae07, 32'h4296d08e, 32'hc1414e16, 32'hc29bf165, 32'hc09bed3c, 32'h42b9d0b1, 32'hc2c633aa};
test_output[14688:14695] = '{32'h425efc14, 32'h41a9ae07, 32'h4296d08e, 32'h0, 32'h0, 32'h0, 32'h42b9d0b1, 32'h0};
test_input[14696:14703] = '{32'h42adb0a6, 32'h4238cdf1, 32'hc07f54e2, 32'hc09605a3, 32'hc28d2ec1, 32'hc22f60f8, 32'hc0eb0fc8, 32'h424cec7b};
test_output[14696:14703] = '{32'h42adb0a6, 32'h4238cdf1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h424cec7b};
test_input[14704:14711] = '{32'hc1c051ee, 32'hc2c4bf7b, 32'hc25dcf46, 32'hc2a2130f, 32'hc0344ff3, 32'h42be61bc, 32'hc27f3cdb, 32'h400e15b6};
test_output[14704:14711] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42be61bc, 32'h0, 32'h400e15b6};
test_input[14712:14719] = '{32'hc2b4bd4d, 32'h4289f6ab, 32'h417a0afb, 32'hc28e3ad4, 32'hc26ebf70, 32'hc17a945b, 32'hc29b46bf, 32'hc2a4ac2e};
test_output[14712:14719] = '{32'h0, 32'h4289f6ab, 32'h417a0afb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14720:14727] = '{32'h40cd8e78, 32'hc178bb83, 32'h429fbe81, 32'hc2a39c6e, 32'h41d9628c, 32'h42a5c16a, 32'h428df844, 32'hc1af0c92};
test_output[14720:14727] = '{32'h40cd8e78, 32'h0, 32'h429fbe81, 32'h0, 32'h41d9628c, 32'h42a5c16a, 32'h428df844, 32'h0};
test_input[14728:14735] = '{32'hbfb1ca3a, 32'hc2b62c51, 32'hc227e0ba, 32'h41df5df9, 32'h422b6760, 32'hc092a243, 32'hc1a3c3fa, 32'hc2740bb0};
test_output[14728:14735] = '{32'h0, 32'h0, 32'h0, 32'h41df5df9, 32'h422b6760, 32'h0, 32'h0, 32'h0};
test_input[14736:14743] = '{32'hc1cd1f02, 32'hbfd7fc72, 32'h427dcb65, 32'h42b5ccde, 32'h420fd290, 32'h428ec15e, 32'hc28ea35e, 32'hc2bb7220};
test_output[14736:14743] = '{32'h0, 32'h0, 32'h427dcb65, 32'h42b5ccde, 32'h420fd290, 32'h428ec15e, 32'h0, 32'h0};
test_input[14744:14751] = '{32'hc1772fd1, 32'h3f56e8e5, 32'hc27b33ae, 32'h42818b8c, 32'h423348f5, 32'h42aba744, 32'h42aa8669, 32'hc2746049};
test_output[14744:14751] = '{32'h0, 32'h3f56e8e5, 32'h0, 32'h42818b8c, 32'h423348f5, 32'h42aba744, 32'h42aa8669, 32'h0};
test_input[14752:14759] = '{32'h42a45fc4, 32'h41ea15fd, 32'h426b0646, 32'h42a1f147, 32'hc2b8e5e3, 32'hc28e97d6, 32'hc15d3aa2, 32'h40c9fdd2};
test_output[14752:14759] = '{32'h42a45fc4, 32'h41ea15fd, 32'h426b0646, 32'h42a1f147, 32'h0, 32'h0, 32'h0, 32'h40c9fdd2};
test_input[14760:14767] = '{32'h424f0845, 32'h4107012d, 32'hc20235c3, 32'h418f19c8, 32'hc24fe5c3, 32'hc286b33a, 32'hc2a49972, 32'h42a9f581};
test_output[14760:14767] = '{32'h424f0845, 32'h4107012d, 32'h0, 32'h418f19c8, 32'h0, 32'h0, 32'h0, 32'h42a9f581};
test_input[14768:14775] = '{32'h41b822a4, 32'hc1c9a8f2, 32'hc1d558a6, 32'hc22286ee, 32'hc25300dc, 32'h41d48f0f, 32'hc24e0e04, 32'hc166443a};
test_output[14768:14775] = '{32'h41b822a4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41d48f0f, 32'h0, 32'h0};
test_input[14776:14783] = '{32'hc1a8a6e8, 32'h41afa499, 32'hc28407bc, 32'hc2bc31d5, 32'hc2a8de1f, 32'hc0aea5a5, 32'hc1b30fee, 32'hc1d9627e};
test_output[14776:14783] = '{32'h0, 32'h41afa499, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14784:14791] = '{32'hc256efd3, 32'hc27f8404, 32'hc1f2738d, 32'h422664d9, 32'h42c7413e, 32'hc2ba1393, 32'hc2bfd7f8, 32'hc21d5cd2};
test_output[14784:14791] = '{32'h0, 32'h0, 32'h0, 32'h422664d9, 32'h42c7413e, 32'h0, 32'h0, 32'h0};
test_input[14792:14799] = '{32'h4292bbb7, 32'hc2c7cf08, 32'hc09a18ad, 32'hc238052d, 32'h4202f9f8, 32'h4251ada5, 32'hc25df428, 32'h40d982e1};
test_output[14792:14799] = '{32'h4292bbb7, 32'h0, 32'h0, 32'h0, 32'h4202f9f8, 32'h4251ada5, 32'h0, 32'h40d982e1};
test_input[14800:14807] = '{32'hc225e677, 32'hc22af59e, 32'hc27671b3, 32'h416ff708, 32'h41b9e5b8, 32'hc203c359, 32'h41e1fba6, 32'hc23bcb97};
test_output[14800:14807] = '{32'h0, 32'h0, 32'h0, 32'h416ff708, 32'h41b9e5b8, 32'h0, 32'h41e1fba6, 32'h0};
test_input[14808:14815] = '{32'h3fda0116, 32'h427dfc29, 32'hc29eb80b, 32'hc28fb847, 32'h42c74a6e, 32'hc23f49bf, 32'hc295e8f5, 32'h42ab3501};
test_output[14808:14815] = '{32'h3fda0116, 32'h427dfc29, 32'h0, 32'h0, 32'h42c74a6e, 32'h0, 32'h0, 32'h42ab3501};
test_input[14816:14823] = '{32'hc13562d8, 32'hc2a85082, 32'hc2a60f97, 32'hc27d29f2, 32'hc2b89c24, 32'h41b8ebda, 32'h413b0503, 32'h42171b8f};
test_output[14816:14823] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b8ebda, 32'h413b0503, 32'h42171b8f};
test_input[14824:14831] = '{32'hc1b29f14, 32'hc2931bbe, 32'hc14af202, 32'h422731b3, 32'hc285d142, 32'h4260b189, 32'h40d96209, 32'hc2c7e3ae};
test_output[14824:14831] = '{32'h0, 32'h0, 32'h0, 32'h422731b3, 32'h0, 32'h4260b189, 32'h40d96209, 32'h0};
test_input[14832:14839] = '{32'h4200254c, 32'h425ee128, 32'hc1dcb793, 32'hc290571b, 32'h42b73210, 32'h42bfad22, 32'h3ffacf10, 32'h42c00574};
test_output[14832:14839] = '{32'h4200254c, 32'h425ee128, 32'h0, 32'h0, 32'h42b73210, 32'h42bfad22, 32'h3ffacf10, 32'h42c00574};
test_input[14840:14847] = '{32'h419823b2, 32'hc25c08dd, 32'h4248f52d, 32'hc2701ca2, 32'h41e6ea16, 32'hc2c5bfb7, 32'h42a91a90, 32'hc227395a};
test_output[14840:14847] = '{32'h419823b2, 32'h0, 32'h4248f52d, 32'h0, 32'h41e6ea16, 32'h0, 32'h42a91a90, 32'h0};
test_input[14848:14855] = '{32'hc2c2f9e8, 32'hc2388dc6, 32'h429e3ef8, 32'hc29aa0bc, 32'h428dfcbf, 32'hc1de8f82, 32'hc24685d9, 32'h42bd2a37};
test_output[14848:14855] = '{32'h0, 32'h0, 32'h429e3ef8, 32'h0, 32'h428dfcbf, 32'h0, 32'h0, 32'h42bd2a37};
test_input[14856:14863] = '{32'h42b62348, 32'hc2013423, 32'h423b844b, 32'hc1836ad2, 32'hc1e5ac6d, 32'h428d2809, 32'h41fc094a, 32'h4276193d};
test_output[14856:14863] = '{32'h42b62348, 32'h0, 32'h423b844b, 32'h0, 32'h0, 32'h428d2809, 32'h41fc094a, 32'h4276193d};
test_input[14864:14871] = '{32'h42211540, 32'h42a2184a, 32'hc2bd65b4, 32'hc20051d2, 32'h42a319e3, 32'hc2a84414, 32'h4209e4e3, 32'h423e097f};
test_output[14864:14871] = '{32'h42211540, 32'h42a2184a, 32'h0, 32'h0, 32'h42a319e3, 32'h0, 32'h4209e4e3, 32'h423e097f};
test_input[14872:14879] = '{32'hc2204a52, 32'hc2b4979a, 32'h42b1cbb7, 32'h410ddddd, 32'h42b4b8eb, 32'h429a3e26, 32'hc1c82374, 32'hc2127716};
test_output[14872:14879] = '{32'h0, 32'h0, 32'h42b1cbb7, 32'h410ddddd, 32'h42b4b8eb, 32'h429a3e26, 32'h0, 32'h0};
test_input[14880:14887] = '{32'h4287fc98, 32'hc200a765, 32'h428ef0f3, 32'hc2741966, 32'h42b1093d, 32'hc2c43a6e, 32'hc263a837, 32'hc2b7afa9};
test_output[14880:14887] = '{32'h4287fc98, 32'h0, 32'h428ef0f3, 32'h0, 32'h42b1093d, 32'h0, 32'h0, 32'h0};
test_input[14888:14895] = '{32'hc1e4a655, 32'hc24bbc3c, 32'hc114de80, 32'h41f25f2f, 32'h41d03190, 32'hc27384bc, 32'h416c74f3, 32'hc253896f};
test_output[14888:14895] = '{32'h0, 32'h0, 32'h0, 32'h41f25f2f, 32'h41d03190, 32'h0, 32'h416c74f3, 32'h0};
test_input[14896:14903] = '{32'h428f4d0b, 32'h4252160a, 32'hc28cfa18, 32'hc258bae7, 32'h41bcf96a, 32'h4121299f, 32'hc2a1cc2c, 32'hc2bd2209};
test_output[14896:14903] = '{32'h428f4d0b, 32'h4252160a, 32'h0, 32'h0, 32'h41bcf96a, 32'h4121299f, 32'h0, 32'h0};
test_input[14904:14911] = '{32'hc2158b71, 32'h4127687a, 32'hc1bbfc11, 32'hc2bceda5, 32'h425bb88e, 32'h41991122, 32'hc2c3e013, 32'h41df952f};
test_output[14904:14911] = '{32'h0, 32'h4127687a, 32'h0, 32'h0, 32'h425bb88e, 32'h41991122, 32'h0, 32'h41df952f};
test_input[14912:14919] = '{32'h42ac1ff2, 32'h41d835e2, 32'h423444fe, 32'h429472cc, 32'hc2a6d482, 32'h421dc944, 32'h40663a75, 32'hc294c4ad};
test_output[14912:14919] = '{32'h42ac1ff2, 32'h41d835e2, 32'h423444fe, 32'h429472cc, 32'h0, 32'h421dc944, 32'h40663a75, 32'h0};
test_input[14920:14927] = '{32'h42060ac2, 32'h429ea792, 32'hc2997319, 32'h428474f8, 32'hc26332c2, 32'hc1ded14b, 32'hc1dee52c, 32'hc22c4c23};
test_output[14920:14927] = '{32'h42060ac2, 32'h429ea792, 32'h0, 32'h428474f8, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14928:14935] = '{32'hc0afdb0d, 32'hc084acf9, 32'h4214fb99, 32'hc244e66a, 32'hc0f80881, 32'hc287f012, 32'hc28ffb97, 32'hc2b00c2c};
test_output[14928:14935] = '{32'h0, 32'h0, 32'h4214fb99, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14936:14943] = '{32'hc259e6bb, 32'h423e325c, 32'h427f7d76, 32'h42b5e0c8, 32'hc105c023, 32'hc20a9eda, 32'hc1bc1a80, 32'h4182a3c5};
test_output[14936:14943] = '{32'h0, 32'h423e325c, 32'h427f7d76, 32'h42b5e0c8, 32'h0, 32'h0, 32'h0, 32'h4182a3c5};
test_input[14944:14951] = '{32'h42b11ae9, 32'hc16986c6, 32'hc288eedd, 32'hc21715ae, 32'h42b11df9, 32'h4281fd22, 32'hc26b8ffe, 32'h41842439};
test_output[14944:14951] = '{32'h42b11ae9, 32'h0, 32'h0, 32'h0, 32'h42b11df9, 32'h4281fd22, 32'h0, 32'h41842439};
test_input[14952:14959] = '{32'h42ac4a0c, 32'hc2b5a8dc, 32'h41ea3875, 32'h420dec4e, 32'hc27a0c1a, 32'h42c30834, 32'h429fd715, 32'hc2288eed};
test_output[14952:14959] = '{32'h42ac4a0c, 32'h0, 32'h41ea3875, 32'h420dec4e, 32'h0, 32'h42c30834, 32'h429fd715, 32'h0};
test_input[14960:14967] = '{32'hc1866537, 32'h425a74cc, 32'h42c74354, 32'hc296a410, 32'h42bb1ce3, 32'hc1e8cf54, 32'hc2aaa9b2, 32'hc293ea62};
test_output[14960:14967] = '{32'h0, 32'h425a74cc, 32'h42c74354, 32'h0, 32'h42bb1ce3, 32'h0, 32'h0, 32'h0};
test_input[14968:14975] = '{32'h42c2e73b, 32'hc2b76346, 32'h41a86069, 32'h4208fb64, 32'hc2aa356a, 32'h422042c1, 32'hc2b2addf, 32'hc200d7da};
test_output[14968:14975] = '{32'h42c2e73b, 32'h0, 32'h41a86069, 32'h4208fb64, 32'h0, 32'h422042c1, 32'h0, 32'h0};
test_input[14976:14983] = '{32'hc274fedc, 32'h4253ccd4, 32'hc29e46ff, 32'h40de7109, 32'h4266958e, 32'hc2611858, 32'hc1ee286b, 32'hc1f33206};
test_output[14976:14983] = '{32'h0, 32'h4253ccd4, 32'h0, 32'h40de7109, 32'h4266958e, 32'h0, 32'h0, 32'h0};
test_input[14984:14991] = '{32'h42bc8363, 32'hc2721127, 32'h42532120, 32'h41a649dd, 32'hc0b998ab, 32'hc28f94da, 32'h42630231, 32'h42b77da5};
test_output[14984:14991] = '{32'h42bc8363, 32'h0, 32'h42532120, 32'h41a649dd, 32'h0, 32'h0, 32'h42630231, 32'h42b77da5};
test_input[14992:14999] = '{32'hc28eac1f, 32'h3fee5e83, 32'hc2c0e61e, 32'h418db41e, 32'h4255f48d, 32'h42a22472, 32'h4208650e, 32'h4219bc3e};
test_output[14992:14999] = '{32'h0, 32'h3fee5e83, 32'h0, 32'h418db41e, 32'h4255f48d, 32'h42a22472, 32'h4208650e, 32'h4219bc3e};
test_input[15000:15007] = '{32'hc298e4b4, 32'h425ffeca, 32'hc0e3643c, 32'h4257fa60, 32'hc1bc329c, 32'hc27dc4c2, 32'h42717460, 32'hc293d15b};
test_output[15000:15007] = '{32'h0, 32'h425ffeca, 32'h0, 32'h4257fa60, 32'h0, 32'h0, 32'h42717460, 32'h0};
test_input[15008:15015] = '{32'hc23c5a3c, 32'h42608794, 32'h413cbb98, 32'h42191c47, 32'h42119309, 32'hc15783e5, 32'h428e09bd, 32'hc203d836};
test_output[15008:15015] = '{32'h0, 32'h42608794, 32'h413cbb98, 32'h42191c47, 32'h42119309, 32'h0, 32'h428e09bd, 32'h0};
test_input[15016:15023] = '{32'hc28eec9d, 32'h427ac58e, 32'h41f80278, 32'hc2566773, 32'h42c54940, 32'h4284061c, 32'hc28161d8, 32'h426cf91b};
test_output[15016:15023] = '{32'h0, 32'h427ac58e, 32'h41f80278, 32'h0, 32'h42c54940, 32'h4284061c, 32'h0, 32'h426cf91b};
test_input[15024:15031] = '{32'h428fe3bb, 32'hc2099324, 32'hc26a45df, 32'hc2856d1a, 32'h42b28334, 32'hc166d273, 32'hc2848248, 32'h428293fc};
test_output[15024:15031] = '{32'h428fe3bb, 32'h0, 32'h0, 32'h0, 32'h42b28334, 32'h0, 32'h0, 32'h428293fc};
test_input[15032:15039] = '{32'hc2699410, 32'h4283269c, 32'h4192fc62, 32'hc29d29a3, 32'h41bba309, 32'h41acf294, 32'hc2c623aa, 32'h429cc199};
test_output[15032:15039] = '{32'h0, 32'h4283269c, 32'h4192fc62, 32'h0, 32'h41bba309, 32'h41acf294, 32'h0, 32'h429cc199};
test_input[15040:15047] = '{32'h41fd5106, 32'h4288648d, 32'h429b120e, 32'hc29928ed, 32'h42a36319, 32'h42c75aec, 32'h41bf8e59, 32'h4277128f};
test_output[15040:15047] = '{32'h41fd5106, 32'h4288648d, 32'h429b120e, 32'h0, 32'h42a36319, 32'h42c75aec, 32'h41bf8e59, 32'h4277128f};
test_input[15048:15055] = '{32'h423bd65a, 32'hc272ee6e, 32'hc291f00d, 32'h42857d11, 32'hc263ec4c, 32'hc20aa38f, 32'hc2a011ea, 32'h41e6b38e};
test_output[15048:15055] = '{32'h423bd65a, 32'h0, 32'h0, 32'h42857d11, 32'h0, 32'h0, 32'h0, 32'h41e6b38e};
test_input[15056:15063] = '{32'hc14bb032, 32'hc1d94400, 32'h424ae703, 32'h42a3ef3a, 32'hc206c272, 32'h422ac69e, 32'h4215bdb0, 32'hc22d83a2};
test_output[15056:15063] = '{32'h0, 32'h0, 32'h424ae703, 32'h42a3ef3a, 32'h0, 32'h422ac69e, 32'h4215bdb0, 32'h0};
test_input[15064:15071] = '{32'hc1f16d17, 32'hc27f4744, 32'h42a899a6, 32'h42628c1e, 32'h426215f2, 32'h4164146c, 32'hc26ac387, 32'hc2c553a0};
test_output[15064:15071] = '{32'h0, 32'h0, 32'h42a899a6, 32'h42628c1e, 32'h426215f2, 32'h4164146c, 32'h0, 32'h0};
test_input[15072:15079] = '{32'h422cf091, 32'h4104f3a4, 32'h42a1bf40, 32'h4228b3dc, 32'hc2b0f962, 32'hc2ab584a, 32'hc2b55377, 32'hc16b6d7e};
test_output[15072:15079] = '{32'h422cf091, 32'h4104f3a4, 32'h42a1bf40, 32'h4228b3dc, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15080:15087] = '{32'hc2325e23, 32'hc08f8724, 32'hc287659f, 32'hc253868d, 32'hc2420e58, 32'hc241a785, 32'h41e6c94a, 32'hc17bdc41};
test_output[15080:15087] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41e6c94a, 32'h0};
test_input[15088:15095] = '{32'h40795d22, 32'h42a8e86a, 32'hc24aeb8e, 32'h4295f7ae, 32'h411c576b, 32'hc273daae, 32'hc263ce7f, 32'hc2aa969f};
test_output[15088:15095] = '{32'h40795d22, 32'h42a8e86a, 32'h0, 32'h4295f7ae, 32'h411c576b, 32'h0, 32'h0, 32'h0};
test_input[15096:15103] = '{32'hc2ae66df, 32'hc296b64c, 32'h413839a0, 32'hc280b478, 32'hc27e5410, 32'hc2b51a75, 32'h4258a943, 32'h409ff71e};
test_output[15096:15103] = '{32'h0, 32'h0, 32'h413839a0, 32'h0, 32'h0, 32'h0, 32'h4258a943, 32'h409ff71e};
test_input[15104:15111] = '{32'h408974e2, 32'hc2aac136, 32'h4267e3a1, 32'h4193022c, 32'h4264c14b, 32'h42b632b5, 32'hc297358b, 32'hc26d3d9f};
test_output[15104:15111] = '{32'h408974e2, 32'h0, 32'h4267e3a1, 32'h4193022c, 32'h4264c14b, 32'h42b632b5, 32'h0, 32'h0};
test_input[15112:15119] = '{32'h410d22a5, 32'h42943032, 32'h424536b7, 32'hc17c55ec, 32'hc2697974, 32'h42c676ee, 32'h41c01567, 32'hbfc2e792};
test_output[15112:15119] = '{32'h410d22a5, 32'h42943032, 32'h424536b7, 32'h0, 32'h0, 32'h42c676ee, 32'h41c01567, 32'h0};
test_input[15120:15127] = '{32'h4147f76f, 32'h42a76b62, 32'h429e4c2f, 32'h4289481b, 32'hc25796d2, 32'hc1cce97a, 32'h42bd1d09, 32'hc2830a3c};
test_output[15120:15127] = '{32'h4147f76f, 32'h42a76b62, 32'h429e4c2f, 32'h4289481b, 32'h0, 32'h0, 32'h42bd1d09, 32'h0};
test_input[15128:15135] = '{32'hc20d7385, 32'hc0348f98, 32'h4287a69a, 32'hc2624283, 32'hc1da767b, 32'h42399b12, 32'hc129ddd5, 32'h4208a427};
test_output[15128:15135] = '{32'h0, 32'h0, 32'h4287a69a, 32'h0, 32'h0, 32'h42399b12, 32'h0, 32'h4208a427};
test_input[15136:15143] = '{32'hc270771b, 32'h421ff99a, 32'hc2a63cb5, 32'h4265c13e, 32'hc13ffcdc, 32'hc2c41bdc, 32'hc2c44d4b, 32'h42b8d20f};
test_output[15136:15143] = '{32'h0, 32'h421ff99a, 32'h0, 32'h4265c13e, 32'h0, 32'h0, 32'h0, 32'h42b8d20f};
test_input[15144:15151] = '{32'h42b9ea88, 32'hc0ee4253, 32'h427d5aa0, 32'hc22e13b5, 32'hc2b4b483, 32'h429e2a21, 32'hc1b4c1c6, 32'h42061e90};
test_output[15144:15151] = '{32'h42b9ea88, 32'h0, 32'h427d5aa0, 32'h0, 32'h0, 32'h429e2a21, 32'h0, 32'h42061e90};
test_input[15152:15159] = '{32'h42a2e55a, 32'h4255590f, 32'h41d536e6, 32'h4230640c, 32'h42a41216, 32'h42ad5c1d, 32'hc28dad1a, 32'hc2985401};
test_output[15152:15159] = '{32'h42a2e55a, 32'h4255590f, 32'h41d536e6, 32'h4230640c, 32'h42a41216, 32'h42ad5c1d, 32'h0, 32'h0};
test_input[15160:15167] = '{32'hc24166a5, 32'h4123e793, 32'hc2c39a1f, 32'h423b611c, 32'h42558276, 32'hc2954a2e, 32'hc20b6464, 32'h4212757c};
test_output[15160:15167] = '{32'h0, 32'h4123e793, 32'h0, 32'h423b611c, 32'h42558276, 32'h0, 32'h0, 32'h4212757c};
test_input[15168:15175] = '{32'hc25780cb, 32'hc2367c4e, 32'h4203f5ff, 32'hc1d1e312, 32'hc2c24a58, 32'h42c6ec6e, 32'h42809019, 32'h422ef969};
test_output[15168:15175] = '{32'h0, 32'h0, 32'h4203f5ff, 32'h0, 32'h0, 32'h42c6ec6e, 32'h42809019, 32'h422ef969};
test_input[15176:15183] = '{32'h429c858c, 32'hc2c69144, 32'hc1afe308, 32'hc22e8be8, 32'h41711bbd, 32'hc29ace33, 32'h41de437a, 32'hc26ad7c6};
test_output[15176:15183] = '{32'h429c858c, 32'h0, 32'h0, 32'h0, 32'h41711bbd, 32'h0, 32'h41de437a, 32'h0};
test_input[15184:15191] = '{32'h42c47d00, 32'hc1f39cf2, 32'hc0e61d8c, 32'hc254b8b9, 32'hc2b08440, 32'hc2740642, 32'h4267ef32, 32'h4244695e};
test_output[15184:15191] = '{32'h42c47d00, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4267ef32, 32'h4244695e};
test_input[15192:15199] = '{32'hc27fa49b, 32'h42626631, 32'h41dc68b7, 32'hc255eb47, 32'hc2b1fbf7, 32'hc26c6a91, 32'hc111f153, 32'h42b92dc8};
test_output[15192:15199] = '{32'h0, 32'h42626631, 32'h41dc68b7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b92dc8};
test_input[15200:15207] = '{32'h420f1d8e, 32'hc09d22b5, 32'h419a117b, 32'h42104cbf, 32'hc1e7706d, 32'h429e9a68, 32'hc2ad9cbb, 32'hc2842e48};
test_output[15200:15207] = '{32'h420f1d8e, 32'h0, 32'h419a117b, 32'h42104cbf, 32'h0, 32'h429e9a68, 32'h0, 32'h0};
test_input[15208:15215] = '{32'hc1c7a529, 32'hc201d5d7, 32'hc2b72340, 32'h40bca7c3, 32'h425ed706, 32'h42ae6fe4, 32'h425f419e, 32'h4083f196};
test_output[15208:15215] = '{32'h0, 32'h0, 32'h0, 32'h40bca7c3, 32'h425ed706, 32'h42ae6fe4, 32'h425f419e, 32'h4083f196};
test_input[15216:15223] = '{32'h41fa0239, 32'hc29509d4, 32'hc269b019, 32'h41d6b058, 32'h42c266a9, 32'h429dff18, 32'h41aec58a, 32'h429df350};
test_output[15216:15223] = '{32'h41fa0239, 32'h0, 32'h0, 32'h41d6b058, 32'h42c266a9, 32'h429dff18, 32'h41aec58a, 32'h429df350};
test_input[15224:15231] = '{32'h41c893c3, 32'hc1862944, 32'h4216fe85, 32'hc267ef90, 32'h4195685d, 32'hc2021acb, 32'h4280e8bf, 32'h416c741f};
test_output[15224:15231] = '{32'h41c893c3, 32'h0, 32'h4216fe85, 32'h0, 32'h4195685d, 32'h0, 32'h4280e8bf, 32'h416c741f};
test_input[15232:15239] = '{32'h4297775a, 32'h41af3bc3, 32'hc23b15af, 32'hc28810ee, 32'hc2759715, 32'hc2913a9d, 32'hc23afb27, 32'hc26ca4c0};
test_output[15232:15239] = '{32'h4297775a, 32'h41af3bc3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15240:15247] = '{32'hc28a026a, 32'hc1874055, 32'h42a06f95, 32'hc29d26f6, 32'h4181f582, 32'hc205dfda, 32'hc29a890a, 32'h41dd6919};
test_output[15240:15247] = '{32'h0, 32'h0, 32'h42a06f95, 32'h0, 32'h4181f582, 32'h0, 32'h0, 32'h41dd6919};
test_input[15248:15255] = '{32'hc1517dc0, 32'hc2965c04, 32'hc2c5e02d, 32'hc2936f27, 32'h42b8e356, 32'hc0b61198, 32'h420fa66d, 32'h4226ac9b};
test_output[15248:15255] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42b8e356, 32'h0, 32'h420fa66d, 32'h4226ac9b};
test_input[15256:15263] = '{32'hc21f4c6d, 32'hc04dfce0, 32'h4083bbb0, 32'h41f9266f, 32'h41ee5fe5, 32'h42720f44, 32'h418bec8d, 32'hc15869e4};
test_output[15256:15263] = '{32'h0, 32'h0, 32'h4083bbb0, 32'h41f9266f, 32'h41ee5fe5, 32'h42720f44, 32'h418bec8d, 32'h0};
test_input[15264:15271] = '{32'hc259742d, 32'h423d3ad0, 32'h4228c4d1, 32'h42baf2a4, 32'hc2464270, 32'hc0185b8c, 32'h418443c4, 32'h42928ba3};
test_output[15264:15271] = '{32'h0, 32'h423d3ad0, 32'h4228c4d1, 32'h42baf2a4, 32'h0, 32'h0, 32'h418443c4, 32'h42928ba3};
test_input[15272:15279] = '{32'hc2acd91c, 32'h4283b5b1, 32'hc2a665ec, 32'h426d3a8c, 32'h423c6a15, 32'h429dad0b, 32'h428cddee, 32'hc1f582f1};
test_output[15272:15279] = '{32'h0, 32'h4283b5b1, 32'h0, 32'h426d3a8c, 32'h423c6a15, 32'h429dad0b, 32'h428cddee, 32'h0};
test_input[15280:15287] = '{32'hc2bcd0ca, 32'h412a8cc6, 32'h42bb113c, 32'h421c77c6, 32'h414ddd99, 32'h42042d28, 32'h411210de, 32'h415e8c12};
test_output[15280:15287] = '{32'h0, 32'h412a8cc6, 32'h42bb113c, 32'h421c77c6, 32'h414ddd99, 32'h42042d28, 32'h411210de, 32'h415e8c12};
test_input[15288:15295] = '{32'h413eb73d, 32'h42ac0b20, 32'hc2107b1a, 32'hc19a007c, 32'hc2be30ed, 32'hc04cd499, 32'h426b55f4, 32'h41dc1e76};
test_output[15288:15295] = '{32'h413eb73d, 32'h42ac0b20, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426b55f4, 32'h41dc1e76};
test_input[15296:15303] = '{32'hc2c23525, 32'hc2b877fb, 32'h41437d7e, 32'h42ac7d28, 32'hc1099b89, 32'hc116ea31, 32'hc008c060, 32'hc1b87f2e};
test_output[15296:15303] = '{32'h0, 32'h0, 32'h41437d7e, 32'h42ac7d28, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15304:15311] = '{32'hc2a3b678, 32'h425ffb73, 32'hc29fbbdf, 32'hc22aae35, 32'h42ac29c7, 32'hc11edf03, 32'hc243340e, 32'hc2adbee3};
test_output[15304:15311] = '{32'h0, 32'h425ffb73, 32'h0, 32'h0, 32'h42ac29c7, 32'h0, 32'h0, 32'h0};
test_input[15312:15319] = '{32'hc2a5f9b3, 32'hc2b5f497, 32'hc26ce0a3, 32'h40980c91, 32'h4170627a, 32'h42bfe06d, 32'hc25558ab, 32'h4215f87f};
test_output[15312:15319] = '{32'h0, 32'h0, 32'h0, 32'h40980c91, 32'h4170627a, 32'h42bfe06d, 32'h0, 32'h4215f87f};
test_input[15320:15327] = '{32'hc21f9184, 32'h413d0d1b, 32'h423bc7f2, 32'hc1ec753d, 32'hc1c4284b, 32'h415a5005, 32'hc17e6bf1, 32'h428d09ad};
test_output[15320:15327] = '{32'h0, 32'h413d0d1b, 32'h423bc7f2, 32'h0, 32'h0, 32'h415a5005, 32'h0, 32'h428d09ad};
test_input[15328:15335] = '{32'hc27ad2f6, 32'hc27b2fa5, 32'h4215f254, 32'hc29a5d83, 32'h42549e3e, 32'hc1ffaf9c, 32'hc26be342, 32'h4233fde1};
test_output[15328:15335] = '{32'h0, 32'h0, 32'h4215f254, 32'h0, 32'h42549e3e, 32'h0, 32'h0, 32'h4233fde1};
test_input[15336:15343] = '{32'h426ff498, 32'hc0f93cc3, 32'hc16e38aa, 32'h42132727, 32'h42135a50, 32'hc22ad682, 32'h421a0d8d, 32'h42548fbc};
test_output[15336:15343] = '{32'h426ff498, 32'h0, 32'h0, 32'h42132727, 32'h42135a50, 32'h0, 32'h421a0d8d, 32'h42548fbc};
test_input[15344:15351] = '{32'h42a53053, 32'h41cd74c5, 32'h422778c3, 32'h41904ecd, 32'h42879c91, 32'h406a2c91, 32'hc2bd038b, 32'h42a9497d};
test_output[15344:15351] = '{32'h42a53053, 32'h41cd74c5, 32'h422778c3, 32'h41904ecd, 32'h42879c91, 32'h406a2c91, 32'h0, 32'h42a9497d};
test_input[15352:15359] = '{32'hc2837dca, 32'hc2c3339f, 32'hc25dfa03, 32'h42838389, 32'h4227a5e7, 32'h4259ff12, 32'hc2a634fd, 32'h42a1a668};
test_output[15352:15359] = '{32'h0, 32'h0, 32'h0, 32'h42838389, 32'h4227a5e7, 32'h4259ff12, 32'h0, 32'h42a1a668};
test_input[15360:15367] = '{32'h42c15880, 32'h4251e21d, 32'hc29a9a5f, 32'hc2303f00, 32'hc2884525, 32'hc25a7c23, 32'hc2aee055, 32'hc291978f};
test_output[15360:15367] = '{32'h42c15880, 32'h4251e21d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15368:15375] = '{32'h3ff78e80, 32'h424ad0bd, 32'h426283d6, 32'hc1e21bad, 32'hc2bf0061, 32'hc208b49f, 32'h423da8a1, 32'h41f8efbc};
test_output[15368:15375] = '{32'h3ff78e80, 32'h424ad0bd, 32'h426283d6, 32'h0, 32'h0, 32'h0, 32'h423da8a1, 32'h41f8efbc};
test_input[15376:15383] = '{32'hc17423f0, 32'h428012d5, 32'h41f6752d, 32'hc28ac207, 32'h4218bad3, 32'h4249fb22, 32'hc139d329, 32'h42bceffe};
test_output[15376:15383] = '{32'h0, 32'h428012d5, 32'h41f6752d, 32'h0, 32'h4218bad3, 32'h4249fb22, 32'h0, 32'h42bceffe};
test_input[15384:15391] = '{32'h40482e9b, 32'hc251aa2b, 32'h42c36823, 32'h41f6f41e, 32'hc2129fb4, 32'hc1bc6d53, 32'hc1a511f0, 32'hc21221ef};
test_output[15384:15391] = '{32'h40482e9b, 32'h0, 32'h42c36823, 32'h41f6f41e, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15392:15399] = '{32'h428be353, 32'hc1153ee0, 32'hc2c5d74f, 32'hc26e28bd, 32'h42a9e8bc, 32'hc1eb0179, 32'h423d70db, 32'h422dd280};
test_output[15392:15399] = '{32'h428be353, 32'h0, 32'h0, 32'h0, 32'h42a9e8bc, 32'h0, 32'h423d70db, 32'h422dd280};
test_input[15400:15407] = '{32'h42820638, 32'h427b778f, 32'h41c87148, 32'hc2b89a78, 32'h406b9249, 32'h42666810, 32'hc28dab2d, 32'h41fe347d};
test_output[15400:15407] = '{32'h42820638, 32'h427b778f, 32'h41c87148, 32'h0, 32'h406b9249, 32'h42666810, 32'h0, 32'h41fe347d};
test_input[15408:15415] = '{32'hc2b6d0d8, 32'hc1d7ef4a, 32'hc1f18e86, 32'hc2955a75, 32'hc287a7f1, 32'hc1172d9d, 32'h428e0d08, 32'hc2aa21a7};
test_output[15408:15415] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428e0d08, 32'h0};
test_input[15416:15423] = '{32'hc2c51183, 32'hc2bb09b4, 32'hc1d5566c, 32'hc24fcca6, 32'hc279ffba, 32'hc27c2c59, 32'h42534c9c, 32'h423411a2};
test_output[15416:15423] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42534c9c, 32'h423411a2};
test_input[15424:15431] = '{32'hc2322e7a, 32'hc1a65c85, 32'hc1c572dc, 32'h42935291, 32'hc204b855, 32'hc2a06c5b, 32'hc291bdb9, 32'hc19781e4};
test_output[15424:15431] = '{32'h0, 32'h0, 32'h0, 32'h42935291, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15432:15439] = '{32'h42216ee1, 32'hc18c33f9, 32'hc2960e8d, 32'hc1ce2a3f, 32'h403297c3, 32'hc23f55a9, 32'hc22d06f2, 32'h42acb86c};
test_output[15432:15439] = '{32'h42216ee1, 32'h0, 32'h0, 32'h0, 32'h403297c3, 32'h0, 32'h0, 32'h42acb86c};
test_input[15440:15447] = '{32'h41a75c4b, 32'hc1ac2020, 32'h42724eec, 32'hc2ab4f14, 32'hbf2d9d1f, 32'hc24c8253, 32'h429243f1, 32'h41d7209c};
test_output[15440:15447] = '{32'h41a75c4b, 32'h0, 32'h42724eec, 32'h0, 32'h0, 32'h0, 32'h429243f1, 32'h41d7209c};
test_input[15448:15455] = '{32'hc2432917, 32'h4122a05c, 32'hc2a4c607, 32'h41df074c, 32'hc14d8b4c, 32'h41cbaf1f, 32'hc12eb156, 32'h42b74eb9};
test_output[15448:15455] = '{32'h0, 32'h4122a05c, 32'h0, 32'h41df074c, 32'h0, 32'h41cbaf1f, 32'h0, 32'h42b74eb9};
test_input[15456:15463] = '{32'hc2a70e5f, 32'h428b40ad, 32'h4125fc11, 32'h3f8b9444, 32'h422cd743, 32'hbfc952e7, 32'hc1d7e8d4, 32'h42156ed5};
test_output[15456:15463] = '{32'h0, 32'h428b40ad, 32'h4125fc11, 32'h3f8b9444, 32'h422cd743, 32'h0, 32'h0, 32'h42156ed5};
test_input[15464:15471] = '{32'hc239aefd, 32'hc2aca0cc, 32'hc201556b, 32'h42035973, 32'hc218181f, 32'hc2a1b19e, 32'hc2008c2a, 32'h41a160d4};
test_output[15464:15471] = '{32'h0, 32'h0, 32'h0, 32'h42035973, 32'h0, 32'h0, 32'h0, 32'h41a160d4};
test_input[15472:15479] = '{32'h4278a5ca, 32'hc2b4728d, 32'hc1124707, 32'hc2c2ab83, 32'hc21bd235, 32'hc1d1e8da, 32'h4253a2a6, 32'hc283e1bb};
test_output[15472:15479] = '{32'h4278a5ca, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4253a2a6, 32'h0};
test_input[15480:15487] = '{32'hc1dbd7d5, 32'hc211e4c6, 32'h423bb69f, 32'hc14bf519, 32'hc2af4fad, 32'h42c0d005, 32'h42c014e5, 32'h4295e3b9};
test_output[15480:15487] = '{32'h0, 32'h0, 32'h423bb69f, 32'h0, 32'h0, 32'h42c0d005, 32'h42c014e5, 32'h4295e3b9};
test_input[15488:15495] = '{32'hc2212fbc, 32'hc1e6bea5, 32'hc2abf3ea, 32'h406a56a0, 32'hc2ac4453, 32'h428e059c, 32'h426f21dd, 32'hc10a9ae1};
test_output[15488:15495] = '{32'h0, 32'h0, 32'h0, 32'h406a56a0, 32'h0, 32'h428e059c, 32'h426f21dd, 32'h0};
test_input[15496:15503] = '{32'hc2a3c815, 32'h4299b1c2, 32'h4236ebb1, 32'hc06c6474, 32'h4237b451, 32'h41f4dacc, 32'h42068edd, 32'h424a3ea4};
test_output[15496:15503] = '{32'h0, 32'h4299b1c2, 32'h4236ebb1, 32'h0, 32'h4237b451, 32'h41f4dacc, 32'h42068edd, 32'h424a3ea4};
test_input[15504:15511] = '{32'h42133ab2, 32'hc1b0e5cb, 32'h42b88e51, 32'h3e304850, 32'h40c90c5c, 32'hc27d8f00, 32'hbf93744e, 32'h42856475};
test_output[15504:15511] = '{32'h42133ab2, 32'h0, 32'h42b88e51, 32'h3e304850, 32'h40c90c5c, 32'h0, 32'h0, 32'h42856475};
test_input[15512:15519] = '{32'h426d1410, 32'hc2aa122c, 32'h424aa1da, 32'hbf8c0397, 32'h418c52f5, 32'h41dfd213, 32'hc26db303, 32'hc1d40eee};
test_output[15512:15519] = '{32'h426d1410, 32'h0, 32'h424aa1da, 32'h0, 32'h418c52f5, 32'h41dfd213, 32'h0, 32'h0};
test_input[15520:15527] = '{32'h4201b7ad, 32'h3f1c3df4, 32'h409fc5b1, 32'hc12c71ea, 32'h420d9e7a, 32'h415d58b9, 32'hc241cda3, 32'hc242510d};
test_output[15520:15527] = '{32'h4201b7ad, 32'h3f1c3df4, 32'h409fc5b1, 32'h0, 32'h420d9e7a, 32'h415d58b9, 32'h0, 32'h0};
test_input[15528:15535] = '{32'h42a8b0ca, 32'hc1db0900, 32'hc28e6b6d, 32'hc29cbe35, 32'h41fe5afb, 32'hbf9d9844, 32'h41729e26, 32'hc0a2cb08};
test_output[15528:15535] = '{32'h42a8b0ca, 32'h0, 32'h0, 32'h0, 32'h41fe5afb, 32'h0, 32'h41729e26, 32'h0};
test_input[15536:15543] = '{32'h4296c4e4, 32'h4202f36f, 32'hc21c0b26, 32'hc281b07e, 32'h42b589b6, 32'hc211b7ae, 32'hc2ae9436, 32'hc21d19e1};
test_output[15536:15543] = '{32'h4296c4e4, 32'h4202f36f, 32'h0, 32'h0, 32'h42b589b6, 32'h0, 32'h0, 32'h0};
test_input[15544:15551] = '{32'hc1f01118, 32'hc291ced4, 32'hc18b42dd, 32'h4161d33e, 32'hc10c4916, 32'hc2288ae1, 32'h419d4d0c, 32'hc0daa0e2};
test_output[15544:15551] = '{32'h0, 32'h0, 32'h0, 32'h4161d33e, 32'h0, 32'h0, 32'h419d4d0c, 32'h0};
test_input[15552:15559] = '{32'hc19d985e, 32'hc1ea996b, 32'hc1be0d65, 32'h4217735e, 32'hc23ecb3c, 32'hc1a9b6f2, 32'hc28e8c75, 32'h422c8b4c};
test_output[15552:15559] = '{32'h0, 32'h0, 32'h0, 32'h4217735e, 32'h0, 32'h0, 32'h0, 32'h422c8b4c};
test_input[15560:15567] = '{32'h419b4c95, 32'hc2400c70, 32'hc1fe0fa5, 32'hc2927a34, 32'h422ae06c, 32'hc2b18686, 32'hc15c709b, 32'h425a7916};
test_output[15560:15567] = '{32'h419b4c95, 32'h0, 32'h0, 32'h0, 32'h422ae06c, 32'h0, 32'h0, 32'h425a7916};
test_input[15568:15575] = '{32'h407750cc, 32'h4284f9ca, 32'hc209c390, 32'h425e1cb6, 32'hc27ef91a, 32'h42a21d7c, 32'h42b086db, 32'h42c09e22};
test_output[15568:15575] = '{32'h407750cc, 32'h4284f9ca, 32'h0, 32'h425e1cb6, 32'h0, 32'h42a21d7c, 32'h42b086db, 32'h42c09e22};
test_input[15576:15583] = '{32'h4142d9df, 32'hc24d6151, 32'h42368cb3, 32'h420fd324, 32'h41a93d09, 32'h42aed4c9, 32'hc2561031, 32'hc287e29d};
test_output[15576:15583] = '{32'h4142d9df, 32'h0, 32'h42368cb3, 32'h420fd324, 32'h41a93d09, 32'h42aed4c9, 32'h0, 32'h0};
test_input[15584:15591] = '{32'h422f9a88, 32'h41d45056, 32'hc2240a45, 32'h403b6358, 32'h40b8ed06, 32'h42b7e569, 32'h42a52b90, 32'h4270d2ea};
test_output[15584:15591] = '{32'h422f9a88, 32'h41d45056, 32'h0, 32'h403b6358, 32'h40b8ed06, 32'h42b7e569, 32'h42a52b90, 32'h4270d2ea};
test_input[15592:15599] = '{32'hc0b65dd4, 32'hc19c7d7e, 32'h428a9ef7, 32'h42a5acc1, 32'h424bc447, 32'hc2a43de1, 32'hc29050d5, 32'h4259246a};
test_output[15592:15599] = '{32'h0, 32'h0, 32'h428a9ef7, 32'h42a5acc1, 32'h424bc447, 32'h0, 32'h0, 32'h4259246a};
test_input[15600:15607] = '{32'h42c50668, 32'hc0e00541, 32'h41af1770, 32'hc20cec78, 32'hc1ef5392, 32'hc216e30d, 32'h42b46ce2, 32'hc1b1fe3f};
test_output[15600:15607] = '{32'h42c50668, 32'h0, 32'h41af1770, 32'h0, 32'h0, 32'h0, 32'h42b46ce2, 32'h0};
test_input[15608:15615] = '{32'h42b5949f, 32'h420f4947, 32'h4291f9a7, 32'h427046e5, 32'hc24e629c, 32'h42a5aaf4, 32'hbf78ed72, 32'h42b3c6ab};
test_output[15608:15615] = '{32'h42b5949f, 32'h420f4947, 32'h4291f9a7, 32'h427046e5, 32'h0, 32'h42a5aaf4, 32'h0, 32'h42b3c6ab};
test_input[15616:15623] = '{32'h42412452, 32'hc2c0cb3a, 32'h3ef20501, 32'hc1b7c9c2, 32'h420742a3, 32'h41c95375, 32'hc1962f55, 32'h4126ec85};
test_output[15616:15623] = '{32'h42412452, 32'h0, 32'h3ef20501, 32'h0, 32'h420742a3, 32'h41c95375, 32'h0, 32'h4126ec85};
test_input[15624:15631] = '{32'hc0c7ec13, 32'h42c458e5, 32'h4223a275, 32'hc2a9e9e2, 32'hc21a0df2, 32'h42a1abe5, 32'h42b0789d, 32'h427ee28b};
test_output[15624:15631] = '{32'h0, 32'h42c458e5, 32'h4223a275, 32'h0, 32'h0, 32'h42a1abe5, 32'h42b0789d, 32'h427ee28b};
test_input[15632:15639] = '{32'hc2766685, 32'h42894814, 32'h42593b24, 32'hc2c0cb93, 32'hc241c798, 32'h424662c4, 32'hc1506a94, 32'h4139c31d};
test_output[15632:15639] = '{32'h0, 32'h42894814, 32'h42593b24, 32'h0, 32'h0, 32'h424662c4, 32'h0, 32'h4139c31d};
test_input[15640:15647] = '{32'h4290878e, 32'hc250bbf4, 32'hc29211d7, 32'h427ddc06, 32'hc221ae57, 32'h414f7256, 32'hc23fd428, 32'h4298304e};
test_output[15640:15647] = '{32'h4290878e, 32'h0, 32'h0, 32'h427ddc06, 32'h0, 32'h414f7256, 32'h0, 32'h4298304e};
test_input[15648:15655] = '{32'h41f46591, 32'hc256a370, 32'hc2a4b31a, 32'hc209bfb7, 32'h42890bbb, 32'hbe88bcf1, 32'hc2656283, 32'hc1e242ef};
test_output[15648:15655] = '{32'h41f46591, 32'h0, 32'h0, 32'h0, 32'h42890bbb, 32'h0, 32'h0, 32'h0};
test_input[15656:15663] = '{32'hc210e52a, 32'h4220e20b, 32'hc2b9d1e3, 32'h426f5ac1, 32'h4274d3ff, 32'h424cc1b0, 32'h4298d496, 32'hc112ae21};
test_output[15656:15663] = '{32'h0, 32'h4220e20b, 32'h0, 32'h426f5ac1, 32'h4274d3ff, 32'h424cc1b0, 32'h4298d496, 32'h0};
test_input[15664:15671] = '{32'hc2524c3c, 32'hc1d17aa9, 32'h421ffd20, 32'h423c9ed2, 32'h4298d24d, 32'h42ac576a, 32'h429b7517, 32'h41382aef};
test_output[15664:15671] = '{32'h0, 32'h0, 32'h421ffd20, 32'h423c9ed2, 32'h4298d24d, 32'h42ac576a, 32'h429b7517, 32'h41382aef};
test_input[15672:15679] = '{32'h426d130f, 32'hc1871e13, 32'h428349ae, 32'h4297b5c6, 32'hc2bf685b, 32'hc2a50843, 32'h429ba774, 32'hc21d9981};
test_output[15672:15679] = '{32'h426d130f, 32'h0, 32'h428349ae, 32'h4297b5c6, 32'h0, 32'h0, 32'h429ba774, 32'h0};
test_input[15680:15687] = '{32'h42540312, 32'h41e8fc16, 32'h42c18655, 32'h41a1d8ca, 32'hc25d625e, 32'hc2b73d54, 32'hc27da790, 32'h416a6abd};
test_output[15680:15687] = '{32'h42540312, 32'h41e8fc16, 32'h42c18655, 32'h41a1d8ca, 32'h0, 32'h0, 32'h0, 32'h416a6abd};
test_input[15688:15695] = '{32'hc191c752, 32'hc28f3aa3, 32'h41d0ad24, 32'h42525fb1, 32'h422d0fcf, 32'hc2c6facb, 32'h418535ef, 32'hc250e25e};
test_output[15688:15695] = '{32'h0, 32'h0, 32'h41d0ad24, 32'h42525fb1, 32'h422d0fcf, 32'h0, 32'h418535ef, 32'h0};
test_input[15696:15703] = '{32'h42042050, 32'h4203d9d1, 32'h417e9ad7, 32'h4266d5ca, 32'h41fa3cb3, 32'hc1d70fb3, 32'h406596e7, 32'hc2bd13a8};
test_output[15696:15703] = '{32'h42042050, 32'h4203d9d1, 32'h417e9ad7, 32'h4266d5ca, 32'h41fa3cb3, 32'h0, 32'h406596e7, 32'h0};
test_input[15704:15711] = '{32'hc0811f73, 32'h427ccd33, 32'hc2c00249, 32'h41d0dc9a, 32'hc1a8263e, 32'h42498294, 32'h416f8629, 32'hc2062bd9};
test_output[15704:15711] = '{32'h0, 32'h427ccd33, 32'h0, 32'h41d0dc9a, 32'h0, 32'h42498294, 32'h416f8629, 32'h0};
test_input[15712:15719] = '{32'hc2c79adc, 32'hc2c7234d, 32'hc226c04f, 32'h424fc5e6, 32'h42650372, 32'hc188d05f, 32'hc0d1379c, 32'hc2b7c2cf};
test_output[15712:15719] = '{32'h0, 32'h0, 32'h0, 32'h424fc5e6, 32'h42650372, 32'h0, 32'h0, 32'h0};
test_input[15720:15727] = '{32'h40fa3912, 32'h42abe85e, 32'h4299392e, 32'hc29a3922, 32'h41dc3572, 32'h41c54387, 32'h424699a2, 32'hc2080cd7};
test_output[15720:15727] = '{32'h40fa3912, 32'h42abe85e, 32'h4299392e, 32'h0, 32'h41dc3572, 32'h41c54387, 32'h424699a2, 32'h0};
test_input[15728:15735] = '{32'hc2ae010d, 32'h40ddf617, 32'h42116e20, 32'h42427833, 32'h42045ab9, 32'hc29c6263, 32'hbfe31d04, 32'hc22007bc};
test_output[15728:15735] = '{32'h0, 32'h40ddf617, 32'h42116e20, 32'h42427833, 32'h42045ab9, 32'h0, 32'h0, 32'h0};
test_input[15736:15743] = '{32'hc18e6b92, 32'h41deb05a, 32'h4115771e, 32'h42b62835, 32'hc0f748af, 32'hc28c7c26, 32'hc2a54219, 32'h42c0db04};
test_output[15736:15743] = '{32'h0, 32'h41deb05a, 32'h4115771e, 32'h42b62835, 32'h0, 32'h0, 32'h0, 32'h42c0db04};
test_input[15744:15751] = '{32'hc2473fc0, 32'h418c4f47, 32'hc21bfd37, 32'hc1f30172, 32'h41d30910, 32'hc2947b5d, 32'h41aa30ac, 32'h41f185ac};
test_output[15744:15751] = '{32'h0, 32'h418c4f47, 32'h0, 32'h0, 32'h41d30910, 32'h0, 32'h41aa30ac, 32'h41f185ac};
test_input[15752:15759] = '{32'h42616353, 32'h4263cec3, 32'hc21c024c, 32'h41692634, 32'h42269a55, 32'h40a08c74, 32'hc2948ce6, 32'h4195e647};
test_output[15752:15759] = '{32'h42616353, 32'h4263cec3, 32'h0, 32'h41692634, 32'h42269a55, 32'h40a08c74, 32'h0, 32'h4195e647};
test_input[15760:15767] = '{32'hc2b417cd, 32'hc2aef28e, 32'hc17a94da, 32'h41dc5572, 32'hc1b47e83, 32'hc25c7acb, 32'hc1e64703, 32'hc28270cc};
test_output[15760:15767] = '{32'h0, 32'h0, 32'h0, 32'h41dc5572, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15768:15775] = '{32'h42593934, 32'hc282be86, 32'h42afac4c, 32'hc235e7dc, 32'h421a2b59, 32'hc1d2d88f, 32'hc19ff761, 32'h42053588};
test_output[15768:15775] = '{32'h42593934, 32'h0, 32'h42afac4c, 32'h0, 32'h421a2b59, 32'h0, 32'h0, 32'h42053588};
test_input[15776:15783] = '{32'h420ecd0f, 32'h42076e58, 32'h42833a23, 32'h4297f1b1, 32'hc23a7fab, 32'h4016c757, 32'hc2608deb, 32'h420369de};
test_output[15776:15783] = '{32'h420ecd0f, 32'h42076e58, 32'h42833a23, 32'h4297f1b1, 32'h0, 32'h4016c757, 32'h0, 32'h420369de};
test_input[15784:15791] = '{32'h42bf6dbe, 32'hc1dc5c96, 32'hc1bbf53f, 32'hc2831098, 32'hc0a24ac1, 32'hc2944d77, 32'h4258a627, 32'h4286790c};
test_output[15784:15791] = '{32'h42bf6dbe, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4258a627, 32'h4286790c};
test_input[15792:15799] = '{32'h42a51d7b, 32'hc29c8c53, 32'h4288cebd, 32'h420d7331, 32'h4283520c, 32'h42a5f252, 32'hc2331c97, 32'h4273402e};
test_output[15792:15799] = '{32'h42a51d7b, 32'h0, 32'h4288cebd, 32'h420d7331, 32'h4283520c, 32'h42a5f252, 32'h0, 32'h4273402e};
test_input[15800:15807] = '{32'h4282efa6, 32'h42a1cff9, 32'hc2b36b90, 32'h42c70467, 32'hc25a2be1, 32'h421f7a28, 32'h423bc53f, 32'h419fa281};
test_output[15800:15807] = '{32'h4282efa6, 32'h42a1cff9, 32'h0, 32'h42c70467, 32'h0, 32'h421f7a28, 32'h423bc53f, 32'h419fa281};
test_input[15808:15815] = '{32'hc1856138, 32'h4200a00f, 32'h4281901e, 32'hc245ec09, 32'h42c633af, 32'hc283c9df, 32'h411c3593, 32'hc290c55b};
test_output[15808:15815] = '{32'h0, 32'h4200a00f, 32'h4281901e, 32'h0, 32'h42c633af, 32'h0, 32'h411c3593, 32'h0};
test_input[15816:15823] = '{32'h42af60b4, 32'h4103fecc, 32'h40fa1706, 32'h41ca7814, 32'hc15febdf, 32'hbe9087c7, 32'hc289d491, 32'hc2a03d85};
test_output[15816:15823] = '{32'h42af60b4, 32'h4103fecc, 32'h40fa1706, 32'h41ca7814, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15824:15831] = '{32'h429a0711, 32'hc288ce52, 32'h4270e5b4, 32'hc1ac7657, 32'h429d6a9a, 32'h400183d8, 32'hc21c9608, 32'hc2bcf10c};
test_output[15824:15831] = '{32'h429a0711, 32'h0, 32'h4270e5b4, 32'h0, 32'h429d6a9a, 32'h400183d8, 32'h0, 32'h0};
test_input[15832:15839] = '{32'h429a946d, 32'h421155a4, 32'h416ca402, 32'h415722f8, 32'h428e9fee, 32'hc1bbd7f8, 32'hc1830a4b, 32'hc1bdf956};
test_output[15832:15839] = '{32'h429a946d, 32'h421155a4, 32'h416ca402, 32'h415722f8, 32'h428e9fee, 32'h0, 32'h0, 32'h0};
test_input[15840:15847] = '{32'hc121c9ca, 32'hc2c2b6b2, 32'hc26ba658, 32'hc1fe5103, 32'hc157e83e, 32'h42086852, 32'hc22b992c, 32'h4209653f};
test_output[15840:15847] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42086852, 32'h0, 32'h4209653f};
test_input[15848:15855] = '{32'hc21b8a67, 32'hbf7c3017, 32'hc2c61411, 32'hc1c779db, 32'hc29c8c27, 32'h41af0dc0, 32'hc181b82b, 32'hc279cc17};
test_output[15848:15855] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41af0dc0, 32'h0, 32'h0};
test_input[15856:15863] = '{32'h40b46b4a, 32'hc296ec80, 32'hc050137c, 32'hc2c71577, 32'hc23e7a0d, 32'h42543a20, 32'hc2a1cf9c, 32'hc1f59cc9};
test_output[15856:15863] = '{32'h40b46b4a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42543a20, 32'h0, 32'h0};
test_input[15864:15871] = '{32'hc1941df1, 32'h42002ba4, 32'hc0377105, 32'h42c6f0e3, 32'hc1ed1aae, 32'h4287083e, 32'hc108c4f5, 32'hc10f5609};
test_output[15864:15871] = '{32'h0, 32'h42002ba4, 32'h0, 32'h42c6f0e3, 32'h0, 32'h4287083e, 32'h0, 32'h0};
test_input[15872:15879] = '{32'h420be175, 32'hc27bcb9b, 32'h42977f36, 32'hc110c82d, 32'h424b0e5e, 32'hc2b79ff6, 32'h4216466f, 32'h42b26deb};
test_output[15872:15879] = '{32'h420be175, 32'h0, 32'h42977f36, 32'h0, 32'h424b0e5e, 32'h0, 32'h4216466f, 32'h42b26deb};
test_input[15880:15887] = '{32'hc22ae272, 32'hc2a37ba9, 32'h424e4ec2, 32'h42417d7c, 32'hc2686e36, 32'hc1cd796b, 32'hc24b6721, 32'h410ccc15};
test_output[15880:15887] = '{32'h0, 32'h0, 32'h424e4ec2, 32'h42417d7c, 32'h0, 32'h0, 32'h0, 32'h410ccc15};
test_input[15888:15895] = '{32'h426833e6, 32'hc2394d0e, 32'hc2b4cc49, 32'hc2baf543, 32'hc299a84c, 32'hc2b62589, 32'hc29eda75, 32'hc239dd06};
test_output[15888:15895] = '{32'h426833e6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15896:15903] = '{32'hc219bf01, 32'h42a6051b, 32'hbffa30d7, 32'h42b3dc40, 32'h425de056, 32'h42b4899e, 32'hc1c500e2, 32'h419f8572};
test_output[15896:15903] = '{32'h0, 32'h42a6051b, 32'h0, 32'h42b3dc40, 32'h425de056, 32'h42b4899e, 32'h0, 32'h419f8572};
test_input[15904:15911] = '{32'hc26f0d2e, 32'hc1771f71, 32'h412c6290, 32'h42571cd6, 32'hc25d77d8, 32'h40b27900, 32'hc2171736, 32'h423e481f};
test_output[15904:15911] = '{32'h0, 32'h0, 32'h412c6290, 32'h42571cd6, 32'h0, 32'h40b27900, 32'h0, 32'h423e481f};
test_input[15912:15919] = '{32'h402d358c, 32'h42046644, 32'h4229bc70, 32'h417c9d8b, 32'h425cc4f7, 32'h42089351, 32'hc22ae152, 32'hc25ccd73};
test_output[15912:15919] = '{32'h402d358c, 32'h42046644, 32'h4229bc70, 32'h417c9d8b, 32'h425cc4f7, 32'h42089351, 32'h0, 32'h0};
test_input[15920:15927] = '{32'h41c0c5c6, 32'hc2a47a1d, 32'hc1dd52e2, 32'hc26344f1, 32'h41e6e630, 32'h4169690f, 32'hc2454767, 32'h41c94f5e};
test_output[15920:15927] = '{32'h41c0c5c6, 32'h0, 32'h0, 32'h0, 32'h41e6e630, 32'h4169690f, 32'h0, 32'h41c94f5e};
test_input[15928:15935] = '{32'h42a9d702, 32'h40029959, 32'h41aa5bfa, 32'h422eedcd, 32'h41409ad4, 32'hc1a6aa5a, 32'hc2c30ec9, 32'hc271fb37};
test_output[15928:15935] = '{32'h42a9d702, 32'h40029959, 32'h41aa5bfa, 32'h422eedcd, 32'h41409ad4, 32'h0, 32'h0, 32'h0};
test_input[15936:15943] = '{32'hc297dc69, 32'h4266e424, 32'hc260f044, 32'h42198814, 32'hc2130b34, 32'hc2c40b74, 32'hc27f3edb, 32'h416d0fd7};
test_output[15936:15943] = '{32'h0, 32'h4266e424, 32'h0, 32'h42198814, 32'h0, 32'h0, 32'h0, 32'h416d0fd7};
test_input[15944:15951] = '{32'h414b8abb, 32'h42a31a46, 32'h4271e12e, 32'h418aa35a, 32'hc2878690, 32'hc1d890f6, 32'h419eb01a, 32'h429023c1};
test_output[15944:15951] = '{32'h414b8abb, 32'h42a31a46, 32'h4271e12e, 32'h418aa35a, 32'h0, 32'h0, 32'h419eb01a, 32'h429023c1};
test_input[15952:15959] = '{32'hc28f5694, 32'h42bcfd2d, 32'hc0352bb8, 32'h4215ce96, 32'hc252d3d9, 32'h4257c6e5, 32'hc2165141, 32'hc26be50e};
test_output[15952:15959] = '{32'h0, 32'h42bcfd2d, 32'h0, 32'h4215ce96, 32'h0, 32'h4257c6e5, 32'h0, 32'h0};
test_input[15960:15967] = '{32'h41ad1fef, 32'h41fc7a10, 32'hc2c1b98c, 32'h42411f5f, 32'h41b46fcc, 32'h428458e7, 32'hc254bb82, 32'hc2c3e439};
test_output[15960:15967] = '{32'h41ad1fef, 32'h41fc7a10, 32'h0, 32'h42411f5f, 32'h41b46fcc, 32'h428458e7, 32'h0, 32'h0};
test_input[15968:15975] = '{32'h422c028e, 32'hc13d0cb9, 32'hc2375d7d, 32'h42938827, 32'h4223f62f, 32'hc2a2cf66, 32'hc2b2de13, 32'hc03a56cc};
test_output[15968:15975] = '{32'h422c028e, 32'h0, 32'h0, 32'h42938827, 32'h4223f62f, 32'h0, 32'h0, 32'h0};
test_input[15976:15983] = '{32'h4221f08b, 32'h41050be9, 32'h42256d03, 32'h42337ab2, 32'hc29624e4, 32'hc1d5ab40, 32'hc13235fe, 32'hc266c3a8};
test_output[15976:15983] = '{32'h4221f08b, 32'h41050be9, 32'h42256d03, 32'h42337ab2, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15984:15991] = '{32'h4295f1dd, 32'hc24bf8b1, 32'h4298236e, 32'h42b3376c, 32'hc2ae0de2, 32'hc270ebb0, 32'h41ba1418, 32'h400f4a41};
test_output[15984:15991] = '{32'h4295f1dd, 32'h0, 32'h4298236e, 32'h42b3376c, 32'h0, 32'h0, 32'h41ba1418, 32'h400f4a41};
test_input[15992:15999] = '{32'hc2a4c7a7, 32'hc29d9b87, 32'h42b1743e, 32'h41985779, 32'h42806953, 32'hc2a0ea86, 32'h41fe2006, 32'h42c113d2};
test_output[15992:15999] = '{32'h0, 32'h0, 32'h42b1743e, 32'h41985779, 32'h42806953, 32'h0, 32'h41fe2006, 32'h42c113d2};
test_input[16000:16007] = '{32'hc20e3fee, 32'h415748cf, 32'hbfbfb43f, 32'h41904a51, 32'h415b76be, 32'h41b21ae7, 32'h42b80681, 32'hc28814d5};
test_output[16000:16007] = '{32'h0, 32'h415748cf, 32'h0, 32'h41904a51, 32'h415b76be, 32'h41b21ae7, 32'h42b80681, 32'h0};
test_input[16008:16015] = '{32'h424b5a8e, 32'h41a3f9f1, 32'h4193d1eb, 32'hc2b979c5, 32'h420604ad, 32'hc2502a5e, 32'h4283ad10, 32'h4180c4a6};
test_output[16008:16015] = '{32'h424b5a8e, 32'h41a3f9f1, 32'h4193d1eb, 32'h0, 32'h420604ad, 32'h0, 32'h4283ad10, 32'h4180c4a6};
test_input[16016:16023] = '{32'h42544c38, 32'hc10bc89e, 32'h41d19a2e, 32'h420cebff, 32'hc169e9be, 32'h42906cfe, 32'h4284b3c3, 32'hc2a5c6cb};
test_output[16016:16023] = '{32'h42544c38, 32'h0, 32'h41d19a2e, 32'h420cebff, 32'h0, 32'h42906cfe, 32'h4284b3c3, 32'h0};
test_input[16024:16031] = '{32'h426261cf, 32'h420a795d, 32'hbf18864e, 32'h41883976, 32'h426649df, 32'hc249fb81, 32'h40f84db3, 32'hc21e03d9};
test_output[16024:16031] = '{32'h426261cf, 32'h420a795d, 32'h0, 32'h41883976, 32'h426649df, 32'h0, 32'h40f84db3, 32'h0};
test_input[16032:16039] = '{32'h4238ad88, 32'hc224ef97, 32'h41724fe8, 32'hc23210d6, 32'h423fffbc, 32'hc2b9069c, 32'hc2be3598, 32'hc28c3aa3};
test_output[16032:16039] = '{32'h4238ad88, 32'h0, 32'h41724fe8, 32'h0, 32'h423fffbc, 32'h0, 32'h0, 32'h0};
test_input[16040:16047] = '{32'h42136a53, 32'hc20831bc, 32'hc2959071, 32'hc28c02f0, 32'hc1a25efd, 32'hc0b83ca2, 32'h423beaad, 32'hc0afd42b};
test_output[16040:16047] = '{32'h42136a53, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423beaad, 32'h0};
test_input[16048:16055] = '{32'hc2ae5b2c, 32'h42b7c528, 32'h42032f1e, 32'h4205b378, 32'h42b9d382, 32'hc28ce000, 32'hc29cd28b, 32'hc2c1bd90};
test_output[16048:16055] = '{32'h0, 32'h42b7c528, 32'h42032f1e, 32'h4205b378, 32'h42b9d382, 32'h0, 32'h0, 32'h0};
test_input[16056:16063] = '{32'hc1efe9ba, 32'hc25329b1, 32'hc2a23673, 32'hc0e5f15d, 32'h4249d558, 32'hc1e8ee5f, 32'hc2b9668a, 32'h420c6a96};
test_output[16056:16063] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4249d558, 32'h0, 32'h0, 32'h420c6a96};
test_input[16064:16071] = '{32'hc28afb28, 32'hc250249e, 32'hc1293048, 32'h42972afb, 32'hc2aa36be, 32'h42a60756, 32'h42a63cf4, 32'h405d9800};
test_output[16064:16071] = '{32'h0, 32'h0, 32'h0, 32'h42972afb, 32'h0, 32'h42a60756, 32'h42a63cf4, 32'h405d9800};
test_input[16072:16079] = '{32'h429c5e13, 32'h41a01495, 32'h42ac1c26, 32'hc21a2c88, 32'h427425f4, 32'hc29dd3d7, 32'hc2914a3e, 32'h42467e22};
test_output[16072:16079] = '{32'h429c5e13, 32'h41a01495, 32'h42ac1c26, 32'h0, 32'h427425f4, 32'h0, 32'h0, 32'h42467e22};
test_input[16080:16087] = '{32'h42405894, 32'hbf9c1811, 32'hc227dba2, 32'h41b46490, 32'h41c91aa1, 32'h422f5ad3, 32'h3f0634c5, 32'h4253666a};
test_output[16080:16087] = '{32'h42405894, 32'h0, 32'h0, 32'h41b46490, 32'h41c91aa1, 32'h422f5ad3, 32'h3f0634c5, 32'h4253666a};
test_input[16088:16095] = '{32'h429a4e0d, 32'hc2c4fc0e, 32'hc1640a95, 32'hc2944bc0, 32'hc23e4c52, 32'hc29499c8, 32'hc28894b7, 32'h4206aa76};
test_output[16088:16095] = '{32'h429a4e0d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4206aa76};
test_input[16096:16103] = '{32'h3fd4c259, 32'h429c3e1f, 32'hc2a49729, 32'h42c3c66d, 32'hc0586a2d, 32'h4292bfc6, 32'hc29b41ef, 32'h425133d9};
test_output[16096:16103] = '{32'h3fd4c259, 32'h429c3e1f, 32'h0, 32'h42c3c66d, 32'h0, 32'h4292bfc6, 32'h0, 32'h425133d9};
test_input[16104:16111] = '{32'h42c20c36, 32'h4262ed00, 32'hc121fbeb, 32'hc2ac3724, 32'h42acf7cd, 32'h42a4ab2c, 32'h4280a818, 32'h41e0ec3f};
test_output[16104:16111] = '{32'h42c20c36, 32'h4262ed00, 32'h0, 32'h0, 32'h42acf7cd, 32'h42a4ab2c, 32'h4280a818, 32'h41e0ec3f};
test_input[16112:16119] = '{32'h4261c048, 32'h42ae3df2, 32'h4071408b, 32'hc1cde512, 32'hc246ecde, 32'hc295d51d, 32'hc130dfd9, 32'h41587dc0};
test_output[16112:16119] = '{32'h4261c048, 32'h42ae3df2, 32'h4071408b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41587dc0};
test_input[16120:16127] = '{32'h428ac8d2, 32'h42048e35, 32'h40f75707, 32'h42664e75, 32'hc10bd9ed, 32'h424fa7b5, 32'hc2bf06b6, 32'h4203bc58};
test_output[16120:16127] = '{32'h428ac8d2, 32'h42048e35, 32'h40f75707, 32'h42664e75, 32'h0, 32'h424fa7b5, 32'h0, 32'h4203bc58};
test_input[16128:16135] = '{32'h42b97b63, 32'hc2626faf, 32'hc225de30, 32'h42512075, 32'h426e554f, 32'h4225ccb8, 32'h42956f27, 32'h41cde9df};
test_output[16128:16135] = '{32'h42b97b63, 32'h0, 32'h0, 32'h42512075, 32'h426e554f, 32'h4225ccb8, 32'h42956f27, 32'h41cde9df};
test_input[16136:16143] = '{32'h42603ac8, 32'hc2718a27, 32'hc2bda371, 32'h429c6f9b, 32'h4201be1b, 32'h426aa6d5, 32'hc2a391da, 32'h4284bd7d};
test_output[16136:16143] = '{32'h42603ac8, 32'h0, 32'h0, 32'h429c6f9b, 32'h4201be1b, 32'h426aa6d5, 32'h0, 32'h4284bd7d};
test_input[16144:16151] = '{32'hc22a65db, 32'hc12031fe, 32'hc2296552, 32'hc19a49d6, 32'hc19d6830, 32'h4212bc6d, 32'hc1a097a0, 32'hc27d2a0d};
test_output[16144:16151] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4212bc6d, 32'h0, 32'h0};
test_input[16152:16159] = '{32'hc288caa8, 32'h427d4214, 32'hbf9fef56, 32'hc220c46b, 32'hc278aa33, 32'h40e17f61, 32'h4101889a, 32'hc277a1f1};
test_output[16152:16159] = '{32'h0, 32'h427d4214, 32'h0, 32'h0, 32'h0, 32'h40e17f61, 32'h4101889a, 32'h0};
test_input[16160:16167] = '{32'h42114b69, 32'hc24f8a6d, 32'h42c72c20, 32'hc23595d8, 32'h427e803f, 32'hc02653d9, 32'h427a94bf, 32'h421295a7};
test_output[16160:16167] = '{32'h42114b69, 32'h0, 32'h42c72c20, 32'h0, 32'h427e803f, 32'h0, 32'h427a94bf, 32'h421295a7};
test_input[16168:16175] = '{32'h428423cb, 32'hc28d442e, 32'h42a8f7b9, 32'h422c40c1, 32'h4251f863, 32'h413f2e07, 32'h41fa49ee, 32'h41615a9a};
test_output[16168:16175] = '{32'h428423cb, 32'h0, 32'h42a8f7b9, 32'h422c40c1, 32'h4251f863, 32'h413f2e07, 32'h41fa49ee, 32'h41615a9a};
test_input[16176:16183] = '{32'h40b5cca5, 32'hbfa6a5b4, 32'h42ada81a, 32'hc1b81b48, 32'hc2c5e996, 32'h4216e165, 32'hc256478a, 32'h428b4d40};
test_output[16176:16183] = '{32'h40b5cca5, 32'h0, 32'h42ada81a, 32'h0, 32'h0, 32'h4216e165, 32'h0, 32'h428b4d40};
test_input[16184:16191] = '{32'hc1d8a7a8, 32'hc28a506b, 32'h427553d3, 32'hc204f176, 32'h41971bc3, 32'h41fd3995, 32'hc11c5111, 32'hc228838b};
test_output[16184:16191] = '{32'h0, 32'h0, 32'h427553d3, 32'h0, 32'h41971bc3, 32'h41fd3995, 32'h0, 32'h0};
test_input[16192:16199] = '{32'h42b7bbe6, 32'hc2794f7a, 32'h42b8137e, 32'hc2448e81, 32'hc2a3c26d, 32'h41c3bf2c, 32'hc244baa6, 32'h428e1663};
test_output[16192:16199] = '{32'h42b7bbe6, 32'h0, 32'h42b8137e, 32'h0, 32'h0, 32'h41c3bf2c, 32'h0, 32'h428e1663};
test_input[16200:16207] = '{32'h42703d01, 32'h4285144f, 32'h421c56ce, 32'hc2858e6a, 32'hc118619f, 32'hc263bea3, 32'h41a33916, 32'hc25e57aa};
test_output[16200:16207] = '{32'h42703d01, 32'h4285144f, 32'h421c56ce, 32'h0, 32'h0, 32'h0, 32'h41a33916, 32'h0};
test_input[16208:16215] = '{32'hc20dddf0, 32'hc294247a, 32'hc2a25d81, 32'hc29e7415, 32'h42a11b34, 32'hc1ef7313, 32'h41a50d64, 32'h41af6ead};
test_output[16208:16215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a11b34, 32'h0, 32'h41a50d64, 32'h41af6ead};
test_input[16216:16223] = '{32'h429f7a08, 32'hc28d4cf3, 32'hc20fae84, 32'hc194ab5d, 32'h41cc7887, 32'h41c4cc33, 32'hc1aa0cb0, 32'h41b259de};
test_output[16216:16223] = '{32'h429f7a08, 32'h0, 32'h0, 32'h0, 32'h41cc7887, 32'h41c4cc33, 32'h0, 32'h41b259de};
test_input[16224:16231] = '{32'h4257b74a, 32'h413246df, 32'hc22dde09, 32'h416b2b71, 32'hc26d8027, 32'h4219db23, 32'hc28d2f2a, 32'hc1cfc6f9};
test_output[16224:16231] = '{32'h4257b74a, 32'h413246df, 32'h0, 32'h416b2b71, 32'h0, 32'h4219db23, 32'h0, 32'h0};
test_input[16232:16239] = '{32'h425fcdbd, 32'h42aa9b27, 32'hc0ee0ab1, 32'h41db9e58, 32'hc2c0cbc1, 32'h40c7372e, 32'h42193b2e, 32'h42472332};
test_output[16232:16239] = '{32'h425fcdbd, 32'h42aa9b27, 32'h0, 32'h41db9e58, 32'h0, 32'h40c7372e, 32'h42193b2e, 32'h42472332};
test_input[16240:16247] = '{32'hc287750d, 32'hc194b172, 32'hc275f12d, 32'hc2996b22, 32'h4242c14f, 32'h427b6f81, 32'h40b080be, 32'h42a127d3};
test_output[16240:16247] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4242c14f, 32'h427b6f81, 32'h40b080be, 32'h42a127d3};
test_input[16248:16255] = '{32'h42ba233b, 32'h422ed3cf, 32'h41f57596, 32'hc13c5f24, 32'hc1b2e0cb, 32'hc28a7bd8, 32'hc24a0eb3, 32'hc280a878};
test_output[16248:16255] = '{32'h42ba233b, 32'h422ed3cf, 32'h41f57596, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16256:16263] = '{32'h42b877d2, 32'hc1a5a53d, 32'h42a04b2a, 32'h42bbcd55, 32'h424aaeb4, 32'hc213c980, 32'hc2a68146, 32'hc2638b3d};
test_output[16256:16263] = '{32'h42b877d2, 32'h0, 32'h42a04b2a, 32'h42bbcd55, 32'h424aaeb4, 32'h0, 32'h0, 32'h0};
test_input[16264:16271] = '{32'hc2bda90c, 32'hc2a53dbd, 32'hc2c2543f, 32'h41359f4a, 32'hc112a983, 32'hc190d9df, 32'h4290cccb, 32'h422aab66};
test_output[16264:16271] = '{32'h0, 32'h0, 32'h0, 32'h41359f4a, 32'h0, 32'h0, 32'h4290cccb, 32'h422aab66};
test_input[16272:16279] = '{32'h41a492aa, 32'hc18a0893, 32'hc26e8225, 32'h406ec018, 32'hc27616e7, 32'hc1f50b36, 32'h42c57ec4, 32'hc22c0bf5};
test_output[16272:16279] = '{32'h41a492aa, 32'h0, 32'h0, 32'h406ec018, 32'h0, 32'h0, 32'h42c57ec4, 32'h0};
test_input[16280:16287] = '{32'hc2872c5f, 32'h402702f6, 32'h42a00872, 32'hc2ba9824, 32'h41d36f02, 32'h42222e24, 32'hc280b3e6, 32'h4278611c};
test_output[16280:16287] = '{32'h0, 32'h402702f6, 32'h42a00872, 32'h0, 32'h41d36f02, 32'h42222e24, 32'h0, 32'h4278611c};
test_input[16288:16295] = '{32'h42b19c4d, 32'hc21ecca6, 32'h40cd35f0, 32'h41cd26b9, 32'h429d1d43, 32'h41984515, 32'h42826409, 32'h40c18296};
test_output[16288:16295] = '{32'h42b19c4d, 32'h0, 32'h40cd35f0, 32'h41cd26b9, 32'h429d1d43, 32'h41984515, 32'h42826409, 32'h40c18296};
test_input[16296:16303] = '{32'h4220f9ac, 32'hc266a472, 32'h42b243a2, 32'hc28841b7, 32'hc2c5c89f, 32'hc2bbac77, 32'hc28d71f7, 32'hc114942c};
test_output[16296:16303] = '{32'h4220f9ac, 32'h0, 32'h42b243a2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16304:16311] = '{32'h4282c78b, 32'h42bab114, 32'h413c41e9, 32'h413fbb29, 32'hc2bf35b5, 32'hc1e82c50, 32'h41a71c1b, 32'hc21fa73f};
test_output[16304:16311] = '{32'h4282c78b, 32'h42bab114, 32'h413c41e9, 32'h413fbb29, 32'h0, 32'h0, 32'h41a71c1b, 32'h0};
test_input[16312:16319] = '{32'h4285f836, 32'hc292542a, 32'hc235957b, 32'h42552d98, 32'h42afadd4, 32'h419d1d16, 32'h429fcd75, 32'hc237cb1c};
test_output[16312:16319] = '{32'h4285f836, 32'h0, 32'h0, 32'h42552d98, 32'h42afadd4, 32'h419d1d16, 32'h429fcd75, 32'h0};
test_input[16320:16327] = '{32'hc2a53d86, 32'hc1cfe57b, 32'hc193fc8b, 32'hc1aff47d, 32'hc2965283, 32'hc2b2c035, 32'hc2a19f44, 32'h4241a6ae};
test_output[16320:16327] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4241a6ae};
test_input[16328:16335] = '{32'h42b49b17, 32'h42154abf, 32'h427524d8, 32'h424846ca, 32'hc1398ab5, 32'hc290d6cc, 32'h424f9130, 32'h42bf8452};
test_output[16328:16335] = '{32'h42b49b17, 32'h42154abf, 32'h427524d8, 32'h424846ca, 32'h0, 32'h0, 32'h424f9130, 32'h42bf8452};
test_input[16336:16343] = '{32'h4287b58e, 32'h42093d88, 32'hc24356cb, 32'h425300d0, 32'hc1edcccc, 32'h42998c5d, 32'h40c98643, 32'h427bde8a};
test_output[16336:16343] = '{32'h4287b58e, 32'h42093d88, 32'h0, 32'h425300d0, 32'h0, 32'h42998c5d, 32'h40c98643, 32'h427bde8a};
test_input[16344:16351] = '{32'h42095c48, 32'h4293a476, 32'hc29328a3, 32'hc279a881, 32'h423158db, 32'hc2752625, 32'hc19c09aa, 32'hc16f85b7};
test_output[16344:16351] = '{32'h42095c48, 32'h4293a476, 32'h0, 32'h0, 32'h423158db, 32'h0, 32'h0, 32'h0};
test_input[16352:16359] = '{32'h42868dab, 32'hc2b06514, 32'h418ce2a1, 32'h4272e70b, 32'hc15e1901, 32'hc267dedf, 32'h4288d0e0, 32'h427f3fd7};
test_output[16352:16359] = '{32'h42868dab, 32'h0, 32'h418ce2a1, 32'h4272e70b, 32'h0, 32'h0, 32'h4288d0e0, 32'h427f3fd7};
test_input[16360:16367] = '{32'hc29d5e70, 32'h423f8cf3, 32'hc1b14c44, 32'hc2b789ff, 32'hc266b117, 32'hc2828ba5, 32'h42ac0b99, 32'h3f727b7b};
test_output[16360:16367] = '{32'h0, 32'h423f8cf3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ac0b99, 32'h3f727b7b};
test_input[16368:16375] = '{32'hc2955b5e, 32'h42b5090c, 32'h41854c94, 32'h41824aab, 32'h42b6eb56, 32'hc25c3342, 32'hbfcd7f19, 32'h40fd6d69};
test_output[16368:16375] = '{32'h0, 32'h42b5090c, 32'h41854c94, 32'h41824aab, 32'h42b6eb56, 32'h0, 32'h0, 32'h40fd6d69};
test_input[16376:16383] = '{32'hc21df288, 32'h41748780, 32'h42294dc8, 32'h42b7ba55, 32'hc16cb069, 32'hc2a9b572, 32'h42c5b4d4, 32'hc18f586a};
test_output[16376:16383] = '{32'h0, 32'h41748780, 32'h42294dc8, 32'h42b7ba55, 32'h0, 32'h0, 32'h42c5b4d4, 32'h0};
test_input[16384:16391] = '{32'h418485cf, 32'h4256a6d6, 32'hc1960902, 32'hc25081cb, 32'h429a078e, 32'h3ff232de, 32'hc1c97895, 32'h4281189e};
test_output[16384:16391] = '{32'h418485cf, 32'h4256a6d6, 32'h0, 32'h0, 32'h429a078e, 32'h3ff232de, 32'h0, 32'h4281189e};
test_input[16392:16399] = '{32'hc2abca78, 32'hc27b2a8e, 32'hc1b4b480, 32'hc2b967a9, 32'hc1247cc8, 32'h4247d2c7, 32'h42be3a4d, 32'hc181fe7e};
test_output[16392:16399] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4247d2c7, 32'h42be3a4d, 32'h0};
test_input[16400:16407] = '{32'hc29ca51c, 32'h42c0a14a, 32'hc2a279d5, 32'hc1e54509, 32'h4147725d, 32'hc1e9f8ec, 32'h423f0594, 32'hc2943914};
test_output[16400:16407] = '{32'h0, 32'h42c0a14a, 32'h0, 32'h0, 32'h4147725d, 32'h0, 32'h423f0594, 32'h0};
test_input[16408:16415] = '{32'h41b5d953, 32'h41dc9866, 32'h418fefaa, 32'h41b40751, 32'h420a3462, 32'hc2b46ba7, 32'hc1df1529, 32'hc22f3db3};
test_output[16408:16415] = '{32'h41b5d953, 32'h41dc9866, 32'h418fefaa, 32'h41b40751, 32'h420a3462, 32'h0, 32'h0, 32'h0};
test_input[16416:16423] = '{32'h42117725, 32'hc210b2d4, 32'h407e726d, 32'h42ba4b2c, 32'h424644e5, 32'h422691a8, 32'hc2b654ee, 32'hc2297a73};
test_output[16416:16423] = '{32'h42117725, 32'h0, 32'h407e726d, 32'h42ba4b2c, 32'h424644e5, 32'h422691a8, 32'h0, 32'h0};
test_input[16424:16431] = '{32'hc2b41172, 32'hc283ece4, 32'hbf8a571f, 32'h42b0d7ee, 32'h3fea8bc1, 32'hc28b8ac7, 32'h42b2a5f0, 32'h401be33a};
test_output[16424:16431] = '{32'h0, 32'h0, 32'h0, 32'h42b0d7ee, 32'h3fea8bc1, 32'h0, 32'h42b2a5f0, 32'h401be33a};
test_input[16432:16439] = '{32'hc0819ae9, 32'h41d7a47f, 32'hc17c2433, 32'hc0d00176, 32'h422bf77a, 32'h42b8a5c3, 32'hc2c4c5a9, 32'hc2285dcc};
test_output[16432:16439] = '{32'h0, 32'h41d7a47f, 32'h0, 32'h0, 32'h422bf77a, 32'h42b8a5c3, 32'h0, 32'h0};
test_input[16440:16447] = '{32'h42969e61, 32'h41a1524d, 32'h42c6e076, 32'hc18cee03, 32'hc25cddca, 32'hc22f1c6d, 32'hc1cff03d, 32'hc2828d4d};
test_output[16440:16447] = '{32'h42969e61, 32'h41a1524d, 32'h42c6e076, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16448:16455] = '{32'h42379ad5, 32'hc2973350, 32'hc2805883, 32'hc21fa7ba, 32'hc1211d2f, 32'hc116d440, 32'h42826d5e, 32'h429558eb};
test_output[16448:16455] = '{32'h42379ad5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42826d5e, 32'h429558eb};
test_input[16456:16463] = '{32'h4048d998, 32'hc29963f7, 32'hc2a13ba5, 32'hc1cae370, 32'hc2030b74, 32'hc22a7956, 32'h41965411, 32'hc1d597ba};
test_output[16456:16463] = '{32'h4048d998, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41965411, 32'h0};
test_input[16464:16471] = '{32'h42c7dc64, 32'hc2b472a2, 32'hc0f56af1, 32'hc2bd5d64, 32'h425202dd, 32'h42785220, 32'h4243ff53, 32'h4270d210};
test_output[16464:16471] = '{32'h42c7dc64, 32'h0, 32'h0, 32'h0, 32'h425202dd, 32'h42785220, 32'h4243ff53, 32'h4270d210};
test_input[16472:16479] = '{32'hc2b195dd, 32'h42088c78, 32'h42188b75, 32'h415b1791, 32'h4183e2d0, 32'hc2b270c5, 32'hc156ec7e, 32'h428dbbb7};
test_output[16472:16479] = '{32'h0, 32'h42088c78, 32'h42188b75, 32'h415b1791, 32'h4183e2d0, 32'h0, 32'h0, 32'h428dbbb7};
test_input[16480:16487] = '{32'hc1993b34, 32'h41ee0bff, 32'h4243e24c, 32'hc2a16c93, 32'hc1ff7f51, 32'hc25db11c, 32'h41a486c6, 32'hc29b23f3};
test_output[16480:16487] = '{32'h0, 32'h41ee0bff, 32'h4243e24c, 32'h0, 32'h0, 32'h0, 32'h41a486c6, 32'h0};
test_input[16488:16495] = '{32'h41bdc0c3, 32'h42305729, 32'hc2ae82e8, 32'hbf56722d, 32'h42b123f6, 32'hc1fae604, 32'h42895003, 32'hc06c1fec};
test_output[16488:16495] = '{32'h41bdc0c3, 32'h42305729, 32'h0, 32'h0, 32'h42b123f6, 32'h0, 32'h42895003, 32'h0};
test_input[16496:16503] = '{32'h426f1770, 32'h4142efe5, 32'h41e8f7d0, 32'h42371ded, 32'h42c6eaef, 32'hc287a93b, 32'h429bf9de, 32'hc25f810a};
test_output[16496:16503] = '{32'h426f1770, 32'h4142efe5, 32'h41e8f7d0, 32'h42371ded, 32'h42c6eaef, 32'h0, 32'h429bf9de, 32'h0};
test_input[16504:16511] = '{32'h429bd318, 32'hc2c35353, 32'h42832dee, 32'h4222b3d7, 32'hc1d8eabd, 32'h42905744, 32'hc2a5034b, 32'hc18a2333};
test_output[16504:16511] = '{32'h429bd318, 32'h0, 32'h42832dee, 32'h4222b3d7, 32'h0, 32'h42905744, 32'h0, 32'h0};
test_input[16512:16519] = '{32'hc24285ff, 32'h429d03ef, 32'h41aac222, 32'hc2628c38, 32'h42c491a5, 32'h414e8f4e, 32'h427bc584, 32'hc20bcd4c};
test_output[16512:16519] = '{32'h0, 32'h429d03ef, 32'h41aac222, 32'h0, 32'h42c491a5, 32'h414e8f4e, 32'h427bc584, 32'h0};
test_input[16520:16527] = '{32'hc28bba0a, 32'h42182251, 32'h41475162, 32'hc25d3679, 32'hc28f153f, 32'hc255aeca, 32'h422dcdaa, 32'hc17387e6};
test_output[16520:16527] = '{32'h0, 32'h42182251, 32'h41475162, 32'h0, 32'h0, 32'h0, 32'h422dcdaa, 32'h0};
test_input[16528:16535] = '{32'hc26de4e0, 32'h4261239b, 32'hc29d5858, 32'h425d21ee, 32'hc2b140ee, 32'h426103e4, 32'h418af4a3, 32'hc1bdb030};
test_output[16528:16535] = '{32'h0, 32'h4261239b, 32'h0, 32'h425d21ee, 32'h0, 32'h426103e4, 32'h418af4a3, 32'h0};
test_input[16536:16543] = '{32'hc22aa14d, 32'h416809e8, 32'h411391af, 32'h42b7b82c, 32'hc1c3f4d7, 32'h427096ff, 32'h41ce66f1, 32'h42b3f3a0};
test_output[16536:16543] = '{32'h0, 32'h416809e8, 32'h411391af, 32'h42b7b82c, 32'h0, 32'h427096ff, 32'h41ce66f1, 32'h42b3f3a0};
test_input[16544:16551] = '{32'h42bab7a2, 32'hc09656e6, 32'hc2a44dc2, 32'hc14fe644, 32'hc2acc347, 32'h41edab7a, 32'hc159967d, 32'hc17442aa};
test_output[16544:16551] = '{32'h42bab7a2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41edab7a, 32'h0, 32'h0};
test_input[16552:16559] = '{32'h42120c44, 32'h41ba1bf5, 32'h42c4283a, 32'h4220dc7c, 32'hc2013b5e, 32'h40120185, 32'hc25242aa, 32'hc24b29de};
test_output[16552:16559] = '{32'h42120c44, 32'h41ba1bf5, 32'h42c4283a, 32'h4220dc7c, 32'h0, 32'h40120185, 32'h0, 32'h0};
test_input[16560:16567] = '{32'h41013ab8, 32'hc2c1973d, 32'h410bd7f2, 32'h4285573b, 32'h42b693a9, 32'hc281bcbd, 32'hc2414ddc, 32'hc00a137b};
test_output[16560:16567] = '{32'h41013ab8, 32'h0, 32'h410bd7f2, 32'h4285573b, 32'h42b693a9, 32'h0, 32'h0, 32'h0};
test_input[16568:16575] = '{32'h41a98f49, 32'h424964b5, 32'h41e270f9, 32'h429bccd6, 32'h411ba8cf, 32'hc2b78746, 32'h42bda654, 32'hc280fc12};
test_output[16568:16575] = '{32'h41a98f49, 32'h424964b5, 32'h41e270f9, 32'h429bccd6, 32'h411ba8cf, 32'h0, 32'h42bda654, 32'h0};
test_input[16576:16583] = '{32'h4294ebc8, 32'h42343be1, 32'hc1b875d4, 32'hc29275ae, 32'h4285d4ff, 32'hc2b383ed, 32'hc1ef81b4, 32'hc12a4d82};
test_output[16576:16583] = '{32'h4294ebc8, 32'h42343be1, 32'h0, 32'h0, 32'h4285d4ff, 32'h0, 32'h0, 32'h0};
test_input[16584:16591] = '{32'h41f9bb4e, 32'h420d5389, 32'h42a8d050, 32'hbeb9732c, 32'h411028bb, 32'h41dc034b, 32'hc28b8092, 32'hc21a2f4a};
test_output[16584:16591] = '{32'h41f9bb4e, 32'h420d5389, 32'h42a8d050, 32'h0, 32'h411028bb, 32'h41dc034b, 32'h0, 32'h0};
test_input[16592:16599] = '{32'hc25e271c, 32'hc23b7242, 32'hc2704183, 32'hc11e2ea7, 32'h40a46e00, 32'hc28750de, 32'hc1e79f93, 32'h4190a0a2};
test_output[16592:16599] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40a46e00, 32'h0, 32'h0, 32'h4190a0a2};
test_input[16600:16607] = '{32'h4297e11f, 32'hc24d5afd, 32'hc0d41b48, 32'h4181c196, 32'h409dced2, 32'hc298a50b, 32'h4144a2b3, 32'h422ba4d5};
test_output[16600:16607] = '{32'h4297e11f, 32'h0, 32'h0, 32'h4181c196, 32'h409dced2, 32'h0, 32'h4144a2b3, 32'h422ba4d5};
test_input[16608:16615] = '{32'hc2b55ae8, 32'hc28e6009, 32'h40830ea4, 32'hc28e097e, 32'hc156350a, 32'h429fab8f, 32'hc2232e3d, 32'hc2b7c600};
test_output[16608:16615] = '{32'h0, 32'h0, 32'h40830ea4, 32'h0, 32'h0, 32'h429fab8f, 32'h0, 32'h0};
test_input[16616:16623] = '{32'hc22a0417, 32'hc1cccddf, 32'hc2af4ee5, 32'h42b67e65, 32'hc2b42ec6, 32'h4296d4ad, 32'h428b785a, 32'hc29f256a};
test_output[16616:16623] = '{32'h0, 32'h0, 32'h0, 32'h42b67e65, 32'h0, 32'h4296d4ad, 32'h428b785a, 32'h0};
test_input[16624:16631] = '{32'h428b65a3, 32'h42b0f0b0, 32'h42943583, 32'h41662e61, 32'h4167157f, 32'hc2633ebe, 32'h423ec4af, 32'hc2c5f88c};
test_output[16624:16631] = '{32'h428b65a3, 32'h42b0f0b0, 32'h42943583, 32'h41662e61, 32'h4167157f, 32'h0, 32'h423ec4af, 32'h0};
test_input[16632:16639] = '{32'h42bf246f, 32'hc280dfa2, 32'hc274d5c5, 32'hc297b3d4, 32'h408b358d, 32'hc1e679cb, 32'hc29ada13, 32'hc21d305e};
test_output[16632:16639] = '{32'h42bf246f, 32'h0, 32'h0, 32'h0, 32'h408b358d, 32'h0, 32'h0, 32'h0};
test_input[16640:16647] = '{32'h42af064b, 32'h42b00c55, 32'h42404e42, 32'h42853b97, 32'hc1c4eb45, 32'hc1f4428a, 32'h424a3c1a, 32'h42bc0faa};
test_output[16640:16647] = '{32'h42af064b, 32'h42b00c55, 32'h42404e42, 32'h42853b97, 32'h0, 32'h0, 32'h424a3c1a, 32'h42bc0faa};
test_input[16648:16655] = '{32'hc0fa3d6a, 32'h416ac486, 32'hbfd12159, 32'h419dfc80, 32'h422ce682, 32'hc23e361e, 32'h422ac545, 32'h4197360c};
test_output[16648:16655] = '{32'h0, 32'h416ac486, 32'h0, 32'h419dfc80, 32'h422ce682, 32'h0, 32'h422ac545, 32'h4197360c};
test_input[16656:16663] = '{32'hc21b6716, 32'h42b913cd, 32'h3ebabd7a, 32'hc29d56e9, 32'hc2933118, 32'h42998d61, 32'h40fa9833, 32'hc2a13e99};
test_output[16656:16663] = '{32'h0, 32'h42b913cd, 32'h3ebabd7a, 32'h0, 32'h0, 32'h42998d61, 32'h40fa9833, 32'h0};
test_input[16664:16671] = '{32'hbfb42dfc, 32'h42c15211, 32'h42a83272, 32'h42c5a864, 32'hc1915f1f, 32'hc264607b, 32'hc21e0868, 32'hbefe53cd};
test_output[16664:16671] = '{32'h0, 32'h42c15211, 32'h42a83272, 32'h42c5a864, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16672:16679] = '{32'hc2a91323, 32'hc2a80bf1, 32'h42bde4ec, 32'h42a52bbd, 32'hc2902832, 32'hc1678fd9, 32'hc1efae20, 32'hc2130031};
test_output[16672:16679] = '{32'h0, 32'h0, 32'h42bde4ec, 32'h42a52bbd, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16680:16687] = '{32'hc2a3b63c, 32'h42a2794b, 32'hc1004620, 32'hc2ad09c0, 32'h418e3710, 32'h42928a3b, 32'hc261ad4a, 32'h418d694b};
test_output[16680:16687] = '{32'h0, 32'h42a2794b, 32'h0, 32'h0, 32'h418e3710, 32'h42928a3b, 32'h0, 32'h418d694b};
test_input[16688:16695] = '{32'h411347db, 32'h3fe47bdb, 32'hc04bd0eb, 32'hc283bd99, 32'h4294f17d, 32'hc22fdf78, 32'hc2378cc9, 32'h41f3d018};
test_output[16688:16695] = '{32'h411347db, 32'h3fe47bdb, 32'h0, 32'h0, 32'h4294f17d, 32'h0, 32'h0, 32'h41f3d018};
test_input[16696:16703] = '{32'hc230c2d5, 32'hc28842e1, 32'hc2afcb2f, 32'hc1319f59, 32'hc0065de4, 32'hc2924945, 32'hc25854ef, 32'hc14649df};
test_output[16696:16703] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16704:16711] = '{32'hc2458eaa, 32'h429620cf, 32'hbfbece85, 32'hbfd5985d, 32'h426cb004, 32'h41fb07ed, 32'h4261c107, 32'h42bdf4ce};
test_output[16704:16711] = '{32'h0, 32'h429620cf, 32'h0, 32'h0, 32'h426cb004, 32'h41fb07ed, 32'h4261c107, 32'h42bdf4ce};
test_input[16712:16719] = '{32'h4289baca, 32'h4213656e, 32'h41d9b929, 32'hc1c83c42, 32'h42425b94, 32'h42bb2825, 32'h4281c270, 32'h427cff81};
test_output[16712:16719] = '{32'h4289baca, 32'h4213656e, 32'h41d9b929, 32'h0, 32'h42425b94, 32'h42bb2825, 32'h4281c270, 32'h427cff81};
test_input[16720:16727] = '{32'h42722bd0, 32'hc10ac928, 32'hc1ad31e3, 32'hc22cbf8e, 32'h42a90c4e, 32'hc167460c, 32'hc19caa7d, 32'hc25098e8};
test_output[16720:16727] = '{32'h42722bd0, 32'h0, 32'h0, 32'h0, 32'h42a90c4e, 32'h0, 32'h0, 32'h0};
test_input[16728:16735] = '{32'hc28b8a0e, 32'h418e61d8, 32'h420f2a76, 32'h418f2242, 32'hc094681d, 32'hc2a5d9bb, 32'hc0cad88b, 32'hbf883b0d};
test_output[16728:16735] = '{32'h0, 32'h418e61d8, 32'h420f2a76, 32'h418f2242, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16736:16743] = '{32'hc1c8172a, 32'h42c1afcd, 32'hc0644044, 32'hc27a77ea, 32'hc1d6eab3, 32'h424d6374, 32'hc01d5ede, 32'h4276fb74};
test_output[16736:16743] = '{32'h0, 32'h42c1afcd, 32'h0, 32'h0, 32'h0, 32'h424d6374, 32'h0, 32'h4276fb74};
test_input[16744:16751] = '{32'h42ad71e1, 32'h412a6a3b, 32'h413e1c77, 32'h42b102ad, 32'hc288cb46, 32'h4211f76a, 32'hc14a733e, 32'hc18affcc};
test_output[16744:16751] = '{32'h42ad71e1, 32'h412a6a3b, 32'h413e1c77, 32'h42b102ad, 32'h0, 32'h4211f76a, 32'h0, 32'h0};
test_input[16752:16759] = '{32'h42851e53, 32'h429cf723, 32'hc15ab5dc, 32'hc28be55a, 32'h424c783d, 32'hc28e6940, 32'hc2b14ced, 32'h418ef6bd};
test_output[16752:16759] = '{32'h42851e53, 32'h429cf723, 32'h0, 32'h0, 32'h424c783d, 32'h0, 32'h0, 32'h418ef6bd};
test_input[16760:16767] = '{32'hc1aae859, 32'hc2a0134c, 32'hc2a8d819, 32'h40e2e590, 32'hc2c739b5, 32'hc2b3e07c, 32'h42c10a08, 32'hc295f01b};
test_output[16760:16767] = '{32'h0, 32'h0, 32'h0, 32'h40e2e590, 32'h0, 32'h0, 32'h42c10a08, 32'h0};
test_input[16768:16775] = '{32'hc1fc774e, 32'hc29c4f19, 32'h4217ec47, 32'hc28ba340, 32'hc007f48e, 32'hc2a20203, 32'hc2969343, 32'h4241d819};
test_output[16768:16775] = '{32'h0, 32'h0, 32'h4217ec47, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4241d819};
test_input[16776:16783] = '{32'hbf645f59, 32'h425a3cd1, 32'hc18760a3, 32'hc14acd96, 32'h428f90e1, 32'h428c1b4f, 32'h420b73e5, 32'hc2bcf4bb};
test_output[16776:16783] = '{32'h0, 32'h425a3cd1, 32'h0, 32'h0, 32'h428f90e1, 32'h428c1b4f, 32'h420b73e5, 32'h0};
test_input[16784:16791] = '{32'h42ba7fc6, 32'hc25285cf, 32'h4107cf0c, 32'h42beff96, 32'hc278cd84, 32'h4247bb90, 32'h429b7d43, 32'h4267586f};
test_output[16784:16791] = '{32'h42ba7fc6, 32'h0, 32'h4107cf0c, 32'h42beff96, 32'h0, 32'h4247bb90, 32'h429b7d43, 32'h4267586f};
test_input[16792:16799] = '{32'h423dd9ce, 32'hc2c76ff4, 32'h42c4e797, 32'h40929cea, 32'hc2557c4a, 32'h429ea725, 32'hc24a4fc0, 32'h41901e14};
test_output[16792:16799] = '{32'h423dd9ce, 32'h0, 32'h42c4e797, 32'h40929cea, 32'h0, 32'h429ea725, 32'h0, 32'h41901e14};
test_input[16800:16807] = '{32'h41d4dc48, 32'hc2726630, 32'h4284cf32, 32'h413eedcf, 32'hc2523b1c, 32'h41930254, 32'hc1d89044, 32'h405658d7};
test_output[16800:16807] = '{32'h41d4dc48, 32'h0, 32'h4284cf32, 32'h413eedcf, 32'h0, 32'h41930254, 32'h0, 32'h405658d7};
test_input[16808:16815] = '{32'hc26ada6f, 32'hc26de631, 32'hc2846db7, 32'hc191ba64, 32'h42122d91, 32'h4299fbb5, 32'h4185fd43, 32'hc19b5d7f};
test_output[16808:16815] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42122d91, 32'h4299fbb5, 32'h4185fd43, 32'h0};
test_input[16816:16823] = '{32'h423773f4, 32'hc1ab8240, 32'hc1964061, 32'h421982d6, 32'hc28c9373, 32'h421b6f1e, 32'hc1310b79, 32'hc2c3fa09};
test_output[16816:16823] = '{32'h423773f4, 32'h0, 32'h0, 32'h421982d6, 32'h0, 32'h421b6f1e, 32'h0, 32'h0};
test_input[16824:16831] = '{32'h428d7b3f, 32'hc2c140c3, 32'hc164e9ae, 32'hc1c00b64, 32'hc2286079, 32'h41c3d22a, 32'h42bfd473, 32'hc24652ec};
test_output[16824:16831] = '{32'h428d7b3f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41c3d22a, 32'h42bfd473, 32'h0};
test_input[16832:16839] = '{32'h428799d3, 32'hc0f62b64, 32'hc1178c97, 32'hc1d65689, 32'h41ee5aa2, 32'h4295a1af, 32'hc284ccca, 32'hc278f530};
test_output[16832:16839] = '{32'h428799d3, 32'h0, 32'h0, 32'h0, 32'h41ee5aa2, 32'h4295a1af, 32'h0, 32'h0};
test_input[16840:16847] = '{32'h42076919, 32'h423f182c, 32'h41806980, 32'hc2764142, 32'h428925fd, 32'hc29e4354, 32'h42ba9cd6, 32'h42846aa2};
test_output[16840:16847] = '{32'h42076919, 32'h423f182c, 32'h41806980, 32'h0, 32'h428925fd, 32'h0, 32'h42ba9cd6, 32'h42846aa2};
test_input[16848:16855] = '{32'hc271bec0, 32'hc265dabb, 32'hc1731a96, 32'hc20609f9, 32'h41443e8e, 32'h428530fd, 32'hc1f31f77, 32'h42875412};
test_output[16848:16855] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41443e8e, 32'h428530fd, 32'h0, 32'h42875412};
test_input[16856:16863] = '{32'h42ab2457, 32'h42b003b8, 32'h3e8e2ded, 32'h4272e58f, 32'h42921fd7, 32'hc1bec907, 32'hc2c214aa, 32'hc2835190};
test_output[16856:16863] = '{32'h42ab2457, 32'h42b003b8, 32'h3e8e2ded, 32'h4272e58f, 32'h42921fd7, 32'h0, 32'h0, 32'h0};
test_input[16864:16871] = '{32'h429bca45, 32'h42adfeed, 32'hc1679bc0, 32'h41cdfec1, 32'h3f8db3db, 32'hc1dff959, 32'hc28eff9f, 32'hc126c12e};
test_output[16864:16871] = '{32'h429bca45, 32'h42adfeed, 32'h0, 32'h41cdfec1, 32'h3f8db3db, 32'h0, 32'h0, 32'h0};
test_input[16872:16879] = '{32'hc1ad4e68, 32'h42b9d1f0, 32'hc2c261a1, 32'h4231f8cd, 32'hc24e9e41, 32'hc265fe39, 32'h42b8d38e, 32'h42396749};
test_output[16872:16879] = '{32'h0, 32'h42b9d1f0, 32'h0, 32'h4231f8cd, 32'h0, 32'h0, 32'h42b8d38e, 32'h42396749};
test_input[16880:16887] = '{32'h42074745, 32'h3f0a15c2, 32'hc28af20d, 32'h40a58b6d, 32'hc20b9036, 32'hc23a659e, 32'hc2b93bd2, 32'hc29c10b9};
test_output[16880:16887] = '{32'h42074745, 32'h3f0a15c2, 32'h0, 32'h40a58b6d, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16888:16895] = '{32'h41cc3f02, 32'h424e8ce7, 32'hc2c7d1d3, 32'h42bb94b8, 32'h42c44da9, 32'h42a35b68, 32'hc0f305f8, 32'hc1d62fcd};
test_output[16888:16895] = '{32'h41cc3f02, 32'h424e8ce7, 32'h0, 32'h42bb94b8, 32'h42c44da9, 32'h42a35b68, 32'h0, 32'h0};
test_input[16896:16903] = '{32'hc2aabfa0, 32'h4268b2b2, 32'h423b002e, 32'h42244378, 32'h42c3bcba, 32'hc28e2428, 32'hc237d17a, 32'h41f93f39};
test_output[16896:16903] = '{32'h0, 32'h4268b2b2, 32'h423b002e, 32'h42244378, 32'h42c3bcba, 32'h0, 32'h0, 32'h41f93f39};
test_input[16904:16911] = '{32'h41d3cf2f, 32'h4255061a, 32'hc2585b0a, 32'h3eadf2b6, 32'hc1306143, 32'hc06d9947, 32'hc142d6bc, 32'hbfe937a1};
test_output[16904:16911] = '{32'h41d3cf2f, 32'h4255061a, 32'h0, 32'h3eadf2b6, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16912:16919] = '{32'h4227639b, 32'h4204afc5, 32'hc1a02d3b, 32'hbf3338f8, 32'h42b572e9, 32'h3fabe79a, 32'h41d1f65e, 32'hc2ae1ea9};
test_output[16912:16919] = '{32'h4227639b, 32'h4204afc5, 32'h0, 32'h0, 32'h42b572e9, 32'h3fabe79a, 32'h41d1f65e, 32'h0};
test_input[16920:16927] = '{32'hc2287005, 32'h4290329e, 32'hc1ee20d8, 32'hc2936ac4, 32'h41801042, 32'hc01c2edd, 32'h426ad28a, 32'h4299f613};
test_output[16920:16927] = '{32'h0, 32'h4290329e, 32'h0, 32'h0, 32'h41801042, 32'h0, 32'h426ad28a, 32'h4299f613};
test_input[16928:16935] = '{32'hc295d6cb, 32'hc29684ec, 32'h3dead61f, 32'h428ba455, 32'h4287db97, 32'h4196a962, 32'hc297c2f6, 32'h425f7042};
test_output[16928:16935] = '{32'h0, 32'h0, 32'h3dead61f, 32'h428ba455, 32'h4287db97, 32'h4196a962, 32'h0, 32'h425f7042};
test_input[16936:16943] = '{32'hc2b7d6ce, 32'h42a8140e, 32'hc1b9c02b, 32'h40fcc7e7, 32'hc14d9fd2, 32'hc2a36f62, 32'hc2446c60, 32'h429741e7};
test_output[16936:16943] = '{32'h0, 32'h42a8140e, 32'h0, 32'h40fcc7e7, 32'h0, 32'h0, 32'h0, 32'h429741e7};
test_input[16944:16951] = '{32'h3f03389f, 32'h420d6cc4, 32'hc20010cc, 32'h41a9f829, 32'h42aa16a4, 32'h4241b11d, 32'h4297be6d, 32'h41efafde};
test_output[16944:16951] = '{32'h3f03389f, 32'h420d6cc4, 32'h0, 32'h41a9f829, 32'h42aa16a4, 32'h4241b11d, 32'h4297be6d, 32'h41efafde};
test_input[16952:16959] = '{32'hc217036d, 32'hc187f9cf, 32'h42646b67, 32'hc1e29329, 32'hc263777d, 32'h411c2b65, 32'h4287b2cc, 32'hc241a43c};
test_output[16952:16959] = '{32'h0, 32'h0, 32'h42646b67, 32'h0, 32'h0, 32'h411c2b65, 32'h4287b2cc, 32'h0};
test_input[16960:16967] = '{32'h42734fbc, 32'h422b2fb0, 32'h41e0e0e6, 32'hc2be38fa, 32'hc2343df1, 32'h41fc6075, 32'hc2b7df47, 32'h420bf206};
test_output[16960:16967] = '{32'h42734fbc, 32'h422b2fb0, 32'h41e0e0e6, 32'h0, 32'h0, 32'h41fc6075, 32'h0, 32'h420bf206};
test_input[16968:16975] = '{32'hc1522bbb, 32'hc2a5ad64, 32'h42a8e9ca, 32'hc1f7d618, 32'h42a1cdff, 32'hc2909eb4, 32'hc1bba327, 32'hc2352cc2};
test_output[16968:16975] = '{32'h0, 32'h0, 32'h42a8e9ca, 32'h0, 32'h42a1cdff, 32'h0, 32'h0, 32'h0};
test_input[16976:16983] = '{32'h3fbfd35c, 32'hc2c32a32, 32'h428c42b1, 32'h42bca1c1, 32'hc2a787b9, 32'hc1bf71c6, 32'h426e4831, 32'h40d03bef};
test_output[16976:16983] = '{32'h3fbfd35c, 32'h0, 32'h428c42b1, 32'h42bca1c1, 32'h0, 32'h0, 32'h426e4831, 32'h40d03bef};
test_input[16984:16991] = '{32'hc2b05eec, 32'hc2a33c01, 32'h42795eca, 32'h42acad20, 32'h423c1cdc, 32'h40f96b3d, 32'hc1b41c9c, 32'h423d6481};
test_output[16984:16991] = '{32'h0, 32'h0, 32'h42795eca, 32'h42acad20, 32'h423c1cdc, 32'h40f96b3d, 32'h0, 32'h423d6481};
test_input[16992:16999] = '{32'h422be92a, 32'hc2324466, 32'h42095c91, 32'h422fbf94, 32'hc1fc996f, 32'hc2882f16, 32'hc063f66b, 32'h4106aa9e};
test_output[16992:16999] = '{32'h422be92a, 32'h0, 32'h42095c91, 32'h422fbf94, 32'h0, 32'h0, 32'h0, 32'h4106aa9e};
test_input[17000:17007] = '{32'h42a2e1ec, 32'h42bd6af1, 32'h3f31ca6f, 32'h40e52034, 32'hc10e6124, 32'hc2c0a169, 32'h41500ec7, 32'h41f6ad31};
test_output[17000:17007] = '{32'h42a2e1ec, 32'h42bd6af1, 32'h3f31ca6f, 32'h40e52034, 32'h0, 32'h0, 32'h41500ec7, 32'h41f6ad31};
test_input[17008:17015] = '{32'h42121cd9, 32'h4288d314, 32'hc2c50fbb, 32'h410162b2, 32'hc222063c, 32'h428c640f, 32'hc22b94e3, 32'hc2692717};
test_output[17008:17015] = '{32'h42121cd9, 32'h4288d314, 32'h0, 32'h410162b2, 32'h0, 32'h428c640f, 32'h0, 32'h0};
test_input[17016:17023] = '{32'hc2407751, 32'hc28076e2, 32'h41ed483e, 32'h422bfcff, 32'h40ef98b8, 32'hc29f38cc, 32'h42464524, 32'hc28bebd0};
test_output[17016:17023] = '{32'h0, 32'h0, 32'h41ed483e, 32'h422bfcff, 32'h40ef98b8, 32'h0, 32'h42464524, 32'h0};
test_input[17024:17031] = '{32'hc236f515, 32'h426d9375, 32'h4193d12e, 32'hc1b13e91, 32'h42988ccb, 32'h42b7a88a, 32'hc2406385, 32'h41a08d69};
test_output[17024:17031] = '{32'h0, 32'h426d9375, 32'h4193d12e, 32'h0, 32'h42988ccb, 32'h42b7a88a, 32'h0, 32'h41a08d69};
test_input[17032:17039] = '{32'h3fc5988f, 32'hc1852657, 32'h41a59b7a, 32'h421628e1, 32'hc2736aeb, 32'hc29fa639, 32'hc2704efc, 32'hc2159475};
test_output[17032:17039] = '{32'h3fc5988f, 32'h0, 32'h41a59b7a, 32'h421628e1, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[17040:17047] = '{32'hc210c2a3, 32'hc2971ce6, 32'hc0003f0d, 32'hc214db75, 32'h42190348, 32'h4261f448, 32'hc05e708a, 32'hc107d14f};
test_output[17040:17047] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42190348, 32'h4261f448, 32'h0, 32'h0};
test_input[17048:17055] = '{32'hc25cb6c1, 32'h4257435e, 32'h4271c43d, 32'hc25e2513, 32'hc2c6c814, 32'h427d20e1, 32'h42605ee8, 32'h4216bbb8};
test_output[17048:17055] = '{32'h0, 32'h4257435e, 32'h4271c43d, 32'h0, 32'h0, 32'h427d20e1, 32'h42605ee8, 32'h4216bbb8};
test_input[17056:17063] = '{32'h41a9ce1c, 32'hc1cd00f2, 32'h42612acc, 32'h422f25fa, 32'h41ab7517, 32'h418207be, 32'h421ebccb, 32'h4280abd7};
test_output[17056:17063] = '{32'h41a9ce1c, 32'h0, 32'h42612acc, 32'h422f25fa, 32'h41ab7517, 32'h418207be, 32'h421ebccb, 32'h4280abd7};
test_input[17064:17071] = '{32'h42ac7a57, 32'hc21d34d3, 32'hc03dd3bb, 32'hc20a15ff, 32'hc2ac2856, 32'h418b1c72, 32'h4247ed1b, 32'h42a207c3};
test_output[17064:17071] = '{32'h42ac7a57, 32'h0, 32'h0, 32'h0, 32'h0, 32'h418b1c72, 32'h4247ed1b, 32'h42a207c3};
test_input[17072:17079] = '{32'hc258ec3d, 32'hc2b5d200, 32'hc205a5ed, 32'h4287a7e0, 32'h42a8827b, 32'hc2be1459, 32'h41b00da3, 32'h3f67dafb};
test_output[17072:17079] = '{32'h0, 32'h0, 32'h0, 32'h4287a7e0, 32'h42a8827b, 32'h0, 32'h41b00da3, 32'h3f67dafb};
test_input[17080:17087] = '{32'hc2a4dee3, 32'hc1c99d9a, 32'h4283d02f, 32'h4246ef62, 32'hc295b594, 32'hc0d189b3, 32'h4213251a, 32'h425f7c0a};
test_output[17080:17087] = '{32'h0, 32'h0, 32'h4283d02f, 32'h4246ef62, 32'h0, 32'h0, 32'h4213251a, 32'h425f7c0a};
test_input[17088:17095] = '{32'h4297e7e9, 32'h40cf6c54, 32'h428bc91a, 32'h42c547e4, 32'h4252b054, 32'h406a72b5, 32'h426ad6e9, 32'hc2b769a0};
test_output[17088:17095] = '{32'h4297e7e9, 32'h40cf6c54, 32'h428bc91a, 32'h42c547e4, 32'h4252b054, 32'h406a72b5, 32'h426ad6e9, 32'h0};
test_input[17096:17103] = '{32'h42a6f738, 32'hc2bdcedc, 32'hc2209f59, 32'hc1eb3c5c, 32'hc26aaa92, 32'h42a1cb70, 32'h41f73e14, 32'hc295f97d};
test_output[17096:17103] = '{32'h42a6f738, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a1cb70, 32'h41f73e14, 32'h0};
test_input[17104:17111] = '{32'hc28da9bc, 32'h42ba79b0, 32'hc2ba8a6d, 32'h42748eb1, 32'h41c4add2, 32'h42793d7c, 32'h42c6aee6, 32'h428bbdf8};
test_output[17104:17111] = '{32'h0, 32'h42ba79b0, 32'h0, 32'h42748eb1, 32'h41c4add2, 32'h42793d7c, 32'h42c6aee6, 32'h428bbdf8};
test_input[17112:17119] = '{32'hc2037620, 32'h40d6c29d, 32'h422192aa, 32'h428d3d83, 32'hc02e880c, 32'hc2637ed2, 32'h4275478c, 32'hc249e7c6};
test_output[17112:17119] = '{32'h0, 32'h40d6c29d, 32'h422192aa, 32'h428d3d83, 32'h0, 32'h0, 32'h4275478c, 32'h0};
test_input[17120:17127] = '{32'hbfdb828d, 32'hc18569ae, 32'h4297ef40, 32'hc25c0a8b, 32'hc191c850, 32'h41c214e3, 32'hc1bfcdfb, 32'h42ac95c8};
test_output[17120:17127] = '{32'h0, 32'h0, 32'h4297ef40, 32'h0, 32'h0, 32'h41c214e3, 32'h0, 32'h42ac95c8};
test_input[17128:17135] = '{32'hc167fffd, 32'hc296ff72, 32'hc1c4e577, 32'h425ea971, 32'h415c8326, 32'h42908992, 32'hc2602816, 32'h4286704d};
test_output[17128:17135] = '{32'h0, 32'h0, 32'h0, 32'h425ea971, 32'h415c8326, 32'h42908992, 32'h0, 32'h4286704d};
test_input[17136:17143] = '{32'hc1be2e6c, 32'h429a1bb9, 32'hc1ad321b, 32'hc2a78582, 32'h428f46d9, 32'h42c74833, 32'hc2bdc3aa, 32'h41c53ac9};
test_output[17136:17143] = '{32'h0, 32'h429a1bb9, 32'h0, 32'h0, 32'h428f46d9, 32'h42c74833, 32'h0, 32'h41c53ac9};
test_input[17144:17151] = '{32'h42b2924e, 32'hc2be11fe, 32'h41adf880, 32'h42c71ca3, 32'hc2841559, 32'hbeab414e, 32'hc286c0a7, 32'h3e7742dc};
test_output[17144:17151] = '{32'h42b2924e, 32'h0, 32'h41adf880, 32'h42c71ca3, 32'h0, 32'h0, 32'h0, 32'h3e7742dc};
test_input[17152:17159] = '{32'h4014e79c, 32'h4267a69b, 32'hc26a316d, 32'h41cba6fa, 32'hc0854787, 32'hc2c08003, 32'hc2415e11, 32'hc2984b3e};
test_output[17152:17159] = '{32'h4014e79c, 32'h4267a69b, 32'h0, 32'h41cba6fa, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[17160:17167] = '{32'hc16fad04, 32'h41d0b5f1, 32'h41e4a113, 32'h422d5cb9, 32'hc2ba5e6d, 32'h429f17d0, 32'hc299e330, 32'h4264cfd6};
test_output[17160:17167] = '{32'h0, 32'h41d0b5f1, 32'h41e4a113, 32'h422d5cb9, 32'h0, 32'h429f17d0, 32'h0, 32'h4264cfd6};
test_input[17168:17175] = '{32'hc2bb8d5f, 32'hc167ffec, 32'hc17b1de2, 32'hc17a09b1, 32'h429dd0be, 32'h42918e86, 32'hc26e484e, 32'h41eae710};
test_output[17168:17175] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429dd0be, 32'h42918e86, 32'h0, 32'h41eae710};
test_input[17176:17183] = '{32'h4297a3df, 32'h42b2299b, 32'hc2b4546b, 32'hc2388fff, 32'hc29bad00, 32'h428a858a, 32'hc1d07e95, 32'h429b691b};
test_output[17176:17183] = '{32'h4297a3df, 32'h42b2299b, 32'h0, 32'h0, 32'h0, 32'h428a858a, 32'h0, 32'h429b691b};
test_input[17184:17191] = '{32'h42c60264, 32'h3fa25f58, 32'h42413c81, 32'hc29626c1, 32'hc2266021, 32'h42060cd5, 32'h4291953d, 32'h4287efd9};
test_output[17184:17191] = '{32'h42c60264, 32'h3fa25f58, 32'h42413c81, 32'h0, 32'h0, 32'h42060cd5, 32'h4291953d, 32'h4287efd9};
test_input[17192:17199] = '{32'hc24f5193, 32'hc1d3b56d, 32'h422b32ac, 32'hc2469639, 32'h421f2ea1, 32'hbfec6720, 32'h42a63ee0, 32'h427279cf};
test_output[17192:17199] = '{32'h0, 32'h0, 32'h422b32ac, 32'h0, 32'h421f2ea1, 32'h0, 32'h42a63ee0, 32'h427279cf};
test_input[17200:17207] = '{32'hc2970466, 32'hc22dde9e, 32'hc172f8c8, 32'h41fa7ef0, 32'hc2c13699, 32'h428a24c0, 32'hc2680a1c, 32'h429e32ca};
test_output[17200:17207] = '{32'h0, 32'h0, 32'h0, 32'h41fa7ef0, 32'h0, 32'h428a24c0, 32'h0, 32'h429e32ca};
test_input[17208:17215] = '{32'h429e42dd, 32'h426c491e, 32'h423f347f, 32'h41d7da83, 32'h4298420e, 32'h425decd5, 32'hc2b97ae7, 32'hc28ae75f};
test_output[17208:17215] = '{32'h429e42dd, 32'h426c491e, 32'h423f347f, 32'h41d7da83, 32'h4298420e, 32'h425decd5, 32'h0, 32'h0};
test_input[17216:17223] = '{32'hc2aec95e, 32'hc2893b3c, 32'h42b52a2a, 32'h42c5ca6f, 32'h4217f741, 32'hc217ac37, 32'hc1dc9e1e, 32'hc26bbfc1};
test_output[17216:17223] = '{32'h0, 32'h0, 32'h42b52a2a, 32'h42c5ca6f, 32'h4217f741, 32'h0, 32'h0, 32'h0};
test_input[17224:17231] = '{32'h4256c212, 32'h4242efdb, 32'h42820153, 32'hc2abfcf4, 32'h427d21e4, 32'h424589e9, 32'hc2b4b0ee, 32'h4218fd34};
test_output[17224:17231] = '{32'h4256c212, 32'h4242efdb, 32'h42820153, 32'h0, 32'h427d21e4, 32'h424589e9, 32'h0, 32'h4218fd34};
test_input[17232:17239] = '{32'hc1c3f10e, 32'h413358ee, 32'hc2c4d301, 32'hc23f4374, 32'hc19498c5, 32'h41b9eee8, 32'h42aa12fd, 32'hc1d29d88};
test_output[17232:17239] = '{32'h0, 32'h413358ee, 32'h0, 32'h0, 32'h0, 32'h41b9eee8, 32'h42aa12fd, 32'h0};
test_input[17240:17247] = '{32'h4151a15a, 32'hc2c1162e, 32'h428235d9, 32'hc07a45c2, 32'h42a3a078, 32'h41ee1286, 32'hc2268771, 32'h424cd4f7};
test_output[17240:17247] = '{32'h4151a15a, 32'h0, 32'h428235d9, 32'h0, 32'h42a3a078, 32'h41ee1286, 32'h0, 32'h424cd4f7};
test_input[17248:17255] = '{32'hc29d0106, 32'hc2abca67, 32'h41f91508, 32'h42996dba, 32'h41c7cbd2, 32'hc1fd62e1, 32'h3f308b5f, 32'h427d5da6};
test_output[17248:17255] = '{32'h0, 32'h0, 32'h41f91508, 32'h42996dba, 32'h41c7cbd2, 32'h0, 32'h3f308b5f, 32'h427d5da6};
test_input[17256:17263] = '{32'h42bb7641, 32'h417e541b, 32'h428b3fe0, 32'h408ee51e, 32'hc279787e, 32'hc2914c86, 32'h42173bcf, 32'hc2943b6d};
test_output[17256:17263] = '{32'h42bb7641, 32'h417e541b, 32'h428b3fe0, 32'h408ee51e, 32'h0, 32'h0, 32'h42173bcf, 32'h0};
test_input[17264:17271] = '{32'h42af7d19, 32'h4292ff37, 32'h4199a7cf, 32'hc28a91e7, 32'h41cd4399, 32'h426f208c, 32'h41930425, 32'hc1b44d0d};
test_output[17264:17271] = '{32'h42af7d19, 32'h4292ff37, 32'h4199a7cf, 32'h0, 32'h41cd4399, 32'h426f208c, 32'h41930425, 32'h0};
test_input[17272:17279] = '{32'h42770615, 32'h4233f665, 32'hc22b3691, 32'hc114b442, 32'h4218829d, 32'hc27e21c9, 32'hc1035df6, 32'h40768a5e};
test_output[17272:17279] = '{32'h42770615, 32'h4233f665, 32'h0, 32'h0, 32'h4218829d, 32'h0, 32'h0, 32'h40768a5e};
test_input[17280:17287] = '{32'h422c89b8, 32'hc1e101ec, 32'h42bc7a73, 32'h40d30603, 32'hc1103851, 32'h428017bb, 32'hc24b6e47, 32'h3fb3cacf};
test_output[17280:17287] = '{32'h422c89b8, 32'h0, 32'h42bc7a73, 32'h40d30603, 32'h0, 32'h428017bb, 32'h0, 32'h3fb3cacf};
test_input[17288:17295] = '{32'hc1cd552f, 32'hc202a550, 32'h4245ff4b, 32'hc2948a8c, 32'h425dc89d, 32'hc2739b53, 32'hc2686418, 32'hc23a7243};
test_output[17288:17295] = '{32'h0, 32'h0, 32'h4245ff4b, 32'h0, 32'h425dc89d, 32'h0, 32'h0, 32'h0};
test_input[17296:17303] = '{32'hc193e176, 32'h4255a332, 32'h41de35b3, 32'hc2953eca, 32'h4265f74f, 32'hc12781f8, 32'h42489a57, 32'hc249548b};
test_output[17296:17303] = '{32'h0, 32'h4255a332, 32'h41de35b3, 32'h0, 32'h4265f74f, 32'h0, 32'h42489a57, 32'h0};
test_input[17304:17311] = '{32'h42bca2dd, 32'hc1e047c7, 32'h423afa6a, 32'h423c0c5f, 32'h4277e401, 32'hc128b883, 32'hc1b98ad2, 32'h42bfe5dc};
test_output[17304:17311] = '{32'h42bca2dd, 32'h0, 32'h423afa6a, 32'h423c0c5f, 32'h4277e401, 32'h0, 32'h0, 32'h42bfe5dc};
test_input[17312:17319] = '{32'h42a580e1, 32'hc2c7e131, 32'hc1df393e, 32'h41a8c290, 32'h42a73d0a, 32'hc20da6e2, 32'h4283d945, 32'h421b2af8};
test_output[17312:17319] = '{32'h42a580e1, 32'h0, 32'h0, 32'h41a8c290, 32'h42a73d0a, 32'h0, 32'h4283d945, 32'h421b2af8};
test_input[17320:17327] = '{32'hc1442d7a, 32'h427ddcb2, 32'h41b4800f, 32'hc2bc802a, 32'h4264f14d, 32'hc275dd5c, 32'h412f1a1f, 32'hc2b99db1};
test_output[17320:17327] = '{32'h0, 32'h427ddcb2, 32'h41b4800f, 32'h0, 32'h4264f14d, 32'h0, 32'h412f1a1f, 32'h0};
test_input[17328:17335] = '{32'h414049af, 32'h42967daa, 32'hc2b7ee1a, 32'hc2269fa0, 32'hc23fbbad, 32'hc29767f9, 32'hc29ddcb6, 32'h426060ff};
test_output[17328:17335] = '{32'h414049af, 32'h42967daa, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426060ff};
test_input[17336:17343] = '{32'hc294fa19, 32'h421250ca, 32'hc2ae0a5b, 32'hc25cf620, 32'hbf749a1d, 32'hc26e0947, 32'h41bad093, 32'hc219d35d};
test_output[17336:17343] = '{32'h0, 32'h421250ca, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41bad093, 32'h0};
test_input[17344:17351] = '{32'hc087622c, 32'hc081f416, 32'hc2c74ba0, 32'hc28c088f, 32'h428df6ed, 32'h421f76f2, 32'h40e8244a, 32'h428d607f};
test_output[17344:17351] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h428df6ed, 32'h421f76f2, 32'h40e8244a, 32'h428d607f};
test_input[17352:17359] = '{32'hc2897612, 32'h41f163b4, 32'hc2babd75, 32'hc227cadf, 32'h421c4aed, 32'h427c773f, 32'hc2b527b2, 32'hc27f366f};
test_output[17352:17359] = '{32'h0, 32'h41f163b4, 32'h0, 32'h0, 32'h421c4aed, 32'h427c773f, 32'h0, 32'h0};
test_input[17360:17367] = '{32'h4230e98b, 32'h42785d28, 32'hc2bd26bd, 32'h42136433, 32'hc2878c69, 32'hbf85bcc6, 32'h428aca1c, 32'hc2965c78};
test_output[17360:17367] = '{32'h4230e98b, 32'h42785d28, 32'h0, 32'h42136433, 32'h0, 32'h0, 32'h428aca1c, 32'h0};
test_input[17368:17375] = '{32'hc282cf1d, 32'hc1cdb988, 32'hc2926e7e, 32'h426ae8c2, 32'h42946e00, 32'hc226398f, 32'hc225b24b, 32'h408a7c72};
test_output[17368:17375] = '{32'h0, 32'h0, 32'h0, 32'h426ae8c2, 32'h42946e00, 32'h0, 32'h0, 32'h408a7c72};
test_input[17376:17383] = '{32'hc26bf744, 32'hc27293b7, 32'hc29d86f6, 32'hc0a78cf3, 32'hc28673ba, 32'hbf015cda, 32'hc1672594, 32'h42a6b6e7};
test_output[17376:17383] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a6b6e7};
test_input[17384:17391] = '{32'hc2802097, 32'hc1db7296, 32'hc295da24, 32'h418b1151, 32'h42bf54ae, 32'h42210d11, 32'hbf9b982e, 32'h4294f36c};
test_output[17384:17391] = '{32'h0, 32'h0, 32'h0, 32'h418b1151, 32'h42bf54ae, 32'h42210d11, 32'h0, 32'h4294f36c};
test_input[17392:17399] = '{32'hc185699d, 32'hc2a13280, 32'hc1099c1f, 32'h425ed844, 32'h42860558, 32'h429b6794, 32'hc2ba536a, 32'hc2965747};
test_output[17392:17399] = '{32'h0, 32'h0, 32'h0, 32'h425ed844, 32'h42860558, 32'h429b6794, 32'h0, 32'h0};
test_input[17400:17407] = '{32'h42b47698, 32'h42c66d25, 32'hc1940424, 32'h42b1cc0e, 32'hc21a544f, 32'h42399d6d, 32'hc2429712, 32'h41815202};
test_output[17400:17407] = '{32'h42b47698, 32'h42c66d25, 32'h0, 32'h42b1cc0e, 32'h0, 32'h42399d6d, 32'h0, 32'h41815202};
test_input[17408:17415] = '{32'hc2672bb6, 32'hc29c6c7f, 32'hc28d2e17, 32'h41440684, 32'hc21fef62, 32'h42473a54, 32'h422dabea, 32'hc24281f0};
test_output[17408:17415] = '{32'h0, 32'h0, 32'h0, 32'h41440684, 32'h0, 32'h42473a54, 32'h422dabea, 32'h0};
test_input[17416:17423] = '{32'hc2c79cc0, 32'h422b9a52, 32'h42612530, 32'h41304c1a, 32'h42af33e5, 32'h41ebdbaf, 32'h408c09fa, 32'h428d2cbf};
test_output[17416:17423] = '{32'h0, 32'h422b9a52, 32'h42612530, 32'h41304c1a, 32'h42af33e5, 32'h41ebdbaf, 32'h408c09fa, 32'h428d2cbf};
test_input[17424:17431] = '{32'hc18a8509, 32'hc0eec3be, 32'hc2b134fc, 32'h42a8a27e, 32'hc2c7f6fd, 32'h42bbf642, 32'hc1d6f651, 32'hc174871e};
test_output[17424:17431] = '{32'h0, 32'h0, 32'h0, 32'h42a8a27e, 32'h0, 32'h42bbf642, 32'h0, 32'h0};
test_input[17432:17439] = '{32'h423faa4d, 32'h42224a73, 32'h41aecc9a, 32'h418aed55, 32'hc1ff9e96, 32'hc2bfdecb, 32'h4257fed3, 32'h4257677a};
test_output[17432:17439] = '{32'h423faa4d, 32'h42224a73, 32'h41aecc9a, 32'h418aed55, 32'h0, 32'h0, 32'h4257fed3, 32'h4257677a};
test_input[17440:17447] = '{32'h420e387c, 32'h42ac6270, 32'h421a77d4, 32'hc2436aa2, 32'hc22d909e, 32'h41d19a18, 32'hc19dcd74, 32'hc20976ec};
test_output[17440:17447] = '{32'h420e387c, 32'h42ac6270, 32'h421a77d4, 32'h0, 32'h0, 32'h41d19a18, 32'h0, 32'h0};
test_input[17448:17455] = '{32'hc2913a91, 32'hc2846315, 32'hc1796f19, 32'hc2244924, 32'h42a17285, 32'h410a997c, 32'hc2281f47, 32'h40a2a262};
test_output[17448:17455] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a17285, 32'h410a997c, 32'h0, 32'h40a2a262};
test_input[17456:17463] = '{32'h42751415, 32'hc2905891, 32'h423cb926, 32'hc2852ecd, 32'hc1ccc400, 32'h425073ec, 32'hc2afe9a6, 32'h41d6aa95};
test_output[17456:17463] = '{32'h42751415, 32'h0, 32'h423cb926, 32'h0, 32'h0, 32'h425073ec, 32'h0, 32'h41d6aa95};
test_input[17464:17471] = '{32'h414c65f9, 32'hc2b574be, 32'hc2567c6a, 32'h42aa4041, 32'hc1eda5ee, 32'hc1a3cb63, 32'h422adf66, 32'h420d2e35};
test_output[17464:17471] = '{32'h414c65f9, 32'h0, 32'h0, 32'h42aa4041, 32'h0, 32'h0, 32'h422adf66, 32'h420d2e35};
test_input[17472:17479] = '{32'hc1e470b8, 32'hc21ef05e, 32'hc01f2a64, 32'h4213c785, 32'hc0166fc3, 32'hc28f9c12, 32'hc198898b, 32'h42aa22c6};
test_output[17472:17479] = '{32'h0, 32'h0, 32'h0, 32'h4213c785, 32'h0, 32'h0, 32'h0, 32'h42aa22c6};
test_input[17480:17487] = '{32'hc1d416fa, 32'hc0e5d16b, 32'hc2a7984b, 32'h42429a13, 32'h42c6999f, 32'hc2c4d9cf, 32'h4272907b, 32'h422b0b0c};
test_output[17480:17487] = '{32'h0, 32'h0, 32'h0, 32'h42429a13, 32'h42c6999f, 32'h0, 32'h4272907b, 32'h422b0b0c};
test_input[17488:17495] = '{32'hc1f378e2, 32'hc2a8fdeb, 32'h42a92b49, 32'hc261217f, 32'h4199036c, 32'h4257fefc, 32'h42adf5e4, 32'h3d2f7035};
test_output[17488:17495] = '{32'h0, 32'h0, 32'h42a92b49, 32'h0, 32'h4199036c, 32'h4257fefc, 32'h42adf5e4, 32'h3d2f7035};
test_input[17496:17503] = '{32'h4201f54c, 32'hc2802fd5, 32'hc1e2763c, 32'h42a7f742, 32'hc224d334, 32'h4284ec77, 32'h41f4ab72, 32'h42902eee};
test_output[17496:17503] = '{32'h4201f54c, 32'h0, 32'h0, 32'h42a7f742, 32'h0, 32'h4284ec77, 32'h41f4ab72, 32'h42902eee};
test_input[17504:17511] = '{32'h4218b6df, 32'hc2b94033, 32'hc297c65a, 32'hc258b82a, 32'hc292a51c, 32'h428af138, 32'h42567467, 32'hc1c851c1};
test_output[17504:17511] = '{32'h4218b6df, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428af138, 32'h42567467, 32'h0};
test_input[17512:17519] = '{32'hc1f06852, 32'hc204265c, 32'hc20d6b5a, 32'h4187629a, 32'hc2812b4b, 32'hc2965173, 32'hc14308c1, 32'hc2305c56};
test_output[17512:17519] = '{32'h0, 32'h0, 32'h0, 32'h4187629a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[17520:17527] = '{32'hc147fc54, 32'hc2961f1e, 32'h4228685f, 32'hc1d912fe, 32'h4293cbb2, 32'hc1ba9c83, 32'hc207cdfb, 32'hc26c8433};
test_output[17520:17527] = '{32'h0, 32'h0, 32'h4228685f, 32'h0, 32'h4293cbb2, 32'h0, 32'h0, 32'h0};
test_input[17528:17535] = '{32'h42485775, 32'h428b6f44, 32'hc10dc248, 32'h423e68a0, 32'hbe25eea0, 32'hc25e9fd3, 32'h4242bf99, 32'hc2b9b0d8};
test_output[17528:17535] = '{32'h42485775, 32'h428b6f44, 32'h0, 32'h423e68a0, 32'h0, 32'h0, 32'h4242bf99, 32'h0};
test_input[17536:17543] = '{32'h40e7d15f, 32'hc17f1adb, 32'h42b5a19d, 32'hbfb539ef, 32'h423de485, 32'h418d8cc1, 32'hc1809ae8, 32'hc1f09462};
test_output[17536:17543] = '{32'h40e7d15f, 32'h0, 32'h42b5a19d, 32'h0, 32'h423de485, 32'h418d8cc1, 32'h0, 32'h0};
test_input[17544:17551] = '{32'hc22b7cd3, 32'hc1a0d733, 32'hc1e25244, 32'hc2c797a1, 32'h41a71869, 32'h4295b4d6, 32'h42471e01, 32'h42a4d210};
test_output[17544:17551] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41a71869, 32'h4295b4d6, 32'h42471e01, 32'h42a4d210};
test_input[17552:17559] = '{32'h420df3f5, 32'hc263211e, 32'hc2c128aa, 32'hc2ada99f, 32'hc1f15f9e, 32'hc2a0537b, 32'h41aa5ea4, 32'hc0ef1982};
test_output[17552:17559] = '{32'h420df3f5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41aa5ea4, 32'h0};
test_input[17560:17567] = '{32'hc2768338, 32'h42922c00, 32'hc17472b6, 32'hc25b6782, 32'hc2634873, 32'h42a8cace, 32'h41def0f3, 32'h42b30675};
test_output[17560:17567] = '{32'h0, 32'h42922c00, 32'h0, 32'h0, 32'h0, 32'h42a8cace, 32'h41def0f3, 32'h42b30675};
test_input[17568:17575] = '{32'h41840841, 32'hc0269f16, 32'hc2b367df, 32'h42a6e389, 32'h429eb077, 32'hc285439e, 32'h42887391, 32'h422ba278};
test_output[17568:17575] = '{32'h41840841, 32'h0, 32'h0, 32'h42a6e389, 32'h429eb077, 32'h0, 32'h42887391, 32'h422ba278};
test_input[17576:17583] = '{32'hc29aa9d3, 32'hc20fca03, 32'h429f0473, 32'hc2ad075a, 32'hc1ae7231, 32'hc26cfde6, 32'h4152e2a6, 32'h3f013d45};
test_output[17576:17583] = '{32'h0, 32'h0, 32'h429f0473, 32'h0, 32'h0, 32'h0, 32'h4152e2a6, 32'h3f013d45};
test_input[17584:17591] = '{32'hc297b52d, 32'h42202dfd, 32'h4282b234, 32'hc1380bec, 32'h416f0ba9, 32'hc2a113fb, 32'h427cea59, 32'hc01452e8};
test_output[17584:17591] = '{32'h0, 32'h42202dfd, 32'h4282b234, 32'h0, 32'h416f0ba9, 32'h0, 32'h427cea59, 32'h0};
test_input[17592:17599] = '{32'hc22d4092, 32'hc209934e, 32'hc213ae5f, 32'h42a13aac, 32'hc2278d95, 32'h42988183, 32'hc2a26c96, 32'h42b0a502};
test_output[17592:17599] = '{32'h0, 32'h0, 32'h0, 32'h42a13aac, 32'h0, 32'h42988183, 32'h0, 32'h42b0a502};
test_input[17600:17607] = '{32'h42a0498b, 32'h4255597d, 32'h42922fdc, 32'h3ff688c9, 32'h41a1278d, 32'hc2624a9d, 32'hc242b751, 32'hc0a9069f};
test_output[17600:17607] = '{32'h42a0498b, 32'h4255597d, 32'h42922fdc, 32'h3ff688c9, 32'h41a1278d, 32'h0, 32'h0, 32'h0};
test_input[17608:17615] = '{32'hc202b325, 32'h42bd48fd, 32'hc23817e6, 32'hc2b36f6d, 32'h42894841, 32'hc2ae69dd, 32'hc2736d03, 32'h42ba1343};
test_output[17608:17615] = '{32'h0, 32'h42bd48fd, 32'h0, 32'h0, 32'h42894841, 32'h0, 32'h0, 32'h42ba1343};
test_input[17616:17623] = '{32'hc08a259c, 32'h425fc381, 32'hc202165f, 32'h42409fad, 32'hc2c74eee, 32'hc2ac098c, 32'hc297733e, 32'h41903b82};
test_output[17616:17623] = '{32'h0, 32'h425fc381, 32'h0, 32'h42409fad, 32'h0, 32'h0, 32'h0, 32'h41903b82};
test_input[17624:17631] = '{32'hc2c34cd7, 32'h3f0e9aab, 32'hc28d1ac5, 32'h421a5c9d, 32'hc0f9b271, 32'h41cf4c9a, 32'hc2b9bb98, 32'hc2c1a4c4};
test_output[17624:17631] = '{32'h0, 32'h3f0e9aab, 32'h0, 32'h421a5c9d, 32'h0, 32'h41cf4c9a, 32'h0, 32'h0};
test_input[17632:17639] = '{32'hc287bce4, 32'h408b3bce, 32'hc2baaebe, 32'hc21a55fb, 32'h42af4e36, 32'hc28d9534, 32'hc2334ad2, 32'h4298c93d};
test_output[17632:17639] = '{32'h0, 32'h408b3bce, 32'h0, 32'h0, 32'h42af4e36, 32'h0, 32'h0, 32'h4298c93d};
test_input[17640:17647] = '{32'hc27c1d23, 32'hc210c6fa, 32'hc2bf0a4c, 32'h42a767db, 32'h42b5bc17, 32'hc2a00390, 32'h427f63ce, 32'h407b428e};
test_output[17640:17647] = '{32'h0, 32'h0, 32'h0, 32'h42a767db, 32'h42b5bc17, 32'h0, 32'h427f63ce, 32'h407b428e};
test_input[17648:17655] = '{32'h42bfa14a, 32'hc15238e1, 32'hc23c6c2d, 32'hc0f5283f, 32'hc2992aa4, 32'h422c0909, 32'hc25d63d7, 32'h4217b3f9};
test_output[17648:17655] = '{32'h42bfa14a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422c0909, 32'h0, 32'h4217b3f9};
test_input[17656:17663] = '{32'hc24acc5a, 32'hc27a7887, 32'hc1fe0a43, 32'h419d0b1d, 32'h42c4c9e3, 32'h42956d57, 32'h428f3a3a, 32'hc20be79c};
test_output[17656:17663] = '{32'h0, 32'h0, 32'h0, 32'h419d0b1d, 32'h42c4c9e3, 32'h42956d57, 32'h428f3a3a, 32'h0};
test_input[17664:17671] = '{32'hc2c322a2, 32'hc2aaa229, 32'hc2c639d2, 32'hc249398b, 32'hc24c516a, 32'h4152ced9, 32'hc236021d, 32'h4242b5ba};
test_output[17664:17671] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4152ced9, 32'h0, 32'h4242b5ba};
test_input[17672:17679] = '{32'h422d91ec, 32'h41d0d7e3, 32'hc0984521, 32'hc24d8f1c, 32'h4006e9c2, 32'h412ae918, 32'h425441c7, 32'hc21227b4};
test_output[17672:17679] = '{32'h422d91ec, 32'h41d0d7e3, 32'h0, 32'h0, 32'h4006e9c2, 32'h412ae918, 32'h425441c7, 32'h0};
test_input[17680:17687] = '{32'hc198e64f, 32'h42aeb6d1, 32'h429b7269, 32'h42896cba, 32'hc12a9fd8, 32'hc2a97cc0, 32'hc2a966a6, 32'h42b6056a};
test_output[17680:17687] = '{32'h0, 32'h42aeb6d1, 32'h429b7269, 32'h42896cba, 32'h0, 32'h0, 32'h0, 32'h42b6056a};
test_input[17688:17695] = '{32'h41ad7e9a, 32'h41eb3af2, 32'h428e47b8, 32'h428ed402, 32'h426e26f7, 32'hc1f6da34, 32'hc1abef5b, 32'h42adb90b};
test_output[17688:17695] = '{32'h41ad7e9a, 32'h41eb3af2, 32'h428e47b8, 32'h428ed402, 32'h426e26f7, 32'h0, 32'h0, 32'h42adb90b};
test_input[17696:17703] = '{32'h429d184c, 32'hc1505472, 32'h429f2155, 32'hc2850081, 32'hc29d6511, 32'hc2132b83, 32'h4236e72c, 32'h42c4643e};
test_output[17696:17703] = '{32'h429d184c, 32'h0, 32'h429f2155, 32'h0, 32'h0, 32'h0, 32'h4236e72c, 32'h42c4643e};
test_input[17704:17711] = '{32'hc2947a15, 32'h424c2358, 32'hc1813a40, 32'hc2bb1a98, 32'hc15d284b, 32'hc0ccee6d, 32'h4280d456, 32'hc22aaf31};
test_output[17704:17711] = '{32'h0, 32'h424c2358, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4280d456, 32'h0};
test_input[17712:17719] = '{32'hc1d7f66e, 32'h424f97c9, 32'h41fdb9b0, 32'hc02d1420, 32'hc2b3484e, 32'h42bc80fb, 32'hc29681d5, 32'h41946a73};
test_output[17712:17719] = '{32'h0, 32'h424f97c9, 32'h41fdb9b0, 32'h0, 32'h0, 32'h42bc80fb, 32'h0, 32'h41946a73};
test_input[17720:17727] = '{32'hc28ca84b, 32'h41c9a902, 32'h3f4f224d, 32'h429f8d44, 32'h42232ebb, 32'hc2043e5a, 32'hc204f4d7, 32'h4271387b};
test_output[17720:17727] = '{32'h0, 32'h41c9a902, 32'h3f4f224d, 32'h429f8d44, 32'h42232ebb, 32'h0, 32'h0, 32'h4271387b};
test_input[17728:17735] = '{32'hc162d01f, 32'hc00bf84d, 32'h41e7f964, 32'h42bb8cde, 32'h4296d16d, 32'h426eb4ab, 32'hc13ebe5c, 32'h42a6c34e};
test_output[17728:17735] = '{32'h0, 32'h0, 32'h41e7f964, 32'h42bb8cde, 32'h4296d16d, 32'h426eb4ab, 32'h0, 32'h42a6c34e};
test_input[17736:17743] = '{32'h42a214a9, 32'hc19f72bf, 32'hc2234ef8, 32'hc28b9998, 32'h42281fd8, 32'hc1aff0ac, 32'h401b0d71, 32'hc0a44438};
test_output[17736:17743] = '{32'h42a214a9, 32'h0, 32'h0, 32'h0, 32'h42281fd8, 32'h0, 32'h401b0d71, 32'h0};
test_input[17744:17751] = '{32'hc22e62b8, 32'h41c4fcf2, 32'hc016310a, 32'hc2a4de6e, 32'hc28dcce7, 32'h403b20e1, 32'hc2996662, 32'h415d461b};
test_output[17744:17751] = '{32'h0, 32'h41c4fcf2, 32'h0, 32'h0, 32'h0, 32'h403b20e1, 32'h0, 32'h415d461b};
test_input[17752:17759] = '{32'hc235d6c6, 32'hc23df784, 32'hc1897784, 32'h4287438b, 32'hc2465f37, 32'hc26cba4b, 32'hc29fb083, 32'h41520f93};
test_output[17752:17759] = '{32'h0, 32'h0, 32'h0, 32'h4287438b, 32'h0, 32'h0, 32'h0, 32'h41520f93};
test_input[17760:17767] = '{32'h4252428a, 32'hc257fe3d, 32'h42c03d63, 32'hc05e6c49, 32'hc1a73216, 32'hc29354b7, 32'hc26dcc29, 32'hc188c9d1};
test_output[17760:17767] = '{32'h4252428a, 32'h0, 32'h42c03d63, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[17768:17775] = '{32'h42ac040c, 32'h419e9802, 32'h3f37b74a, 32'h4128e92a, 32'h42b63748, 32'h41e5fcee, 32'hc2b005f9, 32'h41fdb23a};
test_output[17768:17775] = '{32'h42ac040c, 32'h419e9802, 32'h3f37b74a, 32'h4128e92a, 32'h42b63748, 32'h41e5fcee, 32'h0, 32'h41fdb23a};
test_input[17776:17783] = '{32'hc294ec6a, 32'h40adca17, 32'h42af2a53, 32'hc1804773, 32'hc297e98d, 32'h428326d6, 32'hc05de96c, 32'h41789e2b};
test_output[17776:17783] = '{32'h0, 32'h40adca17, 32'h42af2a53, 32'h0, 32'h0, 32'h428326d6, 32'h0, 32'h41789e2b};
test_input[17784:17791] = '{32'hc22b3356, 32'h42a363fd, 32'hc2a6adb9, 32'hc2519e0d, 32'h428321d6, 32'hc29f6864, 32'h40ebe4bd, 32'hc242586a};
test_output[17784:17791] = '{32'h0, 32'h42a363fd, 32'h0, 32'h0, 32'h428321d6, 32'h0, 32'h40ebe4bd, 32'h0};
test_input[17792:17799] = '{32'h42ab3acb, 32'h419a2df4, 32'h42321993, 32'h429d29c8, 32'h424ce3c9, 32'hc25f3dc9, 32'hc159bc08, 32'h4187c4d3};
test_output[17792:17799] = '{32'h42ab3acb, 32'h419a2df4, 32'h42321993, 32'h429d29c8, 32'h424ce3c9, 32'h0, 32'h0, 32'h4187c4d3};
test_input[17800:17807] = '{32'h42c335d1, 32'hc1ed36bd, 32'h42603afa, 32'h41a9d32d, 32'hc2b50024, 32'hc2b73da6, 32'hc1e17b9e, 32'hc2bd6ced};
test_output[17800:17807] = '{32'h42c335d1, 32'h0, 32'h42603afa, 32'h41a9d32d, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[17808:17815] = '{32'h42b35090, 32'h42992d04, 32'h41e096ee, 32'h4242ee36, 32'hc2474421, 32'h420382f5, 32'hc2be610f, 32'hc2158843};
test_output[17808:17815] = '{32'h42b35090, 32'h42992d04, 32'h41e096ee, 32'h4242ee36, 32'h0, 32'h420382f5, 32'h0, 32'h0};
test_input[17816:17823] = '{32'h429943f4, 32'hc1cabeac, 32'h42c74124, 32'h40b908fc, 32'h42baf810, 32'h428e5373, 32'hc0bf7f2c, 32'h41e9752c};
test_output[17816:17823] = '{32'h429943f4, 32'h0, 32'h42c74124, 32'h40b908fc, 32'h42baf810, 32'h428e5373, 32'h0, 32'h41e9752c};
test_input[17824:17831] = '{32'h42a9f613, 32'hc111433c, 32'h42830cb6, 32'hc2826abf, 32'h41fa7c35, 32'hc29ffa5c, 32'h42841344, 32'hc2326b37};
test_output[17824:17831] = '{32'h42a9f613, 32'h0, 32'h42830cb6, 32'h0, 32'h41fa7c35, 32'h0, 32'h42841344, 32'h0};
test_input[17832:17839] = '{32'h413da27c, 32'hc2a00755, 32'h42375839, 32'h42171a54, 32'hc2c73c9b, 32'h42ae8115, 32'hc2a2d11f, 32'hc0fab41a};
test_output[17832:17839] = '{32'h413da27c, 32'h0, 32'h42375839, 32'h42171a54, 32'h0, 32'h42ae8115, 32'h0, 32'h0};
test_input[17840:17847] = '{32'hc22d592a, 32'hc2a06e99, 32'hc29645f1, 32'hc141f526, 32'h4236d331, 32'h42a2fcf4, 32'hc2adc57f, 32'hc1c6ab93};
test_output[17840:17847] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4236d331, 32'h42a2fcf4, 32'h0, 32'h0};
test_input[17848:17855] = '{32'hc282a11e, 32'hc28aa965, 32'h42ad7e7a, 32'hc27ad165, 32'hc23fb72a, 32'hc2c76f52, 32'hc22f8007, 32'h42b0df47};
test_output[17848:17855] = '{32'h0, 32'h0, 32'h42ad7e7a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b0df47};
test_input[17856:17863] = '{32'h423dd19c, 32'hc2149546, 32'hc2b33e24, 32'hc2057e62, 32'h424a9964, 32'hc2b5aa30, 32'h42145081, 32'hc2a9fa3a};
test_output[17856:17863] = '{32'h423dd19c, 32'h0, 32'h0, 32'h0, 32'h424a9964, 32'h0, 32'h42145081, 32'h0};
test_input[17864:17871] = '{32'hc22fac1d, 32'hc096dfe7, 32'hc14f08ca, 32'h41e1b293, 32'h3ebb0e51, 32'h424fc013, 32'hc1e6ed7d, 32'h4249554d};
test_output[17864:17871] = '{32'h0, 32'h0, 32'h0, 32'h41e1b293, 32'h3ebb0e51, 32'h424fc013, 32'h0, 32'h4249554d};
test_input[17872:17879] = '{32'h418cdd33, 32'hc24ea5ae, 32'h41afd179, 32'h423f1c7f, 32'h424e16e8, 32'hc2b11a9a, 32'hc1083857, 32'h42be1010};
test_output[17872:17879] = '{32'h418cdd33, 32'h0, 32'h41afd179, 32'h423f1c7f, 32'h424e16e8, 32'h0, 32'h0, 32'h42be1010};
test_input[17880:17887] = '{32'h42a108c6, 32'hc2362f88, 32'hc297f549, 32'h42354856, 32'h4286acbf, 32'h408e0efc, 32'hc23ee801, 32'hc2b89036};
test_output[17880:17887] = '{32'h42a108c6, 32'h0, 32'h0, 32'h42354856, 32'h4286acbf, 32'h408e0efc, 32'h0, 32'h0};
test_input[17888:17895] = '{32'hc1f29498, 32'hc202ea1b, 32'h42979604, 32'h41f4b2cd, 32'hc2b83a45, 32'hc23c7e93, 32'h427cf297, 32'h421fe3cf};
test_output[17888:17895] = '{32'h0, 32'h0, 32'h42979604, 32'h41f4b2cd, 32'h0, 32'h0, 32'h427cf297, 32'h421fe3cf};
test_input[17896:17903] = '{32'h40fbd412, 32'hc2a6fd00, 32'hc298c43e, 32'hbec3a36c, 32'hc272ae92, 32'hc2a781b4, 32'h42088b70, 32'h41d40815};
test_output[17896:17903] = '{32'h40fbd412, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42088b70, 32'h41d40815};
test_input[17904:17911] = '{32'h42877f97, 32'hc1067d50, 32'h424efbed, 32'h425daef5, 32'h429cd747, 32'hc20d4c20, 32'h40a57e20, 32'h42b527e2};
test_output[17904:17911] = '{32'h42877f97, 32'h0, 32'h424efbed, 32'h425daef5, 32'h429cd747, 32'h0, 32'h40a57e20, 32'h42b527e2};
test_input[17912:17919] = '{32'hc1d30fa7, 32'h41fb5808, 32'h41c004c3, 32'h41b7d74f, 32'hc218357e, 32'h42c09217, 32'hc1f1db86, 32'h42b52ed0};
test_output[17912:17919] = '{32'h0, 32'h41fb5808, 32'h41c004c3, 32'h41b7d74f, 32'h0, 32'h42c09217, 32'h0, 32'h42b52ed0};
test_input[17920:17927] = '{32'h4255e2ba, 32'hbf38431c, 32'hc1e8f45e, 32'h41fdbf85, 32'hc01bd0a9, 32'hc28527e2, 32'hc2400dd3, 32'hc289d422};
test_output[17920:17927] = '{32'h4255e2ba, 32'h0, 32'h0, 32'h41fdbf85, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[17928:17935] = '{32'hc189b47d, 32'h42af4379, 32'h41eed74b, 32'hc284c7a2, 32'h41d0d414, 32'h4214a1e8, 32'hc25f96f8, 32'hc2998dc4};
test_output[17928:17935] = '{32'h0, 32'h42af4379, 32'h41eed74b, 32'h0, 32'h41d0d414, 32'h4214a1e8, 32'h0, 32'h0};
test_input[17936:17943] = '{32'hc1f0a7d9, 32'hc2990e11, 32'hc2796063, 32'h42af31bf, 32'hc1256a62, 32'hc1f0d6cf, 32'hc1d58f45, 32'h40bedc01};
test_output[17936:17943] = '{32'h0, 32'h0, 32'h0, 32'h42af31bf, 32'h0, 32'h0, 32'h0, 32'h40bedc01};
test_input[17944:17951] = '{32'hc22e82fa, 32'h4106bddf, 32'h428ea621, 32'h4274a235, 32'h4283d50b, 32'hc287f10f, 32'h417f7c73, 32'hc24fa8af};
test_output[17944:17951] = '{32'h0, 32'h4106bddf, 32'h428ea621, 32'h4274a235, 32'h4283d50b, 32'h0, 32'h417f7c73, 32'h0};
test_input[17952:17959] = '{32'hc27382cf, 32'h421b6cb0, 32'h42018600, 32'h427cd422, 32'h42ba29e9, 32'h42a13e4a, 32'h42a37e9a, 32'h415f6bd9};
test_output[17952:17959] = '{32'h0, 32'h421b6cb0, 32'h42018600, 32'h427cd422, 32'h42ba29e9, 32'h42a13e4a, 32'h42a37e9a, 32'h415f6bd9};
test_input[17960:17967] = '{32'hc2358e72, 32'h423da13d, 32'h422e102d, 32'h42359a5c, 32'h41da0c31, 32'hc1efefc9, 32'h4256e519, 32'hc238052c};
test_output[17960:17967] = '{32'h0, 32'h423da13d, 32'h422e102d, 32'h42359a5c, 32'h41da0c31, 32'h0, 32'h4256e519, 32'h0};
test_input[17968:17975] = '{32'hc2567a84, 32'hc1a9c41f, 32'hc2ac34b7, 32'hc1e082eb, 32'hc1990d3d, 32'h417ee41f, 32'hc0217d04, 32'hc23449f7};
test_output[17968:17975] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h417ee41f, 32'h0, 32'h0};
test_input[17976:17983] = '{32'h41e53b64, 32'h4030f3b2, 32'hc2801ea7, 32'hc22a8fc8, 32'h41b4cd32, 32'h4277ac43, 32'h42ac6d1e, 32'hc1f4edae};
test_output[17976:17983] = '{32'h41e53b64, 32'h4030f3b2, 32'h0, 32'h0, 32'h41b4cd32, 32'h4277ac43, 32'h42ac6d1e, 32'h0};
test_input[17984:17991] = '{32'hc2362b6b, 32'hc1d153f7, 32'hc2968d8b, 32'hc2a51d26, 32'h41c02e96, 32'h41a11300, 32'hc2881cde, 32'h41dfc7d0};
test_output[17984:17991] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41c02e96, 32'h41a11300, 32'h0, 32'h41dfc7d0};
test_input[17992:17999] = '{32'hc1add015, 32'h428ddb28, 32'h42228f63, 32'h42a85b17, 32'hc225242d, 32'hc253755d, 32'h42c2f8e5, 32'h41cb3873};
test_output[17992:17999] = '{32'h0, 32'h428ddb28, 32'h42228f63, 32'h42a85b17, 32'h0, 32'h0, 32'h42c2f8e5, 32'h41cb3873};
test_input[18000:18007] = '{32'hc1972785, 32'hc29177dd, 32'h4072c2c9, 32'hc27ed29e, 32'h4277e9e3, 32'hc2440627, 32'hc2bb36ab, 32'h4296483d};
test_output[18000:18007] = '{32'h0, 32'h0, 32'h4072c2c9, 32'h0, 32'h4277e9e3, 32'h0, 32'h0, 32'h4296483d};
test_input[18008:18015] = '{32'hc2910f0e, 32'hbfe10e6e, 32'h41d18b8c, 32'h41bd3d6f, 32'hc28724b5, 32'hc2b0d519, 32'h41b96101, 32'h426bf84a};
test_output[18008:18015] = '{32'h0, 32'h0, 32'h41d18b8c, 32'h41bd3d6f, 32'h0, 32'h0, 32'h41b96101, 32'h426bf84a};
test_input[18016:18023] = '{32'hc1287615, 32'h42acf3c0, 32'hc0872fb2, 32'hc176e52a, 32'h4170bbce, 32'h4050334a, 32'h4284ca44, 32'hc2b6a84a};
test_output[18016:18023] = '{32'h0, 32'h42acf3c0, 32'h0, 32'h0, 32'h4170bbce, 32'h4050334a, 32'h4284ca44, 32'h0};
test_input[18024:18031] = '{32'hc256a91a, 32'hc19b10d2, 32'h42236428, 32'hc2b05430, 32'hc2a00408, 32'h427f332a, 32'h4177b797, 32'h40966978};
test_output[18024:18031] = '{32'h0, 32'h0, 32'h42236428, 32'h0, 32'h0, 32'h427f332a, 32'h4177b797, 32'h40966978};
test_input[18032:18039] = '{32'hc24fe952, 32'hc2acf582, 32'h425941fd, 32'h41827fc9, 32'hc2238c76, 32'h42959f78, 32'h427e4160, 32'hc1d83b1b};
test_output[18032:18039] = '{32'h0, 32'h0, 32'h425941fd, 32'h41827fc9, 32'h0, 32'h42959f78, 32'h427e4160, 32'h0};
test_input[18040:18047] = '{32'hc2a61234, 32'hc1d27c66, 32'h41267ed8, 32'hc172e2e8, 32'h4096eedd, 32'h4100795d, 32'hc2863215, 32'hc10cfdcf};
test_output[18040:18047] = '{32'h0, 32'h0, 32'h41267ed8, 32'h0, 32'h4096eedd, 32'h4100795d, 32'h0, 32'h0};
test_input[18048:18055] = '{32'h40ba5239, 32'hc1c7a4de, 32'hc08a6be6, 32'hc29aa59d, 32'hc2ad1068, 32'h428bdaa0, 32'hc288ebbd, 32'h420f06d9};
test_output[18048:18055] = '{32'h40ba5239, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428bdaa0, 32'h0, 32'h420f06d9};
test_input[18056:18063] = '{32'h41b023aa, 32'h42be2bc9, 32'h428a0c09, 32'h418d4c5f, 32'hc216d15c, 32'hc29b9617, 32'hc11ad4eb, 32'hc22ae559};
test_output[18056:18063] = '{32'h41b023aa, 32'h42be2bc9, 32'h428a0c09, 32'h418d4c5f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18064:18071] = '{32'hc2a82231, 32'hc263de1a, 32'h4152c749, 32'hc034b733, 32'hc2a20efd, 32'h42337c85, 32'hc2c2f936, 32'h41fb4dad};
test_output[18064:18071] = '{32'h0, 32'h0, 32'h4152c749, 32'h0, 32'h0, 32'h42337c85, 32'h0, 32'h41fb4dad};
test_input[18072:18079] = '{32'hc28e9168, 32'h42a2b717, 32'hc21d02fe, 32'h4288f938, 32'hc2031bb7, 32'hc1fa2123, 32'h4232190f, 32'hc1c58698};
test_output[18072:18079] = '{32'h0, 32'h42a2b717, 32'h0, 32'h4288f938, 32'h0, 32'h0, 32'h4232190f, 32'h0};
test_input[18080:18087] = '{32'hc29299e7, 32'hc25a16e4, 32'hc287f366, 32'h42b32afd, 32'h42ba4254, 32'h42282c4a, 32'h421ecaa3, 32'hc2b24ed9};
test_output[18080:18087] = '{32'h0, 32'h0, 32'h0, 32'h42b32afd, 32'h42ba4254, 32'h42282c4a, 32'h421ecaa3, 32'h0};
test_input[18088:18095] = '{32'hc1c24aa3, 32'h42b21b21, 32'hc102db9d, 32'hc1e11271, 32'hc29fde4f, 32'hc283e6a9, 32'h42635715, 32'h426ffbe7};
test_output[18088:18095] = '{32'h0, 32'h42b21b21, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42635715, 32'h426ffbe7};
test_input[18096:18103] = '{32'h429bf63a, 32'h41417ba3, 32'h42bcc29e, 32'h427b8005, 32'hc1fb2bbc, 32'hc1edbd9e, 32'hc16a6692, 32'h41d07e89};
test_output[18096:18103] = '{32'h429bf63a, 32'h41417ba3, 32'h42bcc29e, 32'h427b8005, 32'h0, 32'h0, 32'h0, 32'h41d07e89};
test_input[18104:18111] = '{32'h428e87f4, 32'hc24a9e6a, 32'h42bfbc24, 32'hc01422a7, 32'hc29a65e7, 32'hc2c2ad71, 32'hc1ca6e8f, 32'hc22bc1d9};
test_output[18104:18111] = '{32'h428e87f4, 32'h0, 32'h42bfbc24, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18112:18119] = '{32'hc26850a0, 32'hc2455126, 32'h42339d89, 32'hc166f689, 32'h42bb8410, 32'hc1529da7, 32'hc2863f50, 32'h425602c3};
test_output[18112:18119] = '{32'h0, 32'h0, 32'h42339d89, 32'h0, 32'h42bb8410, 32'h0, 32'h0, 32'h425602c3};
test_input[18120:18127] = '{32'hc2a5b389, 32'h422f1263, 32'h42b976f5, 32'hc2c79779, 32'hc27713a7, 32'h423ff23f, 32'h42abc473, 32'h42993328};
test_output[18120:18127] = '{32'h0, 32'h422f1263, 32'h42b976f5, 32'h0, 32'h0, 32'h423ff23f, 32'h42abc473, 32'h42993328};
test_input[18128:18135] = '{32'h428c09fe, 32'hbfe6bf10, 32'hc2bf6f38, 32'h4276682c, 32'hc2806c99, 32'h423abd15, 32'h42a54beb, 32'hc08cb1df};
test_output[18128:18135] = '{32'h428c09fe, 32'h0, 32'h0, 32'h4276682c, 32'h0, 32'h423abd15, 32'h42a54beb, 32'h0};
test_input[18136:18143] = '{32'hc2a2d33f, 32'hc2b879f6, 32'hc2220b2d, 32'hc2a2980b, 32'h4250c544, 32'hc2a639ca, 32'h42a51f8f, 32'h428c8e53};
test_output[18136:18143] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4250c544, 32'h0, 32'h42a51f8f, 32'h428c8e53};
test_input[18144:18151] = '{32'h424404d8, 32'hc29ff694, 32'hc0d5f6b2, 32'h42872587, 32'h42a34f24, 32'h42a42ec9, 32'hc05aa3ff, 32'hc169bf5b};
test_output[18144:18151] = '{32'h424404d8, 32'h0, 32'h0, 32'h42872587, 32'h42a34f24, 32'h42a42ec9, 32'h0, 32'h0};
test_input[18152:18159] = '{32'h42af5aad, 32'hc2965c0b, 32'hc0a41ebe, 32'hc21afa71, 32'h42b7210a, 32'h4218ca28, 32'h419c5280, 32'hc20b04b3};
test_output[18152:18159] = '{32'h42af5aad, 32'h0, 32'h0, 32'h0, 32'h42b7210a, 32'h4218ca28, 32'h419c5280, 32'h0};
test_input[18160:18167] = '{32'hc2020e29, 32'h42c09ba8, 32'h42598a21, 32'h4150dd4a, 32'hc2a2b3e6, 32'hc202642c, 32'hc245af77, 32'h422ea4d3};
test_output[18160:18167] = '{32'h0, 32'h42c09ba8, 32'h42598a21, 32'h4150dd4a, 32'h0, 32'h0, 32'h0, 32'h422ea4d3};
test_input[18168:18175] = '{32'h426097ea, 32'h429175ff, 32'h41ca714a, 32'hc0cec6bb, 32'hc2c20841, 32'hc284a157, 32'h423cf84a, 32'hc2401fa1};
test_output[18168:18175] = '{32'h426097ea, 32'h429175ff, 32'h41ca714a, 32'h0, 32'h0, 32'h0, 32'h423cf84a, 32'h0};
test_input[18176:18183] = '{32'hc28ddec5, 32'hc2ad4df0, 32'h42a31db7, 32'hc23368c0, 32'h41cd566a, 32'h42a9dcda, 32'h4297de40, 32'hc256ccc4};
test_output[18176:18183] = '{32'h0, 32'h0, 32'h42a31db7, 32'h0, 32'h41cd566a, 32'h42a9dcda, 32'h4297de40, 32'h0};
test_input[18184:18191] = '{32'hc138a056, 32'hc2904791, 32'h4076ad05, 32'h4149734c, 32'h403d03f8, 32'hc27f1710, 32'h42997f82, 32'h42639804};
test_output[18184:18191] = '{32'h0, 32'h0, 32'h4076ad05, 32'h4149734c, 32'h403d03f8, 32'h0, 32'h42997f82, 32'h42639804};
test_input[18192:18199] = '{32'h4227676b, 32'hc26844cc, 32'hc2a59acd, 32'h42bad6b6, 32'h42c56423, 32'h414d1f26, 32'hc0518bce, 32'h42c7330b};
test_output[18192:18199] = '{32'h4227676b, 32'h0, 32'h0, 32'h42bad6b6, 32'h42c56423, 32'h414d1f26, 32'h0, 32'h42c7330b};
test_input[18200:18207] = '{32'hc26ee6cb, 32'hc2812691, 32'hc2c3e4b4, 32'h41ea49c3, 32'h427242dd, 32'h418c66ad, 32'hc2a92949, 32'hc2177cf2};
test_output[18200:18207] = '{32'h0, 32'h0, 32'h0, 32'h41ea49c3, 32'h427242dd, 32'h418c66ad, 32'h0, 32'h0};
test_input[18208:18215] = '{32'h429437ac, 32'hc293c4f6, 32'h42c56f4e, 32'h42a64254, 32'h42a13d36, 32'hc1324b63, 32'h42c0c0cb, 32'hc249fe44};
test_output[18208:18215] = '{32'h429437ac, 32'h0, 32'h42c56f4e, 32'h42a64254, 32'h42a13d36, 32'h0, 32'h42c0c0cb, 32'h0};
test_input[18216:18223] = '{32'hc1ba48be, 32'h422fd3be, 32'h42ba75d5, 32'hc2094c76, 32'h41048636, 32'hc2561613, 32'hc10545d5, 32'h41bbfe51};
test_output[18216:18223] = '{32'h0, 32'h422fd3be, 32'h42ba75d5, 32'h0, 32'h41048636, 32'h0, 32'h0, 32'h41bbfe51};
test_input[18224:18231] = '{32'hc2ba3469, 32'hc29f23d9, 32'hc2b0d2a3, 32'h4047675a, 32'h41c75777, 32'h42a68043, 32'hc0896813, 32'h4268691f};
test_output[18224:18231] = '{32'h0, 32'h0, 32'h0, 32'h4047675a, 32'h41c75777, 32'h42a68043, 32'h0, 32'h4268691f};
test_input[18232:18239] = '{32'h422cf351, 32'h423484ae, 32'hc2af0adc, 32'hc2b64796, 32'h4284afeb, 32'h42b3d9d2, 32'hc1e9d937, 32'h4283770a};
test_output[18232:18239] = '{32'h422cf351, 32'h423484ae, 32'h0, 32'h0, 32'h4284afeb, 32'h42b3d9d2, 32'h0, 32'h4283770a};
test_input[18240:18247] = '{32'hc2aaa7f5, 32'hc1ba3e72, 32'hc2b13dd6, 32'hc2af6e9e, 32'hc1ad4d3d, 32'hc29639e7, 32'h427eda59, 32'h41c191ea};
test_output[18240:18247] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427eda59, 32'h41c191ea};
test_input[18248:18255] = '{32'hc10320e2, 32'h427d43f1, 32'hc1d1d3d1, 32'h42c6d251, 32'h42407a7d, 32'hc2998dfa, 32'hc1d9b16e, 32'hc2c7d27b};
test_output[18248:18255] = '{32'h0, 32'h427d43f1, 32'h0, 32'h42c6d251, 32'h42407a7d, 32'h0, 32'h0, 32'h0};
test_input[18256:18263] = '{32'h42b69f99, 32'h425ea2e4, 32'hc27422d1, 32'hc295a270, 32'h41f99e32, 32'hc2834e98, 32'hc25673c8, 32'h41d5aa84};
test_output[18256:18263] = '{32'h42b69f99, 32'h425ea2e4, 32'h0, 32'h0, 32'h41f99e32, 32'h0, 32'h0, 32'h41d5aa84};
test_input[18264:18271] = '{32'hc25e32d9, 32'hc2c22f9e, 32'h4139eb59, 32'h429991bf, 32'hc210c9ed, 32'hc2c4432e, 32'hc2b42347, 32'hc1ef0362};
test_output[18264:18271] = '{32'h0, 32'h0, 32'h4139eb59, 32'h429991bf, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18272:18279] = '{32'h41f1975f, 32'hbf7f1655, 32'hc2651ffb, 32'hc1d8ff8a, 32'hc2b52e49, 32'h42b5c7fc, 32'hc2563c4a, 32'h4204002c};
test_output[18272:18279] = '{32'h41f1975f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b5c7fc, 32'h0, 32'h4204002c};
test_input[18280:18287] = '{32'hc2112992, 32'hc2ba2d52, 32'h4162326b, 32'h4167a258, 32'h422c6123, 32'h41a95923, 32'hc250ccbb, 32'h4279796d};
test_output[18280:18287] = '{32'h0, 32'h0, 32'h4162326b, 32'h4167a258, 32'h422c6123, 32'h41a95923, 32'h0, 32'h4279796d};
test_input[18288:18295] = '{32'h4238ec2e, 32'h426e72fe, 32'h4224bf70, 32'h421bb22c, 32'hc1f2b13d, 32'h4097a9f8, 32'hc1ffee3d, 32'hc2c3db76};
test_output[18288:18295] = '{32'h4238ec2e, 32'h426e72fe, 32'h4224bf70, 32'h421bb22c, 32'h0, 32'h4097a9f8, 32'h0, 32'h0};
test_input[18296:18303] = '{32'hc2780939, 32'h41ec5136, 32'hc245c3a3, 32'hc254ede4, 32'hc06ae2e2, 32'h41cb148a, 32'hc2bff58a, 32'h4272bfbf};
test_output[18296:18303] = '{32'h0, 32'h41ec5136, 32'h0, 32'h0, 32'h0, 32'h41cb148a, 32'h0, 32'h4272bfbf};
test_input[18304:18311] = '{32'h429d0cd3, 32'h42546411, 32'h429010a7, 32'h4249d65d, 32'hc219286d, 32'hc26fc812, 32'hc2b1ea8a, 32'hc0793f3e};
test_output[18304:18311] = '{32'h429d0cd3, 32'h42546411, 32'h429010a7, 32'h4249d65d, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18312:18319] = '{32'hc1a164bc, 32'hc1751457, 32'hc1afd646, 32'hc1f1a193, 32'h421fb189, 32'hc28879b1, 32'h4212f579, 32'h41a2f407};
test_output[18312:18319] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h421fb189, 32'h0, 32'h4212f579, 32'h41a2f407};
test_input[18320:18327] = '{32'hc2951e90, 32'hc013834f, 32'hc26c4ae8, 32'hc1dc1540, 32'hc18e566a, 32'hc2a7ee32, 32'hbf500618, 32'hc268a84f};
test_output[18320:18327] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18328:18335] = '{32'hc2c1e5be, 32'h4207470b, 32'hc1d42146, 32'hc2beaba5, 32'h428dcb83, 32'h4201e6fe, 32'hc2b724d6, 32'h4263e4d4};
test_output[18328:18335] = '{32'h0, 32'h4207470b, 32'h0, 32'h0, 32'h428dcb83, 32'h4201e6fe, 32'h0, 32'h4263e4d4};
test_input[18336:18343] = '{32'hc1caa5d7, 32'hc25d1737, 32'h425f8e3d, 32'hc24717eb, 32'h42b2f982, 32'h425e7441, 32'h42b5f6fd, 32'hc2bff4d8};
test_output[18336:18343] = '{32'h0, 32'h0, 32'h425f8e3d, 32'h0, 32'h42b2f982, 32'h425e7441, 32'h42b5f6fd, 32'h0};
test_input[18344:18351] = '{32'hc2a6f419, 32'h42a3730e, 32'h418ff92e, 32'h42c411b8, 32'hc2205f79, 32'h42c0728a, 32'hc2955e9f, 32'h41de672b};
test_output[18344:18351] = '{32'h0, 32'h42a3730e, 32'h418ff92e, 32'h42c411b8, 32'h0, 32'h42c0728a, 32'h0, 32'h41de672b};
test_input[18352:18359] = '{32'hc25baa34, 32'h429dd16f, 32'hc2c48121, 32'h4208813e, 32'h425383b2, 32'hc1cb30b3, 32'hc2c00481, 32'hc2137c7a};
test_output[18352:18359] = '{32'h0, 32'h429dd16f, 32'h0, 32'h4208813e, 32'h425383b2, 32'h0, 32'h0, 32'h0};
test_input[18360:18367] = '{32'hc2b1bfde, 32'h405386a4, 32'hc2be8265, 32'hc1df40fb, 32'h42a0cb4d, 32'h42729add, 32'hc256776e, 32'hc2c0900b};
test_output[18360:18367] = '{32'h0, 32'h405386a4, 32'h0, 32'h0, 32'h42a0cb4d, 32'h42729add, 32'h0, 32'h0};
test_input[18368:18375] = '{32'hc21c8100, 32'hc218d395, 32'h41d233b5, 32'hc2984da5, 32'h417f3ac5, 32'hc29b03bb, 32'hc26b29aa, 32'h4266e13f};
test_output[18368:18375] = '{32'h0, 32'h0, 32'h41d233b5, 32'h0, 32'h417f3ac5, 32'h0, 32'h0, 32'h4266e13f};
test_input[18376:18383] = '{32'hc2901de8, 32'h42b67dd0, 32'hc2854f73, 32'h4298b17c, 32'h41e76b2d, 32'hc2723cd1, 32'h42ae1bf3, 32'hc28c3c76};
test_output[18376:18383] = '{32'h0, 32'h42b67dd0, 32'h0, 32'h4298b17c, 32'h41e76b2d, 32'h0, 32'h42ae1bf3, 32'h0};
test_input[18384:18391] = '{32'h40b85fd8, 32'h4209025b, 32'hc11c48df, 32'hc2c740c2, 32'h418665f8, 32'hc06f5516, 32'hc1a652d8, 32'h42b0c94d};
test_output[18384:18391] = '{32'h40b85fd8, 32'h4209025b, 32'h0, 32'h0, 32'h418665f8, 32'h0, 32'h0, 32'h42b0c94d};
test_input[18392:18399] = '{32'hc1b28e78, 32'h409b06f4, 32'hc1d40c6b, 32'hc2400eda, 32'hc2b47123, 32'h427c66da, 32'hc1ae0a8c, 32'h41d59ed6};
test_output[18392:18399] = '{32'h0, 32'h409b06f4, 32'h0, 32'h0, 32'h0, 32'h427c66da, 32'h0, 32'h41d59ed6};
test_input[18400:18407] = '{32'h41868a56, 32'hc1f10697, 32'h4268e1be, 32'hc285b72b, 32'h426837aa, 32'h41d8b041, 32'hc246f843, 32'hc03f41f4};
test_output[18400:18407] = '{32'h41868a56, 32'h0, 32'h4268e1be, 32'h0, 32'h426837aa, 32'h41d8b041, 32'h0, 32'h0};
test_input[18408:18415] = '{32'hc0d1b692, 32'h4125a780, 32'hc185d155, 32'h41dcc223, 32'h4295cd25, 32'hc18986e4, 32'hc2a0e4e0, 32'hc18ee8ec};
test_output[18408:18415] = '{32'h0, 32'h4125a780, 32'h0, 32'h41dcc223, 32'h4295cd25, 32'h0, 32'h0, 32'h0};
test_input[18416:18423] = '{32'hc20f3ef3, 32'hc178718d, 32'h4267cb56, 32'hc1f3647a, 32'h41099e6f, 32'h41942755, 32'hc18ed1f5, 32'hc1673dcb};
test_output[18416:18423] = '{32'h0, 32'h0, 32'h4267cb56, 32'h0, 32'h41099e6f, 32'h41942755, 32'h0, 32'h0};
test_input[18424:18431] = '{32'h420b6630, 32'h423f348c, 32'hc2486418, 32'hc28b7383, 32'hc13cfc45, 32'h42739424, 32'h4245b09c, 32'h4123c72d};
test_output[18424:18431] = '{32'h420b6630, 32'h423f348c, 32'h0, 32'h0, 32'h0, 32'h42739424, 32'h4245b09c, 32'h4123c72d};
test_input[18432:18439] = '{32'hc2524dac, 32'hc2844e9c, 32'hc11298e2, 32'hc1e6bfb1, 32'h422640f9, 32'hc0c32895, 32'h40f86336, 32'h4102e186};
test_output[18432:18439] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h422640f9, 32'h0, 32'h40f86336, 32'h4102e186};
test_input[18440:18447] = '{32'hc2b53402, 32'h425aa3f6, 32'h41a6fbd7, 32'h42217a16, 32'hc215af32, 32'h42ac39a7, 32'hc0da2619, 32'hc2bd4778};
test_output[18440:18447] = '{32'h0, 32'h425aa3f6, 32'h41a6fbd7, 32'h42217a16, 32'h0, 32'h42ac39a7, 32'h0, 32'h0};
test_input[18448:18455] = '{32'h4223fcf0, 32'h42c1027f, 32'hc297e8a1, 32'hc1297413, 32'hc288d755, 32'h429f034f, 32'h423e584f, 32'hc18bd62e};
test_output[18448:18455] = '{32'h4223fcf0, 32'h42c1027f, 32'h0, 32'h0, 32'h0, 32'h429f034f, 32'h423e584f, 32'h0};
test_input[18456:18463] = '{32'h42a07b31, 32'hc2a55cae, 32'h42b464ea, 32'h42a3ef50, 32'hc1bb7132, 32'h428e2c52, 32'h42859492, 32'h429e7086};
test_output[18456:18463] = '{32'h42a07b31, 32'h0, 32'h42b464ea, 32'h42a3ef50, 32'h0, 32'h428e2c52, 32'h42859492, 32'h429e7086};
test_input[18464:18471] = '{32'hc1961bd6, 32'hc2018cbf, 32'h425b1486, 32'h42bd1990, 32'hc293d609, 32'h42baff25, 32'h42833ef5, 32'hc2b4c88c};
test_output[18464:18471] = '{32'h0, 32'h0, 32'h425b1486, 32'h42bd1990, 32'h0, 32'h42baff25, 32'h42833ef5, 32'h0};
test_input[18472:18479] = '{32'hc2571b0c, 32'h4218b9c1, 32'h42acbc18, 32'hc2bf632c, 32'h4216d9ae, 32'hc2804267, 32'h42c45884, 32'h429eec52};
test_output[18472:18479] = '{32'h0, 32'h4218b9c1, 32'h42acbc18, 32'h0, 32'h4216d9ae, 32'h0, 32'h42c45884, 32'h429eec52};
test_input[18480:18487] = '{32'h4208240f, 32'h429e8378, 32'h423b1dc3, 32'hc2401127, 32'hc237350b, 32'hc29f5a0e, 32'h42b8f2ce, 32'h40aead2e};
test_output[18480:18487] = '{32'h4208240f, 32'h429e8378, 32'h423b1dc3, 32'h0, 32'h0, 32'h0, 32'h42b8f2ce, 32'h40aead2e};
test_input[18488:18495] = '{32'h404bf7dd, 32'hc25294ce, 32'h42b3146d, 32'hc272390a, 32'h410b7489, 32'h42b32f0f, 32'hc26ab614, 32'h42364015};
test_output[18488:18495] = '{32'h404bf7dd, 32'h0, 32'h42b3146d, 32'h0, 32'h410b7489, 32'h42b32f0f, 32'h0, 32'h42364015};
test_input[18496:18503] = '{32'hc23c0ad7, 32'h40ed08e5, 32'h4249fc07, 32'h425a069e, 32'hc2abdce7, 32'hc2912a6c, 32'h42a9829c, 32'hc2166da4};
test_output[18496:18503] = '{32'h0, 32'h40ed08e5, 32'h4249fc07, 32'h425a069e, 32'h0, 32'h0, 32'h42a9829c, 32'h0};
test_input[18504:18511] = '{32'hbf900f52, 32'h41f0ccb9, 32'h41356d13, 32'h41a47ea7, 32'h41cbeb5f, 32'hc20c49f3, 32'hc291ff73, 32'hc18a6734};
test_output[18504:18511] = '{32'h0, 32'h41f0ccb9, 32'h41356d13, 32'h41a47ea7, 32'h41cbeb5f, 32'h0, 32'h0, 32'h0};
test_input[18512:18519] = '{32'hc2b84017, 32'hc0cd38e1, 32'hc2497b24, 32'h4277cb56, 32'hc28d7ab5, 32'hc29068a0, 32'h4220a777, 32'h4187a5bd};
test_output[18512:18519] = '{32'h0, 32'h0, 32'h0, 32'h4277cb56, 32'h0, 32'h0, 32'h4220a777, 32'h4187a5bd};
test_input[18520:18527] = '{32'hc040c428, 32'hc1b28609, 32'h428689b5, 32'hc2add686, 32'h42a02dd6, 32'h42162bba, 32'h41caed13, 32'hc202f786};
test_output[18520:18527] = '{32'h0, 32'h0, 32'h428689b5, 32'h0, 32'h42a02dd6, 32'h42162bba, 32'h41caed13, 32'h0};
test_input[18528:18535] = '{32'hc29a2f7d, 32'h422ded08, 32'hc255384a, 32'h42c102f0, 32'hc2bd4cc4, 32'h42b5248b, 32'hc258dea2, 32'h40bc3dfb};
test_output[18528:18535] = '{32'h0, 32'h422ded08, 32'h0, 32'h42c102f0, 32'h0, 32'h42b5248b, 32'h0, 32'h40bc3dfb};
test_input[18536:18543] = '{32'hc2278677, 32'hc2b4448d, 32'hc2b65dd5, 32'hc2a341b7, 32'hc1c329b1, 32'hc26123b6, 32'hc2729c36, 32'hc25af276};
test_output[18536:18543] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18544:18551] = '{32'hc247fb6e, 32'h4290f820, 32'hc14aeca0, 32'hc26ee41f, 32'hc2138704, 32'hc2759ea5, 32'hc26f72cd, 32'h42bcae5e};
test_output[18544:18551] = '{32'h0, 32'h4290f820, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bcae5e};
test_input[18552:18559] = '{32'hc23b49eb, 32'hc2878b2c, 32'hc2c13773, 32'h41d08258, 32'h429266f1, 32'h4262edaf, 32'h4287bd63, 32'h4126842f};
test_output[18552:18559] = '{32'h0, 32'h0, 32'h0, 32'h41d08258, 32'h429266f1, 32'h4262edaf, 32'h4287bd63, 32'h4126842f};
test_input[18560:18567] = '{32'hc1fc1a34, 32'hc2adf296, 32'hc2119edf, 32'hc16ee0da, 32'hc2781ab8, 32'h42c2eb4d, 32'h416b14d2, 32'h41c63bc4};
test_output[18560:18567] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c2eb4d, 32'h416b14d2, 32'h41c63bc4};
test_input[18568:18575] = '{32'hc2948e41, 32'h42b973ad, 32'hc2b516f2, 32'h4156bafa, 32'hc27894d5, 32'h42c4a0ea, 32'h42b5d29b, 32'hc2a33e8d};
test_output[18568:18575] = '{32'h0, 32'h42b973ad, 32'h0, 32'h4156bafa, 32'h0, 32'h42c4a0ea, 32'h42b5d29b, 32'h0};
test_input[18576:18583] = '{32'h41580dad, 32'hc256b504, 32'hc2b2e28e, 32'h41a21231, 32'hc26ac926, 32'h40944824, 32'h4287731a, 32'h42721c50};
test_output[18576:18583] = '{32'h41580dad, 32'h0, 32'h0, 32'h41a21231, 32'h0, 32'h40944824, 32'h4287731a, 32'h42721c50};
test_input[18584:18591] = '{32'h422bba65, 32'h42966f24, 32'h41bc5877, 32'h409ac20a, 32'hc234a8a7, 32'hc21e0941, 32'hc1244ddd, 32'h41d2c07a};
test_output[18584:18591] = '{32'h422bba65, 32'h42966f24, 32'h41bc5877, 32'h409ac20a, 32'h0, 32'h0, 32'h0, 32'h41d2c07a};
test_input[18592:18599] = '{32'h42a74e51, 32'hc272e754, 32'hc17ecf1d, 32'h429bf060, 32'hc1b13640, 32'hc2b7615b, 32'h42552322, 32'hc29d5383};
test_output[18592:18599] = '{32'h42a74e51, 32'h0, 32'h0, 32'h429bf060, 32'h0, 32'h0, 32'h42552322, 32'h0};
test_input[18600:18607] = '{32'h42b69be2, 32'hc093bf0d, 32'h42807857, 32'h40849c28, 32'hc23574c5, 32'h4267e5ea, 32'hc273dbd6, 32'hc28375ac};
test_output[18600:18607] = '{32'h42b69be2, 32'h0, 32'h42807857, 32'h40849c28, 32'h0, 32'h4267e5ea, 32'h0, 32'h0};
test_input[18608:18615] = '{32'hc20689dd, 32'h42b6ee26, 32'hc2b4fea6, 32'hc1a505ad, 32'hc1b2a4b9, 32'h421ccd5f, 32'hc215ec8e, 32'hc2a27f48};
test_output[18608:18615] = '{32'h0, 32'h42b6ee26, 32'h0, 32'h0, 32'h0, 32'h421ccd5f, 32'h0, 32'h0};
test_input[18616:18623] = '{32'h42c5ff8d, 32'h4298dd80, 32'h4253fa53, 32'hc28598d9, 32'hc0a61c53, 32'h42bf4160, 32'h4245557a, 32'hbecfb250};
test_output[18616:18623] = '{32'h42c5ff8d, 32'h4298dd80, 32'h4253fa53, 32'h0, 32'h0, 32'h42bf4160, 32'h4245557a, 32'h0};
test_input[18624:18631] = '{32'hc1a9a7d4, 32'h41b134cc, 32'hc27fc355, 32'hc270ea60, 32'hc10e7eb4, 32'h42afb5a4, 32'hc2b7abbf, 32'hc18c06d5};
test_output[18624:18631] = '{32'h0, 32'h41b134cc, 32'h0, 32'h0, 32'h0, 32'h42afb5a4, 32'h0, 32'h0};
test_input[18632:18639] = '{32'hc29f192e, 32'hc217bb62, 32'hc2c0724c, 32'hc1f8cb7b, 32'hc2b24d96, 32'h429ecf75, 32'hc21a4985, 32'h42bb46c0};
test_output[18632:18639] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429ecf75, 32'h0, 32'h42bb46c0};
test_input[18640:18647] = '{32'h4150d706, 32'hc24fd3f1, 32'hc215e065, 32'hc232cee1, 32'h41926891, 32'h425d52a3, 32'h42b8e088, 32'h428ad4fb};
test_output[18640:18647] = '{32'h4150d706, 32'h0, 32'h0, 32'h0, 32'h41926891, 32'h425d52a3, 32'h42b8e088, 32'h428ad4fb};
test_input[18648:18655] = '{32'hbe72cc81, 32'h4289a493, 32'hc2b5a360, 32'h42221c12, 32'h42bd45d4, 32'h4250a31f, 32'h41f93aaa, 32'hc12dea31};
test_output[18648:18655] = '{32'h0, 32'h4289a493, 32'h0, 32'h42221c12, 32'h42bd45d4, 32'h4250a31f, 32'h41f93aaa, 32'h0};
test_input[18656:18663] = '{32'h42ad02e1, 32'h40ae3c46, 32'hc2a3a6e7, 32'h414eae81, 32'h41edbfed, 32'h428516ef, 32'hc1dd6773, 32'h41034570};
test_output[18656:18663] = '{32'h42ad02e1, 32'h40ae3c46, 32'h0, 32'h414eae81, 32'h41edbfed, 32'h428516ef, 32'h0, 32'h41034570};
test_input[18664:18671] = '{32'h4193b56e, 32'hc039be87, 32'hc2c54eac, 32'h4234299f, 32'hc29b69b3, 32'hc27e4973, 32'hc29e80d9, 32'hc136d732};
test_output[18664:18671] = '{32'h4193b56e, 32'h0, 32'h0, 32'h4234299f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18672:18679] = '{32'h41576b67, 32'hc1bbd413, 32'hc25fd1a1, 32'h42b91a8f, 32'h42af2eef, 32'hc2344bbc, 32'h41c71624, 32'hc2a1b0e7};
test_output[18672:18679] = '{32'h41576b67, 32'h0, 32'h0, 32'h42b91a8f, 32'h42af2eef, 32'h0, 32'h41c71624, 32'h0};
test_input[18680:18687] = '{32'h41c88cfa, 32'h4271226b, 32'h42bb4a1c, 32'h42b0bf93, 32'hc1b84119, 32'h426dc3fe, 32'hc0dba215, 32'h4258ec16};
test_output[18680:18687] = '{32'h41c88cfa, 32'h4271226b, 32'h42bb4a1c, 32'h42b0bf93, 32'h0, 32'h426dc3fe, 32'h0, 32'h4258ec16};
test_input[18688:18695] = '{32'h41c68f36, 32'hc25a397c, 32'hc280b2fa, 32'h427d1337, 32'h4281fb90, 32'h4179506d, 32'hc075f3fa, 32'hc294d55e};
test_output[18688:18695] = '{32'h41c68f36, 32'h0, 32'h0, 32'h427d1337, 32'h4281fb90, 32'h4179506d, 32'h0, 32'h0};
test_input[18696:18703] = '{32'h418dcc0a, 32'hc2909f03, 32'hc0a847f6, 32'hc1f366f6, 32'h424b1a7d, 32'h42948f32, 32'hc204ddd7, 32'h41939eb2};
test_output[18696:18703] = '{32'h418dcc0a, 32'h0, 32'h0, 32'h0, 32'h424b1a7d, 32'h42948f32, 32'h0, 32'h41939eb2};
test_input[18704:18711] = '{32'hc2c3a5b9, 32'hc221dc97, 32'hc0d0c3f1, 32'h427e8619, 32'h42b8342c, 32'hc1a584a3, 32'h41fdb0b0, 32'h3e75ed9c};
test_output[18704:18711] = '{32'h0, 32'h0, 32'h0, 32'h427e8619, 32'h42b8342c, 32'h0, 32'h41fdb0b0, 32'h3e75ed9c};
test_input[18712:18719] = '{32'h421b27a4, 32'hc20f91e8, 32'h4285b920, 32'h421b6223, 32'h41bd3f00, 32'h4224479a, 32'hc230a76a, 32'hc2939dcf};
test_output[18712:18719] = '{32'h421b27a4, 32'h0, 32'h4285b920, 32'h421b6223, 32'h41bd3f00, 32'h4224479a, 32'h0, 32'h0};
test_input[18720:18727] = '{32'hc21b3b5c, 32'hc19d0d45, 32'hc2c33701, 32'hc23bfdbf, 32'hc2459c43, 32'h429a450f, 32'h424744d5, 32'hc218136f};
test_output[18720:18727] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429a450f, 32'h424744d5, 32'h0};
test_input[18728:18735] = '{32'hc20daec4, 32'h4272fd74, 32'h415420b7, 32'hc273c264, 32'hc24263d5, 32'hc2af260b, 32'hc29b2b7a, 32'h428aaeb6};
test_output[18728:18735] = '{32'h0, 32'h4272fd74, 32'h415420b7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428aaeb6};
test_input[18736:18743] = '{32'hc28e0c3e, 32'h41caf497, 32'hc2170f3c, 32'h41103c11, 32'hc2455882, 32'h420a9300, 32'h42b3ab2b, 32'hc2597c31};
test_output[18736:18743] = '{32'h0, 32'h41caf497, 32'h0, 32'h41103c11, 32'h0, 32'h420a9300, 32'h42b3ab2b, 32'h0};
test_input[18744:18751] = '{32'hc2c223cb, 32'hc20350cf, 32'h42b04946, 32'h4254fdb6, 32'h41abf4e9, 32'h4294925d, 32'hc21c4689, 32'hc246a7b8};
test_output[18744:18751] = '{32'h0, 32'h0, 32'h42b04946, 32'h4254fdb6, 32'h41abf4e9, 32'h4294925d, 32'h0, 32'h0};
test_input[18752:18759] = '{32'h42bae221, 32'h42276238, 32'h4219cb80, 32'hc17b3b6c, 32'hc23cca44, 32'h41c8d605, 32'hc21eadbf, 32'hc2bcb4aa};
test_output[18752:18759] = '{32'h42bae221, 32'h42276238, 32'h4219cb80, 32'h0, 32'h0, 32'h41c8d605, 32'h0, 32'h0};
test_input[18760:18767] = '{32'h426738ea, 32'h424fd570, 32'hc1f628f2, 32'h426cbeb6, 32'hc1f8db8c, 32'h4211b372, 32'hc26f567a, 32'h429b2e77};
test_output[18760:18767] = '{32'h426738ea, 32'h424fd570, 32'h0, 32'h426cbeb6, 32'h0, 32'h4211b372, 32'h0, 32'h429b2e77};
test_input[18768:18775] = '{32'hc0075aad, 32'hc2ba2d3f, 32'h4156f04e, 32'hc1af0906, 32'h40f0542b, 32'hc167ce23, 32'hc2c73de9, 32'hc14c15db};
test_output[18768:18775] = '{32'h0, 32'h0, 32'h4156f04e, 32'h0, 32'h40f0542b, 32'h0, 32'h0, 32'h0};
test_input[18776:18783] = '{32'hc2acd2e2, 32'h4206dc64, 32'h419e1b30, 32'h42ae2da1, 32'hc2ae5c5f, 32'h42845a55, 32'hc1c96b76, 32'hc21cc322};
test_output[18776:18783] = '{32'h0, 32'h4206dc64, 32'h419e1b30, 32'h42ae2da1, 32'h0, 32'h42845a55, 32'h0, 32'h0};
test_input[18784:18791] = '{32'hc2c35e9b, 32'h42938bd3, 32'hbe996d04, 32'hc227584c, 32'hc10a9651, 32'h414855da, 32'hc28c0872, 32'hc2999e3e};
test_output[18784:18791] = '{32'h0, 32'h42938bd3, 32'h0, 32'h0, 32'h0, 32'h414855da, 32'h0, 32'h0};
test_input[18792:18799] = '{32'hc265a490, 32'h4206dff6, 32'h419b0b5a, 32'hc258d907, 32'hc17ed8a7, 32'hc1d3b494, 32'hc2aaa4ab, 32'hc2875fdb};
test_output[18792:18799] = '{32'h0, 32'h4206dff6, 32'h419b0b5a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18800:18807] = '{32'hc241ab36, 32'hc2831503, 32'hc182b226, 32'h419433f5, 32'hbf37ddd6, 32'hc21e40ac, 32'h41b03bbf, 32'hc04a2b8b};
test_output[18800:18807] = '{32'h0, 32'h0, 32'h0, 32'h419433f5, 32'h0, 32'h0, 32'h41b03bbf, 32'h0};
test_input[18808:18815] = '{32'hc09be739, 32'h4290bb7b, 32'h40846db5, 32'h42a3ecec, 32'h42b3779d, 32'h41790e3d, 32'h4136e52f, 32'hc1cdc300};
test_output[18808:18815] = '{32'h0, 32'h4290bb7b, 32'h40846db5, 32'h42a3ecec, 32'h42b3779d, 32'h41790e3d, 32'h4136e52f, 32'h0};
test_input[18816:18823] = '{32'h4287c9f4, 32'h42b8eb46, 32'h423774e5, 32'hc1f5b60b, 32'h427422c3, 32'hc2c420e5, 32'h423810c2, 32'h4226a200};
test_output[18816:18823] = '{32'h4287c9f4, 32'h42b8eb46, 32'h423774e5, 32'h0, 32'h427422c3, 32'h0, 32'h423810c2, 32'h4226a200};
test_input[18824:18831] = '{32'hc258e41d, 32'h4162742d, 32'h42c4771c, 32'hc263e23d, 32'hc29a9527, 32'hc1b4c40d, 32'hc21e5707, 32'hc2664655};
test_output[18824:18831] = '{32'h0, 32'h4162742d, 32'h42c4771c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18832:18839] = '{32'h425010fb, 32'hc1f17363, 32'hc0b82b06, 32'hc0dd0ad9, 32'h424ad0e2, 32'hc22b1aae, 32'hc2434039, 32'hc2178090};
test_output[18832:18839] = '{32'h425010fb, 32'h0, 32'h0, 32'h0, 32'h424ad0e2, 32'h0, 32'h0, 32'h0};
test_input[18840:18847] = '{32'h41f3af61, 32'h42951150, 32'hc28caf4d, 32'h42ad2f92, 32'h4263f955, 32'h429c15d8, 32'hc283ead9, 32'hc228039c};
test_output[18840:18847] = '{32'h41f3af61, 32'h42951150, 32'h0, 32'h42ad2f92, 32'h4263f955, 32'h429c15d8, 32'h0, 32'h0};
test_input[18848:18855] = '{32'hc2971dfe, 32'h4295a0db, 32'hc28bf22d, 32'h4226bb22, 32'hc299d1b1, 32'hc2071475, 32'hc2531be3, 32'hc2b6de3a};
test_output[18848:18855] = '{32'h0, 32'h4295a0db, 32'h0, 32'h4226bb22, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18856:18863] = '{32'h4283a615, 32'hc1edd759, 32'hc207e641, 32'hc1d2cd67, 32'hc20fc0c9, 32'hc2ae462a, 32'hc29e3dc1, 32'hc2997919};
test_output[18856:18863] = '{32'h4283a615, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18864:18871] = '{32'h429e9264, 32'h42988429, 32'h41ad7515, 32'hc2503af7, 32'h42be2aae, 32'h414ebb3c, 32'hc281f86d, 32'h4244fb33};
test_output[18864:18871] = '{32'h429e9264, 32'h42988429, 32'h41ad7515, 32'h0, 32'h42be2aae, 32'h414ebb3c, 32'h0, 32'h4244fb33};
test_input[18872:18879] = '{32'h42922842, 32'h42061d9e, 32'hc14c0e5f, 32'h428da7d5, 32'h41b9ee9e, 32'hc1ccad2d, 32'hc27980c3, 32'hc1061afb};
test_output[18872:18879] = '{32'h42922842, 32'h42061d9e, 32'h0, 32'h428da7d5, 32'h41b9ee9e, 32'h0, 32'h0, 32'h0};
test_input[18880:18887] = '{32'h42312e03, 32'h41e55857, 32'hc0bf6e18, 32'h42a10c58, 32'hc011b7f2, 32'hc00f8cd4, 32'hc1469aaf, 32'h424255dd};
test_output[18880:18887] = '{32'h42312e03, 32'h41e55857, 32'h0, 32'h42a10c58, 32'h0, 32'h0, 32'h0, 32'h424255dd};
test_input[18888:18895] = '{32'h40e00235, 32'hc2c0880d, 32'hc2522827, 32'h41fe8a95, 32'h42030a74, 32'h421f317e, 32'h4293e0ec, 32'hc220341e};
test_output[18888:18895] = '{32'h40e00235, 32'h0, 32'h0, 32'h41fe8a95, 32'h42030a74, 32'h421f317e, 32'h4293e0ec, 32'h0};
test_input[18896:18903] = '{32'h4216ef79, 32'hc2447b0e, 32'hc0a49db9, 32'hc23eb87c, 32'h420e156e, 32'hc29a82d7, 32'h41adfa86, 32'hc185392a};
test_output[18896:18903] = '{32'h4216ef79, 32'h0, 32'h0, 32'h0, 32'h420e156e, 32'h0, 32'h41adfa86, 32'h0};
test_input[18904:18911] = '{32'h3f8069dc, 32'hc22612c2, 32'hc27a5ea3, 32'hc1dbc889, 32'h428b139c, 32'hc2b49052, 32'hc2b4a48e, 32'h42c7816b};
test_output[18904:18911] = '{32'h3f8069dc, 32'h0, 32'h0, 32'h0, 32'h428b139c, 32'h0, 32'h0, 32'h42c7816b};
test_input[18912:18919] = '{32'hc2a8bc74, 32'hc1a70179, 32'h42b469c6, 32'hc22c1e33, 32'hc1971de1, 32'hc266a171, 32'h4186dd85, 32'h42c34d3f};
test_output[18912:18919] = '{32'h0, 32'h0, 32'h42b469c6, 32'h0, 32'h0, 32'h0, 32'h4186dd85, 32'h42c34d3f};
test_input[18920:18927] = '{32'h41aef436, 32'h41c6f021, 32'hc27a1da8, 32'h42b0725b, 32'h417885b0, 32'h41c048e3, 32'h40c43cc6, 32'hc1b739d9};
test_output[18920:18927] = '{32'h41aef436, 32'h41c6f021, 32'h0, 32'h42b0725b, 32'h417885b0, 32'h41c048e3, 32'h40c43cc6, 32'h0};
test_input[18928:18935] = '{32'h41d262c6, 32'h4294e3c1, 32'h42c77b65, 32'hc26bdcaf, 32'hc283f004, 32'hc25c5444, 32'hc24894db, 32'h4222e225};
test_output[18928:18935] = '{32'h41d262c6, 32'h4294e3c1, 32'h42c77b65, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4222e225};
test_input[18936:18943] = '{32'hc2b1a990, 32'h42418a7b, 32'hc224dd10, 32'hc0ba7c56, 32'hc28a4cd5, 32'h41f33d00, 32'hc20cd1f7, 32'hc0a61ed5};
test_output[18936:18943] = '{32'h0, 32'h42418a7b, 32'h0, 32'h0, 32'h0, 32'h41f33d00, 32'h0, 32'h0};
test_input[18944:18951] = '{32'h42658efe, 32'h4223116f, 32'hc2438280, 32'hc277ab8c, 32'hc289952f, 32'hc2533c69, 32'hc2038bcc, 32'hc1c6e2b0};
test_output[18944:18951] = '{32'h42658efe, 32'h4223116f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18952:18959] = '{32'hc204cfcb, 32'h414933c5, 32'hc283a846, 32'h42ac3160, 32'h428642d4, 32'hc2b407a7, 32'h42636c61, 32'h42255853};
test_output[18952:18959] = '{32'h0, 32'h414933c5, 32'h0, 32'h42ac3160, 32'h428642d4, 32'h0, 32'h42636c61, 32'h42255853};
test_input[18960:18967] = '{32'h42baed50, 32'h41c7203c, 32'h41c05cd8, 32'hc1aba1d7, 32'h423a1118, 32'hc2397df6, 32'hc2a7a3b6, 32'h4289fcc2};
test_output[18960:18967] = '{32'h42baed50, 32'h41c7203c, 32'h41c05cd8, 32'h0, 32'h423a1118, 32'h0, 32'h0, 32'h4289fcc2};
test_input[18968:18975] = '{32'hc276fd23, 32'h4140afb7, 32'h42929975, 32'h42831e7a, 32'h4126f876, 32'hc2aeed2c, 32'h42a6a447, 32'h41dbb73a};
test_output[18968:18975] = '{32'h0, 32'h4140afb7, 32'h42929975, 32'h42831e7a, 32'h4126f876, 32'h0, 32'h42a6a447, 32'h41dbb73a};
test_input[18976:18983] = '{32'hc263d6b9, 32'hc17ab122, 32'h4177bb38, 32'hc27ef5f1, 32'h421c2817, 32'h4164f1a5, 32'hc1af457d, 32'hc1db4681};
test_output[18976:18983] = '{32'h0, 32'h0, 32'h4177bb38, 32'h0, 32'h421c2817, 32'h4164f1a5, 32'h0, 32'h0};
test_input[18984:18991] = '{32'hbfcd0edb, 32'hc147a971, 32'hc2c10b7a, 32'h414dfc8d, 32'hc2b68432, 32'hc2b8e538, 32'h426f7d84, 32'h42a93437};
test_output[18984:18991] = '{32'h0, 32'h0, 32'h0, 32'h414dfc8d, 32'h0, 32'h0, 32'h426f7d84, 32'h42a93437};
test_input[18992:18999] = '{32'h42319cc1, 32'h42858d6d, 32'h400337c2, 32'h41a41890, 32'h42c7b7a6, 32'h41bb5f13, 32'h42592a0e, 32'h4092bbf4};
test_output[18992:18999] = '{32'h42319cc1, 32'h42858d6d, 32'h400337c2, 32'h41a41890, 32'h42c7b7a6, 32'h41bb5f13, 32'h42592a0e, 32'h4092bbf4};
test_input[19000:19007] = '{32'hc1b3066b, 32'h42c4fd02, 32'hc21b964e, 32'hc291bfbb, 32'h4219a2f9, 32'hc16f2f82, 32'hc2b33c44, 32'hc2aa37a3};
test_output[19000:19007] = '{32'h0, 32'h42c4fd02, 32'h0, 32'h0, 32'h4219a2f9, 32'h0, 32'h0, 32'h0};
test_input[19008:19015] = '{32'hc2a536a5, 32'h42554ed7, 32'h42b9f618, 32'h418a158b, 32'h42555415, 32'h421ff9d4, 32'hc1dabb98, 32'h423ddf65};
test_output[19008:19015] = '{32'h0, 32'h42554ed7, 32'h42b9f618, 32'h418a158b, 32'h42555415, 32'h421ff9d4, 32'h0, 32'h423ddf65};
test_input[19016:19023] = '{32'h427464e9, 32'hc2b09fb1, 32'hc2a1e272, 32'hc2b5e23b, 32'hc2bf6ec7, 32'h4228d229, 32'h42bcf4ab, 32'h42955974};
test_output[19016:19023] = '{32'h427464e9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4228d229, 32'h42bcf4ab, 32'h42955974};
test_input[19024:19031] = '{32'hc286e612, 32'hc0c23898, 32'hc28d150c, 32'h425f936b, 32'h42540810, 32'hc2a367cf, 32'hc1eaa3ad, 32'h42954455};
test_output[19024:19031] = '{32'h0, 32'h0, 32'h0, 32'h425f936b, 32'h42540810, 32'h0, 32'h0, 32'h42954455};
test_input[19032:19039] = '{32'h41aefb05, 32'h41084642, 32'hc2944779, 32'hc2a83f71, 32'hc219f7a7, 32'h421b2c67, 32'h4278b9c1, 32'hc2bb18c0};
test_output[19032:19039] = '{32'h41aefb05, 32'h41084642, 32'h0, 32'h0, 32'h0, 32'h421b2c67, 32'h4278b9c1, 32'h0};
test_input[19040:19047] = '{32'h417e2af4, 32'h41e94d3e, 32'hc268c07b, 32'hc18a5a1f, 32'h424aaf3d, 32'h41d45139, 32'hc2aa7609, 32'hc2bf0bb3};
test_output[19040:19047] = '{32'h417e2af4, 32'h41e94d3e, 32'h0, 32'h0, 32'h424aaf3d, 32'h41d45139, 32'h0, 32'h0};
test_input[19048:19055] = '{32'hc1cdb81f, 32'h42529686, 32'h4253c8a3, 32'h4205c965, 32'h411dd82e, 32'hc2900a2b, 32'hc2b1b4d3, 32'h42bd4bb1};
test_output[19048:19055] = '{32'h0, 32'h42529686, 32'h4253c8a3, 32'h4205c965, 32'h411dd82e, 32'h0, 32'h0, 32'h42bd4bb1};
test_input[19056:19063] = '{32'h425f98e3, 32'hc1888ce5, 32'h42acf7a1, 32'hc2c41514, 32'hc26500a9, 32'h426244b8, 32'h42927037, 32'hc2ab6635};
test_output[19056:19063] = '{32'h425f98e3, 32'h0, 32'h42acf7a1, 32'h0, 32'h0, 32'h426244b8, 32'h42927037, 32'h0};
test_input[19064:19071] = '{32'hc23fadcc, 32'hc292028c, 32'hc2bca012, 32'hc2b20ecd, 32'hc1cc0543, 32'hc26d0878, 32'hc2b80128, 32'hc0feab47};
test_output[19064:19071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19072:19079] = '{32'h42991485, 32'hc252bbb1, 32'h428ec7f9, 32'hc073d338, 32'hc299e969, 32'h422b711e, 32'hc270e68c, 32'h4285426d};
test_output[19072:19079] = '{32'h42991485, 32'h0, 32'h428ec7f9, 32'h0, 32'h0, 32'h422b711e, 32'h0, 32'h4285426d};
test_input[19080:19087] = '{32'h42ae626c, 32'h429e8015, 32'hc2226684, 32'h42c12b91, 32'hc2be6570, 32'h426675e4, 32'h421fccbb, 32'hc2a1eac0};
test_output[19080:19087] = '{32'h42ae626c, 32'h429e8015, 32'h0, 32'h42c12b91, 32'h0, 32'h426675e4, 32'h421fccbb, 32'h0};
test_input[19088:19095] = '{32'hc2ac497f, 32'hc225476f, 32'hc2280169, 32'h41c0f1c6, 32'h42432a48, 32'hc20e5bfd, 32'h4282c22c, 32'h40825b43};
test_output[19088:19095] = '{32'h0, 32'h0, 32'h0, 32'h41c0f1c6, 32'h42432a48, 32'h0, 32'h4282c22c, 32'h40825b43};
test_input[19096:19103] = '{32'hc2c7e6bf, 32'h427301e1, 32'hc2264f9c, 32'hc21c595b, 32'hc2babf49, 32'hc2a6f2ba, 32'hc2964a7b, 32'hc2848b98};
test_output[19096:19103] = '{32'h0, 32'h427301e1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19104:19111] = '{32'hc0e6258f, 32'h4248c3cf, 32'h42bd3725, 32'h418517b7, 32'hc0672bcb, 32'h4028775d, 32'hc20ca4c4, 32'hc2c5cc7b};
test_output[19104:19111] = '{32'h0, 32'h4248c3cf, 32'h42bd3725, 32'h418517b7, 32'h0, 32'h4028775d, 32'h0, 32'h0};
test_input[19112:19119] = '{32'h41f8c3fa, 32'h406e38c1, 32'h42568fed, 32'hc2af9689, 32'h429dc01c, 32'hc0fadacf, 32'h42858e88, 32'h3f9d832c};
test_output[19112:19119] = '{32'h41f8c3fa, 32'h406e38c1, 32'h42568fed, 32'h0, 32'h429dc01c, 32'h0, 32'h42858e88, 32'h3f9d832c};
test_input[19120:19127] = '{32'hc295aed5, 32'h428f39ab, 32'hc2760e29, 32'h42af101c, 32'hc183f9d4, 32'hc29a944b, 32'hc2521148, 32'h4286ac19};
test_output[19120:19127] = '{32'h0, 32'h428f39ab, 32'h0, 32'h42af101c, 32'h0, 32'h0, 32'h0, 32'h4286ac19};
test_input[19128:19135] = '{32'h41a82eea, 32'hc2692f6a, 32'hc28ce4ad, 32'hc27320d5, 32'h426d19f1, 32'h4159ed37, 32'hc297b0eb, 32'h41766a2e};
test_output[19128:19135] = '{32'h41a82eea, 32'h0, 32'h0, 32'h0, 32'h426d19f1, 32'h4159ed37, 32'h0, 32'h41766a2e};
test_input[19136:19143] = '{32'hc29357e9, 32'hc2a9dcb1, 32'h427b8976, 32'h419519b2, 32'hc1c5fe1b, 32'hc26f43b3, 32'h410cb8ec, 32'h428fdd9a};
test_output[19136:19143] = '{32'h0, 32'h0, 32'h427b8976, 32'h419519b2, 32'h0, 32'h0, 32'h410cb8ec, 32'h428fdd9a};
test_input[19144:19151] = '{32'hc2a59c54, 32'h4293bcf2, 32'hc2088996, 32'hc1ac0e87, 32'h419e0fe9, 32'h4289c22d, 32'h426d7179, 32'hc1c997bc};
test_output[19144:19151] = '{32'h0, 32'h4293bcf2, 32'h0, 32'h0, 32'h419e0fe9, 32'h4289c22d, 32'h426d7179, 32'h0};
test_input[19152:19159] = '{32'h420d3cdc, 32'h40ca7aaa, 32'hc280d884, 32'h42c5c919, 32'hc23fbba0, 32'hc1d25ca4, 32'hc23faedb, 32'h426827b7};
test_output[19152:19159] = '{32'h420d3cdc, 32'h40ca7aaa, 32'h0, 32'h42c5c919, 32'h0, 32'h0, 32'h0, 32'h426827b7};
test_input[19160:19167] = '{32'hc2979ecb, 32'h42aa1101, 32'hc1bdec33, 32'h42365e86, 32'hc137c064, 32'hc20729c2, 32'h429e47c6, 32'h42c79ec7};
test_output[19160:19167] = '{32'h0, 32'h42aa1101, 32'h0, 32'h42365e86, 32'h0, 32'h0, 32'h429e47c6, 32'h42c79ec7};
test_input[19168:19175] = '{32'hc2ab960b, 32'hc22eb7c1, 32'h42a31933, 32'h40e9a154, 32'hc2b08569, 32'hc2826a3e, 32'h42c1e5f8, 32'h4246335b};
test_output[19168:19175] = '{32'h0, 32'h0, 32'h42a31933, 32'h40e9a154, 32'h0, 32'h0, 32'h42c1e5f8, 32'h4246335b};
test_input[19176:19183] = '{32'hc286a209, 32'hc0994e8c, 32'h42c716ac, 32'hc0f2fed7, 32'h428818e3, 32'h424f0c34, 32'h423c8e9b, 32'h42b34f66};
test_output[19176:19183] = '{32'h0, 32'h0, 32'h42c716ac, 32'h0, 32'h428818e3, 32'h424f0c34, 32'h423c8e9b, 32'h42b34f66};
test_input[19184:19191] = '{32'hc15f6437, 32'hc2b4c8da, 32'hc2a5d3f1, 32'h42028d1c, 32'hc2041732, 32'hc1ed5598, 32'h42745e61, 32'h42b000d8};
test_output[19184:19191] = '{32'h0, 32'h0, 32'h0, 32'h42028d1c, 32'h0, 32'h0, 32'h42745e61, 32'h42b000d8};
test_input[19192:19199] = '{32'hc28f63fb, 32'h412a6766, 32'hc20fc637, 32'h407bdb17, 32'hc2a84bc6, 32'h4273188c, 32'h4259406f, 32'h42106d42};
test_output[19192:19199] = '{32'h0, 32'h412a6766, 32'h0, 32'h407bdb17, 32'h0, 32'h4273188c, 32'h4259406f, 32'h42106d42};
test_input[19200:19207] = '{32'hc291548d, 32'hc0e43300, 32'h419a4dc4, 32'hc2ae2f81, 32'hc242deb5, 32'hc1e71cba, 32'h425c350a, 32'h4292febf};
test_output[19200:19207] = '{32'h0, 32'h0, 32'h419a4dc4, 32'h0, 32'h0, 32'h0, 32'h425c350a, 32'h4292febf};
test_input[19208:19215] = '{32'hc1616ae7, 32'hc2b4f81c, 32'h42c54649, 32'hc26613af, 32'hc282ea70, 32'hc09467d2, 32'hc08e12d7, 32'h42a95638};
test_output[19208:19215] = '{32'h0, 32'h0, 32'h42c54649, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a95638};
test_input[19216:19223] = '{32'h429961ac, 32'hc1852584, 32'hc19cb618, 32'h419ba73e, 32'hc2b1a3eb, 32'hc03fcf14, 32'hc2b785ff, 32'hc20ea556};
test_output[19216:19223] = '{32'h429961ac, 32'h0, 32'h0, 32'h419ba73e, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19224:19231] = '{32'h42a5a16e, 32'h429dcf84, 32'h42c3c5ed, 32'h41541ffa, 32'h3e4a9651, 32'hc297acca, 32'hc2860a50, 32'hc2821857};
test_output[19224:19231] = '{32'h42a5a16e, 32'h429dcf84, 32'h42c3c5ed, 32'h41541ffa, 32'h3e4a9651, 32'h0, 32'h0, 32'h0};
test_input[19232:19239] = '{32'h4257e016, 32'h3f6f4f3d, 32'hc1246576, 32'h428b545c, 32'h42832996, 32'hc221ba15, 32'hc16ef32f, 32'hc284555a};
test_output[19232:19239] = '{32'h4257e016, 32'h3f6f4f3d, 32'h0, 32'h428b545c, 32'h42832996, 32'h0, 32'h0, 32'h0};
test_input[19240:19247] = '{32'h423d70b7, 32'hc1514b90, 32'h41bd053d, 32'hc179e708, 32'h429478b2, 32'hc1dc6816, 32'h418ebba2, 32'h429af059};
test_output[19240:19247] = '{32'h423d70b7, 32'h0, 32'h41bd053d, 32'h0, 32'h429478b2, 32'h0, 32'h418ebba2, 32'h429af059};
test_input[19248:19255] = '{32'h42aeef3f, 32'h4221d652, 32'hc26ece04, 32'hc29044ce, 32'h412fbfb7, 32'hc2a8caf0, 32'h42899487, 32'hc0aaa7cc};
test_output[19248:19255] = '{32'h42aeef3f, 32'h4221d652, 32'h0, 32'h0, 32'h412fbfb7, 32'h0, 32'h42899487, 32'h0};
test_input[19256:19263] = '{32'h418a5226, 32'h424ded13, 32'hc22f254c, 32'hc17a09f2, 32'h428225c6, 32'h41e94b33, 32'h41530e18, 32'h415cef8f};
test_output[19256:19263] = '{32'h418a5226, 32'h424ded13, 32'h0, 32'h0, 32'h428225c6, 32'h41e94b33, 32'h41530e18, 32'h415cef8f};
test_input[19264:19271] = '{32'hc28e0ea0, 32'hc26b7ee7, 32'h429510da, 32'hc2265503, 32'h3ec7dc8e, 32'hc2651727, 32'hc0751a4e, 32'hc22c4962};
test_output[19264:19271] = '{32'h0, 32'h0, 32'h429510da, 32'h0, 32'h3ec7dc8e, 32'h0, 32'h0, 32'h0};
test_input[19272:19279] = '{32'h40fe7316, 32'h42032712, 32'hc07bfd5b, 32'h421241c0, 32'h42338960, 32'h41e58e00, 32'h42b8da0e, 32'hc083576d};
test_output[19272:19279] = '{32'h40fe7316, 32'h42032712, 32'h0, 32'h421241c0, 32'h42338960, 32'h41e58e00, 32'h42b8da0e, 32'h0};
test_input[19280:19287] = '{32'h42337dc9, 32'hc2849b2e, 32'hc2891781, 32'hc22c8d74, 32'h411c60c8, 32'h41edd0b6, 32'h4200c4d0, 32'hc29746d9};
test_output[19280:19287] = '{32'h42337dc9, 32'h0, 32'h0, 32'h0, 32'h411c60c8, 32'h41edd0b6, 32'h4200c4d0, 32'h0};
test_input[19288:19295] = '{32'h42ad9d53, 32'hc282897f, 32'h42abafcc, 32'hc2053387, 32'hc294e70c, 32'h4068e707, 32'h4182039a, 32'h4257ad8b};
test_output[19288:19295] = '{32'h42ad9d53, 32'h0, 32'h42abafcc, 32'h0, 32'h0, 32'h4068e707, 32'h4182039a, 32'h4257ad8b};
test_input[19296:19303] = '{32'h428c4e4e, 32'hc02152ee, 32'h4291790a, 32'h4005168f, 32'h422fa445, 32'h41d06880, 32'hc2697b3a, 32'h42a0b074};
test_output[19296:19303] = '{32'h428c4e4e, 32'h0, 32'h4291790a, 32'h4005168f, 32'h422fa445, 32'h41d06880, 32'h0, 32'h42a0b074};
test_input[19304:19311] = '{32'h40bdfb1c, 32'h419c8754, 32'h428c1466, 32'h3ff9d91c, 32'h42aa934f, 32'h426653c8, 32'h4297e7a2, 32'hc182a956};
test_output[19304:19311] = '{32'h40bdfb1c, 32'h419c8754, 32'h428c1466, 32'h3ff9d91c, 32'h42aa934f, 32'h426653c8, 32'h4297e7a2, 32'h0};
test_input[19312:19319] = '{32'hc2485b9e, 32'h421830ca, 32'h4278a5f8, 32'h42a42460, 32'hc2a58e99, 32'hc20fdb4b, 32'hc23a07c5, 32'hc16c5329};
test_output[19312:19319] = '{32'h0, 32'h421830ca, 32'h4278a5f8, 32'h42a42460, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19320:19327] = '{32'h4296d8dc, 32'h41c9fab8, 32'h401ac014, 32'h41ef9258, 32'hc28d3ea2, 32'h42acad32, 32'hc29cdd01, 32'h421ff085};
test_output[19320:19327] = '{32'h4296d8dc, 32'h41c9fab8, 32'h401ac014, 32'h41ef9258, 32'h0, 32'h42acad32, 32'h0, 32'h421ff085};
test_input[19328:19335] = '{32'hc2a1399d, 32'hc284f767, 32'h42aea252, 32'h42bbc0f5, 32'h412fec6e, 32'h41c5233f, 32'hc2b255f0, 32'h418ca255};
test_output[19328:19335] = '{32'h0, 32'h0, 32'h42aea252, 32'h42bbc0f5, 32'h412fec6e, 32'h41c5233f, 32'h0, 32'h418ca255};
test_input[19336:19343] = '{32'h414addc1, 32'hc2adeaca, 32'hc2b25079, 32'hc225a048, 32'hc19072c6, 32'hc1419249, 32'hc2c13970, 32'hc0a5111b};
test_output[19336:19343] = '{32'h414addc1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19344:19351] = '{32'hc2090e0c, 32'h417caaa2, 32'hc2956c0a, 32'h41c76196, 32'h405ae53a, 32'hc21028bb, 32'h4164bf01, 32'hc1800e7a};
test_output[19344:19351] = '{32'h0, 32'h417caaa2, 32'h0, 32'h41c76196, 32'h405ae53a, 32'h0, 32'h4164bf01, 32'h0};
test_input[19352:19359] = '{32'h40568a82, 32'hc0fa6eed, 32'hc2931136, 32'hc135f50b, 32'h42bab854, 32'h421cfc52, 32'hc2bb0a42, 32'h41ed58a6};
test_output[19352:19359] = '{32'h40568a82, 32'h0, 32'h0, 32'h0, 32'h42bab854, 32'h421cfc52, 32'h0, 32'h41ed58a6};
test_input[19360:19367] = '{32'hc21bd0ad, 32'hc286f039, 32'h410d129a, 32'h42690061, 32'h414376ed, 32'hc26bcdd1, 32'h42b25e95, 32'h413f5bbc};
test_output[19360:19367] = '{32'h0, 32'h0, 32'h410d129a, 32'h42690061, 32'h414376ed, 32'h0, 32'h42b25e95, 32'h413f5bbc};
test_input[19368:19375] = '{32'h42a979e4, 32'h3fca46a8, 32'h40b605b2, 32'h428d249f, 32'h4232362c, 32'hc27e1652, 32'h42b3ab91, 32'hc1ed1a92};
test_output[19368:19375] = '{32'h42a979e4, 32'h3fca46a8, 32'h40b605b2, 32'h428d249f, 32'h4232362c, 32'h0, 32'h42b3ab91, 32'h0};
test_input[19376:19383] = '{32'hc28123eb, 32'hbf836eb3, 32'h4296f256, 32'h428381ed, 32'hc24d6738, 32'h4192c121, 32'hc11d7205, 32'h42bccab2};
test_output[19376:19383] = '{32'h0, 32'h0, 32'h4296f256, 32'h428381ed, 32'h0, 32'h4192c121, 32'h0, 32'h42bccab2};
test_input[19384:19391] = '{32'hc2824b44, 32'hc069e111, 32'hc2b10f27, 32'hc27f7e90, 32'h4206ee72, 32'hc2b90513, 32'hc2042427, 32'hc14fcd2f};
test_output[19384:19391] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4206ee72, 32'h0, 32'h0, 32'h0};
test_input[19392:19399] = '{32'h4257fc28, 32'h42b77052, 32'h4084a7c4, 32'h40af15cd, 32'hc16e5f4a, 32'h41c2d171, 32'hc2b27a44, 32'h4281d921};
test_output[19392:19399] = '{32'h4257fc28, 32'h42b77052, 32'h4084a7c4, 32'h40af15cd, 32'h0, 32'h41c2d171, 32'h0, 32'h4281d921};
test_input[19400:19407] = '{32'hc23139c3, 32'h42a846ed, 32'h424a73b1, 32'hc2be5b7f, 32'hc2146c07, 32'hc225956d, 32'hc22df982, 32'hc2915791};
test_output[19400:19407] = '{32'h0, 32'h42a846ed, 32'h424a73b1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19408:19415] = '{32'hc280be88, 32'hc2ad20a4, 32'hc2a5ed30, 32'hc2b5e666, 32'h41ef83a3, 32'h42a78b8b, 32'h4278e575, 32'h4212b4a9};
test_output[19408:19415] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41ef83a3, 32'h42a78b8b, 32'h4278e575, 32'h4212b4a9};
test_input[19416:19423] = '{32'h3f9a50a1, 32'h3fc8d3e9, 32'h4231134f, 32'h428cef89, 32'hc2297cad, 32'hc1575575, 32'hc081dc4e, 32'hc2a9afb0};
test_output[19416:19423] = '{32'h3f9a50a1, 32'h3fc8d3e9, 32'h4231134f, 32'h428cef89, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19424:19431] = '{32'hc2a7df26, 32'h42c76dc6, 32'h42b9056f, 32'h429c8402, 32'h42a5b614, 32'h41925fa4, 32'hc219ba77, 32'hc1b79eac};
test_output[19424:19431] = '{32'h0, 32'h42c76dc6, 32'h42b9056f, 32'h429c8402, 32'h42a5b614, 32'h41925fa4, 32'h0, 32'h0};
test_input[19432:19439] = '{32'h426bab3b, 32'hc269c175, 32'h41e09f54, 32'hc2862b2e, 32'h42422e2e, 32'hc25e9d70, 32'hc29d7b87, 32'hc2b9c96f};
test_output[19432:19439] = '{32'h426bab3b, 32'h0, 32'h41e09f54, 32'h0, 32'h42422e2e, 32'h0, 32'h0, 32'h0};
test_input[19440:19447] = '{32'hc2b5d33b, 32'hc248600e, 32'h41a41cba, 32'hc189a4d5, 32'h41e1073e, 32'hc0e82ef9, 32'h42b609e0, 32'hc200d0ab};
test_output[19440:19447] = '{32'h0, 32'h0, 32'h41a41cba, 32'h0, 32'h41e1073e, 32'h0, 32'h42b609e0, 32'h0};
test_input[19448:19455] = '{32'hc09acc2a, 32'h4274e460, 32'h4229f910, 32'h4272388e, 32'h4181c61f, 32'hc26eaf4b, 32'hc27fe21e, 32'h42287bd6};
test_output[19448:19455] = '{32'h0, 32'h4274e460, 32'h4229f910, 32'h4272388e, 32'h4181c61f, 32'h0, 32'h0, 32'h42287bd6};
test_input[19456:19463] = '{32'hc242fa80, 32'h41cd2999, 32'h421480f0, 32'h427fadda, 32'h427e8e9c, 32'hc1c15762, 32'hc22b56a4, 32'h40dfb32d};
test_output[19456:19463] = '{32'h0, 32'h41cd2999, 32'h421480f0, 32'h427fadda, 32'h427e8e9c, 32'h0, 32'h0, 32'h40dfb32d};
test_input[19464:19471] = '{32'h424c03c2, 32'hbf9ad5c2, 32'hc28f5030, 32'h42c11adf, 32'h42857360, 32'h408294e6, 32'h40088c34, 32'h40e8b030};
test_output[19464:19471] = '{32'h424c03c2, 32'h0, 32'h0, 32'h42c11adf, 32'h42857360, 32'h408294e6, 32'h40088c34, 32'h40e8b030};
test_input[19472:19479] = '{32'h427011e0, 32'h41eab9b6, 32'h424b0805, 32'hc1ddeec7, 32'hc1eda375, 32'h424de97c, 32'hc220fbd9, 32'h4287eb17};
test_output[19472:19479] = '{32'h427011e0, 32'h41eab9b6, 32'h424b0805, 32'h0, 32'h0, 32'h424de97c, 32'h0, 32'h4287eb17};
test_input[19480:19487] = '{32'hc29d22c4, 32'hc2872347, 32'h428d0ce7, 32'h41482816, 32'hc113f0a9, 32'hc220684b, 32'h42b80233, 32'hc29eba4e};
test_output[19480:19487] = '{32'h0, 32'h0, 32'h428d0ce7, 32'h41482816, 32'h0, 32'h0, 32'h42b80233, 32'h0};
test_input[19488:19495] = '{32'hc1abc69e, 32'h42a4a30f, 32'h3fa9b335, 32'h4233a475, 32'h419409dc, 32'h4272db38, 32'h422d2948, 32'h413156b0};
test_output[19488:19495] = '{32'h0, 32'h42a4a30f, 32'h3fa9b335, 32'h4233a475, 32'h419409dc, 32'h4272db38, 32'h422d2948, 32'h413156b0};
test_input[19496:19503] = '{32'h41e67954, 32'h42c25818, 32'h4282dc03, 32'hc103d2b2, 32'h41287531, 32'hc20e3cbe, 32'h425ace00, 32'hc2af867d};
test_output[19496:19503] = '{32'h41e67954, 32'h42c25818, 32'h4282dc03, 32'h0, 32'h41287531, 32'h0, 32'h425ace00, 32'h0};
test_input[19504:19511] = '{32'hc217b25e, 32'hc2a73674, 32'h41acbc35, 32'h425ce2e0, 32'h429edf0d, 32'hc2986fbc, 32'hc1a0ca76, 32'h427fd64d};
test_output[19504:19511] = '{32'h0, 32'h0, 32'h41acbc35, 32'h425ce2e0, 32'h429edf0d, 32'h0, 32'h0, 32'h427fd64d};
test_input[19512:19519] = '{32'hc1d6fc70, 32'hc255a77d, 32'hc20ef4a2, 32'hc1a13902, 32'hc2afe466, 32'hc2b68ea7, 32'hc2adc8bc, 32'h4221c417};
test_output[19512:19519] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4221c417};
test_input[19520:19527] = '{32'h428f778f, 32'h4284f50c, 32'h41f17acc, 32'hc1f33774, 32'hc283ff2d, 32'hc2132a4f, 32'h423ac8d9, 32'hc203e704};
test_output[19520:19527] = '{32'h428f778f, 32'h4284f50c, 32'h41f17acc, 32'h0, 32'h0, 32'h0, 32'h423ac8d9, 32'h0};
test_input[19528:19535] = '{32'hc2843480, 32'h4245c667, 32'h41b64947, 32'hc20176f1, 32'h40131d21, 32'hc296557b, 32'h422dee6f, 32'h42769501};
test_output[19528:19535] = '{32'h0, 32'h4245c667, 32'h41b64947, 32'h0, 32'h40131d21, 32'h0, 32'h422dee6f, 32'h42769501};
test_input[19536:19543] = '{32'h42b1ba49, 32'h429e4c8f, 32'h42828dd8, 32'h425a631a, 32'h4232ce56, 32'h41df7569, 32'hc205edf6, 32'hc20ce6a3};
test_output[19536:19543] = '{32'h42b1ba49, 32'h429e4c8f, 32'h42828dd8, 32'h425a631a, 32'h4232ce56, 32'h41df7569, 32'h0, 32'h0};
test_input[19544:19551] = '{32'h41aa83fa, 32'h4232d2d1, 32'h42374be3, 32'h41c59307, 32'hc0143cca, 32'hc0f0f240, 32'h402fcbd9, 32'h40e39f49};
test_output[19544:19551] = '{32'h41aa83fa, 32'h4232d2d1, 32'h42374be3, 32'h41c59307, 32'h0, 32'h0, 32'h402fcbd9, 32'h40e39f49};
test_input[19552:19559] = '{32'hc28bb1ba, 32'hc207a7eb, 32'h41e6559c, 32'hc289719b, 32'hc27080c1, 32'hbf483620, 32'hc1da5b0c, 32'h42c573c5};
test_output[19552:19559] = '{32'h0, 32'h0, 32'h41e6559c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c573c5};
test_input[19560:19567] = '{32'h41505fa1, 32'h40759c74, 32'hc26cdd00, 32'h424a6245, 32'h403ddbb9, 32'h429fddd3, 32'hc1c6ac74, 32'h4186c5c5};
test_output[19560:19567] = '{32'h41505fa1, 32'h40759c74, 32'h0, 32'h424a6245, 32'h403ddbb9, 32'h429fddd3, 32'h0, 32'h4186c5c5};
test_input[19568:19575] = '{32'h428f2dc0, 32'hc2c684ce, 32'h42a09b39, 32'hc27de43c, 32'h4175f252, 32'h42448841, 32'h411da58a, 32'h41cf3356};
test_output[19568:19575] = '{32'h428f2dc0, 32'h0, 32'h42a09b39, 32'h0, 32'h4175f252, 32'h42448841, 32'h411da58a, 32'h41cf3356};
test_input[19576:19583] = '{32'h41279fb9, 32'hc25bc652, 32'hc227bf75, 32'h4292ceca, 32'hc2c25b86, 32'h42ac31d0, 32'h42adc87f, 32'h417aca6b};
test_output[19576:19583] = '{32'h41279fb9, 32'h0, 32'h0, 32'h4292ceca, 32'h0, 32'h42ac31d0, 32'h42adc87f, 32'h417aca6b};
test_input[19584:19591] = '{32'hc24236db, 32'h42be4e3a, 32'h42ba9431, 32'h42397037, 32'hc1db41f6, 32'h429879b0, 32'h424380a2, 32'h424087e4};
test_output[19584:19591] = '{32'h0, 32'h42be4e3a, 32'h42ba9431, 32'h42397037, 32'h0, 32'h429879b0, 32'h424380a2, 32'h424087e4};
test_input[19592:19599] = '{32'hc297d849, 32'h41aa4df7, 32'hc223f6ae, 32'h42a45dd9, 32'h4227ba83, 32'hc18f8b0f, 32'hc205c238, 32'hc28a2f93};
test_output[19592:19599] = '{32'h0, 32'h41aa4df7, 32'h0, 32'h42a45dd9, 32'h4227ba83, 32'h0, 32'h0, 32'h0};
test_input[19600:19607] = '{32'hc26eccc5, 32'h422e2b14, 32'hc0c680c1, 32'h427ef5c0, 32'hc2148bb4, 32'h429fcc0e, 32'h423ca368, 32'h423aa677};
test_output[19600:19607] = '{32'h0, 32'h422e2b14, 32'h0, 32'h427ef5c0, 32'h0, 32'h429fcc0e, 32'h423ca368, 32'h423aa677};
test_input[19608:19615] = '{32'hc273bda2, 32'h42a9d4b8, 32'h4141278b, 32'hc0dfbed6, 32'hc22e0198, 32'h42c0dd01, 32'h427065a3, 32'h4298f88d};
test_output[19608:19615] = '{32'h0, 32'h42a9d4b8, 32'h4141278b, 32'h0, 32'h0, 32'h42c0dd01, 32'h427065a3, 32'h4298f88d};
test_input[19616:19623] = '{32'hc296cdaf, 32'h4260e886, 32'h42c61e1a, 32'hc11f3145, 32'h42321b36, 32'h401d10f2, 32'h42b6b044, 32'hc2026ca2};
test_output[19616:19623] = '{32'h0, 32'h4260e886, 32'h42c61e1a, 32'h0, 32'h42321b36, 32'h401d10f2, 32'h42b6b044, 32'h0};
test_input[19624:19631] = '{32'h4144cfcb, 32'h415b9e4d, 32'hc1e47c60, 32'hc15d556d, 32'h418b8d1f, 32'hc29a8254, 32'h4277f28d, 32'hc254349e};
test_output[19624:19631] = '{32'h4144cfcb, 32'h415b9e4d, 32'h0, 32'h0, 32'h418b8d1f, 32'h0, 32'h4277f28d, 32'h0};
test_input[19632:19639] = '{32'hc23df3b5, 32'hc2b5fe27, 32'h41b3e355, 32'h42873613, 32'h414649db, 32'hc278b4fb, 32'h4285c9e9, 32'hc299a3d9};
test_output[19632:19639] = '{32'h0, 32'h0, 32'h41b3e355, 32'h42873613, 32'h414649db, 32'h0, 32'h4285c9e9, 32'h0};
test_input[19640:19647] = '{32'h42a629d0, 32'h4261251c, 32'h4133ac95, 32'h42a9b79a, 32'h424e2a8b, 32'h4268aa4d, 32'h4101aed3, 32'h42bacbc6};
test_output[19640:19647] = '{32'h42a629d0, 32'h4261251c, 32'h4133ac95, 32'h42a9b79a, 32'h424e2a8b, 32'h4268aa4d, 32'h4101aed3, 32'h42bacbc6};
test_input[19648:19655] = '{32'hbfda32fe, 32'h423c324f, 32'hc24c7b6f, 32'hc21b3d14, 32'h424374da, 32'hc2419437, 32'h414818a7, 32'h424ef82c};
test_output[19648:19655] = '{32'h0, 32'h423c324f, 32'h0, 32'h0, 32'h424374da, 32'h0, 32'h414818a7, 32'h424ef82c};
test_input[19656:19663] = '{32'h4292388e, 32'h42b3b533, 32'hc281344a, 32'hc07835a4, 32'h42a331a2, 32'h4205bb90, 32'hc2b33403, 32'hc214173f};
test_output[19656:19663] = '{32'h4292388e, 32'h42b3b533, 32'h0, 32'h0, 32'h42a331a2, 32'h4205bb90, 32'h0, 32'h0};
test_input[19664:19671] = '{32'hc21e4270, 32'h42a95a4e, 32'h42ae179a, 32'h3fd36052, 32'hc28d93dc, 32'h4282d9ed, 32'h425bb2d7, 32'h425934bb};
test_output[19664:19671] = '{32'h0, 32'h42a95a4e, 32'h42ae179a, 32'h3fd36052, 32'h0, 32'h4282d9ed, 32'h425bb2d7, 32'h425934bb};
test_input[19672:19679] = '{32'h4289f03c, 32'hc2a192c9, 32'hc2072882, 32'h41273d86, 32'h429c706d, 32'hc228cefb, 32'h42180383, 32'h42544cc2};
test_output[19672:19679] = '{32'h4289f03c, 32'h0, 32'h0, 32'h41273d86, 32'h429c706d, 32'h0, 32'h42180383, 32'h42544cc2};
test_input[19680:19687] = '{32'h42a46c28, 32'h41b8b465, 32'h42715a54, 32'h425835ca, 32'hc1ac00d2, 32'hc2184a67, 32'hc2829a03, 32'hc12d9450};
test_output[19680:19687] = '{32'h42a46c28, 32'h41b8b465, 32'h42715a54, 32'h425835ca, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19688:19695] = '{32'h42b8a1fc, 32'hc2354a93, 32'h42202b09, 32'h4226fc39, 32'hc24612cd, 32'h42811ad8, 32'h412dfae5, 32'hc20b82a6};
test_output[19688:19695] = '{32'h42b8a1fc, 32'h0, 32'h42202b09, 32'h4226fc39, 32'h0, 32'h42811ad8, 32'h412dfae5, 32'h0};
test_input[19696:19703] = '{32'h42b77b39, 32'h42962522, 32'h42847d48, 32'h41d3301c, 32'hc293b451, 32'hc21b9cc3, 32'h4297a39e, 32'hc1c94fe3};
test_output[19696:19703] = '{32'h42b77b39, 32'h42962522, 32'h42847d48, 32'h41d3301c, 32'h0, 32'h0, 32'h4297a39e, 32'h0};
test_input[19704:19711] = '{32'hc2324d13, 32'h428325a0, 32'hc03d1054, 32'hc2b0b76c, 32'h4290ce22, 32'h428dc82a, 32'h41ea6658, 32'hc2c79141};
test_output[19704:19711] = '{32'h0, 32'h428325a0, 32'h0, 32'h0, 32'h4290ce22, 32'h428dc82a, 32'h41ea6658, 32'h0};
test_input[19712:19719] = '{32'hc0588db0, 32'h40cb07c9, 32'h421efa2b, 32'hc2128e38, 32'h41416206, 32'h40e17a7c, 32'hc2a1043b, 32'hc125671b};
test_output[19712:19719] = '{32'h0, 32'h40cb07c9, 32'h421efa2b, 32'h0, 32'h41416206, 32'h40e17a7c, 32'h0, 32'h0};
test_input[19720:19727] = '{32'hc23e8018, 32'h41a0a351, 32'hc2b632c3, 32'hc2666c0e, 32'h429a7c81, 32'hc19f3372, 32'h41cc495c, 32'hc226be2f};
test_output[19720:19727] = '{32'h0, 32'h41a0a351, 32'h0, 32'h0, 32'h429a7c81, 32'h0, 32'h41cc495c, 32'h0};
test_input[19728:19735] = '{32'h426d3680, 32'hc230c1d5, 32'h423f34bc, 32'hc2399e61, 32'h425fb76e, 32'h418c9020, 32'h42a7b0b8, 32'hc21b1225};
test_output[19728:19735] = '{32'h426d3680, 32'h0, 32'h423f34bc, 32'h0, 32'h425fb76e, 32'h418c9020, 32'h42a7b0b8, 32'h0};
test_input[19736:19743] = '{32'hc1eb560e, 32'hc29ede01, 32'hc2716f4b, 32'hc0c8b918, 32'h41edc6c6, 32'hc1caab17, 32'hc2c76e99, 32'hc2747022};
test_output[19736:19743] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41edc6c6, 32'h0, 32'h0, 32'h0};
test_input[19744:19751] = '{32'hc229e898, 32'h42ad7c33, 32'hc1d1efe1, 32'hc25c271f, 32'hc266f2db, 32'h42b667bd, 32'hc1eaaa35, 32'h429fc17a};
test_output[19744:19751] = '{32'h0, 32'h42ad7c33, 32'h0, 32'h0, 32'h0, 32'h42b667bd, 32'h0, 32'h429fc17a};
test_input[19752:19759] = '{32'h42347dd0, 32'h423d0374, 32'h41296c7c, 32'h42bfa7fa, 32'h4233d2f4, 32'h42bc8626, 32'hc191ec6e, 32'hc1b2e00e};
test_output[19752:19759] = '{32'h42347dd0, 32'h423d0374, 32'h41296c7c, 32'h42bfa7fa, 32'h4233d2f4, 32'h42bc8626, 32'h0, 32'h0};
test_input[19760:19767] = '{32'hc27c4963, 32'h4036e967, 32'hc29dfcf3, 32'h4280894d, 32'hc28e796c, 32'hc28cfac3, 32'h42b8943c, 32'hc2adc419};
test_output[19760:19767] = '{32'h0, 32'h4036e967, 32'h0, 32'h4280894d, 32'h0, 32'h0, 32'h42b8943c, 32'h0};
test_input[19768:19775] = '{32'hbfbdf950, 32'h41909a6f, 32'hc28cd362, 32'hc2a99258, 32'hc119094c, 32'h424f42fd, 32'h41dc7f00, 32'h42906fb1};
test_output[19768:19775] = '{32'h0, 32'h41909a6f, 32'h0, 32'h0, 32'h0, 32'h424f42fd, 32'h41dc7f00, 32'h42906fb1};
test_input[19776:19783] = '{32'hc2448675, 32'h42833174, 32'h42795043, 32'h4174c9bc, 32'hc1d8d450, 32'hc29a1036, 32'h424c8a98, 32'hc291a5ca};
test_output[19776:19783] = '{32'h0, 32'h42833174, 32'h42795043, 32'h4174c9bc, 32'h0, 32'h0, 32'h424c8a98, 32'h0};
test_input[19784:19791] = '{32'hc2b473f7, 32'hc1341c39, 32'h42598354, 32'hc2c224d3, 32'h42b893b6, 32'hc19f1abe, 32'h429a3b2f, 32'h409fdd6e};
test_output[19784:19791] = '{32'h0, 32'h0, 32'h42598354, 32'h0, 32'h42b893b6, 32'h0, 32'h429a3b2f, 32'h409fdd6e};
test_input[19792:19799] = '{32'h42642899, 32'hc1092b01, 32'hc1cbd733, 32'hc2484e35, 32'hc1b52d13, 32'hc228b27b, 32'hc1f01657, 32'h41f5eb69};
test_output[19792:19799] = '{32'h42642899, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f5eb69};
test_input[19800:19807] = '{32'h4227bdff, 32'hc228b998, 32'hc28ca70d, 32'h42a89cc8, 32'h421d5d8c, 32'h40d917c2, 32'h41a054f8, 32'h428f1bd2};
test_output[19800:19807] = '{32'h4227bdff, 32'h0, 32'h0, 32'h42a89cc8, 32'h421d5d8c, 32'h40d917c2, 32'h41a054f8, 32'h428f1bd2};
test_input[19808:19815] = '{32'hc289a1ad, 32'h4187f53f, 32'h42c26ff5, 32'h4291be39, 32'hc2c2097c, 32'hc284dc52, 32'hc1b65e17, 32'h42c69814};
test_output[19808:19815] = '{32'h0, 32'h4187f53f, 32'h42c26ff5, 32'h4291be39, 32'h0, 32'h0, 32'h0, 32'h42c69814};
test_input[19816:19823] = '{32'hc1f35d52, 32'hc29a9e92, 32'h429203c1, 32'h4185cc04, 32'hc1ce457f, 32'h429455a8, 32'hc194ffd6, 32'h421a8b49};
test_output[19816:19823] = '{32'h0, 32'h0, 32'h429203c1, 32'h4185cc04, 32'h0, 32'h429455a8, 32'h0, 32'h421a8b49};
test_input[19824:19831] = '{32'h4043aafb, 32'hc04b7108, 32'h42a5f535, 32'h41e8a857, 32'hc2b81d7d, 32'h420870d9, 32'h40fa5bcf, 32'h4167f9ee};
test_output[19824:19831] = '{32'h4043aafb, 32'h0, 32'h42a5f535, 32'h41e8a857, 32'h0, 32'h420870d9, 32'h40fa5bcf, 32'h4167f9ee};
test_input[19832:19839] = '{32'hc28c6a79, 32'hc22e9242, 32'hc0917983, 32'h41cebda7, 32'hc2c524d5, 32'h42c51b69, 32'h4286bcf1, 32'hc2984e3d};
test_output[19832:19839] = '{32'h0, 32'h0, 32'h0, 32'h41cebda7, 32'h0, 32'h42c51b69, 32'h4286bcf1, 32'h0};
test_input[19840:19847] = '{32'hc216d084, 32'hc28b02bd, 32'h41d251fb, 32'hc23126b2, 32'h41b5b576, 32'hc11f7c0e, 32'hc1edb3ff, 32'hc2c6864f};
test_output[19840:19847] = '{32'h0, 32'h0, 32'h41d251fb, 32'h0, 32'h41b5b576, 32'h0, 32'h0, 32'h0};
test_input[19848:19855] = '{32'h42c78267, 32'hc233dab0, 32'h41dfb090, 32'h42b0684f, 32'h42abb43a, 32'h42490294, 32'h42b10af8, 32'hc0a86061};
test_output[19848:19855] = '{32'h42c78267, 32'h0, 32'h41dfb090, 32'h42b0684f, 32'h42abb43a, 32'h42490294, 32'h42b10af8, 32'h0};
test_input[19856:19863] = '{32'h40e0b008, 32'h42533446, 32'hc253df40, 32'h41182e93, 32'h429470b4, 32'h4215719b, 32'h4204da6b, 32'hc239fee5};
test_output[19856:19863] = '{32'h40e0b008, 32'h42533446, 32'h0, 32'h41182e93, 32'h429470b4, 32'h4215719b, 32'h4204da6b, 32'h0};
test_input[19864:19871] = '{32'hc1962362, 32'h409ea885, 32'h4288c121, 32'h41f1bc88, 32'h4220e587, 32'h425fd5f6, 32'hc28aea67, 32'hc27f1c5e};
test_output[19864:19871] = '{32'h0, 32'h409ea885, 32'h4288c121, 32'h41f1bc88, 32'h4220e587, 32'h425fd5f6, 32'h0, 32'h0};
test_input[19872:19879] = '{32'hc29cbf1a, 32'h4282d65c, 32'hc120fb10, 32'hc23dd049, 32'hc10495a4, 32'hc289de7c, 32'h4299de76, 32'hc103687b};
test_output[19872:19879] = '{32'h0, 32'h4282d65c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4299de76, 32'h0};
test_input[19880:19887] = '{32'h4199c3b0, 32'hc2b10654, 32'hc2ad9b55, 32'h420f4dfd, 32'hc1313156, 32'h420486a9, 32'hc2334d2e, 32'hc2aa6444};
test_output[19880:19887] = '{32'h4199c3b0, 32'h0, 32'h0, 32'h420f4dfd, 32'h0, 32'h420486a9, 32'h0, 32'h0};
test_input[19888:19895] = '{32'h42228e0d, 32'h429ee437, 32'h42335ca5, 32'h42c4a5aa, 32'h4267823f, 32'h42031ba2, 32'h41ba4158, 32'hc2c6d3d2};
test_output[19888:19895] = '{32'h42228e0d, 32'h429ee437, 32'h42335ca5, 32'h42c4a5aa, 32'h4267823f, 32'h42031ba2, 32'h41ba4158, 32'h0};
test_input[19896:19903] = '{32'hc2c69a2c, 32'hc1bec4ae, 32'hc215a7d5, 32'h42288c52, 32'h426189d6, 32'hc20ec9b5, 32'hc2866a2a, 32'h428769a1};
test_output[19896:19903] = '{32'h0, 32'h0, 32'h0, 32'h42288c52, 32'h426189d6, 32'h0, 32'h0, 32'h428769a1};
test_input[19904:19911] = '{32'hc29dfda2, 32'h42749bab, 32'hc1c3f145, 32'h4139dac2, 32'h429399d3, 32'h41e7a4c9, 32'h424da4cb, 32'h4252f730};
test_output[19904:19911] = '{32'h0, 32'h42749bab, 32'h0, 32'h4139dac2, 32'h429399d3, 32'h41e7a4c9, 32'h424da4cb, 32'h4252f730};
test_input[19912:19919] = '{32'h42950167, 32'h412bd196, 32'h412d7947, 32'h42492765, 32'hc1a02c2d, 32'hc255be8a, 32'hc20d5859, 32'hc2b46b90};
test_output[19912:19919] = '{32'h42950167, 32'h412bd196, 32'h412d7947, 32'h42492765, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19920:19927] = '{32'h427b86e7, 32'h4284c5fd, 32'h41c98ac6, 32'h41afea42, 32'hc1a24b39, 32'h42a56f50, 32'h4125f5d8, 32'hc2ab80ad};
test_output[19920:19927] = '{32'h427b86e7, 32'h4284c5fd, 32'h41c98ac6, 32'h41afea42, 32'h0, 32'h42a56f50, 32'h4125f5d8, 32'h0};
test_input[19928:19935] = '{32'hc2aca69e, 32'hc196b7e8, 32'hc11c8249, 32'h418ffa9b, 32'h42987052, 32'hc08b950f, 32'h415f9de7, 32'h4274c91b};
test_output[19928:19935] = '{32'h0, 32'h0, 32'h0, 32'h418ffa9b, 32'h42987052, 32'h0, 32'h415f9de7, 32'h4274c91b};
test_input[19936:19943] = '{32'h42a12077, 32'hc19576f6, 32'h42483555, 32'hc288e505, 32'h425e4c0f, 32'hc211c037, 32'h420d9e27, 32'h42b3d66f};
test_output[19936:19943] = '{32'h42a12077, 32'h0, 32'h42483555, 32'h0, 32'h425e4c0f, 32'h0, 32'h420d9e27, 32'h42b3d66f};
test_input[19944:19951] = '{32'h429ce536, 32'hc22169c3, 32'h42a6a16d, 32'h426ae466, 32'h41c1d2a3, 32'h42bc83a4, 32'h41e33e6a, 32'hc0525555};
test_output[19944:19951] = '{32'h429ce536, 32'h0, 32'h42a6a16d, 32'h426ae466, 32'h41c1d2a3, 32'h42bc83a4, 32'h41e33e6a, 32'h0};
test_input[19952:19959] = '{32'hc2ba7aff, 32'hc222d787, 32'h42660b0a, 32'hc231d54a, 32'hc23f3551, 32'h42a01da2, 32'hc20fdda1, 32'hc24424e7};
test_output[19952:19959] = '{32'h0, 32'h0, 32'h42660b0a, 32'h0, 32'h0, 32'h42a01da2, 32'h0, 32'h0};
test_input[19960:19967] = '{32'hc2c6d7d7, 32'h4182bbcc, 32'hc21aa940, 32'hc1fa2477, 32'h41af13c7, 32'hc25a48d9, 32'hc236c7b4, 32'h4214a61c};
test_output[19960:19967] = '{32'h0, 32'h4182bbcc, 32'h0, 32'h0, 32'h41af13c7, 32'h0, 32'h0, 32'h4214a61c};
test_input[19968:19975] = '{32'h41a09e32, 32'hc2078492, 32'hc280c6bb, 32'hc127efaf, 32'h422dbd86, 32'h414047f4, 32'hc20082d4, 32'h4295ad94};
test_output[19968:19975] = '{32'h41a09e32, 32'h0, 32'h0, 32'h0, 32'h422dbd86, 32'h414047f4, 32'h0, 32'h4295ad94};
test_input[19976:19983] = '{32'h41925131, 32'h42b5fd6f, 32'h41aa4bd0, 32'h427c1f08, 32'h427c94a8, 32'h4112e33c, 32'hc18ff288, 32'h41a5b501};
test_output[19976:19983] = '{32'h41925131, 32'h42b5fd6f, 32'h41aa4bd0, 32'h427c1f08, 32'h427c94a8, 32'h4112e33c, 32'h0, 32'h41a5b501};
test_input[19984:19991] = '{32'h40ed387b, 32'h4058386a, 32'h423e3a15, 32'h42034cc7, 32'h4294a68d, 32'h420a3971, 32'hc2a434fd, 32'hc2175681};
test_output[19984:19991] = '{32'h40ed387b, 32'h4058386a, 32'h423e3a15, 32'h42034cc7, 32'h4294a68d, 32'h420a3971, 32'h0, 32'h0};
test_input[19992:19999] = '{32'hc29d466a, 32'hc2a90c2d, 32'h4290ae8b, 32'hc10fffc9, 32'hc2a02458, 32'hc22b8213, 32'hc23cc22c, 32'hc1e7c885};
test_output[19992:19999] = '{32'h0, 32'h0, 32'h4290ae8b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20000:20007] = '{32'hc1c0e8dc, 32'hc12ad414, 32'h41fdcd3e, 32'hc2b90099, 32'h42764056, 32'hc27cd682, 32'hc0da99f8, 32'h42413ba0};
test_output[20000:20007] = '{32'h0, 32'h0, 32'h41fdcd3e, 32'h0, 32'h42764056, 32'h0, 32'h0, 32'h42413ba0};
test_input[20008:20015] = '{32'hc1239089, 32'hc17cb87c, 32'h41f2bb18, 32'h42af3339, 32'h42bda65d, 32'hc1cee8fb, 32'hc227559a, 32'hc28f84cb};
test_output[20008:20015] = '{32'h0, 32'h0, 32'h41f2bb18, 32'h42af3339, 32'h42bda65d, 32'h0, 32'h0, 32'h0};
test_input[20016:20023] = '{32'h42bc4e54, 32'hc2592e1f, 32'h3e0ebcfa, 32'hc2096ccc, 32'hc235a355, 32'hc293ba01, 32'hc2a2e52c, 32'h42556c31};
test_output[20016:20023] = '{32'h42bc4e54, 32'h0, 32'h3e0ebcfa, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42556c31};
test_input[20024:20031] = '{32'h422a80c6, 32'hc28dcadd, 32'h42c7383b, 32'hc12bdfdc, 32'hc18337a5, 32'hc1f8d671, 32'hc218073a, 32'h426bdbc9};
test_output[20024:20031] = '{32'h422a80c6, 32'h0, 32'h42c7383b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426bdbc9};
test_input[20032:20039] = '{32'hc24eed3f, 32'hc04779e0, 32'hc231efb8, 32'hc2580232, 32'hc283fe31, 32'hc18b6b78, 32'h428796fc, 32'h413d490f};
test_output[20032:20039] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428796fc, 32'h413d490f};
test_input[20040:20047] = '{32'h42a067df, 32'hc277e6cd, 32'h424e41a8, 32'hc1d08444, 32'h428d3460, 32'hc22a4219, 32'h42be5fd5, 32'h420008ba};
test_output[20040:20047] = '{32'h42a067df, 32'h0, 32'h424e41a8, 32'h0, 32'h428d3460, 32'h0, 32'h42be5fd5, 32'h420008ba};
test_input[20048:20055] = '{32'h42b2f91c, 32'hc20ff447, 32'hc2b998de, 32'hc246180d, 32'h427553ea, 32'hc2a59c54, 32'hc2943c19, 32'hc16217af};
test_output[20048:20055] = '{32'h42b2f91c, 32'h0, 32'h0, 32'h0, 32'h427553ea, 32'h0, 32'h0, 32'h0};
test_input[20056:20063] = '{32'hc1f33eae, 32'h4294c212, 32'hc01319d5, 32'hc1951cf7, 32'hc211258f, 32'hc2ad8512, 32'h42310f1d, 32'hc0f849fb};
test_output[20056:20063] = '{32'h0, 32'h4294c212, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42310f1d, 32'h0};
test_input[20064:20071] = '{32'hc298951c, 32'hc1e48988, 32'h42a7aef6, 32'hc2bedf81, 32'hc1f06014, 32'hc2008afa, 32'hbfd9dc20, 32'hc16a4f6d};
test_output[20064:20071] = '{32'h0, 32'h0, 32'h42a7aef6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20072:20079] = '{32'h4249279b, 32'h42c7a70a, 32'h42ae4605, 32'h423dedb2, 32'h41ec0c92, 32'h41d9c684, 32'hc2a4e7ba, 32'hc2b81862};
test_output[20072:20079] = '{32'h4249279b, 32'h42c7a70a, 32'h42ae4605, 32'h423dedb2, 32'h41ec0c92, 32'h41d9c684, 32'h0, 32'h0};
test_input[20080:20087] = '{32'hc237e9f1, 32'hc111777a, 32'hc1542e22, 32'h4293d2fb, 32'h419843a1, 32'hc2593ea2, 32'hc1f99e57, 32'hc2b21855};
test_output[20080:20087] = '{32'h0, 32'h0, 32'h0, 32'h4293d2fb, 32'h419843a1, 32'h0, 32'h0, 32'h0};
test_input[20088:20095] = '{32'h4240b782, 32'h42640df6, 32'hc291cd1c, 32'hc2bdec80, 32'h40defd28, 32'h4211b0fc, 32'h41f251ef, 32'h42b4346c};
test_output[20088:20095] = '{32'h4240b782, 32'h42640df6, 32'h0, 32'h0, 32'h40defd28, 32'h4211b0fc, 32'h41f251ef, 32'h42b4346c};
test_input[20096:20103] = '{32'hc29bd8d6, 32'h42196626, 32'hc2bf8940, 32'hc2795781, 32'hc192bf1c, 32'hc180b117, 32'h42194aa6, 32'h42afcef5};
test_output[20096:20103] = '{32'h0, 32'h42196626, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42194aa6, 32'h42afcef5};
test_input[20104:20111] = '{32'hc2aa90ce, 32'h42220a20, 32'hc1b98b7a, 32'h42890d5e, 32'hc2ba5ec9, 32'h429cf039, 32'hc2a3d13f, 32'hc18355db};
test_output[20104:20111] = '{32'h0, 32'h42220a20, 32'h0, 32'h42890d5e, 32'h0, 32'h429cf039, 32'h0, 32'h0};
test_input[20112:20119] = '{32'h42302466, 32'h425d69a8, 32'h426f6985, 32'hc2a3cc3a, 32'hc243b4a6, 32'hc2b30003, 32'hc19a992f, 32'hc185468e};
test_output[20112:20119] = '{32'h42302466, 32'h425d69a8, 32'h426f6985, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20120:20127] = '{32'hc03382f8, 32'h42937e50, 32'hc29841a4, 32'h41ccc8d6, 32'h41b0a28c, 32'h42059e83, 32'hc242069c, 32'h42c6a20b};
test_output[20120:20127] = '{32'h0, 32'h42937e50, 32'h0, 32'h41ccc8d6, 32'h41b0a28c, 32'h42059e83, 32'h0, 32'h42c6a20b};
test_input[20128:20135] = '{32'h41bf3b5a, 32'h41837530, 32'hc2b64fe7, 32'hc2153611, 32'hc1c1f2da, 32'h4113509a, 32'hc2243d71, 32'hc244069b};
test_output[20128:20135] = '{32'h41bf3b5a, 32'h41837530, 32'h0, 32'h0, 32'h0, 32'h4113509a, 32'h0, 32'h0};
test_input[20136:20143] = '{32'hc2ad5fcd, 32'h4262cd32, 32'hc2c3926e, 32'h420c7c89, 32'h41fe57fd, 32'hc17396f9, 32'h40ed7230, 32'hc19c7262};
test_output[20136:20143] = '{32'h0, 32'h4262cd32, 32'h0, 32'h420c7c89, 32'h41fe57fd, 32'h0, 32'h40ed7230, 32'h0};
test_input[20144:20151] = '{32'h42b7b060, 32'h4131150d, 32'h42a26c64, 32'h401d8280, 32'hc2800772, 32'h41ac7402, 32'hc2b7b630, 32'h410808dd};
test_output[20144:20151] = '{32'h42b7b060, 32'h4131150d, 32'h42a26c64, 32'h401d8280, 32'h0, 32'h41ac7402, 32'h0, 32'h410808dd};
test_input[20152:20159] = '{32'hc0295089, 32'hc1f86a46, 32'h40e7e695, 32'h427decb3, 32'h42b4bd69, 32'hc2a5f4e4, 32'h4235a0b6, 32'hc0fd6278};
test_output[20152:20159] = '{32'h0, 32'h0, 32'h40e7e695, 32'h427decb3, 32'h42b4bd69, 32'h0, 32'h4235a0b6, 32'h0};
test_input[20160:20167] = '{32'h422a563c, 32'hc251226b, 32'h426ca3ca, 32'h423dc8d4, 32'h429ff31c, 32'hc2c10873, 32'h42bb96b2, 32'hc0e2eef4};
test_output[20160:20167] = '{32'h422a563c, 32'h0, 32'h426ca3ca, 32'h423dc8d4, 32'h429ff31c, 32'h0, 32'h42bb96b2, 32'h0};
test_input[20168:20175] = '{32'hc204b935, 32'h41e0330d, 32'h40b15bb7, 32'hc0fdc0aa, 32'h42aeb382, 32'hc223e9bc, 32'hc1d8504b, 32'hc13e5071};
test_output[20168:20175] = '{32'h0, 32'h41e0330d, 32'h40b15bb7, 32'h0, 32'h42aeb382, 32'h0, 32'h0, 32'h0};
test_input[20176:20183] = '{32'hc1e86e80, 32'hc2a2d06e, 32'hc147d114, 32'h4295f1ac, 32'hc158581f, 32'h419a94be, 32'h420c2f5c, 32'h42ad4f39};
test_output[20176:20183] = '{32'h0, 32'h0, 32'h0, 32'h4295f1ac, 32'h0, 32'h419a94be, 32'h420c2f5c, 32'h42ad4f39};
test_input[20184:20191] = '{32'h40fa94da, 32'h4294c1eb, 32'hc03f4b0f, 32'h42375339, 32'h428e76ed, 32'h42a58e85, 32'h429faf59, 32'h42a442b5};
test_output[20184:20191] = '{32'h40fa94da, 32'h4294c1eb, 32'h0, 32'h42375339, 32'h428e76ed, 32'h42a58e85, 32'h429faf59, 32'h42a442b5};
test_input[20192:20199] = '{32'h429d04dc, 32'h42823191, 32'h429572b8, 32'hc204a6d2, 32'hc2b8c260, 32'h423fbadc, 32'hc29436d2, 32'hc25bcba1};
test_output[20192:20199] = '{32'h429d04dc, 32'h42823191, 32'h429572b8, 32'h0, 32'h0, 32'h423fbadc, 32'h0, 32'h0};
test_input[20200:20207] = '{32'h40b684b1, 32'hc1be8bca, 32'h42a3577f, 32'hc29cb252, 32'hc218808c, 32'hc29745ae, 32'h428f807f, 32'h41c0481b};
test_output[20200:20207] = '{32'h40b684b1, 32'h0, 32'h42a3577f, 32'h0, 32'h0, 32'h0, 32'h428f807f, 32'h41c0481b};
test_input[20208:20215] = '{32'h4256ece5, 32'h40cf0859, 32'h4180eefc, 32'hc29d4dd6, 32'hc0241a5f, 32'hc284c71b, 32'h409f928a, 32'h41d527d2};
test_output[20208:20215] = '{32'h4256ece5, 32'h40cf0859, 32'h4180eefc, 32'h0, 32'h0, 32'h0, 32'h409f928a, 32'h41d527d2};
test_input[20216:20223] = '{32'h41b5dc1f, 32'hc28a1196, 32'h4232912d, 32'hc1e8ba1a, 32'h42c63fae, 32'hc2c36fdb, 32'hc235f46e, 32'h4185cd38};
test_output[20216:20223] = '{32'h41b5dc1f, 32'h0, 32'h4232912d, 32'h0, 32'h42c63fae, 32'h0, 32'h0, 32'h4185cd38};
test_input[20224:20231] = '{32'hc2042c02, 32'h42be5b44, 32'h42367fe0, 32'hbe0ced79, 32'h42926b58, 32'h41a44c98, 32'hc2369264, 32'hc2bca958};
test_output[20224:20231] = '{32'h0, 32'h42be5b44, 32'h42367fe0, 32'h0, 32'h42926b58, 32'h41a44c98, 32'h0, 32'h0};
test_input[20232:20239] = '{32'h4139f2f2, 32'h42af0213, 32'h41a3886f, 32'h4240ca1c, 32'h426cea2a, 32'hc20877f2, 32'h418a0194, 32'h41d2994c};
test_output[20232:20239] = '{32'h4139f2f2, 32'h42af0213, 32'h41a3886f, 32'h4240ca1c, 32'h426cea2a, 32'h0, 32'h418a0194, 32'h41d2994c};
test_input[20240:20247] = '{32'h4257fc84, 32'hc28be591, 32'hc23ba254, 32'hc21ba3ce, 32'hc2adafe3, 32'hc11fd9ec, 32'hc2097ca3, 32'hc2bd6d44};
test_output[20240:20247] = '{32'h4257fc84, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20248:20255] = '{32'hc2694f39, 32'hc28bea24, 32'hc26230db, 32'h40dfc44f, 32'hc1d4c1f8, 32'hc28daedb, 32'h408f80af, 32'hc2251987};
test_output[20248:20255] = '{32'h0, 32'h0, 32'h0, 32'h40dfc44f, 32'h0, 32'h0, 32'h408f80af, 32'h0};
test_input[20256:20263] = '{32'hc17804f4, 32'hc2224443, 32'hc281b12e, 32'hc238c906, 32'hc2308cb0, 32'hc19b205d, 32'h4194383a, 32'hc23390b1};
test_output[20256:20263] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4194383a, 32'h0};
test_input[20264:20271] = '{32'hc203f182, 32'h42613bf9, 32'hc2917341, 32'hc20e21e1, 32'h40ef9d0d, 32'hc27712b0, 32'hc2bc9a46, 32'h4251ad3e};
test_output[20264:20271] = '{32'h0, 32'h42613bf9, 32'h0, 32'h0, 32'h40ef9d0d, 32'h0, 32'h0, 32'h4251ad3e};
test_input[20272:20279] = '{32'hc2c690f4, 32'h42a926e9, 32'h427f3afb, 32'h42b23fad, 32'hc2bf933b, 32'h410d8742, 32'h41ae4a23, 32'h41ff9709};
test_output[20272:20279] = '{32'h0, 32'h42a926e9, 32'h427f3afb, 32'h42b23fad, 32'h0, 32'h410d8742, 32'h41ae4a23, 32'h41ff9709};
test_input[20280:20287] = '{32'h42c76faf, 32'h428ea0ab, 32'h4288cbf0, 32'hc0893403, 32'h42110ce3, 32'hc1ba2c2a, 32'hc24f5db1, 32'hc22ec071};
test_output[20280:20287] = '{32'h42c76faf, 32'h428ea0ab, 32'h4288cbf0, 32'h0, 32'h42110ce3, 32'h0, 32'h0, 32'h0};
test_input[20288:20295] = '{32'hc164b99b, 32'h410ad7bc, 32'h4295d106, 32'hc29443d9, 32'hc1b2832d, 32'hc1878396, 32'h41b18eee, 32'hbfaeae05};
test_output[20288:20295] = '{32'h0, 32'h410ad7bc, 32'h4295d106, 32'h0, 32'h0, 32'h0, 32'h41b18eee, 32'h0};
test_input[20296:20303] = '{32'hc28485e5, 32'h42c50341, 32'h4295125d, 32'h42bd8eef, 32'h4295a7d4, 32'hc27728e0, 32'h42816db9, 32'hc28af1d6};
test_output[20296:20303] = '{32'h0, 32'h42c50341, 32'h4295125d, 32'h42bd8eef, 32'h4295a7d4, 32'h0, 32'h42816db9, 32'h0};
test_input[20304:20311] = '{32'h41badd30, 32'hc1e7a859, 32'h42807357, 32'hc1511b46, 32'hc2a74177, 32'hc2816106, 32'hc16f014c, 32'hc184b69f};
test_output[20304:20311] = '{32'h41badd30, 32'h0, 32'h42807357, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20312:20319] = '{32'h40cd5f7e, 32'hc22cd084, 32'h41aafc95, 32'h429a0a92, 32'hc2a6ba39, 32'h4296a869, 32'h426a297e, 32'hc287cd5c};
test_output[20312:20319] = '{32'h40cd5f7e, 32'h0, 32'h41aafc95, 32'h429a0a92, 32'h0, 32'h4296a869, 32'h426a297e, 32'h0};
test_input[20320:20327] = '{32'hc2bc860b, 32'hc29a239d, 32'hc256d82d, 32'hc1d249e9, 32'hc28b88a6, 32'h40e2882d, 32'hc2c3ea70, 32'h41c2a770};
test_output[20320:20327] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40e2882d, 32'h0, 32'h41c2a770};
test_input[20328:20335] = '{32'hc1d85176, 32'h4264fb8d, 32'hc2672fe3, 32'hc2232a7f, 32'hbd8f1939, 32'h42a33783, 32'hc2c1cdc6, 32'h423809bb};
test_output[20328:20335] = '{32'h0, 32'h4264fb8d, 32'h0, 32'h0, 32'h0, 32'h42a33783, 32'h0, 32'h423809bb};
test_input[20336:20343] = '{32'h41c938c5, 32'hc18ddec6, 32'h404e6e25, 32'h40b92230, 32'h42abe784, 32'hc2c60226, 32'hc296312e, 32'h424c2d79};
test_output[20336:20343] = '{32'h41c938c5, 32'h0, 32'h404e6e25, 32'h40b92230, 32'h42abe784, 32'h0, 32'h0, 32'h424c2d79};
test_input[20344:20351] = '{32'h42510b92, 32'h416435c3, 32'h426b5c5d, 32'h429c53ed, 32'h42326c04, 32'hc26ca71d, 32'hc28887da, 32'hc2a8a0a3};
test_output[20344:20351] = '{32'h42510b92, 32'h416435c3, 32'h426b5c5d, 32'h429c53ed, 32'h42326c04, 32'h0, 32'h0, 32'h0};
test_input[20352:20359] = '{32'hc27619ca, 32'h415a6a83, 32'h422a3a29, 32'h42bb310b, 32'h41e5df74, 32'hc227f39e, 32'hc297a13e, 32'h425b6e79};
test_output[20352:20359] = '{32'h0, 32'h415a6a83, 32'h422a3a29, 32'h42bb310b, 32'h41e5df74, 32'h0, 32'h0, 32'h425b6e79};
test_input[20360:20367] = '{32'hc1d8da48, 32'hc2718637, 32'hc2c233a8, 32'hc22e884c, 32'h420c318d, 32'hc256bbf7, 32'hc033ceef, 32'h424b99dc};
test_output[20360:20367] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h420c318d, 32'h0, 32'h0, 32'h424b99dc};
test_input[20368:20375] = '{32'h41c71a86, 32'hc2875d93, 32'hc134e040, 32'hc277ad52, 32'hc2aaa82a, 32'h425588c5, 32'h41d2d856, 32'h422b88e8};
test_output[20368:20375] = '{32'h41c71a86, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425588c5, 32'h41d2d856, 32'h422b88e8};
test_input[20376:20383] = '{32'h41c2bd28, 32'hc299a397, 32'hc29babb0, 32'h42bad38e, 32'h41477fa8, 32'hc24389ec, 32'h428a58f1, 32'hc17003e1};
test_output[20376:20383] = '{32'h41c2bd28, 32'h0, 32'h0, 32'h42bad38e, 32'h41477fa8, 32'h0, 32'h428a58f1, 32'h0};
test_input[20384:20391] = '{32'h423e9a45, 32'h42bcca66, 32'h42bb1359, 32'h413780c6, 32'h41d6cd0c, 32'h421e8d63, 32'hc2ae95f7, 32'hc24d84cd};
test_output[20384:20391] = '{32'h423e9a45, 32'h42bcca66, 32'h42bb1359, 32'h413780c6, 32'h41d6cd0c, 32'h421e8d63, 32'h0, 32'h0};
test_input[20392:20399] = '{32'h4239fb9b, 32'hc2798946, 32'h41cc3b8e, 32'hc25779d2, 32'hc2931489, 32'h42b5eb49, 32'h421e8ab5, 32'hc20683cf};
test_output[20392:20399] = '{32'h4239fb9b, 32'h0, 32'h41cc3b8e, 32'h0, 32'h0, 32'h42b5eb49, 32'h421e8ab5, 32'h0};
test_input[20400:20407] = '{32'h4101f793, 32'hc1d5e5ff, 32'hc1476f72, 32'hc25af3aa, 32'hc286342b, 32'h42b31c3a, 32'hc01a0449, 32'hc2bb1ee8};
test_output[20400:20407] = '{32'h4101f793, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b31c3a, 32'h0, 32'h0};
test_input[20408:20415] = '{32'h42acbc96, 32'h4180ea07, 32'h42363733, 32'hc267e3fb, 32'h428c416f, 32'hc2b903a0, 32'hc15113d2, 32'hc25b7ad0};
test_output[20408:20415] = '{32'h42acbc96, 32'h4180ea07, 32'h42363733, 32'h0, 32'h428c416f, 32'h0, 32'h0, 32'h0};
test_input[20416:20423] = '{32'hc1f1100c, 32'hc2b62209, 32'hc23025d3, 32'h429d15e3, 32'h42a075f9, 32'hc2baa3c3, 32'hc28b287c, 32'hc239093e};
test_output[20416:20423] = '{32'h0, 32'h0, 32'h0, 32'h429d15e3, 32'h42a075f9, 32'h0, 32'h0, 32'h0};
test_input[20424:20431] = '{32'h42b79a5b, 32'hc1528b5d, 32'h4113c5fb, 32'hc2a47a75, 32'hc2765ce6, 32'hc2526aff, 32'h4288253a, 32'h429fb44c};
test_output[20424:20431] = '{32'h42b79a5b, 32'h0, 32'h4113c5fb, 32'h0, 32'h0, 32'h0, 32'h4288253a, 32'h429fb44c};
test_input[20432:20439] = '{32'hc2147f17, 32'hc19eccff, 32'h4282cb84, 32'h4290779e, 32'hc2446335, 32'hc25c3407, 32'h4208d369, 32'hc2c40fd3};
test_output[20432:20439] = '{32'h0, 32'h0, 32'h4282cb84, 32'h4290779e, 32'h0, 32'h0, 32'h4208d369, 32'h0};
test_input[20440:20447] = '{32'h3f27ce9e, 32'h423533b3, 32'hc2725385, 32'hc29f2f0a, 32'hc0dccb04, 32'hc2b2c8db, 32'h42904401, 32'h42929290};
test_output[20440:20447] = '{32'h3f27ce9e, 32'h423533b3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42904401, 32'h42929290};
test_input[20448:20455] = '{32'h40021d59, 32'hc20eb414, 32'hc1f6c548, 32'h428d0b6b, 32'hc2565285, 32'hc28f8fcd, 32'hc21b309e, 32'h4215abce};
test_output[20448:20455] = '{32'h40021d59, 32'h0, 32'h0, 32'h428d0b6b, 32'h0, 32'h0, 32'h0, 32'h4215abce};
test_input[20456:20463] = '{32'h422a949f, 32'hc294c931, 32'h424a8d47, 32'hc117a6a6, 32'hc2a8f8a9, 32'h3f877da8, 32'hc2919fbc, 32'h42c11d97};
test_output[20456:20463] = '{32'h422a949f, 32'h0, 32'h424a8d47, 32'h0, 32'h0, 32'h3f877da8, 32'h0, 32'h42c11d97};
test_input[20464:20471] = '{32'h420e7b12, 32'hc285735d, 32'h42368ad7, 32'hc13a6c46, 32'hc267fc5e, 32'hc29eeb64, 32'hc2a55797, 32'h428259f2};
test_output[20464:20471] = '{32'h420e7b12, 32'h0, 32'h42368ad7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428259f2};
test_input[20472:20479] = '{32'hc237609b, 32'hc220d46b, 32'h428f6125, 32'h416a66b1, 32'h42c0a074, 32'hc1f98921, 32'h41c2b65d, 32'h41d2663d};
test_output[20472:20479] = '{32'h0, 32'h0, 32'h428f6125, 32'h416a66b1, 32'h42c0a074, 32'h0, 32'h41c2b65d, 32'h41d2663d};
test_input[20480:20487] = '{32'hc1ff7987, 32'hc27fe3a4, 32'h427a42bf, 32'h422e6ce9, 32'hc1469764, 32'hc27fc636, 32'h4161e751, 32'hc14714c8};
test_output[20480:20487] = '{32'h0, 32'h0, 32'h427a42bf, 32'h422e6ce9, 32'h0, 32'h0, 32'h4161e751, 32'h0};
test_input[20488:20495] = '{32'h427cd458, 32'h41d60921, 32'hc264ea89, 32'h4114e078, 32'h42654605, 32'h42b43861, 32'h41af26d8, 32'h41ae2a2c};
test_output[20488:20495] = '{32'h427cd458, 32'h41d60921, 32'h0, 32'h4114e078, 32'h42654605, 32'h42b43861, 32'h41af26d8, 32'h41ae2a2c};
test_input[20496:20503] = '{32'hc1a0d641, 32'hc237c06c, 32'hc2bad6c0, 32'hc2c55140, 32'h41e36c1c, 32'hc1709d59, 32'hc2b9378c, 32'hc2be6dd1};
test_output[20496:20503] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41e36c1c, 32'h0, 32'h0, 32'h0};
test_input[20504:20511] = '{32'hc149f508, 32'h4232abaf, 32'h4289dbf5, 32'hc29cd7e0, 32'hc292fbff, 32'h412edcb8, 32'h40aab998, 32'hc2967300};
test_output[20504:20511] = '{32'h0, 32'h4232abaf, 32'h4289dbf5, 32'h0, 32'h0, 32'h412edcb8, 32'h40aab998, 32'h0};
test_input[20512:20519] = '{32'h41dc8d09, 32'hc2a8284d, 32'h42a2c269, 32'h42c20bd7, 32'h42a8d376, 32'h4195d1f6, 32'h41c143f9, 32'hc27177bf};
test_output[20512:20519] = '{32'h41dc8d09, 32'h0, 32'h42a2c269, 32'h42c20bd7, 32'h42a8d376, 32'h4195d1f6, 32'h41c143f9, 32'h0};
test_input[20520:20527] = '{32'h41ea4ca5, 32'hc0473a2c, 32'h4295e93d, 32'h40e8c50c, 32'h429898ca, 32'h4283b6b6, 32'hc1c2fc9b, 32'hc08fbd1b};
test_output[20520:20527] = '{32'h41ea4ca5, 32'h0, 32'h4295e93d, 32'h40e8c50c, 32'h429898ca, 32'h4283b6b6, 32'h0, 32'h0};
test_input[20528:20535] = '{32'hc2407e56, 32'h42c7fc3c, 32'hc2849acd, 32'hc2b56b69, 32'hc24bfe5a, 32'h424059ba, 32'hc283a2f9, 32'h42ac8cfb};
test_output[20528:20535] = '{32'h0, 32'h42c7fc3c, 32'h0, 32'h0, 32'h0, 32'h424059ba, 32'h0, 32'h42ac8cfb};
test_input[20536:20543] = '{32'h427db0a2, 32'h42832867, 32'hc0c86c65, 32'hc2014eb1, 32'hc2bad3ef, 32'hc25a76b6, 32'hc21f4bcc, 32'hc1f7ed07};
test_output[20536:20543] = '{32'h427db0a2, 32'h42832867, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20544:20551] = '{32'hc280ff64, 32'hc02366a7, 32'h426aa521, 32'h425895fc, 32'hc294d4f6, 32'hc10d99b8, 32'h41565fcd, 32'h42067d1e};
test_output[20544:20551] = '{32'h0, 32'h0, 32'h426aa521, 32'h425895fc, 32'h0, 32'h0, 32'h41565fcd, 32'h42067d1e};
test_input[20552:20559] = '{32'hc2161df3, 32'hc1feab45, 32'h41dcd994, 32'hc2b51442, 32'hc261bb5d, 32'hc29c7cec, 32'h42130879, 32'hc15c57ff};
test_output[20552:20559] = '{32'h0, 32'h0, 32'h41dcd994, 32'h0, 32'h0, 32'h0, 32'h42130879, 32'h0};
test_input[20560:20567] = '{32'h42782d04, 32'hc07ebfcd, 32'h3df7b5e5, 32'hc01358b7, 32'h4233d597, 32'h4205b273, 32'hc2a2e563, 32'h42c0b0c7};
test_output[20560:20567] = '{32'h42782d04, 32'h0, 32'h3df7b5e5, 32'h0, 32'h4233d597, 32'h4205b273, 32'h0, 32'h42c0b0c7};
test_input[20568:20575] = '{32'hc2522c9b, 32'h4245972c, 32'hc2a0e28f, 32'h423cee9d, 32'h41d2a175, 32'hc279be1e, 32'h42aa9931, 32'hc2996285};
test_output[20568:20575] = '{32'h0, 32'h4245972c, 32'h0, 32'h423cee9d, 32'h41d2a175, 32'h0, 32'h42aa9931, 32'h0};
test_input[20576:20583] = '{32'h42c78985, 32'h42a47142, 32'h427c52c2, 32'hc221a704, 32'h42281c84, 32'h428de414, 32'hc23521d9, 32'hc1014e67};
test_output[20576:20583] = '{32'h42c78985, 32'h42a47142, 32'h427c52c2, 32'h0, 32'h42281c84, 32'h428de414, 32'h0, 32'h0};
test_input[20584:20591] = '{32'hc1e8717c, 32'hc14a0aa1, 32'h427bc919, 32'h42b6f655, 32'h405506e7, 32'hc2966125, 32'h41d004a0, 32'hc2bd6b25};
test_output[20584:20591] = '{32'h0, 32'h0, 32'h427bc919, 32'h42b6f655, 32'h405506e7, 32'h0, 32'h41d004a0, 32'h0};
test_input[20592:20599] = '{32'hc1d60722, 32'h41bb324d, 32'hc2ab2f10, 32'hc28f6361, 32'hc240f47f, 32'hc29de79c, 32'h429bd239, 32'h42241156};
test_output[20592:20599] = '{32'h0, 32'h41bb324d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429bd239, 32'h42241156};
test_input[20600:20607] = '{32'h420a9a92, 32'h41cd2313, 32'hc166335a, 32'h4299d7c9, 32'h42768ad4, 32'hc21e7342, 32'hc20cc079, 32'hc087aea1};
test_output[20600:20607] = '{32'h420a9a92, 32'h41cd2313, 32'h0, 32'h4299d7c9, 32'h42768ad4, 32'h0, 32'h0, 32'h0};
test_input[20608:20615] = '{32'hc24c5ece, 32'hc2a5f094, 32'h422f3944, 32'hc1178454, 32'h42767e27, 32'hc2ae7029, 32'h426a8857, 32'hc290a02c};
test_output[20608:20615] = '{32'h0, 32'h0, 32'h422f3944, 32'h0, 32'h42767e27, 32'h0, 32'h426a8857, 32'h0};
test_input[20616:20623] = '{32'hc2a8fb61, 32'h419696ae, 32'hc1897fe9, 32'h4199593b, 32'h4228cbfa, 32'hc28b357b, 32'hc29b01c6, 32'hc24026c8};
test_output[20616:20623] = '{32'h0, 32'h419696ae, 32'h0, 32'h4199593b, 32'h4228cbfa, 32'h0, 32'h0, 32'h0};
test_input[20624:20631] = '{32'h42c130a7, 32'h40ac133b, 32'hc2a1de99, 32'h40f3e7a9, 32'hc25bf943, 32'hc1f9de40, 32'h41876e41, 32'hc2c33679};
test_output[20624:20631] = '{32'h42c130a7, 32'h40ac133b, 32'h0, 32'h40f3e7a9, 32'h0, 32'h0, 32'h41876e41, 32'h0};
test_input[20632:20639] = '{32'h419a120d, 32'hc2a16c66, 32'h4294a9cc, 32'h40758cc4, 32'hc057900f, 32'h419f8d42, 32'h41d9d90c, 32'hc24b9bef};
test_output[20632:20639] = '{32'h419a120d, 32'h0, 32'h4294a9cc, 32'h40758cc4, 32'h0, 32'h419f8d42, 32'h41d9d90c, 32'h0};
test_input[20640:20647] = '{32'hc2a8c51a, 32'h41546460, 32'hc219cf56, 32'hc22e1c92, 32'hc19241fa, 32'h42aeedb4, 32'h42b5a8c4, 32'hc285346d};
test_output[20640:20647] = '{32'h0, 32'h41546460, 32'h0, 32'h0, 32'h0, 32'h42aeedb4, 32'h42b5a8c4, 32'h0};
test_input[20648:20655] = '{32'h422eaffb, 32'hc2000db4, 32'h42770143, 32'h41e01c91, 32'h413bd29d, 32'hc10ddbba, 32'h41808962, 32'hc2c612ee};
test_output[20648:20655] = '{32'h422eaffb, 32'h0, 32'h42770143, 32'h41e01c91, 32'h413bd29d, 32'h0, 32'h41808962, 32'h0};
test_input[20656:20663] = '{32'h42b80375, 32'h4188d005, 32'hc2b1bd34, 32'hc28676c0, 32'h4297a76a, 32'h42a2c306, 32'h42588735, 32'hc261e0c3};
test_output[20656:20663] = '{32'h42b80375, 32'h4188d005, 32'h0, 32'h0, 32'h4297a76a, 32'h42a2c306, 32'h42588735, 32'h0};
test_input[20664:20671] = '{32'h418bdc70, 32'hc08c908d, 32'hc1dd67d6, 32'h41efd4df, 32'hc28660f7, 32'hc2b7d1aa, 32'h429bd00a, 32'hc1fd5eec};
test_output[20664:20671] = '{32'h418bdc70, 32'h0, 32'h0, 32'h41efd4df, 32'h0, 32'h0, 32'h429bd00a, 32'h0};
test_input[20672:20679] = '{32'h417a5b02, 32'h4205946a, 32'h42b2dc37, 32'hbfdbb228, 32'h42944847, 32'h422ab7e7, 32'hc0b0200b, 32'h42817ba7};
test_output[20672:20679] = '{32'h417a5b02, 32'h4205946a, 32'h42b2dc37, 32'h0, 32'h42944847, 32'h422ab7e7, 32'h0, 32'h42817ba7};
test_input[20680:20687] = '{32'hc29b0b35, 32'hc282f9d7, 32'hc2575474, 32'hc17e622c, 32'hc0ec1f01, 32'hc2c18ac4, 32'hc2ae61b5, 32'h411364db};
test_output[20680:20687] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h411364db};
test_input[20688:20695] = '{32'hc29f8a46, 32'h42ac5b92, 32'h422eb767, 32'h42a6e9b7, 32'hc294bb98, 32'hc2564164, 32'hc011e2ca, 32'h4291085a};
test_output[20688:20695] = '{32'h0, 32'h42ac5b92, 32'h422eb767, 32'h42a6e9b7, 32'h0, 32'h0, 32'h0, 32'h4291085a};
test_input[20696:20703] = '{32'h423588ce, 32'h42491018, 32'h4211562c, 32'h42863e45, 32'hc1d875b8, 32'hc2893f14, 32'hc145cc0d, 32'h4255f99f};
test_output[20696:20703] = '{32'h423588ce, 32'h42491018, 32'h4211562c, 32'h42863e45, 32'h0, 32'h0, 32'h0, 32'h4255f99f};
test_input[20704:20711] = '{32'h41ace73d, 32'hc1ccce0a, 32'hc151b161, 32'hc20aaf25, 32'h42a489df, 32'h417808b4, 32'hc22897b0, 32'h4266d31b};
test_output[20704:20711] = '{32'h41ace73d, 32'h0, 32'h0, 32'h0, 32'h42a489df, 32'h417808b4, 32'h0, 32'h4266d31b};
test_input[20712:20719] = '{32'hc29fb046, 32'h41843034, 32'hc231648b, 32'hc285fcee, 32'hc224f4c0, 32'hc1f244bc, 32'hbfbe733a, 32'hc18b3923};
test_output[20712:20719] = '{32'h0, 32'h41843034, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20720:20727] = '{32'h42779b14, 32'hc23420e3, 32'hc27b23fb, 32'h42506a8c, 32'h428e532d, 32'h4289590e, 32'hc2b6e000, 32'hc1bb5b19};
test_output[20720:20727] = '{32'h42779b14, 32'h0, 32'h0, 32'h42506a8c, 32'h428e532d, 32'h4289590e, 32'h0, 32'h0};
test_input[20728:20735] = '{32'hc2799067, 32'h429a0732, 32'hc0ef2a80, 32'hc0ca1473, 32'h42a1548f, 32'h4299c5ae, 32'h42ae78fb, 32'h41bc8057};
test_output[20728:20735] = '{32'h0, 32'h429a0732, 32'h0, 32'h0, 32'h42a1548f, 32'h4299c5ae, 32'h42ae78fb, 32'h41bc8057};
test_input[20736:20743] = '{32'hc1319cb3, 32'hc2a2c61c, 32'h42346f6e, 32'h42c79990, 32'h3d3b80cc, 32'h429bc2f5, 32'h428a2e4a, 32'hc2b4ae50};
test_output[20736:20743] = '{32'h0, 32'h0, 32'h42346f6e, 32'h42c79990, 32'h3d3b80cc, 32'h429bc2f5, 32'h428a2e4a, 32'h0};
test_input[20744:20751] = '{32'h4191eeef, 32'h42b3fe57, 32'hc23c2ea8, 32'hc12dd0eb, 32'h42b2ef92, 32'h4219e988, 32'h42377519, 32'h42a53a8b};
test_output[20744:20751] = '{32'h4191eeef, 32'h42b3fe57, 32'h0, 32'h0, 32'h42b2ef92, 32'h4219e988, 32'h42377519, 32'h42a53a8b};
test_input[20752:20759] = '{32'hc2b8031e, 32'h42bf29ab, 32'hc21ce6ba, 32'hc1d43642, 32'hc22a02e7, 32'h4213d832, 32'h4263d983, 32'hc1c83307};
test_output[20752:20759] = '{32'h0, 32'h42bf29ab, 32'h0, 32'h0, 32'h0, 32'h4213d832, 32'h4263d983, 32'h0};
test_input[20760:20767] = '{32'h423e54d3, 32'h4293f265, 32'hc16f19b1, 32'hc2a3c111, 32'h42b9290d, 32'hc16d0a24, 32'h4290556b, 32'h42834b7e};
test_output[20760:20767] = '{32'h423e54d3, 32'h4293f265, 32'h0, 32'h0, 32'h42b9290d, 32'h0, 32'h4290556b, 32'h42834b7e};
test_input[20768:20775] = '{32'h4199d611, 32'h41f71da6, 32'hc244b1f2, 32'h40645672, 32'hc2aef0be, 32'hc299f200, 32'h426ef807, 32'h41aef422};
test_output[20768:20775] = '{32'h4199d611, 32'h41f71da6, 32'h0, 32'h40645672, 32'h0, 32'h0, 32'h426ef807, 32'h41aef422};
test_input[20776:20783] = '{32'h42b9399a, 32'hc12099f9, 32'h42ad12fb, 32'h427191a1, 32'h4167c7a9, 32'h428ec517, 32'h42a83a19, 32'hc2a61b3e};
test_output[20776:20783] = '{32'h42b9399a, 32'h0, 32'h42ad12fb, 32'h427191a1, 32'h4167c7a9, 32'h428ec517, 32'h42a83a19, 32'h0};
test_input[20784:20791] = '{32'hbf9379fd, 32'hc1688042, 32'h42a58049, 32'h428887c2, 32'h40ceb2c3, 32'h42c28ed5, 32'hc1f6ebf6, 32'h409df683};
test_output[20784:20791] = '{32'h0, 32'h0, 32'h42a58049, 32'h428887c2, 32'h40ceb2c3, 32'h42c28ed5, 32'h0, 32'h409df683};
test_input[20792:20799] = '{32'hc2988d05, 32'hc2abb55c, 32'h414f8588, 32'hc2978b24, 32'h4198f912, 32'hc20ea0d1, 32'h422e0961, 32'hc1887d4e};
test_output[20792:20799] = '{32'h0, 32'h0, 32'h414f8588, 32'h0, 32'h4198f912, 32'h0, 32'h422e0961, 32'h0};
test_input[20800:20807] = '{32'h4259766b, 32'h418ff947, 32'hc1352fb7, 32'hc1d106a9, 32'h427ae396, 32'hc2c69318, 32'h4036eb22, 32'h4181dc70};
test_output[20800:20807] = '{32'h4259766b, 32'h418ff947, 32'h0, 32'h0, 32'h427ae396, 32'h0, 32'h4036eb22, 32'h4181dc70};
test_input[20808:20815] = '{32'hc291bff2, 32'hc1de4a3d, 32'h42093c4b, 32'hc2b3d5b3, 32'hc28f5cb0, 32'h422fbe7f, 32'h41598b5d, 32'hc2912e7c};
test_output[20808:20815] = '{32'h0, 32'h0, 32'h42093c4b, 32'h0, 32'h0, 32'h422fbe7f, 32'h41598b5d, 32'h0};
test_input[20816:20823] = '{32'hc2928845, 32'h42acd55f, 32'h3ff31d26, 32'hc23305d5, 32'h428cd3f2, 32'hc2ae3267, 32'hc19a7594, 32'hc2192cc7};
test_output[20816:20823] = '{32'h0, 32'h42acd55f, 32'h3ff31d26, 32'h0, 32'h428cd3f2, 32'h0, 32'h0, 32'h0};
test_input[20824:20831] = '{32'h421a83a8, 32'h40ea2fc7, 32'h41cab5e2, 32'h42abce9f, 32'h41f85918, 32'h42bd3865, 32'hc1d3888a, 32'h3f3b8411};
test_output[20824:20831] = '{32'h421a83a8, 32'h40ea2fc7, 32'h41cab5e2, 32'h42abce9f, 32'h41f85918, 32'h42bd3865, 32'h0, 32'h3f3b8411};
test_input[20832:20839] = '{32'hc2c58af6, 32'hc2baadb6, 32'hc1b4ee76, 32'h42443271, 32'hc2a92ec8, 32'hc27aeb53, 32'hc29c362b, 32'hc25e24e2};
test_output[20832:20839] = '{32'h0, 32'h0, 32'h0, 32'h42443271, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20840:20847] = '{32'hc2ad6f69, 32'hc2a8bc78, 32'h42a216f7, 32'hc1b433d9, 32'h426853bf, 32'hc24f0643, 32'h42662c5e, 32'hc297d72b};
test_output[20840:20847] = '{32'h0, 32'h0, 32'h42a216f7, 32'h0, 32'h426853bf, 32'h0, 32'h42662c5e, 32'h0};
test_input[20848:20855] = '{32'hc233c428, 32'h42024bba, 32'hc2c7d7a8, 32'hc1cd65a3, 32'h4192e8af, 32'h42617bcf, 32'hc1c7609b, 32'h41c8fb1b};
test_output[20848:20855] = '{32'h0, 32'h42024bba, 32'h0, 32'h0, 32'h4192e8af, 32'h42617bcf, 32'h0, 32'h41c8fb1b};
test_input[20856:20863] = '{32'h425bec4a, 32'hc0fef3b6, 32'hc292646a, 32'h420f6553, 32'hc1ee6b03, 32'hc282355c, 32'hc0d54c64, 32'h429da1b1};
test_output[20856:20863] = '{32'h425bec4a, 32'h0, 32'h0, 32'h420f6553, 32'h0, 32'h0, 32'h0, 32'h429da1b1};
test_input[20864:20871] = '{32'hc21e9eec, 32'hc289970e, 32'h42c14db9, 32'hc1ad73cb, 32'h417420ee, 32'h42b4fa96, 32'h42545bb8, 32'hc2bc2129};
test_output[20864:20871] = '{32'h0, 32'h0, 32'h42c14db9, 32'h0, 32'h417420ee, 32'h42b4fa96, 32'h42545bb8, 32'h0};
test_input[20872:20879] = '{32'h420ddec6, 32'h4163d8fc, 32'h40b2b1bf, 32'hc26406e8, 32'hc23365db, 32'h426751a2, 32'h4236f661, 32'h42854c26};
test_output[20872:20879] = '{32'h420ddec6, 32'h4163d8fc, 32'h40b2b1bf, 32'h0, 32'h0, 32'h426751a2, 32'h4236f661, 32'h42854c26};
test_input[20880:20887] = '{32'h42653fb3, 32'hc2ad5c39, 32'hc200358f, 32'h423c8392, 32'h40db2581, 32'h4112344d, 32'h40a2ec11, 32'hc219f2c9};
test_output[20880:20887] = '{32'h42653fb3, 32'h0, 32'h0, 32'h423c8392, 32'h40db2581, 32'h4112344d, 32'h40a2ec11, 32'h0};
test_input[20888:20895] = '{32'hc2ae6fb1, 32'h42323765, 32'hc1e09c1a, 32'hc1fac57b, 32'hc1967eec, 32'hc238bf77, 32'h42ad1437, 32'h41fde198};
test_output[20888:20895] = '{32'h0, 32'h42323765, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ad1437, 32'h41fde198};
test_input[20896:20903] = '{32'hc137886a, 32'h4171d93d, 32'hc252ade2, 32'hc04f711c, 32'h429d466e, 32'hc233556c, 32'h42b77296, 32'h4261ba90};
test_output[20896:20903] = '{32'h0, 32'h4171d93d, 32'h0, 32'h0, 32'h429d466e, 32'h0, 32'h42b77296, 32'h4261ba90};
test_input[20904:20911] = '{32'hc1596d58, 32'h425bf623, 32'h415171ba, 32'hc26e2a02, 32'hc01d6dac, 32'h40920904, 32'h42a51968, 32'h4256af8f};
test_output[20904:20911] = '{32'h0, 32'h425bf623, 32'h415171ba, 32'h0, 32'h0, 32'h40920904, 32'h42a51968, 32'h4256af8f};
test_input[20912:20919] = '{32'h421b393b, 32'hc290b0b1, 32'hc251f5f1, 32'hc28d2ef8, 32'hc1cf30fe, 32'hc1d0b25a, 32'hc288dd54, 32'hc161ccf6};
test_output[20912:20919] = '{32'h421b393b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20920:20927] = '{32'hc2003503, 32'h42babaec, 32'hbf751d93, 32'hc1ce8769, 32'hc294f597, 32'h4202a702, 32'h41964293, 32'h420a1622};
test_output[20920:20927] = '{32'h0, 32'h42babaec, 32'h0, 32'h0, 32'h0, 32'h4202a702, 32'h41964293, 32'h420a1622};
test_input[20928:20935] = '{32'hc272a023, 32'hc2199447, 32'hc12e4921, 32'hbfaa4424, 32'h42134945, 32'h42aa34c3, 32'hc201e928, 32'h41e00284};
test_output[20928:20935] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42134945, 32'h42aa34c3, 32'h0, 32'h41e00284};
test_input[20936:20943] = '{32'hc2444547, 32'hc2b5f642, 32'h414f3ccf, 32'h40eeed8b, 32'h420539b6, 32'h424eefbe, 32'h42723fa5, 32'h42b420e2};
test_output[20936:20943] = '{32'h0, 32'h0, 32'h414f3ccf, 32'h40eeed8b, 32'h420539b6, 32'h424eefbe, 32'h42723fa5, 32'h42b420e2};
test_input[20944:20951] = '{32'hc1dad543, 32'hc18bb0c4, 32'h42b51dfb, 32'hc18717f5, 32'hc2ab7d01, 32'h4245b75e, 32'hc2c7d93d, 32'h4136461d};
test_output[20944:20951] = '{32'h0, 32'h0, 32'h42b51dfb, 32'h0, 32'h0, 32'h4245b75e, 32'h0, 32'h4136461d};
test_input[20952:20959] = '{32'h415e1cdb, 32'hc28e0c5f, 32'hc226e5de, 32'h429b3470, 32'h429cb1eb, 32'h4213163b, 32'h41bde692, 32'hc2c1425b};
test_output[20952:20959] = '{32'h415e1cdb, 32'h0, 32'h0, 32'h429b3470, 32'h429cb1eb, 32'h4213163b, 32'h41bde692, 32'h0};
test_input[20960:20967] = '{32'h418011b1, 32'h418006c9, 32'hc1e3f6ee, 32'h42b497d5, 32'hc2c51fd9, 32'hc2a5c169, 32'hc2b70a71, 32'h426400ab};
test_output[20960:20967] = '{32'h418011b1, 32'h418006c9, 32'h0, 32'h42b497d5, 32'h0, 32'h0, 32'h0, 32'h426400ab};
test_input[20968:20975] = '{32'h40fba5c7, 32'hc1a4f1e8, 32'h4230552d, 32'hc112c6b7, 32'h42a94382, 32'hc218b609, 32'h421e1d66, 32'h4282f9e0};
test_output[20968:20975] = '{32'h40fba5c7, 32'h0, 32'h4230552d, 32'h0, 32'h42a94382, 32'h0, 32'h421e1d66, 32'h4282f9e0};
test_input[20976:20983] = '{32'h42754f26, 32'h422bd5fb, 32'h42362604, 32'hc1d521c1, 32'hc22fbf6b, 32'h42aac05e, 32'hc0cc34f7, 32'h41f89340};
test_output[20976:20983] = '{32'h42754f26, 32'h422bd5fb, 32'h42362604, 32'h0, 32'h0, 32'h42aac05e, 32'h0, 32'h41f89340};
test_input[20984:20991] = '{32'h41443f5f, 32'hc2bb7a45, 32'hc26f5a10, 32'hc2ac9995, 32'h418ff05c, 32'hc2bae8f9, 32'h4259d135, 32'hbf69effa};
test_output[20984:20991] = '{32'h41443f5f, 32'h0, 32'h0, 32'h0, 32'h418ff05c, 32'h0, 32'h4259d135, 32'h0};
test_input[20992:20999] = '{32'h4134f409, 32'hc2a45546, 32'h427d601d, 32'hc26213e1, 32'h429e4706, 32'hc2ba7343, 32'h423c84f1, 32'hc1000e72};
test_output[20992:20999] = '{32'h4134f409, 32'h0, 32'h427d601d, 32'h0, 32'h429e4706, 32'h0, 32'h423c84f1, 32'h0};
test_input[21000:21007] = '{32'h429014e9, 32'hc1b74644, 32'hc2166327, 32'h3e60c93e, 32'hc2c5fa2c, 32'h41e17c21, 32'hc283dcc9, 32'hc2b88598};
test_output[21000:21007] = '{32'h429014e9, 32'h0, 32'h0, 32'h3e60c93e, 32'h0, 32'h41e17c21, 32'h0, 32'h0};
test_input[21008:21015] = '{32'hc261c93d, 32'hc10c9e67, 32'h429dbbbe, 32'hc29704b2, 32'h429b7e26, 32'hc1f09d6a, 32'hc1efa433, 32'h42c4d674};
test_output[21008:21015] = '{32'h0, 32'h0, 32'h429dbbbe, 32'h0, 32'h429b7e26, 32'h0, 32'h0, 32'h42c4d674};
test_input[21016:21023] = '{32'hc295301a, 32'h41bfa7a8, 32'h4198efa1, 32'hc2c54e74, 32'hc2619c6f, 32'h423f5770, 32'hc1ddc451, 32'hc0d6c293};
test_output[21016:21023] = '{32'h0, 32'h41bfa7a8, 32'h4198efa1, 32'h0, 32'h0, 32'h423f5770, 32'h0, 32'h0};
test_input[21024:21031] = '{32'h42a73b47, 32'hc264bfe4, 32'hc1c59470, 32'hc286418c, 32'h41cfa43a, 32'hc20f047b, 32'h402c7452, 32'hc114cb54};
test_output[21024:21031] = '{32'h42a73b47, 32'h0, 32'h0, 32'h0, 32'h41cfa43a, 32'h0, 32'h402c7452, 32'h0};
test_input[21032:21039] = '{32'h42aeba08, 32'hc2642377, 32'hc209fcf8, 32'h426ba752, 32'h414520f9, 32'hc294264a, 32'h428d00df, 32'h42a4ed68};
test_output[21032:21039] = '{32'h42aeba08, 32'h0, 32'h0, 32'h426ba752, 32'h414520f9, 32'h0, 32'h428d00df, 32'h42a4ed68};
test_input[21040:21047] = '{32'hc29ed864, 32'hc298cf1e, 32'h424794e2, 32'h42b06a55, 32'hc2b127cc, 32'h42871938, 32'h42badaab, 32'h42a4cc62};
test_output[21040:21047] = '{32'h0, 32'h0, 32'h424794e2, 32'h42b06a55, 32'h0, 32'h42871938, 32'h42badaab, 32'h42a4cc62};
test_input[21048:21055] = '{32'h41b65de6, 32'h42779c36, 32'h42869696, 32'hc26aba65, 32'hc2a7fd76, 32'h420f47e0, 32'h42178aa4, 32'h408b9458};
test_output[21048:21055] = '{32'h41b65de6, 32'h42779c36, 32'h42869696, 32'h0, 32'h0, 32'h420f47e0, 32'h42178aa4, 32'h408b9458};
test_input[21056:21063] = '{32'h427bcbcf, 32'h424aab61, 32'h3fb8ecc1, 32'h4201c3db, 32'hc23796a6, 32'hc1493890, 32'h42bb3a00, 32'h42a93152};
test_output[21056:21063] = '{32'h427bcbcf, 32'h424aab61, 32'h3fb8ecc1, 32'h4201c3db, 32'h0, 32'h0, 32'h42bb3a00, 32'h42a93152};
test_input[21064:21071] = '{32'h429d5a09, 32'h40b33c19, 32'hc1fbd084, 32'h40fde8d9, 32'hc1045cbf, 32'h428f3af3, 32'h42b5eb9b, 32'h40f03a10};
test_output[21064:21071] = '{32'h429d5a09, 32'h40b33c19, 32'h0, 32'h40fde8d9, 32'h0, 32'h428f3af3, 32'h42b5eb9b, 32'h40f03a10};
test_input[21072:21079] = '{32'hc1e23ab8, 32'hc2b5f6f4, 32'hc18b6a42, 32'hc2a824f9, 32'h4125d0c4, 32'h42b368f8, 32'h42be6d56, 32'h4217d51c};
test_output[21072:21079] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4125d0c4, 32'h42b368f8, 32'h42be6d56, 32'h4217d51c};
test_input[21080:21087] = '{32'h42bf59ca, 32'h41df22cb, 32'h42aece48, 32'hc262ce45, 32'h41a59d2f, 32'hc2a776e0, 32'hc1c8d554, 32'hc2887de2};
test_output[21080:21087] = '{32'h42bf59ca, 32'h41df22cb, 32'h42aece48, 32'h0, 32'h41a59d2f, 32'h0, 32'h0, 32'h0};
test_input[21088:21095] = '{32'hbff2fba4, 32'hc2b5106c, 32'h42ba7ab6, 32'h426499f6, 32'h4292f7d2, 32'h42c79a1e, 32'hc28d4456, 32'hc2864115};
test_output[21088:21095] = '{32'h0, 32'h0, 32'h42ba7ab6, 32'h426499f6, 32'h4292f7d2, 32'h42c79a1e, 32'h0, 32'h0};
test_input[21096:21103] = '{32'h4297481e, 32'h42b9a883, 32'h4117ec13, 32'hc21a547b, 32'h412fafe3, 32'h4267805d, 32'hc187a9c7, 32'hc26eb8ed};
test_output[21096:21103] = '{32'h4297481e, 32'h42b9a883, 32'h4117ec13, 32'h0, 32'h412fafe3, 32'h4267805d, 32'h0, 32'h0};
test_input[21104:21111] = '{32'h427c1a6e, 32'hc21a1d79, 32'hc2b562e8, 32'hc2b8b689, 32'h407ebc51, 32'hc1d5c23b, 32'hc2bda643, 32'h42104708};
test_output[21104:21111] = '{32'h427c1a6e, 32'h0, 32'h0, 32'h0, 32'h407ebc51, 32'h0, 32'h0, 32'h42104708};
test_input[21112:21119] = '{32'h428362be, 32'hc24c9d48, 32'hc28c8d5f, 32'hc22701ce, 32'hc29f6b8a, 32'h4239a564, 32'h42b71326, 32'h42854d10};
test_output[21112:21119] = '{32'h428362be, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4239a564, 32'h42b71326, 32'h42854d10};
test_input[21120:21127] = '{32'hc1807f77, 32'hc1f90626, 32'hc293f88b, 32'h41b1bda8, 32'h41bd7928, 32'hc2504640, 32'h422f607a, 32'hbe93723f};
test_output[21120:21127] = '{32'h0, 32'h0, 32'h0, 32'h41b1bda8, 32'h41bd7928, 32'h0, 32'h422f607a, 32'h0};
test_input[21128:21135] = '{32'hc21bf5a2, 32'h4144b41d, 32'h40f60d68, 32'h4265c68c, 32'h41e5b2a2, 32'h41ee90b8, 32'hc2c56468, 32'hc1c352df};
test_output[21128:21135] = '{32'h0, 32'h4144b41d, 32'h40f60d68, 32'h4265c68c, 32'h41e5b2a2, 32'h41ee90b8, 32'h0, 32'h0};
test_input[21136:21143] = '{32'hc01ae0d6, 32'h42bc02d0, 32'h429d197d, 32'h429ca118, 32'h42adf18d, 32'h419b30fb, 32'hc19d1d6c, 32'h421fa7a6};
test_output[21136:21143] = '{32'h0, 32'h42bc02d0, 32'h429d197d, 32'h429ca118, 32'h42adf18d, 32'h419b30fb, 32'h0, 32'h421fa7a6};
test_input[21144:21151] = '{32'h40e4b2d3, 32'hc290029f, 32'h417cc04d, 32'h42b36347, 32'h41900909, 32'h428bfab3, 32'hc0b1643e, 32'h426ee517};
test_output[21144:21151] = '{32'h40e4b2d3, 32'h0, 32'h417cc04d, 32'h42b36347, 32'h41900909, 32'h428bfab3, 32'h0, 32'h426ee517};
test_input[21152:21159] = '{32'hc2802bb4, 32'h41c34b39, 32'hc2accf11, 32'h420dc502, 32'h41e973d1, 32'hc230b223, 32'hc27100f6, 32'hc1e802f3};
test_output[21152:21159] = '{32'h0, 32'h41c34b39, 32'h0, 32'h420dc502, 32'h41e973d1, 32'h0, 32'h0, 32'h0};
test_input[21160:21167] = '{32'h40a56b93, 32'h40192afc, 32'h42c70a21, 32'h424b687c, 32'h426581d1, 32'h423f8354, 32'h4200422a, 32'hc25e74cd};
test_output[21160:21167] = '{32'h40a56b93, 32'h40192afc, 32'h42c70a21, 32'h424b687c, 32'h426581d1, 32'h423f8354, 32'h4200422a, 32'h0};
test_input[21168:21175] = '{32'h41029064, 32'h3ee55151, 32'h423bd5f5, 32'h4299db62, 32'h428764c3, 32'hc2805630, 32'h41d7b3ee, 32'h4204f486};
test_output[21168:21175] = '{32'h41029064, 32'h3ee55151, 32'h423bd5f5, 32'h4299db62, 32'h428764c3, 32'h0, 32'h41d7b3ee, 32'h4204f486};
test_input[21176:21183] = '{32'hc209aa33, 32'hc2c56518, 32'hc25d2fc1, 32'hc2a3aced, 32'h4153dd3b, 32'h42a70ddf, 32'h42254583, 32'h42bfb434};
test_output[21176:21183] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4153dd3b, 32'h42a70ddf, 32'h42254583, 32'h42bfb434};
test_input[21184:21191] = '{32'hc29df507, 32'h42ac2125, 32'hc23520be, 32'hc2c78340, 32'hc2c4d509, 32'hbe43f81f, 32'h4295ebb2, 32'h42a66342};
test_output[21184:21191] = '{32'h0, 32'h42ac2125, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4295ebb2, 32'h42a66342};
test_input[21192:21199] = '{32'hc254d881, 32'h41dfc46d, 32'hc2b24c72, 32'hc2c42a8d, 32'hbf4f06c8, 32'hc235dbcf, 32'hc262cdb1, 32'hc0a1659b};
test_output[21192:21199] = '{32'h0, 32'h41dfc46d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21200:21207] = '{32'hc1d18db4, 32'h42b07bc5, 32'hc2a8d02a, 32'hc2b596cc, 32'h423d1fb4, 32'h4289f13d, 32'h4290736a, 32'h42b1f074};
test_output[21200:21207] = '{32'h0, 32'h42b07bc5, 32'h0, 32'h0, 32'h423d1fb4, 32'h4289f13d, 32'h4290736a, 32'h42b1f074};
test_input[21208:21215] = '{32'h402b3b78, 32'h41bfab3f, 32'hc2a078e2, 32'h427d98a6, 32'hc2350dd2, 32'hc14c866b, 32'hc0e3b8e8, 32'hc2306506};
test_output[21208:21215] = '{32'h402b3b78, 32'h41bfab3f, 32'h0, 32'h427d98a6, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21216:21223] = '{32'hc294141c, 32'h42881fb0, 32'h42748fcb, 32'hc2065b06, 32'hc14c31da, 32'hc296d7df, 32'h41860108, 32'h42b0dc87};
test_output[21216:21223] = '{32'h0, 32'h42881fb0, 32'h42748fcb, 32'h0, 32'h0, 32'h0, 32'h41860108, 32'h42b0dc87};
test_input[21224:21231] = '{32'hc2b09d61, 32'h3fdeb203, 32'h42163fca, 32'hc18cb0e4, 32'hc1eb875c, 32'hbfc25763, 32'hc08fbc59, 32'hc24e1a52};
test_output[21224:21231] = '{32'h0, 32'h3fdeb203, 32'h42163fca, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21232:21239] = '{32'hc2a50dee, 32'h426f364d, 32'h42c02165, 32'hc138611c, 32'h42bafaf3, 32'h425b5a93, 32'h419b0135, 32'hc2a7527b};
test_output[21232:21239] = '{32'h0, 32'h426f364d, 32'h42c02165, 32'h0, 32'h42bafaf3, 32'h425b5a93, 32'h419b0135, 32'h0};
test_input[21240:21247] = '{32'h42578bbc, 32'hc288cf44, 32'h4104bbfe, 32'hc187aecb, 32'h40bf3b03, 32'h42bd316f, 32'hc21c763b, 32'h42130fb6};
test_output[21240:21247] = '{32'h42578bbc, 32'h0, 32'h4104bbfe, 32'h0, 32'h40bf3b03, 32'h42bd316f, 32'h0, 32'h42130fb6};
test_input[21248:21255] = '{32'hc2799957, 32'hc12d9039, 32'h41eea18f, 32'h421eba7b, 32'hc29ca4a8, 32'hc03ca55a, 32'hc2980acd, 32'h428bdd32};
test_output[21248:21255] = '{32'h0, 32'h0, 32'h41eea18f, 32'h421eba7b, 32'h0, 32'h0, 32'h0, 32'h428bdd32};
test_input[21256:21263] = '{32'h42a82f59, 32'h40de18f4, 32'h426f217e, 32'h428716cd, 32'hc25226d3, 32'hc2b28b01, 32'h420cd404, 32'hc20a5164};
test_output[21256:21263] = '{32'h42a82f59, 32'h40de18f4, 32'h426f217e, 32'h428716cd, 32'h0, 32'h0, 32'h420cd404, 32'h0};
test_input[21264:21271] = '{32'h4275af32, 32'hc28b3d64, 32'h42102682, 32'hc1d2ac82, 32'hc2a219f2, 32'hc2aed2f5, 32'hc1dc132b, 32'hc223ff42};
test_output[21264:21271] = '{32'h4275af32, 32'h0, 32'h42102682, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21272:21279] = '{32'h41dffb00, 32'hc29312d1, 32'h41b0c193, 32'hc2a863f7, 32'hc24be5dc, 32'hc2bb258a, 32'h428c381b, 32'hc282e3f1};
test_output[21272:21279] = '{32'h41dffb00, 32'h0, 32'h41b0c193, 32'h0, 32'h0, 32'h0, 32'h428c381b, 32'h0};
test_input[21280:21287] = '{32'h42b3b690, 32'hc23d943c, 32'h40bce463, 32'h42c532e5, 32'hc2556f64, 32'h423242a5, 32'h41c7ce79, 32'hc29ffb46};
test_output[21280:21287] = '{32'h42b3b690, 32'h0, 32'h40bce463, 32'h42c532e5, 32'h0, 32'h423242a5, 32'h41c7ce79, 32'h0};
test_input[21288:21295] = '{32'h41a94dc1, 32'h41cae0c0, 32'h4142fc8d, 32'hc20b6925, 32'hc19fd23a, 32'hc1f0c5ea, 32'h4152463a, 32'h42a224b6};
test_output[21288:21295] = '{32'h41a94dc1, 32'h41cae0c0, 32'h4142fc8d, 32'h0, 32'h0, 32'h0, 32'h4152463a, 32'h42a224b6};
test_input[21296:21303] = '{32'hc2472ccd, 32'hc294d91e, 32'h42b7bce8, 32'hc1e230a0, 32'hc0f09598, 32'hc288d8a3, 32'hc278ab73, 32'hc249de7e};
test_output[21296:21303] = '{32'h0, 32'h0, 32'h42b7bce8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21304:21311] = '{32'hc14a0bd0, 32'h42190e43, 32'h4224da5e, 32'hc299cfaa, 32'h4219bcde, 32'h4111d631, 32'hc22f5c88, 32'hc27d4616};
test_output[21304:21311] = '{32'h0, 32'h42190e43, 32'h4224da5e, 32'h0, 32'h4219bcde, 32'h4111d631, 32'h0, 32'h0};
test_input[21312:21319] = '{32'hc290af3e, 32'h42a8a2d3, 32'hc2a5571c, 32'hc25db5c6, 32'hc28b4bcd, 32'h4249937c, 32'hc241d078, 32'h429e07d9};
test_output[21312:21319] = '{32'h0, 32'h42a8a2d3, 32'h0, 32'h0, 32'h0, 32'h4249937c, 32'h0, 32'h429e07d9};
test_input[21320:21327] = '{32'h41e04f74, 32'h421320ee, 32'hc276be25, 32'hc29a1376, 32'hbe13cfd1, 32'hc2abdee1, 32'hc1b1ca4c, 32'hc17b48c1};
test_output[21320:21327] = '{32'h41e04f74, 32'h421320ee, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21328:21335] = '{32'h41aa245a, 32'h428d2d86, 32'hc2a32183, 32'h41f6a25e, 32'h420bdd24, 32'hc23b34a3, 32'h4285b9ed, 32'h42123755};
test_output[21328:21335] = '{32'h41aa245a, 32'h428d2d86, 32'h0, 32'h41f6a25e, 32'h420bdd24, 32'h0, 32'h4285b9ed, 32'h42123755};
test_input[21336:21343] = '{32'hc24b13a0, 32'h4232fd1d, 32'hc28e920a, 32'h420629a0, 32'hc20a1068, 32'hc2141744, 32'h414cbec3, 32'h4218dc47};
test_output[21336:21343] = '{32'h0, 32'h4232fd1d, 32'h0, 32'h420629a0, 32'h0, 32'h0, 32'h414cbec3, 32'h4218dc47};
test_input[21344:21351] = '{32'hc2887e89, 32'hc2270c58, 32'h41ebb1c4, 32'hc2b7a788, 32'hbfec88a6, 32'h3fbda207, 32'h428f40a1, 32'hc2c3c631};
test_output[21344:21351] = '{32'h0, 32'h0, 32'h41ebb1c4, 32'h0, 32'h0, 32'h3fbda207, 32'h428f40a1, 32'h0};
test_input[21352:21359] = '{32'hc255943d, 32'h420f17f1, 32'h42b1a2d6, 32'h42b8bad2, 32'h428dd4fa, 32'hc133d1f7, 32'h4130d3e0, 32'hc28e3074};
test_output[21352:21359] = '{32'h0, 32'h420f17f1, 32'h42b1a2d6, 32'h42b8bad2, 32'h428dd4fa, 32'h0, 32'h4130d3e0, 32'h0};
test_input[21360:21367] = '{32'hc211b227, 32'h41ae8f2b, 32'h42bd7018, 32'hc24e83e4, 32'hc299aea8, 32'h4076bcc0, 32'h404b2aa1, 32'hc2930ffb};
test_output[21360:21367] = '{32'h0, 32'h41ae8f2b, 32'h42bd7018, 32'h0, 32'h0, 32'h4076bcc0, 32'h404b2aa1, 32'h0};
test_input[21368:21375] = '{32'h41bfc383, 32'h419c9e94, 32'h42b7176b, 32'hc218ead7, 32'hc21f6887, 32'hc23caa16, 32'hc2b0f0d1, 32'hc0af3dbd};
test_output[21368:21375] = '{32'h41bfc383, 32'h419c9e94, 32'h42b7176b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21376:21383] = '{32'hc2a60579, 32'hc277c9c2, 32'h429e0247, 32'hc1d0c233, 32'h41ced5d3, 32'h429b894d, 32'hc2a6b3fc, 32'hc217f8c0};
test_output[21376:21383] = '{32'h0, 32'h0, 32'h429e0247, 32'h0, 32'h41ced5d3, 32'h429b894d, 32'h0, 32'h0};
test_input[21384:21391] = '{32'h4245441f, 32'hc1d069ae, 32'h414f1c46, 32'hc28b6d81, 32'h4269d5a9, 32'h427ea0b8, 32'h4286df51, 32'hc2a9e149};
test_output[21384:21391] = '{32'h4245441f, 32'h0, 32'h414f1c46, 32'h0, 32'h4269d5a9, 32'h427ea0b8, 32'h4286df51, 32'h0};
test_input[21392:21399] = '{32'hc1f6e3da, 32'h4249022d, 32'hc287d213, 32'hc292c7df, 32'h423f95f0, 32'h42083c00, 32'h42749c21, 32'hc2965d9d};
test_output[21392:21399] = '{32'h0, 32'h4249022d, 32'h0, 32'h0, 32'h423f95f0, 32'h42083c00, 32'h42749c21, 32'h0};
test_input[21400:21407] = '{32'h42b818e8, 32'h41c94c14, 32'h4249696d, 32'h41c8b7d7, 32'hc04ec4ef, 32'hc112e642, 32'h4217dd76, 32'h41e4f23f};
test_output[21400:21407] = '{32'h42b818e8, 32'h41c94c14, 32'h4249696d, 32'h41c8b7d7, 32'h0, 32'h0, 32'h4217dd76, 32'h41e4f23f};
test_input[21408:21415] = '{32'h419a97fd, 32'hc1e9962b, 32'hc2be35d5, 32'h414f4ce3, 32'h42882ba2, 32'hc1a33b55, 32'hc03d2050, 32'h4289a54f};
test_output[21408:21415] = '{32'h419a97fd, 32'h0, 32'h0, 32'h414f4ce3, 32'h42882ba2, 32'h0, 32'h0, 32'h4289a54f};
test_input[21416:21423] = '{32'hc221fa3b, 32'h42964a68, 32'h40d95a82, 32'h42718df2, 32'h428d8531, 32'h42c40339, 32'h4208446b, 32'hc2146c19};
test_output[21416:21423] = '{32'h0, 32'h42964a68, 32'h40d95a82, 32'h42718df2, 32'h428d8531, 32'h42c40339, 32'h4208446b, 32'h0};
test_input[21424:21431] = '{32'hc250bf6d, 32'h4290c90d, 32'h42b2d21e, 32'h4131db0c, 32'h423c4c59, 32'hc2a31c8f, 32'h429bd050, 32'h429bb0af};
test_output[21424:21431] = '{32'h0, 32'h4290c90d, 32'h42b2d21e, 32'h4131db0c, 32'h423c4c59, 32'h0, 32'h429bd050, 32'h429bb0af};
test_input[21432:21439] = '{32'h412ab8ee, 32'h42207a2e, 32'hc242197e, 32'h4274f64a, 32'h421c5834, 32'h42585bb2, 32'hc21b08a7, 32'hc2af6781};
test_output[21432:21439] = '{32'h412ab8ee, 32'h42207a2e, 32'h0, 32'h4274f64a, 32'h421c5834, 32'h42585bb2, 32'h0, 32'h0};
test_input[21440:21447] = '{32'h42a8190a, 32'h42bdc00d, 32'hc2a20286, 32'hc0cbf866, 32'h41b65587, 32'h4263fb34, 32'h4243a159, 32'h40dd5190};
test_output[21440:21447] = '{32'h42a8190a, 32'h42bdc00d, 32'h0, 32'h0, 32'h41b65587, 32'h4263fb34, 32'h4243a159, 32'h40dd5190};
test_input[21448:21455] = '{32'hc262d3c0, 32'hc293f82b, 32'h42c438f2, 32'h42b62178, 32'hc11096d0, 32'hc27fb82c, 32'h4231f008, 32'h425d244f};
test_output[21448:21455] = '{32'h0, 32'h0, 32'h42c438f2, 32'h42b62178, 32'h0, 32'h0, 32'h4231f008, 32'h425d244f};
test_input[21456:21463] = '{32'hbfba0118, 32'hc26f5f2f, 32'h426fbd21, 32'hc2861850, 32'hc2c3d193, 32'h41c26ed0, 32'h4240ca66, 32'h4089f22f};
test_output[21456:21463] = '{32'h0, 32'h0, 32'h426fbd21, 32'h0, 32'h0, 32'h41c26ed0, 32'h4240ca66, 32'h4089f22f};
test_input[21464:21471] = '{32'h42bf6bc7, 32'h42105dfd, 32'hc2b303a7, 32'hc1e3c8e1, 32'hc1e958a2, 32'hc23d625c, 32'hc2813cdf, 32'hc29f6e8c};
test_output[21464:21471] = '{32'h42bf6bc7, 32'h42105dfd, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21472:21479] = '{32'h41a46004, 32'hc1cb91bb, 32'h41455cb6, 32'h42593ddc, 32'h427b25a2, 32'h429dcae3, 32'hc2b56d15, 32'hc25c6ffc};
test_output[21472:21479] = '{32'h41a46004, 32'h0, 32'h41455cb6, 32'h42593ddc, 32'h427b25a2, 32'h429dcae3, 32'h0, 32'h0};
test_input[21480:21487] = '{32'hc249c94b, 32'h42a4435b, 32'hc18a7d01, 32'h42c74aa1, 32'h421c423f, 32'h429f6bb2, 32'hc216e357, 32'h3e8913c8};
test_output[21480:21487] = '{32'h0, 32'h42a4435b, 32'h0, 32'h42c74aa1, 32'h421c423f, 32'h429f6bb2, 32'h0, 32'h3e8913c8};
test_input[21488:21495] = '{32'hc14a82d6, 32'h42ab5b4f, 32'hc27c017a, 32'h4287a1fc, 32'hc26f298a, 32'hc1848a58, 32'hc1b62da2, 32'h42b16eed};
test_output[21488:21495] = '{32'h0, 32'h42ab5b4f, 32'h0, 32'h4287a1fc, 32'h0, 32'h0, 32'h0, 32'h42b16eed};
test_input[21496:21503] = '{32'h40c74244, 32'hc1510a26, 32'hc254284c, 32'h421106e0, 32'h42b60606, 32'hc2a7551a, 32'hc29168b8, 32'hc260d3a0};
test_output[21496:21503] = '{32'h40c74244, 32'h0, 32'h0, 32'h421106e0, 32'h42b60606, 32'h0, 32'h0, 32'h0};
test_input[21504:21511] = '{32'hc1b51079, 32'hc2805279, 32'h42a0a653, 32'h42a06f69, 32'hc1b575ca, 32'h41d5a7a1, 32'hc243ec21, 32'h42a4358b};
test_output[21504:21511] = '{32'h0, 32'h0, 32'h42a0a653, 32'h42a06f69, 32'h0, 32'h41d5a7a1, 32'h0, 32'h42a4358b};
test_input[21512:21519] = '{32'h4282e6f1, 32'h42167c29, 32'h41a240b8, 32'hc0b454ca, 32'h420214b7, 32'h42219b44, 32'h429f8709, 32'hc25909fb};
test_output[21512:21519] = '{32'h4282e6f1, 32'h42167c29, 32'h41a240b8, 32'h0, 32'h420214b7, 32'h42219b44, 32'h429f8709, 32'h0};
test_input[21520:21527] = '{32'h427eb0e9, 32'hc2a03d79, 32'hc2a0efce, 32'hc2649c58, 32'h427c4fe9, 32'hc1204da0, 32'h4111669d, 32'h41c2b116};
test_output[21520:21527] = '{32'h427eb0e9, 32'h0, 32'h0, 32'h0, 32'h427c4fe9, 32'h0, 32'h4111669d, 32'h41c2b116};
test_input[21528:21535] = '{32'h4282a405, 32'h429b5def, 32'hc28dbfcd, 32'h4297afc7, 32'hc2a29658, 32'hc21a43cf, 32'hc237bfca, 32'hc1cdce67};
test_output[21528:21535] = '{32'h4282a405, 32'h429b5def, 32'h0, 32'h4297afc7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21536:21543] = '{32'hc2be025f, 32'h4204dafc, 32'hc0657df9, 32'h42bec0e4, 32'hc1103610, 32'h426ac409, 32'h4080610b, 32'hc0072de5};
test_output[21536:21543] = '{32'h0, 32'h4204dafc, 32'h0, 32'h42bec0e4, 32'h0, 32'h426ac409, 32'h4080610b, 32'h0};
test_input[21544:21551] = '{32'hc26e545a, 32'h428279ae, 32'h413cee8d, 32'h42b0b4ef, 32'h42170c1a, 32'hc182b285, 32'hc2024fc0, 32'hc2806fb7};
test_output[21544:21551] = '{32'h0, 32'h428279ae, 32'h413cee8d, 32'h42b0b4ef, 32'h42170c1a, 32'h0, 32'h0, 32'h0};
test_input[21552:21559] = '{32'h41e99bee, 32'h418d21a7, 32'hc1c81e0f, 32'hc247b975, 32'h416502c4, 32'h429e5f51, 32'hc16fce5f, 32'h42927ed9};
test_output[21552:21559] = '{32'h41e99bee, 32'h418d21a7, 32'h0, 32'h0, 32'h416502c4, 32'h429e5f51, 32'h0, 32'h42927ed9};
test_input[21560:21567] = '{32'hc1950423, 32'hc1bddc7c, 32'h41b0bfc3, 32'hc29dabfa, 32'h41070c7a, 32'h42a7e1f8, 32'h42986cbc, 32'h421aa45c};
test_output[21560:21567] = '{32'h0, 32'h0, 32'h41b0bfc3, 32'h0, 32'h41070c7a, 32'h42a7e1f8, 32'h42986cbc, 32'h421aa45c};
test_input[21568:21575] = '{32'hc2275d8e, 32'h40a78b65, 32'h427dd8c8, 32'hc23a138d, 32'hc168e898, 32'hc2984cfd, 32'h42a97add, 32'h4218a3ac};
test_output[21568:21575] = '{32'h0, 32'h40a78b65, 32'h427dd8c8, 32'h0, 32'h0, 32'h0, 32'h42a97add, 32'h4218a3ac};
test_input[21576:21583] = '{32'h42c78007, 32'h4210a91a, 32'h41a62533, 32'h42b79d25, 32'h42340bd5, 32'hc2746c46, 32'h42a0238f, 32'hc2a54ba2};
test_output[21576:21583] = '{32'h42c78007, 32'h4210a91a, 32'h41a62533, 32'h42b79d25, 32'h42340bd5, 32'h0, 32'h42a0238f, 32'h0};
test_input[21584:21591] = '{32'h426828f2, 32'h41354156, 32'h42989822, 32'h4293c8cf, 32'h42bee15c, 32'hc2815c85, 32'h42053aa1, 32'h42b50629};
test_output[21584:21591] = '{32'h426828f2, 32'h41354156, 32'h42989822, 32'h4293c8cf, 32'h42bee15c, 32'h0, 32'h42053aa1, 32'h42b50629};
test_input[21592:21599] = '{32'hc1d922e7, 32'h4217a4fd, 32'hc0276918, 32'h424591f0, 32'h42688f64, 32'hc2aac54e, 32'hc293f40f, 32'h41f7e846};
test_output[21592:21599] = '{32'h0, 32'h4217a4fd, 32'h0, 32'h424591f0, 32'h42688f64, 32'h0, 32'h0, 32'h41f7e846};
test_input[21600:21607] = '{32'h42b4976f, 32'hc2bd5b22, 32'hc144c04e, 32'h3e8ca0e4, 32'h428a7794, 32'h4117f44f, 32'h42360b97, 32'hc2a57031};
test_output[21600:21607] = '{32'h42b4976f, 32'h0, 32'h0, 32'h3e8ca0e4, 32'h428a7794, 32'h4117f44f, 32'h42360b97, 32'h0};
test_input[21608:21615] = '{32'h41a66160, 32'h4148ff51, 32'h41bb3580, 32'h424bd8db, 32'h42c7dae0, 32'h428266a9, 32'h41bbd5c8, 32'hc267d7ee};
test_output[21608:21615] = '{32'h41a66160, 32'h4148ff51, 32'h41bb3580, 32'h424bd8db, 32'h42c7dae0, 32'h428266a9, 32'h41bbd5c8, 32'h0};
test_input[21616:21623] = '{32'h428b7fee, 32'hc100a7a8, 32'hc1b93e35, 32'hc2b11666, 32'hc230907a, 32'hc2aa2999, 32'h4253a4a9, 32'h42b36868};
test_output[21616:21623] = '{32'h428b7fee, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4253a4a9, 32'h42b36868};
test_input[21624:21631] = '{32'hc2893a3d, 32'h428d1c1e, 32'hc1f53d5c, 32'h42b49f8d, 32'h4207ef97, 32'hc22a5c16, 32'h427e9261, 32'hc20b34ee};
test_output[21624:21631] = '{32'h0, 32'h428d1c1e, 32'h0, 32'h42b49f8d, 32'h4207ef97, 32'h0, 32'h427e9261, 32'h0};
test_input[21632:21639] = '{32'hc16abe33, 32'hc2837780, 32'hc26e9de7, 32'h419e29d7, 32'hc24381cb, 32'h428b9d1e, 32'h42299827, 32'h418eb181};
test_output[21632:21639] = '{32'h0, 32'h0, 32'h0, 32'h419e29d7, 32'h0, 32'h428b9d1e, 32'h42299827, 32'h418eb181};
test_input[21640:21647] = '{32'h42980009, 32'hc29a249a, 32'hc2aa3993, 32'h428b2e35, 32'h428c1b85, 32'hbff35a14, 32'h404a97c9, 32'h42a7a77a};
test_output[21640:21647] = '{32'h42980009, 32'h0, 32'h0, 32'h428b2e35, 32'h428c1b85, 32'h0, 32'h404a97c9, 32'h42a7a77a};
test_input[21648:21655] = '{32'h42309748, 32'hc212a80f, 32'h3fa04947, 32'h422bd4dd, 32'h42c61abd, 32'hc2259f62, 32'hc2a8c8c6, 32'h42beec61};
test_output[21648:21655] = '{32'h42309748, 32'h0, 32'h3fa04947, 32'h422bd4dd, 32'h42c61abd, 32'h0, 32'h0, 32'h42beec61};
test_input[21656:21663] = '{32'hc12222a3, 32'hc229dafa, 32'h4252a3d6, 32'h423f6e30, 32'hc18c1046, 32'h42a5fc4d, 32'hc1c9bed2, 32'hc2c5d2a2};
test_output[21656:21663] = '{32'h0, 32'h0, 32'h4252a3d6, 32'h423f6e30, 32'h0, 32'h42a5fc4d, 32'h0, 32'h0};
test_input[21664:21671] = '{32'h42aea595, 32'h42c7c863, 32'h42c097a0, 32'hc29f9de9, 32'hc27a93cc, 32'hc285ecbf, 32'hc2a30bec, 32'hc297501d};
test_output[21664:21671] = '{32'h42aea595, 32'h42c7c863, 32'h42c097a0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21672:21679] = '{32'h42936fff, 32'hc20ef26e, 32'h42c77b35, 32'hc288cb96, 32'hc1e3ce54, 32'hc2295ad2, 32'hc23d94df, 32'h425fd78e};
test_output[21672:21679] = '{32'h42936fff, 32'h0, 32'h42c77b35, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425fd78e};
test_input[21680:21687] = '{32'hc27fcccd, 32'h40aa0e96, 32'h4240c1e9, 32'h42387440, 32'h4207adff, 32'hc2ae105f, 32'h41a180a0, 32'hc2355f7a};
test_output[21680:21687] = '{32'h0, 32'h40aa0e96, 32'h4240c1e9, 32'h42387440, 32'h4207adff, 32'h0, 32'h41a180a0, 32'h0};
test_input[21688:21695] = '{32'h4282820e, 32'h423e7d15, 32'hc096e996, 32'hc29cde0b, 32'hc1c27e78, 32'h425934c9, 32'hc2577c87, 32'h40b7fa47};
test_output[21688:21695] = '{32'h4282820e, 32'h423e7d15, 32'h0, 32'h0, 32'h0, 32'h425934c9, 32'h0, 32'h40b7fa47};
test_input[21696:21703] = '{32'hc2942532, 32'h42c11b14, 32'h42a84d40, 32'hc2bbb56e, 32'hc2a06833, 32'h421efff9, 32'hc21a4185, 32'h3ea9a90d};
test_output[21696:21703] = '{32'h0, 32'h42c11b14, 32'h42a84d40, 32'h0, 32'h0, 32'h421efff9, 32'h0, 32'h3ea9a90d};
test_input[21704:21711] = '{32'h4076403b, 32'h42a72076, 32'hc2a3f355, 32'hc24e7a6f, 32'h4220bf34, 32'h42a9d770, 32'hc254f839, 32'h42b9ee26};
test_output[21704:21711] = '{32'h4076403b, 32'h42a72076, 32'h0, 32'h0, 32'h4220bf34, 32'h42a9d770, 32'h0, 32'h42b9ee26};
test_input[21712:21719] = '{32'h429da61c, 32'hc26d3ec4, 32'hc1c1047d, 32'hc27d5a55, 32'hc2b61963, 32'h3f91176d, 32'hc257fa97, 32'hc1c71777};
test_output[21712:21719] = '{32'h429da61c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3f91176d, 32'h0, 32'h0};
test_input[21720:21727] = '{32'hc090698b, 32'h42baaf26, 32'h4231b3ea, 32'h42bc5f69, 32'h415c25c4, 32'hc09916bb, 32'hc03d8031, 32'hc210ee3e};
test_output[21720:21727] = '{32'h0, 32'h42baaf26, 32'h4231b3ea, 32'h42bc5f69, 32'h415c25c4, 32'h0, 32'h0, 32'h0};
test_input[21728:21735] = '{32'h427ba955, 32'h42a9ffcd, 32'h42855c32, 32'h41ce4129, 32'hc2be90cf, 32'hc28172a1, 32'h426f1c79, 32'hc28e0f3f};
test_output[21728:21735] = '{32'h427ba955, 32'h42a9ffcd, 32'h42855c32, 32'h41ce4129, 32'h0, 32'h0, 32'h426f1c79, 32'h0};
test_input[21736:21743] = '{32'hc1e26a71, 32'hc1be2962, 32'h4172ac20, 32'hc224297a, 32'h419b986f, 32'hc1b483b1, 32'h42b2791b, 32'h3fcb3ec9};
test_output[21736:21743] = '{32'h0, 32'h0, 32'h4172ac20, 32'h0, 32'h419b986f, 32'h0, 32'h42b2791b, 32'h3fcb3ec9};
test_input[21744:21751] = '{32'hc202804d, 32'h42c4721d, 32'h4294b3b2, 32'hc242dc42, 32'h42c015ce, 32'h4149b8d2, 32'hc1820a00, 32'h42aa1f49};
test_output[21744:21751] = '{32'h0, 32'h42c4721d, 32'h4294b3b2, 32'h0, 32'h42c015ce, 32'h4149b8d2, 32'h0, 32'h42aa1f49};
test_input[21752:21759] = '{32'hc226277d, 32'h41a8f930, 32'hc268e9dd, 32'hc219b3a1, 32'hc2265477, 32'h42bc620a, 32'h424cb92c, 32'hc0ac9c96};
test_output[21752:21759] = '{32'h0, 32'h41a8f930, 32'h0, 32'h0, 32'h0, 32'h42bc620a, 32'h424cb92c, 32'h0};
test_input[21760:21767] = '{32'hc2b7e127, 32'hc2204348, 32'h4163dc42, 32'hc210ad38, 32'h42b4da56, 32'hc29053d6, 32'hc0ba40ac, 32'hc286b809};
test_output[21760:21767] = '{32'h0, 32'h0, 32'h4163dc42, 32'h0, 32'h42b4da56, 32'h0, 32'h0, 32'h0};
test_input[21768:21775] = '{32'h424f9319, 32'h4202cb1e, 32'h41f277a9, 32'h41495583, 32'h40a2f735, 32'h42a61c30, 32'hc283f536, 32'hc172aebb};
test_output[21768:21775] = '{32'h424f9319, 32'h4202cb1e, 32'h41f277a9, 32'h41495583, 32'h40a2f735, 32'h42a61c30, 32'h0, 32'h0};
test_input[21776:21783] = '{32'hc12258e5, 32'h4194791c, 32'h428c9446, 32'hc1853b4d, 32'h418b9476, 32'hc1cfaa24, 32'h40722844, 32'h42bd492d};
test_output[21776:21783] = '{32'h0, 32'h4194791c, 32'h428c9446, 32'h0, 32'h418b9476, 32'h0, 32'h40722844, 32'h42bd492d};
test_input[21784:21791] = '{32'h427577bf, 32'h41720de9, 32'h421e80c9, 32'hc1f154a2, 32'h42ae2f18, 32'h414b67f9, 32'h42a861c6, 32'hc0addeb0};
test_output[21784:21791] = '{32'h427577bf, 32'h41720de9, 32'h421e80c9, 32'h0, 32'h42ae2f18, 32'h414b67f9, 32'h42a861c6, 32'h0};
test_input[21792:21799] = '{32'h41edbb6e, 32'hc28b7c22, 32'h42b67224, 32'hc2728405, 32'hc2453351, 32'h424a19e8, 32'hc199c913, 32'h429d493b};
test_output[21792:21799] = '{32'h41edbb6e, 32'h0, 32'h42b67224, 32'h0, 32'h0, 32'h424a19e8, 32'h0, 32'h429d493b};
test_input[21800:21807] = '{32'h42c6afb2, 32'hc23ac274, 32'h42a7008d, 32'h42316ab7, 32'h429eca6a, 32'h4278eaca, 32'h413ed515, 32'h41eb7dd5};
test_output[21800:21807] = '{32'h42c6afb2, 32'h0, 32'h42a7008d, 32'h42316ab7, 32'h429eca6a, 32'h4278eaca, 32'h413ed515, 32'h41eb7dd5};
test_input[21808:21815] = '{32'h41e4a09e, 32'h402cb0ea, 32'h4298a848, 32'hc2b85349, 32'hc14a3f41, 32'h42c1f13a, 32'h42a11670, 32'h41947903};
test_output[21808:21815] = '{32'h41e4a09e, 32'h402cb0ea, 32'h4298a848, 32'h0, 32'h0, 32'h42c1f13a, 32'h42a11670, 32'h41947903};
test_input[21816:21823] = '{32'hc2c74d63, 32'h42a73058, 32'h3fe7ba6e, 32'h42c39e03, 32'h42815743, 32'hc29e43d3, 32'h42820578, 32'h42c41b80};
test_output[21816:21823] = '{32'h0, 32'h42a73058, 32'h3fe7ba6e, 32'h42c39e03, 32'h42815743, 32'h0, 32'h42820578, 32'h42c41b80};
test_input[21824:21831] = '{32'h429566e7, 32'hc29e4927, 32'h3f8f1c84, 32'hc2850e36, 32'h410dc34d, 32'h429d136d, 32'h421c5efe, 32'h42841f22};
test_output[21824:21831] = '{32'h429566e7, 32'h0, 32'h3f8f1c84, 32'h0, 32'h410dc34d, 32'h429d136d, 32'h421c5efe, 32'h42841f22};
test_input[21832:21839] = '{32'h40db5ada, 32'h40e1255a, 32'h42a614ee, 32'hc240df99, 32'h41ca5e29, 32'hc01c35ca, 32'hc249cede, 32'hc2920d2e};
test_output[21832:21839] = '{32'h40db5ada, 32'h40e1255a, 32'h42a614ee, 32'h0, 32'h41ca5e29, 32'h0, 32'h0, 32'h0};
test_input[21840:21847] = '{32'h42bc829b, 32'h42a23c61, 32'h42923907, 32'hc21f7674, 32'hc2baa5ef, 32'h4286df36, 32'hc1c4d95e, 32'hc1a442db};
test_output[21840:21847] = '{32'h42bc829b, 32'h42a23c61, 32'h42923907, 32'h0, 32'h0, 32'h4286df36, 32'h0, 32'h0};
test_input[21848:21855] = '{32'h428f006f, 32'hc2a6b44e, 32'hc1f35830, 32'hc2290094, 32'hc2c34e5b, 32'h42b51535, 32'hc209c680, 32'h42535f16};
test_output[21848:21855] = '{32'h428f006f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b51535, 32'h0, 32'h42535f16};
test_input[21856:21863] = '{32'hc1b528d0, 32'hc23ce8d0, 32'h42700c22, 32'hc2c39393, 32'h4220b3e0, 32'hc1a0b349, 32'h427f5567, 32'hc2b97b66};
test_output[21856:21863] = '{32'h0, 32'h0, 32'h42700c22, 32'h0, 32'h4220b3e0, 32'h0, 32'h427f5567, 32'h0};
test_input[21864:21871] = '{32'h4251583f, 32'h41412356, 32'hc2c0237a, 32'h42be36d8, 32'h428fc4cd, 32'hc221deab, 32'h42862dc8, 32'h4294cb8c};
test_output[21864:21871] = '{32'h4251583f, 32'h41412356, 32'h0, 32'h42be36d8, 32'h428fc4cd, 32'h0, 32'h42862dc8, 32'h4294cb8c};
test_input[21872:21879] = '{32'hc2a7669d, 32'h414509b9, 32'h41a33930, 32'hc19bafd1, 32'hbfccede1, 32'hc18a3704, 32'hc257eab5, 32'h42bcdc6a};
test_output[21872:21879] = '{32'h0, 32'h414509b9, 32'h41a33930, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bcdc6a};
test_input[21880:21887] = '{32'hc2c7dce0, 32'hc25783b8, 32'hc2a43d7b, 32'hc2237b21, 32'h415c4ecb, 32'h40528d48, 32'hc2b59bdf, 32'hc2113b42};
test_output[21880:21887] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h415c4ecb, 32'h40528d48, 32'h0, 32'h0};
test_input[21888:21895] = '{32'h4256698f, 32'h4194387f, 32'hc2b3b499, 32'hc2b8f4be, 32'hc216caaa, 32'hc1668614, 32'hc2c3ffe4, 32'hc2c4ebe6};
test_output[21888:21895] = '{32'h4256698f, 32'h4194387f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21896:21903] = '{32'hc13b473c, 32'h427e5dd1, 32'h422e28d9, 32'hc212315b, 32'hc10c684b, 32'h426af4da, 32'hc2010619, 32'h429e3a28};
test_output[21896:21903] = '{32'h0, 32'h427e5dd1, 32'h422e28d9, 32'h0, 32'h0, 32'h426af4da, 32'h0, 32'h429e3a28};
test_input[21904:21911] = '{32'hc1c4f83d, 32'h41ed5acf, 32'hc26e633f, 32'h42761557, 32'hc229eadb, 32'h42a484ab, 32'hc2be224f, 32'h421f419f};
test_output[21904:21911] = '{32'h0, 32'h41ed5acf, 32'h0, 32'h42761557, 32'h0, 32'h42a484ab, 32'h0, 32'h421f419f};
test_input[21912:21919] = '{32'h422e6948, 32'hc29c1c05, 32'h41c43632, 32'hc1d03f93, 32'hc29ecbe7, 32'hc12e4f3f, 32'hc289b205, 32'h413f68e7};
test_output[21912:21919] = '{32'h422e6948, 32'h0, 32'h41c43632, 32'h0, 32'h0, 32'h0, 32'h0, 32'h413f68e7};
test_input[21920:21927] = '{32'hc293f09c, 32'hc2841641, 32'hc287e0a8, 32'h4296af42, 32'h4224438e, 32'hc2a087ed, 32'hc27fde97, 32'h42bfde65};
test_output[21920:21927] = '{32'h0, 32'h0, 32'h0, 32'h4296af42, 32'h4224438e, 32'h0, 32'h0, 32'h42bfde65};
test_input[21928:21935] = '{32'hc0d5188c, 32'h42325d0f, 32'hc28ac5a0, 32'h42ae504a, 32'h42453739, 32'hc238c78d, 32'h41e9a637, 32'hc13b045c};
test_output[21928:21935] = '{32'h0, 32'h42325d0f, 32'h0, 32'h42ae504a, 32'h42453739, 32'h0, 32'h41e9a637, 32'h0};
test_input[21936:21943] = '{32'h4095e962, 32'hc17437a0, 32'hc23fcb18, 32'h41cfa5d2, 32'h3f9d5e3c, 32'hc21c81c4, 32'hc2a9a5b9, 32'h421779b2};
test_output[21936:21943] = '{32'h4095e962, 32'h0, 32'h0, 32'h41cfa5d2, 32'h3f9d5e3c, 32'h0, 32'h0, 32'h421779b2};
test_input[21944:21951] = '{32'hc2b1f8f7, 32'hc28eb7f2, 32'h42c478f4, 32'h40baab0e, 32'h42b495a4, 32'h41fbbf06, 32'h418d7c98, 32'hc2540173};
test_output[21944:21951] = '{32'h0, 32'h0, 32'h42c478f4, 32'h40baab0e, 32'h42b495a4, 32'h41fbbf06, 32'h418d7c98, 32'h0};
test_input[21952:21959] = '{32'h42a3b70a, 32'h428bf6f0, 32'hc2828e1e, 32'hc2b886a7, 32'hc2aa6312, 32'hc2a2f105, 32'h425eef13, 32'hc2c2f285};
test_output[21952:21959] = '{32'h42a3b70a, 32'h428bf6f0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425eef13, 32'h0};
test_input[21960:21967] = '{32'hc251c81a, 32'h42158b3d, 32'hc202c756, 32'hc222178f, 32'hc2a2edf2, 32'hc2beec64, 32'hc2399397, 32'hc23156a6};
test_output[21960:21967] = '{32'h0, 32'h42158b3d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21968:21975] = '{32'hc2a27643, 32'h4226133c, 32'hc2952118, 32'h42c3d578, 32'h42c3d654, 32'h421e8248, 32'h42921719, 32'h4139ce0d};
test_output[21968:21975] = '{32'h0, 32'h4226133c, 32'h0, 32'h42c3d578, 32'h42c3d654, 32'h421e8248, 32'h42921719, 32'h4139ce0d};
test_input[21976:21983] = '{32'h41eac42c, 32'hc2389098, 32'hc2a5f07a, 32'h42ad65ab, 32'h41047d36, 32'hc130c8cd, 32'h42ba1b7f, 32'h4200b568};
test_output[21976:21983] = '{32'h41eac42c, 32'h0, 32'h0, 32'h42ad65ab, 32'h41047d36, 32'h0, 32'h42ba1b7f, 32'h4200b568};
test_input[21984:21991] = '{32'h42574fe1, 32'h429d0332, 32'hc2991381, 32'hc2b48674, 32'h41b045fe, 32'h4259ddc9, 32'h41fac5bb, 32'hc2aa033b};
test_output[21984:21991] = '{32'h42574fe1, 32'h429d0332, 32'h0, 32'h0, 32'h41b045fe, 32'h4259ddc9, 32'h41fac5bb, 32'h0};
test_input[21992:21999] = '{32'h4250a650, 32'h42b806ba, 32'hc2a28e90, 32'hc277e432, 32'h425fe82d, 32'hc1dd1920, 32'hc1b203ba, 32'h42936e60};
test_output[21992:21999] = '{32'h4250a650, 32'h42b806ba, 32'h0, 32'h0, 32'h425fe82d, 32'h0, 32'h0, 32'h42936e60};
test_input[22000:22007] = '{32'h42c2b1b6, 32'h42879f1f, 32'h41269f69, 32'h429908dd, 32'hbeb9e8d4, 32'hc2ab0453, 32'h41f78bce, 32'h42bdf64c};
test_output[22000:22007] = '{32'h42c2b1b6, 32'h42879f1f, 32'h41269f69, 32'h429908dd, 32'h0, 32'h0, 32'h41f78bce, 32'h42bdf64c};
test_input[22008:22015] = '{32'h42b1af51, 32'h42a2ef88, 32'hc2ad5891, 32'h42b62125, 32'h418f70f2, 32'hc2a9882b, 32'h421438eb, 32'hc20070cc};
test_output[22008:22015] = '{32'h42b1af51, 32'h42a2ef88, 32'h0, 32'h42b62125, 32'h418f70f2, 32'h0, 32'h421438eb, 32'h0};
test_input[22016:22023] = '{32'h425df33b, 32'h41fe596b, 32'hc23832a7, 32'hc2839a82, 32'h4211edb3, 32'h429abff8, 32'hc2adc388, 32'hc01b0da5};
test_output[22016:22023] = '{32'h425df33b, 32'h41fe596b, 32'h0, 32'h0, 32'h4211edb3, 32'h429abff8, 32'h0, 32'h0};
test_input[22024:22031] = '{32'hc18e9664, 32'hc2a8ded4, 32'h42b6533c, 32'hc2504875, 32'h411c07e0, 32'hc0b2ea8d, 32'h42c27498, 32'h4113dac3};
test_output[22024:22031] = '{32'h0, 32'h0, 32'h42b6533c, 32'h0, 32'h411c07e0, 32'h0, 32'h42c27498, 32'h4113dac3};
test_input[22032:22039] = '{32'hc2a7aacd, 32'h42c3ef18, 32'h42ad6a29, 32'hc22e7532, 32'hc1cd007b, 32'hc2a1b816, 32'hc034fb5e, 32'h4291e2d9};
test_output[22032:22039] = '{32'h0, 32'h42c3ef18, 32'h42ad6a29, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4291e2d9};
test_input[22040:22047] = '{32'hc2a6d73a, 32'h42009776, 32'hc2c37bb7, 32'h4290c2a3, 32'h429fdbfb, 32'hc291a393, 32'h40866960, 32'h4136eddc};
test_output[22040:22047] = '{32'h0, 32'h42009776, 32'h0, 32'h4290c2a3, 32'h429fdbfb, 32'h0, 32'h40866960, 32'h4136eddc};
test_input[22048:22055] = '{32'h41d9846f, 32'h428b8ef5, 32'hc0c10381, 32'hc200997a, 32'h427f9e11, 32'h4260e5df, 32'h42c26620, 32'hc29e742d};
test_output[22048:22055] = '{32'h41d9846f, 32'h428b8ef5, 32'h0, 32'h0, 32'h427f9e11, 32'h4260e5df, 32'h42c26620, 32'h0};
test_input[22056:22063] = '{32'hc2270da9, 32'hc2b86424, 32'hc248d255, 32'h4215fb75, 32'hc21f49d9, 32'hbd7676ce, 32'hc28adb44, 32'h422ee397};
test_output[22056:22063] = '{32'h0, 32'h0, 32'h0, 32'h4215fb75, 32'h0, 32'h0, 32'h0, 32'h422ee397};
test_input[22064:22071] = '{32'h40bfac03, 32'hc2729e71, 32'h429b6a16, 32'hc1199761, 32'hc126199d, 32'hc2454480, 32'h429776ce, 32'h4272d702};
test_output[22064:22071] = '{32'h40bfac03, 32'h0, 32'h429b6a16, 32'h0, 32'h0, 32'h0, 32'h429776ce, 32'h4272d702};
test_input[22072:22079] = '{32'h428f468b, 32'h40e17cd8, 32'hc227a69b, 32'h3ffc16ca, 32'h42bb4207, 32'h41b3ef06, 32'hc21d68e5, 32'hc2165d51};
test_output[22072:22079] = '{32'h428f468b, 32'h40e17cd8, 32'h0, 32'h3ffc16ca, 32'h42bb4207, 32'h41b3ef06, 32'h0, 32'h0};
test_input[22080:22087] = '{32'h42950b51, 32'h426bc7ae, 32'hc0649a7d, 32'hc2659b39, 32'h4222ef1a, 32'hc1ed6cc1, 32'h41daad68, 32'h4085f602};
test_output[22080:22087] = '{32'h42950b51, 32'h426bc7ae, 32'h0, 32'h0, 32'h4222ef1a, 32'h0, 32'h41daad68, 32'h4085f602};
test_input[22088:22095] = '{32'h4299a441, 32'hc2486190, 32'hc24d13d2, 32'h414f2469, 32'hc2c637de, 32'hc2185682, 32'hc29075aa, 32'h429ec6bd};
test_output[22088:22095] = '{32'h4299a441, 32'h0, 32'h0, 32'h414f2469, 32'h0, 32'h0, 32'h0, 32'h429ec6bd};
test_input[22096:22103] = '{32'hc24eb8b7, 32'h422f90f4, 32'h428db51c, 32'h3fc21112, 32'h42210fd3, 32'h413b4452, 32'h418914a6, 32'hbfb604d7};
test_output[22096:22103] = '{32'h0, 32'h422f90f4, 32'h428db51c, 32'h3fc21112, 32'h42210fd3, 32'h413b4452, 32'h418914a6, 32'h0};
test_input[22104:22111] = '{32'h41f5aeac, 32'h429f6b0a, 32'h42c4f72d, 32'h42754708, 32'hc2535d2b, 32'hc213e5ec, 32'h42bc8928, 32'h42708e68};
test_output[22104:22111] = '{32'h41f5aeac, 32'h429f6b0a, 32'h42c4f72d, 32'h42754708, 32'h0, 32'h0, 32'h42bc8928, 32'h42708e68};
test_input[22112:22119] = '{32'hc293d0c3, 32'hc1dac629, 32'h40996c28, 32'h41dba348, 32'hc264dd47, 32'h4271988e, 32'hc2185b3c, 32'hc0378c6a};
test_output[22112:22119] = '{32'h0, 32'h0, 32'h40996c28, 32'h41dba348, 32'h0, 32'h4271988e, 32'h0, 32'h0};
test_input[22120:22127] = '{32'hc12ea61c, 32'h41ce14d0, 32'hc18a88fb, 32'hc2405e69, 32'h411915a6, 32'h42a88b96, 32'hc226ef72, 32'h42909200};
test_output[22120:22127] = '{32'h0, 32'h41ce14d0, 32'h0, 32'h0, 32'h411915a6, 32'h42a88b96, 32'h0, 32'h42909200};
test_input[22128:22135] = '{32'h42b3b1f4, 32'h422d7b13, 32'hc2918339, 32'h42993250, 32'h410df8b7, 32'hc0d7cf08, 32'hc230554b, 32'h42bf451a};
test_output[22128:22135] = '{32'h42b3b1f4, 32'h422d7b13, 32'h0, 32'h42993250, 32'h410df8b7, 32'h0, 32'h0, 32'h42bf451a};
test_input[22136:22143] = '{32'hc238aeec, 32'hc106622d, 32'h425f10e5, 32'hc25670fb, 32'hc2bddf9c, 32'hc24ec0a0, 32'hc2827ba7, 32'h42932d94};
test_output[22136:22143] = '{32'h0, 32'h0, 32'h425f10e5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42932d94};
test_input[22144:22151] = '{32'hc2bc4234, 32'hc09ad69a, 32'h41df1ec7, 32'h4192d36e, 32'hc1d46227, 32'h41fdf853, 32'hc2602a40, 32'hc1c74475};
test_output[22144:22151] = '{32'h0, 32'h0, 32'h41df1ec7, 32'h4192d36e, 32'h0, 32'h41fdf853, 32'h0, 32'h0};
test_input[22152:22159] = '{32'h42699277, 32'hc25eefaa, 32'hc20bbd01, 32'h413924a9, 32'h429c1e01, 32'hc06a2a0f, 32'h427c5091, 32'h42377a84};
test_output[22152:22159] = '{32'h42699277, 32'h0, 32'h0, 32'h413924a9, 32'h429c1e01, 32'h0, 32'h427c5091, 32'h42377a84};
test_input[22160:22167] = '{32'h428df575, 32'hc297b592, 32'hc1706855, 32'h4281ee09, 32'h42988aec, 32'hc0b55551, 32'h42b6b674, 32'h420db0fb};
test_output[22160:22167] = '{32'h428df575, 32'h0, 32'h0, 32'h4281ee09, 32'h42988aec, 32'h0, 32'h42b6b674, 32'h420db0fb};
test_input[22168:22175] = '{32'h42a71021, 32'hc2511ad1, 32'hc2ae598d, 32'hc225198d, 32'h42aff2ce, 32'hc2bba87a, 32'hc24bb15b, 32'h424d7c37};
test_output[22168:22175] = '{32'h42a71021, 32'h0, 32'h0, 32'h0, 32'h42aff2ce, 32'h0, 32'h0, 32'h424d7c37};
test_input[22176:22183] = '{32'h4293e270, 32'hc15fbb10, 32'h428885ff, 32'hc2b7bba3, 32'h41e708b7, 32'h429c2eeb, 32'hc2c4914a, 32'h428863d4};
test_output[22176:22183] = '{32'h4293e270, 32'h0, 32'h428885ff, 32'h0, 32'h41e708b7, 32'h429c2eeb, 32'h0, 32'h428863d4};
test_input[22184:22191] = '{32'h41f5957c, 32'h42655d46, 32'hc135a0ca, 32'hc1c9093f, 32'hc2a1172b, 32'hc27bd31d, 32'h413d0b09, 32'h40b7d2b2};
test_output[22184:22191] = '{32'h41f5957c, 32'h42655d46, 32'h0, 32'h0, 32'h0, 32'h0, 32'h413d0b09, 32'h40b7d2b2};
test_input[22192:22199] = '{32'h425121c1, 32'h41ba05a8, 32'h42bf9287, 32'hc2346c96, 32'hc255cf32, 32'h42894c5d, 32'h429f8ff5, 32'hc29d91d2};
test_output[22192:22199] = '{32'h425121c1, 32'h41ba05a8, 32'h42bf9287, 32'h0, 32'h0, 32'h42894c5d, 32'h429f8ff5, 32'h0};
test_input[22200:22207] = '{32'h424b984e, 32'hc1d7b714, 32'h42a0b451, 32'hc2126fb2, 32'h4211f559, 32'h42c0a855, 32'hc21deab2, 32'hc23a32bf};
test_output[22200:22207] = '{32'h424b984e, 32'h0, 32'h42a0b451, 32'h0, 32'h4211f559, 32'h42c0a855, 32'h0, 32'h0};
test_input[22208:22215] = '{32'hc27fc0e2, 32'h429fa67d, 32'hc219cf93, 32'h414277f9, 32'h42632803, 32'hc249fd83, 32'h42be494d, 32'h4286d26e};
test_output[22208:22215] = '{32'h0, 32'h429fa67d, 32'h0, 32'h414277f9, 32'h42632803, 32'h0, 32'h42be494d, 32'h4286d26e};
test_input[22216:22223] = '{32'h428c2bf8, 32'hc2386005, 32'h405b23cf, 32'hc2c76579, 32'h4267ea28, 32'hc2c0b8d1, 32'h40ae85f2, 32'hbeeaf634};
test_output[22216:22223] = '{32'h428c2bf8, 32'h0, 32'h405b23cf, 32'h0, 32'h4267ea28, 32'h0, 32'h40ae85f2, 32'h0};
test_input[22224:22231] = '{32'h420a2132, 32'h42aa67e7, 32'h40acedf6, 32'hc272e2d4, 32'hc25a6ad8, 32'hc29f7c56, 32'hc19d6919, 32'hc1ea18d8};
test_output[22224:22231] = '{32'h420a2132, 32'h42aa67e7, 32'h40acedf6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22232:22239] = '{32'hc0368b5f, 32'h410bd352, 32'h42c5f5b6, 32'h40dd8653, 32'hc2381c3a, 32'h425369a8, 32'h410764c2, 32'hc2aedea0};
test_output[22232:22239] = '{32'h0, 32'h410bd352, 32'h42c5f5b6, 32'h40dd8653, 32'h0, 32'h425369a8, 32'h410764c2, 32'h0};
test_input[22240:22247] = '{32'h4223d574, 32'hc21b27ae, 32'hc0ec2171, 32'hc23e70b1, 32'hc118aa26, 32'hc1d65078, 32'hc29fc77f, 32'h4270afb5};
test_output[22240:22247] = '{32'h4223d574, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4270afb5};
test_input[22248:22255] = '{32'h41cb46f7, 32'hc194c381, 32'h42a0331b, 32'h42a754dc, 32'h42632b48, 32'hc2b6f9eb, 32'hbfd59377, 32'hc2618aa5};
test_output[22248:22255] = '{32'h41cb46f7, 32'h0, 32'h42a0331b, 32'h42a754dc, 32'h42632b48, 32'h0, 32'h0, 32'h0};
test_input[22256:22263] = '{32'h42819ce6, 32'h4227d1b3, 32'hc1990dda, 32'h405e699a, 32'h411f95da, 32'hc29bc9c7, 32'h41c79400, 32'h40b46ca3};
test_output[22256:22263] = '{32'h42819ce6, 32'h4227d1b3, 32'h0, 32'h405e699a, 32'h411f95da, 32'h0, 32'h41c79400, 32'h40b46ca3};
test_input[22264:22271] = '{32'h42a4d6d7, 32'hc2adb514, 32'h42c2e0fa, 32'hc1628228, 32'hc1dcb041, 32'h41ad6fde, 32'h42bb2656, 32'h4283ff15};
test_output[22264:22271] = '{32'h42a4d6d7, 32'h0, 32'h42c2e0fa, 32'h0, 32'h0, 32'h41ad6fde, 32'h42bb2656, 32'h4283ff15};
test_input[22272:22279] = '{32'hc280f54a, 32'hc25ebb77, 32'h42998912, 32'h42182c77, 32'h42b7b05c, 32'hc1db3342, 32'hc2a52934, 32'h42bfa1ae};
test_output[22272:22279] = '{32'h0, 32'h0, 32'h42998912, 32'h42182c77, 32'h42b7b05c, 32'h0, 32'h0, 32'h42bfa1ae};
test_input[22280:22287] = '{32'hc281a740, 32'h42165285, 32'hc2b85a76, 32'h402a1a49, 32'hc23d9ded, 32'h422df190, 32'h41bdc1c1, 32'h4281c3da};
test_output[22280:22287] = '{32'h0, 32'h42165285, 32'h0, 32'h402a1a49, 32'h0, 32'h422df190, 32'h41bdc1c1, 32'h4281c3da};
test_input[22288:22295] = '{32'hc23401ca, 32'hc2c3f7c3, 32'h4141e25e, 32'h42c54671, 32'h42960d3a, 32'h428d77b2, 32'h4270af9b, 32'h42ba3bbf};
test_output[22288:22295] = '{32'h0, 32'h0, 32'h4141e25e, 32'h42c54671, 32'h42960d3a, 32'h428d77b2, 32'h4270af9b, 32'h42ba3bbf};
test_input[22296:22303] = '{32'h42bf7d82, 32'hc2310597, 32'hbfde521e, 32'hc293c25a, 32'hc26fece4, 32'h42a9e338, 32'hc2254fba, 32'h40688cbd};
test_output[22296:22303] = '{32'h42bf7d82, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a9e338, 32'h0, 32'h40688cbd};
test_input[22304:22311] = '{32'hc1e09dfd, 32'hc25880f3, 32'hc2460a8d, 32'hc1585bfa, 32'h42120f6b, 32'h42c19303, 32'h420ec73f, 32'hc2934109};
test_output[22304:22311] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42120f6b, 32'h42c19303, 32'h420ec73f, 32'h0};
test_input[22312:22319] = '{32'hc2c50860, 32'hc2a97e97, 32'hc2871408, 32'h42875d43, 32'hbfeb1675, 32'h41f5574b, 32'h4166a2d8, 32'hbf0e2766};
test_output[22312:22319] = '{32'h0, 32'h0, 32'h0, 32'h42875d43, 32'h0, 32'h41f5574b, 32'h4166a2d8, 32'h0};
test_input[22320:22327] = '{32'hc1bb514c, 32'hc2318900, 32'h422c9886, 32'h41f3de0e, 32'hc23f38e7, 32'h41ea6859, 32'h416a5bca, 32'h41665d4e};
test_output[22320:22327] = '{32'h0, 32'h0, 32'h422c9886, 32'h41f3de0e, 32'h0, 32'h41ea6859, 32'h416a5bca, 32'h41665d4e};
test_input[22328:22335] = '{32'h41ce19fc, 32'hc1f7e8c8, 32'h42872be2, 32'h4238f5f9, 32'h42a240fa, 32'h419ca97a, 32'hc246129e, 32'hc2b24e4d};
test_output[22328:22335] = '{32'h41ce19fc, 32'h0, 32'h42872be2, 32'h4238f5f9, 32'h42a240fa, 32'h419ca97a, 32'h0, 32'h0};
test_input[22336:22343] = '{32'hc2984e98, 32'h41b52ea8, 32'h41adc15b, 32'h4298ca59, 32'hc28c014f, 32'h42b0557c, 32'hc20dfa5f, 32'h42c0096d};
test_output[22336:22343] = '{32'h0, 32'h41b52ea8, 32'h41adc15b, 32'h4298ca59, 32'h0, 32'h42b0557c, 32'h0, 32'h42c0096d};
test_input[22344:22351] = '{32'hc2420eeb, 32'h41dd127b, 32'h4236e507, 32'h423722bc, 32'hc188cfb8, 32'hc28170b8, 32'h40858e25, 32'hc1ddf563};
test_output[22344:22351] = '{32'h0, 32'h41dd127b, 32'h4236e507, 32'h423722bc, 32'h0, 32'h0, 32'h40858e25, 32'h0};
test_input[22352:22359] = '{32'h426de592, 32'hc229fa9f, 32'hc287648b, 32'hc205ca94, 32'hc2c3bad4, 32'hc19d36cb, 32'h422961c7, 32'h411d8be0};
test_output[22352:22359] = '{32'h426de592, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422961c7, 32'h411d8be0};
test_input[22360:22367] = '{32'hc1d1840f, 32'h41704936, 32'h41797ade, 32'hc16c2e82, 32'h420af776, 32'h42c3fea9, 32'h424e1e7b, 32'h41fba913};
test_output[22360:22367] = '{32'h0, 32'h41704936, 32'h41797ade, 32'h0, 32'h420af776, 32'h42c3fea9, 32'h424e1e7b, 32'h41fba913};
test_input[22368:22375] = '{32'h427b171b, 32'h418071ad, 32'hc28af863, 32'hc22db339, 32'hc1d3af29, 32'h429e4339, 32'hc23c86d4, 32'h409c1d40};
test_output[22368:22375] = '{32'h427b171b, 32'h418071ad, 32'h0, 32'h0, 32'h0, 32'h429e4339, 32'h0, 32'h409c1d40};
test_input[22376:22383] = '{32'h429c3918, 32'hc227314e, 32'hc23a1cd8, 32'h416447aa, 32'hc1be7377, 32'h42aa4b40, 32'h4237d0ca, 32'h41584bc3};
test_output[22376:22383] = '{32'h429c3918, 32'h0, 32'h0, 32'h416447aa, 32'h0, 32'h42aa4b40, 32'h4237d0ca, 32'h41584bc3};
test_input[22384:22391] = '{32'h423a530e, 32'hbfd42f0f, 32'h42b38f53, 32'hbff8fd5e, 32'hc1d70101, 32'hc227c2c0, 32'h41d675c6, 32'hc189bde6};
test_output[22384:22391] = '{32'h423a530e, 32'h0, 32'h42b38f53, 32'h0, 32'h0, 32'h0, 32'h41d675c6, 32'h0};
test_input[22392:22399] = '{32'hc26f7eae, 32'hc20f6ce6, 32'hc2ad6472, 32'h42423e6c, 32'hc1894af7, 32'hc10cea31, 32'hc2a626e2, 32'hc2b8f96c};
test_output[22392:22399] = '{32'h0, 32'h0, 32'h0, 32'h42423e6c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22400:22407] = '{32'hc18d9967, 32'h4175b77a, 32'h4290c6b7, 32'hc22514cd, 32'hc2085374, 32'hc2abbae7, 32'h40abeb5c, 32'hc2a92ab8};
test_output[22400:22407] = '{32'h0, 32'h4175b77a, 32'h4290c6b7, 32'h0, 32'h0, 32'h0, 32'h40abeb5c, 32'h0};
test_input[22408:22415] = '{32'h41f4422e, 32'h3f5182a6, 32'h41d67055, 32'hc2c3c80e, 32'hc2b1b535, 32'h41255c14, 32'hc25d0e11, 32'h41969f5d};
test_output[22408:22415] = '{32'h41f4422e, 32'h3f5182a6, 32'h41d67055, 32'h0, 32'h0, 32'h41255c14, 32'h0, 32'h41969f5d};
test_input[22416:22423] = '{32'hc17164e5, 32'h428681f0, 32'hc24a6268, 32'h425cd8c5, 32'h41fad3d7, 32'h42aed4b4, 32'h4295e244, 32'hc2b04ba2};
test_output[22416:22423] = '{32'h0, 32'h428681f0, 32'h0, 32'h425cd8c5, 32'h41fad3d7, 32'h42aed4b4, 32'h4295e244, 32'h0};
test_input[22424:22431] = '{32'h40c71f95, 32'h429d1434, 32'h426159f5, 32'h4258bccd, 32'hc111426d, 32'hc2c038bd, 32'hc2246db2, 32'h427b0a72};
test_output[22424:22431] = '{32'h40c71f95, 32'h429d1434, 32'h426159f5, 32'h4258bccd, 32'h0, 32'h0, 32'h0, 32'h427b0a72};
test_input[22432:22439] = '{32'hc1ec7343, 32'hc1c4eb89, 32'h42bf67c6, 32'h41597447, 32'h414fc014, 32'h3e980df8, 32'hc28dce4c, 32'hc235d78a};
test_output[22432:22439] = '{32'h0, 32'h0, 32'h42bf67c6, 32'h41597447, 32'h414fc014, 32'h3e980df8, 32'h0, 32'h0};
test_input[22440:22447] = '{32'hc2c6b722, 32'h4219cdc4, 32'h41d3adcc, 32'hc2a75ff6, 32'h41992314, 32'hc296d896, 32'h4158a468, 32'h42818052};
test_output[22440:22447] = '{32'h0, 32'h4219cdc4, 32'h41d3adcc, 32'h0, 32'h41992314, 32'h0, 32'h4158a468, 32'h42818052};
test_input[22448:22455] = '{32'hc134cd0c, 32'h4293bcd9, 32'hc1d01efc, 32'h42a5fefc, 32'h42b2ede1, 32'hc2c15e3e, 32'h42a5f4d7, 32'hc1b91abb};
test_output[22448:22455] = '{32'h0, 32'h4293bcd9, 32'h0, 32'h42a5fefc, 32'h42b2ede1, 32'h0, 32'h42a5f4d7, 32'h0};
test_input[22456:22463] = '{32'h41a392a0, 32'hc20954bc, 32'hc2b43832, 32'h4177e097, 32'hc09a5d84, 32'hc27e341f, 32'h41f5e4c3, 32'hc29b8516};
test_output[22456:22463] = '{32'h41a392a0, 32'h0, 32'h0, 32'h4177e097, 32'h0, 32'h0, 32'h41f5e4c3, 32'h0};
test_input[22464:22471] = '{32'hc231786a, 32'hc105da36, 32'h41577ea7, 32'h415675db, 32'hc2b3f9e2, 32'h42c29272, 32'hc2c3b515, 32'h41a31aff};
test_output[22464:22471] = '{32'h0, 32'h0, 32'h41577ea7, 32'h415675db, 32'h0, 32'h42c29272, 32'h0, 32'h41a31aff};
test_input[22472:22479] = '{32'h429daa2d, 32'h42a032a8, 32'h42450b31, 32'hc230ee6c, 32'hc197b6df, 32'h415fde3d, 32'h41ff559c, 32'hc203bd50};
test_output[22472:22479] = '{32'h429daa2d, 32'h42a032a8, 32'h42450b31, 32'h0, 32'h0, 32'h415fde3d, 32'h41ff559c, 32'h0};
test_input[22480:22487] = '{32'hc287dde8, 32'h41dcb3d7, 32'hc20755fa, 32'hc292646a, 32'h42c5f510, 32'hc2019485, 32'hc1a50def, 32'hc2823910};
test_output[22480:22487] = '{32'h0, 32'h41dcb3d7, 32'h0, 32'h0, 32'h42c5f510, 32'h0, 32'h0, 32'h0};
test_input[22488:22495] = '{32'hc03b73d7, 32'h4191435a, 32'h4274c620, 32'hc2b73f69, 32'hc1a43ae9, 32'h42856815, 32'h4256c656, 32'h42aa0980};
test_output[22488:22495] = '{32'h0, 32'h4191435a, 32'h4274c620, 32'h0, 32'h0, 32'h42856815, 32'h4256c656, 32'h42aa0980};
test_input[22496:22503] = '{32'hc27c0fc7, 32'hc29e7b75, 32'hc2a79353, 32'h41ab7028, 32'hc26fec82, 32'h3feb8590, 32'hc2313ec3, 32'h4251e4e1};
test_output[22496:22503] = '{32'h0, 32'h0, 32'h0, 32'h41ab7028, 32'h0, 32'h3feb8590, 32'h0, 32'h4251e4e1};
test_input[22504:22511] = '{32'hc200e0cc, 32'h3fd84f09, 32'hc189353d, 32'hc0860ec2, 32'hc0fde60f, 32'hc1986d97, 32'h4231458d, 32'h421cf7a1};
test_output[22504:22511] = '{32'h0, 32'h3fd84f09, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4231458d, 32'h421cf7a1};
test_input[22512:22519] = '{32'hc27a1732, 32'h429de037, 32'h42b55791, 32'h4251eef3, 32'h42b18efb, 32'hc2871069, 32'h429e83c3, 32'h3f904394};
test_output[22512:22519] = '{32'h0, 32'h429de037, 32'h42b55791, 32'h4251eef3, 32'h42b18efb, 32'h0, 32'h429e83c3, 32'h3f904394};
test_input[22520:22527] = '{32'h4227e3aa, 32'h425ac079, 32'h4291cb85, 32'hc1dada92, 32'h420bddca, 32'h42be7990, 32'hc24f0327, 32'h42b54fd7};
test_output[22520:22527] = '{32'h4227e3aa, 32'h425ac079, 32'h4291cb85, 32'h0, 32'h420bddca, 32'h42be7990, 32'h0, 32'h42b54fd7};
test_input[22528:22535] = '{32'hc28a7e49, 32'hc1d535f8, 32'hc2c466c7, 32'h41f4308b, 32'h4205fdc2, 32'hc227aa06, 32'h42bfe120, 32'h41dbf6c1};
test_output[22528:22535] = '{32'h0, 32'h0, 32'h0, 32'h41f4308b, 32'h4205fdc2, 32'h0, 32'h42bfe120, 32'h41dbf6c1};
test_input[22536:22543] = '{32'hc2551c29, 32'h41a0ccae, 32'hc1ba8498, 32'h4182a53f, 32'h3fa0cb78, 32'hc28e61bb, 32'hc260ae12, 32'h4172af9e};
test_output[22536:22543] = '{32'h0, 32'h41a0ccae, 32'h0, 32'h4182a53f, 32'h3fa0cb78, 32'h0, 32'h0, 32'h4172af9e};
test_input[22544:22551] = '{32'hc1164e48, 32'hc1873385, 32'h429ca7c8, 32'h41b7c8eb, 32'hc295af36, 32'h41c18533, 32'hc2977a02, 32'h429f246a};
test_output[22544:22551] = '{32'h0, 32'h0, 32'h429ca7c8, 32'h41b7c8eb, 32'h0, 32'h41c18533, 32'h0, 32'h429f246a};
test_input[22552:22559] = '{32'h41c06dd6, 32'hc21ac000, 32'h42950912, 32'hc10c36a8, 32'hc2a155d0, 32'hc1f13ef3, 32'h42abd85a, 32'hc2b376ca};
test_output[22552:22559] = '{32'h41c06dd6, 32'h0, 32'h42950912, 32'h0, 32'h0, 32'h0, 32'h42abd85a, 32'h0};
test_input[22560:22567] = '{32'hc29c275b, 32'hc2b531f3, 32'h42924395, 32'hc109b9c5, 32'hc1bcc873, 32'hc267c8a8, 32'hc1c2a1a9, 32'h41a86c54};
test_output[22560:22567] = '{32'h0, 32'h0, 32'h42924395, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41a86c54};
test_input[22568:22575] = '{32'h42946a77, 32'hc2be07ca, 32'h40991b53, 32'h41927e66, 32'h42841bd6, 32'h40aab866, 32'h42b504fc, 32'hc1ae416f};
test_output[22568:22575] = '{32'h42946a77, 32'h0, 32'h40991b53, 32'h41927e66, 32'h42841bd6, 32'h40aab866, 32'h42b504fc, 32'h0};
test_input[22576:22583] = '{32'h42836812, 32'hc255b6a8, 32'hc2b224ec, 32'hc24e30f9, 32'h41cb6cf0, 32'h3f4bbbf8, 32'h42b8cb8f, 32'hc1305693};
test_output[22576:22583] = '{32'h42836812, 32'h0, 32'h0, 32'h0, 32'h41cb6cf0, 32'h3f4bbbf8, 32'h42b8cb8f, 32'h0};
test_input[22584:22591] = '{32'hc267f2fd, 32'h423e090d, 32'hc22d7984, 32'h42b86f85, 32'h4258b897, 32'h42762d07, 32'h41aa0863, 32'hc0d06b9b};
test_output[22584:22591] = '{32'h0, 32'h423e090d, 32'h0, 32'h42b86f85, 32'h4258b897, 32'h42762d07, 32'h41aa0863, 32'h0};
test_input[22592:22599] = '{32'hc17296bb, 32'h42946de4, 32'hc09fbe48, 32'h42358d1e, 32'h4208df54, 32'h4151ccbc, 32'h425ab3dc, 32'hc2334848};
test_output[22592:22599] = '{32'h0, 32'h42946de4, 32'h0, 32'h42358d1e, 32'h4208df54, 32'h4151ccbc, 32'h425ab3dc, 32'h0};
test_input[22600:22607] = '{32'h427e6f22, 32'h4291ab79, 32'hc2684f42, 32'h429d2ebe, 32'h42c062b7, 32'h4263f0db, 32'h4234e0c0, 32'h4203f168};
test_output[22600:22607] = '{32'h427e6f22, 32'h4291ab79, 32'h0, 32'h429d2ebe, 32'h42c062b7, 32'h4263f0db, 32'h4234e0c0, 32'h4203f168};
test_input[22608:22615] = '{32'h42807e46, 32'hbcfaf557, 32'h4198d87e, 32'hc0b99d90, 32'h41a448f3, 32'h41ac292f, 32'hc2b10e04, 32'h41eb3d40};
test_output[22608:22615] = '{32'h42807e46, 32'h0, 32'h4198d87e, 32'h0, 32'h41a448f3, 32'h41ac292f, 32'h0, 32'h41eb3d40};
test_input[22616:22623] = '{32'hc1ceb259, 32'h4286bd9c, 32'h42a3ba34, 32'h42c382be, 32'h417dfdf7, 32'h41bece74, 32'hc11b387f, 32'h3ed9108b};
test_output[22616:22623] = '{32'h0, 32'h4286bd9c, 32'h42a3ba34, 32'h42c382be, 32'h417dfdf7, 32'h41bece74, 32'h0, 32'h3ed9108b};
test_input[22624:22631] = '{32'h4220d16d, 32'hc2c72f70, 32'hc1d29a02, 32'hc118450f, 32'hc25fdc84, 32'hc2039204, 32'hbf66cdae, 32'h42749749};
test_output[22624:22631] = '{32'h4220d16d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42749749};
test_input[22632:22639] = '{32'h42afa164, 32'h42c40d3a, 32'hc10f8305, 32'h423da4af, 32'h4202c7ee, 32'h41bfaae7, 32'hc2c481e0, 32'h416d3385};
test_output[22632:22639] = '{32'h42afa164, 32'h42c40d3a, 32'h0, 32'h423da4af, 32'h4202c7ee, 32'h41bfaae7, 32'h0, 32'h416d3385};
test_input[22640:22647] = '{32'h4282c6a0, 32'hc2c06bf8, 32'h42099fa9, 32'h4235c1d3, 32'hc279317e, 32'h4267174a, 32'h429a9cfd, 32'h41a15b01};
test_output[22640:22647] = '{32'h4282c6a0, 32'h0, 32'h42099fa9, 32'h4235c1d3, 32'h0, 32'h4267174a, 32'h429a9cfd, 32'h41a15b01};
test_input[22648:22655] = '{32'hc2ae812e, 32'h423aaa8b, 32'hc1cd9b8b, 32'hc2bcba5d, 32'h42b2a4c4, 32'h40a47e17, 32'hc2b3a996, 32'h422e05ad};
test_output[22648:22655] = '{32'h0, 32'h423aaa8b, 32'h0, 32'h0, 32'h42b2a4c4, 32'h40a47e17, 32'h0, 32'h422e05ad};
test_input[22656:22663] = '{32'hc2850d8f, 32'hc297f5dc, 32'h42a5a597, 32'h428b4603, 32'hc2bc9023, 32'h42b3cea6, 32'h421c035a, 32'hc23b2edc};
test_output[22656:22663] = '{32'h0, 32'h0, 32'h42a5a597, 32'h428b4603, 32'h0, 32'h42b3cea6, 32'h421c035a, 32'h0};
test_input[22664:22671] = '{32'hc2118156, 32'h426638b0, 32'hc202657f, 32'h428d259a, 32'h428517d6, 32'h42919091, 32'h426b5da4, 32'hc2039dc9};
test_output[22664:22671] = '{32'h0, 32'h426638b0, 32'h0, 32'h428d259a, 32'h428517d6, 32'h42919091, 32'h426b5da4, 32'h0};
test_input[22672:22679] = '{32'h4230042b, 32'h42a558ba, 32'hc2739712, 32'hc2070b68, 32'h4295b1b9, 32'hc1aa73a6, 32'h420cef7d, 32'h423cf227};
test_output[22672:22679] = '{32'h4230042b, 32'h42a558ba, 32'h0, 32'h0, 32'h4295b1b9, 32'h0, 32'h420cef7d, 32'h423cf227};
test_input[22680:22687] = '{32'hc1e19b7c, 32'hc2a18582, 32'h429a70d9, 32'hc206f103, 32'hc27a3c07, 32'hc2ad960d, 32'hc2aa6b2d, 32'hc2433364};
test_output[22680:22687] = '{32'h0, 32'h0, 32'h429a70d9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22688:22695] = '{32'h42bc76ae, 32'hc1f49ea0, 32'hc205509a, 32'hc208b078, 32'h425361f5, 32'h41aa28b0, 32'hc1880211, 32'hc083e555};
test_output[22688:22695] = '{32'h42bc76ae, 32'h0, 32'h0, 32'h0, 32'h425361f5, 32'h41aa28b0, 32'h0, 32'h0};
test_input[22696:22703] = '{32'hc223e90a, 32'h42068c26, 32'hc2a330b2, 32'h42441b79, 32'h41505685, 32'h41f1fbbf, 32'hc1e2c7eb, 32'h421289d5};
test_output[22696:22703] = '{32'h0, 32'h42068c26, 32'h0, 32'h42441b79, 32'h41505685, 32'h41f1fbbf, 32'h0, 32'h421289d5};
test_input[22704:22711] = '{32'h42100e75, 32'h427eeabb, 32'h429efd64, 32'h3fcb8e96, 32'hc2be0030, 32'h4211edc9, 32'hc2967b9d, 32'hc1085fe7};
test_output[22704:22711] = '{32'h42100e75, 32'h427eeabb, 32'h429efd64, 32'h3fcb8e96, 32'h0, 32'h4211edc9, 32'h0, 32'h0};
test_input[22712:22719] = '{32'h42195636, 32'h4280fb04, 32'h41e0bb3a, 32'hc1e66c68, 32'h427a5b41, 32'hc2688ded, 32'hc2285362, 32'hc20312e3};
test_output[22712:22719] = '{32'h42195636, 32'h4280fb04, 32'h41e0bb3a, 32'h0, 32'h427a5b41, 32'h0, 32'h0, 32'h0};
test_input[22720:22727] = '{32'hc2b3d0f7, 32'hc26072ea, 32'hc2c0e619, 32'hc187de73, 32'h40ac24b3, 32'h41eb6db3, 32'h4290a6f3, 32'h40d39a2b};
test_output[22720:22727] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40ac24b3, 32'h41eb6db3, 32'h4290a6f3, 32'h40d39a2b};
test_input[22728:22735] = '{32'hc2904f3c, 32'hc239f1be, 32'h421d0921, 32'h41639f7f, 32'h429e0d56, 32'h42a1351a, 32'hc1605a9a, 32'hc1f5ac4e};
test_output[22728:22735] = '{32'h0, 32'h0, 32'h421d0921, 32'h41639f7f, 32'h429e0d56, 32'h42a1351a, 32'h0, 32'h0};
test_input[22736:22743] = '{32'hc1b7d93d, 32'h42a0d3f1, 32'hc0b06d90, 32'h42a217ec, 32'hc1d6db8d, 32'h423d0d53, 32'hc28266cf, 32'hc22d04c5};
test_output[22736:22743] = '{32'h0, 32'h42a0d3f1, 32'h0, 32'h42a217ec, 32'h0, 32'h423d0d53, 32'h0, 32'h0};
test_input[22744:22751] = '{32'hc26cf0f1, 32'h42b63c37, 32'h422126e8, 32'hc2356c7c, 32'h41086edb, 32'h428ec71e, 32'hc23c1a08, 32'hc23e3479};
test_output[22744:22751] = '{32'h0, 32'h42b63c37, 32'h422126e8, 32'h0, 32'h41086edb, 32'h428ec71e, 32'h0, 32'h0};
test_input[22752:22759] = '{32'hc1b1e9eb, 32'hc1ecfb2b, 32'hc279b6d1, 32'hc2171bd2, 32'h411e9c6e, 32'h425e6036, 32'hc2734449, 32'h41853ba1};
test_output[22752:22759] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h411e9c6e, 32'h425e6036, 32'h0, 32'h41853ba1};
test_input[22760:22767] = '{32'hc28dacbc, 32'h425c977f, 32'hc272e6f2, 32'h428bb2d4, 32'h42900755, 32'hc2398fb6, 32'hc2378dfb, 32'hc2c5534c};
test_output[22760:22767] = '{32'h0, 32'h425c977f, 32'h0, 32'h428bb2d4, 32'h42900755, 32'h0, 32'h0, 32'h0};
test_input[22768:22775] = '{32'hc140b9e6, 32'hc29f19c2, 32'hc249362b, 32'h41bc6736, 32'h42a95638, 32'h42b17c8b, 32'hc29d6d49, 32'hc28f3f8b};
test_output[22768:22775] = '{32'h0, 32'h0, 32'h0, 32'h41bc6736, 32'h42a95638, 32'h42b17c8b, 32'h0, 32'h0};
test_input[22776:22783] = '{32'hc2acdf2c, 32'hc214e718, 32'hc1407115, 32'h4209e219, 32'h412af706, 32'h409b6bee, 32'h4251f77c, 32'hc21d3184};
test_output[22776:22783] = '{32'h0, 32'h0, 32'h0, 32'h4209e219, 32'h412af706, 32'h409b6bee, 32'h4251f77c, 32'h0};
test_input[22784:22791] = '{32'h41b18bf6, 32'h428d4939, 32'hc29fab95, 32'hc13b482f, 32'hc09fc4df, 32'hc233dfd6, 32'h41aad38a, 32'h4246785a};
test_output[22784:22791] = '{32'h41b18bf6, 32'h428d4939, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41aad38a, 32'h4246785a};
test_input[22792:22799] = '{32'hc2c4740d, 32'h4282c61e, 32'h42413448, 32'hc23d4033, 32'hc0057f62, 32'h42b169c1, 32'h4204dd24, 32'hc01f46cd};
test_output[22792:22799] = '{32'h0, 32'h4282c61e, 32'h42413448, 32'h0, 32'h0, 32'h42b169c1, 32'h4204dd24, 32'h0};
test_input[22800:22807] = '{32'h4249ad22, 32'hc28550a4, 32'hc294adcb, 32'hc2b837a7, 32'h428bb3a6, 32'h429205d8, 32'h4160e93c, 32'hc2a0bce5};
test_output[22800:22807] = '{32'h4249ad22, 32'h0, 32'h0, 32'h0, 32'h428bb3a6, 32'h429205d8, 32'h4160e93c, 32'h0};
test_input[22808:22815] = '{32'h41d876e1, 32'hc2a07718, 32'h4194c499, 32'h411a2b5f, 32'h4221db48, 32'hc1e76d1e, 32'hc207e8a4, 32'hc2b4cce4};
test_output[22808:22815] = '{32'h41d876e1, 32'h0, 32'h4194c499, 32'h411a2b5f, 32'h4221db48, 32'h0, 32'h0, 32'h0};
test_input[22816:22823] = '{32'h4207ab32, 32'hc2a64029, 32'h42a95560, 32'hc244819d, 32'hc1ec3359, 32'hc2513814, 32'hc1319a75, 32'hc158aa29};
test_output[22816:22823] = '{32'h4207ab32, 32'h0, 32'h42a95560, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22824:22831] = '{32'h42b5d856, 32'hc29da621, 32'h403bbd7d, 32'h428463ef, 32'h40f7da7e, 32'hc28181a0, 32'hc25e3cbc, 32'hc21d70f2};
test_output[22824:22831] = '{32'h42b5d856, 32'h0, 32'h403bbd7d, 32'h428463ef, 32'h40f7da7e, 32'h0, 32'h0, 32'h0};
test_input[22832:22839] = '{32'h41ca0c40, 32'h41718d60, 32'h418aa502, 32'h42a5d8e2, 32'h41ced251, 32'hc24a3ba7, 32'h429341f4, 32'h420d35ae};
test_output[22832:22839] = '{32'h41ca0c40, 32'h41718d60, 32'h418aa502, 32'h42a5d8e2, 32'h41ced251, 32'h0, 32'h429341f4, 32'h420d35ae};
test_input[22840:22847] = '{32'hc223fef0, 32'h4220e947, 32'hc1d2f838, 32'h4171ef6c, 32'hc20095cb, 32'hc2757977, 32'h41c6d419, 32'h4116ca86};
test_output[22840:22847] = '{32'h0, 32'h4220e947, 32'h0, 32'h4171ef6c, 32'h0, 32'h0, 32'h41c6d419, 32'h4116ca86};
test_input[22848:22855] = '{32'h4186bd66, 32'hc2a239bb, 32'h41b34909, 32'hc280204d, 32'hc2632bec, 32'hc0f9120a, 32'hc1310536, 32'hc2b92735};
test_output[22848:22855] = '{32'h4186bd66, 32'h0, 32'h41b34909, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22856:22863] = '{32'hc2249e80, 32'hc1e7d7be, 32'hc27b8bec, 32'h42bc00ce, 32'h42c0b07a, 32'hc1488285, 32'h4296b630, 32'hc1c135b4};
test_output[22856:22863] = '{32'h0, 32'h0, 32'h0, 32'h42bc00ce, 32'h42c0b07a, 32'h0, 32'h4296b630, 32'h0};
test_input[22864:22871] = '{32'hc164ef38, 32'hc27e50db, 32'h42c64ccb, 32'hc28c2c10, 32'h4224aac7, 32'hc1965f92, 32'hc2a80309, 32'h40e75c90};
test_output[22864:22871] = '{32'h0, 32'h0, 32'h42c64ccb, 32'h0, 32'h4224aac7, 32'h0, 32'h0, 32'h40e75c90};
test_input[22872:22879] = '{32'hc1b3c31c, 32'h42b67a34, 32'hc26ce047, 32'h4262ac1b, 32'hc0e3488e, 32'hc2514928, 32'hc23ef9ec, 32'h424c37d5};
test_output[22872:22879] = '{32'h0, 32'h42b67a34, 32'h0, 32'h4262ac1b, 32'h0, 32'h0, 32'h0, 32'h424c37d5};
test_input[22880:22887] = '{32'hc29f9dbc, 32'h41dfab68, 32'h422374e2, 32'hc21ea7a0, 32'hc26fb038, 32'hc25e9d07, 32'h41003825, 32'hc271aa57};
test_output[22880:22887] = '{32'h0, 32'h41dfab68, 32'h422374e2, 32'h0, 32'h0, 32'h0, 32'h41003825, 32'h0};
test_input[22888:22895] = '{32'h422f1c1b, 32'hc295d11e, 32'h42b68257, 32'hc24c45b9, 32'hc1c033e4, 32'hc09bfab3, 32'hbff0f164, 32'h422ed7e7};
test_output[22888:22895] = '{32'h422f1c1b, 32'h0, 32'h42b68257, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422ed7e7};
test_input[22896:22903] = '{32'h41ae27b3, 32'h42552a4d, 32'h419075e3, 32'hc1ead479, 32'hc14e959f, 32'h42555906, 32'hc291f645, 32'h421c69ac};
test_output[22896:22903] = '{32'h41ae27b3, 32'h42552a4d, 32'h419075e3, 32'h0, 32'h0, 32'h42555906, 32'h0, 32'h421c69ac};
test_input[22904:22911] = '{32'hc22d2cbc, 32'h42907a20, 32'hc2c01e18, 32'hc28267c9, 32'hc1ccf4ab, 32'h42bfab39, 32'hc253ed2e, 32'h41f68578};
test_output[22904:22911] = '{32'h0, 32'h42907a20, 32'h0, 32'h0, 32'h0, 32'h42bfab39, 32'h0, 32'h41f68578};
test_input[22912:22919] = '{32'hc28db91d, 32'hc21a5184, 32'h3f835090, 32'hc271342e, 32'hc2766add, 32'hc29283df, 32'h426104e4, 32'hc20f0281};
test_output[22912:22919] = '{32'h0, 32'h0, 32'h3f835090, 32'h0, 32'h0, 32'h0, 32'h426104e4, 32'h0};
test_input[22920:22927] = '{32'h422223be, 32'hc1855262, 32'h42a44bc7, 32'h4237cbca, 32'hc29fcf3e, 32'h42306188, 32'hc28209b4, 32'h42a72a0b};
test_output[22920:22927] = '{32'h422223be, 32'h0, 32'h42a44bc7, 32'h4237cbca, 32'h0, 32'h42306188, 32'h0, 32'h42a72a0b};
test_input[22928:22935] = '{32'hc26ee4f1, 32'h4200de49, 32'h427f1b62, 32'hc243b9ac, 32'hc2b61e45, 32'hc17186b3, 32'h4092165d, 32'hc2ab06c1};
test_output[22928:22935] = '{32'h0, 32'h4200de49, 32'h427f1b62, 32'h0, 32'h0, 32'h0, 32'h4092165d, 32'h0};
test_input[22936:22943] = '{32'h427860dc, 32'h428ece22, 32'h42b2e585, 32'hc0c2e7e4, 32'h428b758d, 32'hc26bf6e5, 32'hc093c49c, 32'hc2706f35};
test_output[22936:22943] = '{32'h427860dc, 32'h428ece22, 32'h42b2e585, 32'h0, 32'h428b758d, 32'h0, 32'h0, 32'h0};
test_input[22944:22951] = '{32'h425cb035, 32'hc2a093a4, 32'h41960dbf, 32'h42b533fc, 32'hc27021ad, 32'h420f2aa0, 32'h42086d55, 32'h4261cd87};
test_output[22944:22951] = '{32'h425cb035, 32'h0, 32'h41960dbf, 32'h42b533fc, 32'h0, 32'h420f2aa0, 32'h42086d55, 32'h4261cd87};
test_input[22952:22959] = '{32'h41bf2099, 32'h424814a0, 32'h41f78e79, 32'h42a44ac0, 32'h421c369c, 32'hc1d0016c, 32'hc22f0931, 32'hc2955b92};
test_output[22952:22959] = '{32'h41bf2099, 32'h424814a0, 32'h41f78e79, 32'h42a44ac0, 32'h421c369c, 32'h0, 32'h0, 32'h0};
test_input[22960:22967] = '{32'h40e0b9c9, 32'hc1b3bfab, 32'h421b4b8d, 32'hc2a40e91, 32'h423da296, 32'h41b75e36, 32'h42b13703, 32'h42ae5994};
test_output[22960:22967] = '{32'h40e0b9c9, 32'h0, 32'h421b4b8d, 32'h0, 32'h423da296, 32'h41b75e36, 32'h42b13703, 32'h42ae5994};
test_input[22968:22975] = '{32'hc186d159, 32'hc2a09d97, 32'h426f589d, 32'hc1248f4e, 32'hc22b1564, 32'hc20a0bbc, 32'hc1bb86cb, 32'h41560a64};
test_output[22968:22975] = '{32'h0, 32'h0, 32'h426f589d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41560a64};
test_input[22976:22983] = '{32'hc1a2b467, 32'h42781319, 32'h41aeb7a8, 32'h41f0339c, 32'hc2444677, 32'h4075be26, 32'h42662ff3, 32'h42c12834};
test_output[22976:22983] = '{32'h0, 32'h42781319, 32'h41aeb7a8, 32'h41f0339c, 32'h0, 32'h4075be26, 32'h42662ff3, 32'h42c12834};
test_input[22984:22991] = '{32'h424220ef, 32'h427d3fdd, 32'hc275422f, 32'hc2a53980, 32'hc2194e46, 32'hbffb384a, 32'h4227ab25, 32'hc29bd919};
test_output[22984:22991] = '{32'h424220ef, 32'h427d3fdd, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4227ab25, 32'h0};
test_input[22992:22999] = '{32'h42b72c21, 32'hc0b3c91b, 32'hc2b59dde, 32'hc1cbbad2, 32'h4164a5da, 32'h40d3f5b8, 32'hc283cf72, 32'h4255c533};
test_output[22992:22999] = '{32'h42b72c21, 32'h0, 32'h0, 32'h0, 32'h4164a5da, 32'h40d3f5b8, 32'h0, 32'h4255c533};
test_input[23000:23007] = '{32'hc2441ccb, 32'h40803cb5, 32'h429e5a13, 32'h4299fff5, 32'h422d1d2a, 32'h42aa79be, 32'hc1271113, 32'h41c9e24e};
test_output[23000:23007] = '{32'h0, 32'h40803cb5, 32'h429e5a13, 32'h4299fff5, 32'h422d1d2a, 32'h42aa79be, 32'h0, 32'h41c9e24e};
test_input[23008:23015] = '{32'hc268c25b, 32'h426925ac, 32'h429b63aa, 32'h4220740d, 32'hc21a4063, 32'hc298618e, 32'hc23d3cbc, 32'hc21e8da0};
test_output[23008:23015] = '{32'h0, 32'h426925ac, 32'h429b63aa, 32'h4220740d, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23016:23023] = '{32'h4212260f, 32'h42834aae, 32'h42007662, 32'hc2062c1f, 32'h429de29f, 32'h424e5efd, 32'hc2a4a60f, 32'hc21f52e2};
test_output[23016:23023] = '{32'h4212260f, 32'h42834aae, 32'h42007662, 32'h0, 32'h429de29f, 32'h424e5efd, 32'h0, 32'h0};
test_input[23024:23031] = '{32'h429a6011, 32'h40d2277f, 32'h42bda0fb, 32'hc2c0b5b1, 32'h428849b9, 32'hc28eccd1, 32'hc28b0b58, 32'hc25a241b};
test_output[23024:23031] = '{32'h429a6011, 32'h40d2277f, 32'h42bda0fb, 32'h0, 32'h428849b9, 32'h0, 32'h0, 32'h0};
test_input[23032:23039] = '{32'h41db8c26, 32'h407b1979, 32'h4205a883, 32'h4241ac2f, 32'hc275643d, 32'hc2bb18a6, 32'hc27e7486, 32'h42877581};
test_output[23032:23039] = '{32'h41db8c26, 32'h407b1979, 32'h4205a883, 32'h4241ac2f, 32'h0, 32'h0, 32'h0, 32'h42877581};
test_input[23040:23047] = '{32'h4296002f, 32'hc20f06de, 32'h41d1261c, 32'h42c4a788, 32'h40d10963, 32'hc27ff257, 32'hc1ae7cb7, 32'h42420281};
test_output[23040:23047] = '{32'h4296002f, 32'h0, 32'h41d1261c, 32'h42c4a788, 32'h40d10963, 32'h0, 32'h0, 32'h42420281};
test_input[23048:23055] = '{32'h42377907, 32'h42451d84, 32'hc1fb1cb6, 32'h427fd330, 32'h4284a4a0, 32'hc2854c0d, 32'hc29e9253, 32'hc2aa9432};
test_output[23048:23055] = '{32'h42377907, 32'h42451d84, 32'h0, 32'h427fd330, 32'h4284a4a0, 32'h0, 32'h0, 32'h0};
test_input[23056:23063] = '{32'h42c38716, 32'hc07058c2, 32'h41bd91c9, 32'h424e1475, 32'h40d577c7, 32'hc1d3805f, 32'hc015c414, 32'hc2bc2a1e};
test_output[23056:23063] = '{32'h42c38716, 32'h0, 32'h41bd91c9, 32'h424e1475, 32'h40d577c7, 32'h0, 32'h0, 32'h0};
test_input[23064:23071] = '{32'h41237a84, 32'hc220e29e, 32'hc231e7b7, 32'hc1b01e9d, 32'h4204d2bb, 32'hc181d6a0, 32'hc26c0210, 32'hc293637f};
test_output[23064:23071] = '{32'h41237a84, 32'h0, 32'h0, 32'h0, 32'h4204d2bb, 32'h0, 32'h0, 32'h0};
test_input[23072:23079] = '{32'hc256cf76, 32'h4130297e, 32'h4280a675, 32'hc14f7076, 32'h4282fbee, 32'hc18db17f, 32'hc2483762, 32'hc1d2669b};
test_output[23072:23079] = '{32'h0, 32'h4130297e, 32'h4280a675, 32'h0, 32'h4282fbee, 32'h0, 32'h0, 32'h0};
test_input[23080:23087] = '{32'h4291e28b, 32'h41e33ac7, 32'hc09debbf, 32'hc29939e8, 32'hc2b966d8, 32'hc2792afa, 32'hc2ba06b7, 32'hc0e9987c};
test_output[23080:23087] = '{32'h4291e28b, 32'h41e33ac7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23088:23095] = '{32'hc2a0bbc2, 32'h428938a2, 32'h424839f1, 32'hc1b0d11f, 32'hc224d0ed, 32'hc229c409, 32'h42aa6ccc, 32'h424f776f};
test_output[23088:23095] = '{32'h0, 32'h428938a2, 32'h424839f1, 32'h0, 32'h0, 32'h0, 32'h42aa6ccc, 32'h424f776f};
test_input[23096:23103] = '{32'hc2457f22, 32'hc266b17b, 32'h422eee2c, 32'h4233f930, 32'h42377e13, 32'hc2160bb7, 32'h42c45c23, 32'h42008c10};
test_output[23096:23103] = '{32'h0, 32'h0, 32'h422eee2c, 32'h4233f930, 32'h42377e13, 32'h0, 32'h42c45c23, 32'h42008c10};
test_input[23104:23111] = '{32'h4184d835, 32'hc200d8b7, 32'hc2b23199, 32'h42705b7a, 32'h41e5c5c6, 32'hc0c3844f, 32'hc0f80912, 32'h42b75173};
test_output[23104:23111] = '{32'h4184d835, 32'h0, 32'h0, 32'h42705b7a, 32'h41e5c5c6, 32'h0, 32'h0, 32'h42b75173};
test_input[23112:23119] = '{32'h42b0ec4f, 32'h42b02514, 32'hc0f3887c, 32'h42345b8e, 32'hc020b9f7, 32'h42145e53, 32'hc226db17, 32'hc29938a8};
test_output[23112:23119] = '{32'h42b0ec4f, 32'h42b02514, 32'h0, 32'h42345b8e, 32'h0, 32'h42145e53, 32'h0, 32'h0};
test_input[23120:23127] = '{32'h41c5ff5a, 32'hc235153e, 32'h428a4e7a, 32'hc1c51f70, 32'hc2ade6d2, 32'hc187c809, 32'h42c29d92, 32'h425de4ff};
test_output[23120:23127] = '{32'h41c5ff5a, 32'h0, 32'h428a4e7a, 32'h0, 32'h0, 32'h0, 32'h42c29d92, 32'h425de4ff};
test_input[23128:23135] = '{32'h41daceca, 32'h42bf85d5, 32'h420f8cbb, 32'h419ab316, 32'hc28a5af6, 32'hc2af7f0f, 32'hc20ae360, 32'h41d38afe};
test_output[23128:23135] = '{32'h41daceca, 32'h42bf85d5, 32'h420f8cbb, 32'h419ab316, 32'h0, 32'h0, 32'h0, 32'h41d38afe};
test_input[23136:23143] = '{32'hc1e4f7c2, 32'hc28f7a32, 32'h427dd5da, 32'hc27be06b, 32'hc1d8e1e4, 32'h41f1bc22, 32'h42b69538, 32'h4293eadf};
test_output[23136:23143] = '{32'h0, 32'h0, 32'h427dd5da, 32'h0, 32'h0, 32'h41f1bc22, 32'h42b69538, 32'h4293eadf};
test_input[23144:23151] = '{32'hc234fc4e, 32'h41fd61d5, 32'hc233c4ea, 32'h41d2ce3d, 32'h425548de, 32'hc2050659, 32'h41acef0a, 32'hc1f60c6d};
test_output[23144:23151] = '{32'h0, 32'h41fd61d5, 32'h0, 32'h41d2ce3d, 32'h425548de, 32'h0, 32'h41acef0a, 32'h0};
test_input[23152:23159] = '{32'h4293fcce, 32'hc20b3128, 32'h41a3910e, 32'h423313fa, 32'hc2840ebd, 32'h41c5ee27, 32'hc2a33215, 32'hc095f516};
test_output[23152:23159] = '{32'h4293fcce, 32'h0, 32'h41a3910e, 32'h423313fa, 32'h0, 32'h41c5ee27, 32'h0, 32'h0};
test_input[23160:23167] = '{32'h42a51d7b, 32'h418aabc0, 32'hc2b64546, 32'h4120af05, 32'h41ab9c67, 32'hc2c273ed, 32'hc24c1323, 32'hc2acd3e0};
test_output[23160:23167] = '{32'h42a51d7b, 32'h418aabc0, 32'h0, 32'h4120af05, 32'h41ab9c67, 32'h0, 32'h0, 32'h0};
test_input[23168:23175] = '{32'hc2a9b208, 32'h42b5c1a7, 32'h41c63b91, 32'h42692be7, 32'hc216e464, 32'h42b97c53, 32'h42563cf2, 32'hc2a8e236};
test_output[23168:23175] = '{32'h0, 32'h42b5c1a7, 32'h41c63b91, 32'h42692be7, 32'h0, 32'h42b97c53, 32'h42563cf2, 32'h0};
test_input[23176:23183] = '{32'hc2831f4a, 32'hc21ee6cb, 32'h428190cf, 32'hc26e871c, 32'hc05cb190, 32'h4237dbed, 32'h422bb717, 32'hc208e0ae};
test_output[23176:23183] = '{32'h0, 32'h0, 32'h428190cf, 32'h0, 32'h0, 32'h4237dbed, 32'h422bb717, 32'h0};
test_input[23184:23191] = '{32'h41da0068, 32'hc2c1c977, 32'h41cd5dee, 32'h41c29f43, 32'hc2b10663, 32'h42065a7f, 32'h4239be91, 32'h429c3e44};
test_output[23184:23191] = '{32'h41da0068, 32'h0, 32'h41cd5dee, 32'h41c29f43, 32'h0, 32'h42065a7f, 32'h4239be91, 32'h429c3e44};
test_input[23192:23199] = '{32'h4271ffd1, 32'h42c63701, 32'h4199d323, 32'hc2724d15, 32'hc1360915, 32'h421845ee, 32'hc28e2abe, 32'h426e6816};
test_output[23192:23199] = '{32'h4271ffd1, 32'h42c63701, 32'h4199d323, 32'h0, 32'h0, 32'h421845ee, 32'h0, 32'h426e6816};
test_input[23200:23207] = '{32'hc234c58a, 32'h42718595, 32'h4239d54d, 32'h42626a42, 32'h4290584b, 32'h425d6c61, 32'h40c91b76, 32'h41a97e25};
test_output[23200:23207] = '{32'h0, 32'h42718595, 32'h4239d54d, 32'h42626a42, 32'h4290584b, 32'h425d6c61, 32'h40c91b76, 32'h41a97e25};
test_input[23208:23215] = '{32'h4201572c, 32'h42729f0c, 32'hc14d7a8e, 32'h428f453e, 32'hc1ecd46d, 32'h3e689a7d, 32'hbebd2f17, 32'hc2915957};
test_output[23208:23215] = '{32'h4201572c, 32'h42729f0c, 32'h0, 32'h428f453e, 32'h0, 32'h3e689a7d, 32'h0, 32'h0};
test_input[23216:23223] = '{32'hc2907897, 32'h42852111, 32'hc2bc3eb6, 32'h42bc3a69, 32'h4233512d, 32'h4258c075, 32'hc212f90b, 32'hc2ae901e};
test_output[23216:23223] = '{32'h0, 32'h42852111, 32'h0, 32'h42bc3a69, 32'h4233512d, 32'h4258c075, 32'h0, 32'h0};
test_input[23224:23231] = '{32'hc12376ee, 32'h410dff09, 32'hc249f3db, 32'h42c34c20, 32'h4249936d, 32'h428664e8, 32'hc0a59d0a, 32'hc225b665};
test_output[23224:23231] = '{32'h0, 32'h410dff09, 32'h0, 32'h42c34c20, 32'h4249936d, 32'h428664e8, 32'h0, 32'h0};
test_input[23232:23239] = '{32'h42c7e411, 32'hc2c7686b, 32'h40d4c3a1, 32'h428ccda0, 32'h41b5f864, 32'hc2bbb814, 32'hc1e20ef8, 32'hc282c8d4};
test_output[23232:23239] = '{32'h42c7e411, 32'h0, 32'h40d4c3a1, 32'h428ccda0, 32'h41b5f864, 32'h0, 32'h0, 32'h0};
test_input[23240:23247] = '{32'h41ff247f, 32'hc1955aa2, 32'hc272763c, 32'h4291589c, 32'h42739d1e, 32'hc1e0fb01, 32'hc2b3436c, 32'h41a3492f};
test_output[23240:23247] = '{32'h41ff247f, 32'h0, 32'h0, 32'h4291589c, 32'h42739d1e, 32'h0, 32'h0, 32'h41a3492f};
test_input[23248:23255] = '{32'h40c2c67c, 32'h41e31c2d, 32'h4146698f, 32'h42aea9da, 32'h4268ec58, 32'hc2b56363, 32'hc11c3faa, 32'h40c50b80};
test_output[23248:23255] = '{32'h40c2c67c, 32'h41e31c2d, 32'h4146698f, 32'h42aea9da, 32'h4268ec58, 32'h0, 32'h0, 32'h40c50b80};
test_input[23256:23263] = '{32'hc18a6da9, 32'hc23c55fc, 32'hc2560eea, 32'h4293da67, 32'h424460cb, 32'hc2a8024d, 32'hc25c6471, 32'h41db40ee};
test_output[23256:23263] = '{32'h0, 32'h0, 32'h0, 32'h4293da67, 32'h424460cb, 32'h0, 32'h0, 32'h41db40ee};
test_input[23264:23271] = '{32'h42c58470, 32'h42aae88e, 32'hc113a9c5, 32'h422cf73e, 32'hc0831dd7, 32'hc2b8c46e, 32'hc2aa0fb6, 32'hc29ed067};
test_output[23264:23271] = '{32'h42c58470, 32'h42aae88e, 32'h0, 32'h422cf73e, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23272:23279] = '{32'h42a959b0, 32'h418e9e3e, 32'h42999b53, 32'h424eeec8, 32'h41e76fbb, 32'hc2b2827b, 32'hc222a40a, 32'hc22f7702};
test_output[23272:23279] = '{32'h42a959b0, 32'h418e9e3e, 32'h42999b53, 32'h424eeec8, 32'h41e76fbb, 32'h0, 32'h0, 32'h0};
test_input[23280:23287] = '{32'h41d95bf5, 32'h42bf8330, 32'h3f797a0a, 32'h42266306, 32'h420bf4a5, 32'h42350787, 32'hc1bac60b, 32'hc24affc8};
test_output[23280:23287] = '{32'h41d95bf5, 32'h42bf8330, 32'h3f797a0a, 32'h42266306, 32'h420bf4a5, 32'h42350787, 32'h0, 32'h0};
test_input[23288:23295] = '{32'h418086e3, 32'h4213c275, 32'h42896fc8, 32'hc2c69360, 32'hc21643df, 32'h42b3453c, 32'h42559a75, 32'hc1dd747a};
test_output[23288:23295] = '{32'h418086e3, 32'h4213c275, 32'h42896fc8, 32'h0, 32'h0, 32'h42b3453c, 32'h42559a75, 32'h0};
test_input[23296:23303] = '{32'hc19bc151, 32'h423ee6a9, 32'hc2c28027, 32'hc228b895, 32'h4288a505, 32'h42702023, 32'hc27390ad, 32'h42c5dca5};
test_output[23296:23303] = '{32'h0, 32'h423ee6a9, 32'h0, 32'h0, 32'h4288a505, 32'h42702023, 32'h0, 32'h42c5dca5};
test_input[23304:23311] = '{32'h41fd16f9, 32'hc0ff8485, 32'hc2c49730, 32'hc205a054, 32'h4132a954, 32'hc2aa01cf, 32'h424e2c94, 32'h427891d9};
test_output[23304:23311] = '{32'h41fd16f9, 32'h0, 32'h0, 32'h0, 32'h4132a954, 32'h0, 32'h424e2c94, 32'h427891d9};
test_input[23312:23319] = '{32'h4287c56f, 32'hc1c907ac, 32'h41696fb1, 32'h41a7338b, 32'h40d1fa86, 32'hc215d77b, 32'hc11243aa, 32'hc2c4bca6};
test_output[23312:23319] = '{32'h4287c56f, 32'h0, 32'h41696fb1, 32'h41a7338b, 32'h40d1fa86, 32'h0, 32'h0, 32'h0};
test_input[23320:23327] = '{32'h41d7f3ce, 32'hc223dcb5, 32'h4176ade2, 32'hc11ea8ca, 32'h3ff59c7d, 32'hc25d6102, 32'hc1f8618d, 32'h42579bd1};
test_output[23320:23327] = '{32'h41d7f3ce, 32'h0, 32'h4176ade2, 32'h0, 32'h3ff59c7d, 32'h0, 32'h0, 32'h42579bd1};
test_input[23328:23335] = '{32'h421e64b7, 32'hc25624e0, 32'hc21b495b, 32'hc28b3a61, 32'h42a8035e, 32'hc2c60554, 32'hc2c2db37, 32'hc0588b70};
test_output[23328:23335] = '{32'h421e64b7, 32'h0, 32'h0, 32'h0, 32'h42a8035e, 32'h0, 32'h0, 32'h0};
test_input[23336:23343] = '{32'hc179902a, 32'hc2af7179, 32'hc2885126, 32'h4289145a, 32'h42a9b9aa, 32'h4249f6bf, 32'h41fe5876, 32'h422b78ef};
test_output[23336:23343] = '{32'h0, 32'h0, 32'h0, 32'h4289145a, 32'h42a9b9aa, 32'h4249f6bf, 32'h41fe5876, 32'h422b78ef};
test_input[23344:23351] = '{32'hc1ee0d0e, 32'h41ded410, 32'hc2470365, 32'hc1a8e78c, 32'h429fe118, 32'hc26d3380, 32'h42b5d2ac, 32'h41a47ac6};
test_output[23344:23351] = '{32'h0, 32'h41ded410, 32'h0, 32'h0, 32'h429fe118, 32'h0, 32'h42b5d2ac, 32'h41a47ac6};
test_input[23352:23359] = '{32'hc2b1e89b, 32'hc19b494e, 32'hc23e9efa, 32'h405dfef3, 32'h42515db3, 32'h3fbd9568, 32'h41794f84, 32'hc2a52459};
test_output[23352:23359] = '{32'h0, 32'h0, 32'h0, 32'h405dfef3, 32'h42515db3, 32'h3fbd9568, 32'h41794f84, 32'h0};
test_input[23360:23367] = '{32'hc1a154c7, 32'hc1d294c8, 32'hc1877e81, 32'h402a9e4f, 32'h42540e45, 32'h428cce01, 32'hc1fefad3, 32'hc29e6a96};
test_output[23360:23367] = '{32'h0, 32'h0, 32'h0, 32'h402a9e4f, 32'h42540e45, 32'h428cce01, 32'h0, 32'h0};
test_input[23368:23375] = '{32'hc14207cf, 32'h427ae509, 32'hc28776ba, 32'hc2079fa7, 32'h429e2bb0, 32'h4207aadb, 32'hc2af1ee6, 32'hc2476903};
test_output[23368:23375] = '{32'h0, 32'h427ae509, 32'h0, 32'h0, 32'h429e2bb0, 32'h4207aadb, 32'h0, 32'h0};
test_input[23376:23383] = '{32'hc1abb2b0, 32'h428e1703, 32'hc1e6583b, 32'hc2817fb5, 32'hc2b01b3d, 32'hc23e0df9, 32'hc2afb15f, 32'hc1b8b985};
test_output[23376:23383] = '{32'h0, 32'h428e1703, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23384:23391] = '{32'h41bc4cb4, 32'hc27e92d8, 32'h425eee82, 32'h422ce870, 32'hc229a522, 32'h427daafa, 32'hc2c4ac78, 32'h42bb8920};
test_output[23384:23391] = '{32'h41bc4cb4, 32'h0, 32'h425eee82, 32'h422ce870, 32'h0, 32'h427daafa, 32'h0, 32'h42bb8920};
test_input[23392:23399] = '{32'h428afd4d, 32'hc0450547, 32'h4235ea1c, 32'hc2b7c8b3, 32'h41873d28, 32'hc204564e, 32'h413a0db0, 32'hc241532c};
test_output[23392:23399] = '{32'h428afd4d, 32'h0, 32'h4235ea1c, 32'h0, 32'h41873d28, 32'h0, 32'h413a0db0, 32'h0};
test_input[23400:23407] = '{32'h3e445f32, 32'hc2b7b105, 32'hc1853cd3, 32'hc2412fbd, 32'hc2c2c2bb, 32'hc2a1f6a3, 32'hbf2222c9, 32'h42574493};
test_output[23400:23407] = '{32'h3e445f32, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42574493};
test_input[23408:23415] = '{32'hc22882d2, 32'hc21af2ac, 32'hc2a128b8, 32'hc2246840, 32'hc2c79d68, 32'h4231159d, 32'hc21de09b, 32'hc2c4318f};
test_output[23408:23415] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4231159d, 32'h0, 32'h0};
test_input[23416:23423] = '{32'hc29c24af, 32'h4292f629, 32'h427c3e7b, 32'hc2a9366c, 32'hc2572c7e, 32'h40fb0b8b, 32'h3fd82a39, 32'h41d97056};
test_output[23416:23423] = '{32'h0, 32'h4292f629, 32'h427c3e7b, 32'h0, 32'h0, 32'h40fb0b8b, 32'h3fd82a39, 32'h41d97056};
test_input[23424:23431] = '{32'h41eda175, 32'h4261e1ac, 32'h428a84e0, 32'hc2734e61, 32'h42a6a916, 32'h42bd630c, 32'hc2ac071c, 32'h428bf54b};
test_output[23424:23431] = '{32'h41eda175, 32'h4261e1ac, 32'h428a84e0, 32'h0, 32'h42a6a916, 32'h42bd630c, 32'h0, 32'h428bf54b};
test_input[23432:23439] = '{32'h429b3e3c, 32'hc2a9a013, 32'hc2961164, 32'h42b1f91d, 32'h41a1294a, 32'h42015dab, 32'hc2b8ccb9, 32'hc205ffd1};
test_output[23432:23439] = '{32'h429b3e3c, 32'h0, 32'h0, 32'h42b1f91d, 32'h41a1294a, 32'h42015dab, 32'h0, 32'h0};
test_input[23440:23447] = '{32'hc26ee95b, 32'hc2217d59, 32'h42b69dce, 32'hc1094063, 32'hbfbe258c, 32'hc2951641, 32'hc2a616a6, 32'hc27c1625};
test_output[23440:23447] = '{32'h0, 32'h0, 32'h42b69dce, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23448:23455] = '{32'hc2915e00, 32'h420ba545, 32'h4282bcd0, 32'h419d03e0, 32'hc2c45d59, 32'hc25cc9d1, 32'hc1ce40a3, 32'hc250f6fb};
test_output[23448:23455] = '{32'h0, 32'h420ba545, 32'h4282bcd0, 32'h419d03e0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23456:23463] = '{32'hc2b199ba, 32'h4282daf3, 32'hc297bcc1, 32'hc29cad8e, 32'h41ae86f8, 32'h4181a70d, 32'h42a9cd9e, 32'hc284d843};
test_output[23456:23463] = '{32'h0, 32'h4282daf3, 32'h0, 32'h0, 32'h41ae86f8, 32'h4181a70d, 32'h42a9cd9e, 32'h0};
test_input[23464:23471] = '{32'hc201f0e9, 32'h42a58f74, 32'h418087c9, 32'hc1adee53, 32'h426cbba5, 32'h4224f661, 32'hc21bb90a, 32'h42942ac9};
test_output[23464:23471] = '{32'h0, 32'h42a58f74, 32'h418087c9, 32'h0, 32'h426cbba5, 32'h4224f661, 32'h0, 32'h42942ac9};
test_input[23472:23479] = '{32'hc1f839f0, 32'hc2b4d14e, 32'h42bc6436, 32'hc2a9ecff, 32'hc2be6714, 32'h42a4beca, 32'h42b2e1a3, 32'hc1a69bec};
test_output[23472:23479] = '{32'h0, 32'h0, 32'h42bc6436, 32'h0, 32'h0, 32'h42a4beca, 32'h42b2e1a3, 32'h0};
test_input[23480:23487] = '{32'hc138f6f0, 32'hc26120b4, 32'hc2787b98, 32'hc1228d9e, 32'hc24ec5d7, 32'hc1d1c0e9, 32'hc2a43732, 32'hc2579a97};
test_output[23480:23487] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23488:23495] = '{32'h4211b1f0, 32'hc2b4067a, 32'hc16910b0, 32'h410da099, 32'h42ab1487, 32'h423e983d, 32'h4014e086, 32'hc20edb7c};
test_output[23488:23495] = '{32'h4211b1f0, 32'h0, 32'h0, 32'h410da099, 32'h42ab1487, 32'h423e983d, 32'h4014e086, 32'h0};
test_input[23496:23503] = '{32'hc2abc517, 32'hbee24ac3, 32'h4265ffa3, 32'h41ac6c20, 32'h40a8d839, 32'hc29c72c4, 32'h421a349d, 32'h428e193b};
test_output[23496:23503] = '{32'h0, 32'h0, 32'h4265ffa3, 32'h41ac6c20, 32'h40a8d839, 32'h0, 32'h421a349d, 32'h428e193b};
test_input[23504:23511] = '{32'hc2b768f4, 32'hc0ce464f, 32'h423dfbfe, 32'hc1fc5c05, 32'h4285e642, 32'h41265def, 32'hc2c7cdaf, 32'hc1faa5bb};
test_output[23504:23511] = '{32'h0, 32'h0, 32'h423dfbfe, 32'h0, 32'h4285e642, 32'h41265def, 32'h0, 32'h0};
test_input[23512:23519] = '{32'h425186df, 32'hc2713e73, 32'hc289b003, 32'h409949f5, 32'h428deed6, 32'hc1fd0150, 32'h42423a8e, 32'h4296257b};
test_output[23512:23519] = '{32'h425186df, 32'h0, 32'h0, 32'h409949f5, 32'h428deed6, 32'h0, 32'h42423a8e, 32'h4296257b};
test_input[23520:23527] = '{32'hc1e3c179, 32'h4293e6cc, 32'h424d1bff, 32'h42193341, 32'h425176b9, 32'h42c0d7b0, 32'hc28228f6, 32'h4251b7f0};
test_output[23520:23527] = '{32'h0, 32'h4293e6cc, 32'h424d1bff, 32'h42193341, 32'h425176b9, 32'h42c0d7b0, 32'h0, 32'h4251b7f0};
test_input[23528:23535] = '{32'hc2acd060, 32'hc2abda46, 32'hc19ceb32, 32'hc1478f96, 32'hc2b72e9a, 32'h41d5fde8, 32'h4290dc7a, 32'h41cdcd56};
test_output[23528:23535] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41d5fde8, 32'h4290dc7a, 32'h41cdcd56};
test_input[23536:23543] = '{32'h41421124, 32'h42177574, 32'h421877d1, 32'h428ac134, 32'hc22c1938, 32'h42996716, 32'h4288b6ca, 32'hc27735ca};
test_output[23536:23543] = '{32'h41421124, 32'h42177574, 32'h421877d1, 32'h428ac134, 32'h0, 32'h42996716, 32'h4288b6ca, 32'h0};
test_input[23544:23551] = '{32'h414f17de, 32'h42b6bfe8, 32'h42051402, 32'h42c184b6, 32'h424aba08, 32'hc20d4f4e, 32'h428dd332, 32'h420d538c};
test_output[23544:23551] = '{32'h414f17de, 32'h42b6bfe8, 32'h42051402, 32'h42c184b6, 32'h424aba08, 32'h0, 32'h428dd332, 32'h420d538c};
test_input[23552:23559] = '{32'hc1e35b02, 32'hc1467912, 32'hc285e720, 32'hc2b4ac91, 32'hbf7591a7, 32'h41c12952, 32'h42407111, 32'h42a546a0};
test_output[23552:23559] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41c12952, 32'h42407111, 32'h42a546a0};
test_input[23560:23567] = '{32'hc2728c0c, 32'hc1c1c056, 32'hc1f62c4b, 32'hc1aa654b, 32'hc0a4140a, 32'h41b1123d, 32'hc1238580, 32'h42012c81};
test_output[23560:23567] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b1123d, 32'h0, 32'h42012c81};
test_input[23568:23575] = '{32'hc259427d, 32'h41e098c4, 32'h426e8505, 32'h423192d9, 32'hc261d24d, 32'hc234b80e, 32'h42bdac98, 32'h42ac4ed0};
test_output[23568:23575] = '{32'h0, 32'h41e098c4, 32'h426e8505, 32'h423192d9, 32'h0, 32'h0, 32'h42bdac98, 32'h42ac4ed0};
test_input[23576:23583] = '{32'h41fe2e18, 32'h42bcddd1, 32'h40db5550, 32'h42987100, 32'h40b2b895, 32'h42c5111c, 32'hc244c69c, 32'h428234f8};
test_output[23576:23583] = '{32'h41fe2e18, 32'h42bcddd1, 32'h40db5550, 32'h42987100, 32'h40b2b895, 32'h42c5111c, 32'h0, 32'h428234f8};
test_input[23584:23591] = '{32'h41939705, 32'h4268b68a, 32'hc28162a3, 32'hc233ccb7, 32'hc244ea56, 32'hc1941cbf, 32'hc2232e81, 32'h422f4631};
test_output[23584:23591] = '{32'h41939705, 32'h4268b68a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422f4631};
test_input[23592:23599] = '{32'hc2262e42, 32'h42c2a095, 32'hc272456f, 32'h42c49377, 32'h42c1b1a0, 32'hc241348a, 32'h40def6a0, 32'h424207ec};
test_output[23592:23599] = '{32'h0, 32'h42c2a095, 32'h0, 32'h42c49377, 32'h42c1b1a0, 32'h0, 32'h40def6a0, 32'h424207ec};
test_input[23600:23607] = '{32'h42c4afb2, 32'h41684a5d, 32'hc16940bf, 32'h42b1f094, 32'h42b10043, 32'h4223e241, 32'hc117cd99, 32'h426dc43a};
test_output[23600:23607] = '{32'h42c4afb2, 32'h41684a5d, 32'h0, 32'h42b1f094, 32'h42b10043, 32'h4223e241, 32'h0, 32'h426dc43a};
test_input[23608:23615] = '{32'hc2658064, 32'h42a8ac18, 32'hc2a48648, 32'hc295181d, 32'h4288234d, 32'hc2267872, 32'hc0884555, 32'hc2b87db0};
test_output[23608:23615] = '{32'h0, 32'h42a8ac18, 32'h0, 32'h0, 32'h4288234d, 32'h0, 32'h0, 32'h0};
test_input[23616:23623] = '{32'h4184c112, 32'hc1fc0389, 32'hc2829ce1, 32'h3fe39c3d, 32'h427d1faa, 32'hc2aee489, 32'hc240602f, 32'h422de35c};
test_output[23616:23623] = '{32'h4184c112, 32'h0, 32'h0, 32'h3fe39c3d, 32'h427d1faa, 32'h0, 32'h0, 32'h422de35c};
test_input[23624:23631] = '{32'hc2bc46e9, 32'hc2b3239e, 32'h42635b1c, 32'h424a75e4, 32'hc1b5b506, 32'h404943d0, 32'hc286c01c, 32'h42889e48};
test_output[23624:23631] = '{32'h0, 32'h0, 32'h42635b1c, 32'h424a75e4, 32'h0, 32'h404943d0, 32'h0, 32'h42889e48};
test_input[23632:23639] = '{32'hc212c98e, 32'h42b85d1a, 32'hc2b0bec2, 32'h422827b8, 32'hc1f2d3f9, 32'hc26a3373, 32'h425348c3, 32'hc2aad2bd};
test_output[23632:23639] = '{32'h0, 32'h42b85d1a, 32'h0, 32'h422827b8, 32'h0, 32'h0, 32'h425348c3, 32'h0};
test_input[23640:23647] = '{32'h428911bd, 32'h41b7099f, 32'h4261416b, 32'hc2805171, 32'h41cbd8a5, 32'h42b7545a, 32'hc1f13321, 32'hc1c1acad};
test_output[23640:23647] = '{32'h428911bd, 32'h41b7099f, 32'h4261416b, 32'h0, 32'h41cbd8a5, 32'h42b7545a, 32'h0, 32'h0};
test_input[23648:23655] = '{32'h429160de, 32'hc24e3088, 32'hbe621399, 32'h42895b77, 32'h4251dc4f, 32'h427a1f5d, 32'h42b87fb3, 32'hc1f70ace};
test_output[23648:23655] = '{32'h429160de, 32'h0, 32'h0, 32'h42895b77, 32'h4251dc4f, 32'h427a1f5d, 32'h42b87fb3, 32'h0};
test_input[23656:23663] = '{32'hc2b9cfa0, 32'hc23f0e5f, 32'h425731d9, 32'h41612196, 32'h422efd9b, 32'h4293df05, 32'h41aa2ef3, 32'h41a70555};
test_output[23656:23663] = '{32'h0, 32'h0, 32'h425731d9, 32'h41612196, 32'h422efd9b, 32'h4293df05, 32'h41aa2ef3, 32'h41a70555};
test_input[23664:23671] = '{32'h4208e07c, 32'hc20c59ab, 32'hc22551f9, 32'hc2c6bd6b, 32'h42694977, 32'h427f3269, 32'hc2c265d4, 32'hc0b52131};
test_output[23664:23671] = '{32'h4208e07c, 32'h0, 32'h0, 32'h0, 32'h42694977, 32'h427f3269, 32'h0, 32'h0};
test_input[23672:23679] = '{32'hc284b3ed, 32'h4252ea84, 32'h429f62fd, 32'h41497987, 32'hc2a72426, 32'hc298f68d, 32'h41f7335f, 32'hc2186aac};
test_output[23672:23679] = '{32'h0, 32'h4252ea84, 32'h429f62fd, 32'h41497987, 32'h0, 32'h0, 32'h41f7335f, 32'h0};
test_input[23680:23687] = '{32'hc08b3ee6, 32'h4296e073, 32'h42c546f1, 32'h42919b44, 32'hc2a8f7ce, 32'h42bc7473, 32'h428965d6, 32'hc29a7624};
test_output[23680:23687] = '{32'h0, 32'h4296e073, 32'h42c546f1, 32'h42919b44, 32'h0, 32'h42bc7473, 32'h428965d6, 32'h0};
test_input[23688:23695] = '{32'h40454478, 32'h42ade478, 32'h423ae639, 32'hc2a4e030, 32'hc13405b1, 32'hc25fd4f3, 32'hc27e7edb, 32'hc235ebeb};
test_output[23688:23695] = '{32'h40454478, 32'h42ade478, 32'h423ae639, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23696:23703] = '{32'h42248198, 32'h42a3e3f8, 32'hc2712051, 32'hc27939e1, 32'h42955783, 32'h429b0552, 32'hc1a80b38, 32'h4224f632};
test_output[23696:23703] = '{32'h42248198, 32'h42a3e3f8, 32'h0, 32'h0, 32'h42955783, 32'h429b0552, 32'h0, 32'h4224f632};
test_input[23704:23711] = '{32'h42846e1b, 32'h41875d58, 32'h422ef38d, 32'hc2a76bf9, 32'hc297da1e, 32'h42c77861, 32'h4291a701, 32'h41f4d9a4};
test_output[23704:23711] = '{32'h42846e1b, 32'h41875d58, 32'h422ef38d, 32'h0, 32'h0, 32'h42c77861, 32'h4291a701, 32'h41f4d9a4};
test_input[23712:23719] = '{32'h4293d4fa, 32'hc17d2273, 32'hc1c829e1, 32'hc28cc54a, 32'h42c54f44, 32'h42bcadc6, 32'h429af25f, 32'h42911daa};
test_output[23712:23719] = '{32'h4293d4fa, 32'h0, 32'h0, 32'h0, 32'h42c54f44, 32'h42bcadc6, 32'h429af25f, 32'h42911daa};
test_input[23720:23727] = '{32'h42ab8e4a, 32'hc2248b71, 32'h4272ac3e, 32'hc21c5c07, 32'h42258e66, 32'hc2c7d9c8, 32'h4176890d, 32'h42963a1f};
test_output[23720:23727] = '{32'h42ab8e4a, 32'h0, 32'h4272ac3e, 32'h0, 32'h42258e66, 32'h0, 32'h4176890d, 32'h42963a1f};
test_input[23728:23735] = '{32'hbcc834d5, 32'h4294e828, 32'hc1fdc9d9, 32'h4288d4e8, 32'h42bd03dc, 32'h41d977e0, 32'hc2bacd8d, 32'h42b9a065};
test_output[23728:23735] = '{32'h0, 32'h4294e828, 32'h0, 32'h4288d4e8, 32'h42bd03dc, 32'h41d977e0, 32'h0, 32'h42b9a065};
test_input[23736:23743] = '{32'h420fb318, 32'hc2290e3d, 32'hc2c44be9, 32'hc2336ec6, 32'h4222d12b, 32'hc26dda5b, 32'h4269d578, 32'hc289b057};
test_output[23736:23743] = '{32'h420fb318, 32'h0, 32'h0, 32'h0, 32'h4222d12b, 32'h0, 32'h4269d578, 32'h0};
test_input[23744:23751] = '{32'h41b29791, 32'h42aa923f, 32'hc25482ba, 32'h40b422e3, 32'h42b99dd5, 32'hc18f67f0, 32'h402f3216, 32'h41c1dcb5};
test_output[23744:23751] = '{32'h41b29791, 32'h42aa923f, 32'h0, 32'h40b422e3, 32'h42b99dd5, 32'h0, 32'h402f3216, 32'h41c1dcb5};
test_input[23752:23759] = '{32'h41bb6c14, 32'hc29eb950, 32'hc25dc91d, 32'hc28b21eb, 32'hc25f2d65, 32'hc21cd384, 32'h424a4b7b, 32'h426384c4};
test_output[23752:23759] = '{32'h41bb6c14, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h424a4b7b, 32'h426384c4};
test_input[23760:23767] = '{32'h425d8dc7, 32'hc249b1be, 32'h3ef7885c, 32'h4284f507, 32'h4211a607, 32'h422127dd, 32'hc21f57d2, 32'h426bf0c6};
test_output[23760:23767] = '{32'h425d8dc7, 32'h0, 32'h3ef7885c, 32'h4284f507, 32'h4211a607, 32'h422127dd, 32'h0, 32'h426bf0c6};
test_input[23768:23775] = '{32'hc29cc817, 32'h429bc354, 32'hc26d3d08, 32'h426ad96b, 32'hc2b62f7d, 32'h42660b04, 32'hc22cb528, 32'h41833ba2};
test_output[23768:23775] = '{32'h0, 32'h429bc354, 32'h0, 32'h426ad96b, 32'h0, 32'h42660b04, 32'h0, 32'h41833ba2};
test_input[23776:23783] = '{32'h42a00371, 32'h429cca88, 32'hc28982f9, 32'hc1f2d8c8, 32'hc2256e9b, 32'hc1fa15c9, 32'hc234ef5d, 32'h42a33869};
test_output[23776:23783] = '{32'h42a00371, 32'h429cca88, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a33869};
test_input[23784:23791] = '{32'h41024cf9, 32'h42390244, 32'hc0791965, 32'hc25e551a, 32'h424b7d88, 32'h419eb82e, 32'h4166c33e, 32'hc202ee7f};
test_output[23784:23791] = '{32'h41024cf9, 32'h42390244, 32'h0, 32'h0, 32'h424b7d88, 32'h419eb82e, 32'h4166c33e, 32'h0};
test_input[23792:23799] = '{32'h421a97b0, 32'hc2167acd, 32'hc16783bd, 32'hc26e1951, 32'h428abed8, 32'hc28accfa, 32'h41ed8646, 32'h41dbe3ae};
test_output[23792:23799] = '{32'h421a97b0, 32'h0, 32'h0, 32'h0, 32'h428abed8, 32'h0, 32'h41ed8646, 32'h41dbe3ae};
test_input[23800:23807] = '{32'hc2932fbe, 32'h42004aeb, 32'hc2168e5d, 32'h41fa82ea, 32'hc233d446, 32'h41e2a4d3, 32'h4186605f, 32'h429d69b6};
test_output[23800:23807] = '{32'h0, 32'h42004aeb, 32'h0, 32'h41fa82ea, 32'h0, 32'h41e2a4d3, 32'h4186605f, 32'h429d69b6};
test_input[23808:23815] = '{32'h42819391, 32'hc232f3ab, 32'h42154c37, 32'h424f3f98, 32'hc2608f9f, 32'hc2bf4d55, 32'h42955ade, 32'h4219e72c};
test_output[23808:23815] = '{32'h42819391, 32'h0, 32'h42154c37, 32'h424f3f98, 32'h0, 32'h0, 32'h42955ade, 32'h4219e72c};
test_input[23816:23823] = '{32'hc1b9cb0e, 32'hc293176f, 32'hc294545a, 32'hc12db77b, 32'hc1c48693, 32'hc2555330, 32'hbec5728c, 32'h40d0b95b};
test_output[23816:23823] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40d0b95b};
test_input[23824:23831] = '{32'h42bc45af, 32'hc2b92b77, 32'h42a50086, 32'h426bab7b, 32'hc254d5fb, 32'hc2c3e0ee, 32'h425f8fe6, 32'hc2810fc2};
test_output[23824:23831] = '{32'h42bc45af, 32'h0, 32'h42a50086, 32'h426bab7b, 32'h0, 32'h0, 32'h425f8fe6, 32'h0};
test_input[23832:23839] = '{32'h428adff2, 32'hc2a55a29, 32'hc292d9d2, 32'hc2b45412, 32'hc211f8e6, 32'h4105cd23, 32'hc27da065, 32'h41c1d3ce};
test_output[23832:23839] = '{32'h428adff2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4105cd23, 32'h0, 32'h41c1d3ce};
test_input[23840:23847] = '{32'h4297d6ae, 32'hc1b0cbd3, 32'hc2433aa0, 32'h4240707c, 32'hc27d2ea7, 32'hc258a183, 32'h41fa8cf9, 32'hc2b66dd2};
test_output[23840:23847] = '{32'h4297d6ae, 32'h0, 32'h0, 32'h4240707c, 32'h0, 32'h0, 32'h41fa8cf9, 32'h0};
test_input[23848:23855] = '{32'h429c8fe6, 32'h42c0248f, 32'hc2900401, 32'hc2b6ac19, 32'hc1b128ba, 32'hbf197c4e, 32'hc2421bda, 32'hc29eb6ab};
test_output[23848:23855] = '{32'h429c8fe6, 32'h42c0248f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23856:23863] = '{32'h41b90bca, 32'h42902a1f, 32'hc1a87713, 32'h4230daf5, 32'h428847c0, 32'hc13f2d24, 32'hc2706b05, 32'hc2955fdc};
test_output[23856:23863] = '{32'h41b90bca, 32'h42902a1f, 32'h0, 32'h4230daf5, 32'h428847c0, 32'h0, 32'h0, 32'h0};
test_input[23864:23871] = '{32'h42602131, 32'hc1a54303, 32'hc2a9eaea, 32'hc29e8d15, 32'h41b97b71, 32'hc22fc330, 32'h42234250, 32'hc0b710cc};
test_output[23864:23871] = '{32'h42602131, 32'h0, 32'h0, 32'h0, 32'h41b97b71, 32'h0, 32'h42234250, 32'h0};
test_input[23872:23879] = '{32'h3f1623ab, 32'h423d1695, 32'hbef95949, 32'h4115201d, 32'h42a7d28c, 32'hc26e7593, 32'h4287f28c, 32'h42a1a4c2};
test_output[23872:23879] = '{32'h3f1623ab, 32'h423d1695, 32'h0, 32'h4115201d, 32'h42a7d28c, 32'h0, 32'h4287f28c, 32'h42a1a4c2};
test_input[23880:23887] = '{32'h427aeca4, 32'hc193ea51, 32'hc28bfa23, 32'h42acb048, 32'h42909949, 32'hc2854acc, 32'hc21e735d, 32'h4281c4a2};
test_output[23880:23887] = '{32'h427aeca4, 32'h0, 32'h0, 32'h42acb048, 32'h42909949, 32'h0, 32'h0, 32'h4281c4a2};
test_input[23888:23895] = '{32'h42970457, 32'h3e7fbab3, 32'hc290952c, 32'hc2352b7d, 32'hc217d82a, 32'h42a40d07, 32'h41f4d5d3, 32'hc284a581};
test_output[23888:23895] = '{32'h42970457, 32'h3e7fbab3, 32'h0, 32'h0, 32'h0, 32'h42a40d07, 32'h41f4d5d3, 32'h0};
test_input[23896:23903] = '{32'h428d27f3, 32'hc20e9277, 32'h426b574d, 32'h4207920a, 32'h42a99e55, 32'hc256ecbb, 32'hc295d9d1, 32'h428d1972};
test_output[23896:23903] = '{32'h428d27f3, 32'h0, 32'h426b574d, 32'h4207920a, 32'h42a99e55, 32'h0, 32'h0, 32'h428d1972};
test_input[23904:23911] = '{32'h426f97ab, 32'hc288378f, 32'hc26bff6b, 32'hc2249198, 32'h428f07a0, 32'hc2b02df9, 32'hc2bee390, 32'h41409061};
test_output[23904:23911] = '{32'h426f97ab, 32'h0, 32'h0, 32'h0, 32'h428f07a0, 32'h0, 32'h0, 32'h41409061};
test_input[23912:23919] = '{32'h4272b3b1, 32'hc2c31b29, 32'h419795ea, 32'hc21027f8, 32'hc28db3bf, 32'hc25ce71f, 32'h4232ab9a, 32'h424d79c5};
test_output[23912:23919] = '{32'h4272b3b1, 32'h0, 32'h419795ea, 32'h0, 32'h0, 32'h0, 32'h4232ab9a, 32'h424d79c5};
test_input[23920:23927] = '{32'h415c1d0a, 32'h42af89e8, 32'hc233e303, 32'h40a04564, 32'hc0597308, 32'h429500b2, 32'hc1b73e79, 32'hc2a60a45};
test_output[23920:23927] = '{32'h415c1d0a, 32'h42af89e8, 32'h0, 32'h40a04564, 32'h0, 32'h429500b2, 32'h0, 32'h0};
test_input[23928:23935] = '{32'h42b7d186, 32'hc0539266, 32'h414eaa36, 32'hc161502d, 32'hc19243e2, 32'hc2c7171d, 32'hc2a928b2, 32'hc28ccb12};
test_output[23928:23935] = '{32'h42b7d186, 32'h0, 32'h414eaa36, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23936:23943] = '{32'h429ec88f, 32'hc1983c26, 32'hc2070978, 32'h4141a4b7, 32'h4296d1c6, 32'hc281c991, 32'hc25180a5, 32'hc230ddea};
test_output[23936:23943] = '{32'h429ec88f, 32'h0, 32'h0, 32'h4141a4b7, 32'h4296d1c6, 32'h0, 32'h0, 32'h0};
test_input[23944:23951] = '{32'h42884f44, 32'h41302f24, 32'h42a7d3ea, 32'h40ab3eb7, 32'hc1c98f48, 32'hc273c374, 32'hc22d2073, 32'hc240f66e};
test_output[23944:23951] = '{32'h42884f44, 32'h41302f24, 32'h42a7d3ea, 32'h40ab3eb7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23952:23959] = '{32'h40e6bd1d, 32'hc2b153e7, 32'h415bca4c, 32'hc1f2ec00, 32'h4292f5cf, 32'hc1c82ac8, 32'h41bb3c0c, 32'h423be529};
test_output[23952:23959] = '{32'h40e6bd1d, 32'h0, 32'h415bca4c, 32'h0, 32'h4292f5cf, 32'h0, 32'h41bb3c0c, 32'h423be529};
test_input[23960:23967] = '{32'h42854796, 32'hc2974857, 32'h428e191e, 32'h410e4296, 32'hc2821338, 32'hc26d716c, 32'hc2c126d4, 32'hc2c7b3c8};
test_output[23960:23967] = '{32'h42854796, 32'h0, 32'h428e191e, 32'h410e4296, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23968:23975] = '{32'h4268dae2, 32'h4241abc0, 32'h41c5f954, 32'hc283d5c7, 32'h41cf5704, 32'hc2880bf3, 32'h41d0585e, 32'hc10daba1};
test_output[23968:23975] = '{32'h4268dae2, 32'h4241abc0, 32'h41c5f954, 32'h0, 32'h41cf5704, 32'h0, 32'h41d0585e, 32'h0};
test_input[23976:23983] = '{32'h41e44568, 32'h42517247, 32'h42842856, 32'h42a84323, 32'hbe3affb8, 32'hc231d2fe, 32'hc251975a, 32'h421f5387};
test_output[23976:23983] = '{32'h41e44568, 32'h42517247, 32'h42842856, 32'h42a84323, 32'h0, 32'h0, 32'h0, 32'h421f5387};
test_input[23984:23991] = '{32'h4245f4c1, 32'h4285e15e, 32'hc21479d9, 32'h408d8f1e, 32'hc2b2ce65, 32'h429dfd86, 32'h41bf820a, 32'h42a56e06};
test_output[23984:23991] = '{32'h4245f4c1, 32'h4285e15e, 32'h0, 32'h408d8f1e, 32'h0, 32'h429dfd86, 32'h41bf820a, 32'h42a56e06};
test_input[23992:23999] = '{32'h4033093a, 32'hc2be6901, 32'h42189e6e, 32'h429b8c3b, 32'h42979787, 32'h417b2f6a, 32'h417c62e8, 32'hc2b4ed62};
test_output[23992:23999] = '{32'h4033093a, 32'h0, 32'h42189e6e, 32'h429b8c3b, 32'h42979787, 32'h417b2f6a, 32'h417c62e8, 32'h0};
test_input[24000:24007] = '{32'hc2ba3080, 32'h425f1b5e, 32'h426ceb72, 32'hc1e6c2a8, 32'hc20ab703, 32'hc19dd0ec, 32'h40368c52, 32'h42ab8a19};
test_output[24000:24007] = '{32'h0, 32'h425f1b5e, 32'h426ceb72, 32'h0, 32'h0, 32'h0, 32'h40368c52, 32'h42ab8a19};
test_input[24008:24015] = '{32'hc2051559, 32'hc1656bf6, 32'hc0fdf830, 32'h4114fe4e, 32'h42901447, 32'h4174e5d5, 32'h424a351e, 32'hc2a4bbb6};
test_output[24008:24015] = '{32'h0, 32'h0, 32'h0, 32'h4114fe4e, 32'h42901447, 32'h4174e5d5, 32'h424a351e, 32'h0};
test_input[24016:24023] = '{32'h41f30571, 32'hc2604a21, 32'hc212e449, 32'hc1a032be, 32'hc29f3697, 32'h42b5bbb9, 32'hc224f6e0, 32'hc289f765};
test_output[24016:24023] = '{32'h41f30571, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b5bbb9, 32'h0, 32'h0};
test_input[24024:24031] = '{32'hc25f294e, 32'hc2526f07, 32'h42a0c1cf, 32'h4124e883, 32'hc19103c0, 32'h42552806, 32'hc0816653, 32'h42b31857};
test_output[24024:24031] = '{32'h0, 32'h0, 32'h42a0c1cf, 32'h4124e883, 32'h0, 32'h42552806, 32'h0, 32'h42b31857};
test_input[24032:24039] = '{32'hc1926dca, 32'hc272f408, 32'h41525331, 32'hc18dae55, 32'h41352b54, 32'h414036bd, 32'h41a740b8, 32'hc136064f};
test_output[24032:24039] = '{32'h0, 32'h0, 32'h41525331, 32'h0, 32'h41352b54, 32'h414036bd, 32'h41a740b8, 32'h0};
test_input[24040:24047] = '{32'h426883e5, 32'hc1d96036, 32'h422aa1c5, 32'h4222c788, 32'h4289bc9b, 32'h4275d76c, 32'h41e5d842, 32'h4278e37f};
test_output[24040:24047] = '{32'h426883e5, 32'h0, 32'h422aa1c5, 32'h4222c788, 32'h4289bc9b, 32'h4275d76c, 32'h41e5d842, 32'h4278e37f};
test_input[24048:24055] = '{32'hc18fc7e7, 32'h42b84741, 32'h41891c21, 32'h41213422, 32'h42263c2a, 32'hc2c11c79, 32'h42789601, 32'h40a6dfe0};
test_output[24048:24055] = '{32'h0, 32'h42b84741, 32'h41891c21, 32'h41213422, 32'h42263c2a, 32'h0, 32'h42789601, 32'h40a6dfe0};
test_input[24056:24063] = '{32'h420c2aa3, 32'hc2a369b6, 32'h42942cc3, 32'h4269c03f, 32'h41885e6d, 32'h4293d23f, 32'h4206399f, 32'hc234fdba};
test_output[24056:24063] = '{32'h420c2aa3, 32'h0, 32'h42942cc3, 32'h4269c03f, 32'h41885e6d, 32'h4293d23f, 32'h4206399f, 32'h0};
test_input[24064:24071] = '{32'hc2942ea5, 32'hc2823954, 32'h41a4a0bd, 32'h410cd51c, 32'h408db7b5, 32'hc2a66209, 32'h42891544, 32'h42b65c54};
test_output[24064:24071] = '{32'h0, 32'h0, 32'h41a4a0bd, 32'h410cd51c, 32'h408db7b5, 32'h0, 32'h42891544, 32'h42b65c54};
test_input[24072:24079] = '{32'h41d334e2, 32'h42555f77, 32'hc257aa13, 32'h42725121, 32'hc11847a0, 32'hc1e6170c, 32'hc2a76263, 32'hc2b9d212};
test_output[24072:24079] = '{32'h41d334e2, 32'h42555f77, 32'h0, 32'h42725121, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24080:24087] = '{32'h428704c6, 32'h41c59c54, 32'hc2beb269, 32'h42a4ff24, 32'hc2977cf6, 32'hc2839888, 32'hc1f3ad9f, 32'h3f711d24};
test_output[24080:24087] = '{32'h428704c6, 32'h41c59c54, 32'h0, 32'h42a4ff24, 32'h0, 32'h0, 32'h0, 32'h3f711d24};
test_input[24088:24095] = '{32'hbe9cb6aa, 32'h42b9797c, 32'h42c6e18a, 32'hc2819808, 32'hc23df303, 32'h41cb3f73, 32'h4234841d, 32'h4128f1cf};
test_output[24088:24095] = '{32'h0, 32'h42b9797c, 32'h42c6e18a, 32'h0, 32'h0, 32'h41cb3f73, 32'h4234841d, 32'h4128f1cf};
test_input[24096:24103] = '{32'hc24c4c34, 32'hc2523752, 32'hc2bdb73a, 32'hc2488a22, 32'hc036517e, 32'h428fae40, 32'hc22154a2, 32'hc2b34e91};
test_output[24096:24103] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428fae40, 32'h0, 32'h0};
test_input[24104:24111] = '{32'h42c0294b, 32'hc27cf3ec, 32'hc2ba39ea, 32'h4281cf78, 32'h3f997548, 32'hc2b8d6bb, 32'hc11c3f1f, 32'h42aad921};
test_output[24104:24111] = '{32'h42c0294b, 32'h0, 32'h0, 32'h4281cf78, 32'h3f997548, 32'h0, 32'h0, 32'h42aad921};
test_input[24112:24119] = '{32'h420bb01b, 32'h42a4c5ff, 32'h420ed2c8, 32'hc1acb60b, 32'hc0ffccf1, 32'h42abe494, 32'h4126f95d, 32'hc2a794db};
test_output[24112:24119] = '{32'h420bb01b, 32'h42a4c5ff, 32'h420ed2c8, 32'h0, 32'h0, 32'h42abe494, 32'h4126f95d, 32'h0};
test_input[24120:24127] = '{32'hc0ba6d24, 32'h41e37b83, 32'hc260ad5b, 32'h421461c5, 32'hc282ad07, 32'hc28bbf2b, 32'hc29f5b2c, 32'hc14c9a60};
test_output[24120:24127] = '{32'h0, 32'h41e37b83, 32'h0, 32'h421461c5, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24128:24135] = '{32'h42abba84, 32'h429de253, 32'hc267423c, 32'hc1db26df, 32'hc2132013, 32'hc27e3913, 32'h4099e730, 32'h423df9f8};
test_output[24128:24135] = '{32'h42abba84, 32'h429de253, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4099e730, 32'h423df9f8};
test_input[24136:24143] = '{32'h42067aa0, 32'h4219ff6c, 32'h42597110, 32'h42a61720, 32'h428cf1a5, 32'h418b4c7b, 32'hc266690d, 32'hc2707e15};
test_output[24136:24143] = '{32'h42067aa0, 32'h4219ff6c, 32'h42597110, 32'h42a61720, 32'h428cf1a5, 32'h418b4c7b, 32'h0, 32'h0};
test_input[24144:24151] = '{32'h424fc51c, 32'h4241705c, 32'h42545389, 32'h42c39575, 32'h422d9f01, 32'h42bd49ac, 32'h428f5418, 32'h42a110d9};
test_output[24144:24151] = '{32'h424fc51c, 32'h4241705c, 32'h42545389, 32'h42c39575, 32'h422d9f01, 32'h42bd49ac, 32'h428f5418, 32'h42a110d9};
test_input[24152:24159] = '{32'hc252a67d, 32'hc1fe0107, 32'hc2c36fe5, 32'hc0c1e642, 32'hc1040a5c, 32'h420059bc, 32'hc1f2ac20, 32'h41e5ea39};
test_output[24152:24159] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420059bc, 32'h0, 32'h41e5ea39};
test_input[24160:24167] = '{32'h424f29df, 32'h425f2925, 32'h41967398, 32'h4265de89, 32'h425841b8, 32'h42b0d6ac, 32'h42782d82, 32'hc2976275};
test_output[24160:24167] = '{32'h424f29df, 32'h425f2925, 32'h41967398, 32'h4265de89, 32'h425841b8, 32'h42b0d6ac, 32'h42782d82, 32'h0};
test_input[24168:24175] = '{32'hc2976420, 32'hc282f5ea, 32'h42055721, 32'h4186d001, 32'hc17f4de8, 32'hc0f6e8e2, 32'h429db520, 32'hc27fb29d};
test_output[24168:24175] = '{32'h0, 32'h0, 32'h42055721, 32'h4186d001, 32'h0, 32'h0, 32'h429db520, 32'h0};
test_input[24176:24183] = '{32'h42adc93d, 32'hc09ed0cd, 32'hc1b2cbb4, 32'h428d4981, 32'hc1d9df1f, 32'h4266527d, 32'h41e2003d, 32'hc28df760};
test_output[24176:24183] = '{32'h42adc93d, 32'h0, 32'h0, 32'h428d4981, 32'h0, 32'h4266527d, 32'h41e2003d, 32'h0};
test_input[24184:24191] = '{32'hc0f4e5bd, 32'h41bf2b27, 32'hc2af9a95, 32'h424381ef, 32'hc2566c5b, 32'h3ebf90a1, 32'hc29b8a5d, 32'hc1de20f7};
test_output[24184:24191] = '{32'h0, 32'h41bf2b27, 32'h0, 32'h424381ef, 32'h0, 32'h3ebf90a1, 32'h0, 32'h0};
test_input[24192:24199] = '{32'hc1847c49, 32'h42186f03, 32'h42ab41ce, 32'h41f347b3, 32'hc28126b4, 32'hc288fadc, 32'h4093ec10, 32'hc22c8c5f};
test_output[24192:24199] = '{32'h0, 32'h42186f03, 32'h42ab41ce, 32'h41f347b3, 32'h0, 32'h0, 32'h4093ec10, 32'h0};
test_input[24200:24207] = '{32'hc2a00aba, 32'h4197ef4a, 32'hc1514456, 32'hc0b8ecb7, 32'h40aa52c6, 32'h42473966, 32'h421c6bcf, 32'hc2c32f5e};
test_output[24200:24207] = '{32'h0, 32'h4197ef4a, 32'h0, 32'h0, 32'h40aa52c6, 32'h42473966, 32'h421c6bcf, 32'h0};
test_input[24208:24215] = '{32'h42c486ec, 32'h41ca9a2c, 32'h423d9f9f, 32'hc22549e1, 32'hc2c488d5, 32'hc1c4f3bf, 32'h421ce2d8, 32'h421f8a86};
test_output[24208:24215] = '{32'h42c486ec, 32'h41ca9a2c, 32'h423d9f9f, 32'h0, 32'h0, 32'h0, 32'h421ce2d8, 32'h421f8a86};
test_input[24216:24223] = '{32'hc2c76945, 32'h42106ea0, 32'h41fd0daf, 32'hc19189ee, 32'h419fedf5, 32'h4296e1e4, 32'h4227e91b, 32'h421103a8};
test_output[24216:24223] = '{32'h0, 32'h42106ea0, 32'h41fd0daf, 32'h0, 32'h419fedf5, 32'h4296e1e4, 32'h4227e91b, 32'h421103a8};
test_input[24224:24231] = '{32'h42c034df, 32'h42709661, 32'hc26a171c, 32'h42541ae6, 32'hc1854366, 32'h421ce7a1, 32'hc2986e07, 32'hc2007b88};
test_output[24224:24231] = '{32'h42c034df, 32'h42709661, 32'h0, 32'h42541ae6, 32'h0, 32'h421ce7a1, 32'h0, 32'h0};
test_input[24232:24239] = '{32'hc2b005af, 32'hc24663e7, 32'h42a55c23, 32'h429806e8, 32'h41da7c38, 32'h41a0cc9b, 32'hc108473a, 32'hc06f2aa1};
test_output[24232:24239] = '{32'h0, 32'h0, 32'h42a55c23, 32'h429806e8, 32'h41da7c38, 32'h41a0cc9b, 32'h0, 32'h0};
test_input[24240:24247] = '{32'h42525c2c, 32'hc20b6c5c, 32'hc11005b6, 32'h428c3bb4, 32'hc1921abd, 32'hc296ec9f, 32'h42a978e6, 32'h42285ce8};
test_output[24240:24247] = '{32'h42525c2c, 32'h0, 32'h0, 32'h428c3bb4, 32'h0, 32'h0, 32'h42a978e6, 32'h42285ce8};
test_input[24248:24255] = '{32'h42c4489a, 32'h3ff2b369, 32'hc26e610e, 32'h3fce6c93, 32'hc13f1062, 32'h41cadf39, 32'hc1b9951d, 32'hc283a0aa};
test_output[24248:24255] = '{32'h42c4489a, 32'h3ff2b369, 32'h0, 32'h3fce6c93, 32'h0, 32'h41cadf39, 32'h0, 32'h0};
test_input[24256:24263] = '{32'h425631bf, 32'h4229a762, 32'h41d89c7d, 32'hc0d6cd37, 32'hc2b42f34, 32'h42034d16, 32'hc18f41ee, 32'h424a704c};
test_output[24256:24263] = '{32'h425631bf, 32'h4229a762, 32'h41d89c7d, 32'h0, 32'h0, 32'h42034d16, 32'h0, 32'h424a704c};
test_input[24264:24271] = '{32'hc222b627, 32'h41fc90ee, 32'h421bf2c1, 32'hc11bf5ed, 32'h41db72ad, 32'h4206c855, 32'h410a768f, 32'h42a4be1d};
test_output[24264:24271] = '{32'h0, 32'h41fc90ee, 32'h421bf2c1, 32'h0, 32'h41db72ad, 32'h4206c855, 32'h410a768f, 32'h42a4be1d};
test_input[24272:24279] = '{32'hc23ee397, 32'h40b42951, 32'hc20df70e, 32'hc209165a, 32'h428648e6, 32'h4252ae91, 32'h419f91ce, 32'h423b3c0a};
test_output[24272:24279] = '{32'h0, 32'h40b42951, 32'h0, 32'h0, 32'h428648e6, 32'h4252ae91, 32'h419f91ce, 32'h423b3c0a};
test_input[24280:24287] = '{32'hc24c12c4, 32'h4249de67, 32'hc29956ed, 32'h3e470753, 32'h40f5572b, 32'h425ebbd3, 32'hc0e21d61, 32'h42385a00};
test_output[24280:24287] = '{32'h0, 32'h4249de67, 32'h0, 32'h3e470753, 32'h40f5572b, 32'h425ebbd3, 32'h0, 32'h42385a00};
test_input[24288:24295] = '{32'h4280c085, 32'hc2bfefb6, 32'hc2967dcc, 32'hc244d882, 32'h412493e6, 32'h429f991c, 32'hc29b1aef, 32'h40d22fa3};
test_output[24288:24295] = '{32'h4280c085, 32'h0, 32'h0, 32'h0, 32'h412493e6, 32'h429f991c, 32'h0, 32'h40d22fa3};
test_input[24296:24303] = '{32'hc276ae96, 32'hc22c473e, 32'hc2b7c4c3, 32'hc2901705, 32'hc2bfb868, 32'h42b9b670, 32'hc20c590b, 32'hc187fbbe};
test_output[24296:24303] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b9b670, 32'h0, 32'h0};
test_input[24304:24311] = '{32'h429f12d8, 32'h416c83ee, 32'h428a3299, 32'h42a3aabe, 32'hc2557fe9, 32'h423b3539, 32'hc290d457, 32'h4288a4dd};
test_output[24304:24311] = '{32'h429f12d8, 32'h416c83ee, 32'h428a3299, 32'h42a3aabe, 32'h0, 32'h423b3539, 32'h0, 32'h4288a4dd};
test_input[24312:24319] = '{32'hc112caad, 32'hc2c7e8d9, 32'hc133dbf6, 32'h42c79fa9, 32'hc03bf55d, 32'hc27a66ad, 32'h42296f16, 32'hc21e45bb};
test_output[24312:24319] = '{32'h0, 32'h0, 32'h0, 32'h42c79fa9, 32'h0, 32'h0, 32'h42296f16, 32'h0};
test_input[24320:24327] = '{32'hc26cdf08, 32'hc22b8275, 32'h419b6b05, 32'h42ba88e5, 32'hc1fdf1bc, 32'h427d2149, 32'h42b23fd5, 32'h42a75883};
test_output[24320:24327] = '{32'h0, 32'h0, 32'h419b6b05, 32'h42ba88e5, 32'h0, 32'h427d2149, 32'h42b23fd5, 32'h42a75883};
test_input[24328:24335] = '{32'h403d42fe, 32'h41f8dbba, 32'h422b19ca, 32'h42352743, 32'hc0867051, 32'hc26729de, 32'h42bf83b9, 32'hc25a1d6b};
test_output[24328:24335] = '{32'h403d42fe, 32'h41f8dbba, 32'h422b19ca, 32'h42352743, 32'h0, 32'h0, 32'h42bf83b9, 32'h0};
test_input[24336:24343] = '{32'h41cd4858, 32'hc2838769, 32'h425a3a6b, 32'hc1e19d1f, 32'hc1b0a399, 32'h41961009, 32'h41bbb0c8, 32'hc2570d67};
test_output[24336:24343] = '{32'h41cd4858, 32'h0, 32'h425a3a6b, 32'h0, 32'h0, 32'h41961009, 32'h41bbb0c8, 32'h0};
test_input[24344:24351] = '{32'h425e327f, 32'hc287c40a, 32'h4104d379, 32'hc2932cc1, 32'h425748fb, 32'hc270eca0, 32'hc221f988, 32'hc24f559a};
test_output[24344:24351] = '{32'h425e327f, 32'h0, 32'h4104d379, 32'h0, 32'h425748fb, 32'h0, 32'h0, 32'h0};
test_input[24352:24359] = '{32'h417bde09, 32'hc1bbac00, 32'h418b9b1f, 32'h429c8102, 32'hc201b02d, 32'hc2b6efdb, 32'h426b1847, 32'h40e4ec61};
test_output[24352:24359] = '{32'h417bde09, 32'h0, 32'h418b9b1f, 32'h429c8102, 32'h0, 32'h0, 32'h426b1847, 32'h40e4ec61};
test_input[24360:24367] = '{32'hc2527984, 32'h42bd3e1d, 32'hc19ba9f3, 32'h42b778fb, 32'hc2ab18fc, 32'h420ab5ea, 32'hc28f8245, 32'hc2a68a24};
test_output[24360:24367] = '{32'h0, 32'h42bd3e1d, 32'h0, 32'h42b778fb, 32'h0, 32'h420ab5ea, 32'h0, 32'h0};
test_input[24368:24375] = '{32'h41c5406e, 32'h423d17b0, 32'hc2907d75, 32'hc2b551bf, 32'hc22166ff, 32'hc1e17a67, 32'h4283c493, 32'hc21d1d94};
test_output[24368:24375] = '{32'h41c5406e, 32'h423d17b0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4283c493, 32'h0};
test_input[24376:24383] = '{32'hc273e05e, 32'hc2a14c73, 32'h41b52afa, 32'h41be037e, 32'h41822b29, 32'h427ec3a9, 32'hc2c4a5ce, 32'hc188eba1};
test_output[24376:24383] = '{32'h0, 32'h0, 32'h41b52afa, 32'h41be037e, 32'h41822b29, 32'h427ec3a9, 32'h0, 32'h0};
test_input[24384:24391] = '{32'hc22bb591, 32'hc2711177, 32'h411c0741, 32'h42a24ace, 32'h41bbc941, 32'hc2b6df45, 32'hc2bb4b81, 32'h41d99fd1};
test_output[24384:24391] = '{32'h0, 32'h0, 32'h411c0741, 32'h42a24ace, 32'h41bbc941, 32'h0, 32'h0, 32'h41d99fd1};
test_input[24392:24399] = '{32'hc2bc4ca8, 32'hc20f8e8a, 32'h425bf514, 32'hc21dd8b5, 32'hc139f095, 32'hc295a566, 32'hc2128836, 32'h421e6605};
test_output[24392:24399] = '{32'h0, 32'h0, 32'h425bf514, 32'h0, 32'h0, 32'h0, 32'h0, 32'h421e6605};
test_input[24400:24407] = '{32'hc2ab9936, 32'h42514e10, 32'hc24672bd, 32'h42c55e85, 32'h423d8bdb, 32'h3fa55c8f, 32'hc288f8ac, 32'h41affb58};
test_output[24400:24407] = '{32'h0, 32'h42514e10, 32'h0, 32'h42c55e85, 32'h423d8bdb, 32'h3fa55c8f, 32'h0, 32'h41affb58};
test_input[24408:24415] = '{32'h4279aec8, 32'hc2b7e4af, 32'hc19069c3, 32'h4278341e, 32'h41583a6d, 32'h40677880, 32'h40393aea, 32'h423dcfac};
test_output[24408:24415] = '{32'h4279aec8, 32'h0, 32'h0, 32'h4278341e, 32'h41583a6d, 32'h40677880, 32'h40393aea, 32'h423dcfac};
test_input[24416:24423] = '{32'hc236d955, 32'h42961de4, 32'h42b55d63, 32'h428455e9, 32'hc1c39f79, 32'h421723c1, 32'hc1df264f, 32'hc1f77b47};
test_output[24416:24423] = '{32'h0, 32'h42961de4, 32'h42b55d63, 32'h428455e9, 32'h0, 32'h421723c1, 32'h0, 32'h0};
test_input[24424:24431] = '{32'h42aceb88, 32'hc2614581, 32'hc21a6203, 32'hc270f633, 32'hc08d21d3, 32'h42c6aa5d, 32'hc2935a69, 32'h429f8a04};
test_output[24424:24431] = '{32'h42aceb88, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c6aa5d, 32'h0, 32'h429f8a04};
test_input[24432:24439] = '{32'hc2c03c64, 32'hc28eda6d, 32'h424d0696, 32'h4010e56d, 32'h417f4d0f, 32'hc288b2ce, 32'hc148e7b6, 32'hc1cf6a8e};
test_output[24432:24439] = '{32'h0, 32'h0, 32'h424d0696, 32'h4010e56d, 32'h417f4d0f, 32'h0, 32'h0, 32'h0};
test_input[24440:24447] = '{32'hc1a6d3f1, 32'h4214689f, 32'h3f24d869, 32'h423ae5a6, 32'h41d5d92e, 32'hc2117eb9, 32'hc2905246, 32'hc21bbf72};
test_output[24440:24447] = '{32'h0, 32'h4214689f, 32'h3f24d869, 32'h423ae5a6, 32'h41d5d92e, 32'h0, 32'h0, 32'h0};
test_input[24448:24455] = '{32'hc02e3234, 32'hc2bd6b16, 32'hc183d615, 32'hc2c6f857, 32'hc1c9eef7, 32'h422f7fee, 32'h40a6066c, 32'hc22e1483};
test_output[24448:24455] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422f7fee, 32'h40a6066c, 32'h0};
test_input[24456:24463] = '{32'hc2962e1f, 32'h4267b50b, 32'hc2a7905a, 32'hbed425da, 32'h429021db, 32'h4287e434, 32'hc2ad2ce7, 32'h424f97bb};
test_output[24456:24463] = '{32'h0, 32'h4267b50b, 32'h0, 32'h0, 32'h429021db, 32'h4287e434, 32'h0, 32'h424f97bb};
test_input[24464:24471] = '{32'h419c547a, 32'hc2b05d5f, 32'h4205b7f0, 32'h42831c0b, 32'hc25131a0, 32'h4173c594, 32'h4253d4a2, 32'h40be21ba};
test_output[24464:24471] = '{32'h419c547a, 32'h0, 32'h4205b7f0, 32'h42831c0b, 32'h0, 32'h4173c594, 32'h4253d4a2, 32'h40be21ba};
test_input[24472:24479] = '{32'h40689261, 32'hc2877f36, 32'hc2950453, 32'hc20c05b6, 32'h42ac8079, 32'h428711f3, 32'hc2b216f1, 32'hc28430ed};
test_output[24472:24479] = '{32'h40689261, 32'h0, 32'h0, 32'h0, 32'h42ac8079, 32'h428711f3, 32'h0, 32'h0};
test_input[24480:24487] = '{32'h4226c057, 32'h42196c2a, 32'h409c7e57, 32'hc1e859a5, 32'h419a4a24, 32'h4283f73e, 32'hc274f191, 32'hc2935a5c};
test_output[24480:24487] = '{32'h4226c057, 32'h42196c2a, 32'h409c7e57, 32'h0, 32'h419a4a24, 32'h4283f73e, 32'h0, 32'h0};
test_input[24488:24495] = '{32'h42a8be97, 32'hc292c826, 32'hc1dc898e, 32'hc210b7d8, 32'hc2719831, 32'hc100e559, 32'h42349106, 32'h4299aea0};
test_output[24488:24495] = '{32'h42a8be97, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42349106, 32'h4299aea0};
test_input[24496:24503] = '{32'hc22291aa, 32'hc27132ca, 32'h4168ba16, 32'hc297b250, 32'h42bd01bb, 32'hc236e105, 32'h3fbb38ef, 32'h4245b938};
test_output[24496:24503] = '{32'h0, 32'h0, 32'h4168ba16, 32'h0, 32'h42bd01bb, 32'h0, 32'h3fbb38ef, 32'h4245b938};
test_input[24504:24511] = '{32'hc2b07708, 32'hc2266a33, 32'h429edae5, 32'hc2a3fa7a, 32'h41f66b66, 32'hc193f9f2, 32'h4299e3ed, 32'hc2612709};
test_output[24504:24511] = '{32'h0, 32'h0, 32'h429edae5, 32'h0, 32'h41f66b66, 32'h0, 32'h4299e3ed, 32'h0};
test_input[24512:24519] = '{32'hc0dd42ac, 32'h40d6d316, 32'h4231fd8d, 32'h41ec41db, 32'h42b97eea, 32'hc26ee1fb, 32'hc2ab29b9, 32'h406663e2};
test_output[24512:24519] = '{32'h0, 32'h40d6d316, 32'h4231fd8d, 32'h41ec41db, 32'h42b97eea, 32'h0, 32'h0, 32'h406663e2};
test_input[24520:24527] = '{32'h4110e683, 32'hc1f0d1bc, 32'hc249f490, 32'h40a8bd84, 32'h42b15568, 32'h4253cd91, 32'hc222e525, 32'hc27eca61};
test_output[24520:24527] = '{32'h4110e683, 32'h0, 32'h0, 32'h40a8bd84, 32'h42b15568, 32'h4253cd91, 32'h0, 32'h0};
test_input[24528:24535] = '{32'hc2952e31, 32'h4287fb5b, 32'h4263f3da, 32'h4184d4c0, 32'h42abd7a8, 32'h42860612, 32'hc273b7ca, 32'hc2b8c06d};
test_output[24528:24535] = '{32'h0, 32'h4287fb5b, 32'h4263f3da, 32'h4184d4c0, 32'h42abd7a8, 32'h42860612, 32'h0, 32'h0};
test_input[24536:24543] = '{32'h4174b016, 32'hc1f4c632, 32'h4242b373, 32'hc2ab92e6, 32'hc2a3c11d, 32'h42a693c0, 32'h42a6a0fc, 32'hc256e9e2};
test_output[24536:24543] = '{32'h4174b016, 32'h0, 32'h4242b373, 32'h0, 32'h0, 32'h42a693c0, 32'h42a6a0fc, 32'h0};
test_input[24544:24551] = '{32'h42128b18, 32'h4288e40d, 32'h42b67752, 32'hc2a6c061, 32'h4147f52d, 32'hc1213d3c, 32'hc2b0a62c, 32'h42815e3a};
test_output[24544:24551] = '{32'h42128b18, 32'h4288e40d, 32'h42b67752, 32'h0, 32'h4147f52d, 32'h0, 32'h0, 32'h42815e3a};
test_input[24552:24559] = '{32'hc2324b0d, 32'hc281d1ad, 32'h4280d94f, 32'h42bb126e, 32'h42ac24f7, 32'hc2a652b9, 32'h418d6559, 32'h41ddcb1e};
test_output[24552:24559] = '{32'h0, 32'h0, 32'h4280d94f, 32'h42bb126e, 32'h42ac24f7, 32'h0, 32'h418d6559, 32'h41ddcb1e};
test_input[24560:24567] = '{32'hc226ae2e, 32'hc1f4c6c5, 32'h4227fda3, 32'hc2133647, 32'hc2b333e8, 32'h418e726d, 32'h42b825ff, 32'hc2bbe46e};
test_output[24560:24567] = '{32'h0, 32'h0, 32'h4227fda3, 32'h0, 32'h0, 32'h418e726d, 32'h42b825ff, 32'h0};
test_input[24568:24575] = '{32'h428da057, 32'h420faa06, 32'hc2b886ee, 32'h429ebd09, 32'h428d9d1e, 32'h41b6502c, 32'h418a7e0f, 32'hc2baeda2};
test_output[24568:24575] = '{32'h428da057, 32'h420faa06, 32'h0, 32'h429ebd09, 32'h428d9d1e, 32'h41b6502c, 32'h418a7e0f, 32'h0};
test_input[24576:24583] = '{32'h42907c42, 32'hc1b70974, 32'hc12f5cd5, 32'hc04a0443, 32'hc2b46869, 32'h4270bec6, 32'h42b07e2a, 32'hc232ecb0};
test_output[24576:24583] = '{32'h42907c42, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4270bec6, 32'h42b07e2a, 32'h0};
test_input[24584:24591] = '{32'hc2b8b732, 32'h42a22d91, 32'hc2c29a5a, 32'h427a7b1c, 32'h4215035e, 32'hc29a039f, 32'hc1ece55f, 32'h41ae3d84};
test_output[24584:24591] = '{32'h0, 32'h42a22d91, 32'h0, 32'h427a7b1c, 32'h4215035e, 32'h0, 32'h0, 32'h41ae3d84};
test_input[24592:24599] = '{32'hc0e40328, 32'hc2bf8eee, 32'hc28a52fa, 32'h42156df0, 32'h42bd71fd, 32'h421ce7b9, 32'h42b5924e, 32'h417b607f};
test_output[24592:24599] = '{32'h0, 32'h0, 32'h0, 32'h42156df0, 32'h42bd71fd, 32'h421ce7b9, 32'h42b5924e, 32'h417b607f};
test_input[24600:24607] = '{32'h41d50c5f, 32'hc1672091, 32'hc166abd5, 32'h4298cb4c, 32'hc2166054, 32'h42a2441f, 32'h424944d2, 32'h4294ff21};
test_output[24600:24607] = '{32'h41d50c5f, 32'h0, 32'h0, 32'h4298cb4c, 32'h0, 32'h42a2441f, 32'h424944d2, 32'h4294ff21};
test_input[24608:24615] = '{32'hc0ad5b51, 32'hc25e73a1, 32'hc2818b33, 32'hc2c2891f, 32'h42bcd6a0, 32'hc273f365, 32'hc2c1de62, 32'h4275c00b};
test_output[24608:24615] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42bcd6a0, 32'h0, 32'h0, 32'h4275c00b};
test_input[24616:24623] = '{32'h428df016, 32'hc262da44, 32'h422ec8d0, 32'hc249b68f, 32'h3ff080e3, 32'hc275ff09, 32'hc2b31c90, 32'h424fc31c};
test_output[24616:24623] = '{32'h428df016, 32'h0, 32'h422ec8d0, 32'h0, 32'h3ff080e3, 32'h0, 32'h0, 32'h424fc31c};
test_input[24624:24631] = '{32'h429f5956, 32'h4212397a, 32'hc27d7a37, 32'hc1aa23d4, 32'hc243aff4, 32'hc254506d, 32'h421c1c05, 32'hc278703a};
test_output[24624:24631] = '{32'h429f5956, 32'h4212397a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h421c1c05, 32'h0};
test_input[24632:24639] = '{32'h426a12fd, 32'h424d52ec, 32'hc180899e, 32'hc24d70ad, 32'hc2316abd, 32'hc2aa62e5, 32'h412c2610, 32'hc1116442};
test_output[24632:24639] = '{32'h426a12fd, 32'h424d52ec, 32'h0, 32'h0, 32'h0, 32'h0, 32'h412c2610, 32'h0};
test_input[24640:24647] = '{32'h4236960c, 32'hc267601c, 32'h42887ad7, 32'h422897be, 32'hc27224fb, 32'hc2373524, 32'hc26b801e, 32'h42c20ca1};
test_output[24640:24647] = '{32'h4236960c, 32'h0, 32'h42887ad7, 32'h422897be, 32'h0, 32'h0, 32'h0, 32'h42c20ca1};
test_input[24648:24655] = '{32'h42112aba, 32'hc2bc3601, 32'hc22ca533, 32'h42bd67d2, 32'h42bb2561, 32'hc0f779e1, 32'hc1bf99a1, 32'h426f8ef8};
test_output[24648:24655] = '{32'h42112aba, 32'h0, 32'h0, 32'h42bd67d2, 32'h42bb2561, 32'h0, 32'h0, 32'h426f8ef8};
test_input[24656:24663] = '{32'h402a47e4, 32'h417391f5, 32'hc2b32108, 32'hc24f47c0, 32'hc0a20cc2, 32'hc2794f78, 32'hc251afb5, 32'h42a12ba3};
test_output[24656:24663] = '{32'h402a47e4, 32'h417391f5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a12ba3};
test_input[24664:24671] = '{32'h41bb123f, 32'h41207423, 32'h420f8916, 32'h428d98bc, 32'hc287ffda, 32'h426995e1, 32'h4244855a, 32'h4170f5d2};
test_output[24664:24671] = '{32'h41bb123f, 32'h41207423, 32'h420f8916, 32'h428d98bc, 32'h0, 32'h426995e1, 32'h4244855a, 32'h4170f5d2};
test_input[24672:24679] = '{32'h42c75db5, 32'hc290b3eb, 32'h4132cf6f, 32'h41a40238, 32'hc2793485, 32'h4239b0c4, 32'hc29559d8, 32'hc2244762};
test_output[24672:24679] = '{32'h42c75db5, 32'h0, 32'h4132cf6f, 32'h41a40238, 32'h0, 32'h4239b0c4, 32'h0, 32'h0};
test_input[24680:24687] = '{32'h41adab27, 32'h406df058, 32'hc1fcab1d, 32'hc21aa445, 32'hc283a30f, 32'h425cea05, 32'h41c7e59c, 32'hc199490b};
test_output[24680:24687] = '{32'h41adab27, 32'h406df058, 32'h0, 32'h0, 32'h0, 32'h425cea05, 32'h41c7e59c, 32'h0};
test_input[24688:24695] = '{32'hc2544908, 32'h41b2d29d, 32'hc1db1c02, 32'h41f78298, 32'hc219bf0c, 32'hc2ba0915, 32'hc27e2cc2, 32'hc145fedb};
test_output[24688:24695] = '{32'h0, 32'h41b2d29d, 32'h0, 32'h41f78298, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24696:24703] = '{32'hc21939f9, 32'hc23cb040, 32'hc22f65dc, 32'h41d08be2, 32'h4200f546, 32'hc18f502f, 32'hc2845794, 32'hc2a0e427};
test_output[24696:24703] = '{32'h0, 32'h0, 32'h0, 32'h41d08be2, 32'h4200f546, 32'h0, 32'h0, 32'h0};
test_input[24704:24711] = '{32'hc1dc3e44, 32'hc19943bb, 32'h41845aa1, 32'h41bc8d72, 32'hc1a0e6a8, 32'hc1916e5b, 32'hc26e35fc, 32'hc290e588};
test_output[24704:24711] = '{32'h0, 32'h0, 32'h41845aa1, 32'h41bc8d72, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24712:24719] = '{32'h41efd8c2, 32'h42a8abed, 32'hc2875cdc, 32'h41e51c39, 32'h42c12f51, 32'hc1a79016, 32'hc0a46d60, 32'hc193cdc4};
test_output[24712:24719] = '{32'h41efd8c2, 32'h42a8abed, 32'h0, 32'h41e51c39, 32'h42c12f51, 32'h0, 32'h0, 32'h0};
test_input[24720:24727] = '{32'hc215d5dd, 32'hc2a44c74, 32'h41d272b4, 32'hc28fd413, 32'h428f2bf9, 32'h42a7db92, 32'hc2b39d84, 32'h428401a4};
test_output[24720:24727] = '{32'h0, 32'h0, 32'h41d272b4, 32'h0, 32'h428f2bf9, 32'h42a7db92, 32'h0, 32'h428401a4};
test_input[24728:24735] = '{32'hc1e5262c, 32'h421c8b72, 32'hc2399c79, 32'hc2687930, 32'hc284b436, 32'h428ff3c1, 32'hc21faa45, 32'hc2703c5b};
test_output[24728:24735] = '{32'h0, 32'h421c8b72, 32'h0, 32'h0, 32'h0, 32'h428ff3c1, 32'h0, 32'h0};
test_input[24736:24743] = '{32'hc2473f1c, 32'hc299f28b, 32'h42621b0c, 32'h422bcd96, 32'h3ef0f1ef, 32'hc2574405, 32'h4247d48c, 32'h4247f2a6};
test_output[24736:24743] = '{32'h0, 32'h0, 32'h42621b0c, 32'h422bcd96, 32'h3ef0f1ef, 32'h0, 32'h4247d48c, 32'h4247f2a6};
test_input[24744:24751] = '{32'hc24bc48b, 32'h3f1e1a89, 32'h402f506f, 32'hc29a45c6, 32'h42c6d6d4, 32'hc1ac97c0, 32'hc20e14e5, 32'hc1029df2};
test_output[24744:24751] = '{32'h0, 32'h3f1e1a89, 32'h402f506f, 32'h0, 32'h42c6d6d4, 32'h0, 32'h0, 32'h0};
test_input[24752:24759] = '{32'hc252ee94, 32'h42978a4c, 32'h3f80b772, 32'hc2a15574, 32'hc284b71d, 32'hc29abcdc, 32'h42a70d96, 32'hc2acece3};
test_output[24752:24759] = '{32'h0, 32'h42978a4c, 32'h3f80b772, 32'h0, 32'h0, 32'h0, 32'h42a70d96, 32'h0};
test_input[24760:24767] = '{32'hc23c4ebf, 32'hc12ff2f4, 32'hc291ad35, 32'hc0a85504, 32'hc2b2927d, 32'h41eb844d, 32'h4273f45f, 32'h42ab1cf8};
test_output[24760:24767] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41eb844d, 32'h4273f45f, 32'h42ab1cf8};
test_input[24768:24775] = '{32'hc249f293, 32'h411e5ffb, 32'hc22a9a15, 32'h41f4931b, 32'h4206beb5, 32'h42964340, 32'hc2b605d5, 32'hc20a5584};
test_output[24768:24775] = '{32'h0, 32'h411e5ffb, 32'h0, 32'h41f4931b, 32'h4206beb5, 32'h42964340, 32'h0, 32'h0};
test_input[24776:24783] = '{32'hc280509b, 32'h42b6dc48, 32'hc15a0c77, 32'h421b829a, 32'h419b3067, 32'hc28ab394, 32'hc2c50a81, 32'hc252d500};
test_output[24776:24783] = '{32'h0, 32'h42b6dc48, 32'h0, 32'h421b829a, 32'h419b3067, 32'h0, 32'h0, 32'h0};
test_input[24784:24791] = '{32'h420eecd0, 32'h424afc6c, 32'h421232ac, 32'hc23c6869, 32'h414ab74d, 32'hc17f3323, 32'hc2314098, 32'h41f074a4};
test_output[24784:24791] = '{32'h420eecd0, 32'h424afc6c, 32'h421232ac, 32'h0, 32'h414ab74d, 32'h0, 32'h0, 32'h41f074a4};
test_input[24792:24799] = '{32'hc2a3efe3, 32'h42c7efd5, 32'h41938802, 32'h41ecd003, 32'h42b5952c, 32'h3f98a9fb, 32'h4282bc40, 32'hc22b18b0};
test_output[24792:24799] = '{32'h0, 32'h42c7efd5, 32'h41938802, 32'h41ecd003, 32'h42b5952c, 32'h3f98a9fb, 32'h4282bc40, 32'h0};
test_input[24800:24807] = '{32'hc29047de, 32'h42b66068, 32'h41480a65, 32'h41cbed3f, 32'h423dfabe, 32'hc2989da1, 32'h4127754d, 32'hc2262840};
test_output[24800:24807] = '{32'h0, 32'h42b66068, 32'h41480a65, 32'h41cbed3f, 32'h423dfabe, 32'h0, 32'h4127754d, 32'h0};
test_input[24808:24815] = '{32'h4033b5d6, 32'hc20de451, 32'hc1dbdcbf, 32'hc24e7174, 32'hc1b2ab23, 32'h420fc958, 32'hc2c7c2c2, 32'h420c0c1f};
test_output[24808:24815] = '{32'h4033b5d6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420fc958, 32'h0, 32'h420c0c1f};
test_input[24816:24823] = '{32'hc25d9cb7, 32'h42318466, 32'hc0bef92f, 32'hc28ef974, 32'h429032cb, 32'h42648887, 32'hc296d016, 32'h4199c428};
test_output[24816:24823] = '{32'h0, 32'h42318466, 32'h0, 32'h0, 32'h429032cb, 32'h42648887, 32'h0, 32'h4199c428};
test_input[24824:24831] = '{32'h41fefc43, 32'hc11909cf, 32'hc272182d, 32'h42379c6d, 32'hc2861343, 32'h428ec259, 32'hc0dfc539, 32'h420ffe52};
test_output[24824:24831] = '{32'h41fefc43, 32'h0, 32'h0, 32'h42379c6d, 32'h0, 32'h428ec259, 32'h0, 32'h420ffe52};
test_input[24832:24839] = '{32'h40d6e606, 32'h414259c0, 32'h42933d59, 32'hbcee1937, 32'h4205b380, 32'h426ad65c, 32'h41dbc21d, 32'hc0d9b40b};
test_output[24832:24839] = '{32'h40d6e606, 32'h414259c0, 32'h42933d59, 32'h0, 32'h4205b380, 32'h426ad65c, 32'h41dbc21d, 32'h0};
test_input[24840:24847] = '{32'h41d12ae5, 32'h41cba2a9, 32'h41ed989c, 32'h4202483c, 32'h42060b50, 32'h42947582, 32'hc26da7b4, 32'hc21c325a};
test_output[24840:24847] = '{32'h41d12ae5, 32'h41cba2a9, 32'h41ed989c, 32'h4202483c, 32'h42060b50, 32'h42947582, 32'h0, 32'h0};
test_input[24848:24855] = '{32'h4296de82, 32'h41f5de10, 32'hc2826d12, 32'h42c2503c, 32'hc28fdd7d, 32'hc2bb829f, 32'hc1f67638, 32'hc28bcf07};
test_output[24848:24855] = '{32'h4296de82, 32'h41f5de10, 32'h0, 32'h42c2503c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24856:24863] = '{32'h42c3fd01, 32'h4210810b, 32'hc2b546ce, 32'hc22bf89a, 32'h40fdd26a, 32'h419d6d61, 32'h42a97a44, 32'h42950eb6};
test_output[24856:24863] = '{32'h42c3fd01, 32'h4210810b, 32'h0, 32'h0, 32'h40fdd26a, 32'h419d6d61, 32'h42a97a44, 32'h42950eb6};
test_input[24864:24871] = '{32'h428d443a, 32'h42b10748, 32'h4273e894, 32'hc2357262, 32'h42a57863, 32'h4184d026, 32'hc2b13c0b, 32'hc1a69e51};
test_output[24864:24871] = '{32'h428d443a, 32'h42b10748, 32'h4273e894, 32'h0, 32'h42a57863, 32'h4184d026, 32'h0, 32'h0};
test_input[24872:24879] = '{32'hc04b7cb8, 32'hc267bedd, 32'h411c1244, 32'h42c12c18, 32'hc28a1d98, 32'hc2b2f216, 32'h4205af28, 32'hc228c064};
test_output[24872:24879] = '{32'h0, 32'h0, 32'h411c1244, 32'h42c12c18, 32'h0, 32'h0, 32'h4205af28, 32'h0};
test_input[24880:24887] = '{32'hc19b40cd, 32'hc18da5bd, 32'h428cc3d4, 32'hc05c63e9, 32'hc1fe609a, 32'hc22a8c84, 32'hc04ce7e5, 32'hc0cbb77b};
test_output[24880:24887] = '{32'h0, 32'h0, 32'h428cc3d4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24888:24895] = '{32'h4109655b, 32'h4228c8b5, 32'hc28a294b, 32'h42344b83, 32'h428be5dc, 32'h41fed90a, 32'h4236f0a1, 32'hc1e9d808};
test_output[24888:24895] = '{32'h4109655b, 32'h4228c8b5, 32'h0, 32'h42344b83, 32'h428be5dc, 32'h41fed90a, 32'h4236f0a1, 32'h0};
test_input[24896:24903] = '{32'h424726c8, 32'h42449c6c, 32'hc131bbc7, 32'h415c89dd, 32'h4283e1ba, 32'h42212d6b, 32'hc2213590, 32'hc1b2e949};
test_output[24896:24903] = '{32'h424726c8, 32'h42449c6c, 32'h0, 32'h415c89dd, 32'h4283e1ba, 32'h42212d6b, 32'h0, 32'h0};
test_input[24904:24911] = '{32'hc135bd58, 32'hc2ae624b, 32'hc1a212ac, 32'hc288d536, 32'hc0bfcf8b, 32'h429d70eb, 32'hc2895541, 32'hc2b24672};
test_output[24904:24911] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429d70eb, 32'h0, 32'h0};
test_input[24912:24919] = '{32'hc25be13a, 32'h41c2824a, 32'h4223468c, 32'hc2088adf, 32'h40601ded, 32'hc2b332a9, 32'h4195a46e, 32'h42a85907};
test_output[24912:24919] = '{32'h0, 32'h41c2824a, 32'h4223468c, 32'h0, 32'h40601ded, 32'h0, 32'h4195a46e, 32'h42a85907};
test_input[24920:24927] = '{32'h418646c3, 32'hc0d85134, 32'hbeb97dac, 32'hc2798ead, 32'hc16c3271, 32'hc2bf73ae, 32'hbed692eb, 32'hc23791f3};
test_output[24920:24927] = '{32'h418646c3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24928:24935] = '{32'h427d3b22, 32'hc2601d63, 32'h42873526, 32'hc0da6c05, 32'hc24ebe58, 32'hc14a8be1, 32'h4296c220, 32'h408c5a99};
test_output[24928:24935] = '{32'h427d3b22, 32'h0, 32'h42873526, 32'h0, 32'h0, 32'h0, 32'h4296c220, 32'h408c5a99};
test_input[24936:24943] = '{32'h42802bfb, 32'hc2bea30a, 32'h423a7e4f, 32'h42af8a98, 32'h4148dca0, 32'h42b30d33, 32'hc2aecb0a, 32'h423e3138};
test_output[24936:24943] = '{32'h42802bfb, 32'h0, 32'h423a7e4f, 32'h42af8a98, 32'h4148dca0, 32'h42b30d33, 32'h0, 32'h423e3138};
test_input[24944:24951] = '{32'h422e6de5, 32'h414360e1, 32'hc21b756f, 32'h42bcfaf4, 32'h42655d1a, 32'h41f90260, 32'hc2646228, 32'h423950de};
test_output[24944:24951] = '{32'h422e6de5, 32'h414360e1, 32'h0, 32'h42bcfaf4, 32'h42655d1a, 32'h41f90260, 32'h0, 32'h423950de};
test_input[24952:24959] = '{32'hc20aa85b, 32'hc28b0ab0, 32'h42b1070f, 32'h41169c2c, 32'hc1fe5b88, 32'h413ce10a, 32'h423d0824, 32'hbf09d332};
test_output[24952:24959] = '{32'h0, 32'h0, 32'h42b1070f, 32'h41169c2c, 32'h0, 32'h413ce10a, 32'h423d0824, 32'h0};
test_input[24960:24967] = '{32'h4260630b, 32'hc2c5c0a8, 32'h4296c00a, 32'hc28a61aa, 32'h41d55165, 32'h4031d42c, 32'h4102a23c, 32'h41fb949e};
test_output[24960:24967] = '{32'h4260630b, 32'h0, 32'h4296c00a, 32'h0, 32'h41d55165, 32'h4031d42c, 32'h4102a23c, 32'h41fb949e};
test_input[24968:24975] = '{32'h4256b8ff, 32'h426c8f7e, 32'h42977fbe, 32'h4266805d, 32'h419431e5, 32'h428ad64c, 32'h42bf8698, 32'h427fbdaf};
test_output[24968:24975] = '{32'h4256b8ff, 32'h426c8f7e, 32'h42977fbe, 32'h4266805d, 32'h419431e5, 32'h428ad64c, 32'h42bf8698, 32'h427fbdaf};
test_input[24976:24983] = '{32'h42188cae, 32'h424a150b, 32'h423f2f8c, 32'h4221ed03, 32'hc2afebe4, 32'hc277f9af, 32'h420bad88, 32'h41410062};
test_output[24976:24983] = '{32'h42188cae, 32'h424a150b, 32'h423f2f8c, 32'h4221ed03, 32'h0, 32'h0, 32'h420bad88, 32'h41410062};
test_input[24984:24991] = '{32'h42c7e000, 32'hc270ebb0, 32'h418ca0aa, 32'h423a6121, 32'h42a14966, 32'hc288527d, 32'h421d4d56, 32'h42939cd8};
test_output[24984:24991] = '{32'h42c7e000, 32'h0, 32'h418ca0aa, 32'h423a6121, 32'h42a14966, 32'h0, 32'h421d4d56, 32'h42939cd8};
test_input[24992:24999] = '{32'h418f63fc, 32'hc2c043d2, 32'h429485eb, 32'h42972672, 32'h4275ba7e, 32'h42bdb038, 32'hc2aa4c9d, 32'hc29df31e};
test_output[24992:24999] = '{32'h418f63fc, 32'h0, 32'h429485eb, 32'h42972672, 32'h4275ba7e, 32'h42bdb038, 32'h0, 32'h0};
test_input[25000:25007] = '{32'h3f6aea40, 32'hc1d2a794, 32'h426de657, 32'hc088e7ee, 32'h41b03f70, 32'hc2284e66, 32'h42c196b7, 32'hc2c7f37f};
test_output[25000:25007] = '{32'h3f6aea40, 32'h0, 32'h426de657, 32'h0, 32'h41b03f70, 32'h0, 32'h42c196b7, 32'h0};
test_input[25008:25015] = '{32'hc2a1f6dc, 32'hbfa2c379, 32'h4293d923, 32'hc2a197b1, 32'h4159ffa8, 32'hc2a841ac, 32'h427981e2, 32'hc2155d93};
test_output[25008:25015] = '{32'h0, 32'h0, 32'h4293d923, 32'h0, 32'h4159ffa8, 32'h0, 32'h427981e2, 32'h0};
test_input[25016:25023] = '{32'hc2c63723, 32'h42b5da8b, 32'h40c79112, 32'h429c1026, 32'hbf3c5599, 32'h41b930b0, 32'h410b2a28, 32'h4098ddb1};
test_output[25016:25023] = '{32'h0, 32'h42b5da8b, 32'h40c79112, 32'h429c1026, 32'h0, 32'h41b930b0, 32'h410b2a28, 32'h4098ddb1};
test_input[25024:25031] = '{32'h423bb933, 32'h421b88f3, 32'h429c397a, 32'h40b1d0f4, 32'h4268277b, 32'h42585478, 32'h429ab8c2, 32'h41f6d883};
test_output[25024:25031] = '{32'h423bb933, 32'h421b88f3, 32'h429c397a, 32'h40b1d0f4, 32'h4268277b, 32'h42585478, 32'h429ab8c2, 32'h41f6d883};
test_input[25032:25039] = '{32'h4164a647, 32'hc2b26a87, 32'hc1da0aad, 32'hc2c28f74, 32'hc1b7e006, 32'h41123533, 32'h422ed6ad, 32'hc26bbf02};
test_output[25032:25039] = '{32'h4164a647, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41123533, 32'h422ed6ad, 32'h0};
test_input[25040:25047] = '{32'hc2831dd9, 32'hc286e266, 32'hc1dd71bd, 32'hc25a9bda, 32'hbd370f09, 32'hc28b9513, 32'h42514a94, 32'h4096a843};
test_output[25040:25047] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42514a94, 32'h4096a843};
test_input[25048:25055] = '{32'h42b74be8, 32'hc2980c59, 32'h4261ccfa, 32'hc201a54b, 32'hc10a2232, 32'hc2ad5382, 32'hc27609f4, 32'hc2a18f3c};
test_output[25048:25055] = '{32'h42b74be8, 32'h0, 32'h4261ccfa, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25056:25063] = '{32'h423ebd23, 32'hc10bf1f7, 32'hc2ae361d, 32'h41744b89, 32'h42988bf6, 32'hc2829cb3, 32'h4239e6ec, 32'hc167e595};
test_output[25056:25063] = '{32'h423ebd23, 32'h0, 32'h0, 32'h41744b89, 32'h42988bf6, 32'h0, 32'h4239e6ec, 32'h0};
test_input[25064:25071] = '{32'h422b1d0c, 32'hc208991c, 32'hc297f120, 32'h41dd798f, 32'h42c5b65a, 32'h4220e344, 32'hc2ab4987, 32'h40da483a};
test_output[25064:25071] = '{32'h422b1d0c, 32'h0, 32'h0, 32'h41dd798f, 32'h42c5b65a, 32'h4220e344, 32'h0, 32'h40da483a};
test_input[25072:25079] = '{32'h4222bce7, 32'hc1e80a32, 32'hc2744e92, 32'hc2832475, 32'hc22f3d03, 32'hc17866da, 32'hc2006a6c, 32'hc14b9e75};
test_output[25072:25079] = '{32'h4222bce7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25080:25087] = '{32'hc2910044, 32'hc16c6dea, 32'hc28047e2, 32'hc2944b6d, 32'h4287f9f1, 32'h42741a5d, 32'hc2a43c7b, 32'hc237437d};
test_output[25080:25087] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4287f9f1, 32'h42741a5d, 32'h0, 32'h0};
test_input[25088:25095] = '{32'h421fdcb5, 32'hc22b74b0, 32'h42606b41, 32'hc1c017e1, 32'hc220a38f, 32'hc24485df, 32'hc2ab0db0, 32'hc2bcec97};
test_output[25088:25095] = '{32'h421fdcb5, 32'h0, 32'h42606b41, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25096:25103] = '{32'hc02861cf, 32'hc127eba4, 32'hc218468a, 32'h41bd9f41, 32'h420cc319, 32'hc1a8ad00, 32'hc21ec837, 32'h4299978e};
test_output[25096:25103] = '{32'h0, 32'h0, 32'h0, 32'h41bd9f41, 32'h420cc319, 32'h0, 32'h0, 32'h4299978e};
test_input[25104:25111] = '{32'h40ebb748, 32'h428e62ff, 32'h424ae633, 32'h41ed86d4, 32'h42415881, 32'hc1dfde54, 32'h415ee418, 32'hc2abe96b};
test_output[25104:25111] = '{32'h40ebb748, 32'h428e62ff, 32'h424ae633, 32'h41ed86d4, 32'h42415881, 32'h0, 32'h415ee418, 32'h0};
test_input[25112:25119] = '{32'hc2aeb656, 32'h4264b4fd, 32'h42a54dd2, 32'h42a3c4d1, 32'hc18a423a, 32'hc2adf2a7, 32'h428e7590, 32'hc22c3b91};
test_output[25112:25119] = '{32'h0, 32'h4264b4fd, 32'h42a54dd2, 32'h42a3c4d1, 32'h0, 32'h0, 32'h428e7590, 32'h0};
test_input[25120:25127] = '{32'hc0bf7cbf, 32'hc2b65be9, 32'h429bf171, 32'hc2687ee7, 32'h429a35c6, 32'h4269deef, 32'hc1d1ca68, 32'h4151f287};
test_output[25120:25127] = '{32'h0, 32'h0, 32'h429bf171, 32'h0, 32'h429a35c6, 32'h4269deef, 32'h0, 32'h4151f287};
test_input[25128:25135] = '{32'h429b41af, 32'h41e20cbb, 32'h42b125a9, 32'hc1238a65, 32'h420a6037, 32'h41ef2b18, 32'h420ee6d4, 32'hc2ab8023};
test_output[25128:25135] = '{32'h429b41af, 32'h41e20cbb, 32'h42b125a9, 32'h0, 32'h420a6037, 32'h41ef2b18, 32'h420ee6d4, 32'h0};
test_input[25136:25143] = '{32'h429f9276, 32'hc270c0d8, 32'hc2936f02, 32'hc03ce446, 32'h4077d5f2, 32'hc2416614, 32'hc22230e8, 32'h4278f29f};
test_output[25136:25143] = '{32'h429f9276, 32'h0, 32'h0, 32'h0, 32'h4077d5f2, 32'h0, 32'h0, 32'h4278f29f};
test_input[25144:25151] = '{32'h42a0ff6b, 32'hc25f1c35, 32'hc29faa14, 32'hc265a752, 32'hc2a83be8, 32'h414509cd, 32'hc202e025, 32'h41f29ef6};
test_output[25144:25151] = '{32'h42a0ff6b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h414509cd, 32'h0, 32'h41f29ef6};
test_input[25152:25159] = '{32'hc1e3ceae, 32'hc2ba9da5, 32'h4235e0ea, 32'h42428858, 32'hc070d055, 32'hc2093b61, 32'hc2a18d50, 32'h40fbed2e};
test_output[25152:25159] = '{32'h0, 32'h0, 32'h4235e0ea, 32'h42428858, 32'h0, 32'h0, 32'h0, 32'h40fbed2e};
test_input[25160:25167] = '{32'hc026d5e2, 32'hc1e607a9, 32'h4226a0d5, 32'h421cbcee, 32'hc170a325, 32'hc2785d57, 32'hc19c0d8e, 32'hc1b53a6d};
test_output[25160:25167] = '{32'h0, 32'h0, 32'h4226a0d5, 32'h421cbcee, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25168:25175] = '{32'h4225e59f, 32'hc2b97ee4, 32'hc1ad1609, 32'h4171896c, 32'h42b25edc, 32'hc17fe369, 32'hc20254c3, 32'hc2800d94};
test_output[25168:25175] = '{32'h4225e59f, 32'h0, 32'h0, 32'h4171896c, 32'h42b25edc, 32'h0, 32'h0, 32'h0};
test_input[25176:25183] = '{32'h42b4aaae, 32'h42c60b9e, 32'h41a18c0c, 32'h4295af26, 32'h4193de4a, 32'hc2beb91d, 32'hc2488b40, 32'hc29335fc};
test_output[25176:25183] = '{32'h42b4aaae, 32'h42c60b9e, 32'h41a18c0c, 32'h4295af26, 32'h4193de4a, 32'h0, 32'h0, 32'h0};
test_input[25184:25191] = '{32'h41c65935, 32'hc2b596e2, 32'h41fbb6c4, 32'h420140a4, 32'hc29bd426, 32'h4278d024, 32'hc0805485, 32'hc1ccbaf5};
test_output[25184:25191] = '{32'h41c65935, 32'h0, 32'h41fbb6c4, 32'h420140a4, 32'h0, 32'h4278d024, 32'h0, 32'h0};
test_input[25192:25199] = '{32'h42ac59f8, 32'hc23661b2, 32'h41de108b, 32'h42b250be, 32'h418b6751, 32'hc282f613, 32'hc1c10813, 32'h40929cd2};
test_output[25192:25199] = '{32'h42ac59f8, 32'h0, 32'h41de108b, 32'h42b250be, 32'h418b6751, 32'h0, 32'h0, 32'h40929cd2};
test_input[25200:25207] = '{32'h42bc2d64, 32'h3fc21bfe, 32'h3f8d60e9, 32'h40ba0097, 32'h408030d2, 32'h41a8b3e3, 32'h428a5812, 32'hc2aea347};
test_output[25200:25207] = '{32'h42bc2d64, 32'h3fc21bfe, 32'h3f8d60e9, 32'h40ba0097, 32'h408030d2, 32'h41a8b3e3, 32'h428a5812, 32'h0};
test_input[25208:25215] = '{32'hc287865e, 32'hc246a8dc, 32'h418cc880, 32'hc1dfcf94, 32'hc2c6a1f7, 32'hc23e837e, 32'hc294e10a, 32'h4223cf0f};
test_output[25208:25215] = '{32'h0, 32'h0, 32'h418cc880, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4223cf0f};
test_input[25216:25223] = '{32'h42b39cf9, 32'hc18b6514, 32'h408f77db, 32'hc2960cdc, 32'hc284432c, 32'h42a39348, 32'hc29ad6e2, 32'h4110b3e0};
test_output[25216:25223] = '{32'h42b39cf9, 32'h0, 32'h408f77db, 32'h0, 32'h0, 32'h42a39348, 32'h0, 32'h4110b3e0};
test_input[25224:25231] = '{32'h421b9a19, 32'h4292bf75, 32'h42b5a860, 32'hc08d2969, 32'h419161af, 32'h42a6e31d, 32'hc26a7d41, 32'hc192af16};
test_output[25224:25231] = '{32'h421b9a19, 32'h4292bf75, 32'h42b5a860, 32'h0, 32'h419161af, 32'h42a6e31d, 32'h0, 32'h0};
test_input[25232:25239] = '{32'hc279e821, 32'h425368cd, 32'hc26865a3, 32'h422270d9, 32'h42c3b74d, 32'h424cc3d3, 32'hc29c587a, 32'h4212f7b0};
test_output[25232:25239] = '{32'h0, 32'h425368cd, 32'h0, 32'h422270d9, 32'h42c3b74d, 32'h424cc3d3, 32'h0, 32'h4212f7b0};
test_input[25240:25247] = '{32'h4273447d, 32'hc2b4a459, 32'hc1ff409a, 32'hc2ac9025, 32'h42a6ff36, 32'h425a4173, 32'hbf8aec1e, 32'h423afae6};
test_output[25240:25247] = '{32'h4273447d, 32'h0, 32'h0, 32'h0, 32'h42a6ff36, 32'h425a4173, 32'h0, 32'h423afae6};
test_input[25248:25255] = '{32'hc2afa670, 32'hc2600327, 32'h41b03761, 32'h40a8fe92, 32'h429f4ea2, 32'hc26c3cdb, 32'hc1e92560, 32'h428b253b};
test_output[25248:25255] = '{32'h0, 32'h0, 32'h41b03761, 32'h40a8fe92, 32'h429f4ea2, 32'h0, 32'h0, 32'h428b253b};
test_input[25256:25263] = '{32'h426c714c, 32'hc1bbae03, 32'hc28eecda, 32'h411a8d80, 32'hc2a75d52, 32'h4223d63a, 32'hc185d53f, 32'hc28e8488};
test_output[25256:25263] = '{32'h426c714c, 32'h0, 32'h0, 32'h411a8d80, 32'h0, 32'h4223d63a, 32'h0, 32'h0};
test_input[25264:25271] = '{32'hc28d4976, 32'hc2b72944, 32'hc2a9f51f, 32'hc2570c82, 32'hc29379a5, 32'hc28ba6ff, 32'hc1cfe51b, 32'h4217c9a5};
test_output[25264:25271] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4217c9a5};
test_input[25272:25279] = '{32'hc164a11b, 32'h42a2845c, 32'hc2552c64, 32'hc2468d02, 32'hc2aa2357, 32'h42b76f0e, 32'h42392494, 32'hc1e98b96};
test_output[25272:25279] = '{32'h0, 32'h42a2845c, 32'h0, 32'h0, 32'h0, 32'h42b76f0e, 32'h42392494, 32'h0};
test_input[25280:25287] = '{32'hc19a240d, 32'hc14e79cf, 32'h42c5af16, 32'h42331c55, 32'hc1b094e4, 32'h42008fdd, 32'hc2c518fc, 32'h42273cad};
test_output[25280:25287] = '{32'h0, 32'h0, 32'h42c5af16, 32'h42331c55, 32'h0, 32'h42008fdd, 32'h0, 32'h42273cad};
test_input[25288:25295] = '{32'h42763169, 32'hbebeb926, 32'hc2c04fe1, 32'hc2c2650b, 32'hc1b2accb, 32'h429e68c5, 32'hc276cd03, 32'h42217ee7};
test_output[25288:25295] = '{32'h42763169, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429e68c5, 32'h0, 32'h42217ee7};
test_input[25296:25303] = '{32'hc003a6e7, 32'hc0e93247, 32'h42005bbc, 32'h3ece935a, 32'hc29a702f, 32'hc2c50010, 32'h413fdf20, 32'hc241b182};
test_output[25296:25303] = '{32'h0, 32'h0, 32'h42005bbc, 32'h3ece935a, 32'h0, 32'h0, 32'h413fdf20, 32'h0};
test_input[25304:25311] = '{32'hc2b0169d, 32'h41e3b373, 32'hc2b77bdb, 32'h422deacb, 32'h429ffabf, 32'h41737ae1, 32'h41bb4cf6, 32'h421ed304};
test_output[25304:25311] = '{32'h0, 32'h41e3b373, 32'h0, 32'h422deacb, 32'h429ffabf, 32'h41737ae1, 32'h41bb4cf6, 32'h421ed304};
test_input[25312:25319] = '{32'hc291db11, 32'hc2599ec4, 32'hc29e9e7f, 32'hc1fc510b, 32'h40fa192d, 32'hc1d0c2c1, 32'h40e7692e, 32'h4271be6b};
test_output[25312:25319] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40fa192d, 32'h0, 32'h40e7692e, 32'h4271be6b};
test_input[25320:25327] = '{32'hc2bce3fd, 32'hbfe593f6, 32'h41f49210, 32'h42b1911b, 32'hbf999cca, 32'h42bc0a45, 32'h419cd32f, 32'hc24e8a97};
test_output[25320:25327] = '{32'h0, 32'h0, 32'h41f49210, 32'h42b1911b, 32'h0, 32'h42bc0a45, 32'h419cd32f, 32'h0};
test_input[25328:25335] = '{32'h42858643, 32'h410435b9, 32'h42b0f544, 32'h428160aa, 32'h41c83b51, 32'hc10e733b, 32'h42bb496d, 32'h42049832};
test_output[25328:25335] = '{32'h42858643, 32'h410435b9, 32'h42b0f544, 32'h428160aa, 32'h41c83b51, 32'h0, 32'h42bb496d, 32'h42049832};
test_input[25336:25343] = '{32'h41bc18fd, 32'h4281e589, 32'hc189a646, 32'hc23bf00b, 32'hc2641e74, 32'h40b8a2a4, 32'hc23cf42f, 32'hc28f30a6};
test_output[25336:25343] = '{32'h41bc18fd, 32'h4281e589, 32'h0, 32'h0, 32'h0, 32'h40b8a2a4, 32'h0, 32'h0};
test_input[25344:25351] = '{32'hc2a03250, 32'h427c843c, 32'h422f5496, 32'hbedc6cd1, 32'hc23782f9, 32'hc1cbee87, 32'hc2246a9f, 32'h42404b59};
test_output[25344:25351] = '{32'h0, 32'h427c843c, 32'h422f5496, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42404b59};
test_input[25352:25359] = '{32'hc22141ed, 32'h4156096c, 32'hc2a2ec49, 32'hc28fdfcd, 32'h42223bbd, 32'hc22e98f8, 32'hc2b975fb, 32'h42bf77a2};
test_output[25352:25359] = '{32'h0, 32'h4156096c, 32'h0, 32'h0, 32'h42223bbd, 32'h0, 32'h0, 32'h42bf77a2};
test_input[25360:25367] = '{32'h416167ae, 32'h41402f76, 32'hc236494a, 32'h42a7e5a8, 32'hc0a312ba, 32'h4287ba84, 32'h42c73c62, 32'hc28acb27};
test_output[25360:25367] = '{32'h416167ae, 32'h41402f76, 32'h0, 32'h42a7e5a8, 32'h0, 32'h4287ba84, 32'h42c73c62, 32'h0};
test_input[25368:25375] = '{32'h41891ff6, 32'hc2c4147d, 32'hc2c18f6a, 32'hc272a029, 32'h422856c4, 32'hc0cdd756, 32'hc11e1f06, 32'h42b2c84d};
test_output[25368:25375] = '{32'h41891ff6, 32'h0, 32'h0, 32'h0, 32'h422856c4, 32'h0, 32'h0, 32'h42b2c84d};
test_input[25376:25383] = '{32'h426c3598, 32'h4266f26f, 32'hc2219b5d, 32'h42af365c, 32'hc06f0414, 32'h41badcb3, 32'h428b5a0e, 32'h4275c7de};
test_output[25376:25383] = '{32'h426c3598, 32'h4266f26f, 32'h0, 32'h42af365c, 32'h0, 32'h41badcb3, 32'h428b5a0e, 32'h4275c7de};
test_input[25384:25391] = '{32'h41cf4dc1, 32'h4169c633, 32'hc2c07370, 32'hc27308b3, 32'h422327bf, 32'h4123291c, 32'hc20aafaf, 32'hc259661d};
test_output[25384:25391] = '{32'h41cf4dc1, 32'h4169c633, 32'h0, 32'h0, 32'h422327bf, 32'h4123291c, 32'h0, 32'h0};
test_input[25392:25399] = '{32'h4225a0be, 32'h41932159, 32'h421044ab, 32'h427a0265, 32'hc2150b0c, 32'hc134ec1a, 32'hc1adb566, 32'hc261d344};
test_output[25392:25399] = '{32'h4225a0be, 32'h41932159, 32'h421044ab, 32'h427a0265, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25400:25407] = '{32'hc157aed0, 32'h4209aab5, 32'h42c12598, 32'hc11124e7, 32'hc297255d, 32'hc2afddf2, 32'h42a18718, 32'hc2a0bcb7};
test_output[25400:25407] = '{32'h0, 32'h4209aab5, 32'h42c12598, 32'h0, 32'h0, 32'h0, 32'h42a18718, 32'h0};
test_input[25408:25415] = '{32'hc2758e21, 32'h41309e13, 32'hc22ec38c, 32'h42279b02, 32'h41aa3a17, 32'h4197d965, 32'hc166ccf1, 32'hc2799f36};
test_output[25408:25415] = '{32'h0, 32'h41309e13, 32'h0, 32'h42279b02, 32'h41aa3a17, 32'h4197d965, 32'h0, 32'h0};
test_input[25416:25423] = '{32'h42b7ba37, 32'hc233a339, 32'h423a5c87, 32'hc223cd87, 32'h41f93d64, 32'hc29f11bc, 32'hc15ee9f1, 32'h429d9739};
test_output[25416:25423] = '{32'h42b7ba37, 32'h0, 32'h423a5c87, 32'h0, 32'h41f93d64, 32'h0, 32'h0, 32'h429d9739};
test_input[25424:25431] = '{32'h4285408f, 32'hc291911a, 32'h41bf0683, 32'hc2c5707e, 32'h427621e3, 32'h429cb609, 32'h4198a481, 32'hc1d4c329};
test_output[25424:25431] = '{32'h4285408f, 32'h0, 32'h41bf0683, 32'h0, 32'h427621e3, 32'h429cb609, 32'h4198a481, 32'h0};
test_input[25432:25439] = '{32'h4178b5a4, 32'h42b9e9e1, 32'h423c3521, 32'hc1881f5b, 32'h4292e6af, 32'h42160e95, 32'hc267c62f, 32'hc242f7f5};
test_output[25432:25439] = '{32'h4178b5a4, 32'h42b9e9e1, 32'h423c3521, 32'h0, 32'h4292e6af, 32'h42160e95, 32'h0, 32'h0};
test_input[25440:25447] = '{32'hc1ad99e7, 32'hc1da1d87, 32'h42c0d7e5, 32'hc236fefb, 32'h411aae4c, 32'h42b17bd7, 32'h422ea159, 32'hc23a0dfd};
test_output[25440:25447] = '{32'h0, 32'h0, 32'h42c0d7e5, 32'h0, 32'h411aae4c, 32'h42b17bd7, 32'h422ea159, 32'h0};
test_input[25448:25455] = '{32'h42a66ec4, 32'h42c6f10c, 32'hc1b4aebe, 32'hc28fcac3, 32'hc24c883a, 32'h427a3d66, 32'hc2aeaa17, 32'hc1563883};
test_output[25448:25455] = '{32'h42a66ec4, 32'h42c6f10c, 32'h0, 32'h0, 32'h0, 32'h427a3d66, 32'h0, 32'h0};
test_input[25456:25463] = '{32'h42b8b488, 32'hc266ef5c, 32'h4265a644, 32'h418dd832, 32'hc271c93f, 32'h426acaab, 32'hc11d5f94, 32'h42a25a6a};
test_output[25456:25463] = '{32'h42b8b488, 32'h0, 32'h4265a644, 32'h418dd832, 32'h0, 32'h426acaab, 32'h0, 32'h42a25a6a};
test_input[25464:25471] = '{32'hc20c05ce, 32'h41d3b032, 32'hc27ba733, 32'hc19d4b5b, 32'h40f452c6, 32'h42322492, 32'h4247d056, 32'h406d8e0e};
test_output[25464:25471] = '{32'h0, 32'h41d3b032, 32'h0, 32'h0, 32'h40f452c6, 32'h42322492, 32'h4247d056, 32'h406d8e0e};
test_input[25472:25479] = '{32'h42c3b1a4, 32'hc2b8ae27, 32'h42ad1918, 32'hc2978391, 32'h40e2c27a, 32'h41d010e4, 32'h40d27ec5, 32'h4295b9c8};
test_output[25472:25479] = '{32'h42c3b1a4, 32'h0, 32'h42ad1918, 32'h0, 32'h40e2c27a, 32'h41d010e4, 32'h40d27ec5, 32'h4295b9c8};
test_input[25480:25487] = '{32'hc15d7531, 32'hc1820fde, 32'h4196614e, 32'h42099a83, 32'h42a990c4, 32'h428b4bf5, 32'h421d8a7c, 32'hc2b5b9a0};
test_output[25480:25487] = '{32'h0, 32'h0, 32'h4196614e, 32'h42099a83, 32'h42a990c4, 32'h428b4bf5, 32'h421d8a7c, 32'h0};
test_input[25488:25495] = '{32'h42aea392, 32'hc1553741, 32'hc2c574b6, 32'hc2ad29ce, 32'h426f16be, 32'h4231e2f7, 32'hc27284a8, 32'h41c64af9};
test_output[25488:25495] = '{32'h42aea392, 32'h0, 32'h0, 32'h0, 32'h426f16be, 32'h4231e2f7, 32'h0, 32'h41c64af9};
test_input[25496:25503] = '{32'h42b06353, 32'hc2b51d7a, 32'h42899b58, 32'h412762bf, 32'h4284539d, 32'hc1948280, 32'hc28dda6a, 32'hc1885109};
test_output[25496:25503] = '{32'h42b06353, 32'h0, 32'h42899b58, 32'h412762bf, 32'h4284539d, 32'h0, 32'h0, 32'h0};
test_input[25504:25511] = '{32'hc1021826, 32'h4282b11a, 32'hc2a8b2b2, 32'h4281a60c, 32'hc266cdca, 32'hc1bb253e, 32'hc24b676f, 32'hc260edd0};
test_output[25504:25511] = '{32'h0, 32'h4282b11a, 32'h0, 32'h4281a60c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25512:25519] = '{32'hc28b395f, 32'hc247d2de, 32'h428ea821, 32'hc17c9060, 32'h4207d9bf, 32'h41aaabaf, 32'hc26b3897, 32'hc22e23db};
test_output[25512:25519] = '{32'h0, 32'h0, 32'h428ea821, 32'h0, 32'h4207d9bf, 32'h41aaabaf, 32'h0, 32'h0};
test_input[25520:25527] = '{32'h42b7f3d3, 32'hc29951cf, 32'h4233e497, 32'hc2401e6e, 32'hc24ce23c, 32'h425f2e2c, 32'h42c71419, 32'h40f24387};
test_output[25520:25527] = '{32'h42b7f3d3, 32'h0, 32'h4233e497, 32'h0, 32'h0, 32'h425f2e2c, 32'h42c71419, 32'h40f24387};
test_input[25528:25535] = '{32'h428645c2, 32'hc288d8ea, 32'hc298d963, 32'hc2b8aa7a, 32'hc2803e6f, 32'hc24d5933, 32'h4282b38f, 32'h42922998};
test_output[25528:25535] = '{32'h428645c2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4282b38f, 32'h42922998};
test_input[25536:25543] = '{32'hc106a370, 32'hc1aaa245, 32'hc2068236, 32'h4215888f, 32'hc297fa86, 32'h426396fa, 32'h4079f003, 32'hc28e6dee};
test_output[25536:25543] = '{32'h0, 32'h0, 32'h0, 32'h4215888f, 32'h0, 32'h426396fa, 32'h4079f003, 32'h0};
test_input[25544:25551] = '{32'h41135002, 32'hc1400a51, 32'hc1dd86b1, 32'h42698b47, 32'h423b552f, 32'h4293b52d, 32'h42ad6bb1, 32'h42886b95};
test_output[25544:25551] = '{32'h41135002, 32'h0, 32'h0, 32'h42698b47, 32'h423b552f, 32'h4293b52d, 32'h42ad6bb1, 32'h42886b95};
test_input[25552:25559] = '{32'hc13eb369, 32'h42b47825, 32'hc1ff33e9, 32'hc1b11e61, 32'hc155d890, 32'h416888b9, 32'h41e815ef, 32'h429bbc00};
test_output[25552:25559] = '{32'h0, 32'h42b47825, 32'h0, 32'h0, 32'h0, 32'h416888b9, 32'h41e815ef, 32'h429bbc00};
test_input[25560:25567] = '{32'hc1c46bfe, 32'h4263ae80, 32'h4254b14a, 32'h412cf01c, 32'hc29d5bfa, 32'h4287f4a8, 32'h428e2880, 32'hc219e526};
test_output[25560:25567] = '{32'h0, 32'h4263ae80, 32'h4254b14a, 32'h412cf01c, 32'h0, 32'h4287f4a8, 32'h428e2880, 32'h0};
test_input[25568:25575] = '{32'h4280060b, 32'hc2156daf, 32'hc2c72389, 32'hc279db92, 32'hc2bcf507, 32'hc2021c73, 32'h42823924, 32'h41c3b7aa};
test_output[25568:25575] = '{32'h4280060b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42823924, 32'h41c3b7aa};
test_input[25576:25583] = '{32'hc2066064, 32'hc28f478b, 32'hc1801b7c, 32'hc1c07c98, 32'h42aae9ba, 32'h4299bfee, 32'h41c9fb38, 32'hc20f4af4};
test_output[25576:25583] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42aae9ba, 32'h4299bfee, 32'h41c9fb38, 32'h0};
test_input[25584:25591] = '{32'hc29b3e40, 32'hc2a3fda6, 32'hc28f2262, 32'hc2b08c4f, 32'h4208eda7, 32'hc286ca32, 32'h42b5048f, 32'h426b1a04};
test_output[25584:25591] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4208eda7, 32'h0, 32'h42b5048f, 32'h426b1a04};
test_input[25592:25599] = '{32'h41808ad5, 32'h420a2555, 32'hc22a7e3f, 32'h41c20932, 32'h41faa157, 32'hc1554626, 32'hc2ae10ce, 32'hc23c3b44};
test_output[25592:25599] = '{32'h41808ad5, 32'h420a2555, 32'h0, 32'h41c20932, 32'h41faa157, 32'h0, 32'h0, 32'h0};
test_input[25600:25607] = '{32'h4285dd1d, 32'h4280bda0, 32'h42682d0f, 32'hc2960988, 32'hc22d3b3d, 32'h4261c670, 32'h4201ff64, 32'h41b403d8};
test_output[25600:25607] = '{32'h4285dd1d, 32'h4280bda0, 32'h42682d0f, 32'h0, 32'h0, 32'h4261c670, 32'h4201ff64, 32'h41b403d8};
test_input[25608:25615] = '{32'hc18e4287, 32'h42c64e4d, 32'hc2abdfc4, 32'h40f4a01a, 32'h42a3781c, 32'hc22363d2, 32'h423e4789, 32'hc2a20b1a};
test_output[25608:25615] = '{32'h0, 32'h42c64e4d, 32'h0, 32'h40f4a01a, 32'h42a3781c, 32'h0, 32'h423e4789, 32'h0};
test_input[25616:25623] = '{32'hc13a77c1, 32'hc13d37ef, 32'h411f0c80, 32'hc228f0db, 32'hc1523bc4, 32'hc2221bdb, 32'hc1eb6b00, 32'h42664cf6};
test_output[25616:25623] = '{32'h0, 32'h0, 32'h411f0c80, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42664cf6};
test_input[25624:25631] = '{32'hc2bd3d32, 32'hc2a83d66, 32'h41bdbf0d, 32'hc2c7c41f, 32'hc2826018, 32'hc1a214a1, 32'h4227a215, 32'hc20bfe37};
test_output[25624:25631] = '{32'h0, 32'h0, 32'h41bdbf0d, 32'h0, 32'h0, 32'h0, 32'h4227a215, 32'h0};
test_input[25632:25639] = '{32'h42813823, 32'hc20ee9c3, 32'h408598a8, 32'hc2306f52, 32'h423fedef, 32'h4272e1b2, 32'hc283560d, 32'hc12509a6};
test_output[25632:25639] = '{32'h42813823, 32'h0, 32'h408598a8, 32'h0, 32'h423fedef, 32'h4272e1b2, 32'h0, 32'h0};
test_input[25640:25647] = '{32'h429c4b6c, 32'h428f9495, 32'h405c4612, 32'hc14a2748, 32'h3fd5c1ea, 32'h4127b4fe, 32'h41a6147e, 32'h4299abed};
test_output[25640:25647] = '{32'h429c4b6c, 32'h428f9495, 32'h405c4612, 32'h0, 32'h3fd5c1ea, 32'h4127b4fe, 32'h41a6147e, 32'h4299abed};
test_input[25648:25655] = '{32'hc00defc2, 32'hc2c72ce9, 32'h429ad97b, 32'h42052fa8, 32'h42b37006, 32'h42b926f4, 32'hbeb6101a, 32'hc0a7e0c2};
test_output[25648:25655] = '{32'h0, 32'h0, 32'h429ad97b, 32'h42052fa8, 32'h42b37006, 32'h42b926f4, 32'h0, 32'h0};
test_input[25656:25663] = '{32'h3ffffaa6, 32'hc0cc7596, 32'hc2ba363b, 32'hc0db45af, 32'h414c6854, 32'h427c9dd4, 32'hc2a0872e, 32'h429b559c};
test_output[25656:25663] = '{32'h3ffffaa6, 32'h0, 32'h0, 32'h0, 32'h414c6854, 32'h427c9dd4, 32'h0, 32'h429b559c};
test_input[25664:25671] = '{32'hc2a1e509, 32'hc279b2b9, 32'h424f19b1, 32'h42acc2d8, 32'hc295a5ae, 32'hc1716d80, 32'hc0aa9815, 32'h409b4824};
test_output[25664:25671] = '{32'h0, 32'h0, 32'h424f19b1, 32'h42acc2d8, 32'h0, 32'h0, 32'h0, 32'h409b4824};
test_input[25672:25679] = '{32'hc18249f5, 32'hc294cb34, 32'h4116553c, 32'hc1b29c16, 32'h423faffe, 32'h4269d441, 32'h428a29d4, 32'h422cb4b9};
test_output[25672:25679] = '{32'h0, 32'h0, 32'h4116553c, 32'h0, 32'h423faffe, 32'h4269d441, 32'h428a29d4, 32'h422cb4b9};
test_input[25680:25687] = '{32'h427a0e17, 32'hc2afef11, 32'hc226d07b, 32'h4278b671, 32'hc1ecf5af, 32'hc1e70d40, 32'hc2100346, 32'h429ee53a};
test_output[25680:25687] = '{32'h427a0e17, 32'h0, 32'h0, 32'h4278b671, 32'h0, 32'h0, 32'h0, 32'h429ee53a};
test_input[25688:25695] = '{32'hc2a8d2e1, 32'h4228c540, 32'h42c1423d, 32'h429f73d7, 32'h41fc0522, 32'hc200b734, 32'h421bdb4c, 32'h41b514ef};
test_output[25688:25695] = '{32'h0, 32'h4228c540, 32'h42c1423d, 32'h429f73d7, 32'h41fc0522, 32'h0, 32'h421bdb4c, 32'h41b514ef};
test_input[25696:25703] = '{32'h418f823d, 32'h4258a0fb, 32'hc24c9f54, 32'hc27d3c87, 32'h419fcfbf, 32'hc10341b5, 32'hc24adaf4, 32'hc2a54d39};
test_output[25696:25703] = '{32'h418f823d, 32'h4258a0fb, 32'h0, 32'h0, 32'h419fcfbf, 32'h0, 32'h0, 32'h0};
test_input[25704:25711] = '{32'h4202f0ac, 32'h420bc4e7, 32'h42a6a7bf, 32'h42a86605, 32'hc12239f8, 32'h4117a554, 32'h4280a58d, 32'hc0a6214f};
test_output[25704:25711] = '{32'h4202f0ac, 32'h420bc4e7, 32'h42a6a7bf, 32'h42a86605, 32'h0, 32'h4117a554, 32'h4280a58d, 32'h0};
test_input[25712:25719] = '{32'hc1a128f3, 32'hc0d041e7, 32'hc12c7bfc, 32'h42c6b3c5, 32'h40a0acf7, 32'hc0a9455e, 32'h428c64fc, 32'h4232dd71};
test_output[25712:25719] = '{32'h0, 32'h0, 32'h0, 32'h42c6b3c5, 32'h40a0acf7, 32'h0, 32'h428c64fc, 32'h4232dd71};
test_input[25720:25727] = '{32'hc23a2c7d, 32'h42bf2aff, 32'h42927216, 32'h42450d4c, 32'hc246d94e, 32'hc286fdd8, 32'hc244700f, 32'hc2c76d8b};
test_output[25720:25727] = '{32'h0, 32'h42bf2aff, 32'h42927216, 32'h42450d4c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25728:25735] = '{32'h40d39531, 32'h4276fc7b, 32'hc1e0c9cd, 32'h428ac7fe, 32'h41f93cf4, 32'hc264bd4f, 32'h42807991, 32'h42bca65a};
test_output[25728:25735] = '{32'h40d39531, 32'h4276fc7b, 32'h0, 32'h428ac7fe, 32'h41f93cf4, 32'h0, 32'h42807991, 32'h42bca65a};
test_input[25736:25743] = '{32'h42685fd8, 32'hc2594454, 32'hc20a4146, 32'hc2a1a22d, 32'h427d30b1, 32'h400fa9de, 32'h40b1c5a9, 32'hc2918758};
test_output[25736:25743] = '{32'h42685fd8, 32'h0, 32'h0, 32'h0, 32'h427d30b1, 32'h400fa9de, 32'h40b1c5a9, 32'h0};
test_input[25744:25751] = '{32'h41dbf9ed, 32'hc24eadf0, 32'hc15af392, 32'h428a6e45, 32'h41c071d3, 32'hc2203679, 32'hc231b618, 32'hc26f4264};
test_output[25744:25751] = '{32'h41dbf9ed, 32'h0, 32'h0, 32'h428a6e45, 32'h41c071d3, 32'h0, 32'h0, 32'h0};
test_input[25752:25759] = '{32'hc29328c4, 32'hc2a00410, 32'h42a8633c, 32'h427a60f1, 32'hc264d3c8, 32'hc2872d4d, 32'h429232ee, 32'h4222fdc6};
test_output[25752:25759] = '{32'h0, 32'h0, 32'h42a8633c, 32'h427a60f1, 32'h0, 32'h0, 32'h429232ee, 32'h4222fdc6};
test_input[25760:25767] = '{32'h42069e44, 32'hc200985f, 32'hc2923a5e, 32'h42c19c8f, 32'hc29ff238, 32'h42c0322c, 32'h41fb3e96, 32'h4283ceb9};
test_output[25760:25767] = '{32'h42069e44, 32'h0, 32'h0, 32'h42c19c8f, 32'h0, 32'h42c0322c, 32'h41fb3e96, 32'h4283ceb9};
test_input[25768:25775] = '{32'h42589ae5, 32'hbe879346, 32'h41eb37fa, 32'hc281396a, 32'h4271b507, 32'h429a6db3, 32'hc1b87f95, 32'hc1f55b43};
test_output[25768:25775] = '{32'h42589ae5, 32'h0, 32'h41eb37fa, 32'h0, 32'h4271b507, 32'h429a6db3, 32'h0, 32'h0};
test_input[25776:25783] = '{32'hc2508ad5, 32'h42ba21f3, 32'h42896fad, 32'h42679707, 32'hc285d33f, 32'hc1e36661, 32'hbfa7a254, 32'h421821e1};
test_output[25776:25783] = '{32'h0, 32'h42ba21f3, 32'h42896fad, 32'h42679707, 32'h0, 32'h0, 32'h0, 32'h421821e1};
test_input[25784:25791] = '{32'hc2ace426, 32'hc26a26c1, 32'hc2b49990, 32'h4154d29c, 32'h41fa5dff, 32'h428da76b, 32'h411b31b4, 32'h428003cd};
test_output[25784:25791] = '{32'h0, 32'h0, 32'h0, 32'h4154d29c, 32'h41fa5dff, 32'h428da76b, 32'h411b31b4, 32'h428003cd};
test_input[25792:25799] = '{32'h429de059, 32'h42a42055, 32'h4028b016, 32'hc0c8b24c, 32'h411e16fc, 32'h421d3213, 32'hc2b33874, 32'hc2a90f92};
test_output[25792:25799] = '{32'h429de059, 32'h42a42055, 32'h4028b016, 32'h0, 32'h411e16fc, 32'h421d3213, 32'h0, 32'h0};
test_input[25800:25807] = '{32'hc1f98eb4, 32'hc291b953, 32'h429bab94, 32'hc285bc37, 32'hc0ed36a7, 32'h4285d4bb, 32'h425a71b9, 32'hc06b55a4};
test_output[25800:25807] = '{32'h0, 32'h0, 32'h429bab94, 32'h0, 32'h0, 32'h4285d4bb, 32'h425a71b9, 32'h0};
test_input[25808:25815] = '{32'hc246a243, 32'h4243aa9b, 32'h428a7c00, 32'hc2b17cce, 32'hc0178d97, 32'h40c74148, 32'hc2871852, 32'hc2061f9a};
test_output[25808:25815] = '{32'h0, 32'h4243aa9b, 32'h428a7c00, 32'h0, 32'h0, 32'h40c74148, 32'h0, 32'h0};
test_input[25816:25823] = '{32'h423c43ba, 32'h421fdb83, 32'h42601ccb, 32'hc2a80199, 32'h42b23d9b, 32'hc2aff5b5, 32'hc21b4b3b, 32'h42b82ab1};
test_output[25816:25823] = '{32'h423c43ba, 32'h421fdb83, 32'h42601ccb, 32'h0, 32'h42b23d9b, 32'h0, 32'h0, 32'h42b82ab1};
test_input[25824:25831] = '{32'hc2a784aa, 32'h4214e6d5, 32'h42c33af2, 32'hc2ae8c21, 32'hc1c66976, 32'h429188cd, 32'hc1c7fea4, 32'hc153dce0};
test_output[25824:25831] = '{32'h0, 32'h4214e6d5, 32'h42c33af2, 32'h0, 32'h0, 32'h429188cd, 32'h0, 32'h0};
test_input[25832:25839] = '{32'hc1c928bf, 32'hc12809c7, 32'hc25f4ac6, 32'h422c4a00, 32'hc2804e65, 32'hc21ffcff, 32'hc24e5d9f, 32'hc21cffff};
test_output[25832:25839] = '{32'h0, 32'h0, 32'h0, 32'h422c4a00, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25840:25847] = '{32'hc2b941c4, 32'h4213b5b2, 32'h4291ef6f, 32'hc2b2c7ae, 32'hc1991cd8, 32'hc189aa53, 32'hc1712346, 32'h4293f60f};
test_output[25840:25847] = '{32'h0, 32'h4213b5b2, 32'h4291ef6f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4293f60f};
test_input[25848:25855] = '{32'hc267b4d2, 32'hc2959cea, 32'hc2893c92, 32'h42a0c8a1, 32'hc2bcc968, 32'h428ff6a8, 32'hc183d6b8, 32'hc281517c};
test_output[25848:25855] = '{32'h0, 32'h0, 32'h0, 32'h42a0c8a1, 32'h0, 32'h428ff6a8, 32'h0, 32'h0};
test_input[25856:25863] = '{32'hc1ef97bc, 32'h42bb7736, 32'h42457b32, 32'h42b062cd, 32'h42818f83, 32'h4188a280, 32'h428d088e, 32'h4296e4f2};
test_output[25856:25863] = '{32'h0, 32'h42bb7736, 32'h42457b32, 32'h42b062cd, 32'h42818f83, 32'h4188a280, 32'h428d088e, 32'h4296e4f2};
test_input[25864:25871] = '{32'h4199a5ad, 32'hc0c22265, 32'h41550923, 32'hc247bbc6, 32'h4297865c, 32'h42a4db2b, 32'hc266887c, 32'h428afd3f};
test_output[25864:25871] = '{32'h4199a5ad, 32'h0, 32'h41550923, 32'h0, 32'h4297865c, 32'h42a4db2b, 32'h0, 32'h428afd3f};
test_input[25872:25879] = '{32'hc2aa070d, 32'hc23b569e, 32'hc2bf4917, 32'hc259454a, 32'hc274fe95, 32'h42931787, 32'hc1cf3213, 32'h41b8858f};
test_output[25872:25879] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42931787, 32'h0, 32'h41b8858f};
test_input[25880:25887] = '{32'h4210590a, 32'h40d03a62, 32'h42a60aa9, 32'h42215474, 32'h426063e1, 32'h41de5ffc, 32'hc2a1fd6a, 32'h40942fad};
test_output[25880:25887] = '{32'h4210590a, 32'h40d03a62, 32'h42a60aa9, 32'h42215474, 32'h426063e1, 32'h41de5ffc, 32'h0, 32'h40942fad};
test_input[25888:25895] = '{32'hc23add22, 32'hc0c14225, 32'hc286bc30, 32'h429f0ac7, 32'h4090b53a, 32'h42635093, 32'hc17df6eb, 32'hc10f7f42};
test_output[25888:25895] = '{32'h0, 32'h0, 32'h0, 32'h429f0ac7, 32'h4090b53a, 32'h42635093, 32'h0, 32'h0};
test_input[25896:25903] = '{32'hc217ae8f, 32'h421533b0, 32'h4204df44, 32'hbee438cc, 32'hc25737e8, 32'h41bf613c, 32'hc22426a6, 32'hc1735cd3};
test_output[25896:25903] = '{32'h0, 32'h421533b0, 32'h4204df44, 32'h0, 32'h0, 32'h41bf613c, 32'h0, 32'h0};
test_input[25904:25911] = '{32'h42a05580, 32'hc2adfa15, 32'h4273dfc4, 32'hc2b1d62d, 32'hc2aa4947, 32'h41827cd9, 32'hc0b80529, 32'h4130115b};
test_output[25904:25911] = '{32'h42a05580, 32'h0, 32'h4273dfc4, 32'h0, 32'h0, 32'h41827cd9, 32'h0, 32'h4130115b};
test_input[25912:25919] = '{32'hc25759e9, 32'hc2c279ea, 32'h41b26c08, 32'h41c66709, 32'hc2bfcdb3, 32'hc1111bf7, 32'h41b164a5, 32'hc0eb9ed6};
test_output[25912:25919] = '{32'h0, 32'h0, 32'h41b26c08, 32'h41c66709, 32'h0, 32'h0, 32'h41b164a5, 32'h0};
test_input[25920:25927] = '{32'h42968b6e, 32'h42a97eab, 32'hc2334503, 32'hc298a742, 32'h42735e07, 32'hc1b7eb2c, 32'hc0cd03a6, 32'h405cc1e0};
test_output[25920:25927] = '{32'h42968b6e, 32'h42a97eab, 32'h0, 32'h0, 32'h42735e07, 32'h0, 32'h0, 32'h405cc1e0};
test_input[25928:25935] = '{32'hc2a4c6f0, 32'h418a4f3e, 32'hc1b90a5f, 32'hc2248531, 32'hc188f5cb, 32'hc24ef844, 32'hc22d15aa, 32'hc1f75131};
test_output[25928:25935] = '{32'h0, 32'h418a4f3e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25936:25943] = '{32'hc116f1fb, 32'h42736e08, 32'hc178e309, 32'h42af24dc, 32'hc2a0c967, 32'h418644a4, 32'h42aa1f7b, 32'h42b28dd2};
test_output[25936:25943] = '{32'h0, 32'h42736e08, 32'h0, 32'h42af24dc, 32'h0, 32'h418644a4, 32'h42aa1f7b, 32'h42b28dd2};
test_input[25944:25951] = '{32'h4260f0bc, 32'h429159e5, 32'h425bd114, 32'h428011d7, 32'hc27887e6, 32'hc23a38d5, 32'h4237037a, 32'hc2a66c62};
test_output[25944:25951] = '{32'h4260f0bc, 32'h429159e5, 32'h425bd114, 32'h428011d7, 32'h0, 32'h0, 32'h4237037a, 32'h0};
test_input[25952:25959] = '{32'hc1e54233, 32'h427b766e, 32'hc251f6fd, 32'hc2c1c773, 32'hc1563da4, 32'hc26863ad, 32'h42b3a4a5, 32'hc28d5d32};
test_output[25952:25959] = '{32'h0, 32'h427b766e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b3a4a5, 32'h0};
test_input[25960:25967] = '{32'h41ae2b9f, 32'hc199cd5b, 32'hc2c37e62, 32'hc2a48928, 32'hc2c72151, 32'hc1d95e8d, 32'h42895c5c, 32'hc26b206c};
test_output[25960:25967] = '{32'h41ae2b9f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42895c5c, 32'h0};
test_input[25968:25975] = '{32'h42ba1794, 32'hc2969c30, 32'hc2c34be6, 32'h42954430, 32'hc24a8618, 32'h42c1e38a, 32'hc2a243df, 32'hc2642c2b};
test_output[25968:25975] = '{32'h42ba1794, 32'h0, 32'h0, 32'h42954430, 32'h0, 32'h42c1e38a, 32'h0, 32'h0};
test_input[25976:25983] = '{32'h42973546, 32'hc23470ef, 32'h42c23ce7, 32'h42899b03, 32'hbfa4355b, 32'hc2251631, 32'hc1b762e6, 32'hc2856b1a};
test_output[25976:25983] = '{32'h42973546, 32'h0, 32'h42c23ce7, 32'h42899b03, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25984:25991] = '{32'hc1c56803, 32'h42ad5ec4, 32'h42804ae6, 32'h42a0107a, 32'hc2597933, 32'hc249ca04, 32'h42293d0c, 32'h41f90914};
test_output[25984:25991] = '{32'h0, 32'h42ad5ec4, 32'h42804ae6, 32'h42a0107a, 32'h0, 32'h0, 32'h42293d0c, 32'h41f90914};
test_input[25992:25999] = '{32'hc28e3941, 32'h42c5d983, 32'hc1b05b8f, 32'h42b2c373, 32'hc24de674, 32'h4286799e, 32'h424b8ee9, 32'hc2256088};
test_output[25992:25999] = '{32'h0, 32'h42c5d983, 32'h0, 32'h42b2c373, 32'h0, 32'h4286799e, 32'h424b8ee9, 32'h0};
test_input[26000:26007] = '{32'hc2abe791, 32'h42804b8d, 32'hc14b0338, 32'hc2c431f0, 32'h428a8ce9, 32'h41847724, 32'h42ab6888, 32'hc2871280};
test_output[26000:26007] = '{32'h0, 32'h42804b8d, 32'h0, 32'h0, 32'h428a8ce9, 32'h41847724, 32'h42ab6888, 32'h0};
test_input[26008:26015] = '{32'h42114ee5, 32'h42aef416, 32'hc297e3b4, 32'hc1b8d6ce, 32'hc1f06b55, 32'hc2aa296a, 32'hc2bea9c0, 32'h42bcc565};
test_output[26008:26015] = '{32'h42114ee5, 32'h42aef416, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bcc565};
test_input[26016:26023] = '{32'hc244802e, 32'h41be3d06, 32'hc222a1a1, 32'hc27a1efc, 32'hc1301990, 32'hc2aa4730, 32'hc2c658c9, 32'h41abc43b};
test_output[26016:26023] = '{32'h0, 32'h41be3d06, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41abc43b};
test_input[26024:26031] = '{32'h42a7f9b2, 32'h4191a100, 32'hc29ca38e, 32'hc1bfcc40, 32'hc1f8490d, 32'hc2854daa, 32'hc2163ec6, 32'h42a99d40};
test_output[26024:26031] = '{32'h42a7f9b2, 32'h4191a100, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a99d40};
test_input[26032:26039] = '{32'hc27d9866, 32'hc26d7ed8, 32'h4265305e, 32'hc29862f2, 32'h42c505eb, 32'h41dd5081, 32'h41d58e03, 32'h42b69b05};
test_output[26032:26039] = '{32'h0, 32'h0, 32'h4265305e, 32'h0, 32'h42c505eb, 32'h41dd5081, 32'h41d58e03, 32'h42b69b05};
test_input[26040:26047] = '{32'hc2aacb78, 32'h41f30021, 32'hc20de5c8, 32'h42220975, 32'hc206bead, 32'hc0ca4f5a, 32'hc2b000d5, 32'h423c4bd0};
test_output[26040:26047] = '{32'h0, 32'h41f30021, 32'h0, 32'h42220975, 32'h0, 32'h0, 32'h0, 32'h423c4bd0};
test_input[26048:26055] = '{32'hc115edc7, 32'h42b662d6, 32'h42bcc3d6, 32'h429c4127, 32'h422a107d, 32'h42834f6e, 32'h42308e98, 32'hc294bc9f};
test_output[26048:26055] = '{32'h0, 32'h42b662d6, 32'h42bcc3d6, 32'h429c4127, 32'h422a107d, 32'h42834f6e, 32'h42308e98, 32'h0};
test_input[26056:26063] = '{32'h415ced49, 32'h40c8bae6, 32'hc293fef7, 32'hc28c8d93, 32'hc2ac4e52, 32'hc28a6493, 32'h426c442b, 32'h3e13a123};
test_output[26056:26063] = '{32'h415ced49, 32'h40c8bae6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426c442b, 32'h3e13a123};
test_input[26064:26071] = '{32'hc2a7f93e, 32'hc29fec1f, 32'h42a0173a, 32'hc2865090, 32'hc201a768, 32'hc2bff437, 32'hc1252a22, 32'h4287aad0};
test_output[26064:26071] = '{32'h0, 32'h0, 32'h42a0173a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4287aad0};
test_input[26072:26079] = '{32'hbe1f0a22, 32'hc02d95d3, 32'hc2b6540e, 32'h42be9cf7, 32'h42c0fe77, 32'hc2606b59, 32'h4279a210, 32'h419af3cd};
test_output[26072:26079] = '{32'h0, 32'h0, 32'h0, 32'h42be9cf7, 32'h42c0fe77, 32'h0, 32'h4279a210, 32'h419af3cd};
test_input[26080:26087] = '{32'hc2983185, 32'hc2271559, 32'hc2248da5, 32'h42c7b523, 32'hc2014cd1, 32'hc0db20ac, 32'h429f4864, 32'hc2b5b8ad};
test_output[26080:26087] = '{32'h0, 32'h0, 32'h0, 32'h42c7b523, 32'h0, 32'h0, 32'h429f4864, 32'h0};
test_input[26088:26095] = '{32'h4169400c, 32'h41f17e25, 32'h4278a467, 32'h428df644, 32'h420e94c1, 32'hc097ddad, 32'hc28404b6, 32'hc2045666};
test_output[26088:26095] = '{32'h4169400c, 32'h41f17e25, 32'h4278a467, 32'h428df644, 32'h420e94c1, 32'h0, 32'h0, 32'h0};
test_input[26096:26103] = '{32'hc2a54f7f, 32'h41dfc6ac, 32'hbdcd0447, 32'h406e19a8, 32'hc233ccff, 32'hc2900189, 32'h4248d260, 32'h4093c846};
test_output[26096:26103] = '{32'h0, 32'h41dfc6ac, 32'h0, 32'h406e19a8, 32'h0, 32'h0, 32'h4248d260, 32'h4093c846};
test_input[26104:26111] = '{32'hc207be8b, 32'h4186bcd1, 32'hc2973967, 32'h42c770b3, 32'h41b473c4, 32'hc099ed33, 32'h3fd783ed, 32'h42a96251};
test_output[26104:26111] = '{32'h0, 32'h4186bcd1, 32'h0, 32'h42c770b3, 32'h41b473c4, 32'h0, 32'h3fd783ed, 32'h42a96251};
test_input[26112:26119] = '{32'h422b7ee5, 32'hc2bb22ad, 32'h42c636c5, 32'h4194fdea, 32'h42019c24, 32'hc1b45c82, 32'h40acdf1d, 32'hc2c190c6};
test_output[26112:26119] = '{32'h422b7ee5, 32'h0, 32'h42c636c5, 32'h4194fdea, 32'h42019c24, 32'h0, 32'h40acdf1d, 32'h0};
test_input[26120:26127] = '{32'h4210756d, 32'hc1f10d40, 32'hc1aea731, 32'h427c81a6, 32'h42aaf352, 32'h4237cb19, 32'hc1aeeef9, 32'h42989641};
test_output[26120:26127] = '{32'h4210756d, 32'h0, 32'h0, 32'h427c81a6, 32'h42aaf352, 32'h4237cb19, 32'h0, 32'h42989641};
test_input[26128:26135] = '{32'h41cb2a27, 32'h4220942b, 32'h428562c0, 32'hc1a0babe, 32'hc264a6d2, 32'hc1cfea19, 32'h421dd857, 32'hc2951a5e};
test_output[26128:26135] = '{32'h41cb2a27, 32'h4220942b, 32'h428562c0, 32'h0, 32'h0, 32'h0, 32'h421dd857, 32'h0};
test_input[26136:26143] = '{32'hc277a2a2, 32'hc1e3cea1, 32'h414c0b98, 32'hc11fba06, 32'h41c6f200, 32'hc139e426, 32'hc1e471b9, 32'hc138533b};
test_output[26136:26143] = '{32'h0, 32'h0, 32'h414c0b98, 32'h0, 32'h41c6f200, 32'h0, 32'h0, 32'h0};
test_input[26144:26151] = '{32'h428a6bab, 32'h42187faa, 32'h42580337, 32'h428c6598, 32'hc0d32bf5, 32'hc28395f5, 32'hc2bc482e, 32'h4260884e};
test_output[26144:26151] = '{32'h428a6bab, 32'h42187faa, 32'h42580337, 32'h428c6598, 32'h0, 32'h0, 32'h0, 32'h4260884e};
test_input[26152:26159] = '{32'h424935ca, 32'h42be00bf, 32'h428ccc96, 32'hc0411a1d, 32'hc1fca4b9, 32'hc20c7ba8, 32'hbfcc08a0, 32'hc1dc1528};
test_output[26152:26159] = '{32'h424935ca, 32'h42be00bf, 32'h428ccc96, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26160:26167] = '{32'h41fddbc0, 32'hc225a599, 32'h42052808, 32'hc257a7ca, 32'hc269bfda, 32'hc2ba8a58, 32'hc22377e6, 32'h41b6b4f3};
test_output[26160:26167] = '{32'h41fddbc0, 32'h0, 32'h42052808, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b6b4f3};
test_input[26168:26175] = '{32'hc2434615, 32'h429487bd, 32'hc2a5320c, 32'hc1c3420c, 32'hc228b240, 32'hc28ec5eb, 32'hc2657094, 32'hc1cc17d8};
test_output[26168:26175] = '{32'h0, 32'h429487bd, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26176:26183] = '{32'h42322830, 32'hc17576b6, 32'hc14d150d, 32'hc2b5975b, 32'hc2767d1e, 32'h4176f67b, 32'h42bb9a8b, 32'h42705b6b};
test_output[26176:26183] = '{32'h42322830, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4176f67b, 32'h42bb9a8b, 32'h42705b6b};
test_input[26184:26191] = '{32'hc1fd8d4d, 32'hc1ceb0be, 32'h4276c49f, 32'h42293937, 32'hc226f434, 32'hc2a5fadb, 32'hc202fbdf, 32'hc28a959a};
test_output[26184:26191] = '{32'h0, 32'h0, 32'h4276c49f, 32'h42293937, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26192:26199] = '{32'h42c413d5, 32'h4216f042, 32'hc22083d9, 32'hc1c074db, 32'hc25a14e6, 32'hc2adc81f, 32'hbf60628d, 32'h42b1633e};
test_output[26192:26199] = '{32'h42c413d5, 32'h4216f042, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b1633e};
test_input[26200:26207] = '{32'hc2762f50, 32'h41ad5064, 32'h42acc1e2, 32'h429b1070, 32'hc2b925da, 32'hc250c832, 32'h42c63845, 32'h42abcd0e};
test_output[26200:26207] = '{32'h0, 32'h41ad5064, 32'h42acc1e2, 32'h429b1070, 32'h0, 32'h0, 32'h42c63845, 32'h42abcd0e};
test_input[26208:26215] = '{32'hc2751426, 32'hc1a90408, 32'hc29b5541, 32'h4271d1a0, 32'hc2c70708, 32'h4050e527, 32'h42189f78, 32'hbf72f794};
test_output[26208:26215] = '{32'h0, 32'h0, 32'h0, 32'h4271d1a0, 32'h0, 32'h4050e527, 32'h42189f78, 32'h0};
test_input[26216:26223] = '{32'hc2aa3f11, 32'hc1227502, 32'hc20287df, 32'h428c09b6, 32'hc0599a54, 32'hc1fb7f93, 32'hc29a4eca, 32'h418dc612};
test_output[26216:26223] = '{32'h0, 32'h0, 32'h0, 32'h428c09b6, 32'h0, 32'h0, 32'h0, 32'h418dc612};
test_input[26224:26231] = '{32'h42b82654, 32'hbf35e1db, 32'h4297625c, 32'h42460e30, 32'hc26fe2d3, 32'h42192204, 32'h42a8f1af, 32'hc13067d2};
test_output[26224:26231] = '{32'h42b82654, 32'h0, 32'h4297625c, 32'h42460e30, 32'h0, 32'h42192204, 32'h42a8f1af, 32'h0};
test_input[26232:26239] = '{32'h42a05f79, 32'hc29f3e80, 32'hc2a89003, 32'hc2a3c457, 32'h40e30866, 32'h41d97aa2, 32'hc1550809, 32'h42562a06};
test_output[26232:26239] = '{32'h42a05f79, 32'h0, 32'h0, 32'h0, 32'h40e30866, 32'h41d97aa2, 32'h0, 32'h42562a06};
test_input[26240:26247] = '{32'h4295e863, 32'hc25fd175, 32'h42646b58, 32'hc2ab67e2, 32'h42955b14, 32'h425f1969, 32'h427f45ae, 32'hc28d856e};
test_output[26240:26247] = '{32'h4295e863, 32'h0, 32'h42646b58, 32'h0, 32'h42955b14, 32'h425f1969, 32'h427f45ae, 32'h0};
test_input[26248:26255] = '{32'hc1a32051, 32'h426d5421, 32'h427211df, 32'hc2ab643a, 32'h42017d13, 32'h429d4d95, 32'h41c8f09b, 32'h42b63298};
test_output[26248:26255] = '{32'h0, 32'h426d5421, 32'h427211df, 32'h0, 32'h42017d13, 32'h429d4d95, 32'h41c8f09b, 32'h42b63298};
test_input[26256:26263] = '{32'h417b0ac8, 32'hc25412f6, 32'h4254c29f, 32'h417c5d8c, 32'h428b69e4, 32'h42725045, 32'h42501b46, 32'h415eabd9};
test_output[26256:26263] = '{32'h417b0ac8, 32'h0, 32'h4254c29f, 32'h417c5d8c, 32'h428b69e4, 32'h42725045, 32'h42501b46, 32'h415eabd9};
test_input[26264:26271] = '{32'h420cd53c, 32'h424a0270, 32'h42c736ad, 32'hc236197b, 32'h42a78c0f, 32'h41b0f10a, 32'hc28cba8e, 32'hc21ce905};
test_output[26264:26271] = '{32'h420cd53c, 32'h424a0270, 32'h42c736ad, 32'h0, 32'h42a78c0f, 32'h41b0f10a, 32'h0, 32'h0};
test_input[26272:26279] = '{32'hc210d22d, 32'h42a9c601, 32'h425c0496, 32'hc2366f78, 32'hc1bf5b44, 32'hc2be6bd1, 32'hc1ccab92, 32'h42aef353};
test_output[26272:26279] = '{32'h0, 32'h42a9c601, 32'h425c0496, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42aef353};
test_input[26280:26287] = '{32'hc26adc92, 32'h4022e8a1, 32'hc2c3fdb6, 32'hc296df26, 32'h429254bf, 32'hc298f730, 32'hc2a92ea9, 32'hc2a23508};
test_output[26280:26287] = '{32'h0, 32'h4022e8a1, 32'h0, 32'h0, 32'h429254bf, 32'h0, 32'h0, 32'h0};
test_input[26288:26295] = '{32'h42ada51d, 32'h4246b9b1, 32'h42ae7ca5, 32'hc21a184c, 32'h42a1ef25, 32'h41bc3442, 32'h42803afd, 32'h42a26778};
test_output[26288:26295] = '{32'h42ada51d, 32'h4246b9b1, 32'h42ae7ca5, 32'h0, 32'h42a1ef25, 32'h41bc3442, 32'h42803afd, 32'h42a26778};
test_input[26296:26303] = '{32'h42128013, 32'hc2b4e5a5, 32'hc1c4098e, 32'hc221e52c, 32'hc290c2c8, 32'h40c94051, 32'hc1a9bc2a, 32'h424a4ae4};
test_output[26296:26303] = '{32'h42128013, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40c94051, 32'h0, 32'h424a4ae4};
test_input[26304:26311] = '{32'hc2501409, 32'h4239b992, 32'h42508f34, 32'hc21c6fdd, 32'h42c3f58c, 32'h4202af71, 32'h41865e84, 32'hc28c4794};
test_output[26304:26311] = '{32'h0, 32'h4239b992, 32'h42508f34, 32'h0, 32'h42c3f58c, 32'h4202af71, 32'h41865e84, 32'h0};
test_input[26312:26319] = '{32'h420e7d4b, 32'hc2538321, 32'h429486c3, 32'h41c67cf1, 32'h416de3e2, 32'h429e55ec, 32'hc26805e5, 32'hc21830be};
test_output[26312:26319] = '{32'h420e7d4b, 32'h0, 32'h429486c3, 32'h41c67cf1, 32'h416de3e2, 32'h429e55ec, 32'h0, 32'h0};
test_input[26320:26327] = '{32'hc226fef0, 32'h42a68a3d, 32'h42c5174a, 32'h3fe7dcb7, 32'hc2554018, 32'h42ac774a, 32'h426b705b, 32'hc223d773};
test_output[26320:26327] = '{32'h0, 32'h42a68a3d, 32'h42c5174a, 32'h3fe7dcb7, 32'h0, 32'h42ac774a, 32'h426b705b, 32'h0};
test_input[26328:26335] = '{32'hc28adc97, 32'h428106c5, 32'h420ca2a7, 32'h41471375, 32'hc08ffb72, 32'h42524817, 32'hc2c34ecd, 32'hc236f5fd};
test_output[26328:26335] = '{32'h0, 32'h428106c5, 32'h420ca2a7, 32'h41471375, 32'h0, 32'h42524817, 32'h0, 32'h0};
test_input[26336:26343] = '{32'h417c79c1, 32'h421901c3, 32'hc20b730a, 32'h428e5df6, 32'h4257900d, 32'hc1c18fcf, 32'hc1ed099c, 32'h429b4c61};
test_output[26336:26343] = '{32'h417c79c1, 32'h421901c3, 32'h0, 32'h428e5df6, 32'h4257900d, 32'h0, 32'h0, 32'h429b4c61};
test_input[26344:26351] = '{32'h424a93e4, 32'h4086e3d5, 32'h424a0489, 32'h4063fe22, 32'h42392203, 32'hc24c5b3e, 32'h41e10f5e, 32'hc1734eee};
test_output[26344:26351] = '{32'h424a93e4, 32'h4086e3d5, 32'h424a0489, 32'h4063fe22, 32'h42392203, 32'h0, 32'h41e10f5e, 32'h0};
test_input[26352:26359] = '{32'h40687e34, 32'hc2a2e05d, 32'h425ffb09, 32'h42122522, 32'hc2c73e2b, 32'h41b8c1fe, 32'hc2bde088, 32'h4197d136};
test_output[26352:26359] = '{32'h40687e34, 32'h0, 32'h425ffb09, 32'h42122522, 32'h0, 32'h41b8c1fe, 32'h0, 32'h4197d136};
test_input[26360:26367] = '{32'h429c6ae6, 32'hc1f95a26, 32'hc2820e1d, 32'hc2678a59, 32'hc186e224, 32'hc29bd779, 32'h42754e91, 32'h40415497};
test_output[26360:26367] = '{32'h429c6ae6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42754e91, 32'h40415497};
test_input[26368:26375] = '{32'h429a06ca, 32'hc1bc92df, 32'hc2838893, 32'hc182c40d, 32'h4296d018, 32'h42566af3, 32'hc24caca5, 32'hc1b01765};
test_output[26368:26375] = '{32'h429a06ca, 32'h0, 32'h0, 32'h0, 32'h4296d018, 32'h42566af3, 32'h0, 32'h0};
test_input[26376:26383] = '{32'hc0862f48, 32'hc2808e12, 32'hc2b467e6, 32'hc0f821ec, 32'h414f3666, 32'hc20fb617, 32'h4217576b, 32'h4225c4af};
test_output[26376:26383] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h414f3666, 32'h0, 32'h4217576b, 32'h4225c4af};
test_input[26384:26391] = '{32'hc2167ae8, 32'hc1e3c8d1, 32'hc1da23c9, 32'hc0383d63, 32'h401bd10e, 32'h42a14928, 32'h42ba995e, 32'hc2272498};
test_output[26384:26391] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h401bd10e, 32'h42a14928, 32'h42ba995e, 32'h0};
test_input[26392:26399] = '{32'h413bf78f, 32'h422b0cff, 32'h4267caa1, 32'h3fcc15e8, 32'h42a7820d, 32'hc2a20ee0, 32'h42866fbe, 32'hc2076144};
test_output[26392:26399] = '{32'h413bf78f, 32'h422b0cff, 32'h4267caa1, 32'h3fcc15e8, 32'h42a7820d, 32'h0, 32'h42866fbe, 32'h0};
test_input[26400:26407] = '{32'h42304de0, 32'h429e31b6, 32'h4290e4aa, 32'hc295ccda, 32'hc251d286, 32'hc196dec9, 32'hc1df87af, 32'hc239bb78};
test_output[26400:26407] = '{32'h42304de0, 32'h429e31b6, 32'h4290e4aa, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26408:26415] = '{32'hc10586b8, 32'hc1ac703d, 32'hc295acc9, 32'hc28b1938, 32'hc2656272, 32'h42698fd6, 32'h418a50d6, 32'hc197bbe1};
test_output[26408:26415] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42698fd6, 32'h418a50d6, 32'h0};
test_input[26416:26423] = '{32'h42849617, 32'h42290daa, 32'hc22c41fd, 32'hc18f2f85, 32'hc224513f, 32'h42c3c728, 32'hc245bc88, 32'h40359dd7};
test_output[26416:26423] = '{32'h42849617, 32'h42290daa, 32'h0, 32'h0, 32'h0, 32'h42c3c728, 32'h0, 32'h40359dd7};
test_input[26424:26431] = '{32'hc21b6582, 32'hc1fdbbe0, 32'h41b8c2b1, 32'h42c5d75f, 32'h41d00a18, 32'h42b2f34f, 32'hc299bef3, 32'h42b4a955};
test_output[26424:26431] = '{32'h0, 32'h0, 32'h41b8c2b1, 32'h42c5d75f, 32'h41d00a18, 32'h42b2f34f, 32'h0, 32'h42b4a955};
test_input[26432:26439] = '{32'hc08e7b82, 32'h4239d667, 32'hc2c4cea0, 32'h42c088db, 32'h4262a834, 32'hc20e37eb, 32'h423d10c7, 32'hc20c97a6};
test_output[26432:26439] = '{32'h0, 32'h4239d667, 32'h0, 32'h42c088db, 32'h4262a834, 32'h0, 32'h423d10c7, 32'h0};
test_input[26440:26447] = '{32'hc1870ce2, 32'hc235d0d2, 32'hc24504c9, 32'hc1f92745, 32'hc1ac70d9, 32'h41fa1e70, 32'h42bc8fb2, 32'hc0a525a9};
test_output[26440:26447] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41fa1e70, 32'h42bc8fb2, 32'h0};
test_input[26448:26455] = '{32'hc199ee99, 32'hc25afcb3, 32'h422033fc, 32'hc24f1ba1, 32'h42911b6f, 32'hc1cea978, 32'hc14ff806, 32'h42bd8b7d};
test_output[26448:26455] = '{32'h0, 32'h0, 32'h422033fc, 32'h0, 32'h42911b6f, 32'h0, 32'h0, 32'h42bd8b7d};
test_input[26456:26463] = '{32'h429b97ae, 32'hc1e4d30b, 32'hc2a4ebce, 32'hc2009ebb, 32'hc2913f8c, 32'hc2a8b368, 32'h40775b45, 32'h4236bd3a};
test_output[26456:26463] = '{32'h429b97ae, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40775b45, 32'h4236bd3a};
test_input[26464:26471] = '{32'hc25c2ed6, 32'h42927490, 32'h4119f6d9, 32'h428430bd, 32'h429fcba1, 32'hc26ffda5, 32'h42156d1f, 32'hc2829b9f};
test_output[26464:26471] = '{32'h0, 32'h42927490, 32'h4119f6d9, 32'h428430bd, 32'h429fcba1, 32'h0, 32'h42156d1f, 32'h0};
test_input[26472:26479] = '{32'h42c09d0b, 32'hc1f85a12, 32'h426a7da3, 32'hc25de7c1, 32'h428855a4, 32'hc2c03895, 32'h42abc276, 32'h42aecfd3};
test_output[26472:26479] = '{32'h42c09d0b, 32'h0, 32'h426a7da3, 32'h0, 32'h428855a4, 32'h0, 32'h42abc276, 32'h42aecfd3};
test_input[26480:26487] = '{32'hc1d8eee4, 32'hc2928064, 32'h4226740b, 32'hc29e5d36, 32'h42b2e008, 32'h41bf9cc2, 32'hc10e0b8d, 32'hc19918aa};
test_output[26480:26487] = '{32'h0, 32'h0, 32'h4226740b, 32'h0, 32'h42b2e008, 32'h41bf9cc2, 32'h0, 32'h0};
test_input[26488:26495] = '{32'hc226dbed, 32'hc2957284, 32'hc29b7020, 32'hc29628f8, 32'hc259d042, 32'h42c13262, 32'hc201e19d, 32'h4127fbac};
test_output[26488:26495] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c13262, 32'h0, 32'h4127fbac};
test_input[26496:26503] = '{32'h41b56da2, 32'hc280c757, 32'hc1f24139, 32'h42b4043f, 32'h426a0022, 32'hbf8a9ccb, 32'hc23fe6d1, 32'h4280a8c0};
test_output[26496:26503] = '{32'h41b56da2, 32'h0, 32'h0, 32'h42b4043f, 32'h426a0022, 32'h0, 32'h0, 32'h4280a8c0};
test_input[26504:26511] = '{32'h4294d15e, 32'h42acf3e3, 32'h4207b85b, 32'hc295a4ac, 32'h42109ad6, 32'h42b6ca91, 32'hc2a05e61, 32'h42475efc};
test_output[26504:26511] = '{32'h4294d15e, 32'h42acf3e3, 32'h4207b85b, 32'h0, 32'h42109ad6, 32'h42b6ca91, 32'h0, 32'h42475efc};
test_input[26512:26519] = '{32'hc2c140a1, 32'hc2c753e1, 32'h424ba353, 32'hc28a824e, 32'hc178d098, 32'h41303351, 32'hc26c003b, 32'hc2b6a4af};
test_output[26512:26519] = '{32'h0, 32'h0, 32'h424ba353, 32'h0, 32'h0, 32'h41303351, 32'h0, 32'h0};
test_input[26520:26527] = '{32'hc1f2b4a2, 32'h4283e9df, 32'hc291cdaa, 32'h40b6299a, 32'hc0996780, 32'h42727351, 32'hc20219b9, 32'h42c21b98};
test_output[26520:26527] = '{32'h0, 32'h4283e9df, 32'h0, 32'h40b6299a, 32'h0, 32'h42727351, 32'h0, 32'h42c21b98};
test_input[26528:26535] = '{32'h428ea6b9, 32'hc219e2b5, 32'hc2a6686e, 32'h4256a6f2, 32'h421a97b2, 32'hc23276da, 32'hc28e81ea, 32'hc28cf752};
test_output[26528:26535] = '{32'h428ea6b9, 32'h0, 32'h0, 32'h4256a6f2, 32'h421a97b2, 32'h0, 32'h0, 32'h0};
test_input[26536:26543] = '{32'h427466ed, 32'h412abe38, 32'hc17977b9, 32'hc200b923, 32'h4079b8a0, 32'h42be50d2, 32'h425e5d0a, 32'h429ebf07};
test_output[26536:26543] = '{32'h427466ed, 32'h412abe38, 32'h0, 32'h0, 32'h4079b8a0, 32'h42be50d2, 32'h425e5d0a, 32'h429ebf07};
test_input[26544:26551] = '{32'h42654194, 32'hc20056d7, 32'hc14390e9, 32'hc295ae9e, 32'hc20cb95f, 32'hc25ce32a, 32'h42687dfc, 32'h41798a48};
test_output[26544:26551] = '{32'h42654194, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42687dfc, 32'h41798a48};
test_input[26552:26559] = '{32'h429c9e91, 32'hc1ed4ff1, 32'hc2c371df, 32'hc2c4f5e7, 32'hc2bc3727, 32'h429aa60f, 32'h4250dfb5, 32'hc2bd427f};
test_output[26552:26559] = '{32'h429c9e91, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429aa60f, 32'h4250dfb5, 32'h0};
test_input[26560:26567] = '{32'hc1f7b6da, 32'hc1e7fa92, 32'hc299c157, 32'hc2a19fce, 32'h4273cce6, 32'hc0c04452, 32'h42265a55, 32'h423d244d};
test_output[26560:26567] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4273cce6, 32'h0, 32'h42265a55, 32'h423d244d};
test_input[26568:26575] = '{32'hc207d73c, 32'hc21690ab, 32'h429e1816, 32'hc2bdc911, 32'h428d8ab5, 32'hc2bb8be9, 32'h41b148f0, 32'hc27bf63a};
test_output[26568:26575] = '{32'h0, 32'h0, 32'h429e1816, 32'h0, 32'h428d8ab5, 32'h0, 32'h41b148f0, 32'h0};
test_input[26576:26583] = '{32'h424d3a4f, 32'hc1acd2e8, 32'h410389a4, 32'h42a28e30, 32'hc2a56ef7, 32'hc235b7df, 32'hc18fc364, 32'hc298a5a6};
test_output[26576:26583] = '{32'h424d3a4f, 32'h0, 32'h410389a4, 32'h42a28e30, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26584:26591] = '{32'h4294a1fd, 32'hc2aa1f6a, 32'h421310e7, 32'h42a9cb52, 32'h4230253c, 32'h427cb626, 32'hc2bc5814, 32'h42879bc5};
test_output[26584:26591] = '{32'h4294a1fd, 32'h0, 32'h421310e7, 32'h42a9cb52, 32'h4230253c, 32'h427cb626, 32'h0, 32'h42879bc5};
test_input[26592:26599] = '{32'h42acae53, 32'h4280fa56, 32'h3f14f101, 32'hc276db4a, 32'h4214d12e, 32'hc2bccd21, 32'hc2b022f9, 32'h41230de1};
test_output[26592:26599] = '{32'h42acae53, 32'h4280fa56, 32'h3f14f101, 32'h0, 32'h4214d12e, 32'h0, 32'h0, 32'h41230de1};
test_input[26600:26607] = '{32'hc21daf53, 32'hc13e7e78, 32'hc289baf4, 32'h4291d1a6, 32'hc2333850, 32'h41999804, 32'hc2a9b129, 32'hc2ada03f};
test_output[26600:26607] = '{32'h0, 32'h0, 32'h0, 32'h4291d1a6, 32'h0, 32'h41999804, 32'h0, 32'h0};
test_input[26608:26615] = '{32'hc2c15f84, 32'hc27a7752, 32'hc28453dd, 32'hc21da3ff, 32'h427e5a30, 32'hc2849dc3, 32'hc2b23e25, 32'hc29ae90b};
test_output[26608:26615] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h427e5a30, 32'h0, 32'h0, 32'h0};
test_input[26616:26623] = '{32'hc25ffecb, 32'h40544955, 32'h4221d24f, 32'h4124f392, 32'h40eecaa0, 32'hc2c3fd99, 32'hc2193e40, 32'h4275a3c8};
test_output[26616:26623] = '{32'h0, 32'h40544955, 32'h4221d24f, 32'h4124f392, 32'h40eecaa0, 32'h0, 32'h0, 32'h4275a3c8};
test_input[26624:26631] = '{32'hc2b62d18, 32'h40a73072, 32'hc1deb327, 32'hc1a3a448, 32'hc032b5a3, 32'h42c2063c, 32'h429b996d, 32'h42200c0c};
test_output[26624:26631] = '{32'h0, 32'h40a73072, 32'h0, 32'h0, 32'h0, 32'h42c2063c, 32'h429b996d, 32'h42200c0c};
test_input[26632:26639] = '{32'hc23c953a, 32'h4254952e, 32'h4279fc24, 32'h428ab3d5, 32'hc2c4a248, 32'hc2ba4cb3, 32'hc2a758f8, 32'hc28747ab};
test_output[26632:26639] = '{32'h0, 32'h4254952e, 32'h4279fc24, 32'h428ab3d5, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26640:26647] = '{32'h41dbe0ee, 32'hc29b157c, 32'h4222402a, 32'hc2aa1292, 32'hc26ffc9e, 32'hc1c89d37, 32'hc1519cc9, 32'hc2afdbdf};
test_output[26640:26647] = '{32'h41dbe0ee, 32'h0, 32'h4222402a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26648:26655] = '{32'h428ca74a, 32'hc2462159, 32'hc1a4d9f9, 32'h41e7b6c3, 32'h41ca0116, 32'hc196e3e5, 32'hc085cdff, 32'hc2944f4d};
test_output[26648:26655] = '{32'h428ca74a, 32'h0, 32'h0, 32'h41e7b6c3, 32'h41ca0116, 32'h0, 32'h0, 32'h0};
test_input[26656:26663] = '{32'h42bd743c, 32'hc2c05255, 32'hc21cf5df, 32'h42432c56, 32'h420b261f, 32'h4057e732, 32'h42aeae67, 32'h4283ca5a};
test_output[26656:26663] = '{32'h42bd743c, 32'h0, 32'h0, 32'h42432c56, 32'h420b261f, 32'h4057e732, 32'h42aeae67, 32'h4283ca5a};
test_input[26664:26671] = '{32'hc220fa76, 32'hc0403e40, 32'hc2532646, 32'hc2911fae, 32'h420451b7, 32'h42978632, 32'h426bde2e, 32'hc25ca830};
test_output[26664:26671] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h420451b7, 32'h42978632, 32'h426bde2e, 32'h0};
test_input[26672:26679] = '{32'hc2c50454, 32'h427a13f2, 32'h421f7bc0, 32'h42c1760e, 32'hc2846b41, 32'h42b01f14, 32'h423f7c01, 32'hc117378c};
test_output[26672:26679] = '{32'h0, 32'h427a13f2, 32'h421f7bc0, 32'h42c1760e, 32'h0, 32'h42b01f14, 32'h423f7c01, 32'h0};
test_input[26680:26687] = '{32'hc25842dc, 32'h428916da, 32'h4147e5f7, 32'hc2c577f5, 32'h418e86b3, 32'hc29fc092, 32'hc146ced7, 32'hc09a74d0};
test_output[26680:26687] = '{32'h0, 32'h428916da, 32'h4147e5f7, 32'h0, 32'h418e86b3, 32'h0, 32'h0, 32'h0};
test_input[26688:26695] = '{32'h41a25ec0, 32'hc2114be1, 32'h4219c5b0, 32'h40e257f2, 32'hc279082b, 32'hc00f3f43, 32'h42a50b70, 32'hc0cc88a3};
test_output[26688:26695] = '{32'h41a25ec0, 32'h0, 32'h4219c5b0, 32'h40e257f2, 32'h0, 32'h0, 32'h42a50b70, 32'h0};
test_input[26696:26703] = '{32'hc28895a7, 32'hc1b83a1d, 32'hc24df2dd, 32'hc1518ef0, 32'h42c56f6f, 32'hc2468df9, 32'h40afb062, 32'hc2c2ad6f};
test_output[26696:26703] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42c56f6f, 32'h0, 32'h40afb062, 32'h0};
test_input[26704:26711] = '{32'hc15ebad8, 32'hc1eee6b3, 32'hc18d036e, 32'h4098b4e0, 32'hc235de1f, 32'h41291a0e, 32'hc239ff7c, 32'hc0f16f9b};
test_output[26704:26711] = '{32'h0, 32'h0, 32'h0, 32'h4098b4e0, 32'h0, 32'h41291a0e, 32'h0, 32'h0};
test_input[26712:26719] = '{32'hc1e14b95, 32'h426a57fc, 32'hc131dbed, 32'hc299760b, 32'hc0691b32, 32'hc1b8d4c5, 32'hc2328c06, 32'hc2b9121c};
test_output[26712:26719] = '{32'h0, 32'h426a57fc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26720:26727] = '{32'hc2ba0376, 32'hc2907b70, 32'hc2b44628, 32'h40b77845, 32'hbf4233cc, 32'h42c3ac49, 32'hc24973de, 32'hc2832b2d};
test_output[26720:26727] = '{32'h0, 32'h0, 32'h0, 32'h40b77845, 32'h0, 32'h42c3ac49, 32'h0, 32'h0};
test_input[26728:26735] = '{32'h428860c4, 32'hc2571766, 32'hc1f56f66, 32'h3f99572d, 32'hc2aac4a1, 32'h421da20b, 32'hc21869df, 32'hc0acb939};
test_output[26728:26735] = '{32'h428860c4, 32'h0, 32'h0, 32'h3f99572d, 32'h0, 32'h421da20b, 32'h0, 32'h0};
test_input[26736:26743] = '{32'hc246f7e3, 32'h4291ba66, 32'hc241c3ff, 32'hc242d97e, 32'h421bd1d9, 32'h42438acd, 32'h4246a16d, 32'hc0c748df};
test_output[26736:26743] = '{32'h0, 32'h4291ba66, 32'h0, 32'h0, 32'h421bd1d9, 32'h42438acd, 32'h4246a16d, 32'h0};
test_input[26744:26751] = '{32'h42aebb7e, 32'hc1aa3847, 32'hc04f32f7, 32'h419f29e4, 32'h418df78a, 32'hc2743172, 32'h42283df8, 32'h40dae350};
test_output[26744:26751] = '{32'h42aebb7e, 32'h0, 32'h0, 32'h419f29e4, 32'h418df78a, 32'h0, 32'h42283df8, 32'h40dae350};
test_input[26752:26759] = '{32'h429f5814, 32'hc1054614, 32'h4269b731, 32'h42784ec1, 32'hc2b1878c, 32'hc1c8106f, 32'h423eda8b, 32'h40ea175b};
test_output[26752:26759] = '{32'h429f5814, 32'h0, 32'h4269b731, 32'h42784ec1, 32'h0, 32'h0, 32'h423eda8b, 32'h40ea175b};
test_input[26760:26767] = '{32'hc2c2d43a, 32'h420db02f, 32'h42c28ac9, 32'h41fc1cce, 32'h428835c8, 32'h4237a214, 32'h42ba9f13, 32'hc2a51f76};
test_output[26760:26767] = '{32'h0, 32'h420db02f, 32'h42c28ac9, 32'h41fc1cce, 32'h428835c8, 32'h4237a214, 32'h42ba9f13, 32'h0};
test_input[26768:26775] = '{32'h420bd1af, 32'h4265e715, 32'h42a6776e, 32'hc20295c6, 32'hc14f4f21, 32'h422bb7b8, 32'hc1865a60, 32'hc1667c69};
test_output[26768:26775] = '{32'h420bd1af, 32'h4265e715, 32'h42a6776e, 32'h0, 32'h0, 32'h422bb7b8, 32'h0, 32'h0};
test_input[26776:26783] = '{32'hc2291d44, 32'h42789943, 32'h40c9c220, 32'h422dc4cf, 32'h401f69a5, 32'h41f9d94c, 32'hc1ea50b3, 32'hc2c03a05};
test_output[26776:26783] = '{32'h0, 32'h42789943, 32'h40c9c220, 32'h422dc4cf, 32'h401f69a5, 32'h41f9d94c, 32'h0, 32'h0};
test_input[26784:26791] = '{32'hc16ffd37, 32'hc205f0c5, 32'h418437ce, 32'hc280ac76, 32'hc26cc0e8, 32'hbed5e243, 32'h424e2e89, 32'hc29b095e};
test_output[26784:26791] = '{32'h0, 32'h0, 32'h418437ce, 32'h0, 32'h0, 32'h0, 32'h424e2e89, 32'h0};
test_input[26792:26799] = '{32'h42283074, 32'h42a48a7b, 32'h42a9b779, 32'hc2157b38, 32'h4272fb74, 32'h42423141, 32'h429b9032, 32'h4220124d};
test_output[26792:26799] = '{32'h42283074, 32'h42a48a7b, 32'h42a9b779, 32'h0, 32'h4272fb74, 32'h42423141, 32'h429b9032, 32'h4220124d};
test_input[26800:26807] = '{32'h42318d19, 32'hc1817eed, 32'h424cb495, 32'hc2457411, 32'h428ea2a6, 32'hc2ac0bc3, 32'h42195393, 32'h42bab06d};
test_output[26800:26807] = '{32'h42318d19, 32'h0, 32'h424cb495, 32'h0, 32'h428ea2a6, 32'h0, 32'h42195393, 32'h42bab06d};
test_input[26808:26815] = '{32'h40c07fae, 32'h42a9ae5d, 32'h42bc3929, 32'hc20af14d, 32'h41457a01, 32'h42c7818d, 32'hc2069d12, 32'h42b6351d};
test_output[26808:26815] = '{32'h40c07fae, 32'h42a9ae5d, 32'h42bc3929, 32'h0, 32'h41457a01, 32'h42c7818d, 32'h0, 32'h42b6351d};
test_input[26816:26823] = '{32'h42a15992, 32'hc24ed678, 32'hc29549d9, 32'hc0f346be, 32'h421f6eda, 32'hc22163c0, 32'h425e9a8d, 32'h41359c82};
test_output[26816:26823] = '{32'h42a15992, 32'h0, 32'h0, 32'h0, 32'h421f6eda, 32'h0, 32'h425e9a8d, 32'h41359c82};
test_input[26824:26831] = '{32'hc1c17709, 32'hc1d583cc, 32'hc27a825c, 32'hc25e76f5, 32'hbec2bd0d, 32'h4275b32f, 32'h423c70cc, 32'hc1800b9f};
test_output[26824:26831] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4275b32f, 32'h423c70cc, 32'h0};
test_input[26832:26839] = '{32'h424db7e1, 32'hc2972cee, 32'h41da228a, 32'h42500d65, 32'h42c144a4, 32'h429ca43c, 32'h41c5538e, 32'hc2bfc412};
test_output[26832:26839] = '{32'h424db7e1, 32'h0, 32'h41da228a, 32'h42500d65, 32'h42c144a4, 32'h429ca43c, 32'h41c5538e, 32'h0};
test_input[26840:26847] = '{32'h4294398d, 32'h422849c3, 32'hc2b28696, 32'hc20a63a7, 32'h40c87fcd, 32'h42873cb2, 32'hc26d503f, 32'hc2ae671b};
test_output[26840:26847] = '{32'h4294398d, 32'h422849c3, 32'h0, 32'h0, 32'h40c87fcd, 32'h42873cb2, 32'h0, 32'h0};
test_input[26848:26855] = '{32'hc1060ff1, 32'hc1b2eb39, 32'h40faf858, 32'h4170a3ee, 32'h427db148, 32'hc2bfa77f, 32'h416e113b, 32'h426d6f01};
test_output[26848:26855] = '{32'h0, 32'h0, 32'h40faf858, 32'h4170a3ee, 32'h427db148, 32'h0, 32'h416e113b, 32'h426d6f01};
test_input[26856:26863] = '{32'h4223f839, 32'hc245d293, 32'hc1628a22, 32'h4239da40, 32'h4236d3d8, 32'h42b9d84c, 32'h42782cf3, 32'hc2b233f3};
test_output[26856:26863] = '{32'h4223f839, 32'h0, 32'h0, 32'h4239da40, 32'h4236d3d8, 32'h42b9d84c, 32'h42782cf3, 32'h0};
test_input[26864:26871] = '{32'h4248e7fe, 32'hc2c08765, 32'h4197dab8, 32'hc2ad5fe2, 32'hc1f262e5, 32'h42c093e1, 32'hc1d6b67e, 32'hc168eae1};
test_output[26864:26871] = '{32'h4248e7fe, 32'h0, 32'h4197dab8, 32'h0, 32'h0, 32'h42c093e1, 32'h0, 32'h0};
test_input[26872:26879] = '{32'hc2b1af43, 32'h40900605, 32'h423cfc28, 32'hc0ec8e60, 32'h426e20eb, 32'h425f95e4, 32'h42a952e1, 32'hc2ada417};
test_output[26872:26879] = '{32'h0, 32'h40900605, 32'h423cfc28, 32'h0, 32'h426e20eb, 32'h425f95e4, 32'h42a952e1, 32'h0};
test_input[26880:26887] = '{32'h4270829f, 32'hc04db5f2, 32'h4187a0f9, 32'h42951bf6, 32'hc2c407cf, 32'h4199713c, 32'hc2ab4126, 32'h424ec427};
test_output[26880:26887] = '{32'h4270829f, 32'h0, 32'h4187a0f9, 32'h42951bf6, 32'h0, 32'h4199713c, 32'h0, 32'h424ec427};
test_input[26888:26895] = '{32'h41f22428, 32'h426ef051, 32'h4243e4a1, 32'hc2940f72, 32'hc29450b7, 32'h4189b220, 32'h421e8740, 32'h42c6fb30};
test_output[26888:26895] = '{32'h41f22428, 32'h426ef051, 32'h4243e4a1, 32'h0, 32'h0, 32'h4189b220, 32'h421e8740, 32'h42c6fb30};
test_input[26896:26903] = '{32'h427af7bf, 32'hc2c69d99, 32'h429a4519, 32'hc21da7a9, 32'h4210d12c, 32'h415e4a6a, 32'hc1c084df, 32'h42996995};
test_output[26896:26903] = '{32'h427af7bf, 32'h0, 32'h429a4519, 32'h0, 32'h4210d12c, 32'h415e4a6a, 32'h0, 32'h42996995};
test_input[26904:26911] = '{32'hc264fe88, 32'hc25f6f8b, 32'hc1cb7295, 32'h42149c39, 32'hc1964956, 32'h41e80df4, 32'hc28db03b, 32'hc0b71f16};
test_output[26904:26911] = '{32'h0, 32'h0, 32'h0, 32'h42149c39, 32'h0, 32'h41e80df4, 32'h0, 32'h0};
test_input[26912:26919] = '{32'hc1e74408, 32'hbf17dc6c, 32'hc2b23220, 32'hc1e34fe0, 32'hc2ba02ed, 32'hc20d2351, 32'hbfc0eb5d, 32'hc0139806};
test_output[26912:26919] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26920:26927] = '{32'h40216377, 32'hc291a9d3, 32'hc2890a24, 32'h421e82fc, 32'h427ffa85, 32'hc11ce745, 32'hc2bcd870, 32'h4256a7b7};
test_output[26920:26927] = '{32'h40216377, 32'h0, 32'h0, 32'h421e82fc, 32'h427ffa85, 32'h0, 32'h0, 32'h4256a7b7};
test_input[26928:26935] = '{32'h4209e3d4, 32'h40a5cede, 32'hc1deb7a2, 32'hc20a1fdf, 32'h41bf0401, 32'hc16f3c01, 32'h42242576, 32'hbf444808};
test_output[26928:26935] = '{32'h4209e3d4, 32'h40a5cede, 32'h0, 32'h0, 32'h41bf0401, 32'h0, 32'h42242576, 32'h0};
test_input[26936:26943] = '{32'h41985069, 32'hc283d285, 32'h421b06e5, 32'h42bf63a2, 32'h41c529c5, 32'h41e7d8a6, 32'h42ac5573, 32'h4205d644};
test_output[26936:26943] = '{32'h41985069, 32'h0, 32'h421b06e5, 32'h42bf63a2, 32'h41c529c5, 32'h41e7d8a6, 32'h42ac5573, 32'h4205d644};
test_input[26944:26951] = '{32'hc2305bde, 32'h41cb2974, 32'h426943af, 32'h42bfb2bc, 32'hc11fc849, 32'hc189c0d6, 32'hc241726f, 32'hc2120c20};
test_output[26944:26951] = '{32'h0, 32'h41cb2974, 32'h426943af, 32'h42bfb2bc, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26952:26959] = '{32'hc28806ec, 32'h42c7f641, 32'h42a9f6ee, 32'h4290c4fa, 32'h42c350eb, 32'hc20b60e7, 32'hc23cfc2d, 32'hc1cef239};
test_output[26952:26959] = '{32'h0, 32'h42c7f641, 32'h42a9f6ee, 32'h4290c4fa, 32'h42c350eb, 32'h0, 32'h0, 32'h0};
test_input[26960:26967] = '{32'h41901f98, 32'hc2ab1579, 32'h42c669a6, 32'hc295162a, 32'hc0da28b6, 32'h425b19bb, 32'h42a9f9c4, 32'hc1ec788f};
test_output[26960:26967] = '{32'h41901f98, 32'h0, 32'h42c669a6, 32'h0, 32'h0, 32'h425b19bb, 32'h42a9f9c4, 32'h0};
test_input[26968:26975] = '{32'hc29833b2, 32'hbfb5c790, 32'h417f9d0f, 32'hc0de9f85, 32'h414908df, 32'hc203025d, 32'h42468a92, 32'h401b03a0};
test_output[26968:26975] = '{32'h0, 32'h0, 32'h417f9d0f, 32'h0, 32'h414908df, 32'h0, 32'h42468a92, 32'h401b03a0};
test_input[26976:26983] = '{32'h422e06fd, 32'h4286593d, 32'hc1e9eac4, 32'h42b2474f, 32'h428cd935, 32'h4261c999, 32'h42287f42, 32'hc2979a70};
test_output[26976:26983] = '{32'h422e06fd, 32'h4286593d, 32'h0, 32'h42b2474f, 32'h428cd935, 32'h4261c999, 32'h42287f42, 32'h0};
test_input[26984:26991] = '{32'hc151c4e4, 32'h4208de91, 32'hc21305e0, 32'h422eff8e, 32'hc2c5a191, 32'hc296b20e, 32'h4227ad9a, 32'h42b2ade2};
test_output[26984:26991] = '{32'h0, 32'h4208de91, 32'h0, 32'h422eff8e, 32'h0, 32'h0, 32'h4227ad9a, 32'h42b2ade2};
test_input[26992:26999] = '{32'h4287f49c, 32'h42a727bd, 32'h41aee5dc, 32'h428a84e9, 32'hc21d09fc, 32'hc29f07cd, 32'h4243adcb, 32'h4277f4c4};
test_output[26992:26999] = '{32'h4287f49c, 32'h42a727bd, 32'h41aee5dc, 32'h428a84e9, 32'h0, 32'h0, 32'h4243adcb, 32'h4277f4c4};
test_input[27000:27007] = '{32'hc13969a0, 32'hc2ba51c1, 32'h4209dbb6, 32'hc1576d28, 32'hc276933d, 32'hc1861662, 32'h42b6b061, 32'h42428835};
test_output[27000:27007] = '{32'h0, 32'h0, 32'h4209dbb6, 32'h0, 32'h0, 32'h0, 32'h42b6b061, 32'h42428835};
test_input[27008:27015] = '{32'hc0fd9a4e, 32'h415bfb36, 32'h41c49b9b, 32'hc2adafbb, 32'hc0b1d31b, 32'hc2874c8c, 32'h4266a173, 32'h412b0ddf};
test_output[27008:27015] = '{32'h0, 32'h415bfb36, 32'h41c49b9b, 32'h0, 32'h0, 32'h0, 32'h4266a173, 32'h412b0ddf};
test_input[27016:27023] = '{32'hc14213e0, 32'h42c60e32, 32'h426f268e, 32'hc0d36038, 32'hc15f4d96, 32'h42ad8d4b, 32'h41a24c48, 32'h42a786fd};
test_output[27016:27023] = '{32'h0, 32'h42c60e32, 32'h426f268e, 32'h0, 32'h0, 32'h42ad8d4b, 32'h41a24c48, 32'h42a786fd};
test_input[27024:27031] = '{32'h4176e703, 32'h42afd91a, 32'hc2b640e8, 32'h41de6100, 32'h40a2bbf1, 32'hc253e5cc, 32'hc2a28006, 32'h42bfbf51};
test_output[27024:27031] = '{32'h4176e703, 32'h42afd91a, 32'h0, 32'h41de6100, 32'h40a2bbf1, 32'h0, 32'h0, 32'h42bfbf51};
test_input[27032:27039] = '{32'h3f9e4314, 32'hc2c4ced6, 32'h404f9922, 32'h41e92ca3, 32'hc2b0cd72, 32'hc1d893de, 32'hc2a11422, 32'h429ff45b};
test_output[27032:27039] = '{32'h3f9e4314, 32'h0, 32'h404f9922, 32'h41e92ca3, 32'h0, 32'h0, 32'h0, 32'h429ff45b};
test_input[27040:27047] = '{32'hc299281e, 32'h41b75971, 32'h427f1746, 32'h4230d13b, 32'hc26f612c, 32'hc2959cc6, 32'h42580745, 32'h42a2dda8};
test_output[27040:27047] = '{32'h0, 32'h41b75971, 32'h427f1746, 32'h4230d13b, 32'h0, 32'h0, 32'h42580745, 32'h42a2dda8};
test_input[27048:27055] = '{32'hc0acdc72, 32'h42793921, 32'h42af3e0b, 32'hc23f7e0b, 32'hc13dd2fe, 32'hc193baa0, 32'hc159a2ed, 32'hc2c34bd3};
test_output[27048:27055] = '{32'h0, 32'h42793921, 32'h42af3e0b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27056:27063] = '{32'h41eeac29, 32'hc2bd27e8, 32'h422505a2, 32'hc2c70b88, 32'h41b99ad8, 32'h415c1e54, 32'hc1071fbf, 32'h42aaf245};
test_output[27056:27063] = '{32'h41eeac29, 32'h0, 32'h422505a2, 32'h0, 32'h41b99ad8, 32'h415c1e54, 32'h0, 32'h42aaf245};
test_input[27064:27071] = '{32'h427da1e6, 32'h42a06810, 32'hc289220d, 32'hbfae6a34, 32'hc29239bd, 32'h41acb4c4, 32'hc19811a9, 32'h427e5b95};
test_output[27064:27071] = '{32'h427da1e6, 32'h42a06810, 32'h0, 32'h0, 32'h0, 32'h41acb4c4, 32'h0, 32'h427e5b95};
test_input[27072:27079] = '{32'hc29660e4, 32'hc210482b, 32'h42819af8, 32'h426912cb, 32'h42a86974, 32'hc173dfd4, 32'hbec6f5bd, 32'hc176c8d9};
test_output[27072:27079] = '{32'h0, 32'h0, 32'h42819af8, 32'h426912cb, 32'h42a86974, 32'h0, 32'h0, 32'h0};
test_input[27080:27087] = '{32'hc1733856, 32'hc27c63de, 32'hc22ffdf6, 32'h429af2f9, 32'hbf27fe01, 32'h41717877, 32'hc2a1b2eb, 32'h41f97550};
test_output[27080:27087] = '{32'h0, 32'h0, 32'h0, 32'h429af2f9, 32'h0, 32'h41717877, 32'h0, 32'h41f97550};
test_input[27088:27095] = '{32'hc2884abb, 32'h42b8f112, 32'hc2032af3, 32'hc2bb820d, 32'h4282d908, 32'hc2bc62a3, 32'h428da6c7, 32'h42b7b1c8};
test_output[27088:27095] = '{32'h0, 32'h42b8f112, 32'h0, 32'h0, 32'h4282d908, 32'h0, 32'h428da6c7, 32'h42b7b1c8};
test_input[27096:27103] = '{32'hc2a754dd, 32'hc28e008e, 32'h42496914, 32'h42608804, 32'hc1b90518, 32'h40faa5bb, 32'h429f1905, 32'h4207802f};
test_output[27096:27103] = '{32'h0, 32'h0, 32'h42496914, 32'h42608804, 32'h0, 32'h40faa5bb, 32'h429f1905, 32'h4207802f};
test_input[27104:27111] = '{32'h4229071f, 32'h42a541d8, 32'h429cf71d, 32'hc2073f17, 32'h42bd1685, 32'h427a7833, 32'hc2a8a78e, 32'h4100f18e};
test_output[27104:27111] = '{32'h4229071f, 32'h42a541d8, 32'h429cf71d, 32'h0, 32'h42bd1685, 32'h427a7833, 32'h0, 32'h4100f18e};
test_input[27112:27119] = '{32'hc289e34b, 32'hc02b0e40, 32'h422d8d68, 32'h42936082, 32'hc1ca14ec, 32'hc1c6099f, 32'h42891bf9, 32'h419afaf3};
test_output[27112:27119] = '{32'h0, 32'h0, 32'h422d8d68, 32'h42936082, 32'h0, 32'h0, 32'h42891bf9, 32'h419afaf3};
test_input[27120:27127] = '{32'hc1e6347c, 32'hc183138d, 32'h427682fa, 32'h41aaf2dc, 32'h40a79272, 32'h428b78bb, 32'h42c1fa32, 32'h427c1586};
test_output[27120:27127] = '{32'h0, 32'h0, 32'h427682fa, 32'h41aaf2dc, 32'h40a79272, 32'h428b78bb, 32'h42c1fa32, 32'h427c1586};
test_input[27128:27135] = '{32'h425839e4, 32'hc2aaceb2, 32'hc1d9e871, 32'hc25576b2, 32'h41cbfa05, 32'h42477808, 32'hc0ac4760, 32'h4287bbaf};
test_output[27128:27135] = '{32'h425839e4, 32'h0, 32'h0, 32'h0, 32'h41cbfa05, 32'h42477808, 32'h0, 32'h4287bbaf};
test_input[27136:27143] = '{32'h42873654, 32'h42288f6d, 32'hc27400ef, 32'hc2b0ea36, 32'h42a68ff0, 32'hc278ee68, 32'h41934d9e, 32'h3f2235f7};
test_output[27136:27143] = '{32'h42873654, 32'h42288f6d, 32'h0, 32'h0, 32'h42a68ff0, 32'h0, 32'h41934d9e, 32'h3f2235f7};
test_input[27144:27151] = '{32'hc1e33ef8, 32'hc2189ef9, 32'hc1fec728, 32'h41aae628, 32'h422306c3, 32'hc28f99c8, 32'h42af7701, 32'h42ad0299};
test_output[27144:27151] = '{32'h0, 32'h0, 32'h0, 32'h41aae628, 32'h422306c3, 32'h0, 32'h42af7701, 32'h42ad0299};
test_input[27152:27159] = '{32'h42469e38, 32'h42a7bb89, 32'h41ee0cd2, 32'hc1b1bbe7, 32'hc2bba984, 32'hc233cd7d, 32'h4226591e, 32'h4249b436};
test_output[27152:27159] = '{32'h42469e38, 32'h42a7bb89, 32'h41ee0cd2, 32'h0, 32'h0, 32'h0, 32'h4226591e, 32'h4249b436};
test_input[27160:27167] = '{32'h417a2e6f, 32'h42a0854f, 32'h42ada80d, 32'hc2b6a8ee, 32'hc23c8c1a, 32'h42ba4a68, 32'h4166d37e, 32'h4192d7d5};
test_output[27160:27167] = '{32'h417a2e6f, 32'h42a0854f, 32'h42ada80d, 32'h0, 32'h0, 32'h42ba4a68, 32'h4166d37e, 32'h4192d7d5};
test_input[27168:27175] = '{32'h41a4f3b7, 32'hc246b689, 32'hc29ec6ce, 32'hc2206af7, 32'h42862797, 32'hc2996ec4, 32'hc282c4d4, 32'h4150244d};
test_output[27168:27175] = '{32'h41a4f3b7, 32'h0, 32'h0, 32'h0, 32'h42862797, 32'h0, 32'h0, 32'h4150244d};
test_input[27176:27183] = '{32'hc2078737, 32'h41e8733a, 32'hc27d922b, 32'h4224f607, 32'h42072eb3, 32'hc24e3569, 32'hc2285262, 32'hc2a9bbc9};
test_output[27176:27183] = '{32'h0, 32'h41e8733a, 32'h0, 32'h4224f607, 32'h42072eb3, 32'h0, 32'h0, 32'h0};
test_input[27184:27191] = '{32'hc2aee7c2, 32'h4280bc48, 32'h422b0ec3, 32'h41595f8c, 32'h42528b0e, 32'hc155b896, 32'hc19a8364, 32'hc0837372};
test_output[27184:27191] = '{32'h0, 32'h4280bc48, 32'h422b0ec3, 32'h41595f8c, 32'h42528b0e, 32'h0, 32'h0, 32'h0};
test_input[27192:27199] = '{32'h41557730, 32'hc2c72438, 32'h41dd051b, 32'hc24b20f1, 32'hc26a70a6, 32'h4270b6cf, 32'h42b3e685, 32'h413ef627};
test_output[27192:27199] = '{32'h41557730, 32'h0, 32'h41dd051b, 32'h0, 32'h0, 32'h4270b6cf, 32'h42b3e685, 32'h413ef627};
test_input[27200:27207] = '{32'h42904a08, 32'hc13a731b, 32'hc2ac3c04, 32'hc22b5f39, 32'hc23a63ba, 32'hc224d4d1, 32'h3f6f6111, 32'hc294b7d5};
test_output[27200:27207] = '{32'h42904a08, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3f6f6111, 32'h0};
test_input[27208:27215] = '{32'h42925a28, 32'hc288d206, 32'h408f0e80, 32'h423f8633, 32'h428303db, 32'hc2a2b643, 32'h42584730, 32'hc2aa8436};
test_output[27208:27215] = '{32'h42925a28, 32'h0, 32'h408f0e80, 32'h423f8633, 32'h428303db, 32'h0, 32'h42584730, 32'h0};
test_input[27216:27223] = '{32'hc1dd8f2b, 32'h4292a31c, 32'h42ab633e, 32'hc25bc0e8, 32'hc2a1f05a, 32'hc2ac925e, 32'h40f730e5, 32'hc2812216};
test_output[27216:27223] = '{32'h0, 32'h4292a31c, 32'h42ab633e, 32'h0, 32'h0, 32'h0, 32'h40f730e5, 32'h0};
test_input[27224:27231] = '{32'hc23373be, 32'hc23acbc6, 32'h41b2c4e9, 32'hc2389727, 32'hc2c61134, 32'h423fae16, 32'h425fa727, 32'h412da855};
test_output[27224:27231] = '{32'h0, 32'h0, 32'h41b2c4e9, 32'h0, 32'h0, 32'h423fae16, 32'h425fa727, 32'h412da855};
test_input[27232:27239] = '{32'hc2bbd7a0, 32'hc170175d, 32'hc298d572, 32'h41df173b, 32'hc24b3b2d, 32'h4284da15, 32'hc0bb3d6b, 32'hc0187d0a};
test_output[27232:27239] = '{32'h0, 32'h0, 32'h0, 32'h41df173b, 32'h0, 32'h4284da15, 32'h0, 32'h0};
test_input[27240:27247] = '{32'h414c4d00, 32'h42c7523d, 32'h42b15270, 32'hc1a5a618, 32'h41fa09a5, 32'hc2570dba, 32'hc2773dd5, 32'h42ba726c};
test_output[27240:27247] = '{32'h414c4d00, 32'h42c7523d, 32'h42b15270, 32'h0, 32'h41fa09a5, 32'h0, 32'h0, 32'h42ba726c};
test_input[27248:27255] = '{32'hc12ed729, 32'hc06e4e96, 32'h41f787ff, 32'hc26315cb, 32'hc23b1e67, 32'h426f7932, 32'hc238c171, 32'hc20e8064};
test_output[27248:27255] = '{32'h0, 32'h0, 32'h41f787ff, 32'h0, 32'h0, 32'h426f7932, 32'h0, 32'h0};
test_input[27256:27263] = '{32'hc0114757, 32'h4284efe1, 32'hc23774cc, 32'h41f2e6db, 32'h411d840f, 32'h42b9fe7f, 32'h42b58ebf, 32'hc2924af6};
test_output[27256:27263] = '{32'h0, 32'h4284efe1, 32'h0, 32'h41f2e6db, 32'h411d840f, 32'h42b9fe7f, 32'h42b58ebf, 32'h0};
test_input[27264:27271] = '{32'h420c8cd3, 32'h42917eb6, 32'h42a5d686, 32'hc1d41e8a, 32'h4298f088, 32'hc1c39ccb, 32'h4089ea8b, 32'h42c39ddb};
test_output[27264:27271] = '{32'h420c8cd3, 32'h42917eb6, 32'h42a5d686, 32'h0, 32'h4298f088, 32'h0, 32'h4089ea8b, 32'h42c39ddb};
test_input[27272:27279] = '{32'hc20c6c3b, 32'h41ea191b, 32'h4298b8c3, 32'h40097791, 32'h427c82f4, 32'h421e07bd, 32'h42452786, 32'h40062f25};
test_output[27272:27279] = '{32'h0, 32'h41ea191b, 32'h4298b8c3, 32'h40097791, 32'h427c82f4, 32'h421e07bd, 32'h42452786, 32'h40062f25};
test_input[27280:27287] = '{32'hc10d7798, 32'h413e4f65, 32'h417ff138, 32'hc21eaa3c, 32'h42124179, 32'hc2a92963, 32'h3fd30692, 32'hc2863f75};
test_output[27280:27287] = '{32'h0, 32'h413e4f65, 32'h417ff138, 32'h0, 32'h42124179, 32'h0, 32'h3fd30692, 32'h0};
test_input[27288:27295] = '{32'h40902df7, 32'hc2885e64, 32'h42b9a241, 32'hc0825238, 32'h42981ba2, 32'h428ba36c, 32'hc14997e9, 32'hc265a267};
test_output[27288:27295] = '{32'h40902df7, 32'h0, 32'h42b9a241, 32'h0, 32'h42981ba2, 32'h428ba36c, 32'h0, 32'h0};
test_input[27296:27303] = '{32'h42865857, 32'h42c1feab, 32'hc015a00b, 32'h42acf383, 32'h429b812e, 32'h418b4dad, 32'hc2553a01, 32'hc28d940f};
test_output[27296:27303] = '{32'h42865857, 32'h42c1feab, 32'h0, 32'h42acf383, 32'h429b812e, 32'h418b4dad, 32'h0, 32'h0};
test_input[27304:27311] = '{32'h4215267a, 32'h425d74c2, 32'hc2490a75, 32'hc22a9fd4, 32'hc18db01e, 32'hc2941bc6, 32'hc29a7312, 32'h41fe3880};
test_output[27304:27311] = '{32'h4215267a, 32'h425d74c2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41fe3880};
test_input[27312:27319] = '{32'h42a73e80, 32'h41a16cec, 32'h42aa9df5, 32'hc2224a19, 32'h42a1569c, 32'h42ad4612, 32'hc03d8959, 32'h423fa7cf};
test_output[27312:27319] = '{32'h42a73e80, 32'h41a16cec, 32'h42aa9df5, 32'h0, 32'h42a1569c, 32'h42ad4612, 32'h0, 32'h423fa7cf};
test_input[27320:27327] = '{32'hc298a836, 32'h427d8694, 32'h3ffa546d, 32'hc288ac46, 32'h42a9bcbb, 32'hc25f4b9b, 32'h42afb631, 32'hc1acb5b8};
test_output[27320:27327] = '{32'h0, 32'h427d8694, 32'h3ffa546d, 32'h0, 32'h42a9bcbb, 32'h0, 32'h42afb631, 32'h0};
test_input[27328:27335] = '{32'h422a4a8b, 32'hc1a7b533, 32'hc2192418, 32'hc2527664, 32'h42b1b2e0, 32'h428943d1, 32'hc2aeec9a, 32'h421f9f87};
test_output[27328:27335] = '{32'h422a4a8b, 32'h0, 32'h0, 32'h0, 32'h42b1b2e0, 32'h428943d1, 32'h0, 32'h421f9f87};
test_input[27336:27343] = '{32'h4262db7c, 32'hc2231ab0, 32'hc28a7457, 32'hc17e492d, 32'hc27ac3b3, 32'hc202bdfc, 32'h423a8e68, 32'hc25d7598};
test_output[27336:27343] = '{32'h4262db7c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423a8e68, 32'h0};
test_input[27344:27351] = '{32'hc20c7b58, 32'h42ac7e54, 32'h42b633e4, 32'hc1bfec15, 32'hc089c8f6, 32'h42722898, 32'h408bd4ac, 32'h41907008};
test_output[27344:27351] = '{32'h0, 32'h42ac7e54, 32'h42b633e4, 32'h0, 32'h0, 32'h42722898, 32'h408bd4ac, 32'h41907008};
test_input[27352:27359] = '{32'hc2146e61, 32'hc15a6008, 32'hc2c0e350, 32'h42849ccc, 32'h412c5458, 32'h42807c60, 32'hc1e89bd3, 32'h42b61386};
test_output[27352:27359] = '{32'h0, 32'h0, 32'h0, 32'h42849ccc, 32'h412c5458, 32'h42807c60, 32'h0, 32'h42b61386};
test_input[27360:27367] = '{32'hc253e697, 32'h421be33a, 32'hc0ae1e4d, 32'hc278f1dc, 32'h42a6ef38, 32'hc2861caa, 32'h42451671, 32'h42a7d4e5};
test_output[27360:27367] = '{32'h0, 32'h421be33a, 32'h0, 32'h0, 32'h42a6ef38, 32'h0, 32'h42451671, 32'h42a7d4e5};
test_input[27368:27375] = '{32'h40e013bf, 32'h42c1878a, 32'h4277295d, 32'hc13119ae, 32'hc26f455b, 32'hc2b23750, 32'hc19a5ab1, 32'hc26bfd38};
test_output[27368:27375] = '{32'h40e013bf, 32'h42c1878a, 32'h4277295d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27376:27383] = '{32'hc110d8c1, 32'h42b962c1, 32'h422868ef, 32'hc196d740, 32'hc2033eb9, 32'h428861f9, 32'h41438dcc, 32'h410a480a};
test_output[27376:27383] = '{32'h0, 32'h42b962c1, 32'h422868ef, 32'h0, 32'h0, 32'h428861f9, 32'h41438dcc, 32'h410a480a};
test_input[27384:27391] = '{32'h428a7725, 32'h428929d5, 32'h4249017c, 32'hc2c2b9a8, 32'hc29c5512, 32'hc29f7662, 32'hc293411e, 32'h42b8f3ee};
test_output[27384:27391] = '{32'h428a7725, 32'h428929d5, 32'h4249017c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b8f3ee};
test_input[27392:27399] = '{32'h41b2fa7b, 32'h4016d3b4, 32'h4263de59, 32'hc298914a, 32'hc13d1353, 32'h42ba3846, 32'h40577ab9, 32'h42a24d0c};
test_output[27392:27399] = '{32'h41b2fa7b, 32'h4016d3b4, 32'h4263de59, 32'h0, 32'h0, 32'h42ba3846, 32'h40577ab9, 32'h42a24d0c};
test_input[27400:27407] = '{32'hc0025a30, 32'hc1d92c32, 32'hc2b81fc8, 32'hc210bddd, 32'h4264525d, 32'hc0dd9076, 32'hc096d84f, 32'hc24d9654};
test_output[27400:27407] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4264525d, 32'h0, 32'h0, 32'h0};
test_input[27408:27415] = '{32'h410ee18e, 32'h427bf135, 32'h4194825f, 32'hc141c19d, 32'h4182e2ec, 32'h4286bfcd, 32'hc142f46c, 32'h41940840};
test_output[27408:27415] = '{32'h410ee18e, 32'h427bf135, 32'h4194825f, 32'h0, 32'h4182e2ec, 32'h4286bfcd, 32'h0, 32'h41940840};
test_input[27416:27423] = '{32'h42b70dce, 32'h423694f7, 32'h42970cc1, 32'hc0c1ba26, 32'hc207f724, 32'h40ac68df, 32'h4251f941, 32'hc2832502};
test_output[27416:27423] = '{32'h42b70dce, 32'h423694f7, 32'h42970cc1, 32'h0, 32'h0, 32'h40ac68df, 32'h4251f941, 32'h0};
test_input[27424:27431] = '{32'hc299bc38, 32'hc198117c, 32'hc10ec43f, 32'h42ad2c91, 32'h42c4f0e6, 32'hc2a0e086, 32'h426ea449, 32'h428775ce};
test_output[27424:27431] = '{32'h0, 32'h0, 32'h0, 32'h42ad2c91, 32'h42c4f0e6, 32'h0, 32'h426ea449, 32'h428775ce};
test_input[27432:27439] = '{32'h41fff83c, 32'hc2979a33, 32'hc206f002, 32'h41ac233b, 32'h405bf6bb, 32'hc1fd4ec4, 32'hc231a270, 32'h428bd648};
test_output[27432:27439] = '{32'h41fff83c, 32'h0, 32'h0, 32'h41ac233b, 32'h405bf6bb, 32'h0, 32'h0, 32'h428bd648};
test_input[27440:27447] = '{32'hc2c4dd12, 32'hc27d901f, 32'hc2a98761, 32'h42c6f384, 32'hc23ef8d1, 32'hc28666d4, 32'hc2bed25f, 32'hc28bb53a};
test_output[27440:27447] = '{32'h0, 32'h0, 32'h0, 32'h42c6f384, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27448:27455] = '{32'h42422002, 32'h42bac0f8, 32'hc1e1984e, 32'hc211a33c, 32'h429f7fe5, 32'h4283bd4a, 32'hc158c880, 32'hc0c47e1c};
test_output[27448:27455] = '{32'h42422002, 32'h42bac0f8, 32'h0, 32'h0, 32'h429f7fe5, 32'h4283bd4a, 32'h0, 32'h0};
test_input[27456:27463] = '{32'hc1d7b587, 32'h42b18f20, 32'hc1af26e0, 32'hc1054dca, 32'h42619d13, 32'h42bbb4e0, 32'h4160d1b2, 32'hc28a0704};
test_output[27456:27463] = '{32'h0, 32'h42b18f20, 32'h0, 32'h0, 32'h42619d13, 32'h42bbb4e0, 32'h4160d1b2, 32'h0};
test_input[27464:27471] = '{32'hc2893b3f, 32'hc25dc287, 32'h429d0db1, 32'hc1eb0dfe, 32'h425d3b88, 32'hc266d80a, 32'h42953fee, 32'h4223067d};
test_output[27464:27471] = '{32'h0, 32'h0, 32'h429d0db1, 32'h0, 32'h425d3b88, 32'h0, 32'h42953fee, 32'h4223067d};
test_input[27472:27479] = '{32'hc2bec325, 32'h4297d8e7, 32'hc0f54cea, 32'hc247dc90, 32'h420f2c08, 32'hc293811e, 32'h4247b1d1, 32'hc28822cd};
test_output[27472:27479] = '{32'h0, 32'h4297d8e7, 32'h0, 32'h0, 32'h420f2c08, 32'h0, 32'h4247b1d1, 32'h0};
test_input[27480:27487] = '{32'hc212adee, 32'hc1763373, 32'hc28d0629, 32'h41d7858b, 32'hc294ed1f, 32'hc1d7eec7, 32'h4257e977, 32'h425d91b0};
test_output[27480:27487] = '{32'h0, 32'h0, 32'h0, 32'h41d7858b, 32'h0, 32'h0, 32'h4257e977, 32'h425d91b0};
test_input[27488:27495] = '{32'h42ad9d80, 32'hc2081a53, 32'hc1db600b, 32'hc1a27e09, 32'hc1dffcf2, 32'h42903204, 32'hc1619c4d, 32'h42bfbf8f};
test_output[27488:27495] = '{32'h42ad9d80, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42903204, 32'h0, 32'h42bfbf8f};
test_input[27496:27503] = '{32'h4116281f, 32'h42c528f8, 32'hc2a176f8, 32'h428cb54a, 32'h424c2a54, 32'h42aaa8a4, 32'hc222cc3a, 32'h42203481};
test_output[27496:27503] = '{32'h4116281f, 32'h42c528f8, 32'h0, 32'h428cb54a, 32'h424c2a54, 32'h42aaa8a4, 32'h0, 32'h42203481};
test_input[27504:27511] = '{32'hc2488638, 32'hc2aa3e05, 32'h4245793d, 32'h41e3aaad, 32'hc23390a8, 32'hc24365fd, 32'h4189a927, 32'hbf08fbaa};
test_output[27504:27511] = '{32'h0, 32'h0, 32'h4245793d, 32'h41e3aaad, 32'h0, 32'h0, 32'h4189a927, 32'h0};
test_input[27512:27519] = '{32'hc189355f, 32'h42b92ae6, 32'h42972952, 32'h420b3e7e, 32'h429d0858, 32'hc11e1c09, 32'h426e9532, 32'hc21f5d22};
test_output[27512:27519] = '{32'h0, 32'h42b92ae6, 32'h42972952, 32'h420b3e7e, 32'h429d0858, 32'h0, 32'h426e9532, 32'h0};
test_input[27520:27527] = '{32'hc089d66f, 32'hc2663cdd, 32'h3ff138e1, 32'h4280332b, 32'hc28e9e1f, 32'hc2c7cae2, 32'hc250dff1, 32'h41102887};
test_output[27520:27527] = '{32'h0, 32'h0, 32'h3ff138e1, 32'h4280332b, 32'h0, 32'h0, 32'h0, 32'h41102887};
test_input[27528:27535] = '{32'hc1a1fe66, 32'h424b7027, 32'hc228a47f, 32'hc10d0a0e, 32'hc2667466, 32'h42932f46, 32'h428962a9, 32'hc2bf5737};
test_output[27528:27535] = '{32'h0, 32'h424b7027, 32'h0, 32'h0, 32'h0, 32'h42932f46, 32'h428962a9, 32'h0};
test_input[27536:27543] = '{32'h427ada66, 32'hc2a8a18e, 32'h41555d68, 32'hc1241f74, 32'h41430530, 32'h418ecb81, 32'hbf92a008, 32'hc1b46391};
test_output[27536:27543] = '{32'h427ada66, 32'h0, 32'h41555d68, 32'h0, 32'h41430530, 32'h418ecb81, 32'h0, 32'h0};
test_input[27544:27551] = '{32'hc200e035, 32'hc235cdf6, 32'hc2a80fb3, 32'hc020932b, 32'h4295afca, 32'hc1c90153, 32'h429a0838, 32'h42315686};
test_output[27544:27551] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4295afca, 32'h0, 32'h429a0838, 32'h42315686};
test_input[27552:27559] = '{32'h40c1ac9b, 32'hc1d074b8, 32'hc1c93471, 32'hc1e267df, 32'hc199e89a, 32'hc2201215, 32'h429ae2b4, 32'h4291282e};
test_output[27552:27559] = '{32'h40c1ac9b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429ae2b4, 32'h4291282e};
test_input[27560:27567] = '{32'hc2510aac, 32'hc2b39d3f, 32'h4102d71e, 32'hc108f181, 32'h41158690, 32'hc2c4bfed, 32'h42aeefd7, 32'hc18a3204};
test_output[27560:27567] = '{32'h0, 32'h0, 32'h4102d71e, 32'h0, 32'h41158690, 32'h0, 32'h42aeefd7, 32'h0};
test_input[27568:27575] = '{32'h4224d4ed, 32'h424ece0f, 32'hc0428c64, 32'hc2b5f721, 32'h42471a17, 32'hc1ab4c91, 32'h4244c33b, 32'h42789495};
test_output[27568:27575] = '{32'h4224d4ed, 32'h424ece0f, 32'h0, 32'h0, 32'h42471a17, 32'h0, 32'h4244c33b, 32'h42789495};
test_input[27576:27583] = '{32'hc2b0aa98, 32'hc29a4d8a, 32'hc2931a7d, 32'hc224656f, 32'h423a740b, 32'hc208fac7, 32'hc1ac0249, 32'hc1761bae};
test_output[27576:27583] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h423a740b, 32'h0, 32'h0, 32'h0};
test_input[27584:27591] = '{32'hc1e0137c, 32'h40befe04, 32'h423d7f8d, 32'hc242b84a, 32'hc1a0b7a6, 32'hc225c279, 32'hc252c9fb, 32'hc24cbfeb};
test_output[27584:27591] = '{32'h0, 32'h40befe04, 32'h423d7f8d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27592:27599] = '{32'h41111b64, 32'h40aa20e9, 32'hc246bcd9, 32'h41d7d854, 32'hc15f9a41, 32'h42af5d00, 32'h413754fe, 32'h3f9e8a34};
test_output[27592:27599] = '{32'h41111b64, 32'h40aa20e9, 32'h0, 32'h41d7d854, 32'h0, 32'h42af5d00, 32'h413754fe, 32'h3f9e8a34};
test_input[27600:27607] = '{32'h4295868c, 32'hbfef4190, 32'h419f226d, 32'h427c0b7e, 32'h4205ef44, 32'hc2adb375, 32'h428c7dd6, 32'h40793669};
test_output[27600:27607] = '{32'h4295868c, 32'h0, 32'h419f226d, 32'h427c0b7e, 32'h4205ef44, 32'h0, 32'h428c7dd6, 32'h40793669};
test_input[27608:27615] = '{32'hc2c361d7, 32'hc1ea2055, 32'hc2a47ecb, 32'h427f97c7, 32'h421d10c2, 32'hc2a09fcc, 32'h4135908f, 32'h41876102};
test_output[27608:27615] = '{32'h0, 32'h0, 32'h0, 32'h427f97c7, 32'h421d10c2, 32'h0, 32'h4135908f, 32'h41876102};
test_input[27616:27623] = '{32'h422c910e, 32'h42a87fb7, 32'h4105476d, 32'hc1815e2b, 32'hc1f4152b, 32'h42a7ada6, 32'hc1b5a4c7, 32'hc1af9f30};
test_output[27616:27623] = '{32'h422c910e, 32'h42a87fb7, 32'h4105476d, 32'h0, 32'h0, 32'h42a7ada6, 32'h0, 32'h0};
test_input[27624:27631] = '{32'h427802a1, 32'h42a5db6f, 32'hc28900f8, 32'hc290b18d, 32'hc2933eef, 32'hc23b76b3, 32'h3f27ef47, 32'hc29bfe26};
test_output[27624:27631] = '{32'h427802a1, 32'h42a5db6f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3f27ef47, 32'h0};
test_input[27632:27639] = '{32'hc0b379df, 32'hc2379338, 32'h428cbba9, 32'hc25bef95, 32'h41b41eca, 32'hc29da75a, 32'h41c2c00f, 32'hc2419771};
test_output[27632:27639] = '{32'h0, 32'h0, 32'h428cbba9, 32'h0, 32'h41b41eca, 32'h0, 32'h41c2c00f, 32'h0};
test_input[27640:27647] = '{32'h41866e6e, 32'hc1e14291, 32'hc2955003, 32'h42282c50, 32'hc29f3433, 32'h42b5d7eb, 32'h3fe2a15c, 32'hc282ca41};
test_output[27640:27647] = '{32'h41866e6e, 32'h0, 32'h0, 32'h42282c50, 32'h0, 32'h42b5d7eb, 32'h3fe2a15c, 32'h0};
test_input[27648:27655] = '{32'h4243dc36, 32'h3faeaf8a, 32'h42a47850, 32'hc266cdcf, 32'hc28ea121, 32'h41f53033, 32'hbec66404, 32'hbf7853de};
test_output[27648:27655] = '{32'h4243dc36, 32'h3faeaf8a, 32'h42a47850, 32'h0, 32'h0, 32'h41f53033, 32'h0, 32'h0};
test_input[27656:27663] = '{32'h4241d0df, 32'hc291b1e2, 32'h416f610e, 32'h42b34c49, 32'hc20c37e1, 32'h4243d7ab, 32'hc255c715, 32'h42c17517};
test_output[27656:27663] = '{32'h4241d0df, 32'h0, 32'h416f610e, 32'h42b34c49, 32'h0, 32'h4243d7ab, 32'h0, 32'h42c17517};
test_input[27664:27671] = '{32'h419df931, 32'hc2327649, 32'hc20b31d6, 32'h427705bb, 32'h41acc355, 32'h415b30b4, 32'hc28de2b0, 32'hc29226f9};
test_output[27664:27671] = '{32'h419df931, 32'h0, 32'h0, 32'h427705bb, 32'h41acc355, 32'h415b30b4, 32'h0, 32'h0};
test_input[27672:27679] = '{32'hc2bff782, 32'hbf9b680e, 32'h423cbb3a, 32'hc26b9cd8, 32'h426f3395, 32'hc08a6473, 32'h40cdc363, 32'hc22f9840};
test_output[27672:27679] = '{32'h0, 32'h0, 32'h423cbb3a, 32'h0, 32'h426f3395, 32'h0, 32'h40cdc363, 32'h0};
test_input[27680:27687] = '{32'hc2b26c9b, 32'hc29ced27, 32'hc28722a4, 32'h428de666, 32'hc206497f, 32'h42ab11d0, 32'h41ed920e, 32'hc1b9e009};
test_output[27680:27687] = '{32'h0, 32'h0, 32'h0, 32'h428de666, 32'h0, 32'h42ab11d0, 32'h41ed920e, 32'h0};
test_input[27688:27695] = '{32'hc2c02bf1, 32'hc279e1ae, 32'h42607f7d, 32'hc1e39e06, 32'hc132694a, 32'h425abfa5, 32'h412c0a33, 32'hc1c9dc4e};
test_output[27688:27695] = '{32'h0, 32'h0, 32'h42607f7d, 32'h0, 32'h0, 32'h425abfa5, 32'h412c0a33, 32'h0};
test_input[27696:27703] = '{32'h4120432b, 32'h42ba45c3, 32'h4259aa23, 32'hc2c13363, 32'h4242a3da, 32'h42853f58, 32'hc2723dab, 32'hc22fe5cb};
test_output[27696:27703] = '{32'h4120432b, 32'h42ba45c3, 32'h4259aa23, 32'h0, 32'h4242a3da, 32'h42853f58, 32'h0, 32'h0};
test_input[27704:27711] = '{32'hc261a4dd, 32'h42284886, 32'hc1ea4e82, 32'h4291aca1, 32'h3f76fd48, 32'h424c905c, 32'hc2afa330, 32'hc17e5e7b};
test_output[27704:27711] = '{32'h0, 32'h42284886, 32'h0, 32'h4291aca1, 32'h3f76fd48, 32'h424c905c, 32'h0, 32'h0};
test_input[27712:27719] = '{32'h42c3fef8, 32'h42851f96, 32'hc0c9c8a6, 32'hc28c8faf, 32'hc28844b0, 32'hc10ce803, 32'hc26fa08e, 32'hc2147a71};
test_output[27712:27719] = '{32'h42c3fef8, 32'h42851f96, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27720:27727] = '{32'hc294297e, 32'hc29865f7, 32'h42a6c665, 32'h425f1261, 32'h426822b5, 32'hc255cacb, 32'h41286ebd, 32'hc2bd622a};
test_output[27720:27727] = '{32'h0, 32'h0, 32'h42a6c665, 32'h425f1261, 32'h426822b5, 32'h0, 32'h41286ebd, 32'h0};
test_input[27728:27735] = '{32'h42ac8ca8, 32'h409341b0, 32'h4253d3d9, 32'hbf2c01a4, 32'hc212691a, 32'hc2815415, 32'hc1fa7eeb, 32'h42b53a78};
test_output[27728:27735] = '{32'h42ac8ca8, 32'h409341b0, 32'h4253d3d9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b53a78};
test_input[27736:27743] = '{32'h423a9821, 32'hc23236e8, 32'h42b2ba5b, 32'h4254103c, 32'h4211c6d5, 32'h42abc6e2, 32'hc28f2ebb, 32'h41cb3b07};
test_output[27736:27743] = '{32'h423a9821, 32'h0, 32'h42b2ba5b, 32'h4254103c, 32'h4211c6d5, 32'h42abc6e2, 32'h0, 32'h41cb3b07};
test_input[27744:27751] = '{32'hc1fa918d, 32'h419b4260, 32'h428cd33e, 32'hc28f4386, 32'hc23fe7a1, 32'h424b0cb9, 32'h428afdf0, 32'h41467870};
test_output[27744:27751] = '{32'h0, 32'h419b4260, 32'h428cd33e, 32'h0, 32'h0, 32'h424b0cb9, 32'h428afdf0, 32'h41467870};
test_input[27752:27759] = '{32'hc203142d, 32'h42ac19f1, 32'h420f4879, 32'hc225be6b, 32'hc2523a94, 32'h421ea938, 32'h3f0bd9ac, 32'hc272e1b4};
test_output[27752:27759] = '{32'h0, 32'h42ac19f1, 32'h420f4879, 32'h0, 32'h0, 32'h421ea938, 32'h3f0bd9ac, 32'h0};
test_input[27760:27767] = '{32'hc27bca91, 32'h4219b90a, 32'hc084547b, 32'hc13ed983, 32'h4212cc52, 32'hc1fae7ab, 32'hc183b129, 32'hc2a8b0f1};
test_output[27760:27767] = '{32'h0, 32'h4219b90a, 32'h0, 32'h0, 32'h4212cc52, 32'h0, 32'h0, 32'h0};
test_input[27768:27775] = '{32'hc2356bba, 32'hc2b337d5, 32'h41dbb223, 32'hc21e219f, 32'h425f8d7b, 32'hc290d47d, 32'hbf63beb0, 32'h42b45b37};
test_output[27768:27775] = '{32'h0, 32'h0, 32'h41dbb223, 32'h0, 32'h425f8d7b, 32'h0, 32'h0, 32'h42b45b37};
test_input[27776:27783] = '{32'h41242e82, 32'hc1e86855, 32'hc2984c6d, 32'hc2c42ee3, 32'h420ad2b2, 32'h426e9701, 32'h42bb8510, 32'hc2136863};
test_output[27776:27783] = '{32'h41242e82, 32'h0, 32'h0, 32'h0, 32'h420ad2b2, 32'h426e9701, 32'h42bb8510, 32'h0};
test_input[27784:27791] = '{32'hc2a3d009, 32'hc1a36aeb, 32'h41e3e3c6, 32'h41ae1ed7, 32'h4247e0f0, 32'hc1563f8c, 32'h42c2aab3, 32'hc2a0d2b7};
test_output[27784:27791] = '{32'h0, 32'h0, 32'h41e3e3c6, 32'h41ae1ed7, 32'h4247e0f0, 32'h0, 32'h42c2aab3, 32'h0};
test_input[27792:27799] = '{32'hbfd3826b, 32'hc27eb537, 32'h4284f651, 32'h42bc7be3, 32'h421ebbfc, 32'h4174aa41, 32'hc253f90a, 32'hc2950375};
test_output[27792:27799] = '{32'h0, 32'h0, 32'h4284f651, 32'h42bc7be3, 32'h421ebbfc, 32'h4174aa41, 32'h0, 32'h0};
test_input[27800:27807] = '{32'h42c6661d, 32'h402c3ccf, 32'hc23c4368, 32'hc2b4e24a, 32'h42b8f2b6, 32'h419ef0be, 32'hbfb66091, 32'h411c547c};
test_output[27800:27807] = '{32'h42c6661d, 32'h402c3ccf, 32'h0, 32'h0, 32'h42b8f2b6, 32'h419ef0be, 32'h0, 32'h411c547c};
test_input[27808:27815] = '{32'hc13df893, 32'h42a29d8a, 32'hc2a515b1, 32'h418a116c, 32'hc20cccf9, 32'h3f8c7e79, 32'h4243b20a, 32'h4284e462};
test_output[27808:27815] = '{32'h0, 32'h42a29d8a, 32'h0, 32'h418a116c, 32'h0, 32'h3f8c7e79, 32'h4243b20a, 32'h4284e462};
test_input[27816:27823] = '{32'h42945ec4, 32'hc234b6f8, 32'hc101d88a, 32'hc1f2086b, 32'hc2722dbc, 32'hc29e51e8, 32'h42c570ca, 32'hc280ffa9};
test_output[27816:27823] = '{32'h42945ec4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c570ca, 32'h0};
test_input[27824:27831] = '{32'hc26fc69d, 32'h427c3bdb, 32'hc23d3fb1, 32'h42c3e2c5, 32'h41b9a926, 32'h41968f06, 32'hc2aa9ab7, 32'hc218da2a};
test_output[27824:27831] = '{32'h0, 32'h427c3bdb, 32'h0, 32'h42c3e2c5, 32'h41b9a926, 32'h41968f06, 32'h0, 32'h0};
test_input[27832:27839] = '{32'h42b99539, 32'hc2ae6b48, 32'hc29b837a, 32'hc2aaf0b0, 32'h424cf69b, 32'h42c6484d, 32'h41802e4a, 32'h4289cbb3};
test_output[27832:27839] = '{32'h42b99539, 32'h0, 32'h0, 32'h0, 32'h424cf69b, 32'h42c6484d, 32'h41802e4a, 32'h4289cbb3};
test_input[27840:27847] = '{32'hc2bc4461, 32'h41461ad1, 32'h41d0979a, 32'h42938de4, 32'hc1366ecb, 32'h427ee91f, 32'h423199f1, 32'hc2c34d77};
test_output[27840:27847] = '{32'h0, 32'h41461ad1, 32'h41d0979a, 32'h42938de4, 32'h0, 32'h427ee91f, 32'h423199f1, 32'h0};
test_input[27848:27855] = '{32'h423329de, 32'hc2ad8cef, 32'h42c0f464, 32'h42588d54, 32'h42784792, 32'hc29a2961, 32'h42bf9394, 32'h42a53605};
test_output[27848:27855] = '{32'h423329de, 32'h0, 32'h42c0f464, 32'h42588d54, 32'h42784792, 32'h0, 32'h42bf9394, 32'h42a53605};
test_input[27856:27863] = '{32'h40c18c5e, 32'h41ab7b2d, 32'h4247277c, 32'hc2b36503, 32'h42518072, 32'hc0bb6e0e, 32'hc20f8062, 32'h4261fb70};
test_output[27856:27863] = '{32'h40c18c5e, 32'h41ab7b2d, 32'h4247277c, 32'h0, 32'h42518072, 32'h0, 32'h0, 32'h4261fb70};
test_input[27864:27871] = '{32'h426109c2, 32'hc2599f8d, 32'hc1ab40d2, 32'hc1e59807, 32'hc243d107, 32'hc285dfd0, 32'hc28e58fc, 32'hc210f3c6};
test_output[27864:27871] = '{32'h426109c2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27872:27879] = '{32'h42130e3d, 32'h428ed632, 32'hc21797b0, 32'hc20a0740, 32'hc297dd15, 32'h3fdbea9c, 32'hc283adfd, 32'h412d0bfa};
test_output[27872:27879] = '{32'h42130e3d, 32'h428ed632, 32'h0, 32'h0, 32'h0, 32'h3fdbea9c, 32'h0, 32'h412d0bfa};
test_input[27880:27887] = '{32'h42b30b88, 32'hc185fd2f, 32'h42b3907b, 32'hc29b6553, 32'h42845f73, 32'h429507da, 32'h42aeab9c, 32'hc2a2b3b6};
test_output[27880:27887] = '{32'h42b30b88, 32'h0, 32'h42b3907b, 32'h0, 32'h42845f73, 32'h429507da, 32'h42aeab9c, 32'h0};
test_input[27888:27895] = '{32'h4246e927, 32'hc202df3e, 32'h425c1de1, 32'hc2930703, 32'h42184b5f, 32'hc251a770, 32'h4279e20e, 32'hc1aa9be2};
test_output[27888:27895] = '{32'h4246e927, 32'h0, 32'h425c1de1, 32'h0, 32'h42184b5f, 32'h0, 32'h4279e20e, 32'h0};
test_input[27896:27903] = '{32'hc18b8035, 32'h42bcd7a5, 32'hc07dfcc2, 32'h42180427, 32'h41b626ce, 32'hc2b9d41c, 32'h41326a89, 32'h420e848b};
test_output[27896:27903] = '{32'h0, 32'h42bcd7a5, 32'h0, 32'h42180427, 32'h41b626ce, 32'h0, 32'h41326a89, 32'h420e848b};
test_input[27904:27911] = '{32'h429a4dae, 32'h41092736, 32'h4096ea82, 32'hc24d95ce, 32'h42815d0d, 32'h41e306ee, 32'hc0de086b, 32'h425ba90b};
test_output[27904:27911] = '{32'h429a4dae, 32'h41092736, 32'h4096ea82, 32'h0, 32'h42815d0d, 32'h41e306ee, 32'h0, 32'h425ba90b};
test_input[27912:27919] = '{32'hc127e93b, 32'h428dcdf2, 32'hc0fe7fda, 32'h40a5587c, 32'hc2052eb0, 32'hc1ca9f8b, 32'hc0644f45, 32'h4252c566};
test_output[27912:27919] = '{32'h0, 32'h428dcdf2, 32'h0, 32'h40a5587c, 32'h0, 32'h0, 32'h0, 32'h4252c566};
test_input[27920:27927] = '{32'h4245832a, 32'h40beede6, 32'hc0d5739e, 32'h409bbed6, 32'h428179c8, 32'h422e1d98, 32'hc2791ac8, 32'h40e9182b};
test_output[27920:27927] = '{32'h4245832a, 32'h40beede6, 32'h0, 32'h409bbed6, 32'h428179c8, 32'h422e1d98, 32'h0, 32'h40e9182b};
test_input[27928:27935] = '{32'h41a7f2e7, 32'h42a03338, 32'h423fccff, 32'hc29b99c8, 32'hc2888a99, 32'hc2a74801, 32'hc29feb44, 32'hc17c3142};
test_output[27928:27935] = '{32'h41a7f2e7, 32'h42a03338, 32'h423fccff, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27936:27943] = '{32'hc1e27716, 32'hc2b9d780, 32'hc18d3f5c, 32'hc13811f4, 32'h42ae98dd, 32'h41ba056d, 32'h42316c84, 32'hc2a11e81};
test_output[27936:27943] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42ae98dd, 32'h41ba056d, 32'h42316c84, 32'h0};
test_input[27944:27951] = '{32'hc247a3b5, 32'hc1befc24, 32'h42b61790, 32'hc1ce0652, 32'hc2629381, 32'hc20f7303, 32'hc2b599d3, 32'h425b2fc7};
test_output[27944:27951] = '{32'h0, 32'h0, 32'h42b61790, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425b2fc7};
test_input[27952:27959] = '{32'h42be8679, 32'hc2389703, 32'h42c1faef, 32'hc1fab134, 32'h421b4349, 32'h41e93044, 32'h4240dc97, 32'h42aae0eb};
test_output[27952:27959] = '{32'h42be8679, 32'h0, 32'h42c1faef, 32'h0, 32'h421b4349, 32'h41e93044, 32'h4240dc97, 32'h42aae0eb};
test_input[27960:27967] = '{32'hc2621e8c, 32'h42272260, 32'hc2a2cc1f, 32'hc21c1da3, 32'hc200ed47, 32'h41a67efa, 32'hc2beffa0, 32'hc13d9efb};
test_output[27960:27967] = '{32'h0, 32'h42272260, 32'h0, 32'h0, 32'h0, 32'h41a67efa, 32'h0, 32'h0};
test_input[27968:27975] = '{32'hc289d047, 32'h421621e6, 32'hc250d735, 32'hc19dd56a, 32'h415cd0ca, 32'hc138a983, 32'h42c69334, 32'hc2bed94f};
test_output[27968:27975] = '{32'h0, 32'h421621e6, 32'h0, 32'h0, 32'h415cd0ca, 32'h0, 32'h42c69334, 32'h0};
test_input[27976:27983] = '{32'hc2025c91, 32'hc05dce52, 32'hc23a032e, 32'h42840c86, 32'hc197c88d, 32'hbcfa026a, 32'h42851b48, 32'hc2171ff9};
test_output[27976:27983] = '{32'h0, 32'h0, 32'h0, 32'h42840c86, 32'h0, 32'h0, 32'h42851b48, 32'h0};
test_input[27984:27991] = '{32'hc1d9a58d, 32'hc14d21db, 32'h42893c7c, 32'h426b1a37, 32'h42a3fea7, 32'hc0cc8706, 32'hc2357c0b, 32'h427dabf5};
test_output[27984:27991] = '{32'h0, 32'h0, 32'h42893c7c, 32'h426b1a37, 32'h42a3fea7, 32'h0, 32'h0, 32'h427dabf5};
test_input[27992:27999] = '{32'hc1e142b2, 32'hc1a9a983, 32'h41b480ee, 32'hc2b3bb04, 32'h4257843e, 32'h41e96cf6, 32'h41c82baa, 32'h422aa56f};
test_output[27992:27999] = '{32'h0, 32'h0, 32'h41b480ee, 32'h0, 32'h4257843e, 32'h41e96cf6, 32'h41c82baa, 32'h422aa56f};
test_input[28000:28007] = '{32'hc25faead, 32'hc0c3b626, 32'h418e0d8b, 32'h42806c7f, 32'hc29f070e, 32'h40c37ad9, 32'h423badeb, 32'hc263d3f9};
test_output[28000:28007] = '{32'h0, 32'h0, 32'h418e0d8b, 32'h42806c7f, 32'h0, 32'h40c37ad9, 32'h423badeb, 32'h0};
test_input[28008:28015] = '{32'h42c0c4a9, 32'h420cac55, 32'hc2c3b8ff, 32'hc2acfdeb, 32'h428c51d0, 32'h408d525b, 32'h42a61105, 32'hc299c779};
test_output[28008:28015] = '{32'h42c0c4a9, 32'h420cac55, 32'h0, 32'h0, 32'h428c51d0, 32'h408d525b, 32'h42a61105, 32'h0};
test_input[28016:28023] = '{32'hc2c71f2c, 32'hc28e88d7, 32'hc2740454, 32'hc2a91467, 32'hc24c3f55, 32'h41ee420b, 32'hc23bd679, 32'h42a45190};
test_output[28016:28023] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ee420b, 32'h0, 32'h42a45190};
test_input[28024:28031] = '{32'hc17b6829, 32'h421a247d, 32'hc0d0bb47, 32'h40ec4c87, 32'hc2c2755f, 32'h421ce5e8, 32'hc051f771, 32'hc277bf54};
test_output[28024:28031] = '{32'h0, 32'h421a247d, 32'h0, 32'h40ec4c87, 32'h0, 32'h421ce5e8, 32'h0, 32'h0};
test_input[28032:28039] = '{32'h4208e84d, 32'h42195249, 32'hc0b36e0d, 32'h425cd5f3, 32'hc1b4fda9, 32'hc24c6186, 32'hc05e8445, 32'h42a4f7b9};
test_output[28032:28039] = '{32'h4208e84d, 32'h42195249, 32'h0, 32'h425cd5f3, 32'h0, 32'h0, 32'h0, 32'h42a4f7b9};
test_input[28040:28047] = '{32'hc18c9c76, 32'hc2732897, 32'hc1c5c4e7, 32'h4279d879, 32'hc2bec316, 32'hc1b64f7a, 32'h41e5e360, 32'h4232cb45};
test_output[28040:28047] = '{32'h0, 32'h0, 32'h0, 32'h4279d879, 32'h0, 32'h0, 32'h41e5e360, 32'h4232cb45};
test_input[28048:28055] = '{32'hc27f8357, 32'h41a106c7, 32'hc2c44e4f, 32'hc20f6882, 32'hc28d7567, 32'hc28fc55b, 32'hc28adbac, 32'hc2762575};
test_output[28048:28055] = '{32'h0, 32'h41a106c7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28056:28063] = '{32'h4206f672, 32'h42862a0d, 32'h42a19b88, 32'hc233e29e, 32'h3ff80500, 32'h4285a765, 32'h4286b76f, 32'hc0b0d9b4};
test_output[28056:28063] = '{32'h4206f672, 32'h42862a0d, 32'h42a19b88, 32'h0, 32'h3ff80500, 32'h4285a765, 32'h4286b76f, 32'h0};
test_input[28064:28071] = '{32'hc2a0ff65, 32'h41881dc2, 32'hc24db568, 32'hc200c396, 32'h4294813e, 32'hc2adeb0c, 32'h40d32a88, 32'hc233be6d};
test_output[28064:28071] = '{32'h0, 32'h41881dc2, 32'h0, 32'h0, 32'h4294813e, 32'h0, 32'h40d32a88, 32'h0};
test_input[28072:28079] = '{32'hc2ba2b47, 32'h421e5e16, 32'hc28b6329, 32'h428b213d, 32'hc29b8e03, 32'h4148da95, 32'hc15604d1, 32'h4286fbb9};
test_output[28072:28079] = '{32'h0, 32'h421e5e16, 32'h0, 32'h428b213d, 32'h0, 32'h4148da95, 32'h0, 32'h4286fbb9};
test_input[28080:28087] = '{32'hc28ecf2a, 32'h41f68906, 32'hc2a17d98, 32'hc2094d04, 32'hc0a9eb7a, 32'h41bb3a94, 32'h4286aaf7, 32'hc1e95c57};
test_output[28080:28087] = '{32'h0, 32'h41f68906, 32'h0, 32'h0, 32'h0, 32'h41bb3a94, 32'h4286aaf7, 32'h0};
test_input[28088:28095] = '{32'hc20bc608, 32'hc1e3bb11, 32'h42b05f5e, 32'h4274482a, 32'h427b72d8, 32'hc2839f0b, 32'hc2b4ab25, 32'hc24908c2};
test_output[28088:28095] = '{32'h0, 32'h0, 32'h42b05f5e, 32'h4274482a, 32'h427b72d8, 32'h0, 32'h0, 32'h0};
test_input[28096:28103] = '{32'hc1af135d, 32'h42938211, 32'h427f6a77, 32'hbf1b402b, 32'hc2320787, 32'h428cb788, 32'hc1505a7d, 32'hc27d5c45};
test_output[28096:28103] = '{32'h0, 32'h42938211, 32'h427f6a77, 32'h0, 32'h0, 32'h428cb788, 32'h0, 32'h0};
test_input[28104:28111] = '{32'hc228ea88, 32'h4262a2d5, 32'h42a4dd93, 32'hc28d9230, 32'h42bb14e6, 32'h424a64fd, 32'h42b18993, 32'hc244099b};
test_output[28104:28111] = '{32'h0, 32'h4262a2d5, 32'h42a4dd93, 32'h0, 32'h42bb14e6, 32'h424a64fd, 32'h42b18993, 32'h0};
test_input[28112:28119] = '{32'hc252c281, 32'hc290989f, 32'hc2b9c7c8, 32'h4284ca30, 32'hc2a578c6, 32'hc1a5fa63, 32'hc28bac2f, 32'hc04b4c8b};
test_output[28112:28119] = '{32'h0, 32'h0, 32'h0, 32'h4284ca30, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28120:28127] = '{32'h3f1cf029, 32'h429e9da9, 32'hc280120e, 32'h427885da, 32'hc0e22c65, 32'h42695389, 32'h41f7469f, 32'hc22fbe75};
test_output[28120:28127] = '{32'h3f1cf029, 32'h429e9da9, 32'h0, 32'h427885da, 32'h0, 32'h42695389, 32'h41f7469f, 32'h0};
test_input[28128:28135] = '{32'hc28067f6, 32'hc14e58ac, 32'hc2900aa1, 32'hc29114c7, 32'hc0e660b3, 32'hc2b2c736, 32'hc2225cb9, 32'hc1d8e582};
test_output[28128:28135] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28136:28143] = '{32'h42ba2ee3, 32'h42735210, 32'h414381f3, 32'h41369270, 32'h41b6038a, 32'h42674f85, 32'hc2925d2d, 32'hc10ec5b9};
test_output[28136:28143] = '{32'h42ba2ee3, 32'h42735210, 32'h414381f3, 32'h41369270, 32'h41b6038a, 32'h42674f85, 32'h0, 32'h0};
test_input[28144:28151] = '{32'hc1eec88c, 32'hc2476940, 32'h42670cb1, 32'hc252d033, 32'h42c53050, 32'hc2b5aa5d, 32'h426c6c7d, 32'hc21c488e};
test_output[28144:28151] = '{32'h0, 32'h0, 32'h42670cb1, 32'h0, 32'h42c53050, 32'h0, 32'h426c6c7d, 32'h0};
test_input[28152:28159] = '{32'hc117fc57, 32'h42a78d87, 32'h409f3d7c, 32'hc2b2d018, 32'hc29ecf39, 32'h401a9ac9, 32'h4280da97, 32'hc2145ccb};
test_output[28152:28159] = '{32'h0, 32'h42a78d87, 32'h409f3d7c, 32'h0, 32'h0, 32'h401a9ac9, 32'h4280da97, 32'h0};
test_input[28160:28167] = '{32'hc2a1ab97, 32'h42b6f85c, 32'h4241e28a, 32'hc267a77f, 32'h427512dd, 32'h4127f92e, 32'hc1708a9e, 32'h4235df33};
test_output[28160:28167] = '{32'h0, 32'h42b6f85c, 32'h4241e28a, 32'h0, 32'h427512dd, 32'h4127f92e, 32'h0, 32'h4235df33};
test_input[28168:28175] = '{32'h423942a8, 32'hc2906538, 32'h415af3ac, 32'hc28d16ee, 32'hc2bf7825, 32'hc182e2f1, 32'h425117fc, 32'h42291b87};
test_output[28168:28175] = '{32'h423942a8, 32'h0, 32'h415af3ac, 32'h0, 32'h0, 32'h0, 32'h425117fc, 32'h42291b87};
test_input[28176:28183] = '{32'hc2656d94, 32'hc209ed93, 32'h425d4726, 32'hc286c676, 32'h4151db3d, 32'hc23276a3, 32'h429f3ecc, 32'hc2048030};
test_output[28176:28183] = '{32'h0, 32'h0, 32'h425d4726, 32'h0, 32'h4151db3d, 32'h0, 32'h429f3ecc, 32'h0};
test_input[28184:28191] = '{32'h4261b1d8, 32'h4275af64, 32'h4073035e, 32'h4277e7cd, 32'hc297b468, 32'h41a4473d, 32'hc2a727b7, 32'hc2c4d75c};
test_output[28184:28191] = '{32'h4261b1d8, 32'h4275af64, 32'h4073035e, 32'h4277e7cd, 32'h0, 32'h41a4473d, 32'h0, 32'h0};
test_input[28192:28199] = '{32'h4263c239, 32'hc29448b9, 32'h425a393b, 32'h41c12c5e, 32'hc271df84, 32'hc217a2fb, 32'h41e8cf7c, 32'h413c4d74};
test_output[28192:28199] = '{32'h4263c239, 32'h0, 32'h425a393b, 32'h41c12c5e, 32'h0, 32'h0, 32'h41e8cf7c, 32'h413c4d74};
test_input[28200:28207] = '{32'hc28fa108, 32'hc1215603, 32'hc282d372, 32'h40d8c9fa, 32'h420a405f, 32'hc18820bd, 32'h42763e6c, 32'h42b9e99e};
test_output[28200:28207] = '{32'h0, 32'h0, 32'h0, 32'h40d8c9fa, 32'h420a405f, 32'h0, 32'h42763e6c, 32'h42b9e99e};
test_input[28208:28215] = '{32'hc206a264, 32'h426cb2c7, 32'h3ff9b663, 32'h42b6e45a, 32'h42bd3116, 32'h4274d333, 32'h41989008, 32'h428089a5};
test_output[28208:28215] = '{32'h0, 32'h426cb2c7, 32'h3ff9b663, 32'h42b6e45a, 32'h42bd3116, 32'h4274d333, 32'h41989008, 32'h428089a5};
test_input[28216:28223] = '{32'hc283d5a8, 32'hc27a95b0, 32'hc2ade429, 32'hc1b33c89, 32'h41c23fc2, 32'h42c6ba4c, 32'hc23f48a8, 32'h42a909f2};
test_output[28216:28223] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41c23fc2, 32'h42c6ba4c, 32'h0, 32'h42a909f2};
test_input[28224:28231] = '{32'h40174c50, 32'hc17a62c6, 32'h419abefa, 32'hc0377090, 32'h422522a7, 32'h4213551b, 32'hc284f609, 32'h4226e67a};
test_output[28224:28231] = '{32'h40174c50, 32'h0, 32'h419abefa, 32'h0, 32'h422522a7, 32'h4213551b, 32'h0, 32'h4226e67a};
test_input[28232:28239] = '{32'hc14d79f5, 32'h42acf167, 32'h413d72a4, 32'hc2810c5a, 32'hc194d827, 32'hc224cbe5, 32'hc2970fb9, 32'hbf1f60a4};
test_output[28232:28239] = '{32'h0, 32'h42acf167, 32'h413d72a4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28240:28247] = '{32'h41e8a191, 32'h4260892e, 32'h42c5e21b, 32'hc2acfa16, 32'h4260ee1d, 32'h4162190e, 32'hc124be9e, 32'h428d9ea8};
test_output[28240:28247] = '{32'h41e8a191, 32'h4260892e, 32'h42c5e21b, 32'h0, 32'h4260ee1d, 32'h4162190e, 32'h0, 32'h428d9ea8};
test_input[28248:28255] = '{32'h422cbec7, 32'hc2855b6e, 32'h41bd0377, 32'hc295004b, 32'hc24cf92a, 32'hc2b191f1, 32'h4123c0f2, 32'hc1ef03a4};
test_output[28248:28255] = '{32'h422cbec7, 32'h0, 32'h41bd0377, 32'h0, 32'h0, 32'h0, 32'h4123c0f2, 32'h0};
test_input[28256:28263] = '{32'h42630e37, 32'h42130094, 32'h41049b35, 32'h427d0f99, 32'hbfc46b07, 32'hc2031c01, 32'h41b6b985, 32'hc20ed950};
test_output[28256:28263] = '{32'h42630e37, 32'h42130094, 32'h41049b35, 32'h427d0f99, 32'h0, 32'h0, 32'h41b6b985, 32'h0};
test_input[28264:28271] = '{32'h4225a453, 32'hc186b3ff, 32'hc26b9203, 32'h424dcd10, 32'h426356c6, 32'h424c46a2, 32'h42663901, 32'h42a8a65a};
test_output[28264:28271] = '{32'h4225a453, 32'h0, 32'h0, 32'h424dcd10, 32'h426356c6, 32'h424c46a2, 32'h42663901, 32'h42a8a65a};
test_input[28272:28279] = '{32'hc2afb067, 32'hc2af28ae, 32'hc0fd93c2, 32'h3fba3edb, 32'h4283514f, 32'hc2a4a165, 32'hc22b7c1e, 32'h42aad0ed};
test_output[28272:28279] = '{32'h0, 32'h0, 32'h0, 32'h3fba3edb, 32'h4283514f, 32'h0, 32'h0, 32'h42aad0ed};
test_input[28280:28287] = '{32'h428956f3, 32'h42138b32, 32'hc26bd0de, 32'hc2b15f3b, 32'hc277f1dc, 32'h42b60316, 32'h41f60070, 32'h40f1e153};
test_output[28280:28287] = '{32'h428956f3, 32'h42138b32, 32'h0, 32'h0, 32'h0, 32'h42b60316, 32'h41f60070, 32'h40f1e153};
test_input[28288:28295] = '{32'h41594d31, 32'hc29deda7, 32'h424ca4c2, 32'hc2587703, 32'h428e7ef0, 32'hc110eb66, 32'h4133e234, 32'h411abaa0};
test_output[28288:28295] = '{32'h41594d31, 32'h0, 32'h424ca4c2, 32'h0, 32'h428e7ef0, 32'h0, 32'h4133e234, 32'h411abaa0};
test_input[28296:28303] = '{32'hc27ebe3b, 32'hc088a3f9, 32'h40040e57, 32'h40f88779, 32'hc2aa820d, 32'h41e1eb3d, 32'hc27aacc5, 32'hc2243259};
test_output[28296:28303] = '{32'h0, 32'h0, 32'h40040e57, 32'h40f88779, 32'h0, 32'h41e1eb3d, 32'h0, 32'h0};
test_input[28304:28311] = '{32'hc24ca363, 32'h4282c00c, 32'h421811cd, 32'h41f5d1dd, 32'h42bbfeb9, 32'h412eca7a, 32'hc2556a78, 32'h421fe100};
test_output[28304:28311] = '{32'h0, 32'h4282c00c, 32'h421811cd, 32'h41f5d1dd, 32'h42bbfeb9, 32'h412eca7a, 32'h0, 32'h421fe100};
test_input[28312:28319] = '{32'h423f7026, 32'h4268008f, 32'hc242f584, 32'hc2aa62db, 32'hc02487a5, 32'h41caaef9, 32'hc2b765e7, 32'h4299ddc3};
test_output[28312:28319] = '{32'h423f7026, 32'h4268008f, 32'h0, 32'h0, 32'h0, 32'h41caaef9, 32'h0, 32'h4299ddc3};
test_input[28320:28327] = '{32'h4218d1d4, 32'h4249350d, 32'h427fd225, 32'hc2b63d1b, 32'hc238014b, 32'h4130334f, 32'h42b58176, 32'h427a47b1};
test_output[28320:28327] = '{32'h4218d1d4, 32'h4249350d, 32'h427fd225, 32'h0, 32'h0, 32'h4130334f, 32'h42b58176, 32'h427a47b1};
test_input[28328:28335] = '{32'hc1fcc198, 32'h427cce90, 32'h415a0259, 32'hc1ec2086, 32'hc198b100, 32'h4256cbe9, 32'hc2755d2e, 32'hc272038b};
test_output[28328:28335] = '{32'h0, 32'h427cce90, 32'h415a0259, 32'h0, 32'h0, 32'h4256cbe9, 32'h0, 32'h0};
test_input[28336:28343] = '{32'h419aad0d, 32'h41cb40ef, 32'h3e8e1e02, 32'hc2815cdc, 32'hc2873277, 32'hc201d3de, 32'hc18c9fca, 32'hc23eda5d};
test_output[28336:28343] = '{32'h419aad0d, 32'h41cb40ef, 32'h3e8e1e02, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28344:28351] = '{32'h42ba16a0, 32'hc29599fa, 32'hc2a9282a, 32'hc1ea9228, 32'hc1c760dd, 32'hc21a4491, 32'hc2a8a53f, 32'h42ab3ab0};
test_output[28344:28351] = '{32'h42ba16a0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ab3ab0};
test_input[28352:28359] = '{32'h41fe3c0a, 32'h425fa9dd, 32'hc290d251, 32'h42340c6b, 32'hc2c7e0e7, 32'hc2ab84fb, 32'h4232272a, 32'h419f6eeb};
test_output[28352:28359] = '{32'h41fe3c0a, 32'h425fa9dd, 32'h0, 32'h42340c6b, 32'h0, 32'h0, 32'h4232272a, 32'h419f6eeb};
test_input[28360:28367] = '{32'hc2364585, 32'hc2a5cf11, 32'h41cca9c7, 32'h42be1418, 32'hc0a52c87, 32'hc2943517, 32'h4299dfe2, 32'h423e727f};
test_output[28360:28367] = '{32'h0, 32'h0, 32'h41cca9c7, 32'h42be1418, 32'h0, 32'h0, 32'h4299dfe2, 32'h423e727f};
test_input[28368:28375] = '{32'h41dea5c4, 32'h42091d62, 32'hc2113f27, 32'h4245753b, 32'hc0cee7be, 32'hc2a475f8, 32'h429c39f5, 32'hc274679e};
test_output[28368:28375] = '{32'h41dea5c4, 32'h42091d62, 32'h0, 32'h4245753b, 32'h0, 32'h0, 32'h429c39f5, 32'h0};
test_input[28376:28383] = '{32'hc296b495, 32'h41eb5e83, 32'hc11be4c4, 32'h42427dd4, 32'hc2110d5c, 32'h428560ed, 32'hc282206d, 32'hc25a2b9b};
test_output[28376:28383] = '{32'h0, 32'h41eb5e83, 32'h0, 32'h42427dd4, 32'h0, 32'h428560ed, 32'h0, 32'h0};
test_input[28384:28391] = '{32'h427e64bf, 32'hc21ba7dc, 32'h41e8c863, 32'h428ad6cd, 32'hc1ea46f7, 32'hc1874ba6, 32'h403a7541, 32'hc2ad11af};
test_output[28384:28391] = '{32'h427e64bf, 32'h0, 32'h41e8c863, 32'h428ad6cd, 32'h0, 32'h0, 32'h403a7541, 32'h0};
test_input[28392:28399] = '{32'h42b64347, 32'hc1e509eb, 32'h42771785, 32'h42b97f46, 32'hc167a8db, 32'hc24bd46b, 32'hc176ec69, 32'hc24daa49};
test_output[28392:28399] = '{32'h42b64347, 32'h0, 32'h42771785, 32'h42b97f46, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28400:28407] = '{32'hc245489a, 32'hc08adc8c, 32'hc219c1ed, 32'h429dad13, 32'h425f6871, 32'h4293ee7d, 32'h4263544d, 32'hc2c7f5cc};
test_output[28400:28407] = '{32'h0, 32'h0, 32'h0, 32'h429dad13, 32'h425f6871, 32'h4293ee7d, 32'h4263544d, 32'h0};
test_input[28408:28415] = '{32'h4171db5e, 32'hc0b425f4, 32'hc236236f, 32'hc2b5c696, 32'hc0eed85a, 32'hc16fd3a4, 32'hc29f325f, 32'hc2a47013};
test_output[28408:28415] = '{32'h4171db5e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28416:28423] = '{32'hc2b7aae8, 32'h42a3fe89, 32'hc2a148e6, 32'hc2be0381, 32'hc28db08d, 32'h42beb994, 32'hc1a96347, 32'h42bd5fda};
test_output[28416:28423] = '{32'h0, 32'h42a3fe89, 32'h0, 32'h0, 32'h0, 32'h42beb994, 32'h0, 32'h42bd5fda};
test_input[28424:28431] = '{32'h42a42b8e, 32'h41e49e10, 32'hc2827f89, 32'hc164d897, 32'hc103680f, 32'h408d6ef8, 32'h42ada607, 32'h4298a74d};
test_output[28424:28431] = '{32'h42a42b8e, 32'h41e49e10, 32'h0, 32'h0, 32'h0, 32'h408d6ef8, 32'h42ada607, 32'h4298a74d};
test_input[28432:28439] = '{32'hc077cd01, 32'hc2a4dd66, 32'hc058d7ad, 32'hc2c59a21, 32'h42a9a140, 32'hc2b3500c, 32'hc2ab3a8b, 32'hc2af0dc9};
test_output[28432:28439] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a9a140, 32'h0, 32'h0, 32'h0};
test_input[28440:28447] = '{32'hc2900f4b, 32'hc2b64966, 32'hc292d95f, 32'hc258ed74, 32'h41a7abc1, 32'h420ce6bc, 32'hc259469f, 32'hc28b7bd7};
test_output[28440:28447] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41a7abc1, 32'h420ce6bc, 32'h0, 32'h0};
test_input[28448:28455] = '{32'h42738844, 32'hc2b18dfd, 32'hc27f1ea5, 32'h413fd3b8, 32'hc1c3d035, 32'hc23ff62b, 32'hc1d71f9d, 32'h4286c8db};
test_output[28448:28455] = '{32'h42738844, 32'h0, 32'h0, 32'h413fd3b8, 32'h0, 32'h0, 32'h0, 32'h4286c8db};
test_input[28456:28463] = '{32'hc1a03a63, 32'h428e6f44, 32'hc24fecd9, 32'hc09ae4f8, 32'h41f284e4, 32'hc28dcef7, 32'h42c269b3, 32'h42123d2f};
test_output[28456:28463] = '{32'h0, 32'h428e6f44, 32'h0, 32'h0, 32'h41f284e4, 32'h0, 32'h42c269b3, 32'h42123d2f};
test_input[28464:28471] = '{32'h42bea2a6, 32'h42858b20, 32'h425fe3eb, 32'hc161378c, 32'hc2861abe, 32'h412eec67, 32'h428c9b48, 32'h42c1ae77};
test_output[28464:28471] = '{32'h42bea2a6, 32'h42858b20, 32'h425fe3eb, 32'h0, 32'h0, 32'h412eec67, 32'h428c9b48, 32'h42c1ae77};
test_input[28472:28479] = '{32'h412c6bb6, 32'h4246599a, 32'h4245d975, 32'h42b8633f, 32'hc29c6def, 32'hc2ba7f27, 32'hc229bf0b, 32'hc2afb1e8};
test_output[28472:28479] = '{32'h412c6bb6, 32'h4246599a, 32'h4245d975, 32'h42b8633f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28480:28487] = '{32'hc25df8b0, 32'hc21fa7f1, 32'hc1cabd65, 32'h421e76dc, 32'h42b4baf9, 32'hc288fe17, 32'hc27a4a96, 32'h428b22d2};
test_output[28480:28487] = '{32'h0, 32'h0, 32'h0, 32'h421e76dc, 32'h42b4baf9, 32'h0, 32'h0, 32'h428b22d2};
test_input[28488:28495] = '{32'hc1b3bd6a, 32'hc2591095, 32'hc28125bb, 32'h406209cf, 32'hc28b1807, 32'hc2aab0a3, 32'hc29a4070, 32'hc18c4b70};
test_output[28488:28495] = '{32'h0, 32'h0, 32'h0, 32'h406209cf, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28496:28503] = '{32'h42899415, 32'h419d10ca, 32'hc23c736a, 32'hc27b8de0, 32'hc2aff01d, 32'h42376ef7, 32'hc1ce0703, 32'h4239ab16};
test_output[28496:28503] = '{32'h42899415, 32'h419d10ca, 32'h0, 32'h0, 32'h0, 32'h42376ef7, 32'h0, 32'h4239ab16};
test_input[28504:28511] = '{32'hc1de9fdf, 32'h41904495, 32'hc0b932f3, 32'h429ea1f2, 32'hc1efe7f9, 32'h42bdbe2d, 32'hc2930d60, 32'h4114b207};
test_output[28504:28511] = '{32'h0, 32'h41904495, 32'h0, 32'h429ea1f2, 32'h0, 32'h42bdbe2d, 32'h0, 32'h4114b207};
test_input[28512:28519] = '{32'hc2c1cd3c, 32'h427d0640, 32'h41981cbe, 32'hc2042d22, 32'hc2973982, 32'h425d51c6, 32'h40cb5caf, 32'h42afc177};
test_output[28512:28519] = '{32'h0, 32'h427d0640, 32'h41981cbe, 32'h0, 32'h0, 32'h425d51c6, 32'h40cb5caf, 32'h42afc177};
test_input[28520:28527] = '{32'h42bfd7dc, 32'h4189b4e0, 32'h41aded45, 32'hc2261bf0, 32'hc1946ef9, 32'h41cf108b, 32'h41dcd973, 32'h413b7e33};
test_output[28520:28527] = '{32'h42bfd7dc, 32'h4189b4e0, 32'h41aded45, 32'h0, 32'h0, 32'h41cf108b, 32'h41dcd973, 32'h413b7e33};
test_input[28528:28535] = '{32'hc23c88e1, 32'hc2c304b5, 32'hc28d69e6, 32'hc2a380b3, 32'hc212f937, 32'hc200a126, 32'hc2c0a896, 32'h40589307};
test_output[28528:28535] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40589307};
test_input[28536:28543] = '{32'h41f4960c, 32'h4287dac8, 32'h41be8f6e, 32'hc2adb96e, 32'h41a87338, 32'hc1f8bb28, 32'h404ccac3, 32'hc26432bd};
test_output[28536:28543] = '{32'h41f4960c, 32'h4287dac8, 32'h41be8f6e, 32'h0, 32'h41a87338, 32'h0, 32'h404ccac3, 32'h0};
test_input[28544:28551] = '{32'hc27fde3e, 32'hc2a5ec84, 32'h41af28e3, 32'hc2969db2, 32'hc2c190dc, 32'h41899627, 32'hc29615fa, 32'h424b6ec8};
test_output[28544:28551] = '{32'h0, 32'h0, 32'h41af28e3, 32'h0, 32'h0, 32'h41899627, 32'h0, 32'h424b6ec8};
test_input[28552:28559] = '{32'hc1d1cf8a, 32'hc1fe2e0f, 32'hc1c6acaa, 32'hc234814f, 32'hc221c7d0, 32'hc1c9491e, 32'h41f5c851, 32'hc299dc6e};
test_output[28552:28559] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f5c851, 32'h0};
test_input[28560:28567] = '{32'hc222631f, 32'hc06a1a26, 32'h41d788e5, 32'h40983c9e, 32'h40ef10f0, 32'h42a5f782, 32'hc1e92ab8, 32'h3fe54d52};
test_output[28560:28567] = '{32'h0, 32'h0, 32'h41d788e5, 32'h40983c9e, 32'h40ef10f0, 32'h42a5f782, 32'h0, 32'h3fe54d52};
test_input[28568:28575] = '{32'hc0098722, 32'h425683d5, 32'hc24a6e6e, 32'hc215e27b, 32'hc1f61d2c, 32'hbfe08982, 32'hc26a5e33, 32'h4284b3c0};
test_output[28568:28575] = '{32'h0, 32'h425683d5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4284b3c0};
test_input[28576:28583] = '{32'hc2a05003, 32'h42432f72, 32'hc21683a1, 32'hc2b8fcde, 32'hc1b82b7b, 32'h4102d745, 32'hc2b7c532, 32'hc298a0cf};
test_output[28576:28583] = '{32'h0, 32'h42432f72, 32'h0, 32'h0, 32'h0, 32'h4102d745, 32'h0, 32'h0};
test_input[28584:28591] = '{32'h42b416d5, 32'hbfec7551, 32'hc2085c1f, 32'h4028ee47, 32'h4211993d, 32'hc21e2429, 32'hc1723353, 32'hc2af748a};
test_output[28584:28591] = '{32'h42b416d5, 32'h0, 32'h0, 32'h4028ee47, 32'h4211993d, 32'h0, 32'h0, 32'h0};
test_input[28592:28599] = '{32'h42836817, 32'h426543fc, 32'h4283fe1b, 32'h4284c109, 32'hc2b06ac5, 32'h4196deb1, 32'hc2899261, 32'h40d21115};
test_output[28592:28599] = '{32'h42836817, 32'h426543fc, 32'h4283fe1b, 32'h4284c109, 32'h0, 32'h4196deb1, 32'h0, 32'h40d21115};
test_input[28600:28607] = '{32'hc2c6ce8d, 32'hc2a76c9a, 32'h4230d73a, 32'h42c151cd, 32'h42198206, 32'h42065657, 32'h41cb5a34, 32'hc2c32163};
test_output[28600:28607] = '{32'h0, 32'h0, 32'h4230d73a, 32'h42c151cd, 32'h42198206, 32'h42065657, 32'h41cb5a34, 32'h0};
test_input[28608:28615] = '{32'hc2790f49, 32'h42a7e287, 32'hc2424ab5, 32'h42908808, 32'hc233c7f4, 32'h4230b950, 32'hc1757656, 32'hc1d2aad6};
test_output[28608:28615] = '{32'h0, 32'h42a7e287, 32'h0, 32'h42908808, 32'h0, 32'h4230b950, 32'h0, 32'h0};
test_input[28616:28623] = '{32'hc28a2864, 32'h42a5d2bb, 32'h42c062db, 32'hc28347ae, 32'h4232934d, 32'h417532aa, 32'h42a03ff9, 32'h42bc92b7};
test_output[28616:28623] = '{32'h0, 32'h42a5d2bb, 32'h42c062db, 32'h0, 32'h4232934d, 32'h417532aa, 32'h42a03ff9, 32'h42bc92b7};
test_input[28624:28631] = '{32'hc22d90db, 32'hc216170e, 32'h42a204e9, 32'h4228b567, 32'h423b680f, 32'hc19f2d7e, 32'h4166dea2, 32'hc2a9dc24};
test_output[28624:28631] = '{32'h0, 32'h0, 32'h42a204e9, 32'h4228b567, 32'h423b680f, 32'h0, 32'h4166dea2, 32'h0};
test_input[28632:28639] = '{32'hc26b6a2a, 32'h418a8000, 32'hc27a6c46, 32'h427c3c30, 32'hc1b3c9e5, 32'h413ce1fd, 32'hc158ca06, 32'h4140a249};
test_output[28632:28639] = '{32'h0, 32'h418a8000, 32'h0, 32'h427c3c30, 32'h0, 32'h413ce1fd, 32'h0, 32'h4140a249};
test_input[28640:28647] = '{32'hc1cd6fe7, 32'hc254154a, 32'h40256eb3, 32'hc2b68521, 32'hc076fe0c, 32'hc26082f9, 32'hc104d4d9, 32'h42b9314c};
test_output[28640:28647] = '{32'h0, 32'h0, 32'h40256eb3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b9314c};
test_input[28648:28655] = '{32'h42201027, 32'h418b0abb, 32'h4219b5c6, 32'h41bf5291, 32'h415fe39d, 32'h4239983f, 32'hc280d5fd, 32'h429a81e1};
test_output[28648:28655] = '{32'h42201027, 32'h418b0abb, 32'h4219b5c6, 32'h41bf5291, 32'h415fe39d, 32'h4239983f, 32'h0, 32'h429a81e1};
test_input[28656:28663] = '{32'hc294470c, 32'h42af9c23, 32'h40a1526c, 32'h42192da5, 32'h42c55fad, 32'hc28dc5ca, 32'h42a04376, 32'hc2978b6d};
test_output[28656:28663] = '{32'h0, 32'h42af9c23, 32'h40a1526c, 32'h42192da5, 32'h42c55fad, 32'h0, 32'h42a04376, 32'h0};
test_input[28664:28671] = '{32'hc1c8c36c, 32'h4293e5c0, 32'h4232675b, 32'h419ff9c6, 32'h4218fb03, 32'h42be82ba, 32'h42607cec, 32'h41a1cb0d};
test_output[28664:28671] = '{32'h0, 32'h4293e5c0, 32'h4232675b, 32'h419ff9c6, 32'h4218fb03, 32'h42be82ba, 32'h42607cec, 32'h41a1cb0d};
test_input[28672:28679] = '{32'h421a65e2, 32'h42c47342, 32'h425ee023, 32'hc2c7571f, 32'h4281cd2f, 32'hc2855e8a, 32'h41229530, 32'hc2c582e8};
test_output[28672:28679] = '{32'h421a65e2, 32'h42c47342, 32'h425ee023, 32'h0, 32'h4281cd2f, 32'h0, 32'h41229530, 32'h0};
test_input[28680:28687] = '{32'hc2b97682, 32'h4000de52, 32'h4295feb9, 32'h42a66810, 32'hc08b559f, 32'hc2aa698c, 32'h4210595d, 32'h429b2610};
test_output[28680:28687] = '{32'h0, 32'h4000de52, 32'h4295feb9, 32'h42a66810, 32'h0, 32'h0, 32'h4210595d, 32'h429b2610};
test_input[28688:28695] = '{32'h42a907c1, 32'h42876b3a, 32'h4247bddd, 32'h41bd31d6, 32'hc28fa598, 32'hc29e059d, 32'hc27a6ea2, 32'hc2619113};
test_output[28688:28695] = '{32'h42a907c1, 32'h42876b3a, 32'h4247bddd, 32'h41bd31d6, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28696:28703] = '{32'hc058982f, 32'h413290ef, 32'h40698e19, 32'hc2a5ea59, 32'h4269166d, 32'h42c72a98, 32'h42989016, 32'h41f99855};
test_output[28696:28703] = '{32'h0, 32'h413290ef, 32'h40698e19, 32'h0, 32'h4269166d, 32'h42c72a98, 32'h42989016, 32'h41f99855};
test_input[28704:28711] = '{32'h42bdd167, 32'h426bfa7e, 32'hc2c546cd, 32'hc2afb152, 32'hc27b863f, 32'hc0341713, 32'hc27b7d6b, 32'h42af9c74};
test_output[28704:28711] = '{32'h42bdd167, 32'h426bfa7e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42af9c74};
test_input[28712:28719] = '{32'h424bf62b, 32'h42421433, 32'hc1b634fc, 32'hc218f6f3, 32'h423ab566, 32'hc260bb83, 32'hc28167e6, 32'h4134819a};
test_output[28712:28719] = '{32'h424bf62b, 32'h42421433, 32'h0, 32'h0, 32'h423ab566, 32'h0, 32'h0, 32'h4134819a};
test_input[28720:28727] = '{32'h42b4f157, 32'h41e40869, 32'h424fe1de, 32'hc209ae0a, 32'hc20ec3a3, 32'hc23c7d76, 32'h40a9e586, 32'hbf884af9};
test_output[28720:28727] = '{32'h42b4f157, 32'h41e40869, 32'h424fe1de, 32'h0, 32'h0, 32'h0, 32'h40a9e586, 32'h0};
test_input[28728:28735] = '{32'hc275eada, 32'hc2679944, 32'hc2c465c8, 32'h427523de, 32'h42579420, 32'h42395947, 32'hc29f9494, 32'h42842268};
test_output[28728:28735] = '{32'h0, 32'h0, 32'h0, 32'h427523de, 32'h42579420, 32'h42395947, 32'h0, 32'h42842268};
test_input[28736:28743] = '{32'h428d845d, 32'hc16f9577, 32'hc1d1df06, 32'h41574102, 32'hc1ebf713, 32'h416698a1, 32'hc2be3421, 32'h4197fa5e};
test_output[28736:28743] = '{32'h428d845d, 32'h0, 32'h0, 32'h41574102, 32'h0, 32'h416698a1, 32'h0, 32'h4197fa5e};
test_input[28744:28751] = '{32'hc2a4cb49, 32'hc2998f5a, 32'h424b652b, 32'h421e3c6e, 32'hc2805d3b, 32'hc11c6c3d, 32'h40bbbb9d, 32'hbfbb9622};
test_output[28744:28751] = '{32'h0, 32'h0, 32'h424b652b, 32'h421e3c6e, 32'h0, 32'h0, 32'h40bbbb9d, 32'h0};
test_input[28752:28759] = '{32'hc23560e8, 32'hc2ac2c23, 32'h42b9522f, 32'h41e0310c, 32'h4210f376, 32'hc2c13de6, 32'hc0c46dac, 32'h428e2ab3};
test_output[28752:28759] = '{32'h0, 32'h0, 32'h42b9522f, 32'h41e0310c, 32'h4210f376, 32'h0, 32'h0, 32'h428e2ab3};
test_input[28760:28767] = '{32'h42a0e88c, 32'h40eef283, 32'h425bc9ea, 32'hc25f39d2, 32'h424a542f, 32'h424372e3, 32'h420249e0, 32'hc0bcbd1f};
test_output[28760:28767] = '{32'h42a0e88c, 32'h40eef283, 32'h425bc9ea, 32'h0, 32'h424a542f, 32'h424372e3, 32'h420249e0, 32'h0};
test_input[28768:28775] = '{32'h4288c758, 32'hc2725d0e, 32'hc193ec0a, 32'h4292191d, 32'h4248dd52, 32'hc1b48292, 32'h422b1956, 32'hc24df5fc};
test_output[28768:28775] = '{32'h4288c758, 32'h0, 32'h0, 32'h4292191d, 32'h4248dd52, 32'h0, 32'h422b1956, 32'h0};
test_input[28776:28783] = '{32'hc2034939, 32'hc26cf25a, 32'hc2a83394, 32'hc2b72dc0, 32'hc19a3ad1, 32'h4020c5a5, 32'hc1fec710, 32'h428e174b};
test_output[28776:28783] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4020c5a5, 32'h0, 32'h428e174b};
test_input[28784:28791] = '{32'hc2421b96, 32'hc28128ef, 32'hc2a97921, 32'h41687a07, 32'hc291ddd2, 32'h419a75b1, 32'hc2b00c1c, 32'hc2182833};
test_output[28784:28791] = '{32'h0, 32'h0, 32'h0, 32'h41687a07, 32'h0, 32'h419a75b1, 32'h0, 32'h0};
test_input[28792:28799] = '{32'hc2a2671c, 32'h42680674, 32'h425327ed, 32'h41bb433e, 32'hbf85432d, 32'hc25b4cbe, 32'h429bd2d0, 32'h422580e1};
test_output[28792:28799] = '{32'h0, 32'h42680674, 32'h425327ed, 32'h41bb433e, 32'h0, 32'h0, 32'h429bd2d0, 32'h422580e1};
test_input[28800:28807] = '{32'hc2b9e741, 32'hc2c6fce0, 32'h429cd1b2, 32'hc21e682b, 32'hc2c3e5b8, 32'h40eed160, 32'hc18465cd, 32'hc2746ba4};
test_output[28800:28807] = '{32'h0, 32'h0, 32'h429cd1b2, 32'h0, 32'h0, 32'h40eed160, 32'h0, 32'h0};
test_input[28808:28815] = '{32'hc1f717d2, 32'hc2c5ee3a, 32'h42a2d231, 32'hc2a81f4b, 32'hc2af6253, 32'h41f529a0, 32'h419f3b41, 32'hc2a9d42f};
test_output[28808:28815] = '{32'h0, 32'h0, 32'h42a2d231, 32'h0, 32'h0, 32'h41f529a0, 32'h419f3b41, 32'h0};
test_input[28816:28823] = '{32'h4282806c, 32'hc297a614, 32'h42c1b07d, 32'hc1d486a9, 32'h412ce4a8, 32'hc273983c, 32'hc27d69f1, 32'hc1bd1d32};
test_output[28816:28823] = '{32'h4282806c, 32'h0, 32'h42c1b07d, 32'h0, 32'h412ce4a8, 32'h0, 32'h0, 32'h0};
test_input[28824:28831] = '{32'hc22c65c0, 32'hc282494e, 32'h41ca1317, 32'hc2424fae, 32'h423d5fdd, 32'hc12e79bc, 32'h42155dae, 32'h420b17ac};
test_output[28824:28831] = '{32'h0, 32'h0, 32'h41ca1317, 32'h0, 32'h423d5fdd, 32'h0, 32'h42155dae, 32'h420b17ac};
test_input[28832:28839] = '{32'hc0b9ee5b, 32'h3f7ec1ca, 32'hc0c5ac9f, 32'hc1c09378, 32'hc21b4273, 32'hc2b597af, 32'hc17b8ef0, 32'h4198191a};
test_output[28832:28839] = '{32'h0, 32'h3f7ec1ca, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4198191a};
test_input[28840:28847] = '{32'h42701d79, 32'h413c6734, 32'hc2a88732, 32'h420b22c4, 32'hc284817f, 32'hc28bb119, 32'h4155e90d, 32'h415ed470};
test_output[28840:28847] = '{32'h42701d79, 32'h413c6734, 32'h0, 32'h420b22c4, 32'h0, 32'h0, 32'h4155e90d, 32'h415ed470};
test_input[28848:28855] = '{32'h427998b4, 32'h42abd02c, 32'hc2120e5a, 32'h4250882a, 32'h42a2fc09, 32'hc2217080, 32'hc165bfe2, 32'hc29876b5};
test_output[28848:28855] = '{32'h427998b4, 32'h42abd02c, 32'h0, 32'h4250882a, 32'h42a2fc09, 32'h0, 32'h0, 32'h0};
test_input[28856:28863] = '{32'hc1d103dd, 32'h428fcc95, 32'h420414fe, 32'hc272a351, 32'h42b363f0, 32'h421ccaff, 32'h4274736a, 32'hc26dda0d};
test_output[28856:28863] = '{32'h0, 32'h428fcc95, 32'h420414fe, 32'h0, 32'h42b363f0, 32'h421ccaff, 32'h4274736a, 32'h0};
test_input[28864:28871] = '{32'hc16456fe, 32'h428b64f5, 32'h42b184d7, 32'h4236d9cc, 32'h42acb7ab, 32'h42b04b6b, 32'hc2980fab, 32'h41d4e2a6};
test_output[28864:28871] = '{32'h0, 32'h428b64f5, 32'h42b184d7, 32'h4236d9cc, 32'h42acb7ab, 32'h42b04b6b, 32'h0, 32'h41d4e2a6};
test_input[28872:28879] = '{32'h42c5d3c0, 32'hc27d72fd, 32'hc2b2d171, 32'h41f4bff1, 32'h4298def0, 32'h42be3781, 32'hc1c66abd, 32'hc1d7d979};
test_output[28872:28879] = '{32'h42c5d3c0, 32'h0, 32'h0, 32'h41f4bff1, 32'h4298def0, 32'h42be3781, 32'h0, 32'h0};
test_input[28880:28887] = '{32'h41d257d8, 32'h40ee88ae, 32'hc23d5c2c, 32'h4200bada, 32'hc24c4cea, 32'h42c20836, 32'h4207cf2f, 32'h425bd44a};
test_output[28880:28887] = '{32'h41d257d8, 32'h40ee88ae, 32'h0, 32'h4200bada, 32'h0, 32'h42c20836, 32'h4207cf2f, 32'h425bd44a};
test_input[28888:28895] = '{32'hc2b1835a, 32'h42b80a1d, 32'h410ffcee, 32'h41c95d3b, 32'h41e982e3, 32'h421c4170, 32'hc2c47f0c, 32'h42a14e7d};
test_output[28888:28895] = '{32'h0, 32'h42b80a1d, 32'h410ffcee, 32'h41c95d3b, 32'h41e982e3, 32'h421c4170, 32'h0, 32'h42a14e7d};
test_input[28896:28903] = '{32'hc2398d35, 32'hc1bb1c1f, 32'hc132d0f2, 32'hc2b2cbfc, 32'hc2b997e1, 32'hc23c6db3, 32'hc0a27636, 32'h42b33cce};
test_output[28896:28903] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b33cce};
test_input[28904:28911] = '{32'h4206a83f, 32'hc1562939, 32'h423a64a4, 32'h42bfe562, 32'h41c70a06, 32'hc0f82f81, 32'h412af1b5, 32'h427ddae4};
test_output[28904:28911] = '{32'h4206a83f, 32'h0, 32'h423a64a4, 32'h42bfe562, 32'h41c70a06, 32'h0, 32'h412af1b5, 32'h427ddae4};
test_input[28912:28919] = '{32'hc1d96d5f, 32'h4232b796, 32'hc1184ff5, 32'h427ddc8a, 32'hc20ad432, 32'hc2ab5138, 32'h40e89fd4, 32'h42c20be7};
test_output[28912:28919] = '{32'h0, 32'h4232b796, 32'h0, 32'h427ddc8a, 32'h0, 32'h0, 32'h40e89fd4, 32'h42c20be7};
test_input[28920:28927] = '{32'hc2a027f5, 32'h42620a32, 32'h40824907, 32'hc29e2e90, 32'h426e3f2c, 32'h42207539, 32'h42436474, 32'h429218ea};
test_output[28920:28927] = '{32'h0, 32'h42620a32, 32'h40824907, 32'h0, 32'h426e3f2c, 32'h42207539, 32'h42436474, 32'h429218ea};
test_input[28928:28935] = '{32'hc2722cab, 32'h428c1c87, 32'hc0bda893, 32'h41c450ee, 32'hc2b6b943, 32'h4246b629, 32'h42a3fa61, 32'hc2505811};
test_output[28928:28935] = '{32'h0, 32'h428c1c87, 32'h0, 32'h41c450ee, 32'h0, 32'h4246b629, 32'h42a3fa61, 32'h0};
test_input[28936:28943] = '{32'h427b27ea, 32'hc104eeff, 32'h424ad37b, 32'hc2c38b4d, 32'h42b76244, 32'hc2c0fbd1, 32'hc2bc9703, 32'h41e7dfac};
test_output[28936:28943] = '{32'h427b27ea, 32'h0, 32'h424ad37b, 32'h0, 32'h42b76244, 32'h0, 32'h0, 32'h41e7dfac};
test_input[28944:28951] = '{32'h3fa83dc6, 32'hc28ce835, 32'hc24f0fd6, 32'hc2b0fe6b, 32'hc1888981, 32'h40d5de87, 32'h41ae60e3, 32'h423c6725};
test_output[28944:28951] = '{32'h3fa83dc6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40d5de87, 32'h41ae60e3, 32'h423c6725};
test_input[28952:28959] = '{32'hc1645adf, 32'hc1c7bd90, 32'hc100d4da, 32'hc246948e, 32'h41c4cde9, 32'hc21287a3, 32'h41f74514, 32'hc14f49ac};
test_output[28952:28959] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41c4cde9, 32'h0, 32'h41f74514, 32'h0};
test_input[28960:28967] = '{32'hc2803532, 32'hc28c682e, 32'h42acd4c7, 32'h4299e3e9, 32'h41d80106, 32'h429181ae, 32'hc0133fb8, 32'hc229eacd};
test_output[28960:28967] = '{32'h0, 32'h0, 32'h42acd4c7, 32'h4299e3e9, 32'h41d80106, 32'h429181ae, 32'h0, 32'h0};
test_input[28968:28975] = '{32'hc1561103, 32'h40906c8e, 32'hc0879cd8, 32'hc2b8de30, 32'hc20ff95d, 32'hc1132cae, 32'hc2922e20, 32'h428744e0};
test_output[28968:28975] = '{32'h0, 32'h40906c8e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428744e0};
test_input[28976:28983] = '{32'hc2bd544a, 32'h42886fb6, 32'hc29ef31b, 32'h41e3d979, 32'hc249ab43, 32'hc26d5c90, 32'h42beb504, 32'h41ebb585};
test_output[28976:28983] = '{32'h0, 32'h42886fb6, 32'h0, 32'h41e3d979, 32'h0, 32'h0, 32'h42beb504, 32'h41ebb585};
test_input[28984:28991] = '{32'hc2b1216a, 32'h4191a9de, 32'h42a57af0, 32'hc2478bc4, 32'h42b878ee, 32'hc1710903, 32'hc29b32cb, 32'hc2c27015};
test_output[28984:28991] = '{32'h0, 32'h4191a9de, 32'h42a57af0, 32'h0, 32'h42b878ee, 32'h0, 32'h0, 32'h0};
test_input[28992:28999] = '{32'h4104648d, 32'hc2aaa654, 32'h4228ff4e, 32'hc1e88276, 32'h402604c2, 32'hc28e97df, 32'hc236a31c, 32'hc21e600c};
test_output[28992:28999] = '{32'h4104648d, 32'h0, 32'h4228ff4e, 32'h0, 32'h402604c2, 32'h0, 32'h0, 32'h0};
test_input[29000:29007] = '{32'hc2828c61, 32'hc26e79f7, 32'h421fc3d0, 32'h4015bf1a, 32'hc29bc1e8, 32'h42a038bb, 32'hc0578ee8, 32'hc1c96414};
test_output[29000:29007] = '{32'h0, 32'h0, 32'h421fc3d0, 32'h4015bf1a, 32'h0, 32'h42a038bb, 32'h0, 32'h0};
test_input[29008:29015] = '{32'hc210fc90, 32'h425129b0, 32'h41779133, 32'hc1ecd4ac, 32'hc2a44a5d, 32'hc004a378, 32'hc25bbadf, 32'hc2b63585};
test_output[29008:29015] = '{32'h0, 32'h425129b0, 32'h41779133, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29016:29023] = '{32'h42ae987c, 32'h416f507f, 32'h429da466, 32'h3f30861c, 32'hc29885ca, 32'hc2a56d13, 32'h42ab18a9, 32'hc2029c02};
test_output[29016:29023] = '{32'h42ae987c, 32'h416f507f, 32'h429da466, 32'h3f30861c, 32'h0, 32'h0, 32'h42ab18a9, 32'h0};
test_input[29024:29031] = '{32'hc20ca8e9, 32'h4298148a, 32'hc190e5b8, 32'hc20e49c9, 32'hc211a7ec, 32'hc2c12fdc, 32'hc195ed52, 32'hc0d31ed7};
test_output[29024:29031] = '{32'h0, 32'h4298148a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29032:29039] = '{32'hc26d0dce, 32'hc2b80377, 32'hc29ff9b2, 32'hc208c9d0, 32'h42945b46, 32'hc28a3f88, 32'h42708989, 32'hc2a4bde1};
test_output[29032:29039] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42945b46, 32'h0, 32'h42708989, 32'h0};
test_input[29040:29047] = '{32'h42006ebc, 32'h421de22b, 32'h428bc369, 32'hc2379e96, 32'hc2c3eed5, 32'h42c0ff50, 32'hc2b692d4, 32'hc2b97937};
test_output[29040:29047] = '{32'h42006ebc, 32'h421de22b, 32'h428bc369, 32'h0, 32'h0, 32'h42c0ff50, 32'h0, 32'h0};
test_input[29048:29055] = '{32'h412d712a, 32'hc1d5a6bd, 32'h41bc1b4c, 32'h42c2c4c5, 32'h41f18ac1, 32'hc2b1f31b, 32'hc28062e9, 32'hc28fc6a8};
test_output[29048:29055] = '{32'h412d712a, 32'h0, 32'h41bc1b4c, 32'h42c2c4c5, 32'h41f18ac1, 32'h0, 32'h0, 32'h0};
test_input[29056:29063] = '{32'h4288c7d7, 32'hc23bb747, 32'hc2552c2f, 32'h4267d505, 32'hc29d45e2, 32'hc29c534c, 32'hc22703f1, 32'h423a1fda};
test_output[29056:29063] = '{32'h4288c7d7, 32'h0, 32'h0, 32'h4267d505, 32'h0, 32'h0, 32'h0, 32'h423a1fda};
test_input[29064:29071] = '{32'hc1babe8c, 32'hc2b286a7, 32'hc2502f0f, 32'h42979ee6, 32'hc1f77c53, 32'h428e000d, 32'h429f9ba6, 32'hc2adbf68};
test_output[29064:29071] = '{32'h0, 32'h0, 32'h0, 32'h42979ee6, 32'h0, 32'h428e000d, 32'h429f9ba6, 32'h0};
test_input[29072:29079] = '{32'h42a4af08, 32'h42341381, 32'h415f1b69, 32'h42a796ef, 32'h410923d0, 32'hc29ac7dc, 32'h41c509e1, 32'hc2a843b0};
test_output[29072:29079] = '{32'h42a4af08, 32'h42341381, 32'h415f1b69, 32'h42a796ef, 32'h410923d0, 32'h0, 32'h41c509e1, 32'h0};
test_input[29080:29087] = '{32'hc29f733c, 32'h429d6666, 32'h4142b4bc, 32'h42223fc2, 32'h4096bbfb, 32'h42b9d4cf, 32'hc266ac63, 32'hc26df1c9};
test_output[29080:29087] = '{32'h0, 32'h429d6666, 32'h4142b4bc, 32'h42223fc2, 32'h4096bbfb, 32'h42b9d4cf, 32'h0, 32'h0};
test_input[29088:29095] = '{32'h42aa439f, 32'h41267340, 32'h42833619, 32'h3ee19bba, 32'hc23dc97c, 32'hc293e05d, 32'hc156d276, 32'h4225f30a};
test_output[29088:29095] = '{32'h42aa439f, 32'h41267340, 32'h42833619, 32'h3ee19bba, 32'h0, 32'h0, 32'h0, 32'h4225f30a};
test_input[29096:29103] = '{32'hc192486f, 32'h405683d5, 32'h40725b23, 32'hc2353cd1, 32'h41c2cd32, 32'h41dcb653, 32'h42661260, 32'hc1c0e12c};
test_output[29096:29103] = '{32'h0, 32'h405683d5, 32'h40725b23, 32'h0, 32'h41c2cd32, 32'h41dcb653, 32'h42661260, 32'h0};
test_input[29104:29111] = '{32'hc24cd606, 32'h429a60db, 32'hc1bfc40c, 32'hc1c380e9, 32'h4193c798, 32'hc2a8316f, 32'hc29a912b, 32'hc24e9f3c};
test_output[29104:29111] = '{32'h0, 32'h429a60db, 32'h0, 32'h0, 32'h4193c798, 32'h0, 32'h0, 32'h0};
test_input[29112:29119] = '{32'h4123f28f, 32'h4239b7b7, 32'hc21c3b2a, 32'h41966da7, 32'h42b8c670, 32'hc140cfb2, 32'h424fe3e7, 32'h424fa0cf};
test_output[29112:29119] = '{32'h4123f28f, 32'h4239b7b7, 32'h0, 32'h41966da7, 32'h42b8c670, 32'h0, 32'h424fe3e7, 32'h424fa0cf};
test_input[29120:29127] = '{32'h42a3d03f, 32'h427ef9d8, 32'hc286c5ff, 32'hc2b46264, 32'h419afab6, 32'hc294b64c, 32'hc2c167a1, 32'hc2161d46};
test_output[29120:29127] = '{32'h42a3d03f, 32'h427ef9d8, 32'h0, 32'h0, 32'h419afab6, 32'h0, 32'h0, 32'h0};
test_input[29128:29135] = '{32'h421a3af6, 32'h42be6ad6, 32'h4273ac0d, 32'hc272ea00, 32'hc18bd221, 32'hc29083f9, 32'hc1fceef9, 32'hc2bf317e};
test_output[29128:29135] = '{32'h421a3af6, 32'h42be6ad6, 32'h4273ac0d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29136:29143] = '{32'hc20b7a5d, 32'h42bd10cc, 32'h4260e271, 32'h4263a3d9, 32'hc25d2a4a, 32'hc1adb839, 32'hc27ccb87, 32'h41f70a01};
test_output[29136:29143] = '{32'h0, 32'h42bd10cc, 32'h4260e271, 32'h4263a3d9, 32'h0, 32'h0, 32'h0, 32'h41f70a01};
test_input[29144:29151] = '{32'h42b8c230, 32'h41862d36, 32'h42a8e544, 32'hc27fa5c0, 32'hc19e224e, 32'hc230143b, 32'h429d2b09, 32'hc2b6a2ae};
test_output[29144:29151] = '{32'h42b8c230, 32'h41862d36, 32'h42a8e544, 32'h0, 32'h0, 32'h0, 32'h429d2b09, 32'h0};
test_input[29152:29159] = '{32'hc238e541, 32'hc22a79d1, 32'h4244e070, 32'h429d0a20, 32'h42987153, 32'hc08f9253, 32'h4180af27, 32'h41868a0a};
test_output[29152:29159] = '{32'h0, 32'h0, 32'h4244e070, 32'h429d0a20, 32'h42987153, 32'h0, 32'h4180af27, 32'h41868a0a};
test_input[29160:29167] = '{32'h428ad606, 32'hc12a483c, 32'hc120e4b4, 32'hc2c19bb7, 32'hc195c00c, 32'hc26facde, 32'h42c1dbff, 32'h42c7b526};
test_output[29160:29167] = '{32'h428ad606, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c1dbff, 32'h42c7b526};
test_input[29168:29175] = '{32'hc277bb85, 32'hc1298a83, 32'h429a036c, 32'h41e03acd, 32'hbff731f5, 32'hc251f1be, 32'h4254ffcf, 32'hc1d842e1};
test_output[29168:29175] = '{32'h0, 32'h0, 32'h429a036c, 32'h41e03acd, 32'h0, 32'h0, 32'h4254ffcf, 32'h0};
test_input[29176:29183] = '{32'h428d369c, 32'hc2777d25, 32'h423fe963, 32'hc27e65e7, 32'hc0b5efb5, 32'hc20970de, 32'hc29812d9, 32'h42c7f5e1};
test_output[29176:29183] = '{32'h428d369c, 32'h0, 32'h423fe963, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c7f5e1};
test_input[29184:29191] = '{32'h4277a260, 32'h427e7138, 32'hc29b66be, 32'h41cc13dd, 32'h429a718a, 32'hc2a09a0f, 32'h40f4b364, 32'hc27c3fa1};
test_output[29184:29191] = '{32'h4277a260, 32'h427e7138, 32'h0, 32'h41cc13dd, 32'h429a718a, 32'h0, 32'h40f4b364, 32'h0};
test_input[29192:29199] = '{32'h425d87d5, 32'h4149cc97, 32'h404738ef, 32'h42847465, 32'h4291f8ab, 32'h4277ab6c, 32'h429b05ca, 32'h42bb6146};
test_output[29192:29199] = '{32'h425d87d5, 32'h4149cc97, 32'h404738ef, 32'h42847465, 32'h4291f8ab, 32'h4277ab6c, 32'h429b05ca, 32'h42bb6146};
test_input[29200:29207] = '{32'h42a3d973, 32'h426499ed, 32'h42997ea2, 32'h42895e60, 32'h42880fc1, 32'h42c65253, 32'hc232fea3, 32'h42b75fc7};
test_output[29200:29207] = '{32'h42a3d973, 32'h426499ed, 32'h42997ea2, 32'h42895e60, 32'h42880fc1, 32'h42c65253, 32'h0, 32'h42b75fc7};
test_input[29208:29215] = '{32'hc1944a9e, 32'h4291b504, 32'hc0c15c7c, 32'h42293c71, 32'h41adee13, 32'hc28a3cf1, 32'hc26b5a1a, 32'hc257cbf6};
test_output[29208:29215] = '{32'h0, 32'h4291b504, 32'h0, 32'h42293c71, 32'h41adee13, 32'h0, 32'h0, 32'h0};
test_input[29216:29223] = '{32'hc1c6f934, 32'hc26e635b, 32'hc25b3748, 32'h429a25d5, 32'h4232e518, 32'h426a9f59, 32'h41e88825, 32'h420bffd9};
test_output[29216:29223] = '{32'h0, 32'h0, 32'h0, 32'h429a25d5, 32'h4232e518, 32'h426a9f59, 32'h41e88825, 32'h420bffd9};
test_input[29224:29231] = '{32'hc25e83c4, 32'hc2361d6e, 32'h42c4b2d9, 32'h41dd0704, 32'h42866522, 32'hc2179c66, 32'h420534c9, 32'h40e7e4c9};
test_output[29224:29231] = '{32'h0, 32'h0, 32'h42c4b2d9, 32'h41dd0704, 32'h42866522, 32'h0, 32'h420534c9, 32'h40e7e4c9};
test_input[29232:29239] = '{32'hc237c526, 32'h4213ee91, 32'h42bc926e, 32'hc2b6fd0b, 32'h4292c668, 32'hc17b3655, 32'h4208b080, 32'hc02b4cfb};
test_output[29232:29239] = '{32'h0, 32'h4213ee91, 32'h42bc926e, 32'h0, 32'h4292c668, 32'h0, 32'h4208b080, 32'h0};
test_input[29240:29247] = '{32'hc263e639, 32'h423afedc, 32'h42ae8c58, 32'hc1ce2398, 32'hc2bb577c, 32'h41d2a259, 32'hc2a6cdbd, 32'h414bec93};
test_output[29240:29247] = '{32'h0, 32'h423afedc, 32'h42ae8c58, 32'h0, 32'h0, 32'h41d2a259, 32'h0, 32'h414bec93};
test_input[29248:29255] = '{32'hc28bf8fe, 32'h42895f65, 32'hc28a4190, 32'hc1d4ce63, 32'h41d589ec, 32'hc1286d69, 32'h42a391ea, 32'hc27b83db};
test_output[29248:29255] = '{32'h0, 32'h42895f65, 32'h0, 32'h0, 32'h41d589ec, 32'h0, 32'h42a391ea, 32'h0};
test_input[29256:29263] = '{32'h4186fbda, 32'hc1c27d9e, 32'hc28287a2, 32'h4253f868, 32'h42ae9075, 32'h41a11ad2, 32'hc1329918, 32'h427395b5};
test_output[29256:29263] = '{32'h4186fbda, 32'h0, 32'h0, 32'h4253f868, 32'h42ae9075, 32'h41a11ad2, 32'h0, 32'h427395b5};
test_input[29264:29271] = '{32'hc24b0e38, 32'hc2ac04cc, 32'h3f93eab0, 32'hc1acc9ef, 32'hc28fc1ff, 32'h41efa295, 32'hc2a6f694, 32'h4273ab74};
test_output[29264:29271] = '{32'h0, 32'h0, 32'h3f93eab0, 32'h0, 32'h0, 32'h41efa295, 32'h0, 32'h4273ab74};
test_input[29272:29279] = '{32'hc243d8b2, 32'h41f98abd, 32'h415a7920, 32'hc2804c55, 32'h426e69d9, 32'h4146c0a0, 32'h42b51d6e, 32'h41134577};
test_output[29272:29279] = '{32'h0, 32'h41f98abd, 32'h415a7920, 32'h0, 32'h426e69d9, 32'h4146c0a0, 32'h42b51d6e, 32'h41134577};
test_input[29280:29287] = '{32'hc1cd34cf, 32'h42b86dfa, 32'h422cb87b, 32'h42a6b004, 32'hc1adc7b9, 32'h42771773, 32'h403373a0, 32'hc29ca4a2};
test_output[29280:29287] = '{32'h0, 32'h42b86dfa, 32'h422cb87b, 32'h42a6b004, 32'h0, 32'h42771773, 32'h403373a0, 32'h0};
test_input[29288:29295] = '{32'hc2373147, 32'hc2b0da52, 32'hc1639868, 32'h42ad030a, 32'h42b97a5f, 32'hc22657fe, 32'h405b9884, 32'hc1eff293};
test_output[29288:29295] = '{32'h0, 32'h0, 32'h0, 32'h42ad030a, 32'h42b97a5f, 32'h0, 32'h405b9884, 32'h0};
test_input[29296:29303] = '{32'h42aaa6de, 32'h41edc65f, 32'h420e8333, 32'hc2a35926, 32'h4071245d, 32'h42b728c7, 32'h42b62b45, 32'h429e9ad6};
test_output[29296:29303] = '{32'h42aaa6de, 32'h41edc65f, 32'h420e8333, 32'h0, 32'h4071245d, 32'h42b728c7, 32'h42b62b45, 32'h429e9ad6};
test_input[29304:29311] = '{32'h42811a51, 32'h4251b835, 32'hc22eea9d, 32'h42630329, 32'h4281a089, 32'h42a10d14, 32'h41b2ecb1, 32'hc1a0881b};
test_output[29304:29311] = '{32'h42811a51, 32'h4251b835, 32'h0, 32'h42630329, 32'h4281a089, 32'h42a10d14, 32'h41b2ecb1, 32'h0};
test_input[29312:29319] = '{32'hc2a71bbc, 32'hc2ab8fc0, 32'hbfe97678, 32'hc2b82042, 32'hc2ba8d90, 32'h42911a1b, 32'h42c1f0e9, 32'hc27be177};
test_output[29312:29319] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42911a1b, 32'h42c1f0e9, 32'h0};
test_input[29320:29327] = '{32'h42386968, 32'h42084069, 32'h4210a5f5, 32'h41e6c190, 32'h4278824d, 32'hc2727eab, 32'h421db548, 32'h420c35a7};
test_output[29320:29327] = '{32'h42386968, 32'h42084069, 32'h4210a5f5, 32'h41e6c190, 32'h4278824d, 32'h0, 32'h421db548, 32'h420c35a7};
test_input[29328:29335] = '{32'h427d7145, 32'hc272c81a, 32'h42c0e7ce, 32'hc263646a, 32'hc180a47b, 32'hc2a9760d, 32'h42c1752b, 32'h4262e5d8};
test_output[29328:29335] = '{32'h427d7145, 32'h0, 32'h42c0e7ce, 32'h0, 32'h0, 32'h0, 32'h42c1752b, 32'h4262e5d8};
test_input[29336:29343] = '{32'h4190063a, 32'hc200a53a, 32'hc1e8bb6b, 32'h427db9a9, 32'hc215990e, 32'hc243952b, 32'h4115b38b, 32'hc2689dda};
test_output[29336:29343] = '{32'h4190063a, 32'h0, 32'h0, 32'h427db9a9, 32'h0, 32'h0, 32'h4115b38b, 32'h0};
test_input[29344:29351] = '{32'hc29c73b6, 32'h41f4063e, 32'hc1ab1fc2, 32'hc175861c, 32'hc2957b9b, 32'h42949a77, 32'hc2699581, 32'hc157f307};
test_output[29344:29351] = '{32'h0, 32'h41f4063e, 32'h0, 32'h0, 32'h0, 32'h42949a77, 32'h0, 32'h0};
test_input[29352:29359] = '{32'h413b4489, 32'hc1fb9c71, 32'hc26726c6, 32'h4294520f, 32'h42768fb4, 32'h42889cd0, 32'hc1ed90e4, 32'hc2aa2cda};
test_output[29352:29359] = '{32'h413b4489, 32'h0, 32'h0, 32'h4294520f, 32'h42768fb4, 32'h42889cd0, 32'h0, 32'h0};
test_input[29360:29367] = '{32'hc243bb86, 32'h42111fe9, 32'h426c47cc, 32'hc259ca53, 32'hc27706d9, 32'h4225f3a0, 32'hc2619928, 32'h429d0bae};
test_output[29360:29367] = '{32'h0, 32'h42111fe9, 32'h426c47cc, 32'h0, 32'h0, 32'h4225f3a0, 32'h0, 32'h429d0bae};
test_input[29368:29375] = '{32'h416052b8, 32'h42bc35da, 32'hc23184d6, 32'hc29022c1, 32'h42846ee6, 32'hc1e90411, 32'h414af7eb, 32'hc28a815a};
test_output[29368:29375] = '{32'h416052b8, 32'h42bc35da, 32'h0, 32'h0, 32'h42846ee6, 32'h0, 32'h414af7eb, 32'h0};
test_input[29376:29383] = '{32'hc1dc9643, 32'hc2c02e94, 32'h413daa98, 32'hc27b3f4f, 32'hc27844f6, 32'hc28b29ed, 32'h418f1e4c, 32'h422ab850};
test_output[29376:29383] = '{32'h0, 32'h0, 32'h413daa98, 32'h0, 32'h0, 32'h0, 32'h418f1e4c, 32'h422ab850};
test_input[29384:29391] = '{32'hc1f82ff6, 32'h427b1e87, 32'hc1905a69, 32'h42c7bafa, 32'hc2624368, 32'hc24d0bac, 32'hc233277e, 32'hc1bf8515};
test_output[29384:29391] = '{32'h0, 32'h427b1e87, 32'h0, 32'h42c7bafa, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29392:29399] = '{32'h3e39357e, 32'h4291579f, 32'h4219f437, 32'hc2110f35, 32'hc2153974, 32'h424776bc, 32'hc21e1b36, 32'h429b7238};
test_output[29392:29399] = '{32'h3e39357e, 32'h4291579f, 32'h4219f437, 32'h0, 32'h0, 32'h424776bc, 32'h0, 32'h429b7238};
test_input[29400:29407] = '{32'hc2900522, 32'hc0c64c04, 32'hc27b1898, 32'h402ff1da, 32'hc1814b22, 32'h423fdf38, 32'hc211a786, 32'hc27f8c1d};
test_output[29400:29407] = '{32'h0, 32'h0, 32'h0, 32'h402ff1da, 32'h0, 32'h423fdf38, 32'h0, 32'h0};
test_input[29408:29415] = '{32'h412c58b3, 32'h41cdf419, 32'h41813978, 32'h41e87055, 32'hc2b4ec6a, 32'hc257f5bf, 32'hc2c5c171, 32'hc153f283};
test_output[29408:29415] = '{32'h412c58b3, 32'h41cdf419, 32'h41813978, 32'h41e87055, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29416:29423] = '{32'hc248e514, 32'h42bcb013, 32'h4209f7ed, 32'hc2a73eb4, 32'h4214dd14, 32'hc175da0e, 32'h41e7c598, 32'h41b487df};
test_output[29416:29423] = '{32'h0, 32'h42bcb013, 32'h4209f7ed, 32'h0, 32'h4214dd14, 32'h0, 32'h41e7c598, 32'h41b487df};
test_input[29424:29431] = '{32'h42c0fab0, 32'h427eb919, 32'h4241bb89, 32'hc20f5a75, 32'hc22e060a, 32'hc1b9cec2, 32'hc26d86ab, 32'hc1fa5351};
test_output[29424:29431] = '{32'h42c0fab0, 32'h427eb919, 32'h4241bb89, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29432:29439] = '{32'hc11334c1, 32'hc1884e72, 32'hc25d799f, 32'h42a27be1, 32'h41ae1f36, 32'h425f661b, 32'hc144903e, 32'hc0e40ac2};
test_output[29432:29439] = '{32'h0, 32'h0, 32'h0, 32'h42a27be1, 32'h41ae1f36, 32'h425f661b, 32'h0, 32'h0};
test_input[29440:29447] = '{32'hbf209750, 32'hc2c4c14d, 32'hc29205e8, 32'h4198e1da, 32'hc1e48072, 32'hc2c0d2bc, 32'h4237c83a, 32'hc24c13dc};
test_output[29440:29447] = '{32'h0, 32'h0, 32'h0, 32'h4198e1da, 32'h0, 32'h0, 32'h4237c83a, 32'h0};
test_input[29448:29455] = '{32'h41ea483d, 32'h429bb80d, 32'h3f95e763, 32'h41bce30d, 32'hc1b36940, 32'h429373ac, 32'h42bf8641, 32'h4272fbf1};
test_output[29448:29455] = '{32'h41ea483d, 32'h429bb80d, 32'h3f95e763, 32'h41bce30d, 32'h0, 32'h429373ac, 32'h42bf8641, 32'h4272fbf1};
test_input[29456:29463] = '{32'hc105ec09, 32'hc14ec211, 32'hc2273e5f, 32'hc28332b3, 32'h418f040c, 32'h415b395b, 32'hc212fa37, 32'hc1821bd2};
test_output[29456:29463] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h418f040c, 32'h415b395b, 32'h0, 32'h0};
test_input[29464:29471] = '{32'hc1d92e99, 32'h426b119a, 32'hc2a110e1, 32'hc2b2c23d, 32'h4252c24c, 32'h40a95900, 32'h42072b3a, 32'hc2b54f90};
test_output[29464:29471] = '{32'h0, 32'h426b119a, 32'h0, 32'h0, 32'h4252c24c, 32'h40a95900, 32'h42072b3a, 32'h0};
test_input[29472:29479] = '{32'hc19007d6, 32'hc280addd, 32'hc19fc1e3, 32'h42b7fafd, 32'h424de4c6, 32'h42c4ba35, 32'hc28c30b2, 32'hc26c440f};
test_output[29472:29479] = '{32'h0, 32'h0, 32'h0, 32'h42b7fafd, 32'h424de4c6, 32'h42c4ba35, 32'h0, 32'h0};
test_input[29480:29487] = '{32'h428cfe71, 32'h42bba32f, 32'hc285399d, 32'hc0b9c94a, 32'hc20dd952, 32'h428afaff, 32'hc27fa71a, 32'h428ce69e};
test_output[29480:29487] = '{32'h428cfe71, 32'h42bba32f, 32'h0, 32'h0, 32'h0, 32'h428afaff, 32'h0, 32'h428ce69e};
test_input[29488:29495] = '{32'hc2c3c92c, 32'hc2a1cb4b, 32'hc2b40fa3, 32'hc1d0fabc, 32'hc269aa46, 32'h41dc31fa, 32'hc0b25315, 32'h4123b333};
test_output[29488:29495] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41dc31fa, 32'h0, 32'h4123b333};
test_input[29496:29503] = '{32'h4159c91b, 32'h421f0b7b, 32'h41f2f39d, 32'hc1aac78f, 32'h412343dd, 32'h417244d6, 32'h422a3906, 32'h425e5e37};
test_output[29496:29503] = '{32'h4159c91b, 32'h421f0b7b, 32'h41f2f39d, 32'h0, 32'h412343dd, 32'h417244d6, 32'h422a3906, 32'h425e5e37};
test_input[29504:29511] = '{32'hc2aabf62, 32'hc2a97551, 32'hc1828a6e, 32'hc237f752, 32'h42814ac2, 32'h42c3bf14, 32'hc14a9dac, 32'hbff92623};
test_output[29504:29511] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42814ac2, 32'h42c3bf14, 32'h0, 32'h0};
test_input[29512:29519] = '{32'hc23878f3, 32'h427581d3, 32'h42ab305d, 32'hc229beff, 32'h42010d1a, 32'h42ac7d9f, 32'h428a58d1, 32'h3ef82935};
test_output[29512:29519] = '{32'h0, 32'h427581d3, 32'h42ab305d, 32'h0, 32'h42010d1a, 32'h42ac7d9f, 32'h428a58d1, 32'h3ef82935};
test_input[29520:29527] = '{32'h429d7b00, 32'hc23928c5, 32'hc1506de7, 32'h4278d071, 32'hc2980394, 32'hc23b9f51, 32'hc1d95e6b, 32'h421f7ca6};
test_output[29520:29527] = '{32'h429d7b00, 32'h0, 32'h0, 32'h4278d071, 32'h0, 32'h0, 32'h0, 32'h421f7ca6};
test_input[29528:29535] = '{32'h428058f8, 32'h421eaf7e, 32'hc24c4b66, 32'hc188bedf, 32'h42059073, 32'hc29a3ecb, 32'h42afaf3b, 32'hc2625caa};
test_output[29528:29535] = '{32'h428058f8, 32'h421eaf7e, 32'h0, 32'h0, 32'h42059073, 32'h0, 32'h42afaf3b, 32'h0};
test_input[29536:29543] = '{32'hc29c24a6, 32'h4104b916, 32'hc29662af, 32'h42ac42e1, 32'hc19e0f87, 32'hc2450c85, 32'hc2b33056, 32'hc285472e};
test_output[29536:29543] = '{32'h0, 32'h4104b916, 32'h0, 32'h42ac42e1, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29544:29551] = '{32'hc26e1dfe, 32'hc1d73b11, 32'h413a6dc4, 32'h426f31c1, 32'hc208c304, 32'hc27330d8, 32'hc1e928d3, 32'h428933ff};
test_output[29544:29551] = '{32'h0, 32'h0, 32'h413a6dc4, 32'h426f31c1, 32'h0, 32'h0, 32'h0, 32'h428933ff};
test_input[29552:29559] = '{32'hc1b39788, 32'h42abd27c, 32'h428bfc30, 32'hc2b9eac6, 32'hc2b14333, 32'hc2409aca, 32'hc2c59067, 32'hc2744d76};
test_output[29552:29559] = '{32'h0, 32'h42abd27c, 32'h428bfc30, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29560:29567] = '{32'hc284917a, 32'h429e6a22, 32'h4295ed3c, 32'h428e106f, 32'hc2c35346, 32'hc260f4b2, 32'h42556698, 32'h428c62fe};
test_output[29560:29567] = '{32'h0, 32'h429e6a22, 32'h4295ed3c, 32'h428e106f, 32'h0, 32'h0, 32'h42556698, 32'h428c62fe};
test_input[29568:29575] = '{32'h42509377, 32'h40c7d1c8, 32'h427f5610, 32'hc1c2adaa, 32'h4242dff4, 32'h42780d95, 32'h41e715a1, 32'h4241a4c7};
test_output[29568:29575] = '{32'h42509377, 32'h40c7d1c8, 32'h427f5610, 32'h0, 32'h4242dff4, 32'h42780d95, 32'h41e715a1, 32'h4241a4c7};
test_input[29576:29583] = '{32'hc2be7d57, 32'hc29453a8, 32'h41cb5b5d, 32'h42a76113, 32'hc16d5d99, 32'h42b7c523, 32'h42b0cc7a, 32'h42c55fe8};
test_output[29576:29583] = '{32'h0, 32'h0, 32'h41cb5b5d, 32'h42a76113, 32'h0, 32'h42b7c523, 32'h42b0cc7a, 32'h42c55fe8};
test_input[29584:29591] = '{32'h426b2d4c, 32'hc1f75c03, 32'hc2b67c32, 32'h4297cbd8, 32'h417a6a07, 32'hc2908ba0, 32'hc233bace, 32'h416dd4c6};
test_output[29584:29591] = '{32'h426b2d4c, 32'h0, 32'h0, 32'h4297cbd8, 32'h417a6a07, 32'h0, 32'h0, 32'h416dd4c6};
test_input[29592:29599] = '{32'hc23684da, 32'h420fca65, 32'hc1f41e26, 32'h42bffffa, 32'hc245a9bc, 32'hc2b8dc33, 32'hc26ab5e8, 32'h414cf25d};
test_output[29592:29599] = '{32'h0, 32'h420fca65, 32'h0, 32'h42bffffa, 32'h0, 32'h0, 32'h0, 32'h414cf25d};
test_input[29600:29607] = '{32'h420a232b, 32'hc2b26ed2, 32'hc214b05b, 32'h42bae98d, 32'h42b53dc9, 32'h4288f7c3, 32'hc25c2c2d, 32'hc1d27179};
test_output[29600:29607] = '{32'h420a232b, 32'h0, 32'h0, 32'h42bae98d, 32'h42b53dc9, 32'h4288f7c3, 32'h0, 32'h0};
test_input[29608:29615] = '{32'hc23f36d8, 32'h4266fafc, 32'hc25bab16, 32'h4273a85f, 32'hc22d8d23, 32'h42bc8ef6, 32'hc19851ca, 32'h41e89a30};
test_output[29608:29615] = '{32'h0, 32'h4266fafc, 32'h0, 32'h4273a85f, 32'h0, 32'h42bc8ef6, 32'h0, 32'h41e89a30};
test_input[29616:29623] = '{32'hc1e98ad2, 32'hc2a7fbf1, 32'hc2996ba6, 32'hc29f2324, 32'h4086d94b, 32'hc13e5412, 32'h42b5fb65, 32'hc1c54d8e};
test_output[29616:29623] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4086d94b, 32'h0, 32'h42b5fb65, 32'h0};
test_input[29624:29631] = '{32'hc24b5d3c, 32'h426e7cea, 32'hc2a1abd0, 32'h4292b2b9, 32'h4130ef51, 32'h42012515, 32'h41a2fb72, 32'h42b8f9ba};
test_output[29624:29631] = '{32'h0, 32'h426e7cea, 32'h0, 32'h4292b2b9, 32'h4130ef51, 32'h42012515, 32'h41a2fb72, 32'h42b8f9ba};
test_input[29632:29639] = '{32'hc1e9887d, 32'hc15f8605, 32'h421521e7, 32'h42bc241b, 32'h4284e252, 32'hc1ab23fd, 32'h427b8a03, 32'hc2a99fc2};
test_output[29632:29639] = '{32'h0, 32'h0, 32'h421521e7, 32'h42bc241b, 32'h4284e252, 32'h0, 32'h427b8a03, 32'h0};
test_input[29640:29647] = '{32'hc29ef299, 32'h40a1f148, 32'h42a53c0d, 32'h42c058d6, 32'h422e1794, 32'hc16c507a, 32'h4238d20e, 32'h420a15bb};
test_output[29640:29647] = '{32'h0, 32'h40a1f148, 32'h42a53c0d, 32'h42c058d6, 32'h422e1794, 32'h0, 32'h4238d20e, 32'h420a15bb};
test_input[29648:29655] = '{32'h41e18ab8, 32'hc268bfea, 32'hc041980b, 32'hc215a323, 32'hc2a50537, 32'hc253eab8, 32'hc29a16ed, 32'h42a2af29};
test_output[29648:29655] = '{32'h41e18ab8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a2af29};
test_input[29656:29663] = '{32'hc28c87a4, 32'hc2a45484, 32'h41d8286e, 32'hc27ea825, 32'h4294db1f, 32'h42b9a657, 32'hc20a59bb, 32'h42b10d02};
test_output[29656:29663] = '{32'h0, 32'h0, 32'h41d8286e, 32'h0, 32'h4294db1f, 32'h42b9a657, 32'h0, 32'h42b10d02};
test_input[29664:29671] = '{32'h425f2a38, 32'h41dd336b, 32'hc2b86a30, 32'h4223ae9d, 32'h41465939, 32'h41e38218, 32'hc2aeea8e, 32'hc1724e75};
test_output[29664:29671] = '{32'h425f2a38, 32'h41dd336b, 32'h0, 32'h4223ae9d, 32'h41465939, 32'h41e38218, 32'h0, 32'h0};
test_input[29672:29679] = '{32'hc27b131b, 32'h3eb03b44, 32'hc15417a8, 32'hc0cabc9f, 32'hc271c60f, 32'hc2b60cb4, 32'hc192d2c4, 32'h427b5917};
test_output[29672:29679] = '{32'h0, 32'h3eb03b44, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427b5917};
test_input[29680:29687] = '{32'hc1d61b10, 32'h42a1451b, 32'hc2981202, 32'hc1c9c38a, 32'hc207ec45, 32'h4212d84d, 32'h42c46bf1, 32'h42aaf4f5};
test_output[29680:29687] = '{32'h0, 32'h42a1451b, 32'h0, 32'h0, 32'h0, 32'h4212d84d, 32'h42c46bf1, 32'h42aaf4f5};
test_input[29688:29695] = '{32'hc2b354f8, 32'hc2c11df0, 32'h427675ad, 32'h425a3c90, 32'h42b5e8f0, 32'hc280bc05, 32'hc1108c72, 32'hc2a849f1};
test_output[29688:29695] = '{32'h0, 32'h0, 32'h427675ad, 32'h425a3c90, 32'h42b5e8f0, 32'h0, 32'h0, 32'h0};
test_input[29696:29703] = '{32'hc24b1598, 32'hc2b974f6, 32'h42a54697, 32'hc2633e9a, 32'h41b57ae7, 32'h42737ff2, 32'hc2c0a49e, 32'h42c05424};
test_output[29696:29703] = '{32'h0, 32'h0, 32'h42a54697, 32'h0, 32'h41b57ae7, 32'h42737ff2, 32'h0, 32'h42c05424};
test_input[29704:29711] = '{32'h42353ae1, 32'h3e0ba43d, 32'hc0a44dce, 32'hc255d3ec, 32'h423301be, 32'hc2c0716c, 32'h4241c695, 32'hc2c66e27};
test_output[29704:29711] = '{32'h42353ae1, 32'h3e0ba43d, 32'h0, 32'h0, 32'h423301be, 32'h0, 32'h4241c695, 32'h0};
test_input[29712:29719] = '{32'hc2792143, 32'h404e4b0e, 32'hc2b140ce, 32'hc266355b, 32'h425a5895, 32'hc29307af, 32'h42bb93d2, 32'h42a2544d};
test_output[29712:29719] = '{32'h0, 32'h404e4b0e, 32'h0, 32'h0, 32'h425a5895, 32'h0, 32'h42bb93d2, 32'h42a2544d};
test_input[29720:29727] = '{32'h42763a27, 32'h421a760f, 32'hc2b86ef6, 32'h42afa794, 32'h42b9ba5f, 32'hc1467fb3, 32'h41bde495, 32'h4284def3};
test_output[29720:29727] = '{32'h42763a27, 32'h421a760f, 32'h0, 32'h42afa794, 32'h42b9ba5f, 32'h0, 32'h41bde495, 32'h4284def3};
test_input[29728:29735] = '{32'h4263c2dd, 32'hc25ce1f7, 32'hbfa1b1f3, 32'h42456fee, 32'h422ebdf4, 32'h42652820, 32'h4283036d, 32'h4299e6d9};
test_output[29728:29735] = '{32'h4263c2dd, 32'h0, 32'h0, 32'h42456fee, 32'h422ebdf4, 32'h42652820, 32'h4283036d, 32'h4299e6d9};
test_input[29736:29743] = '{32'hc2a8e195, 32'hc2835ad3, 32'hc23d2f2d, 32'h42c7efa9, 32'h42282229, 32'hc2c51e35, 32'hc2abe177, 32'h427332a9};
test_output[29736:29743] = '{32'h0, 32'h0, 32'h0, 32'h42c7efa9, 32'h42282229, 32'h0, 32'h0, 32'h427332a9};
test_input[29744:29751] = '{32'h42871162, 32'hc28a2f97, 32'hc22dbee2, 32'hc27c1d10, 32'hc1d3de61, 32'h4249f9c0, 32'hc2a526b7, 32'h41fd705d};
test_output[29744:29751] = '{32'h42871162, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4249f9c0, 32'h0, 32'h41fd705d};
test_input[29752:29759] = '{32'hc207d072, 32'hc2ba6615, 32'h421e8c0c, 32'h428f07c9, 32'h427b8685, 32'hc272bfb6, 32'hc22a0bfc, 32'h41d0063e};
test_output[29752:29759] = '{32'h0, 32'h0, 32'h421e8c0c, 32'h428f07c9, 32'h427b8685, 32'h0, 32'h0, 32'h41d0063e};
test_input[29760:29767] = '{32'hc297fa35, 32'hc190f618, 32'hc2c2f971, 32'hc2abafeb, 32'hc0ba20a1, 32'h4216dccf, 32'h42a51d1a, 32'h429d4ae0};
test_output[29760:29767] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4216dccf, 32'h42a51d1a, 32'h429d4ae0};
test_input[29768:29775] = '{32'h42290653, 32'hc281998b, 32'hc2938ecb, 32'hc23ddd41, 32'hc2940214, 32'hc17bc2df, 32'hc223f3ee, 32'h41682d84};
test_output[29768:29775] = '{32'h42290653, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41682d84};
test_input[29776:29783] = '{32'h4239691c, 32'h42244670, 32'h422d3e03, 32'h4197b607, 32'hc294154b, 32'h429d4df0, 32'hc1e8a66a, 32'h41f8ddaf};
test_output[29776:29783] = '{32'h4239691c, 32'h42244670, 32'h422d3e03, 32'h4197b607, 32'h0, 32'h429d4df0, 32'h0, 32'h41f8ddaf};
test_input[29784:29791] = '{32'hbe09cc60, 32'h42147fab, 32'h4212264b, 32'h42b3eff8, 32'h3fc228b4, 32'hc287dc42, 32'h429bc0bd, 32'h40744782};
test_output[29784:29791] = '{32'h0, 32'h42147fab, 32'h4212264b, 32'h42b3eff8, 32'h3fc228b4, 32'h0, 32'h429bc0bd, 32'h40744782};
test_input[29792:29799] = '{32'hc1f35013, 32'hbf94b71b, 32'h41fec9e5, 32'hc28b5f02, 32'h428609f8, 32'h42c64c2a, 32'hc293abbc, 32'hc22a0fbf};
test_output[29792:29799] = '{32'h0, 32'h0, 32'h41fec9e5, 32'h0, 32'h428609f8, 32'h42c64c2a, 32'h0, 32'h0};
test_input[29800:29807] = '{32'hc0307f46, 32'hc29ac8ef, 32'hc1275edf, 32'hc20af9d4, 32'h42bb4552, 32'hc18c0cbb, 32'h42603447, 32'hc2289258};
test_output[29800:29807] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42bb4552, 32'h0, 32'h42603447, 32'h0};
test_input[29808:29815] = '{32'hc2857f83, 32'h422686f9, 32'hc2b5c285, 32'h41eb28ec, 32'hc2aeced0, 32'h41abb0de, 32'h41bad0b7, 32'h424df457};
test_output[29808:29815] = '{32'h0, 32'h422686f9, 32'h0, 32'h41eb28ec, 32'h0, 32'h41abb0de, 32'h41bad0b7, 32'h424df457};
test_input[29816:29823] = '{32'h425775d0, 32'h42c4941e, 32'h4235ddd4, 32'h4298e8f0, 32'h42baa802, 32'hc2b7ec4c, 32'hc2c609bc, 32'hc236ac69};
test_output[29816:29823] = '{32'h425775d0, 32'h42c4941e, 32'h4235ddd4, 32'h4298e8f0, 32'h42baa802, 32'h0, 32'h0, 32'h0};
test_input[29824:29831] = '{32'hc29e7d63, 32'h42c045e1, 32'hc162e7c7, 32'h4230d324, 32'hc144b6db, 32'h42c2d808, 32'hc2af744f, 32'hc28deb18};
test_output[29824:29831] = '{32'h0, 32'h42c045e1, 32'h0, 32'h4230d324, 32'h0, 32'h42c2d808, 32'h0, 32'h0};
test_input[29832:29839] = '{32'hc2a45e08, 32'h40fcc568, 32'hc24c8eda, 32'hc22dd4e3, 32'hc21ac401, 32'hc2bddbb3, 32'hc176d9f6, 32'hc20749d0};
test_output[29832:29839] = '{32'h0, 32'h40fcc568, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29840:29847] = '{32'hc28cf7da, 32'h427769f0, 32'h4223ae84, 32'h4141224e, 32'hc231cf16, 32'hc2bef790, 32'hc2b29454, 32'hc25e1a80};
test_output[29840:29847] = '{32'h0, 32'h427769f0, 32'h4223ae84, 32'h4141224e, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29848:29855] = '{32'hc2c414b9, 32'hc29bbd12, 32'h42af92fc, 32'hc2994d55, 32'hc221c5ec, 32'hc21ab571, 32'h4166c185, 32'hc1d13b2d};
test_output[29848:29855] = '{32'h0, 32'h0, 32'h42af92fc, 32'h0, 32'h0, 32'h0, 32'h4166c185, 32'h0};
test_input[29856:29863] = '{32'hc194f5da, 32'hbe458aea, 32'h4296a907, 32'hc2335177, 32'h4245a9ce, 32'hc263d165, 32'hc29a326e, 32'hc2881368};
test_output[29856:29863] = '{32'h0, 32'h0, 32'h4296a907, 32'h0, 32'h4245a9ce, 32'h0, 32'h0, 32'h0};
test_input[29864:29871] = '{32'h3f4f7de7, 32'hc02f9e93, 32'h42aeded4, 32'hc20b894d, 32'h40061d2d, 32'h404da9f5, 32'hc2298e0a, 32'hc2c11297};
test_output[29864:29871] = '{32'h3f4f7de7, 32'h0, 32'h42aeded4, 32'h0, 32'h40061d2d, 32'h404da9f5, 32'h0, 32'h0};
test_input[29872:29879] = '{32'hc2bef0bb, 32'h426158cd, 32'h4296c12a, 32'hc21194c2, 32'h4276f5ab, 32'h42a850f5, 32'hc185fb67, 32'h42bcfd08};
test_output[29872:29879] = '{32'h0, 32'h426158cd, 32'h4296c12a, 32'h0, 32'h4276f5ab, 32'h42a850f5, 32'h0, 32'h42bcfd08};
test_input[29880:29887] = '{32'hc232156e, 32'h414d3549, 32'hc293fccf, 32'h42663f2d, 32'hc1ea4190, 32'h418e3670, 32'hc25093c4, 32'h427cd5b9};
test_output[29880:29887] = '{32'h0, 32'h414d3549, 32'h0, 32'h42663f2d, 32'h0, 32'h418e3670, 32'h0, 32'h427cd5b9};
test_input[29888:29895] = '{32'h42c74873, 32'h42460df2, 32'h42bc0c1e, 32'h428e4151, 32'h4291faf4, 32'h42abceab, 32'h425a1159, 32'hc12068ab};
test_output[29888:29895] = '{32'h42c74873, 32'h42460df2, 32'h42bc0c1e, 32'h428e4151, 32'h4291faf4, 32'h42abceab, 32'h425a1159, 32'h0};
test_input[29896:29903] = '{32'h3fb67ed6, 32'h429ca5a4, 32'h42809f71, 32'hc026e449, 32'hc22c8fdc, 32'hc2708a33, 32'h41da595f, 32'h418e3d9a};
test_output[29896:29903] = '{32'h3fb67ed6, 32'h429ca5a4, 32'h42809f71, 32'h0, 32'h0, 32'h0, 32'h41da595f, 32'h418e3d9a};
test_input[29904:29911] = '{32'h40c4d8ce, 32'h42658bd3, 32'hc2948813, 32'hc27afcbd, 32'hc2003b6f, 32'hc1f5dccf, 32'hc2aa3b69, 32'h429b8861};
test_output[29904:29911] = '{32'h40c4d8ce, 32'h42658bd3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429b8861};
test_input[29912:29919] = '{32'h3fbcb43a, 32'hc20f098a, 32'hc2bca6f6, 32'h4169ce9b, 32'h420e24ab, 32'h42581698, 32'hc29e8e06, 32'hc2c198d5};
test_output[29912:29919] = '{32'h3fbcb43a, 32'h0, 32'h0, 32'h4169ce9b, 32'h420e24ab, 32'h42581698, 32'h0, 32'h0};
test_input[29920:29927] = '{32'h419d4cfd, 32'h42b0bb9b, 32'h42c1e48b, 32'h419e0b8c, 32'hc2bbd714, 32'h42ae6409, 32'hc220ce4d, 32'hc2b404b3};
test_output[29920:29927] = '{32'h419d4cfd, 32'h42b0bb9b, 32'h42c1e48b, 32'h419e0b8c, 32'h0, 32'h42ae6409, 32'h0, 32'h0};
test_input[29928:29935] = '{32'h42197546, 32'h40472164, 32'hc21883cf, 32'hc1e9cc0c, 32'h4275da8e, 32'hc26764c8, 32'hc2059ad4, 32'hc2170086};
test_output[29928:29935] = '{32'h42197546, 32'h40472164, 32'h0, 32'h0, 32'h4275da8e, 32'h0, 32'h0, 32'h0};
test_input[29936:29943] = '{32'h42761f64, 32'h41f72ca3, 32'hc113aa03, 32'h421f60b8, 32'h42abd1b0, 32'hc26dd9b5, 32'h410a77ab, 32'h42340f4e};
test_output[29936:29943] = '{32'h42761f64, 32'h41f72ca3, 32'h0, 32'h421f60b8, 32'h42abd1b0, 32'h0, 32'h410a77ab, 32'h42340f4e};
test_input[29944:29951] = '{32'hc285836c, 32'hc16b22d4, 32'h423c75d0, 32'hc2285b4d, 32'hc2509092, 32'hc2629bdb, 32'hc2903c5b, 32'h4156e435};
test_output[29944:29951] = '{32'h0, 32'h0, 32'h423c75d0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4156e435};
test_input[29952:29959] = '{32'hc1c65c2b, 32'h4248cc61, 32'h422e8ed4, 32'hc294cbf1, 32'hc2708246, 32'hc299f2e1, 32'h41d085ca, 32'hc2adfc62};
test_output[29952:29959] = '{32'h0, 32'h4248cc61, 32'h422e8ed4, 32'h0, 32'h0, 32'h0, 32'h41d085ca, 32'h0};
test_input[29960:29967] = '{32'h429d81fb, 32'hc235b8e1, 32'hc20e4dba, 32'hc28bcac5, 32'hc28f0fe9, 32'hc1b9f329, 32'hc1053188, 32'h42223f43};
test_output[29960:29967] = '{32'h429d81fb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42223f43};
test_input[29968:29975] = '{32'h423a3992, 32'hc1ac4aab, 32'hc1eae29f, 32'h401e5663, 32'h420a3e6d, 32'h418e8664, 32'h428fc5b3, 32'hc2bfb3c6};
test_output[29968:29975] = '{32'h423a3992, 32'h0, 32'h0, 32'h401e5663, 32'h420a3e6d, 32'h418e8664, 32'h428fc5b3, 32'h0};
test_input[29976:29983] = '{32'h4236421a, 32'hc22715f8, 32'h427b2580, 32'h42458fc0, 32'h423840b9, 32'hc1bc8fda, 32'hc13718bd, 32'h400e41bf};
test_output[29976:29983] = '{32'h4236421a, 32'h0, 32'h427b2580, 32'h42458fc0, 32'h423840b9, 32'h0, 32'h0, 32'h400e41bf};
test_input[29984:29991] = '{32'hc1713094, 32'h408a1960, 32'hc1daa0e1, 32'h41fdfcd9, 32'hc2037450, 32'h4204b531, 32'h3f20b710, 32'h41fc7bba};
test_output[29984:29991] = '{32'h0, 32'h408a1960, 32'h0, 32'h41fdfcd9, 32'h0, 32'h4204b531, 32'h3f20b710, 32'h41fc7bba};
test_input[29992:29999] = '{32'hc16d1858, 32'hc22f85a3, 32'h42738cfe, 32'hc2aa8512, 32'hc235636c, 32'h423295b6, 32'h406eb58c, 32'hc24d340b};
test_output[29992:29999] = '{32'h0, 32'h0, 32'h42738cfe, 32'h0, 32'h0, 32'h423295b6, 32'h406eb58c, 32'h0};
test_input[30000:30007] = '{32'hc1ea96ac, 32'hc20550ff, 32'hc2415a70, 32'h42a7dcf9, 32'h41b438cb, 32'hc1a5ce01, 32'hc2ab061d, 32'h41fe11db};
test_output[30000:30007] = '{32'h0, 32'h0, 32'h0, 32'h42a7dcf9, 32'h41b438cb, 32'h0, 32'h0, 32'h41fe11db};
test_input[30008:30015] = '{32'hc1121a33, 32'h422b9941, 32'hc2c505ca, 32'hc20efe38, 32'h4297c451, 32'h41355e76, 32'hc22db92d, 32'h3fce93f2};
test_output[30008:30015] = '{32'h0, 32'h422b9941, 32'h0, 32'h0, 32'h4297c451, 32'h41355e76, 32'h0, 32'h3fce93f2};
test_input[30016:30023] = '{32'hc2abbecb, 32'h42c12d58, 32'h4284aefc, 32'h41569efd, 32'h403d7a86, 32'h41ab4743, 32'hc27d6d62, 32'h42acbbac};
test_output[30016:30023] = '{32'h0, 32'h42c12d58, 32'h4284aefc, 32'h41569efd, 32'h403d7a86, 32'h41ab4743, 32'h0, 32'h42acbbac};
test_input[30024:30031] = '{32'h42992c32, 32'hc298ca6d, 32'h404f9ea5, 32'hc0aab3f6, 32'hc2906212, 32'h4243051b, 32'h419439d6, 32'hc15f416a};
test_output[30024:30031] = '{32'h42992c32, 32'h0, 32'h404f9ea5, 32'h0, 32'h0, 32'h4243051b, 32'h419439d6, 32'h0};
test_input[30032:30039] = '{32'h41e9379a, 32'h427e9028, 32'hc2503b53, 32'h4282a051, 32'h409c304d, 32'hc25c4bc2, 32'h423a1df2, 32'h42a0008a};
test_output[30032:30039] = '{32'h41e9379a, 32'h427e9028, 32'h0, 32'h4282a051, 32'h409c304d, 32'h0, 32'h423a1df2, 32'h42a0008a};
test_input[30040:30047] = '{32'hc2b20fa6, 32'hc099ce07, 32'h4281ed33, 32'h42b1faf8, 32'hc2451aa5, 32'hc28985ea, 32'h423867c5, 32'h41c5599e};
test_output[30040:30047] = '{32'h0, 32'h0, 32'h4281ed33, 32'h42b1faf8, 32'h0, 32'h0, 32'h423867c5, 32'h41c5599e};
test_input[30048:30055] = '{32'h4114796e, 32'hc187dcca, 32'h424f082d, 32'hc290ebb0, 32'hc2c0e73b, 32'h425a902b, 32'h42a8206d, 32'h428f6eff};
test_output[30048:30055] = '{32'h4114796e, 32'h0, 32'h424f082d, 32'h0, 32'h0, 32'h425a902b, 32'h42a8206d, 32'h428f6eff};
test_input[30056:30063] = '{32'h42c0fad6, 32'h425dda9f, 32'h42030dc2, 32'h4207cc92, 32'hc2b8c432, 32'hc093b325, 32'hc2c39945, 32'h41fe03ac};
test_output[30056:30063] = '{32'h42c0fad6, 32'h425dda9f, 32'h42030dc2, 32'h4207cc92, 32'h0, 32'h0, 32'h0, 32'h41fe03ac};
test_input[30064:30071] = '{32'hc12ca1b7, 32'hc2c028ef, 32'hc2c22aca, 32'h423e7b4f, 32'hc29721f4, 32'h42997150, 32'h42219a6c, 32'h42504897};
test_output[30064:30071] = '{32'h0, 32'h0, 32'h0, 32'h423e7b4f, 32'h0, 32'h42997150, 32'h42219a6c, 32'h42504897};
test_input[30072:30079] = '{32'h42629304, 32'h4295bc09, 32'h42c48da9, 32'h41d9a157, 32'hc282bcd9, 32'h42c3a0f6, 32'h4210a512, 32'h41c13356};
test_output[30072:30079] = '{32'h42629304, 32'h4295bc09, 32'h42c48da9, 32'h41d9a157, 32'h0, 32'h42c3a0f6, 32'h4210a512, 32'h41c13356};
test_input[30080:30087] = '{32'h42b37dbe, 32'h4285b418, 32'h42bfecc5, 32'hc262fe34, 32'hc110277b, 32'h422be195, 32'hc1dd2005, 32'hc28ed410};
test_output[30080:30087] = '{32'h42b37dbe, 32'h4285b418, 32'h42bfecc5, 32'h0, 32'h0, 32'h422be195, 32'h0, 32'h0};
test_input[30088:30095] = '{32'hc2a7dd48, 32'h4291a16d, 32'h4294128a, 32'h420718c2, 32'hc2b83b3a, 32'h404e5b7c, 32'hc2957644, 32'hc158a715};
test_output[30088:30095] = '{32'h0, 32'h4291a16d, 32'h4294128a, 32'h420718c2, 32'h0, 32'h404e5b7c, 32'h0, 32'h0};
test_input[30096:30103] = '{32'hc1e3b597, 32'h417adc66, 32'hc24aafa1, 32'h42b1f39d, 32'h42669f1c, 32'hc254255d, 32'h423bf70e, 32'h41eec910};
test_output[30096:30103] = '{32'h0, 32'h417adc66, 32'h0, 32'h42b1f39d, 32'h42669f1c, 32'h0, 32'h423bf70e, 32'h41eec910};
test_input[30104:30111] = '{32'h42ad3e06, 32'h41acc41b, 32'h428cd686, 32'hc14b4804, 32'h41c9a7b9, 32'h41d8e2ff, 32'hc114ce70, 32'h4269c9d8};
test_output[30104:30111] = '{32'h42ad3e06, 32'h41acc41b, 32'h428cd686, 32'h0, 32'h41c9a7b9, 32'h41d8e2ff, 32'h0, 32'h4269c9d8};
test_input[30112:30119] = '{32'h42568b54, 32'h4188b6f8, 32'h42b1d0ac, 32'hc2ba2865, 32'h41f17034, 32'hc1e267eb, 32'hc206e0b7, 32'h4282d9dc};
test_output[30112:30119] = '{32'h42568b54, 32'h4188b6f8, 32'h42b1d0ac, 32'h0, 32'h41f17034, 32'h0, 32'h0, 32'h4282d9dc};
test_input[30120:30127] = '{32'hc1a77886, 32'hc212fc3f, 32'hc2214e9b, 32'h42b29deb, 32'hc23d0813, 32'h41e20dcb, 32'hc28906c0, 32'hc27f6ccd};
test_output[30120:30127] = '{32'h0, 32'h0, 32'h0, 32'h42b29deb, 32'h0, 32'h41e20dcb, 32'h0, 32'h0};
test_input[30128:30135] = '{32'hc223ca71, 32'h41de9a36, 32'hc23348de, 32'h4264213f, 32'hc2c51647, 32'hc269e2f9, 32'h428259be, 32'h42a283f5};
test_output[30128:30135] = '{32'h0, 32'h41de9a36, 32'h0, 32'h4264213f, 32'h0, 32'h0, 32'h428259be, 32'h42a283f5};
test_input[30136:30143] = '{32'hc21afeb8, 32'h4245b473, 32'hc282f091, 32'hc0bb57fe, 32'hc235e636, 32'hc2588d6d, 32'hc2bd7454, 32'h41a1501b};
test_output[30136:30143] = '{32'h0, 32'h4245b473, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41a1501b};
test_input[30144:30151] = '{32'hc14ce2d5, 32'h42a3a113, 32'hc254cc10, 32'hc2a9cd8e, 32'h42b858c4, 32'h40749aa5, 32'hc13fe82d, 32'h40b376b0};
test_output[30144:30151] = '{32'h0, 32'h42a3a113, 32'h0, 32'h0, 32'h42b858c4, 32'h40749aa5, 32'h0, 32'h40b376b0};
test_input[30152:30159] = '{32'hc100a0fa, 32'hc2c70277, 32'h429cd8e1, 32'h428122d8, 32'h42bfd1e0, 32'hc24dc1a6, 32'h42003615, 32'h428e7052};
test_output[30152:30159] = '{32'h0, 32'h0, 32'h429cd8e1, 32'h428122d8, 32'h42bfd1e0, 32'h0, 32'h42003615, 32'h428e7052};
test_input[30160:30167] = '{32'h4239f415, 32'hc23ac345, 32'h429bafa6, 32'h4131a88f, 32'hc206b5bd, 32'h40164d3e, 32'h42ae1e38, 32'hc2c5473f};
test_output[30160:30167] = '{32'h4239f415, 32'h0, 32'h429bafa6, 32'h4131a88f, 32'h0, 32'h40164d3e, 32'h42ae1e38, 32'h0};
test_input[30168:30175] = '{32'h42a06be3, 32'hc1507ff2, 32'hc2b1273d, 32'hc10cd866, 32'hc2a3b47a, 32'h41a0fb3d, 32'h421b07b7, 32'hc2b09f96};
test_output[30168:30175] = '{32'h42a06be3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41a0fb3d, 32'h421b07b7, 32'h0};
test_input[30176:30183] = '{32'h422b96ba, 32'hc22978c3, 32'h422b0c47, 32'hc224a193, 32'hc1ccbd01, 32'h4206121c, 32'h40cc8dfe, 32'hc16e8bbc};
test_output[30176:30183] = '{32'h422b96ba, 32'h0, 32'h422b0c47, 32'h0, 32'h0, 32'h4206121c, 32'h40cc8dfe, 32'h0};
test_input[30184:30191] = '{32'h41f85472, 32'hc1a05230, 32'h41a643f3, 32'h42b2be17, 32'hc2c5a310, 32'hc13f4a6f, 32'h422d7ec2, 32'h429653ca};
test_output[30184:30191] = '{32'h41f85472, 32'h0, 32'h41a643f3, 32'h42b2be17, 32'h0, 32'h0, 32'h422d7ec2, 32'h429653ca};
test_input[30192:30199] = '{32'hc2abb8a8, 32'h4283f6df, 32'hc2040f9c, 32'hc1861d7c, 32'hc14fdb50, 32'h415c8e16, 32'hc2c514b0, 32'h4229fd18};
test_output[30192:30199] = '{32'h0, 32'h4283f6df, 32'h0, 32'h0, 32'h0, 32'h415c8e16, 32'h0, 32'h4229fd18};
test_input[30200:30207] = '{32'hc2369bc3, 32'h4141bc3b, 32'hc2b7e3a1, 32'hc1907961, 32'h42ad61b8, 32'h4215f625, 32'h429db732, 32'hbf1ffa65};
test_output[30200:30207] = '{32'h0, 32'h4141bc3b, 32'h0, 32'h0, 32'h42ad61b8, 32'h4215f625, 32'h429db732, 32'h0};
test_input[30208:30215] = '{32'hc16cebe8, 32'h42498bd0, 32'h42632afd, 32'hc22cd63e, 32'hc1ec6088, 32'h42be7e9f, 32'h42855ed6, 32'hc230706e};
test_output[30208:30215] = '{32'h0, 32'h42498bd0, 32'h42632afd, 32'h0, 32'h0, 32'h42be7e9f, 32'h42855ed6, 32'h0};
test_input[30216:30223] = '{32'h4294b049, 32'hc1be9d31, 32'h424cbf49, 32'h42b5bec6, 32'h422d5941, 32'hc2b66db5, 32'hc2836830, 32'hc208222c};
test_output[30216:30223] = '{32'h4294b049, 32'h0, 32'h424cbf49, 32'h42b5bec6, 32'h422d5941, 32'h0, 32'h0, 32'h0};
test_input[30224:30231] = '{32'hc24fc061, 32'h41b1ef00, 32'h40ba9c8e, 32'h427f6ec0, 32'h41929a7f, 32'h414a82b5, 32'hc23b83cf, 32'h41c547dc};
test_output[30224:30231] = '{32'h0, 32'h41b1ef00, 32'h40ba9c8e, 32'h427f6ec0, 32'h41929a7f, 32'h414a82b5, 32'h0, 32'h41c547dc};
test_input[30232:30239] = '{32'h3f0cce92, 32'h429c09b2, 32'hc27c9703, 32'hc0ed0ab7, 32'hc28a2826, 32'hc296be6d, 32'hc279996b, 32'h42b4e343};
test_output[30232:30239] = '{32'h3f0cce92, 32'h429c09b2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b4e343};
test_input[30240:30247] = '{32'hc2a63bb8, 32'hc2b85a2c, 32'h42745064, 32'hc28e7078, 32'h4275f954, 32'hc12f3a3a, 32'h4117ab34, 32'hc217e4ca};
test_output[30240:30247] = '{32'h0, 32'h0, 32'h42745064, 32'h0, 32'h4275f954, 32'h0, 32'h4117ab34, 32'h0};
test_input[30248:30255] = '{32'hc21b5705, 32'hc22f9149, 32'hc22b5851, 32'hc2b35f0e, 32'hc2823fd1, 32'h4260cb56, 32'hc25ea9fa, 32'h42341538};
test_output[30248:30255] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4260cb56, 32'h0, 32'h42341538};
test_input[30256:30263] = '{32'hc2a7b46f, 32'h4248ed2c, 32'h42af6a5f, 32'h40d8162f, 32'hc0a618f1, 32'hbfc008b7, 32'h42276c28, 32'hc22da942};
test_output[30256:30263] = '{32'h0, 32'h4248ed2c, 32'h42af6a5f, 32'h40d8162f, 32'h0, 32'h0, 32'h42276c28, 32'h0};
test_input[30264:30271] = '{32'h42a0b7a4, 32'h429f6294, 32'hc2978289, 32'hc23e1962, 32'h414dfd1f, 32'h4297e6fa, 32'h41b48eef, 32'h423f89c5};
test_output[30264:30271] = '{32'h42a0b7a4, 32'h429f6294, 32'h0, 32'h0, 32'h414dfd1f, 32'h4297e6fa, 32'h41b48eef, 32'h423f89c5};
test_input[30272:30279] = '{32'h42661036, 32'hc26225cc, 32'hc244c28f, 32'h42525eed, 32'hc14168b0, 32'h410296cf, 32'hc2b94437, 32'hc26de4bb};
test_output[30272:30279] = '{32'h42661036, 32'h0, 32'h0, 32'h42525eed, 32'h0, 32'h410296cf, 32'h0, 32'h0};
test_input[30280:30287] = '{32'h429b9e27, 32'h426e0316, 32'h4188c6b7, 32'h41c745ae, 32'hc1d55a21, 32'hc24b1b4a, 32'hc2571330, 32'hc2bb01c9};
test_output[30280:30287] = '{32'h429b9e27, 32'h426e0316, 32'h4188c6b7, 32'h41c745ae, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30288:30295] = '{32'hc25d669b, 32'h427bde14, 32'hc2803665, 32'h4206d42f, 32'h428f050c, 32'h41108441, 32'hc1605a39, 32'hc1b607e9};
test_output[30288:30295] = '{32'h0, 32'h427bde14, 32'h0, 32'h4206d42f, 32'h428f050c, 32'h41108441, 32'h0, 32'h0};
test_input[30296:30303] = '{32'hc29e4f54, 32'h428a983d, 32'h418e9fbb, 32'h3f8f7697, 32'hc263ad17, 32'h42886754, 32'h42be81da, 32'hc2b201b1};
test_output[30296:30303] = '{32'h0, 32'h428a983d, 32'h418e9fbb, 32'h3f8f7697, 32'h0, 32'h42886754, 32'h42be81da, 32'h0};
test_input[30304:30311] = '{32'h41afd98a, 32'hc26f1489, 32'hc298a7d3, 32'hc271e08b, 32'h42c408c8, 32'hc25f405d, 32'hc26e8567, 32'hc177dda7};
test_output[30304:30311] = '{32'h41afd98a, 32'h0, 32'h0, 32'h0, 32'h42c408c8, 32'h0, 32'h0, 32'h0};
test_input[30312:30319] = '{32'hc29645e1, 32'hc249b2f4, 32'hc1b868aa, 32'hc17ef177, 32'h4280e633, 32'h41d62ff7, 32'h42a8453d, 32'h429aa108};
test_output[30312:30319] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4280e633, 32'h41d62ff7, 32'h42a8453d, 32'h429aa108};
test_input[30320:30327] = '{32'h42739e19, 32'h423b536e, 32'hc076a2a4, 32'h42c6360d, 32'h40dac6b3, 32'h420eaea3, 32'h4182dc3f, 32'h42338b4f};
test_output[30320:30327] = '{32'h42739e19, 32'h423b536e, 32'h0, 32'h42c6360d, 32'h40dac6b3, 32'h420eaea3, 32'h4182dc3f, 32'h42338b4f};
test_input[30328:30335] = '{32'hc1ef3289, 32'hc2b03ddf, 32'hc27bb6d4, 32'hc2c0b59c, 32'h428d6e2c, 32'hc2346602, 32'h429bee96, 32'h42b4fe65};
test_output[30328:30335] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h428d6e2c, 32'h0, 32'h429bee96, 32'h42b4fe65};
test_input[30336:30343] = '{32'h424af116, 32'h42c41915, 32'hc1ac453c, 32'h42645c6b, 32'hc2685698, 32'h421bd119, 32'hc2271ff1, 32'h419e769d};
test_output[30336:30343] = '{32'h424af116, 32'h42c41915, 32'h0, 32'h42645c6b, 32'h0, 32'h421bd119, 32'h0, 32'h419e769d};
test_input[30344:30351] = '{32'hc27ec3a0, 32'h42393998, 32'h41c3d5d8, 32'hc16f7ca8, 32'h4270d434, 32'h4160f478, 32'h42a2c82b, 32'hc1922d47};
test_output[30344:30351] = '{32'h0, 32'h42393998, 32'h41c3d5d8, 32'h0, 32'h4270d434, 32'h4160f478, 32'h42a2c82b, 32'h0};
test_input[30352:30359] = '{32'hc0d4b82c, 32'h40ef710d, 32'hc285043a, 32'h41d5ef49, 32'hc07fbf5e, 32'h428a3924, 32'h40b9523c, 32'h428a8a1b};
test_output[30352:30359] = '{32'h0, 32'h40ef710d, 32'h0, 32'h41d5ef49, 32'h0, 32'h428a3924, 32'h40b9523c, 32'h428a8a1b};
test_input[30360:30367] = '{32'hc1426f97, 32'h4290531d, 32'hc172cdda, 32'h42614ec7, 32'hc2bbc256, 32'hc28085ed, 32'hc1e64df8, 32'hc20e0cf1};
test_output[30360:30367] = '{32'h0, 32'h4290531d, 32'h0, 32'h42614ec7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30368:30375] = '{32'hc2a90150, 32'hc21d0113, 32'h4206a43f, 32'hc2b4e4ed, 32'h42b4ddcf, 32'h428c3fb9, 32'h42c17ac2, 32'h42b988ef};
test_output[30368:30375] = '{32'h0, 32'h0, 32'h4206a43f, 32'h0, 32'h42b4ddcf, 32'h428c3fb9, 32'h42c17ac2, 32'h42b988ef};
test_input[30376:30383] = '{32'h41bf37f2, 32'hc216fa3f, 32'hc27394fb, 32'hc21437bc, 32'h4296e850, 32'hc2722c0d, 32'h405eab42, 32'hc2978322};
test_output[30376:30383] = '{32'h41bf37f2, 32'h0, 32'h0, 32'h0, 32'h4296e850, 32'h0, 32'h405eab42, 32'h0};
test_input[30384:30391] = '{32'h411244b1, 32'h41685c9b, 32'h428baf00, 32'h42b66ccc, 32'hc0ac2316, 32'h428ac2b5, 32'hc14ca0de, 32'h428f3eb5};
test_output[30384:30391] = '{32'h411244b1, 32'h41685c9b, 32'h428baf00, 32'h42b66ccc, 32'h0, 32'h428ac2b5, 32'h0, 32'h428f3eb5};
test_input[30392:30399] = '{32'hc12c3b6c, 32'h42b5d689, 32'hc1b4b414, 32'h42972346, 32'h42612613, 32'hc249419c, 32'hc2ae0e01, 32'h42b37edf};
test_output[30392:30399] = '{32'h0, 32'h42b5d689, 32'h0, 32'h42972346, 32'h42612613, 32'h0, 32'h0, 32'h42b37edf};
test_input[30400:30407] = '{32'hc274da20, 32'h41cd0c79, 32'h422fbdd5, 32'hc18b8917, 32'hc2aa6c17, 32'hc2ace6af, 32'h423de9ac, 32'h42277075};
test_output[30400:30407] = '{32'h0, 32'h41cd0c79, 32'h422fbdd5, 32'h0, 32'h0, 32'h0, 32'h423de9ac, 32'h42277075};
test_input[30408:30415] = '{32'hc1d4ba74, 32'hc1cf139f, 32'hc1202eba, 32'hc2c38dc0, 32'hc2bc07f5, 32'hc1a4410b, 32'h42a9ae0a, 32'hc281881f};
test_output[30408:30415] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a9ae0a, 32'h0};
test_input[30416:30423] = '{32'h42477b9e, 32'hc270cf81, 32'h40a99f69, 32'h426df4da, 32'h4159c148, 32'h3fe4d04b, 32'hc1afea49, 32'h40e203dd};
test_output[30416:30423] = '{32'h42477b9e, 32'h0, 32'h40a99f69, 32'h426df4da, 32'h4159c148, 32'h3fe4d04b, 32'h0, 32'h40e203dd};
test_input[30424:30431] = '{32'hc26fb644, 32'h40c62ff4, 32'hc28f298b, 32'hc198de9e, 32'h426fdffc, 32'h4183b5c9, 32'hc29bd779, 32'h412e0e81};
test_output[30424:30431] = '{32'h0, 32'h40c62ff4, 32'h0, 32'h0, 32'h426fdffc, 32'h4183b5c9, 32'h0, 32'h412e0e81};
test_input[30432:30439] = '{32'h4254e220, 32'h411529a9, 32'hc111c148, 32'hc1c1c78b, 32'hc277bf25, 32'h42a2decb, 32'hc288d088, 32'hc25b77bb};
test_output[30432:30439] = '{32'h4254e220, 32'h411529a9, 32'h0, 32'h0, 32'h0, 32'h42a2decb, 32'h0, 32'h0};
test_input[30440:30447] = '{32'h41c7d6e7, 32'hc17dc905, 32'hc1354767, 32'hc1b53f1f, 32'hc2051d89, 32'hc25c5772, 32'h424ea2e4, 32'h42189a46};
test_output[30440:30447] = '{32'h41c7d6e7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h424ea2e4, 32'h42189a46};
test_input[30448:30455] = '{32'h427ab899, 32'hc27cddef, 32'h416866ef, 32'hc2bef71f, 32'hc2624d51, 32'hc1eca743, 32'h4181e3b9, 32'hc196db97};
test_output[30448:30455] = '{32'h427ab899, 32'h0, 32'h416866ef, 32'h0, 32'h0, 32'h0, 32'h4181e3b9, 32'h0};
test_input[30456:30463] = '{32'h428adf6b, 32'hc24c6c55, 32'h41b74478, 32'hbfc41dde, 32'hc28fd65b, 32'hc2b809f2, 32'hc1c2788f, 32'h42465484};
test_output[30456:30463] = '{32'h428adf6b, 32'h0, 32'h41b74478, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42465484};
test_input[30464:30471] = '{32'h418f7863, 32'h414f7ec8, 32'h42bbcb5c, 32'hc2801b7a, 32'h42874337, 32'h420b9d6d, 32'hc1044458, 32'hc02a28ad};
test_output[30464:30471] = '{32'h418f7863, 32'h414f7ec8, 32'h42bbcb5c, 32'h0, 32'h42874337, 32'h420b9d6d, 32'h0, 32'h0};
test_input[30472:30479] = '{32'h428e3e9c, 32'h4231f19d, 32'h4252e93b, 32'hc2842ad9, 32'h41e0cd86, 32'hc2bbc3de, 32'h42bd6656, 32'h42886893};
test_output[30472:30479] = '{32'h428e3e9c, 32'h4231f19d, 32'h4252e93b, 32'h0, 32'h41e0cd86, 32'h0, 32'h42bd6656, 32'h42886893};
test_input[30480:30487] = '{32'h4231dde0, 32'h4285c459, 32'hc289ba87, 32'hc23c0b75, 32'hc1d8cf06, 32'h42b10c40, 32'hc158099b, 32'hc2c5a157};
test_output[30480:30487] = '{32'h4231dde0, 32'h4285c459, 32'h0, 32'h0, 32'h0, 32'h42b10c40, 32'h0, 32'h0};
test_input[30488:30495] = '{32'h42042341, 32'h42b15d46, 32'h415a0ae2, 32'h411e3ea7, 32'hc290848d, 32'hc276a947, 32'h420a9d7e, 32'hc0d21ea5};
test_output[30488:30495] = '{32'h42042341, 32'h42b15d46, 32'h415a0ae2, 32'h411e3ea7, 32'h0, 32'h0, 32'h420a9d7e, 32'h0};
test_input[30496:30503] = '{32'h4197bd26, 32'hc23b0959, 32'h41ca4678, 32'hc1e10f00, 32'hc2a0dd80, 32'h40f8083a, 32'h42626260, 32'h41aab622};
test_output[30496:30503] = '{32'h4197bd26, 32'h0, 32'h41ca4678, 32'h0, 32'h0, 32'h40f8083a, 32'h42626260, 32'h41aab622};
test_input[30504:30511] = '{32'hc20457ec, 32'h42803169, 32'hc2a5759a, 32'h42ada920, 32'h4285c973, 32'h42b15673, 32'h4234edc1, 32'h4192d8ed};
test_output[30504:30511] = '{32'h0, 32'h42803169, 32'h0, 32'h42ada920, 32'h4285c973, 32'h42b15673, 32'h4234edc1, 32'h4192d8ed};
test_input[30512:30519] = '{32'h4294bf77, 32'hc2a3cf33, 32'h42413ef7, 32'h42c5c010, 32'h42313bfc, 32'hc28aa8ff, 32'h40e699d3, 32'hc1caeb70};
test_output[30512:30519] = '{32'h4294bf77, 32'h0, 32'h42413ef7, 32'h42c5c010, 32'h42313bfc, 32'h0, 32'h40e699d3, 32'h0};
test_input[30520:30527] = '{32'hc28b8db4, 32'hc13c0a1a, 32'h42ad0ec9, 32'h425bc5da, 32'hc160cc82, 32'h41eb5d72, 32'hc2adfb7b, 32'h41cc2d71};
test_output[30520:30527] = '{32'h0, 32'h0, 32'h42ad0ec9, 32'h425bc5da, 32'h0, 32'h41eb5d72, 32'h0, 32'h41cc2d71};
test_input[30528:30535] = '{32'hc2241a43, 32'hc274cce2, 32'hc101bfb6, 32'h424094cb, 32'h42a5af84, 32'hc2800a9f, 32'hc09d36ba, 32'h4216e2ef};
test_output[30528:30535] = '{32'h0, 32'h0, 32'h0, 32'h424094cb, 32'h42a5af84, 32'h0, 32'h0, 32'h4216e2ef};
test_input[30536:30543] = '{32'h40d5b8d1, 32'h42873ef2, 32'h41219a39, 32'hc12aa12b, 32'h429da851, 32'h420545ea, 32'hc12712d6, 32'h422da210};
test_output[30536:30543] = '{32'h40d5b8d1, 32'h42873ef2, 32'h41219a39, 32'h0, 32'h429da851, 32'h420545ea, 32'h0, 32'h422da210};
test_input[30544:30551] = '{32'hc1a6c292, 32'h4286ae68, 32'h41233ec3, 32'hc231f4fe, 32'h419972c1, 32'h427ba65a, 32'h414cbaa6, 32'h41d27846};
test_output[30544:30551] = '{32'h0, 32'h4286ae68, 32'h41233ec3, 32'h0, 32'h419972c1, 32'h427ba65a, 32'h414cbaa6, 32'h41d27846};
test_input[30552:30559] = '{32'h42ad51e8, 32'h425fcfeb, 32'hc28e1dea, 32'h41bb7538, 32'h4254d5d3, 32'h4119f621, 32'h41d346e2, 32'h428ff690};
test_output[30552:30559] = '{32'h42ad51e8, 32'h425fcfeb, 32'h0, 32'h41bb7538, 32'h4254d5d3, 32'h4119f621, 32'h41d346e2, 32'h428ff690};
test_input[30560:30567] = '{32'h4220bf43, 32'h42616ccb, 32'hc1d01366, 32'h42745f81, 32'h4278c017, 32'hc1ef3627, 32'hc29ec5bd, 32'h42c4f54d};
test_output[30560:30567] = '{32'h4220bf43, 32'h42616ccb, 32'h0, 32'h42745f81, 32'h4278c017, 32'h0, 32'h0, 32'h42c4f54d};
test_input[30568:30575] = '{32'hc1a3e97e, 32'hc28c2aba, 32'h42baef09, 32'hc2680e47, 32'hc17296f8, 32'hc1f1face, 32'hc25680b2, 32'h42a23e5f};
test_output[30568:30575] = '{32'h0, 32'h0, 32'h42baef09, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a23e5f};
test_input[30576:30583] = '{32'h42963033, 32'h428bc1d5, 32'hc27d72aa, 32'h42a36496, 32'h42a55f5c, 32'hc2b52d8f, 32'hc2b603b9, 32'hbd28beb1};
test_output[30576:30583] = '{32'h42963033, 32'h428bc1d5, 32'h0, 32'h42a36496, 32'h42a55f5c, 32'h0, 32'h0, 32'h0};
test_input[30584:30591] = '{32'h4297a0b1, 32'h429a892a, 32'hc0807f73, 32'h423af582, 32'hc1dabf9a, 32'h40277966, 32'h42527c4d, 32'h4151be93};
test_output[30584:30591] = '{32'h4297a0b1, 32'h429a892a, 32'h0, 32'h423af582, 32'h0, 32'h40277966, 32'h42527c4d, 32'h4151be93};
test_input[30592:30599] = '{32'h42087131, 32'hc10819bd, 32'hc218c381, 32'h41f7bf2c, 32'hc27b75df, 32'h42939e34, 32'hc2a783b7, 32'h4169de32};
test_output[30592:30599] = '{32'h42087131, 32'h0, 32'h0, 32'h41f7bf2c, 32'h0, 32'h42939e34, 32'h0, 32'h4169de32};
test_input[30600:30607] = '{32'h429c8e60, 32'hc2b4568f, 32'h41d198c1, 32'h42acb4e4, 32'h42a4fcb5, 32'h408b45bd, 32'hc17c670b, 32'hc2a5348e};
test_output[30600:30607] = '{32'h429c8e60, 32'h0, 32'h41d198c1, 32'h42acb4e4, 32'h42a4fcb5, 32'h408b45bd, 32'h0, 32'h0};
test_input[30608:30615] = '{32'hc28e2dee, 32'h424d4b59, 32'h42c219a4, 32'hc21f21e3, 32'h41ba9732, 32'h42967e70, 32'hc281a3dd, 32'h41c670ef};
test_output[30608:30615] = '{32'h0, 32'h424d4b59, 32'h42c219a4, 32'h0, 32'h41ba9732, 32'h42967e70, 32'h0, 32'h41c670ef};
test_input[30616:30623] = '{32'hc15881e5, 32'hc2a79e14, 32'h41c36f67, 32'hc2a14526, 32'hc29b6a2c, 32'hc28c4321, 32'hc2a1ea09, 32'h4226afdd};
test_output[30616:30623] = '{32'h0, 32'h0, 32'h41c36f67, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4226afdd};
test_input[30624:30631] = '{32'h428f8769, 32'h41ef9fb1, 32'h4255e5b9, 32'hc292471d, 32'h4286273d, 32'hc1e785f6, 32'h41edd747, 32'h4273eb4f};
test_output[30624:30631] = '{32'h428f8769, 32'h41ef9fb1, 32'h4255e5b9, 32'h0, 32'h4286273d, 32'h0, 32'h41edd747, 32'h4273eb4f};
test_input[30632:30639] = '{32'h419b7696, 32'hc2544ef1, 32'h42bce5c4, 32'hc2c2f315, 32'h42b2fae1, 32'hc2621790, 32'h42b6684e, 32'h42bfef31};
test_output[30632:30639] = '{32'h419b7696, 32'h0, 32'h42bce5c4, 32'h0, 32'h42b2fae1, 32'h0, 32'h42b6684e, 32'h42bfef31};
test_input[30640:30647] = '{32'hc24b2b10, 32'hc24d1973, 32'hc2b419b2, 32'hc1c1b9bd, 32'h41d5b90b, 32'h42940f7c, 32'hc19998fe, 32'h428748ca};
test_output[30640:30647] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41d5b90b, 32'h42940f7c, 32'h0, 32'h428748ca};
test_input[30648:30655] = '{32'h41f25971, 32'hc23fda84, 32'hc2203cbc, 32'h42b46668, 32'h42b1eb1d, 32'h408cc9b2, 32'h412f3a9c, 32'h4295031a};
test_output[30648:30655] = '{32'h41f25971, 32'h0, 32'h0, 32'h42b46668, 32'h42b1eb1d, 32'h408cc9b2, 32'h412f3a9c, 32'h4295031a};
test_input[30656:30663] = '{32'hc2ad42f5, 32'h428f4538, 32'h424eedbc, 32'hc285fb11, 32'h416b16c5, 32'hc15afd63, 32'hc25c1d43, 32'hc1f5c4c1};
test_output[30656:30663] = '{32'h0, 32'h428f4538, 32'h424eedbc, 32'h0, 32'h416b16c5, 32'h0, 32'h0, 32'h0};
test_input[30664:30671] = '{32'hc206d84c, 32'h42920e1f, 32'h42a9a901, 32'hc2b7dc5c, 32'h427dca52, 32'hc1ccc61c, 32'hc26fa7f3, 32'hc0b6125c};
test_output[30664:30671] = '{32'h0, 32'h42920e1f, 32'h42a9a901, 32'h0, 32'h427dca52, 32'h0, 32'h0, 32'h0};
test_input[30672:30679] = '{32'hc2a8627b, 32'h424ca8a3, 32'hc2815e2c, 32'h426bb936, 32'hc2a5eda2, 32'hc296d4e3, 32'hc299ed9d, 32'hc1cd8214};
test_output[30672:30679] = '{32'h0, 32'h424ca8a3, 32'h0, 32'h426bb936, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30680:30687] = '{32'hc22ff628, 32'hc18bb56f, 32'hc251da34, 32'h42bd7723, 32'hc1a0f914, 32'hc1c9d2ad, 32'hc1014c57, 32'hc203311b};
test_output[30680:30687] = '{32'h0, 32'h0, 32'h0, 32'h42bd7723, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30688:30695] = '{32'h42879aa6, 32'hc21ec1ed, 32'h42c004a3, 32'h4295b1a1, 32'h421a53f5, 32'hc1650ab3, 32'hc1e2306f, 32'hc21a91ce};
test_output[30688:30695] = '{32'h42879aa6, 32'h0, 32'h42c004a3, 32'h4295b1a1, 32'h421a53f5, 32'h0, 32'h0, 32'h0};
test_input[30696:30703] = '{32'hc281040d, 32'hc2560f4b, 32'hc2c3f4c4, 32'hc1bc0180, 32'h42badeb0, 32'hc21e3d9c, 32'hc0cec39b, 32'h42c312d8};
test_output[30696:30703] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42badeb0, 32'h0, 32'h0, 32'h42c312d8};
test_input[30704:30711] = '{32'hc227d6ba, 32'hc2b7618b, 32'hc2a17c4e, 32'hc299c31e, 32'hc2640f1b, 32'h42b955cc, 32'hc2549d2d, 32'h41d856c3};
test_output[30704:30711] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b955cc, 32'h0, 32'h41d856c3};
test_input[30712:30719] = '{32'h41b2d26b, 32'h42ab0d5e, 32'hc2b5c1ad, 32'h42560d21, 32'h424158d5, 32'hc2827ad5, 32'hc21b788b, 32'h42c47760};
test_output[30712:30719] = '{32'h41b2d26b, 32'h42ab0d5e, 32'h0, 32'h42560d21, 32'h424158d5, 32'h0, 32'h0, 32'h42c47760};
test_input[30720:30727] = '{32'h4267cf53, 32'hc2c095cc, 32'h40509e00, 32'hc2c5bd1d, 32'h42a839b1, 32'h418cf56f, 32'h41dc4d2a, 32'hc295997f};
test_output[30720:30727] = '{32'h4267cf53, 32'h0, 32'h40509e00, 32'h0, 32'h42a839b1, 32'h418cf56f, 32'h41dc4d2a, 32'h0};
test_input[30728:30735] = '{32'h42bc7d26, 32'hc0e2a567, 32'hc296f5f0, 32'h400f0d90, 32'h42208086, 32'h42425e28, 32'h420d6959, 32'hc28149f2};
test_output[30728:30735] = '{32'h42bc7d26, 32'h0, 32'h0, 32'h400f0d90, 32'h42208086, 32'h42425e28, 32'h420d6959, 32'h0};
test_input[30736:30743] = '{32'h4202ec5e, 32'h42889ef5, 32'hc2354ba8, 32'h429cca78, 32'h421fde1b, 32'h42b5af1e, 32'hc268db35, 32'h40c78589};
test_output[30736:30743] = '{32'h4202ec5e, 32'h42889ef5, 32'h0, 32'h429cca78, 32'h421fde1b, 32'h42b5af1e, 32'h0, 32'h40c78589};
test_input[30744:30751] = '{32'h42c50059, 32'h41877f57, 32'hc1834ae5, 32'h4228022b, 32'h409351e1, 32'hbdf93ea2, 32'h419e7e46, 32'hc1b3b91d};
test_output[30744:30751] = '{32'h42c50059, 32'h41877f57, 32'h0, 32'h4228022b, 32'h409351e1, 32'h0, 32'h419e7e46, 32'h0};
test_input[30752:30759] = '{32'hc0e5a348, 32'hc1abbb3c, 32'hc188bff5, 32'h42c085fb, 32'hc2b9d7cf, 32'hc2a1b7fa, 32'hc1ccc0a7, 32'h42b919a6};
test_output[30752:30759] = '{32'h0, 32'h0, 32'h0, 32'h42c085fb, 32'h0, 32'h0, 32'h0, 32'h42b919a6};
test_input[30760:30767] = '{32'hc25df3f7, 32'h41d69c5d, 32'h4261f44a, 32'h408baab3, 32'h41ad77be, 32'hc2017771, 32'h42b50dd9, 32'h4265bb7e};
test_output[30760:30767] = '{32'h0, 32'h41d69c5d, 32'h4261f44a, 32'h408baab3, 32'h41ad77be, 32'h0, 32'h42b50dd9, 32'h4265bb7e};
test_input[30768:30775] = '{32'hc292face, 32'hc100a997, 32'hc1540ac8, 32'hc29cb26b, 32'hc104e53d, 32'h42c34042, 32'h41cd92db, 32'h42c7c1ff};
test_output[30768:30775] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c34042, 32'h41cd92db, 32'h42c7c1ff};
test_input[30776:30783] = '{32'hc2282813, 32'hc2a0ee6a, 32'hc2160798, 32'hc25add0b, 32'h41b80b8f, 32'hbfad854f, 32'hc23dd1dc, 32'hc2b427d1};
test_output[30776:30783] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41b80b8f, 32'h0, 32'h0, 32'h0};
test_input[30784:30791] = '{32'h41f17440, 32'h42b9248f, 32'hc1af1a74, 32'h423545d5, 32'hc1e9804f, 32'hc1e1c48b, 32'h42127297, 32'hc1c5fbe1};
test_output[30784:30791] = '{32'h41f17440, 32'h42b9248f, 32'h0, 32'h423545d5, 32'h0, 32'h0, 32'h42127297, 32'h0};
test_input[30792:30799] = '{32'hc21ce719, 32'h424af216, 32'hc2885fa0, 32'h428a9931, 32'hc21fca74, 32'h42b0ec22, 32'h4289c8b4, 32'h423a1cc1};
test_output[30792:30799] = '{32'h0, 32'h424af216, 32'h0, 32'h428a9931, 32'h0, 32'h42b0ec22, 32'h4289c8b4, 32'h423a1cc1};
test_input[30800:30807] = '{32'h424fb433, 32'hc28f0821, 32'hc2c010a0, 32'hc2a29564, 32'h420b1bd9, 32'hc297c155, 32'h41d6aa85, 32'h427cb21a};
test_output[30800:30807] = '{32'h424fb433, 32'h0, 32'h0, 32'h0, 32'h420b1bd9, 32'h0, 32'h41d6aa85, 32'h427cb21a};
test_input[30808:30815] = '{32'h41b372af, 32'hc23c5ed4, 32'hc2735e30, 32'hbf4f8e4c, 32'h42856316, 32'h41b16dd3, 32'hc155525c, 32'h42836cd1};
test_output[30808:30815] = '{32'h41b372af, 32'h0, 32'h0, 32'h0, 32'h42856316, 32'h41b16dd3, 32'h0, 32'h42836cd1};
test_input[30816:30823] = '{32'hc2a05204, 32'h420dcfeb, 32'h41054667, 32'h419b1df5, 32'hc22c92b1, 32'h4164bb28, 32'h41c866a5, 32'h41b939dd};
test_output[30816:30823] = '{32'h0, 32'h420dcfeb, 32'h41054667, 32'h419b1df5, 32'h0, 32'h4164bb28, 32'h41c866a5, 32'h41b939dd};
test_input[30824:30831] = '{32'hc1770098, 32'h427aefba, 32'hc096bd1b, 32'hc12eddd2, 32'h4025ce2f, 32'h4181a07a, 32'h42afc9cc, 32'h41cee2b4};
test_output[30824:30831] = '{32'h0, 32'h427aefba, 32'h0, 32'h0, 32'h4025ce2f, 32'h4181a07a, 32'h42afc9cc, 32'h41cee2b4};
test_input[30832:30839] = '{32'hc2490b67, 32'hc2a9c4f2, 32'h427f25bd, 32'h423bc656, 32'hc291aca9, 32'h42aaade7, 32'hc10647ca, 32'h42ba00f8};
test_output[30832:30839] = '{32'h0, 32'h0, 32'h427f25bd, 32'h423bc656, 32'h0, 32'h42aaade7, 32'h0, 32'h42ba00f8};
test_input[30840:30847] = '{32'h419a908d, 32'hc29ba551, 32'hc28a140b, 32'hc190da90, 32'h41ffa136, 32'h4198e68a, 32'h425f54fb, 32'h429c7340};
test_output[30840:30847] = '{32'h419a908d, 32'h0, 32'h0, 32'h0, 32'h41ffa136, 32'h4198e68a, 32'h425f54fb, 32'h429c7340};
test_input[30848:30855] = '{32'h42a4b941, 32'hc2b993a6, 32'hc20acbee, 32'h4286a57b, 32'h420e4369, 32'h4163b2d1, 32'hc295b97c, 32'h41ca014e};
test_output[30848:30855] = '{32'h42a4b941, 32'h0, 32'h0, 32'h4286a57b, 32'h420e4369, 32'h4163b2d1, 32'h0, 32'h41ca014e};
test_input[30856:30863] = '{32'hc2c28e8b, 32'hc1adcb1e, 32'hc2480f79, 32'h41fcbb34, 32'h422a3c83, 32'h427f2a3f, 32'h42bc42e0, 32'hc19cef83};
test_output[30856:30863] = '{32'h0, 32'h0, 32'h0, 32'h41fcbb34, 32'h422a3c83, 32'h427f2a3f, 32'h42bc42e0, 32'h0};
test_input[30864:30871] = '{32'h41ad5717, 32'h429c97bf, 32'hc2925923, 32'hc1726c1b, 32'hc2c7e1e4, 32'hc18813e3, 32'h426266c0, 32'h42883c86};
test_output[30864:30871] = '{32'h41ad5717, 32'h429c97bf, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426266c0, 32'h42883c86};
test_input[30872:30879] = '{32'h424167d1, 32'hc2c790b8, 32'h420113d2, 32'hc16efa8a, 32'h4285b97e, 32'h414dd8d9, 32'hc2754113, 32'h42668e55};
test_output[30872:30879] = '{32'h424167d1, 32'h0, 32'h420113d2, 32'h0, 32'h4285b97e, 32'h414dd8d9, 32'h0, 32'h42668e55};
test_input[30880:30887] = '{32'h403c3f53, 32'h424ffac7, 32'hc28b916e, 32'hc230c82d, 32'h422e2cec, 32'h42b768d7, 32'h426d4ae5, 32'h42a01bb4};
test_output[30880:30887] = '{32'h403c3f53, 32'h424ffac7, 32'h0, 32'h0, 32'h422e2cec, 32'h42b768d7, 32'h426d4ae5, 32'h42a01bb4};
test_input[30888:30895] = '{32'hc201b8a4, 32'h42145452, 32'h40aa929d, 32'h42789978, 32'h42461fa4, 32'h41dfb458, 32'h40c8388f, 32'hc26d4126};
test_output[30888:30895] = '{32'h0, 32'h42145452, 32'h40aa929d, 32'h42789978, 32'h42461fa4, 32'h41dfb458, 32'h40c8388f, 32'h0};
test_input[30896:30903] = '{32'hc2b71def, 32'h3e6e5497, 32'hc1ba573b, 32'hc21fd22d, 32'h420c6137, 32'h42bba0f6, 32'h41d24354, 32'h40525835};
test_output[30896:30903] = '{32'h0, 32'h3e6e5497, 32'h0, 32'h0, 32'h420c6137, 32'h42bba0f6, 32'h41d24354, 32'h40525835};
test_input[30904:30911] = '{32'hbe7169fe, 32'h40bcf3de, 32'h423d06b5, 32'hc2175f2a, 32'hc2b4e708, 32'hc141d933, 32'h418f7f50, 32'hc214cead};
test_output[30904:30911] = '{32'h0, 32'h40bcf3de, 32'h423d06b5, 32'h0, 32'h0, 32'h0, 32'h418f7f50, 32'h0};
test_input[30912:30919] = '{32'h42aa1255, 32'h4105179e, 32'h422964a9, 32'hc258cc44, 32'hc26f51be, 32'hc2889318, 32'hc2158629, 32'h41cb7754};
test_output[30912:30919] = '{32'h42aa1255, 32'h4105179e, 32'h422964a9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41cb7754};
test_input[30920:30927] = '{32'h4200acd9, 32'h42a2858e, 32'hc2304480, 32'h42af6993, 32'hc280dcd1, 32'h429bf26c, 32'h423b6907, 32'h4155d146};
test_output[30920:30927] = '{32'h4200acd9, 32'h42a2858e, 32'h0, 32'h42af6993, 32'h0, 32'h429bf26c, 32'h423b6907, 32'h4155d146};
test_input[30928:30935] = '{32'h4282cc4c, 32'h42b3a68d, 32'h42c06bc4, 32'h42274087, 32'hc180f15a, 32'hc2ad31af, 32'h42b539cd, 32'h42c14883};
test_output[30928:30935] = '{32'h4282cc4c, 32'h42b3a68d, 32'h42c06bc4, 32'h42274087, 32'h0, 32'h0, 32'h42b539cd, 32'h42c14883};
test_input[30936:30943] = '{32'h42216997, 32'hc259838a, 32'h403d4ea6, 32'h413e15ce, 32'h41391a54, 32'h4252ff9b, 32'h42885c63, 32'hc2b395bb};
test_output[30936:30943] = '{32'h42216997, 32'h0, 32'h403d4ea6, 32'h413e15ce, 32'h41391a54, 32'h4252ff9b, 32'h42885c63, 32'h0};
test_input[30944:30951] = '{32'hc0f81715, 32'h41bef3f1, 32'h42571970, 32'hc2bc8d53, 32'h423346a2, 32'h420ff52d, 32'h406f0901, 32'h41cee471};
test_output[30944:30951] = '{32'h0, 32'h41bef3f1, 32'h42571970, 32'h0, 32'h423346a2, 32'h420ff52d, 32'h406f0901, 32'h41cee471};
test_input[30952:30959] = '{32'h424ad20a, 32'h42c70272, 32'hc1ee898a, 32'hc171b7d6, 32'hc1ce5f3f, 32'h42b6b31d, 32'hc26050b9, 32'h41bb8722};
test_output[30952:30959] = '{32'h424ad20a, 32'h42c70272, 32'h0, 32'h0, 32'h0, 32'h42b6b31d, 32'h0, 32'h41bb8722};
test_input[30960:30967] = '{32'h41c4fe89, 32'hc2221c10, 32'hc19084ce, 32'h424267fa, 32'hc2532ac3, 32'h42a9d08b, 32'hc1f05df4, 32'hc29dee4c};
test_output[30960:30967] = '{32'h41c4fe89, 32'h0, 32'h0, 32'h424267fa, 32'h0, 32'h42a9d08b, 32'h0, 32'h0};
test_input[30968:30975] = '{32'h42965edf, 32'hc237c668, 32'hc2c72807, 32'h403e2691, 32'hc282b157, 32'h4282414d, 32'hc2661ba4, 32'h4119d7ea};
test_output[30968:30975] = '{32'h42965edf, 32'h0, 32'h0, 32'h403e2691, 32'h0, 32'h4282414d, 32'h0, 32'h4119d7ea};
test_input[30976:30983] = '{32'h428c9403, 32'hc2a9c8eb, 32'h421ada89, 32'h41a95369, 32'hc2b2cc59, 32'h420695b3, 32'h4101370b, 32'h42867058};
test_output[30976:30983] = '{32'h428c9403, 32'h0, 32'h421ada89, 32'h41a95369, 32'h0, 32'h420695b3, 32'h4101370b, 32'h42867058};
test_input[30984:30991] = '{32'h3f2a07c7, 32'hc220dac0, 32'h40d1c697, 32'hc089f26b, 32'hc280246f, 32'h4246f38b, 32'h42887b6d, 32'h425855ba};
test_output[30984:30991] = '{32'h3f2a07c7, 32'h0, 32'h40d1c697, 32'h0, 32'h0, 32'h4246f38b, 32'h42887b6d, 32'h425855ba};
test_input[30992:30999] = '{32'h40ae1767, 32'h42841191, 32'hc1fa073b, 32'h41d431c8, 32'h42513ce5, 32'h419fe48b, 32'hc1e0d077, 32'h41c5bdc6};
test_output[30992:30999] = '{32'h40ae1767, 32'h42841191, 32'h0, 32'h41d431c8, 32'h42513ce5, 32'h419fe48b, 32'h0, 32'h41c5bdc6};
test_input[31000:31007] = '{32'hc27e10f4, 32'h4273d9a9, 32'h42628771, 32'h41941aaa, 32'h429201ee, 32'hc24e5014, 32'hc246a2f4, 32'h42bf1f25};
test_output[31000:31007] = '{32'h0, 32'h4273d9a9, 32'h42628771, 32'h41941aaa, 32'h429201ee, 32'h0, 32'h0, 32'h42bf1f25};
test_input[31008:31015] = '{32'h419b0c9b, 32'hc21c6dfa, 32'h420e3738, 32'hc275627e, 32'h418df5f8, 32'h42714550, 32'hc111e6a5, 32'hc2391a54};
test_output[31008:31015] = '{32'h419b0c9b, 32'h0, 32'h420e3738, 32'h0, 32'h418df5f8, 32'h42714550, 32'h0, 32'h0};
test_input[31016:31023] = '{32'hc1f103fa, 32'h42833041, 32'hc2b8375a, 32'hc21282e3, 32'h42419f76, 32'hc21c01b7, 32'hc22d41ea, 32'hc1bea5c3};
test_output[31016:31023] = '{32'h0, 32'h42833041, 32'h0, 32'h0, 32'h42419f76, 32'h0, 32'h0, 32'h0};
test_input[31024:31031] = '{32'hc18a903e, 32'h42a6e623, 32'h4296aa90, 32'h42b84e0a, 32'hc2c38ce7, 32'h4210db29, 32'hc2abcd70, 32'hc2608c60};
test_output[31024:31031] = '{32'h0, 32'h42a6e623, 32'h4296aa90, 32'h42b84e0a, 32'h0, 32'h4210db29, 32'h0, 32'h0};
test_input[31032:31039] = '{32'hc177f9dc, 32'hc0dc861f, 32'hc26837fa, 32'hc1922065, 32'h4281b460, 32'hc2999c1a, 32'h40c40c78, 32'hc1efe227};
test_output[31032:31039] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4281b460, 32'h0, 32'h40c40c78, 32'h0};
test_input[31040:31047] = '{32'h41791393, 32'h425333cd, 32'h41a69ff3, 32'hc268ffbc, 32'hc2b46274, 32'hc2658cdf, 32'hc27d9303, 32'h428de765};
test_output[31040:31047] = '{32'h41791393, 32'h425333cd, 32'h41a69ff3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428de765};
test_input[31048:31055] = '{32'h422ba163, 32'hc2531917, 32'h426ea45b, 32'hc2529399, 32'hc0d783ca, 32'hc15388b9, 32'hc2722aed, 32'h428e4572};
test_output[31048:31055] = '{32'h422ba163, 32'h0, 32'h426ea45b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428e4572};
test_input[31056:31063] = '{32'h42a92c1c, 32'hc23a75f9, 32'h40902fd9, 32'hc28605c3, 32'hc16e1256, 32'hc1ace60b, 32'h40a1051e, 32'hc182c383};
test_output[31056:31063] = '{32'h42a92c1c, 32'h0, 32'h40902fd9, 32'h0, 32'h0, 32'h0, 32'h40a1051e, 32'h0};
test_input[31064:31071] = '{32'hc16cd5b0, 32'h41b9f97b, 32'h423a83ae, 32'hc226e03e, 32'h426f50a1, 32'h41f1b052, 32'h428491c9, 32'h41c4f9bd};
test_output[31064:31071] = '{32'h0, 32'h41b9f97b, 32'h423a83ae, 32'h0, 32'h426f50a1, 32'h41f1b052, 32'h428491c9, 32'h41c4f9bd};
test_input[31072:31079] = '{32'hc261da0a, 32'h42803c82, 32'hc26915c0, 32'h40303dfb, 32'h42983478, 32'h4265cd4c, 32'h41e262b5, 32'hc1937ff8};
test_output[31072:31079] = '{32'h0, 32'h42803c82, 32'h0, 32'h40303dfb, 32'h42983478, 32'h4265cd4c, 32'h41e262b5, 32'h0};
test_input[31080:31087] = '{32'hc22dd940, 32'h42bf64d5, 32'hc1e9d718, 32'h417a131e, 32'h42bd76d8, 32'hc1be019d, 32'h42107c78, 32'hc2b3192c};
test_output[31080:31087] = '{32'h0, 32'h42bf64d5, 32'h0, 32'h417a131e, 32'h42bd76d8, 32'h0, 32'h42107c78, 32'h0};
test_input[31088:31095] = '{32'hc2c0f52f, 32'h42897f0f, 32'hc2092de0, 32'hc2aaa109, 32'hc19559a4, 32'h42a1c079, 32'h42b74e87, 32'h421789bb};
test_output[31088:31095] = '{32'h0, 32'h42897f0f, 32'h0, 32'h0, 32'h0, 32'h42a1c079, 32'h42b74e87, 32'h421789bb};
test_input[31096:31103] = '{32'hc1f85026, 32'h42ab3920, 32'h42c0df1a, 32'h411d652b, 32'hc2a2d30c, 32'hc1e817f8, 32'hc28ac006, 32'hc291e546};
test_output[31096:31103] = '{32'h0, 32'h42ab3920, 32'h42c0df1a, 32'h411d652b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31104:31111] = '{32'hc19637b4, 32'h42a275e6, 32'h42a9eddd, 32'h423eddab, 32'hc2b8eccd, 32'hc288490b, 32'h41c4c6d6, 32'hc238f6e4};
test_output[31104:31111] = '{32'h0, 32'h42a275e6, 32'h42a9eddd, 32'h423eddab, 32'h0, 32'h0, 32'h41c4c6d6, 32'h0};
test_input[31112:31119] = '{32'h42bf0684, 32'hc1963654, 32'hc26c6240, 32'h4287c206, 32'hc25bd4a2, 32'hc28c5c3f, 32'h424ad549, 32'hc1c6cde0};
test_output[31112:31119] = '{32'h42bf0684, 32'h0, 32'h0, 32'h4287c206, 32'h0, 32'h0, 32'h424ad549, 32'h0};
test_input[31120:31127] = '{32'h42b55080, 32'h42b28558, 32'h429b916c, 32'hc21976f0, 32'hc23a9b04, 32'hc1cb2e35, 32'h41b77d90, 32'hc2127fb1};
test_output[31120:31127] = '{32'h42b55080, 32'h42b28558, 32'h429b916c, 32'h0, 32'h0, 32'h0, 32'h41b77d90, 32'h0};
test_input[31128:31135] = '{32'hc1e849c7, 32'h42b2ba50, 32'h4222ad9f, 32'h41a334d4, 32'hc0f45f26, 32'hc2bfb2f5, 32'h41938823, 32'hc29dac70};
test_output[31128:31135] = '{32'h0, 32'h42b2ba50, 32'h4222ad9f, 32'h41a334d4, 32'h0, 32'h0, 32'h41938823, 32'h0};
test_input[31136:31143] = '{32'hc28fcaf4, 32'hc282bb9f, 32'hc29b3662, 32'h3fb8f689, 32'h429a8ef6, 32'h4286e012, 32'hc2620052, 32'h414e13a1};
test_output[31136:31143] = '{32'h0, 32'h0, 32'h0, 32'h3fb8f689, 32'h429a8ef6, 32'h4286e012, 32'h0, 32'h414e13a1};
test_input[31144:31151] = '{32'h42342ad6, 32'h4293db22, 32'hbf62fe66, 32'h42bcce7e, 32'hc1a9f30f, 32'hc24b75e5, 32'hc174d472, 32'h42092860};
test_output[31144:31151] = '{32'h42342ad6, 32'h4293db22, 32'h0, 32'h42bcce7e, 32'h0, 32'h0, 32'h0, 32'h42092860};
test_input[31152:31159] = '{32'hc1e3fec9, 32'hc21c1ffa, 32'h412b6e62, 32'hc13fd8fd, 32'h42bc9b5e, 32'h422816ac, 32'h425a302b, 32'h429b8eda};
test_output[31152:31159] = '{32'h0, 32'h0, 32'h412b6e62, 32'h0, 32'h42bc9b5e, 32'h422816ac, 32'h425a302b, 32'h429b8eda};
test_input[31160:31167] = '{32'h423845d5, 32'h426fd945, 32'h4272a686, 32'hc2817a94, 32'h42c08043, 32'h42a9d1e0, 32'hc0a780c2, 32'h424ff8c4};
test_output[31160:31167] = '{32'h423845d5, 32'h426fd945, 32'h4272a686, 32'h0, 32'h42c08043, 32'h42a9d1e0, 32'h0, 32'h424ff8c4};
test_input[31168:31175] = '{32'h42b8688c, 32'hc18f595e, 32'h4257b3c5, 32'hc0197532, 32'h4150d65f, 32'h419eb5c3, 32'h422503bf, 32'hc25e8402};
test_output[31168:31175] = '{32'h42b8688c, 32'h0, 32'h4257b3c5, 32'h0, 32'h4150d65f, 32'h419eb5c3, 32'h422503bf, 32'h0};
test_input[31176:31183] = '{32'h42529db4, 32'h41af24e0, 32'h4222756b, 32'hc2b5b100, 32'hc2025966, 32'hc2a89665, 32'h42b0e939, 32'h42394f09};
test_output[31176:31183] = '{32'h42529db4, 32'h41af24e0, 32'h4222756b, 32'h0, 32'h0, 32'h0, 32'h42b0e939, 32'h42394f09};
test_input[31184:31191] = '{32'hc2bb1e3f, 32'hc27ece52, 32'h42c741ae, 32'hc1e23a82, 32'h426ef06f, 32'hc1e566b1, 32'hc187b92e, 32'hc2a0c9c6};
test_output[31184:31191] = '{32'h0, 32'h0, 32'h42c741ae, 32'h0, 32'h426ef06f, 32'h0, 32'h0, 32'h0};
test_input[31192:31199] = '{32'h4208b178, 32'hc1dbbcbc, 32'hc2308520, 32'hc0a8e1b0, 32'h423cc4c0, 32'hbf0d9319, 32'hc2762e68, 32'h4287ad53};
test_output[31192:31199] = '{32'h4208b178, 32'h0, 32'h0, 32'h0, 32'h423cc4c0, 32'h0, 32'h0, 32'h4287ad53};
test_input[31200:31207] = '{32'hc2c2c755, 32'hc16afca2, 32'hc2b0fe1d, 32'hc2743a60, 32'h429e8d74, 32'h42c76288, 32'hc2b40d56, 32'hc220d947};
test_output[31200:31207] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429e8d74, 32'h42c76288, 32'h0, 32'h0};
test_input[31208:31215] = '{32'h40c810ff, 32'hc1055a4c, 32'h42aa5e87, 32'h42532d77, 32'hc11f8e38, 32'hc2a966b9, 32'h429edf02, 32'h42ae467f};
test_output[31208:31215] = '{32'h40c810ff, 32'h0, 32'h42aa5e87, 32'h42532d77, 32'h0, 32'h0, 32'h429edf02, 32'h42ae467f};
test_input[31216:31223] = '{32'hc222ebb8, 32'hc296e2b5, 32'hc23783c0, 32'h418a944f, 32'hc2acc7f3, 32'hc1a9d8f0, 32'h4178588e, 32'hc292a1fe};
test_output[31216:31223] = '{32'h0, 32'h0, 32'h0, 32'h418a944f, 32'h0, 32'h0, 32'h4178588e, 32'h0};
test_input[31224:31231] = '{32'h42a50155, 32'hc0e05658, 32'h421a0c91, 32'hc1c60935, 32'h422c12c1, 32'hc2a608f1, 32'hc2858e0c, 32'h4213ca55};
test_output[31224:31231] = '{32'h42a50155, 32'h0, 32'h421a0c91, 32'h0, 32'h422c12c1, 32'h0, 32'h0, 32'h4213ca55};
test_input[31232:31239] = '{32'h42b0983c, 32'h42c74239, 32'hc2096129, 32'h424987d9, 32'h4262fe64, 32'h428fea84, 32'hc0d51ba8, 32'h420db03d};
test_output[31232:31239] = '{32'h42b0983c, 32'h42c74239, 32'h0, 32'h424987d9, 32'h4262fe64, 32'h428fea84, 32'h0, 32'h420db03d};
test_input[31240:31247] = '{32'hc2007d0a, 32'h425c968f, 32'h41c4c395, 32'hc21fd4b5, 32'h424e5e1b, 32'hc18ce9c7, 32'hc290e140, 32'hc2659306};
test_output[31240:31247] = '{32'h0, 32'h425c968f, 32'h41c4c395, 32'h0, 32'h424e5e1b, 32'h0, 32'h0, 32'h0};
test_input[31248:31255] = '{32'hc1f74a22, 32'h4183cb9d, 32'hc180f034, 32'hc28aa142, 32'h42459c9e, 32'h4280a115, 32'h422196ff, 32'hc2250aea};
test_output[31248:31255] = '{32'h0, 32'h4183cb9d, 32'h0, 32'h0, 32'h42459c9e, 32'h4280a115, 32'h422196ff, 32'h0};
test_input[31256:31263] = '{32'hc1244a6d, 32'hc1d2ac78, 32'hc2a6a84e, 32'h42c47b05, 32'h419fbaa1, 32'h429e1069, 32'hc20ded3d, 32'hc29bff39};
test_output[31256:31263] = '{32'h0, 32'h0, 32'h0, 32'h42c47b05, 32'h419fbaa1, 32'h429e1069, 32'h0, 32'h0};
test_input[31264:31271] = '{32'hc19bdb90, 32'hc22c13a8, 32'hc2aa3324, 32'hc2865c1f, 32'hc2a173d7, 32'hc260c4fd, 32'h42c06771, 32'h41eb5d33};
test_output[31264:31271] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c06771, 32'h41eb5d33};
test_input[31272:31279] = '{32'h421a54da, 32'h42791a51, 32'hc265da19, 32'hc28d777b, 32'hc2390209, 32'hc2c380ad, 32'hc11c2c4f, 32'h429b8d52};
test_output[31272:31279] = '{32'h421a54da, 32'h42791a51, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429b8d52};
test_input[31280:31287] = '{32'h4288eab1, 32'h423d7046, 32'h42892e6c, 32'h429b9c01, 32'hc25496d5, 32'h41f13a5c, 32'hc2771a67, 32'hc1256869};
test_output[31280:31287] = '{32'h4288eab1, 32'h423d7046, 32'h42892e6c, 32'h429b9c01, 32'h0, 32'h41f13a5c, 32'h0, 32'h0};
test_input[31288:31295] = '{32'hc2a3b245, 32'h424fd054, 32'hc2052dd7, 32'h41a1102a, 32'h4274f42a, 32'hc2a9a890, 32'h42755512, 32'h41776aa4};
test_output[31288:31295] = '{32'h0, 32'h424fd054, 32'h0, 32'h41a1102a, 32'h4274f42a, 32'h0, 32'h42755512, 32'h41776aa4};
test_input[31296:31303] = '{32'h428f7ba1, 32'hc1d303f8, 32'h41324f1c, 32'h41a53131, 32'hc26da1d0, 32'h42b8d997, 32'hc249421b, 32'h4126dbd2};
test_output[31296:31303] = '{32'h428f7ba1, 32'h0, 32'h41324f1c, 32'h41a53131, 32'h0, 32'h42b8d997, 32'h0, 32'h4126dbd2};
test_input[31304:31311] = '{32'h4146675f, 32'hc1c0d39b, 32'h4296d552, 32'h4235a67b, 32'hc1155c15, 32'h42a1d46e, 32'h42626262, 32'h4112069a};
test_output[31304:31311] = '{32'h4146675f, 32'h0, 32'h4296d552, 32'h4235a67b, 32'h0, 32'h42a1d46e, 32'h42626262, 32'h4112069a};
test_input[31312:31319] = '{32'hc2bfa2b6, 32'h42abe46b, 32'h42a37bad, 32'h422ce75b, 32'hc1bb29bf, 32'hc22914dc, 32'hc1c260a7, 32'h40947b22};
test_output[31312:31319] = '{32'h0, 32'h42abe46b, 32'h42a37bad, 32'h422ce75b, 32'h0, 32'h0, 32'h0, 32'h40947b22};
test_input[31320:31327] = '{32'h4282c396, 32'hc26372d9, 32'h4282f474, 32'hc2360694, 32'h42c1f025, 32'hc299e4b7, 32'h4135b9fb, 32'h422d9a64};
test_output[31320:31327] = '{32'h4282c396, 32'h0, 32'h4282f474, 32'h0, 32'h42c1f025, 32'h0, 32'h4135b9fb, 32'h422d9a64};
test_input[31328:31335] = '{32'hc1804c95, 32'hc19c7532, 32'hc2c11780, 32'hc225aa8e, 32'h41d0c0c6, 32'hc29e6f83, 32'hc28690bb, 32'hc1d73d62};
test_output[31328:31335] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41d0c0c6, 32'h0, 32'h0, 32'h0};
test_input[31336:31343] = '{32'h426544e5, 32'h41f0d2d3, 32'h3fc88223, 32'hc2863348, 32'h420c3aea, 32'h41dc0dfd, 32'hc2246c8f, 32'hc1f9c284};
test_output[31336:31343] = '{32'h426544e5, 32'h41f0d2d3, 32'h3fc88223, 32'h0, 32'h420c3aea, 32'h41dc0dfd, 32'h0, 32'h0};
test_input[31344:31351] = '{32'hc167daae, 32'h429209fb, 32'hc19c6177, 32'h41c6be30, 32'hc1ad377e, 32'h426e9692, 32'hc28dec3c, 32'h414c25be};
test_output[31344:31351] = '{32'h0, 32'h429209fb, 32'h0, 32'h41c6be30, 32'h0, 32'h426e9692, 32'h0, 32'h414c25be};
test_input[31352:31359] = '{32'hc27d1231, 32'hc21bef3f, 32'hc2323e68, 32'hc22e9233, 32'hc1651382, 32'h4299d319, 32'hc2c51a03, 32'hc22b87de};
test_output[31352:31359] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4299d319, 32'h0, 32'h0};
test_input[31360:31367] = '{32'hc19dd88f, 32'hc28a7ca1, 32'hc24c934e, 32'hc283b751, 32'hc027e413, 32'hc2a843dd, 32'hc28dd83e, 32'hc2badd6c};
test_output[31360:31367] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31368:31375] = '{32'hc2aa8aae, 32'h42a17536, 32'h429c1178, 32'hc06b6db3, 32'h4284d182, 32'h41b90eba, 32'hc0f1d04c, 32'hc27f6c8e};
test_output[31368:31375] = '{32'h0, 32'h42a17536, 32'h429c1178, 32'h0, 32'h4284d182, 32'h41b90eba, 32'h0, 32'h0};
test_input[31376:31383] = '{32'hc2287ce1, 32'h4281559f, 32'hc2a5340c, 32'h42c653bc, 32'h428f2f9a, 32'h42a09bf4, 32'h400e781a, 32'h42c39585};
test_output[31376:31383] = '{32'h0, 32'h4281559f, 32'h0, 32'h42c653bc, 32'h428f2f9a, 32'h42a09bf4, 32'h400e781a, 32'h42c39585};
test_input[31384:31391] = '{32'h41853a4f, 32'h41e27b1b, 32'hc1e525a6, 32'h40a39f35, 32'hc28b1c63, 32'hc28a9cf4, 32'hc2172960, 32'hc2935193};
test_output[31384:31391] = '{32'h41853a4f, 32'h41e27b1b, 32'h0, 32'h40a39f35, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31392:31399] = '{32'hc29c0f17, 32'h42824ce8, 32'h42ac92d0, 32'hc2367303, 32'h42c0a582, 32'h42737087, 32'h4269e385, 32'h41e961c0};
test_output[31392:31399] = '{32'h0, 32'h42824ce8, 32'h42ac92d0, 32'h0, 32'h42c0a582, 32'h42737087, 32'h4269e385, 32'h41e961c0};
test_input[31400:31407] = '{32'hc28a25b2, 32'hc2831f37, 32'h42771ed0, 32'hc1596464, 32'hc2b25e89, 32'h424d0bf6, 32'hc2c11c0f, 32'hbf7971e6};
test_output[31400:31407] = '{32'h0, 32'h0, 32'h42771ed0, 32'h0, 32'h0, 32'h424d0bf6, 32'h0, 32'h0};
test_input[31408:31415] = '{32'h42aebd07, 32'h42083079, 32'h4207d016, 32'h426f051b, 32'h4257a0ea, 32'h420c8e1b, 32'h419dbfc3, 32'h42b92bff};
test_output[31408:31415] = '{32'h42aebd07, 32'h42083079, 32'h4207d016, 32'h426f051b, 32'h4257a0ea, 32'h420c8e1b, 32'h419dbfc3, 32'h42b92bff};
test_input[31416:31423] = '{32'h423d20cb, 32'hc281f2fd, 32'hc05ccaea, 32'hc11c274b, 32'hc28d3879, 32'hc23349a6, 32'h42b72d1d, 32'h424ef5b9};
test_output[31416:31423] = '{32'h423d20cb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b72d1d, 32'h424ef5b9};
test_input[31424:31431] = '{32'hc2c08616, 32'hc10fc8bd, 32'hc0e170aa, 32'h42b1088f, 32'h42b8a0a1, 32'h42c70bf7, 32'h429623a1, 32'h41707071};
test_output[31424:31431] = '{32'h0, 32'h0, 32'h0, 32'h42b1088f, 32'h42b8a0a1, 32'h42c70bf7, 32'h429623a1, 32'h41707071};
test_input[31432:31439] = '{32'hc28b3dd8, 32'h42910cb0, 32'hc134a59d, 32'h41d83774, 32'hc28881bc, 32'h42b6a132, 32'hc249c5f4, 32'h42bc571a};
test_output[31432:31439] = '{32'h0, 32'h42910cb0, 32'h0, 32'h41d83774, 32'h0, 32'h42b6a132, 32'h0, 32'h42bc571a};
test_input[31440:31447] = '{32'h42b7af5f, 32'hc20bb62c, 32'h4071b29d, 32'h41926990, 32'hbfdb7231, 32'h42af514e, 32'h425ff379, 32'hc10878b7};
test_output[31440:31447] = '{32'h42b7af5f, 32'h0, 32'h4071b29d, 32'h41926990, 32'h0, 32'h42af514e, 32'h425ff379, 32'h0};
test_input[31448:31455] = '{32'h42201ee8, 32'h42234b7b, 32'h41c796f9, 32'h406ff389, 32'hc23840de, 32'hc1b93ede, 32'hc2a785a2, 32'hc1edbe5c};
test_output[31448:31455] = '{32'h42201ee8, 32'h42234b7b, 32'h41c796f9, 32'h406ff389, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31456:31463] = '{32'hc25bd0c6, 32'h42835e26, 32'hc28d9300, 32'h42c44ef1, 32'h42c221be, 32'hc28aee18, 32'h4213a372, 32'h42abea5d};
test_output[31456:31463] = '{32'h0, 32'h42835e26, 32'h0, 32'h42c44ef1, 32'h42c221be, 32'h0, 32'h4213a372, 32'h42abea5d};
test_input[31464:31471] = '{32'h42544d79, 32'hc18cdf58, 32'h40a278b0, 32'hc21481c6, 32'hc296e868, 32'hc284a683, 32'h423f93bb, 32'h427ac554};
test_output[31464:31471] = '{32'h42544d79, 32'h0, 32'h40a278b0, 32'h0, 32'h0, 32'h0, 32'h423f93bb, 32'h427ac554};
test_input[31472:31479] = '{32'h4256ed70, 32'hc0b55c8e, 32'h4230e0e2, 32'h4179279d, 32'hc23109f0, 32'h4271e627, 32'hc2b3dd9e, 32'h42b1d0ea};
test_output[31472:31479] = '{32'h4256ed70, 32'h0, 32'h4230e0e2, 32'h4179279d, 32'h0, 32'h4271e627, 32'h0, 32'h42b1d0ea};
test_input[31480:31487] = '{32'h429cecc1, 32'h41674c30, 32'h42b2c074, 32'h427280dc, 32'hc1bbb36b, 32'h410f0574, 32'hc2443a34, 32'h42a010b7};
test_output[31480:31487] = '{32'h429cecc1, 32'h41674c30, 32'h42b2c074, 32'h427280dc, 32'h0, 32'h410f0574, 32'h0, 32'h42a010b7};
test_input[31488:31495] = '{32'hc22769a2, 32'h42a21f6d, 32'h427797f9, 32'hc2170e3d, 32'h428b0202, 32'h4209f674, 32'h41689703, 32'hc288eb52};
test_output[31488:31495] = '{32'h0, 32'h42a21f6d, 32'h427797f9, 32'h0, 32'h428b0202, 32'h4209f674, 32'h41689703, 32'h0};
test_input[31496:31503] = '{32'h41602bc5, 32'hc298c3c6, 32'h4293f2f2, 32'hc21c403f, 32'h42c5a1bc, 32'h4282e708, 32'h41eb0697, 32'hc2313ebd};
test_output[31496:31503] = '{32'h41602bc5, 32'h0, 32'h4293f2f2, 32'h0, 32'h42c5a1bc, 32'h4282e708, 32'h41eb0697, 32'h0};
test_input[31504:31511] = '{32'h42bf8450, 32'h421fa16f, 32'hc2904a8d, 32'h42b7ba4f, 32'hc2bde409, 32'hc21f61eb, 32'hc2a6fd58, 32'h41b9d12b};
test_output[31504:31511] = '{32'h42bf8450, 32'h421fa16f, 32'h0, 32'h42b7ba4f, 32'h0, 32'h0, 32'h0, 32'h41b9d12b};
test_input[31512:31519] = '{32'hc2b902cb, 32'hc23e1a94, 32'h42542ef0, 32'hc1a8abd1, 32'hc1cad62f, 32'hc2300c03, 32'h421ab13b, 32'h42225abb};
test_output[31512:31519] = '{32'h0, 32'h0, 32'h42542ef0, 32'h0, 32'h0, 32'h0, 32'h421ab13b, 32'h42225abb};
test_input[31520:31527] = '{32'hc069815c, 32'hc2a1f838, 32'hc2920beb, 32'hc2381b67, 32'hc10d19cc, 32'h41b21894, 32'h4211b568, 32'hc1d9fad6};
test_output[31520:31527] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b21894, 32'h4211b568, 32'h0};
test_input[31528:31535] = '{32'hc221065f, 32'hc1f08473, 32'h42051c7a, 32'h425d3598, 32'hc1a8e592, 32'h42b9f318, 32'hc2b242c3, 32'h4205abbd};
test_output[31528:31535] = '{32'h0, 32'h0, 32'h42051c7a, 32'h425d3598, 32'h0, 32'h42b9f318, 32'h0, 32'h4205abbd};
test_input[31536:31543] = '{32'h424c8070, 32'h41c2ca22, 32'h42ae5583, 32'hc1daff48, 32'h42844736, 32'h42336e11, 32'hc280eee1, 32'hc2712f6d};
test_output[31536:31543] = '{32'h424c8070, 32'h41c2ca22, 32'h42ae5583, 32'h0, 32'h42844736, 32'h42336e11, 32'h0, 32'h0};
test_input[31544:31551] = '{32'hc2541c03, 32'h42a8bb4f, 32'h41b50a11, 32'h41a1b320, 32'h42320fa9, 32'h41cea484, 32'hc1b20044, 32'h4213f602};
test_output[31544:31551] = '{32'h0, 32'h42a8bb4f, 32'h41b50a11, 32'h41a1b320, 32'h42320fa9, 32'h41cea484, 32'h0, 32'h4213f602};
test_input[31552:31559] = '{32'hc2c634a8, 32'hc02aadbc, 32'hc2913206, 32'h4285947f, 32'h42afc726, 32'hc19d6bf0, 32'h426e4dd4, 32'hc163964b};
test_output[31552:31559] = '{32'h0, 32'h0, 32'h0, 32'h4285947f, 32'h42afc726, 32'h0, 32'h426e4dd4, 32'h0};
test_input[31560:31567] = '{32'h419edd5e, 32'h426c6b5d, 32'h4282cf4c, 32'h41e6d67b, 32'hc08b061e, 32'hc230cdbd, 32'hc0cdc9a8, 32'hc170082c};
test_output[31560:31567] = '{32'h419edd5e, 32'h426c6b5d, 32'h4282cf4c, 32'h41e6d67b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31568:31575] = '{32'h41938255, 32'h4288112a, 32'h41b62655, 32'h422cf560, 32'h422ed059, 32'h429910b5, 32'h42c5cd94, 32'h4196873b};
test_output[31568:31575] = '{32'h41938255, 32'h4288112a, 32'h41b62655, 32'h422cf560, 32'h422ed059, 32'h429910b5, 32'h42c5cd94, 32'h4196873b};
test_input[31576:31583] = '{32'h4264b2f1, 32'h42c70114, 32'h427223ba, 32'h42c172a9, 32'hc28c1753, 32'hc23f4549, 32'hc2803a46, 32'hc2c7af2d};
test_output[31576:31583] = '{32'h4264b2f1, 32'h42c70114, 32'h427223ba, 32'h42c172a9, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31584:31591] = '{32'h42c13eea, 32'h41cd038e, 32'h429e9792, 32'hc152f7c6, 32'h423773f3, 32'hc0a0f370, 32'hc22d2ec9, 32'h425f9c41};
test_output[31584:31591] = '{32'h42c13eea, 32'h41cd038e, 32'h429e9792, 32'h0, 32'h423773f3, 32'h0, 32'h0, 32'h425f9c41};
test_input[31592:31599] = '{32'hc0f56311, 32'h4254b52d, 32'h4288a222, 32'h4295bed2, 32'h42c2fb84, 32'hc1750e99, 32'hc25347b3, 32'h424d1ec5};
test_output[31592:31599] = '{32'h0, 32'h4254b52d, 32'h4288a222, 32'h4295bed2, 32'h42c2fb84, 32'h0, 32'h0, 32'h424d1ec5};
test_input[31600:31607] = '{32'h41b0f683, 32'h42832582, 32'h4274f05d, 32'hc2b356d2, 32'h428b20c8, 32'h4297d38a, 32'hc2048249, 32'hc1215062};
test_output[31600:31607] = '{32'h41b0f683, 32'h42832582, 32'h4274f05d, 32'h0, 32'h428b20c8, 32'h4297d38a, 32'h0, 32'h0};
test_input[31608:31615] = '{32'hc287fefb, 32'h42bfd4eb, 32'hc1d0b809, 32'hc2ab11c2, 32'hc2bc9fc2, 32'hbf89a358, 32'h42b79a93, 32'h4216c130};
test_output[31608:31615] = '{32'h0, 32'h42bfd4eb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b79a93, 32'h4216c130};
test_input[31616:31623] = '{32'h42a1309c, 32'hc180c661, 32'h4178e5aa, 32'h42b1fe32, 32'hc2a5f764, 32'hc26c337d, 32'h41196d60, 32'h42384764};
test_output[31616:31623] = '{32'h42a1309c, 32'h0, 32'h4178e5aa, 32'h42b1fe32, 32'h0, 32'h0, 32'h41196d60, 32'h42384764};
test_input[31624:31631] = '{32'h4041430f, 32'hc2c39f44, 32'hc250f6d9, 32'h41bea768, 32'h4218b4b4, 32'hc29400e1, 32'hc2189d79, 32'h42620a0a};
test_output[31624:31631] = '{32'h4041430f, 32'h0, 32'h0, 32'h41bea768, 32'h4218b4b4, 32'h0, 32'h0, 32'h42620a0a};
test_input[31632:31639] = '{32'h418eb18c, 32'hc29d86b0, 32'hc14e81f6, 32'h425481d2, 32'hbed6a179, 32'hc204d47f, 32'h4141b7f9, 32'h414020d9};
test_output[31632:31639] = '{32'h418eb18c, 32'h0, 32'h0, 32'h425481d2, 32'h0, 32'h0, 32'h4141b7f9, 32'h414020d9};
test_input[31640:31647] = '{32'hc1b5e36a, 32'h416156de, 32'h42ab47a4, 32'hc26e834c, 32'hc29c12f9, 32'h42c3738e, 32'h42922052, 32'h42b31d3f};
test_output[31640:31647] = '{32'h0, 32'h416156de, 32'h42ab47a4, 32'h0, 32'h0, 32'h42c3738e, 32'h42922052, 32'h42b31d3f};
test_input[31648:31655] = '{32'h429c97ed, 32'h421b4544, 32'h428385ad, 32'h42af70a2, 32'h425b4989, 32'hc1cf8478, 32'hc2584e2e, 32'h41cad857};
test_output[31648:31655] = '{32'h429c97ed, 32'h421b4544, 32'h428385ad, 32'h42af70a2, 32'h425b4989, 32'h0, 32'h0, 32'h41cad857};
test_input[31656:31663] = '{32'hc229b6db, 32'h4233e450, 32'h42aefab1, 32'h42c08d53, 32'h42929ee9, 32'hc1d23e11, 32'h428c0ef9, 32'hc2947211};
test_output[31656:31663] = '{32'h0, 32'h4233e450, 32'h42aefab1, 32'h42c08d53, 32'h42929ee9, 32'h0, 32'h428c0ef9, 32'h0};
test_input[31664:31671] = '{32'hc2242373, 32'h42b8e204, 32'hc292d90d, 32'h428c9dd3, 32'hc21aa334, 32'hc2b89ffe, 32'h41f02a53, 32'h42b92b6a};
test_output[31664:31671] = '{32'h0, 32'h42b8e204, 32'h0, 32'h428c9dd3, 32'h0, 32'h0, 32'h41f02a53, 32'h42b92b6a};
test_input[31672:31679] = '{32'h42a91e1a, 32'h419b2e86, 32'h429bb775, 32'h426ef5ab, 32'hbf0c62d0, 32'hc1b0fc2e, 32'hc0dd3672, 32'h42a15024};
test_output[31672:31679] = '{32'h42a91e1a, 32'h419b2e86, 32'h429bb775, 32'h426ef5ab, 32'h0, 32'h0, 32'h0, 32'h42a15024};
test_input[31680:31687] = '{32'h408c523f, 32'hc20da098, 32'h42b39b06, 32'hc23398d7, 32'h41a725b1, 32'hc1ba67fa, 32'h42a55572, 32'h42bc201b};
test_output[31680:31687] = '{32'h408c523f, 32'h0, 32'h42b39b06, 32'h0, 32'h41a725b1, 32'h0, 32'h42a55572, 32'h42bc201b};
test_input[31688:31695] = '{32'h41f9f629, 32'h42564859, 32'h42b077e7, 32'hc25ecdf9, 32'h42be0d33, 32'hc213b78f, 32'h4293788c, 32'h425d34c4};
test_output[31688:31695] = '{32'h41f9f629, 32'h42564859, 32'h42b077e7, 32'h0, 32'h42be0d33, 32'h0, 32'h4293788c, 32'h425d34c4};
test_input[31696:31703] = '{32'h415fb143, 32'hc1973275, 32'hc2a2f849, 32'h425be77e, 32'h42976180, 32'hc1a5aca8, 32'hc23c15d0, 32'hc25467d6};
test_output[31696:31703] = '{32'h415fb143, 32'h0, 32'h0, 32'h425be77e, 32'h42976180, 32'h0, 32'h0, 32'h0};
test_input[31704:31711] = '{32'h4284178a, 32'hc282a0d1, 32'hc2bfc579, 32'hc24eff24, 32'hc1274db0, 32'h4209e612, 32'hc1919d7d, 32'h4263c429};
test_output[31704:31711] = '{32'h4284178a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4209e612, 32'h0, 32'h4263c429};
test_input[31712:31719] = '{32'hc1a30fcc, 32'h4060da69, 32'hc1971e71, 32'hc2a26133, 32'h422cec80, 32'hc2c26c97, 32'hc2541d02, 32'hc10a96fb};
test_output[31712:31719] = '{32'h0, 32'h4060da69, 32'h0, 32'h0, 32'h422cec80, 32'h0, 32'h0, 32'h0};
test_input[31720:31727] = '{32'hc243f331, 32'hc226f221, 32'hc2a59012, 32'h40996a6c, 32'h41edd270, 32'h3fcbce4d, 32'hc21f33b1, 32'hc2422c61};
test_output[31720:31727] = '{32'h0, 32'h0, 32'h0, 32'h40996a6c, 32'h41edd270, 32'h3fcbce4d, 32'h0, 32'h0};
test_input[31728:31735] = '{32'h42a9984b, 32'hbfcb2de6, 32'h428969e1, 32'h42a45bfd, 32'h42a9e55b, 32'hc2b3c671, 32'h421a29e8, 32'hc20e6848};
test_output[31728:31735] = '{32'h42a9984b, 32'h0, 32'h428969e1, 32'h42a45bfd, 32'h42a9e55b, 32'h0, 32'h421a29e8, 32'h0};
test_input[31736:31743] = '{32'h42931593, 32'h418707d6, 32'hc2873212, 32'hc2ab1bd1, 32'h42bde830, 32'h42c04bd5, 32'hc25e9ab0, 32'h42bf2352};
test_output[31736:31743] = '{32'h42931593, 32'h418707d6, 32'h0, 32'h0, 32'h42bde830, 32'h42c04bd5, 32'h0, 32'h42bf2352};
test_input[31744:31751] = '{32'h4286c13c, 32'hc1af186d, 32'h428d1478, 32'h418c0a1c, 32'hc2878f5c, 32'hc28ec323, 32'h42868f41, 32'hc2b40e80};
test_output[31744:31751] = '{32'h4286c13c, 32'h0, 32'h428d1478, 32'h418c0a1c, 32'h0, 32'h0, 32'h42868f41, 32'h0};
test_input[31752:31759] = '{32'hc204303c, 32'h40f5a3cd, 32'hc0d983c6, 32'h429d99e2, 32'hc2a4dc17, 32'hc29fd086, 32'h42a4f3de, 32'hc272841c};
test_output[31752:31759] = '{32'h0, 32'h40f5a3cd, 32'h0, 32'h429d99e2, 32'h0, 32'h0, 32'h42a4f3de, 32'h0};
test_input[31760:31767] = '{32'h419bcdf7, 32'hc26eb716, 32'h41440a40, 32'hc27c7277, 32'hc29bd3c3, 32'h3f95a391, 32'h42c43e99, 32'hc1bad82e};
test_output[31760:31767] = '{32'h419bcdf7, 32'h0, 32'h41440a40, 32'h0, 32'h0, 32'h3f95a391, 32'h42c43e99, 32'h0};
test_input[31768:31775] = '{32'h427ca0cb, 32'hc1b94d61, 32'h403c60e2, 32'h42ac771c, 32'h42367f99, 32'h42b5d589, 32'hc2a76fda, 32'hc2818b4b};
test_output[31768:31775] = '{32'h427ca0cb, 32'h0, 32'h403c60e2, 32'h42ac771c, 32'h42367f99, 32'h42b5d589, 32'h0, 32'h0};
test_input[31776:31783] = '{32'hc2947dbf, 32'h425444c3, 32'hc284912d, 32'h40395d12, 32'h429cf91f, 32'hc1badb50, 32'h419f35ad, 32'hc1f55012};
test_output[31776:31783] = '{32'h0, 32'h425444c3, 32'h0, 32'h40395d12, 32'h429cf91f, 32'h0, 32'h419f35ad, 32'h0};
test_input[31784:31791] = '{32'hc1de827f, 32'hc2572462, 32'hc297308e, 32'h418e5c41, 32'h418e37cf, 32'h41d0f545, 32'hc134b7ce, 32'h425ab92a};
test_output[31784:31791] = '{32'h0, 32'h0, 32'h0, 32'h418e5c41, 32'h418e37cf, 32'h41d0f545, 32'h0, 32'h425ab92a};
test_input[31792:31799] = '{32'h41edfd98, 32'h41599e5f, 32'hc231fdfc, 32'h42983f74, 32'h41e7e7e4, 32'hc2a68599, 32'h42187f7d, 32'h42b9ef19};
test_output[31792:31799] = '{32'h41edfd98, 32'h41599e5f, 32'h0, 32'h42983f74, 32'h41e7e7e4, 32'h0, 32'h42187f7d, 32'h42b9ef19};
test_input[31800:31807] = '{32'h41d6bf58, 32'h4296eee8, 32'hc2aeca90, 32'hc2ad2045, 32'hc02fabb3, 32'hc10cbd8c, 32'hc2ab9c78, 32'hc20cc854};
test_output[31800:31807] = '{32'h41d6bf58, 32'h4296eee8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31808:31815] = '{32'hc1ebeddb, 32'hc23af164, 32'h42b1bbda, 32'h425ef7b7, 32'hc26913e4, 32'hc254b00a, 32'h41e4f6ad, 32'h418d0937};
test_output[31808:31815] = '{32'h0, 32'h0, 32'h42b1bbda, 32'h425ef7b7, 32'h0, 32'h0, 32'h41e4f6ad, 32'h418d0937};
test_input[31816:31823] = '{32'hc186df0a, 32'h428b69a7, 32'hc235ada4, 32'h41e26ce8, 32'h42a8dff7, 32'hbf624e75, 32'h415e9223, 32'hc2999e88};
test_output[31816:31823] = '{32'h0, 32'h428b69a7, 32'h0, 32'h41e26ce8, 32'h42a8dff7, 32'h0, 32'h415e9223, 32'h0};
test_input[31824:31831] = '{32'h4246bdaf, 32'h421c99c5, 32'hc26cb9ab, 32'hc28ae426, 32'h424f4b5c, 32'hc2a110a6, 32'hc134abfd, 32'h421029c5};
test_output[31824:31831] = '{32'h4246bdaf, 32'h421c99c5, 32'h0, 32'h0, 32'h424f4b5c, 32'h0, 32'h0, 32'h421029c5};
test_input[31832:31839] = '{32'hc225d3c5, 32'hc2bef45e, 32'hc29b0ea6, 32'h42ad195d, 32'hc1ebd7e6, 32'h42971ab4, 32'h427e4787, 32'h42679706};
test_output[31832:31839] = '{32'h0, 32'h0, 32'h0, 32'h42ad195d, 32'h0, 32'h42971ab4, 32'h427e4787, 32'h42679706};
test_input[31840:31847] = '{32'hc004db0e, 32'hc115699e, 32'hc2a89b0c, 32'hc219f5d6, 32'hc1835fd2, 32'h428a0c84, 32'h417c892e, 32'hc2c19a11};
test_output[31840:31847] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428a0c84, 32'h417c892e, 32'h0};
test_input[31848:31855] = '{32'hc2865f0d, 32'hc12b506a, 32'hc0e8496b, 32'hc2a40776, 32'h4224815c, 32'hc29a4cd5, 32'h41465e25, 32'h42434c85};
test_output[31848:31855] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4224815c, 32'h0, 32'h41465e25, 32'h42434c85};
test_input[31856:31863] = '{32'hc2add8c5, 32'h4282d258, 32'h41fd978b, 32'hc1ea419d, 32'hc28aad91, 32'h4143ac45, 32'h4280dd22, 32'h42ad3dbc};
test_output[31856:31863] = '{32'h0, 32'h4282d258, 32'h41fd978b, 32'h0, 32'h0, 32'h4143ac45, 32'h4280dd22, 32'h42ad3dbc};
test_input[31864:31871] = '{32'hc25a35c4, 32'hc28cfeaa, 32'h412baa43, 32'h42b7cae9, 32'h400709e8, 32'h42b36a8f, 32'hc2b1ddd2, 32'hc2185fc4};
test_output[31864:31871] = '{32'h0, 32'h0, 32'h412baa43, 32'h42b7cae9, 32'h400709e8, 32'h42b36a8f, 32'h0, 32'h0};
test_input[31872:31879] = '{32'hc2bd0453, 32'hc22289f3, 32'hc240af20, 32'hc24c4eb7, 32'h40914db4, 32'hc1f83508, 32'h4213e257, 32'h4026dd07};
test_output[31872:31879] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40914db4, 32'h0, 32'h4213e257, 32'h4026dd07};
test_input[31880:31887] = '{32'h4169e681, 32'hc2270874, 32'hc29e4c5c, 32'h414889fb, 32'hc29b77e0, 32'h42b0701a, 32'hc0ace618, 32'hc2c47d33};
test_output[31880:31887] = '{32'h4169e681, 32'h0, 32'h0, 32'h414889fb, 32'h0, 32'h42b0701a, 32'h0, 32'h0};
test_input[31888:31895] = '{32'h410c404f, 32'hc282d48f, 32'hc2c7ebcd, 32'h42929e02, 32'hc223bfe4, 32'hc2c7e146, 32'hc2749c1c, 32'h41868c84};
test_output[31888:31895] = '{32'h410c404f, 32'h0, 32'h0, 32'h42929e02, 32'h0, 32'h0, 32'h0, 32'h41868c84};
test_input[31896:31903] = '{32'h41e861a6, 32'h4240b5b2, 32'hc28c823e, 32'hc2157ec9, 32'h42a6818a, 32'hc233b6dd, 32'h4195d878, 32'h428882c6};
test_output[31896:31903] = '{32'h41e861a6, 32'h4240b5b2, 32'h0, 32'h0, 32'h42a6818a, 32'h0, 32'h4195d878, 32'h428882c6};
test_input[31904:31911] = '{32'h42aa36fe, 32'h422de3f8, 32'h42a6573f, 32'h4280050f, 32'h428292d1, 32'hc238c070, 32'h4148db45, 32'hc2bdd7ea};
test_output[31904:31911] = '{32'h42aa36fe, 32'h422de3f8, 32'h42a6573f, 32'h4280050f, 32'h428292d1, 32'h0, 32'h4148db45, 32'h0};
test_input[31912:31919] = '{32'hc03e9da7, 32'hc251216e, 32'h426f2b23, 32'hc019dff5, 32'h422783f0, 32'h4027ea59, 32'hc2c21709, 32'h4289c8d7};
test_output[31912:31919] = '{32'h0, 32'h0, 32'h426f2b23, 32'h0, 32'h422783f0, 32'h4027ea59, 32'h0, 32'h4289c8d7};
test_input[31920:31927] = '{32'h421faa9b, 32'h42ac1332, 32'hc188f4ac, 32'hc2ad52ea, 32'h417c7904, 32'h418b2503, 32'hc1e30112, 32'h427ffaff};
test_output[31920:31927] = '{32'h421faa9b, 32'h42ac1332, 32'h0, 32'h0, 32'h417c7904, 32'h418b2503, 32'h0, 32'h427ffaff};
test_input[31928:31935] = '{32'h4254fc21, 32'hc2c60435, 32'h42964557, 32'hc21c9cb8, 32'hc1f346a7, 32'hc0dd45ea, 32'hc17c9112, 32'hc2948178};
test_output[31928:31935] = '{32'h4254fc21, 32'h0, 32'h42964557, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31936:31943] = '{32'h42926afb, 32'h42c45077, 32'h4221bb70, 32'hc11f7bf8, 32'hc1acb860, 32'hc2432d34, 32'h4205ebda, 32'hc19abbb9};
test_output[31936:31943] = '{32'h42926afb, 32'h42c45077, 32'h4221bb70, 32'h0, 32'h0, 32'h0, 32'h4205ebda, 32'h0};
test_input[31944:31951] = '{32'hc0c221f7, 32'h416a94a5, 32'hc20b0c40, 32'h4233ca14, 32'hc18bef58, 32'h41fb8c43, 32'h41ec87ce, 32'h41fdfcdd};
test_output[31944:31951] = '{32'h0, 32'h416a94a5, 32'h0, 32'h4233ca14, 32'h0, 32'h41fb8c43, 32'h41ec87ce, 32'h41fdfcdd};
test_input[31952:31959] = '{32'hc21c9d97, 32'hc2a5e824, 32'hc1e573d8, 32'h42bc0219, 32'h42943c96, 32'h42816157, 32'hc1ad1d4f, 32'h4292d917};
test_output[31952:31959] = '{32'h0, 32'h0, 32'h0, 32'h42bc0219, 32'h42943c96, 32'h42816157, 32'h0, 32'h4292d917};
test_input[31960:31967] = '{32'h42789a3f, 32'h421ff921, 32'h4215b18c, 32'hc2929e4a, 32'hc2aa400d, 32'hc2be9f0f, 32'hc27a5c33, 32'h40e99c7e};
test_output[31960:31967] = '{32'h42789a3f, 32'h421ff921, 32'h4215b18c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40e99c7e};
test_input[31968:31975] = '{32'h4291aef2, 32'hc1e0863a, 32'hc23a963b, 32'hc24a04d3, 32'hc2783d15, 32'hc2790947, 32'h4193f3f1, 32'hc14d8d56};
test_output[31968:31975] = '{32'h4291aef2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4193f3f1, 32'h0};
test_input[31976:31983] = '{32'h42222aff, 32'hc26c13b3, 32'hc20c4eb2, 32'hc22d14c1, 32'hc295a673, 32'hc1d0eda0, 32'h42b276c1, 32'h42486c3f};
test_output[31976:31983] = '{32'h42222aff, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b276c1, 32'h42486c3f};
test_input[31984:31991] = '{32'hc1266270, 32'h41a206af, 32'h41989ef1, 32'h42c49a26, 32'h4268238e, 32'h426eaae8, 32'h420fff41, 32'h4226c296};
test_output[31984:31991] = '{32'h0, 32'h41a206af, 32'h41989ef1, 32'h42c49a26, 32'h4268238e, 32'h426eaae8, 32'h420fff41, 32'h4226c296};
test_input[31992:31999] = '{32'h3eabe276, 32'hc133d198, 32'h42bbd685, 32'hc20d1f17, 32'hc2c61439, 32'h42c2bb3c, 32'hc2a0088d, 32'h421b4701};
test_output[31992:31999] = '{32'h3eabe276, 32'h0, 32'h42bbd685, 32'h0, 32'h0, 32'h42c2bb3c, 32'h0, 32'h421b4701};
end
`endif
