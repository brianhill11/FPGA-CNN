`ifndef CONV_FORWARD_TEST_H
`define CONV_FORWARD_TEST_H
reg [31:0] test_input [32000];
reg [31:0] test_weights [32000];
reg [31:0] test_bias [4000];
reg [31:0] test_output [4000];
initial begin
test_input[0:7] = '{32'hc2b5bcd6, 32'hc1e4293e, 32'h42b85390, 32'h429eea86, 32'h42bfb4b5, 32'hc27dce65, 32'h42838edc, 32'h428ecfe9};
test_weights[0:7] = '{32'h424eadd8, 32'hc2b943ba, 32'hc08888d9, 32'hc2b76173, 32'h4263febc, 32'hc2c3638e, 32'h42a9439b, 32'h41bf92fe};
test_bias[0:0] = '{32'h419983ce};
test_output[0:0] = '{32'h461029d4};
test_input[8:15] = '{32'h418ee06a, 32'hc1f6e9bd, 32'hc0fed321, 32'hc0862694, 32'hc02b649d, 32'hc2adac45, 32'hc23889b2, 32'h4202804c};
test_weights[8:15] = '{32'h41f0e9af, 32'h4283d2ab, 32'h421243f9, 32'hc1a08572, 32'h42bb82ae, 32'h41e6d5b3, 32'hc212697d, 32'hc24c4463};
test_bias[1:1] = '{32'hc2c1e1a9};
test_output[1:1] = '{32'hc58db4a7};
test_input[16:23] = '{32'h42a3e99e, 32'hc0bc70be, 32'h41e7e295, 32'h42421f93, 32'h42807fa4, 32'h4279d8e0, 32'hc23206b6, 32'h42ae114a};
test_weights[16:23] = '{32'h4132f543, 32'h429086f1, 32'h421f7be7, 32'h42474472, 32'h419c9bfe, 32'hc19446ea, 32'h42b5121f, 32'hc177701d};
test_bias[2:2] = '{32'h4286677b};
test_output[2:2] = '{32'hc48ef54f};
test_input[24:31] = '{32'hc1ad1615, 32'h421ab132, 32'hc1859493, 32'hc2b16721, 32'h41b82f47, 32'h42b14ed6, 32'hc2bcb239, 32'h41c51b7f};
test_weights[24:31] = '{32'h4259700f, 32'hc195e1ee, 32'h41ccfbb4, 32'h4250b596, 32'hc2461834, 32'hc18cec60, 32'hc2a494be, 32'h429eeb71};
test_bias[3:3] = '{32'hc24e22e7};
test_output[3:3] = '{32'h4139dfb7};
test_input[32:39] = '{32'hc20ca15a, 32'h423aed03, 32'hc144de7a, 32'hc2662c29, 32'h4295b945, 32'h423a56b7, 32'hc2bf6140, 32'hc2bc545f};
test_weights[32:39] = '{32'h416108f8, 32'hc2918778, 32'h41395d9a, 32'hc29d895e, 32'hc22d1b03, 32'hc2a0861c, 32'h4154c17e, 32'h42729302};
test_bias[4:4] = '{32'h42660532};
test_output[4:4] = '{32'hc65183e4};
test_input[40:47] = '{32'h427a5106, 32'h42809f8c, 32'hc2a7a8ea, 32'h420c2087, 32'hc1e1608a, 32'h428699d5, 32'hc23b11ed, 32'h41e9c8d2};
test_weights[40:47] = '{32'h41e31541, 32'h424c54e1, 32'h4287fb30, 32'h42700ada, 32'h429260ce, 32'hc298c63c, 32'hc2aab28d, 32'hc18179a6};
test_bias[5:5] = '{32'hc22f1493};
test_output[5:5] = '{32'hc50d7c75};
test_input[48:55] = '{32'hc25c8b18, 32'h427ea900, 32'hc20c402a, 32'h427494b7, 32'hc2b00334, 32'hc20ff5d9, 32'hbfb43686, 32'hc033d65e};
test_weights[48:55] = '{32'hc2a1d41a, 32'h42ab81c3, 32'hc28aa7d7, 32'hc2b6afd7, 32'h42697b33, 32'hc1b10a4d, 32'h42b10163, 32'h42500fa4};
test_bias[6:6] = '{32'h4210d5a6};
test_output[6:6] = '{32'h4508f538};
test_input[56:63] = '{32'h4259a376, 32'hc25824b9, 32'hc294e6ee, 32'hc2a46bed, 32'hc2ad98ea, 32'h41ee11a7, 32'hc27c638e, 32'hc27d1335};
test_weights[56:63] = '{32'hc254bd80, 32'hc014832e, 32'h426f2b28, 32'h42c61d75, 32'h428d9bae, 32'h428da446, 32'hc207c3a4, 32'h41a609d2};
test_bias[7:7] = '{32'h428cf1b1};
test_output[7:7] = '{32'hc6908da1};
test_input[64:71] = '{32'h42690849, 32'h4251a359, 32'hc2c07460, 32'hc1e5a503, 32'h42aec944, 32'hc16c033e, 32'h41856e92, 32'h423cabd3};
test_weights[64:71] = '{32'h42442738, 32'h42305482, 32'hc298a433, 32'h417cc1ba, 32'h42ab810c, 32'h42139c64, 32'h41ee33c9, 32'h4209552d};
test_bias[8:8] = '{32'h429ac46d};
test_output[8:8] = '{32'h46a5a235};
test_input[72:79] = '{32'h40ad4d54, 32'hc1baad52, 32'h41d144c7, 32'hc2aa6685, 32'hc2900b90, 32'h4186a684, 32'h42b537c2, 32'hc2c394ca};
test_weights[72:79] = '{32'hc259130f, 32'h420b412d, 32'hc1bcbf7b, 32'h4270f835, 32'hc280bc8d, 32'h41584593, 32'hc05fae27, 32'hc2320ad3};
test_bias[9:9] = '{32'hbff497ab};
test_output[9:9] = '{32'h44ff2ffc};
test_input[80:87] = '{32'hc1839971, 32'h422d6208, 32'hc1603a98, 32'hc220809d, 32'hc2b2b059, 32'h42bfadb0, 32'hc280ef85, 32'hc2b49f2c};
test_weights[80:87] = '{32'h4239824e, 32'hc2a974bf, 32'h3f7557c5, 32'h41d194cb, 32'hc2b2de37, 32'hc245514c, 32'h4282f310, 32'h42bfd87b};
test_bias[10:10] = '{32'h42b0b2c7};
test_output[10:10] = '{32'hc66ae3b4};
test_input[88:95] = '{32'hc1d3ae5b, 32'h4253fb6e, 32'h4253cd1d, 32'h42a5d6ef, 32'h423ea187, 32'hc2b6fc74, 32'hc2a44b99, 32'h3e113bad};
test_weights[88:95] = '{32'hc1a74ca6, 32'h42845196, 32'h42817ba3, 32'h428a874e, 32'hc2a3040b, 32'hc23efc90, 32'h408224e5, 32'hc143bd66};
test_bias[11:11] = '{32'h41e7b269};
test_output[11:11] = '{32'h4651805e};
test_input[96:103] = '{32'h428cd782, 32'hc2a11985, 32'hc2a96490, 32'h42b25e5b, 32'hc294088d, 32'h418c23a6, 32'h418801a7, 32'h42a56baa};
test_weights[96:103] = '{32'h42234a8a, 32'h4266c53c, 32'h42ab9330, 32'h411350fb, 32'h42b1f46f, 32'hc18caf83, 32'h40b1a42e, 32'hc224744e};
test_bias[12:12] = '{32'hc1e0a197};
test_output[12:12] = '{32'hc6901a60};
test_input[104:111] = '{32'hc2a40894, 32'h410daa93, 32'h4217fbb2, 32'h3e552a1a, 32'hc2a9e150, 32'h41f057d2, 32'hc2874746, 32'h421980de};
test_weights[104:111] = '{32'h427f67fa, 32'h420f24a6, 32'hc242c43d, 32'h427dbf07, 32'hc246a1c3, 32'h41dac04a, 32'h425df8c2, 32'hc2be16e3};
test_bias[13:13] = '{32'h422e8f00};
test_output[13:13] = '{32'hc60dcb04};
test_input[112:119] = '{32'h413b14da, 32'h42803516, 32'hc26a880b, 32'hc190ed3d, 32'hc13928f4, 32'hc27acef9, 32'h4120683d, 32'hc286d09a};
test_weights[112:119] = '{32'hc09c2b40, 32'hc2554b4f, 32'h429e9eca, 32'hc23d3c90, 32'h42227617, 32'hc21512cf, 32'hc27260d5, 32'hc2be6d2f};
test_bias[14:14] = '{32'hc2aa5bf0};
test_output[14:14] = '{32'h43a1e1cd};
test_input[120:127] = '{32'hc267693b, 32'h425b6e78, 32'h4223f3bc, 32'hc286eee9, 32'hc1620216, 32'h41c4c1b8, 32'hc26760aa, 32'hc1650de6};
test_weights[120:127] = '{32'hc2ac9721, 32'h4290510f, 32'h429295fb, 32'hc2377faa, 32'hc29b6a4e, 32'h42a310c1, 32'hc1f27165, 32'hc05155fc};
test_bias[15:15] = '{32'h42391acd};
test_output[15:15] = '{32'h469c3e0f};
test_input[128:135] = '{32'hc11a5bbb, 32'h4297c607, 32'h411ff367, 32'hc27ac0ee, 32'hc2908554, 32'hc22830a8, 32'hc1f2bd11, 32'hc2a1fcc2};
test_weights[128:135] = '{32'hc1b78b75, 32'h426a7f80, 32'hc1978fe4, 32'hc2a2a067, 32'hc1a33b13, 32'h42b4fd6e, 32'h42b48c27, 32'hc0ad0de9};
test_bias[16:16] = '{32'h4184e9ca};
test_output[16:16] = '{32'h459b17dc};
test_input[136:143] = '{32'h41fea713, 32'hc22d526e, 32'hc1ea25eb, 32'h42c2fe4b, 32'h3f0647ae, 32'hc2639cbc, 32'h426beb90, 32'hc29a980c};
test_weights[136:143] = '{32'hc28d4243, 32'h4208b88a, 32'hc2c0e457, 32'h42771e87, 32'hc2ba81f3, 32'h412c1833, 32'hc23497b5, 32'hc1f44b7b};
test_bias[17:17] = '{32'h40266d02};
test_output[17:17] = '{32'h4581e095};
test_input[144:151] = '{32'h42c5b01b, 32'h4291e6d2, 32'h428f0edf, 32'h41b5359d, 32'hc219b715, 32'h426067d0, 32'hc2820887, 32'hc2c589d4};
test_weights[144:151] = '{32'h422cc9ac, 32'hc248d25c, 32'hc2bf1f7a, 32'hc289afe6, 32'hc28afc39, 32'h41ac426f, 32'h3f97ff33, 32'hc271d396};
test_bias[18:18] = '{32'hc1a6aa93};
test_output[18:18] = '{32'h44f584d7};
test_input[152:159] = '{32'hc1f6da1f, 32'h42270398, 32'h42b8148f, 32'h3f9684b4, 32'h420b72f0, 32'hc172a386, 32'hc2bb96c8, 32'hc22577ff};
test_weights[152:159] = '{32'hc26027dd, 32'h42056ec7, 32'hc20117e7, 32'h42a44606, 32'hc2a7c6ea, 32'h413677b5, 32'hbfd612bc, 32'hc1db7948};
test_bias[19:19] = '{32'h419d35d8};
test_output[19:19] = '{32'hc4c03ec4};
test_input[160:167] = '{32'hc2c6d42f, 32'hc2bfb29d, 32'hc28322fa, 32'h424fdbdb, 32'h41e9eb52, 32'hc25e48c8, 32'h40817e61, 32'hc1da8a43};
test_weights[160:167] = '{32'h42761e6b, 32'h42916828, 32'h4124e33f, 32'hc14612ac, 32'h42a643d2, 32'h42a61ecf, 32'hc291a6f8, 32'h41eee868};
test_bias[20:20] = '{32'h42103bff};
test_output[20:20] = '{32'hc689ffc9};
test_input[168:175] = '{32'h41feb1b8, 32'h4253f062, 32'h4287cb2d, 32'hc29b4de6, 32'hc20eb456, 32'hc152bdd7, 32'h4263a053, 32'h4259ec3a};
test_weights[168:175] = '{32'h41d4e8df, 32'hc1896ac3, 32'hc290d36b, 32'hc2bb1774, 32'hc221c0d7, 32'h4216e063, 32'h41def7bb, 32'hc2ac4381};
test_bias[21:21] = '{32'h42b133e4};
test_output[21:21] = '{32'h4354955e};
test_input[176:183] = '{32'hc1c23625, 32'h428cec25, 32'hc2b9f211, 32'h3faeeb50, 32'hc2a20687, 32'h41ee5ab4, 32'h421e8bf0, 32'h418fb9ca};
test_weights[176:183] = '{32'hc2b6829a, 32'hc22eca0b, 32'h428f7f61, 32'hc18fafda, 32'hc29eebbd, 32'hc23ebc9a, 32'h41a86b83, 32'hc29a9e0e};
test_bias[22:22] = '{32'h42adaf19};
test_output[22:22] = '{32'hc53c1de6};
test_input[184:191] = '{32'hc2840d79, 32'h4104579f, 32'h42b62a53, 32'h4226d183, 32'h41d3a22a, 32'h428d4fca, 32'h42c7449c, 32'h420fe74a};
test_weights[184:191] = '{32'hc238fe63, 32'hc2a2e3ac, 32'h42848a68, 32'hc1ef375c, 32'h425b408d, 32'h420e5b6f, 32'hc188f1d4, 32'h42a49241};
test_bias[23:23] = '{32'h42bbacc1};
test_output[23:23] = '{32'h464308c8};
test_input[192:199] = '{32'hc227f363, 32'hc2b78a0c, 32'h429b4bff, 32'hc24130db, 32'hc22fba9b, 32'hc103cc64, 32'hc20baa82, 32'h4244c3ae};
test_weights[192:199] = '{32'h4214ab8e, 32'h40c2474e, 32'h41d9fb9f, 32'h42b201b2, 32'h428924be, 32'hc19f1e3a, 32'hc2c15c66, 32'h4293cbf8};
test_bias[24:24] = '{32'h42a3714c};
test_output[24:24] = '{32'hc262c875};
test_input[200:207] = '{32'h41478a84, 32'hc2504517, 32'h418f67c8, 32'h42c26ab8, 32'hc288a236, 32'hc231955e, 32'h427dbf81, 32'h40529c5a};
test_weights[200:207] = '{32'h42aa6d9e, 32'hc1b70d25, 32'hc2afa618, 32'hc23b0e2f, 32'hc259b6cf, 32'hc15d1ba6, 32'h429e0889, 32'hc0be4e13};
test_bias[25:25] = '{32'h42391618};
test_output[25:25] = '{32'h45ac0921};
test_input[208:215] = '{32'hc2a6df08, 32'h425b77dd, 32'h428d5354, 32'h42978cb5, 32'hc26e17ab, 32'hc14cbcb1, 32'hc2542331, 32'h413bcb8c};
test_weights[208:215] = '{32'h42a55359, 32'h4290d1a2, 32'h41fa539b, 32'hc2b5007b, 32'h42315598, 32'h40b7d5e2, 32'hc29e82b7, 32'h422e1527};
test_bias[26:26] = '{32'h4185e0c7};
test_output[26:26] = '{32'hc5ad827a};
test_input[216:223] = '{32'h42764d09, 32'hc1a2e577, 32'hc198c471, 32'hc08b01a3, 32'h4218c77f, 32'h4249fa2e, 32'hc24d431b, 32'hc1f13a6c};
test_weights[216:223] = '{32'hc23f7433, 32'hc1d31654, 32'h426d3fa2, 32'hc2b9651e, 32'h427fd445, 32'hc1ecaf1f, 32'h41b4de72, 32'hc222a9a0};
test_bias[27:27] = '{32'h428ad621};
test_output[27:27] = '{32'hc50077c3};
test_input[224:231] = '{32'hc0cf555e, 32'h3e8443e8, 32'h4102b9ab, 32'h4282d569, 32'hc267aa6a, 32'h4219df2b, 32'hc291ca4e, 32'h41e41b5f};
test_weights[224:231] = '{32'hc231e47e, 32'h42abbdad, 32'h42840e7c, 32'hc28dad21, 32'hc2150792, 32'h424ff3f4, 32'hc28053ee, 32'hc2bf3c72};
test_bias[28:28] = '{32'h42b12532};
test_output[28:28] = '{32'h4516ce95};
test_input[232:239] = '{32'hc2c41a24, 32'h4279bd68, 32'h42c17720, 32'hc08368d4, 32'hc2106250, 32'h427cba40, 32'hc1b632a5, 32'hc2b83fe5};
test_weights[232:239] = '{32'h42777235, 32'hc248bb69, 32'h4166ca62, 32'hc23c0b7c, 32'h4281a600, 32'h41df1fe8, 32'h417ee4d0, 32'hc29272a9};
test_bias[29:29] = '{32'hc2b180eb};
test_output[29:29] = '{32'hc4ecbe48};
test_input[240:247] = '{32'h42353d26, 32'h422a3ad5, 32'h42c7ac7c, 32'h42bfcef1, 32'hc20a5143, 32'h41b925a3, 32'hc26e52ca, 32'h4189f8cf};
test_weights[240:247] = '{32'h41a2b409, 32'hc29d82a6, 32'hc2894ca3, 32'hc28d2233, 32'hc1d77d52, 32'h41f13707, 32'h42205a45, 32'hc178762a};
test_bias[30:30] = '{32'h3d942559};
test_output[30:30] = '{32'hc6856d08};
test_input[248:255] = '{32'h42377e84, 32'h41759c3a, 32'hc1bf4386, 32'hc206c34c, 32'h42910ba7, 32'h42904eda, 32'h42464566, 32'h408d6a6a};
test_weights[248:255] = '{32'h425ad711, 32'h429d24ba, 32'hc2adcb9d, 32'hc29a6847, 32'hc2b4279d, 32'h4250fb91, 32'hc22008c2, 32'h41c284c0};
test_bias[31:31] = '{32'h4200aeda};
test_output[31:31] = '{32'h456cc072};
test_input[256:263] = '{32'hc1bc57f4, 32'h4181d803, 32'h41762ed3, 32'h41b2cbc1, 32'h41b5fd95, 32'h421d5bf0, 32'h4213dc44, 32'h42b087f7};
test_weights[256:263] = '{32'hc2bf3257, 32'hc2a451e3, 32'h427218ca, 32'h42bee64d, 32'h42c58f8e, 32'h4208bcac, 32'hc1b3e204, 32'h416f0f7c};
test_bias[32:32] = '{32'h411078d0};
test_output[32:32] = '{32'h45fc322d};
test_input[264:271] = '{32'h41cd0da4, 32'h42c5abfc, 32'hc1c7b195, 32'hc2ac0cd0, 32'h419c2977, 32'hc2a241da, 32'hc28d6feb, 32'hc2a6dfc1};
test_weights[264:271] = '{32'hc251b896, 32'h42bb7e56, 32'hc074296a, 32'h4287448f, 32'hc289525b, 32'hc23a80d6, 32'hc2b28fdf, 32'h42a47b72};
test_bias[33:33] = '{32'h424b4c5d};
test_output[33:33] = '{32'h45817e68};
test_input[272:279] = '{32'hc2959205, 32'h4295cee8, 32'h4225003c, 32'h423a723e, 32'hc24d98ed, 32'h41bb0866, 32'hc2c0685f, 32'h428902d0};
test_weights[272:279] = '{32'hc262f1fb, 32'hc21c1ac8, 32'h4271977b, 32'h41c996af, 32'h4178fdd0, 32'h4189dbb8, 32'hc197b217, 32'h42736177};
test_bias[34:34] = '{32'hc29eafed};
test_output[34:34] = '{32'h4624178e};
test_input[280:287] = '{32'h42880cfc, 32'hc2aff931, 32'h41217994, 32'h428b18f8, 32'h40d74907, 32'h41e90bc0, 32'h42488ea6, 32'hc08335a7};
test_weights[280:287] = '{32'h42a12383, 32'hc2042caf, 32'h422d9aee, 32'h428bc4f2, 32'hc0e48734, 32'hc21db974, 32'h4076c839, 32'hc16a2510};
test_bias[35:35] = '{32'hc12b0e30};
test_output[35:35] = '{32'h4646f20c};
test_input[288:295] = '{32'hc23ae6ec, 32'hc204353d, 32'h42540ff5, 32'hc0f49897, 32'h42a10926, 32'hc26a5cc2, 32'hc2a10239, 32'hc1096227};
test_weights[288:295] = '{32'h42abb174, 32'h40f83dd5, 32'h42a1b9a1, 32'hc2a877c8, 32'h42142ec8, 32'h42377759, 32'hc2af817b, 32'h42b563fe};
test_bias[36:36] = '{32'hc18076ff};
test_output[36:36] = '{32'h45e1e2f8};
test_input[296:303] = '{32'h4294bd84, 32'h42aad8a4, 32'hc1baef90, 32'h42069deb, 32'h42823517, 32'hc214cab6, 32'h427bdb33, 32'hc0c38966};
test_weights[296:303] = '{32'h419d62ce, 32'h42ac079e, 32'hc2364ab4, 32'h422895c5, 32'h3fa6af6b, 32'hc1d36890, 32'h4229dd66, 32'h41b70cd4};
test_bias[37:37] = '{32'h3f176315};
test_output[37:37] = '{32'h4668c1d5};
test_input[304:311] = '{32'hc23a9176, 32'h42723319, 32'h420a0392, 32'h41eac4cc, 32'h42a7778e, 32'hc2af93fd, 32'h4276229a, 32'h42b1255a};
test_weights[304:311] = '{32'hc2a4774a, 32'hc2400a9c, 32'h42637f56, 32'h4109ae06, 32'hc2b2f051, 32'h42095546, 32'hc2865e0e, 32'hc22978ac};
test_bias[38:38] = '{32'hc1fcc123};
test_output[38:38] = '{32'hc66ec264};
test_input[312:319] = '{32'hc0fc8644, 32'hc20cc09d, 32'hc234fd07, 32'h4093bf1e, 32'h41859d41, 32'hc02ce16d, 32'hc01bd06c, 32'h40f2bd1d};
test_weights[312:319] = '{32'h416395cf, 32'hc1cb3e7e, 32'h42a9557c, 32'hc1c461b5, 32'h4013767d, 32'h41f49f18, 32'hc19077a8, 32'hc25582cc};
test_bias[39:39] = '{32'hc20e683e};
test_output[39:39] = '{32'hc561333e};
test_input[320:327] = '{32'h40603a2b, 32'h41302a52, 32'hc2aa5487, 32'hc2aba88d, 32'h4219b0d7, 32'hc28029bf, 32'h4262eef5, 32'hc2bd17d3};
test_weights[320:327] = '{32'h41d326c5, 32'h4129077c, 32'hc1d0703e, 32'h4199e258, 32'hc298abea, 32'hc2bd98fe, 32'hc1872db3, 32'hc14bcd03};
test_bias[40:40] = '{32'hc1fac6d0};
test_output[40:40] = '{32'h45812749};
test_input[328:335] = '{32'h4224e54b, 32'hc2ab5a7c, 32'hc29cf6a3, 32'h426f333f, 32'hc2b936f8, 32'hc2875ab9, 32'h42644350, 32'hc2b11d21};
test_weights[328:335] = '{32'hc2c69b73, 32'h42974d27, 32'hc294da63, 32'hc2a1458f, 32'h4283c8ac, 32'h4013f145, 32'h42b4efbf, 32'hc29c6512};
test_bias[41:41] = '{32'hc2805763};
test_output[41:41] = '{32'hc56cf3a8};
test_input[336:343] = '{32'h4267b349, 32'h41952845, 32'hc2af25b0, 32'hc2697aaa, 32'hc2375fe1, 32'h4279a54a, 32'hc1a7ff8c, 32'hc2a1e97a};
test_weights[336:343] = '{32'hc240ea97, 32'hc2b7b485, 32'h4181fda6, 32'h41b83d1f, 32'hc057de54, 32'h40d35079, 32'h41847c1e, 32'hc2a7c84d};
test_bias[42:42] = '{32'hc290018c};
test_output[42:42] = '{32'hc3a77adf};
test_input[344:351] = '{32'hc21b9b6d, 32'h4288ee79, 32'hc22e925b, 32'h42a9ff40, 32'hc1bd5461, 32'hc1cbd2d6, 32'h4173f4b2, 32'h41a61337};
test_weights[344:351] = '{32'h420507f9, 32'h4297e9b2, 32'hc282c0ab, 32'hc2b7490c, 32'hc1851d48, 32'hc115cce7, 32'h4286ad01, 32'h418da56f};
test_bias[43:43] = '{32'hc2315166};
test_output[43:43] = '{32'h446e27f3};
test_input[352:359] = '{32'h41acc5c1, 32'hc154e6dc, 32'h428e9126, 32'h42b76bb2, 32'hc24ec6c3, 32'hc2c18176, 32'h4221545d, 32'hc1ae1835};
test_weights[352:359] = '{32'hc189bfdf, 32'hc0238e15, 32'hc1281be9, 32'h42600376, 32'hc24ba218, 32'h42371b4c, 32'hc236ab7b, 32'hc2baf18c};
test_bias[44:44] = '{32'hc2947049};
test_output[44:44] = '{32'h45141ec4};
test_input[360:367] = '{32'hc2ba6d7c, 32'hc2783ac4, 32'h42ac41e1, 32'hc2c65bff, 32'hc2a7b768, 32'h4136d855, 32'h42c08e48, 32'h418bbb82};
test_weights[360:367] = '{32'hc2b7a862, 32'hc24f5138, 32'hc1c67241, 32'hc218b25f, 32'hc28ecc68, 32'hc2256b65, 32'hc218828f, 32'hc1b8f9d7};
test_bias[45:45] = '{32'hc21e9829};
test_output[45:45] = '{32'h4667a8cb};
test_input[368:375] = '{32'h4143280d, 32'hc29e3ed7, 32'hc1649eb2, 32'h42229b24, 32'hc1b5de18, 32'hc2878698, 32'h4273e38c, 32'h42443fe3};
test_weights[368:375] = '{32'h42b84724, 32'hc297d59d, 32'h4277cc41, 32'hbe0d7963, 32'hc21f6d0b, 32'h415de017, 32'h4202ecd2, 32'hc23824ec};
test_bias[46:46] = '{32'hc09eb535};
test_output[46:46] = '{32'h45b9928b};
test_input[376:383] = '{32'hc1a56cdd, 32'hc24c7ddd, 32'h4293646c, 32'hc250b217, 32'hc20cca89, 32'hc2c3c337, 32'hc22bebbe, 32'hc263125a};
test_weights[376:383] = '{32'h420cf078, 32'h421d9a36, 32'h4254629c, 32'h4271e249, 32'hc2104aae, 32'hc28708dc, 32'hc2c71b98, 32'hc249f5b5};
test_bias[47:47] = '{32'hc1f9eae8};
test_output[47:47] = '{32'h464b3d37};
test_input[384:391] = '{32'hc23f4865, 32'hc2bcca27, 32'hc278a069, 32'hc2a292b5, 32'h423e4a0e, 32'hc188f180, 32'hc0a15be1, 32'h42369161};
test_weights[384:391] = '{32'h419dddbd, 32'h416a874a, 32'hc0e76881, 32'hc1b9ac9c, 32'h42766489, 32'h411e5e85, 32'hc23c5bb2, 32'h424c59df};
test_bias[48:48] = '{32'h426cae6b};
test_output[48:48] = '{32'h45a8b0af};
test_input[392:399] = '{32'hc2b7cd6a, 32'h42ab0c70, 32'h4286aaf7, 32'h4221dd2d, 32'hc29d1781, 32'h42526877, 32'hc2c43ba2, 32'hc09d7ffb};
test_weights[392:399] = '{32'hc1ef0b07, 32'hbe84e50f, 32'h4279a573, 32'hc1ae25c0, 32'h42b25e54, 32'h3f296455, 32'h42455e63, 32'hc26375f9};
test_bias[49:49] = '{32'h429d3132};
test_output[49:49] = '{32'hc5a8fd62};
test_input[400:407] = '{32'hc2bd775c, 32'hc24d2644, 32'h423c20d5, 32'h400a703d, 32'hc26962ac, 32'h42111f2b, 32'hc28b40f3, 32'h41359ff1};
test_weights[400:407] = '{32'hc2579cec, 32'hc24886eb, 32'h42531d54, 32'h42b2bb34, 32'h4259e86f, 32'h41b8c5cb, 32'hc295c28e, 32'hc2323b2d};
test_bias[50:50] = '{32'h425193ff};
test_output[50:50] = '{32'h46479344};
test_input[408:415] = '{32'h42985522, 32'hc2ae104b, 32'hc202b7f5, 32'h41dfd1ef, 32'hc1c31577, 32'h40d4641c, 32'hc27dd26a, 32'h4125f7f8};
test_weights[408:415] = '{32'h429c4bc7, 32'h42b0e1bc, 32'hc2304493, 32'hc2be5774, 32'hc2188fa7, 32'hc259a835, 32'hc1a59ff0, 32'hc2079a25};
test_bias[51:51] = '{32'hc29442c0};
test_output[51:51] = '{32'hc4bcd402};
test_input[416:423] = '{32'h42c37c32, 32'h42bfd156, 32'h4281f587, 32'h418ef625, 32'h420bd982, 32'h42b25cdd, 32'hc0af254e, 32'hc29f0e86};
test_weights[416:423] = '{32'hc1718041, 32'hc28aeec8, 32'hc0e235ec, 32'hc26a556e, 32'hc2a8e6a3, 32'hc2949d5a, 32'h41899d6f, 32'h4290f8ef};
test_bias[52:52] = '{32'hc279240a};
test_output[52:52] = '{32'hc6c4711d};
test_input[424:431] = '{32'hc108382e, 32'hc272afe9, 32'hc292e1f0, 32'hc18e0527, 32'h426ab302, 32'h42525386, 32'hc2982e3f, 32'hc13f3cd1};
test_weights[424:431] = '{32'h42c07fcf, 32'h42437220, 32'hc2a2ad52, 32'h41bf8c51, 32'h41a02199, 32'h42c22677, 32'h421e0c9c, 32'h424a31ba};
test_bias[53:53] = '{32'hc0807c89};
test_output[53:53] = '{32'h458a65c5};
test_input[432:439] = '{32'hc2b096e1, 32'h429deac5, 32'h428b2754, 32'h42276c19, 32'h4141328f, 32'h41c6658d, 32'hc23067d5, 32'h427b7028};
test_weights[432:439] = '{32'hc248563a, 32'hc28cd838, 32'hc20fa281, 32'hc294430a, 32'h41682ca7, 32'hc1c45ae6, 32'hc29eacb9, 32'h42871298};
test_bias[54:54] = '{32'h422f1618};
test_output[54:54] = '{32'h4419c09d};
test_input[440:447] = '{32'hc1d7b496, 32'h40c81161, 32'h42162118, 32'hc21d0523, 32'h41e58215, 32'h420cb4bb, 32'h426b22c9, 32'h4293e76f};
test_weights[440:447] = '{32'hc2820ac4, 32'h42bedff3, 32'hc2b324fb, 32'hc2196a6c, 32'hc1b436ed, 32'h42989e5d, 32'hc2a5c04d, 32'h425765d4};
test_bias[55:55] = '{32'hc03ead7d};
test_output[55:55] = '{32'h44cce535};
test_input[448:455] = '{32'h426bcc8b, 32'h429c325a, 32'hc286aef9, 32'h406d9671, 32'hc2311526, 32'hc2370bad, 32'h42a9d879, 32'h422b839c};
test_weights[448:455] = '{32'hc24ccf46, 32'h41c06908, 32'h41a5fd87, 32'h40b7a7d0, 32'h41b4ef99, 32'h41b6e9ba, 32'h4235257e, 32'h424e4ae9};
test_bias[56:56] = '{32'h41db3d63};
test_output[56:56] = '{32'h44be2426};
test_input[456:463] = '{32'h41a00e61, 32'h42a2b131, 32'hc2969702, 32'h421fbe02, 32'h40cd24cf, 32'h427d6c77, 32'h4102e437, 32'hc20efa0f};
test_weights[456:463] = '{32'h42af52ce, 32'hc16232c2, 32'hc0b47538, 32'h4121729e, 32'h428c971f, 32'hc15b1358, 32'h4299c938, 32'h426db613};
test_bias[57:57] = '{32'hc2bed4c5};
test_output[57:57] = '{32'hc4100056};
test_input[464:471] = '{32'h425ae933, 32'h4283e577, 32'h4207511e, 32'h42a67762, 32'hc28f9557, 32'h42744741, 32'h42ad2197, 32'hc23d56ab};
test_weights[464:471] = '{32'hc20b8d3f, 32'h42c18681, 32'h4287de37, 32'h42c4a112, 32'h42b5509b, 32'hc1f051e9, 32'h4096b065, 32'hc1db5e65};
test_bias[58:58] = '{32'h3e99725f};
test_output[58:58] = '{32'h4601f06a};
test_input[472:479] = '{32'hc28d6010, 32'hc1c96f92, 32'h41f6349f, 32'hbeacb1ae, 32'h426e3b1f, 32'h4264420a, 32'hc2b41c53, 32'hc252fd87};
test_weights[472:479] = '{32'hc2ab4932, 32'hc23c32be, 32'h42500f57, 32'h42a78d0c, 32'hc1d2eb69, 32'h429710a4, 32'hc249bac2, 32'h424aa204};
test_bias[59:59] = '{32'hc0854a99};
test_output[59:59] = '{32'h4651a231};
test_input[480:487] = '{32'h426a04b7, 32'h40fe9f8d, 32'hc1c0e73d, 32'hc2105434, 32'h428c18a3, 32'hc1819a9b, 32'h42593fa4, 32'h428c846b};
test_weights[480:487] = '{32'h42743d3e, 32'hc230b1b8, 32'h42ab0e9c, 32'hc1688b3b, 32'h429a1b1e, 32'h41c0c2f5, 32'h421d0a5b, 32'hc2ab9ee2};
test_bias[60:60] = '{32'hc2904958};
test_output[60:60] = '{32'h452a12c6};
test_input[488:495] = '{32'hbf77599d, 32'hc1465517, 32'h424e3c76, 32'hc2c1f287, 32'hc2a317e6, 32'h4248e8b2, 32'hc25e00d5, 32'hc19d26b9};
test_weights[488:495] = '{32'h42bfd7c1, 32'hc25a31cd, 32'hc20a3f07, 32'h42bca0c6, 32'hc1deaf0e, 32'h4294b5a5, 32'h416c9539, 32'hc0c08a81};
test_bias[61:61] = '{32'hc2a99110};
test_output[61:61] = '{32'hc5a03956};
test_input[496:503] = '{32'h425d8aca, 32'h40708435, 32'h417f20fb, 32'hc28bf173, 32'hc2885555, 32'hc11889c9, 32'hc29447cd, 32'h428bb1a1};
test_weights[496:503] = '{32'hc127514e, 32'h42a9ba3c, 32'hc1653616, 32'h4299b105, 32'h428a3c1c, 32'hc1917385, 32'h428ac575, 32'hc2a91e33};
test_bias[62:62] = '{32'h42044296};
test_output[62:62] = '{32'hc6a75a8a};
test_input[504:511] = '{32'h4071a16d, 32'hc24f35bb, 32'hc28b3b42, 32'hc2b2122b, 32'hc2c37cf6, 32'h427f043b, 32'hc2abab1e, 32'hc27ae118};
test_weights[504:511] = '{32'h419dc72f, 32'h429df1e8, 32'h41862af6, 32'h42c3aae6, 32'hc1d92610, 32'hc2a7c171, 32'h425f2568, 32'h42c488fa};
test_bias[63:63] = '{32'hc2a4bfc1};
test_output[63:63] = '{32'hc6d7ce77};
test_input[512:519] = '{32'hc102685d, 32'hc2a353b9, 32'hc1ed0eaf, 32'hc1978070, 32'h426bb544, 32'hc161d189, 32'hc280d73e, 32'hc20e5fa9};
test_weights[512:519] = '{32'h425a719b, 32'h42a2ce21, 32'hc23e1c23, 32'h42a3eede, 32'h4104e819, 32'h42962e32, 32'h4246bc33, 32'h40b9c35b};
test_bias[64:64] = '{32'hbf1d70e5};
test_output[64:64] = '{32'hc62f3b5f};
test_input[520:527] = '{32'hc25f5d16, 32'h425314cf, 32'hc2bba4a4, 32'h420ad6c8, 32'hc289096f, 32'h3fafee03, 32'h410640cd, 32'hc192c5e0};
test_weights[520:527] = '{32'h423284c8, 32'h4298e329, 32'hbfbdd533, 32'hc17a00ac, 32'h421d797f, 32'h42897394, 32'h42a6ca50, 32'h3f95da81};
test_bias[65:65] = '{32'hc2aedc00};
test_output[65:65] = '{32'hc45a6505};
test_input[528:535] = '{32'hc2148893, 32'h41810169, 32'h4285383e, 32'h42028741, 32'h4066e585, 32'hc29af2da, 32'h40f0fd2a, 32'h42088b15};
test_weights[528:535] = '{32'h41cbb90d, 32'hc145d84b, 32'h411dcbd8, 32'h42ba7e79, 32'h423dfb59, 32'hc18fe223, 32'hc1f50c97, 32'hbda6e64f};
test_bias[66:66] = '{32'hc27147f3};
test_output[66:66] = '{32'h456f1bba};
test_input[536:543] = '{32'hc28c88d2, 32'h42c3a834, 32'hc2c44ecc, 32'h42c78121, 32'hc185a54c, 32'hbfc63e5c, 32'h42a9a67f, 32'h4234526c};
test_weights[536:543] = '{32'h42218350, 32'hc224f509, 32'h425dfdd6, 32'h42c7d8d8, 32'h42106964, 32'hc2157e40, 32'h4249798a, 32'hc29f1ad8};
test_bias[67:67] = '{32'h42bb01f8};
test_output[67:67] = '{32'hc5044daf};
test_input[544:551] = '{32'hc254254e, 32'hc2368c04, 32'hc2a70415, 32'h418d21e0, 32'h418ba642, 32'hc21857d4, 32'h42a030b6, 32'h42887883};
test_weights[544:551] = '{32'hc284df22, 32'hc2324030, 32'hbfb258dc, 32'hc0372248, 32'hc226202b, 32'hbf9dcfb6, 32'hc291526e, 32'hc24511e4};
test_bias[68:68] = '{32'h426f89d1};
test_output[68:68] = '{32'hc5828508};
test_input[552:559] = '{32'h40ca7002, 32'hc18ed07f, 32'hc2798715, 32'h42a36953, 32'hc1f03315, 32'hc2933638, 32'h427e81c9, 32'hc2b7d453};
test_weights[552:559] = '{32'h4296ce1b, 32'h42a622a5, 32'h42934db4, 32'hc2513019, 32'h41d90298, 32'hc0c112da, 32'h429c5460, 32'h42a291a0};
test_bias[69:69] = '{32'hc29e3164};
test_output[69:69] = '{32'hc64852dd};
test_input[560:567] = '{32'h418e60da, 32'hbf81a74a, 32'hc239efbe, 32'hc23cd926, 32'h429fbb79, 32'hc208c62f, 32'h4113a674, 32'hc0bf16ff};
test_weights[560:567] = '{32'hc18e5518, 32'h4226e59f, 32'hc2c1e1d5, 32'h429edee8, 32'h40f274c4, 32'h3f1b7e8e, 32'hc2be8b7a, 32'h42230f54};
test_bias[70:70] = '{32'h420d1b79};
test_output[70:70] = '{32'hc2d3f2b5};
test_input[568:575] = '{32'h42a4486e, 32'hc2589852, 32'h42b8b35d, 32'hc14161a3, 32'h41ea9a7d, 32'hc0001614, 32'hc18b4c70, 32'h4224e34e};
test_weights[568:575] = '{32'hc2b09dc2, 32'h429b7083, 32'h41360661, 32'hc2545af7, 32'h40c8f8a3, 32'h421084f1, 32'h42669193, 32'hc269e5ac};
test_bias[71:71] = '{32'hc2a1f0ee};
test_output[71:71] = '{32'hc64d847e};
test_input[576:583] = '{32'h40819fd1, 32'hc25edf6c, 32'hc29b7f63, 32'h419e74c1, 32'h4239ef1f, 32'hc2b5ea79, 32'h42c1957b, 32'hc2491c7b};
test_weights[576:583] = '{32'hc2358a14, 32'hc2a1af57, 32'h42762251, 32'h423a7bda, 32'h410115d0, 32'hc2af6626, 32'h417e79ce, 32'hc23ae799};
test_bias[72:72] = '{32'hc290a871};
test_output[72:72] = '{32'h464550dd};
test_input[584:591] = '{32'h3fa479e3, 32'hc1f71272, 32'hc227f0af, 32'h41079be8, 32'hc0122062, 32'h42b8524a, 32'hc23a5040, 32'hc1e85c18};
test_weights[584:591] = '{32'h421e9d9b, 32'hc2a42c61, 32'hc2811cc7, 32'h42ac7f39, 32'hc228abbc, 32'hc26914f5, 32'h41a709c4, 32'h42b4a37a};
test_bias[73:73] = '{32'hc0cd28a3};
test_output[73:73] = '{32'hc5320ba8};
test_input[592:599] = '{32'h413bdd11, 32'hc2a4a86a, 32'hc0c6497b, 32'hc296f3e1, 32'h4185309c, 32'h41e3080a, 32'hc22af278, 32'hc21c4858};
test_weights[592:599] = '{32'h429177f2, 32'h42ad3f60, 32'h41688f46, 32'hc2992f92, 32'hc2bbccf1, 32'hc09a963e, 32'hc22f54b4, 32'h424950c2};
test_bias[74:74] = '{32'hc24c64f9};
test_output[74:74] = '{32'hc517f602};
test_input[600:607] = '{32'h42275fb2, 32'hc28a4a70, 32'hc1525926, 32'hc24b2bbf, 32'hc28ae17e, 32'h42430cab, 32'hc26416c4, 32'h4259851e};
test_weights[600:607] = '{32'hc22b7b41, 32'h42949f3c, 32'hc20fa8a6, 32'h429a36da, 32'h42a34e9f, 32'h41d03a39, 32'h4252644d, 32'h417d1a1a};
test_bias[75:75] = '{32'hc294991e};
test_output[75:75] = '{32'hc684bd31};
test_input[608:615] = '{32'h42966530, 32'hc205031d, 32'hc218d6c3, 32'h42626f5d, 32'h42944b7c, 32'h41342f61, 32'h424364b8, 32'h423879ee};
test_weights[608:615] = '{32'hc1c221a4, 32'hc2abd54c, 32'hc24715fe, 32'hc2591563, 32'h40a5ce46, 32'hc29fc5a4, 32'hc1c9c595, 32'h425d7fbc};
test_bias[76:76] = '{32'hc2a30d9b};
test_output[76:76] = '{32'h4412a54e};
test_input[616:623] = '{32'hc2a5bdeb, 32'h416254c7, 32'hc292f038, 32'h417dc052, 32'hc227e3df, 32'h425d47a5, 32'hc2bfe117, 32'hc14e33f0};
test_weights[616:623] = '{32'hc204eb74, 32'hc2373f24, 32'h42a4f093, 32'hc25fa0b5, 32'hc1a6b545, 32'h42922123, 32'hc19bf987, 32'h42bd3355};
test_bias[77:77] = '{32'hc2c3215a};
test_output[77:77] = '{32'h441d9e17};
test_input[624:631] = '{32'hc2886e4f, 32'hc0f16f31, 32'hc281104e, 32'hc1d2dcae, 32'h423d4143, 32'hc29f088b, 32'hc2c09629, 32'hc28d5298};
test_weights[624:631] = '{32'hc2a76bf4, 32'hc29dcc01, 32'h42c505db, 32'hc277a513, 32'hc2ae349d, 32'hc2a6da09, 32'h424eccbc, 32'h422833ea};
test_bias[78:78] = '{32'h422094d6};
test_output[78:78] = '{32'hc56e89d5};
test_input[632:639] = '{32'hc1b7fb99, 32'hc1d00572, 32'h41a1528d, 32'hc25a8d3f, 32'hc221ff15, 32'h401ac4a2, 32'h4269e5fa, 32'h41401c06};
test_weights[632:639] = '{32'h4286738c, 32'h42a2ea47, 32'h4244763c, 32'h40a3524f, 32'h42a2beac, 32'h42509d3e, 32'hc1917026, 32'hc27ee3d6};
test_bias[79:79] = '{32'hc0a70dc0};
test_output[79:79] = '{32'hc5f89ae3};
test_input[640:647] = '{32'h428f0b58, 32'h4186f4f1, 32'hc1d9ddd6, 32'h4249b2ec, 32'hc2ac9668, 32'hc2bcca23, 32'h41c9791e, 32'h4224584c};
test_weights[640:647] = '{32'h42bee90f, 32'h42a07f66, 32'hc19e6a01, 32'hc233cd54, 32'hc1378a82, 32'hc2b1657e, 32'hc2806ca3, 32'hbf259eae};
test_bias[80:80] = '{32'h429ea4f7};
test_output[80:80] = '{32'h465eaefa};
test_input[648:655] = '{32'hc2888720, 32'h429a37ee, 32'h428ab067, 32'hc1973e6e, 32'h42aa7b59, 32'h42ac66df, 32'hc040c0a5, 32'hc284abe6};
test_weights[648:655] = '{32'hc119b43f, 32'h410515ae, 32'hc0d365c1, 32'h420d78ba, 32'hc15154b7, 32'hc0c54102, 32'hc131b724, 32'hc229845e};
test_bias[81:81] = '{32'h42a3096c};
test_output[81:81] = '{32'h44b541d2};
test_input[656:663] = '{32'h4252db98, 32'h41185946, 32'hc2809df6, 32'hc2444f34, 32'hc2ba2cfa, 32'h420480b9, 32'hc296b0a4, 32'hc211d5d4};
test_weights[656:663] = '{32'h418f1f81, 32'hc2a2778d, 32'hc295909c, 32'hc1e6a89e, 32'hc1765f94, 32'h4280d6c4, 32'h4289f72d, 32'hc2c1a316};
test_bias[82:82] = '{32'hc238fa83};
test_output[82:82] = '{32'h4600dcec};
test_input[664:671] = '{32'h4103bfe3, 32'hc1a4b2f0, 32'h423c452f, 32'hc2701ffa, 32'hc1a6b573, 32'hc22058ea, 32'hc25ea981, 32'hc24a77e1};
test_weights[664:671] = '{32'h42807779, 32'h418d6550, 32'hc279957b, 32'hc1c561f5, 32'h3e15e6ef, 32'hc18806ea, 32'h42a90617, 32'hc2799891};
test_bias[83:83] = '{32'h428926d8};
test_output[83:83] = '{32'hc5029723};
test_input[672:679] = '{32'hc2726809, 32'h429a790a, 32'hc2b0229d, 32'hc23fde84, 32'h42a0d6f8, 32'h4057a4c5, 32'h41edfb04, 32'hc16cb8fa};
test_weights[672:679] = '{32'h428f0a0d, 32'hc282c678, 32'h42aaff02, 32'h42242135, 32'h41d97e4a, 32'hc24f5133, 32'h3fd4d6a5, 32'h415e6c93};
test_bias[84:84] = '{32'hc28a03dd};
test_output[84:84] = '{32'hc6858fae};
test_input[680:687] = '{32'hc189b0a4, 32'hc12e5593, 32'h42a3a062, 32'hc155cac9, 32'h426eb89c, 32'h42046cd7, 32'hc2873b30, 32'hc2811845};
test_weights[680:687] = '{32'h42ad9bd3, 32'h42358feb, 32'h4288c751, 32'h42a9100f, 32'hc2a39def, 32'h4021111c, 32'h424e899d, 32'h42c1742c};
test_bias[85:85] = '{32'h4298ea4d};
test_output[85:85] = '{32'hc63b311c};
test_input[688:695] = '{32'hc19a25aa, 32'h4270c005, 32'h421ea84f, 32'h3e9ba21f, 32'hc22987a0, 32'h41d9037f, 32'h428cb8f6, 32'hc2aaa074};
test_weights[688:695] = '{32'h428f835c, 32'hc13be57d, 32'hc2968893, 32'h42a2c0a1, 32'h429419c5, 32'hc288d398, 32'hc21d18e5, 32'hc2a96891};
test_bias[86:86] = '{32'h411cc6f7};
test_output[86:86] = '{32'hc5ae1c87};
test_input[696:703] = '{32'h4100079a, 32'hc01a8748, 32'h4025a793, 32'h40d8a954, 32'h41c1f472, 32'hc2c4243f, 32'hc283a2aa, 32'hc25dc5ba};
test_weights[696:703] = '{32'h429cf12a, 32'h4215abb8, 32'hc2345029, 32'h4287039b, 32'h429aad8f, 32'h42512641, 32'hc1cbc89c, 32'hc18c2c32};
test_bias[87:87] = '{32'hc2a5e566};
test_output[87:87] = '{32'h433e33f7};
test_input[704:711] = '{32'hc2c368aa, 32'h4254fc23, 32'hc0087019, 32'hc209eb51, 32'hc22dea39, 32'h425421f5, 32'hc286606b, 32'h421f1bd4};
test_weights[704:711] = '{32'hc2c6c333, 32'hc251756f, 32'hc23a4e1f, 32'h429f3815, 32'hc1d69586, 32'h42b502f6, 32'hc2520586, 32'hc201730f};
test_bias[88:88] = '{32'hc214e06a};
test_output[88:88] = '{32'h464275b1};
test_input[712:719] = '{32'hc2ae23df, 32'hc1750783, 32'h42b15c80, 32'h41f0c2de, 32'hc2c6ee19, 32'h42bfd968, 32'h411a8200, 32'h424c90b8};
test_weights[712:719] = '{32'h41c64b63, 32'h42bf2605, 32'h42ac726f, 32'hc24f7536, 32'hc22ad868, 32'hc1b737ea, 32'hc2217312, 32'hc291402d};
test_bias[89:89] = '{32'h41e06304};
test_output[89:89] = '{32'h43db93fe};
test_input[720:727] = '{32'hc27d709c, 32'hc201c95c, 32'h41184bdb, 32'h42a67905, 32'hc2911711, 32'h41015c65, 32'h40e3b142, 32'hc1a7d22a};
test_weights[720:727] = '{32'h3fcb47dc, 32'hc223d44a, 32'h424ff44f, 32'h424864f4, 32'hc28124c7, 32'hc2bb494d, 32'hc2844cce, 32'h42744923};
test_bias[90:90] = '{32'hc25a929c};
test_output[90:90] = '{32'h45fa6fd5};
test_input[728:735] = '{32'hc29fd6a6, 32'h42c7afe5, 32'hc11a8822, 32'h4224709a, 32'hc2c5d4f4, 32'hc2a12a51, 32'hc11216cd, 32'h429e6d0f};
test_weights[728:735] = '{32'hc2117571, 32'h42b60707, 32'hc0f2ee07, 32'hc2235d86, 32'h413c2d37, 32'hc20043a7, 32'hc258a3f9, 32'hc224a0a6};
test_bias[91:91] = '{32'h42ae9ed6};
test_output[91:91] = '{32'h460ea7ef};
test_input[736:743] = '{32'hc298d2c0, 32'hc1189b88, 32'h42b41818, 32'hc25ee94b, 32'hc17adb62, 32'h42281d19, 32'hc1ef142b, 32'h420deabb};
test_weights[736:743] = '{32'h426bf40d, 32'hc29bb442, 32'h4247d2f4, 32'h427170d6, 32'h429eef18, 32'hc2af20ae, 32'h42a31424, 32'hc218bb82};
test_bias[92:92] = '{32'h41284445};
test_output[92:92] = '{32'hc6312517};
test_input[744:751] = '{32'hc180bc52, 32'h42070138, 32'hc171b70b, 32'hc2654a6b, 32'hc2a578e6, 32'h41f7ed36, 32'hc07dcd5f, 32'h42b2b08c};
test_weights[744:751] = '{32'h42bc6411, 32'hc2958e48, 32'h41119a11, 32'h4289a3ed, 32'hc171494d, 32'hc27fcc50, 32'hc22be330, 32'hc286ddeb};
test_bias[93:93] = '{32'hc2b3e9ad};
test_output[93:93] = '{32'hc667425e};
test_input[752:759] = '{32'hc2ba4557, 32'h424d02c7, 32'hc261d6fc, 32'hc28a93e4, 32'h41982a90, 32'h4295831e, 32'hc2b70c24, 32'h425a211f};
test_weights[752:759] = '{32'hc26a360c, 32'hc1eb520f, 32'h41b14834, 32'hc28188ad, 32'hc1f2b1b1, 32'h41eb0669, 32'h42b96983, 32'hc2702299};
test_bias[94:94] = '{32'hc25c79d6};
test_output[94:94] = '{32'hc53c4582};
test_input[760:767] = '{32'hc23789c5, 32'h420eb9e2, 32'h4230c918, 32'hc2570b19, 32'hc2a2ca85, 32'h427b7716, 32'hc2aa765c, 32'hc283d941};
test_weights[760:767] = '{32'hc2a6aa0a, 32'h42786ba7, 32'h41714645, 32'hc28a9f78, 32'hc17323ce, 32'hc2be3b72, 32'hc2430529, 32'hc23ed1a2};
test_bias[95:95] = '{32'hc29210fb};
test_output[95:95] = '{32'h4649d3fc};
test_input[768:775] = '{32'h42adc68f, 32'hc2b61ce2, 32'h41cb0d7b, 32'hc1b4c449, 32'hc2bbb385, 32'hc21247b1, 32'hc1a10aa4, 32'hc19ed553};
test_weights[768:775] = '{32'h427f551c, 32'hc2c4dc6c, 32'hc159ea31, 32'hc2541c1e, 32'h41301e9f, 32'hc2bf08b9, 32'h3fe9358c, 32'hc26a8339};
test_bias[96:96] = '{32'hc1375280};
test_output[96:96] = '{32'h4693f2e1};
test_input[776:783] = '{32'h41a666a7, 32'h41f4cfd6, 32'h41ba7316, 32'h42891759, 32'h429a0a72, 32'hc257186a, 32'h4262b265, 32'hc1f210bc};
test_weights[776:783] = '{32'hc2333987, 32'hc18596ef, 32'h418953fc, 32'h428d32f3, 32'hc2af9faa, 32'hc2886ed1, 32'hc293bb60, 32'h42598bba};
test_bias[97:97] = '{32'hc26b7353};
test_output[97:97] = '{32'hc5a22ba4};
test_input[784:791] = '{32'hc1c07067, 32'hc2c76a7e, 32'hc1ac7e7c, 32'hc232a093, 32'h42b3f5ed, 32'hc0d8adcc, 32'h42c6581a, 32'hc2a44195};
test_weights[784:791] = '{32'hc1aedc48, 32'h421d1523, 32'h41f60882, 32'hc286c2b7, 32'h419c0ae8, 32'hc177e85e, 32'h4240a39d, 32'h400f08fb};
test_bias[98:98] = '{32'h42c19bae};
test_output[98:98] = '{32'h45ac0b6f};
test_input[792:799] = '{32'hc2ad0ff4, 32'h427400aa, 32'hc0c643a4, 32'h42753969, 32'h429a30d5, 32'h4180238f, 32'hc2bea02e, 32'hc2131cbd};
test_weights[792:799] = '{32'h42870dbc, 32'h406fbb9e, 32'hc293a1cb, 32'h411921f9, 32'h4276b02f, 32'hc2a9d218, 32'hc2b5b1d5, 32'h429bd500};
test_bias[99:99] = '{32'hc1265f3d};
test_output[99:99] = '{32'h458ff769};
test_input[800:807] = '{32'hc2a16fa5, 32'hc27b428e, 32'h426bbb1f, 32'h42a0eafb, 32'hc2b376ac, 32'h42895770, 32'hc2c14f06, 32'hc2c2093d};
test_weights[800:807] = '{32'h4263ca08, 32'hc1d1accd, 32'h427b06d4, 32'hc01d4c5a, 32'h42565716, 32'h42ac20e3, 32'h42ab12bd, 32'h41b8b188};
test_bias[100:100] = '{32'hc1f08f60};
test_output[100:100] = '{32'hc60ad4e6};
test_input[808:815] = '{32'h41b882a1, 32'hc289c015, 32'hc11bdd9a, 32'hc2780288, 32'hc26d65e5, 32'hc11a2155, 32'h42c31e9a, 32'hc19f7cdb};
test_weights[808:815] = '{32'hc2346d26, 32'h4276990b, 32'h42b1a88d, 32'hc1ace922, 32'h418a69c0, 32'hc1806b23, 32'hc2b56778, 32'hc2022fc7};
test_bias[101:101] = '{32'hc0e929d4};
test_output[101:101] = '{32'hc6590cc7};
test_input[816:823] = '{32'hc291476a, 32'h42aa4faf, 32'h3ff351dc, 32'hc2a00343, 32'h41f0ead5, 32'h41fe9939, 32'hc28ca144, 32'hc2265b63};
test_weights[816:823] = '{32'hc2b1447c, 32'h42313a2a, 32'hc28b911b, 32'hc271d561, 32'hc2c56817, 32'h40e57909, 32'hc2c06e3c, 32'h413fb690};
test_bias[102:102] = '{32'hc2b0355a};
test_output[102:102] = '{32'h468f5cdd};
test_input[824:831] = '{32'h4250bdb0, 32'h42a9ee72, 32'h414e00aa, 32'hc28af687, 32'hc29e3edb, 32'h429dc2a8, 32'hc114254b, 32'hc28d60d9};
test_weights[824:831] = '{32'h42547f9d, 32'hc26e46fe, 32'h40a4949f, 32'h4288a2db, 32'h4215caf3, 32'h4116de01, 32'h42a5afb6, 32'hc185765d};
test_bias[103:103] = '{32'h42b0ebea};
test_output[103:103] = '{32'hc607c0b8};
test_input[832:839] = '{32'hc1ab62b5, 32'hc24ee5c7, 32'hc1aadafd, 32'h42a97854, 32'h42b43f86, 32'hc299fe0b, 32'hc21dccdc, 32'h42086183};
test_weights[832:839] = '{32'h419a5ff0, 32'h41c8c2c5, 32'h40854974, 32'hc23d11ce, 32'hc0a4eda6, 32'hc29a5b5c, 32'h42817081, 32'h42b18101};
test_bias[104:104] = '{32'h42a7f242};
test_output[104:104] = '{32'h43652692};
test_input[840:847] = '{32'hc23addde, 32'hc2297634, 32'hc112db73, 32'h42a28ee6, 32'h427e8126, 32'hc2307669, 32'hc23f5cb6, 32'h410ca567};
test_weights[840:847] = '{32'hc0c9208b, 32'h4257eadf, 32'h425faf3d, 32'hc2929d72, 32'hc0a7eb20, 32'h42c5d4e2, 32'h4245dbd0, 32'hc168dcfb};
test_bias[105:105] = '{32'h3e8978f8};
test_output[105:105] = '{32'hc674a247};
test_input[848:855] = '{32'h42b40bf9, 32'h42aa027e, 32'h422a0528, 32'hc2184d8c, 32'h418abda4, 32'hc2b2464f, 32'hc2613db0, 32'h42900954};
test_weights[848:855] = '{32'h41c2822e, 32'h426d4d1e, 32'hc1a367c7, 32'h425a609c, 32'hc2b10aec, 32'hc21bd513, 32'h42a40575, 32'h41b4c4da};
test_bias[106:106] = '{32'h40e58fed};
test_output[106:106] = '{32'h454a6b61};
test_input[856:863] = '{32'h4248eea6, 32'hc12345ae, 32'hc2bf98aa, 32'hc187155e, 32'hc174b7d3, 32'h41ae64bb, 32'h4264b10b, 32'hc23b8c29};
test_weights[856:863] = '{32'h42bdac68, 32'hc0defc97, 32'hc05e54f1, 32'h419fa825, 32'hc2643d0b, 32'hc2a21477, 32'h424c99e3, 32'hc27aad5e};
test_bias[107:107] = '{32'hc285c34f};
test_output[107:107] = '{32'h4618137b};
test_input[864:871] = '{32'hc1c1cb7d, 32'h41156c58, 32'h425e8d63, 32'hc22f78ef, 32'hc29d3b8c, 32'hc14dfe66, 32'hc272c9e9, 32'h42639517};
test_weights[864:871] = '{32'hc1a6578b, 32'h42203f96, 32'h422ff25c, 32'hc2c6db23, 32'h426b42db, 32'hc2926f4d, 32'h4231eb1c, 32'hc229c25f};
test_bias[108:108] = '{32'hbf49b78f};
test_output[108:108] = '{32'hc48ab0e2};
test_input[872:879] = '{32'hc1ac3193, 32'h42b80e9e, 32'h4260be57, 32'hc2017217, 32'hc1cf9906, 32'h4193a43e, 32'h424c5562, 32'hc280ca3d};
test_weights[872:879] = '{32'h414b0c84, 32'h42c4b78a, 32'h423e8161, 32'hc2a86822, 32'hc2b8ec89, 32'h429d5815, 32'hc1a0f9cf, 32'hc212fc2f};
test_bias[109:109] = '{32'h429487a6};
test_output[109:109] = '{32'h4697e6d4};
test_input[880:887] = '{32'h42c75ac8, 32'h42837b7a, 32'h424ff914, 32'hc1febdfb, 32'hc18414f0, 32'hc2364d1a, 32'hc2358335, 32'h421c8fbb};
test_weights[880:887] = '{32'h416c48df, 32'hc27ce079, 32'hc18ccc19, 32'hc2c3934d, 32'hc2adaf4d, 32'hc181fe31, 32'h42ab1344, 32'h41dcff51};
test_bias[110:110] = '{32'hc2b83d27};
test_output[110:110] = '{32'hc4966caf};
test_input[888:895] = '{32'h40d12a6b, 32'hc24b4f7e, 32'h427f71c6, 32'h42a4f55e, 32'hc2afe7e7, 32'h421a0934, 32'h4276f274, 32'hc2541fe9};
test_weights[888:895] = '{32'h4283aaf9, 32'h42c16c79, 32'h421c8034, 32'hc27edc1f, 32'hc2c51690, 32'h425aad18, 32'hc283bfc2, 32'hc2a76d72};
test_bias[111:111] = '{32'h41d66e7e};
test_output[111:111] = '{32'h45759f38};
test_input[896:903] = '{32'hbf8ee309, 32'h41d879c2, 32'hc2093cb6, 32'h41f4f1fd, 32'h413718f6, 32'h42651ec6, 32'h42625ec8, 32'hc2b59bfa};
test_weights[896:903] = '{32'h4178e033, 32'h425bb21b, 32'h41ac28e3, 32'h421420e4, 32'h42afee8a, 32'hbf1dc8f7, 32'h4270d618, 32'hc20f494a};
test_bias[112:112] = '{32'hc256d814};
test_output[112:112] = '{32'h46138899};
test_input[904:911] = '{32'hc27cc315, 32'h42b9815d, 32'h42bc37e7, 32'h420ff69d, 32'hc2aa2c6d, 32'hc2186ce2, 32'hc2c20a41, 32'hc29e7031};
test_weights[904:911] = '{32'h423d224c, 32'h4225fa0c, 32'h42b5bfbd, 32'hc2834897, 32'h4247f4af, 32'h418f45b7, 32'h414f666e, 32'hc291378b};
test_bias[113:113] = '{32'hc2a6a44c};
test_output[113:113] = '{32'h45cbed20};
test_input[912:919] = '{32'hc1729065, 32'h41268ed8, 32'hc2b50dad, 32'hc2a49d01, 32'hc2be2dd9, 32'hc25ac5a4, 32'hc25245ac, 32'h4128e1e7};
test_weights[912:919] = '{32'hc244f5c5, 32'hc27d08e1, 32'h42478a2f, 32'h42417073, 32'h41d969f5, 32'hc10a5519, 32'hc1841497, 32'h4255d2e3};
test_bias[114:114] = '{32'h41d45d95};
test_output[114:114] = '{32'hc60d93d3};
test_input[920:927] = '{32'hc26e0db6, 32'h4296273a, 32'hc2c05189, 32'hc219685a, 32'hc282b8c2, 32'h4151085c, 32'hc2c59237, 32'hc1c7b8dd};
test_weights[920:927] = '{32'hc2811e2c, 32'hc2bedcde, 32'h42bc1c48, 32'hc0be1fd2, 32'h4105125b, 32'h428968b8, 32'h4262e617, 32'h4216180d};
test_bias[115:115] = '{32'hc2248b6e};
test_output[115:115] = '{32'hc68f7cf4};
test_input[928:935] = '{32'h4294a312, 32'h429bab2d, 32'h4132994f, 32'hc20af4ce, 32'hc1c11420, 32'hbf968db1, 32'h41d4743b, 32'h4220beab};
test_weights[928:935] = '{32'hc290a6a4, 32'hc22931cd, 32'hc292c2fb, 32'hc28dda6a, 32'h42af362b, 32'hc1c99bbc, 32'h4269bfd4, 32'h42064953};
test_bias[116:116] = '{32'hc2adb25a};
test_output[116:116] = '{32'hc5c4a904};
test_input[936:943] = '{32'h4285a404, 32'h42ab9719, 32'h4287e874, 32'hc2841475, 32'h41e15b23, 32'hc2830bef, 32'hc2ba5b62, 32'h419a2e9e};
test_weights[936:943] = '{32'hc164e908, 32'h4189ea24, 32'hc2702a2c, 32'h41dc0269, 32'h4221000a, 32'hc2468a55, 32'hc27b8c9f, 32'h40a705c8};
test_bias[117:117] = '{32'h41ee6a82};
test_output[117:117] = '{32'h459c587f};
test_input[944:951] = '{32'h42bbacf1, 32'h42249a77, 32'h42918716, 32'hc195d730, 32'h4295c165, 32'h42c29820, 32'h413fe156, 32'hc1b202c8};
test_weights[944:951] = '{32'h41fa5f11, 32'h429661c2, 32'hc1bf610f, 32'hc28357f3, 32'hc21fe920, 32'hc1a6328c, 32'h428e09d8, 32'hc0fa76d2};
test_bias[118:118] = '{32'hc2b258b5};
test_output[118:118] = '{32'h44b447c8};
test_input[952:959] = '{32'h42aa0afd, 32'hc275d7b7, 32'hc1e13177, 32'h4278c71a, 32'hc11f63a5, 32'hc27d6ea3, 32'hc2a8ba39, 32'h40071f9b};
test_weights[952:959] = '{32'hc274dca0, 32'hc196cee7, 32'hc2984f53, 32'hc1f545b1, 32'h42c5f191, 32'h42b6d5ba, 32'h42a906ee, 32'hbfa47a85};
test_bias[119:119] = '{32'hc2c0a499};
test_output[119:119] = '{32'hc68b3012};
test_input[960:967] = '{32'hc29ccab7, 32'h4284c5e0, 32'h41f13bef, 32'hc27a92d1, 32'hc16785c6, 32'hc26b7d0b, 32'hc21d1f39, 32'hc2a96f8b};
test_weights[960:967] = '{32'h4291c5bd, 32'hc1fe7844, 32'hc229c258, 32'h428a1259, 32'hbff37b14, 32'h426bfea2, 32'hc2a26b02, 32'hc0dfc209};
test_bias[120:120] = '{32'h42c1a1a3};
test_output[120:120] = '{32'hc64b1302};
test_input[968:975] = '{32'h42aab00c, 32'hc1873da9, 32'h4293259b, 32'h42869845, 32'h41e2962d, 32'hc188f262, 32'h3f2fe29a, 32'h42616529};
test_weights[968:975] = '{32'h40b42e2f, 32'hc26d9742, 32'hc2b2502b, 32'h41fd90f9, 32'h422205e1, 32'h40147669, 32'hc0e4238e, 32'h421b26c4};
test_bias[121:121] = '{32'h4084b852};
test_output[121:121] = '{32'h43af4c93};
test_input[976:983] = '{32'h42083264, 32'hc229a741, 32'hc2c740b9, 32'h41eb5944, 32'hc015db87, 32'h423482a9, 32'hc23cbe12, 32'h412d3911};
test_weights[976:983] = '{32'hc20e8090, 32'hc28c06c8, 32'hc22730cf, 32'hc29f9e64, 32'hc2866a43, 32'h4280e6a7, 32'h42590f65, 32'h4085cbda};
test_bias[122:122] = '{32'h4204de6a};
test_output[122:122] = '{32'h4581e485};
test_input[984:991] = '{32'hc24edc1f, 32'h3fba26d7, 32'h42b2ac4b, 32'hc2bfc1c6, 32'hc2015f2b, 32'hc2aaa3f2, 32'h40ad2f51, 32'h428e9ebe};
test_weights[984:991] = '{32'hc291120b, 32'hc226512d, 32'hc003ad26, 32'hc28311a8, 32'hc2a1a647, 32'hc2514cd3, 32'hc234d7f9, 32'hc2afab77};
test_bias[123:123] = '{32'h42aba327};
test_output[123:123] = '{32'h46233963};
test_input[992:999] = '{32'h429c1d22, 32'h42494624, 32'hc20f786a, 32'h41eb8eed, 32'h40fde706, 32'h426c98cf, 32'hc2a20f4b, 32'h429365be};
test_weights[992:999] = '{32'hc146ddb3, 32'hc2962d23, 32'hc2b9a579, 32'h42b1f463, 32'hc187c162, 32'h405879fb, 32'hc26974f5, 32'h41f476a6};
test_bias[124:124] = '{32'h42423b65};
test_output[124:124] = '{32'h4601a047};
test_input[1000:1007] = '{32'hc2b33b15, 32'h4266c37b, 32'hc29e1bf6, 32'hc2b18b92, 32'h42062200, 32'hc222ce3b, 32'hc2ae6848, 32'h421e0e3f};
test_weights[1000:1007] = '{32'hc1918190, 32'hc2a4e81c, 32'h42c425ce, 32'hc278088c, 32'hc128e122, 32'hc25e11ba, 32'h41efa9ce, 32'hc2824bd3};
test_bias[125:125] = '{32'hc2986301};
test_output[125:125] = '{32'hc608726c};
test_input[1008:1015] = '{32'hc278731f, 32'hc29032e8, 32'h428320f3, 32'hc25c2671, 32'hc20bf4d2, 32'h421b6ade, 32'h4223bbf0, 32'h42160e84};
test_weights[1008:1015] = '{32'h423d02b7, 32'hc210fe6d, 32'h42351ab6, 32'hc1c77629, 32'hc28bb254, 32'h42c30647, 32'h42afca43, 32'h417916a6};
test_bias[126:126] = '{32'h42880e7e};
test_output[126:126] = '{32'h4662976e};
test_input[1016:1023] = '{32'hc2c0f42f, 32'h42ac80d9, 32'hc2c7c168, 32'hc28d3a58, 32'h41d02753, 32'hc1c08f9d, 32'h4284cd9c, 32'h42adcd61};
test_weights[1016:1023] = '{32'hc294a06e, 32'h4189a176, 32'h4213635b, 32'h42946e73, 32'hc2080b78, 32'h42a33220, 32'hc2c2aec2, 32'h42ae0627};
test_bias[127:127] = '{32'hc1b3a18a};
test_output[127:127] = '{32'hc4ff2415};
test_input[1024:1031] = '{32'hc26275b3, 32'hc0eeceb5, 32'h4233a616, 32'hc2bfe13d, 32'hc26f2711, 32'hc1ce0f2e, 32'hc2884581, 32'hc0ebef9c};
test_weights[1024:1031] = '{32'hc2b8adce, 32'h427c3c35, 32'h4278a17d, 32'h4221a91f, 32'h4268376e, 32'hc298ab92, 32'hc23f9854, 32'h42bf5b70};
test_bias[128:128] = '{32'hc1f01006};
test_output[128:128] = '{32'h4592b6a6};
test_input[1032:1039] = '{32'hc19062f8, 32'hc23f4d2e, 32'h41d4337f, 32'hc1e60047, 32'h4208cbb5, 32'hc2aad437, 32'h42b8ceff, 32'hc0af092e};
test_weights[1032:1039] = '{32'hc28de9c0, 32'hc2c3aa01, 32'h41dda082, 32'hc259dcf0, 32'hc2595ed9, 32'hc2811c7e, 32'h4111e58e, 32'h40d3d4f4};
test_bias[129:129] = '{32'hc2ad2a0c};
test_output[129:129] = '{32'h46456e40};
test_input[1040:1047] = '{32'hc29610dd, 32'h40d25550, 32'hc2756e08, 32'hc29b8118, 32'hc2b47da3, 32'h4146e48a, 32'h42935337, 32'hc2a8a533};
test_weights[1040:1047] = '{32'hc25dc578, 32'hc11fdfed, 32'h42a2ceea, 32'hc283cfa4, 32'h429bc0fa, 32'h41646e41, 32'h4226d3e6, 32'h42a121a0};
test_bias[130:130] = '{32'h3e9c6dae};
test_output[130:130] = '{32'hc5c65cf0};
test_input[1048:1055] = '{32'h4227138c, 32'h41edc49c, 32'hc2b7a01c, 32'hc2ac7aea, 32'hc261554d, 32'hc2b43b28, 32'hc27037b1, 32'h42ae82f7};
test_weights[1048:1055] = '{32'hc0cd252e, 32'h4245fa98, 32'h4231c749, 32'hc25e9465, 32'hc2b8535f, 32'h42858370, 32'hc2c531ad, 32'h41085227};
test_bias[131:131] = '{32'hc267ed3c};
test_output[131:131] = '{32'h45f0c12c};
test_input[1056:1063] = '{32'h41b5eda2, 32'hc2354326, 32'hc27ec864, 32'hc26112b1, 32'h42387ecd, 32'h4295a4b8, 32'hc239bb0c, 32'h42804694};
test_weights[1056:1063] = '{32'hc29503be, 32'h42234803, 32'h42bd0db1, 32'hc201ee73, 32'hc12d5001, 32'hc1337602, 32'hc25c875a, 32'hc2af5cb7};
test_bias[132:132] = '{32'hc2b8f24a};
test_output[132:132] = '{32'hc63f21aa};
test_input[1064:1071] = '{32'hc29f9aec, 32'h40ed73d7, 32'h42c6664c, 32'h423891c5, 32'hc1ef7c23, 32'hc2b95beb, 32'h42ad81db, 32'h42a0b6da};
test_weights[1064:1071] = '{32'h423fd061, 32'hc26acf23, 32'h42c7cf0a, 32'hc2746520, 32'hc1f2c5eb, 32'hc2557693, 32'hc0525a8e, 32'h42c4f736};
test_bias[133:133] = '{32'h42c6d1de};
test_output[133:133] = '{32'h4680368e};
test_input[1072:1079] = '{32'h40b01d42, 32'h42b7090c, 32'hc282a2bf, 32'hc2509b77, 32'hc0b381d2, 32'hc21da48f, 32'hc25adbb5, 32'hbf42c26d};
test_weights[1072:1079] = '{32'h423d585d, 32'h42c18448, 32'hbfc54e23, 32'hc23a6a75, 32'h415cabfb, 32'hc2b19fbb, 32'hc148d0d5, 32'hbe9928f0};
test_bias[134:134] = '{32'hc281558f};
test_output[134:134] = '{32'h46752f5d};
test_input[1080:1087] = '{32'hc1acd09c, 32'hc22b0b44, 32'h42056e23, 32'hc1cabb7e, 32'hc2b74d38, 32'h413128e6, 32'hc16c3c13, 32'h42ac7f9e};
test_weights[1080:1087] = '{32'h42185f7e, 32'h424aedc0, 32'h3fb425fb, 32'hc081eb9f, 32'h410ef7f1, 32'hbfa8ff03, 32'h42c63813, 32'h42c106f7};
test_bias[135:135] = '{32'hc23dad96};
test_output[135:135] = '{32'h4544182e};
test_input[1088:1095] = '{32'hc278c60e, 32'h42b200f2, 32'hc244a9f9, 32'h3e9428c8, 32'hc2a21f0d, 32'hc2a80431, 32'h42a60b7e, 32'hc1d2a2b6};
test_weights[1088:1095] = '{32'hc2a42202, 32'h419d0a1d, 32'h4181b801, 32'hc258939e, 32'hc12c4ea0, 32'h41fa1e14, 32'h4106e510, 32'hc24573c0};
test_bias[136:136] = '{32'h426dc179};
test_output[136:136] = '{32'h45c63e28};
test_input[1096:1103] = '{32'hc21fc5f1, 32'hc2b76533, 32'hc1825d80, 32'h42b872e0, 32'h424721f1, 32'hc2b3687f, 32'h410a9956, 32'h42a0d927};
test_weights[1096:1103] = '{32'h4087c355, 32'hc28d71b2, 32'hc125ebb6, 32'h41eff0d0, 32'h4214d242, 32'h41cb0645, 32'hc22294ad, 32'h4279ea99};
test_bias[137:137] = '{32'hc14654e1};
test_output[137:137] = '{32'h4652ba95};
test_input[1104:1111] = '{32'h4292ba48, 32'hc1c0e0e9, 32'h42611496, 32'hc2728a05, 32'h4288335e, 32'h42b8d598, 32'h42a680e5, 32'hc1e5941c};
test_weights[1104:1111] = '{32'h420e43f7, 32'h4237d698, 32'hc28d6452, 32'hc28c04a9, 32'h426cdc08, 32'h4196259b, 32'hc199ca5d, 32'h40ccf395};
test_bias[138:138] = '{32'h42a6c49a};
test_output[138:138] = '{32'h45b652f3};
test_input[1112:1119] = '{32'hc2bedecf, 32'hc29e6454, 32'hc14bb8ec, 32'hc1eff1af, 32'hc2b6f87c, 32'hc28e6873, 32'hc28de2aa, 32'h429d66e9};
test_weights[1112:1119] = '{32'hc1e2bb8e, 32'hc2393917, 32'h422bb693, 32'h428db05a, 32'hc282734d, 32'hc19fe1ca, 32'hc16ee3a2, 32'hc0c06d9a};
test_bias[139:139] = '{32'h42616744};
test_output[139:139] = '{32'h46375445};
test_input[1120:1127] = '{32'hc2492f53, 32'hc29e7427, 32'hc2765ec7, 32'hc22edef6, 32'hc292d136, 32'h42bfd126, 32'h42b6976a, 32'h42c44c7e};
test_weights[1120:1127] = '{32'hc21fb068, 32'hc1e51c54, 32'h428ec62f, 32'hc22fae40, 32'hc248011e, 32'h4163c778, 32'hc1468c29, 32'hc2849dd5};
test_bias[140:140] = '{32'h42122f27};
test_output[140:140] = '{32'hc44020e9};
test_input[1128:1135] = '{32'h41de4160, 32'hc220fbce, 32'h4204c1eb, 32'h4187c975, 32'h4291c519, 32'h42844d57, 32'hc25602f9, 32'h41d1fef5};
test_weights[1128:1135] = '{32'hc2ba08af, 32'hc2ae84fb, 32'hc08fc4fc, 32'hc2109188, 32'hc119b136, 32'h429041f1, 32'h417f12dc, 32'h41570d8a};
test_bias[141:141] = '{32'h42b97cd2};
test_output[141:141] = '{32'h456f4fab};
test_input[1136:1143] = '{32'h42b62fda, 32'hbfab799f, 32'h4115593b, 32'h4256cea7, 32'h3f1a4290, 32'hc270d14d, 32'hc0d11f28, 32'h3f2c1a55};
test_weights[1136:1143] = '{32'h42a58f09, 32'h42762c3a, 32'h42a50b16, 32'hc2a08a07, 32'h427bef7a, 32'h421cfb01, 32'h42bdcf0f, 32'hc23a4054};
test_bias[142:142] = '{32'h4283fd30};
test_output[142:142] = '{32'h447be52f};
test_input[1144:1151] = '{32'hc073c438, 32'hc26a9ddd, 32'h40d0752d, 32'h4257288f, 32'hc27e95bb, 32'hc27c7261, 32'hc280f513, 32'h4191b952};
test_weights[1144:1151] = '{32'hc2c30911, 32'hc27ee0cf, 32'hc09d5dab, 32'hc2a7987d, 32'h42ab9b3e, 32'h420c5894, 32'h41ee5b93, 32'hc2911163};
test_bias[143:143] = '{32'h42453b94};
test_output[143:143] = '{32'hc6308c77};
test_input[1152:1159] = '{32'hc1d910ae, 32'h41f5781d, 32'h42bbf2e5, 32'h42c7792f, 32'h4246aa75, 32'hc2ba8e32, 32'hc0af8b68, 32'hc25d8282};
test_weights[1152:1159] = '{32'h429830f1, 32'hc20e09e6, 32'hc260fb5a, 32'h41a333bb, 32'hc2a1f9aa, 32'h41b30219, 32'h421f8185, 32'h420c3312};
test_bias[144:144] = '{32'h4221e198};
test_output[144:144] = '{32'hc664a844};
test_input[1160:1167] = '{32'h424e5c71, 32'h42beab5f, 32'h42bef077, 32'h3fdbaf5b, 32'hc2510a7d, 32'h4113d8ae, 32'hc23577f1, 32'h41be74c0};
test_weights[1160:1167] = '{32'h426705c4, 32'hc14a63c0, 32'hc252a4ae, 32'h42376800, 32'h42493127, 32'h423de273, 32'hc20c7371, 32'h41307efd};
test_bias[145:145] = '{32'h42b93f2e};
test_output[145:145] = '{32'hc5558d72};
test_input[1168:1175] = '{32'h4299f009, 32'h429918d1, 32'hc2963919, 32'hc289a12e, 32'hc21c4c02, 32'hc2398d0f, 32'h42400806, 32'h42449452};
test_weights[1168:1175] = '{32'h41f370ae, 32'h428010e4, 32'hc247aecc, 32'h426a0513, 32'h4241789a, 32'h41bc990d, 32'h42ab2563, 32'hc22d2280};
test_bias[146:146] = '{32'hc2b58dd5};
test_output[146:146] = '{32'h45b790f4};
test_input[1176:1183] = '{32'hc18b1966, 32'h427039b0, 32'hc27a2f6d, 32'hc2a7e030, 32'h428a3dd2, 32'hc242ca85, 32'h42854950, 32'h4278911c};
test_weights[1176:1183] = '{32'hc226d1ed, 32'h423adc33, 32'h4238b054, 32'hbee2cd85, 32'hc186c548, 32'hc29d5a7d, 32'h429068e0, 32'h4280fe19};
test_bias[147:147] = '{32'hc262224a};
test_output[147:147] = '{32'h463d38fa};
test_input[1184:1191] = '{32'hc290fa78, 32'h424e10c2, 32'h4213a0c3, 32'h41ba97dc, 32'h42be79a4, 32'h42af8836, 32'hc0e7dff8, 32'h42b3d8b8};
test_weights[1184:1191] = '{32'hc23368fd, 32'h4192581d, 32'hc2414cd6, 32'h41eea1df, 32'h40bd15c5, 32'h41b18c4c, 32'hc2a1b6ed, 32'hbdfbc1ef};
test_bias[148:148] = '{32'h425bff18};
test_output[148:148] = '{32'h45c332cb};
test_input[1192:1199] = '{32'hc2513e51, 32'hc21655b3, 32'h42bc5894, 32'hc18916ae, 32'h429dcccf, 32'hc2bc2ead, 32'h427b099f, 32'h3f149c65};
test_weights[1192:1199] = '{32'hc2a7d642, 32'hc2bfff71, 32'h428b45f0, 32'hc164da42, 32'h42aa1a29, 32'hc258f88a, 32'hc1c2628b, 32'h42514abd};
test_bias[149:149] = '{32'hc21e3a56};
test_output[149:149] = '{32'h46c3f203};
test_input[1200:1207] = '{32'h421e34b8, 32'hc2a89a9f, 32'h428de544, 32'hc2b48eb3, 32'hc24b9735, 32'h412b0baa, 32'h427c32c6, 32'h42965b3d};
test_weights[1200:1207] = '{32'h410d1fe5, 32'h4110624b, 32'h420c9f04, 32'hc2a9a132, 32'h42745a47, 32'h42c5c00d, 32'h428e87ef, 32'h42b6661e};
test_bias[150:150] = '{32'hc1ae25ae};
test_output[150:150] = '{32'h46948d7e};
test_input[1208:1215] = '{32'hc18223fb, 32'h419675cc, 32'hc2418170, 32'h425e8116, 32'h414f8d14, 32'hc2b8f2c6, 32'hc25dac75, 32'h42330bea};
test_weights[1208:1215] = '{32'hc2ac66c0, 32'h4299f6f0, 32'hc1e41e77, 32'hc2887fb5, 32'h42bbfdbf, 32'hc2bf6e82, 32'hc29ef00e, 32'hc299e005};
test_bias[151:151] = '{32'hc2aa42e7};
test_output[151:151] = '{32'h4631cae9};
test_input[1216:1223] = '{32'hc21f2b55, 32'h418663c5, 32'h3f1869b4, 32'hc21a518c, 32'hc2a66a3c, 32'hc2124310, 32'h42b247b5, 32'h42c32027};
test_weights[1216:1223] = '{32'h4089b4cc, 32'hc29e5784, 32'hc1a1dc4b, 32'hc2aed40b, 32'h427bab57, 32'hc19ea53e, 32'h41c6ed32, 32'hc2339c5d};
test_bias[152:152] = '{32'hc298fd59};
test_output[152:152] = '{32'hc598ddaf};
test_input[1224:1231] = '{32'hc2a66565, 32'h4144628b, 32'hc10bad54, 32'h42bf055a, 32'h4278a2c9, 32'h42c2e9a0, 32'hc2bb8319, 32'hc281f2e4};
test_weights[1224:1231] = '{32'hc2b7fed7, 32'h424527ef, 32'h429f3baa, 32'hc2813791, 32'h413213b1, 32'h42b8e08b, 32'hc2786eec, 32'h428a7b00};
test_bias[153:153] = '{32'hc1e4601d};
test_output[153:153] = '{32'h4641956e};
test_input[1232:1239] = '{32'h42c62b41, 32'hc16ca5e7, 32'h426d4eee, 32'h41efc6c4, 32'h41d3e2d7, 32'hc255c5e8, 32'h414b048b, 32'hc2714e9e};
test_weights[1232:1239] = '{32'h41acba92, 32'hc29db834, 32'hc209bd23, 32'hc1e88ef5, 32'hbf381391, 32'hc1704197, 32'h429e52d1, 32'hc28bce87};
test_bias[154:154] = '{32'h41bfbc3a};
test_output[154:154] = '{32'h45c8a39c};
test_input[1240:1247] = '{32'hc29a44c9, 32'hc2a651b6, 32'h413d727f, 32'hc245c543, 32'h4236491c, 32'h41cc16b1, 32'h424dae17, 32'h41c1782c};
test_weights[1240:1247] = '{32'h42ae04f4, 32'h425f0ceb, 32'hc2ad890c, 32'h4254a086, 32'hc0826bd2, 32'hc1b402e2, 32'hc2172ce0, 32'hc1b5c1f3};
test_bias[155:155] = '{32'hc1919ffd};
test_output[155:155] = '{32'hc68ec5f9};
test_input[1248:1255] = '{32'h424ea107, 32'h42742c7e, 32'h421209a7, 32'h40b7f952, 32'h425aeb35, 32'hc2acda5a, 32'h42c7d07d, 32'h42a3c36c};
test_weights[1248:1255] = '{32'h413728ab, 32'h40f5c484, 32'hc29cbd27, 32'h41d4b636, 32'h42a33d53, 32'hc28645c0, 32'h42a0d70a, 32'h41ceb41c};
test_bias[156:156] = '{32'h413ea6b2};
test_output[156:156] = '{32'h4692be96};
test_input[1256:1263] = '{32'hc22277ee, 32'h42af79f0, 32'h4160cfcf, 32'hc1a4a522, 32'h4286cce5, 32'h41474471, 32'h42a6586f, 32'hc2af6927};
test_weights[1256:1263] = '{32'h428ae7e8, 32'hc26e330b, 32'hc2b17fdd, 32'hc2c52505, 32'h424fa415, 32'h42900ec3, 32'h42be6199, 32'hc1a6858f};
test_bias[157:157] = '{32'h427860cf};
test_output[157:157] = '{32'h45d8c58d};
test_input[1264:1271] = '{32'h42c435c9, 32'h4075214b, 32'hc29189b3, 32'h417e4640, 32'hc1980c48, 32'hc1e58f54, 32'h42b699ef, 32'hc28fa39f};
test_weights[1264:1271] = '{32'h40ee8156, 32'h4137c91e, 32'hc291af87, 32'hc2a3512f, 32'hc2b4486e, 32'h4292db7f, 32'hc2ab6c3e, 32'h42bc3031};
test_bias[158:158] = '{32'h3fb7f3d4};
test_output[158:158] = '{32'hc61f560b};
test_input[1272:1279] = '{32'h42a56475, 32'hc186be34, 32'h420d9733, 32'hc2008ee7, 32'hc2bb2332, 32'hc1ff70e7, 32'h42bed684, 32'h429949c0};
test_weights[1272:1279] = '{32'h419553c3, 32'h42234bad, 32'h42be6f65, 32'h40c2392c, 32'hc20ceeeb, 32'hc239dd04, 32'h4200fb2d, 32'hc1db4469};
test_bias[159:159] = '{32'h41d83e70};
test_output[159:159] = '{32'h46195bdc};
test_input[1280:1287] = '{32'h42a47a8b, 32'hc2bdb1d0, 32'h4258d044, 32'hc18ded57, 32'hc2711ba8, 32'hc12543dc, 32'hc2b0c72c, 32'hc2454c23};
test_weights[1280:1287] = '{32'hc260b02a, 32'hc2b3ee33, 32'h41c86b5c, 32'hc28042aa, 32'hc1601461, 32'hc1a4febf, 32'hc29b02cb, 32'hc23125db};
test_bias[160:160] = '{32'hc2bebbb9};
test_output[160:160] = '{32'h46802beb};
test_input[1288:1295] = '{32'h426e7616, 32'h42585e38, 32'hc213e12c, 32'h420d1920, 32'h411d4d12, 32'h4287828b, 32'hc16e2c4a, 32'hc24ca9bc};
test_weights[1288:1295] = '{32'hc124798d, 32'hc24a8aea, 32'hc1de3228, 32'hc25cedd2, 32'hc275c6b4, 32'hc22bb9cc, 32'hc2837044, 32'h424f421e};
test_bias[161:161] = '{32'hc2a49d33};
test_output[161:161] = '{32'hc6151553};
test_input[1296:1303] = '{32'hc16c71ec, 32'h415c7953, 32'h4266d084, 32'h422d5540, 32'hc18a0960, 32'h420bfc21, 32'h412e8299, 32'hc2805944};
test_weights[1296:1303] = '{32'hc26c3f8a, 32'h4295b0b4, 32'h420b86c3, 32'h406ec782, 32'h41dbb9ff, 32'h4272a2b4, 32'h429a1a45, 32'hc28f6ff8};
test_bias[162:162] = '{32'h42b86687};
test_output[162:162] = '{32'h462ffa80};
test_input[1304:1311] = '{32'h41cb9304, 32'hc1ab754c, 32'h403edac7, 32'h42344d15, 32'hc29f641e, 32'h4274a9ad, 32'h4266e228, 32'h41eb32ce};
test_weights[1304:1311] = '{32'h42423904, 32'h42096755, 32'h4298628c, 32'h419640ba, 32'h42c66042, 32'hc2123323, 32'hc28faba8, 32'h4221e984};
test_bias[163:163] = '{32'h41ea1e9b};
test_output[163:163] = '{32'hc633996f};
test_input[1312:1319] = '{32'h421c58b9, 32'hc213030d, 32'h4259b65a, 32'hc2a1f7d6, 32'hc12fe606, 32'h42740521, 32'hc1a07cce, 32'hc2c075d4};
test_weights[1312:1319] = '{32'h4294530b, 32'h41ac4f13, 32'h418cfd0f, 32'h4243985d, 32'hc2b7c0e5, 32'hc2133b81, 32'h425e544d, 32'h428c1748};
test_bias[164:164] = '{32'hc2be3f0d};
test_output[164:164] = '{32'hc61d7ee3};
test_input[1320:1327] = '{32'h4278bf79, 32'h42840346, 32'h42490fdd, 32'h4286f1ce, 32'h428135d5, 32'hc27c3911, 32'hc20962f0, 32'h41505f4b};
test_weights[1320:1327] = '{32'h42b77cdd, 32'h428f3543, 32'h40713fe2, 32'h42b608fd, 32'h41903f02, 32'h42bf9428, 32'hc2979cf0, 32'h40561ba7};
test_bias[165:165] = '{32'h41ced33a};
test_output[165:165] = '{32'h466380ac};
test_input[1328:1335] = '{32'hc2499be5, 32'hc1d21b82, 32'h42808898, 32'h40f6bbe5, 32'hc1656635, 32'hc286b6a6, 32'h41f60258, 32'hc2ae40cb};
test_weights[1328:1335] = '{32'h421f9cbb, 32'hc0d24ffb, 32'hc283d969, 32'hc14e73a1, 32'hc28d361c, 32'hc288138f, 32'h427e11c9, 32'hbfef1b4f};
test_bias[166:166] = '{32'h4276669f};
test_output[166:166] = '{32'h44c7bc07};
test_input[1336:1343] = '{32'h41ffa159, 32'hc286a35c, 32'h42876c65, 32'hc2a34e05, 32'h42972df9, 32'hc2a7dc58, 32'hc260d185, 32'hc1e21032};
test_weights[1336:1343] = '{32'h41d04e3e, 32'h429be11d, 32'hc23bbd52, 32'h4286ac14, 32'hc2b6b6ef, 32'h41a56976, 32'h4215bb71, 32'hc230c72b};
test_bias[167:167] = '{32'hc262674e};
test_output[167:167] = '{32'hc6b0e776};
test_input[1344:1351] = '{32'h4261c744, 32'hc23f76b6, 32'h414b54d7, 32'h42899d4b, 32'h41eb041b, 32'hc0e8d9b9, 32'h429a78ec, 32'h42958448};
test_weights[1344:1351] = '{32'hc23f9551, 32'hc2a23dcc, 32'h402e19bf, 32'hc1cc1bee, 32'h42851faf, 32'h4241d0c2, 32'h4200fa06, 32'hc24b57e1};
test_bias[168:168] = '{32'hc2b4b232};
test_output[168:168] = '{32'hc3a98268};
test_input[1352:1359] = '{32'h4258f895, 32'hc0a25787, 32'h4299c17b, 32'hc2bb6b67, 32'hc211b860, 32'h426f6afd, 32'hc272066e, 32'h42101898};
test_weights[1352:1359] = '{32'hc2085c82, 32'h42a3f5f6, 32'hc28637c8, 32'hc20a56a4, 32'hc16ea51d, 32'hc28e497d, 32'h42b23634, 32'h422e4eee};
test_bias[169:169] = '{32'hc0d5b67a};
test_output[169:169] = '{32'hc6373a32};
test_input[1360:1367] = '{32'hc2411182, 32'hc24d77e4, 32'hc2177b75, 32'hc25c5be7, 32'hc2078994, 32'h421a60a6, 32'hc21aacc6, 32'h42657046};
test_weights[1360:1367] = '{32'hc1d352ec, 32'hc09ae00e, 32'h4250976e, 32'h4290846c, 32'h424b5440, 32'h41ea5c4b, 32'hc2b7ddd3, 32'h4214186f};
test_bias[170:170] = '{32'hc1e89de9};
test_output[170:170] = '{32'h441c7193};
test_input[1368:1375] = '{32'h417f0009, 32'hc2c53e9e, 32'hc27fca7c, 32'h4251aac6, 32'hc0d6a011, 32'hc2859baa, 32'h42173949, 32'hc2ab115e};
test_weights[1368:1375] = '{32'hc2733b06, 32'hc2b7a4de, 32'h4286901d, 32'hc1a7c11d, 32'hbf92d40a, 32'h42a597ba, 32'hc29accf7, 32'hc1e67d74};
test_bias[171:171] = '{32'h41931dc9};
test_output[171:171] = '{32'hc54d1f6c};
test_input[1376:1383] = '{32'h42b57f61, 32'hc29d5ae8, 32'hc205b845, 32'hc2b95ed2, 32'hc1cb7dc7, 32'h42071224, 32'hc202545e, 32'hc2aa9286};
test_weights[1376:1383] = '{32'h42481bae, 32'h42be8a22, 32'hc29c83d4, 32'hc2718600, 32'hc29e1816, 32'h4285ecf7, 32'h416af30b, 32'hc2b5241c};
test_bias[172:172] = '{32'h42239dbd};
test_output[172:172] = '{32'h46835f27};
test_input[1384:1391] = '{32'h4113623b, 32'h418db1ba, 32'hc1e20929, 32'hc2a0b3a7, 32'h421dba93, 32'h42986233, 32'h42980067, 32'h42bdd45b};
test_weights[1384:1391] = '{32'h4287c9b0, 32'h41905d2e, 32'h41a8316b, 32'h429db1c9, 32'hc157bbeb, 32'hc2321e8e, 32'h4223f200, 32'hc2751d1c};
test_bias[173:173] = '{32'h4171fe69};
test_output[173:173] = '{32'hc644cc2f};
test_input[1392:1399] = '{32'h42a486cf, 32'hc2c4b737, 32'hc2196476, 32'hc2be676b, 32'hbf05a2c6, 32'hc12965a3, 32'hc2903f8b, 32'h42b92f40};
test_weights[1392:1399] = '{32'hc2b54f5e, 32'h427cf05d, 32'h42436600, 32'hc2c4625a, 32'h4292ba6d, 32'hc28a88e2, 32'h41f31088, 32'h41de7833};
test_bias[174:174] = '{32'hc2b04a71};
test_output[174:174] = '{32'hc5a2dfe9};
test_input[1400:1407] = '{32'h423d6907, 32'hc23d77d4, 32'hc1a7aa1a, 32'hc2a6f61a, 32'h424d3db4, 32'hc03ec76e, 32'hc260abda, 32'hc190ac28};
test_weights[1400:1407] = '{32'hc209a546, 32'h42c41b31, 32'hc217976e, 32'h4160b4ed, 32'h413de9ba, 32'h42a4efdd, 32'hc255108e, 32'hc2a205ad};
test_bias[175:175] = '{32'h42ae2af1};
test_output[175:175] = '{32'hc4da1eef};
test_input[1408:1415] = '{32'h42a8d1c0, 32'h42669abf, 32'h41f07079, 32'h4246cd2d, 32'hc2986979, 32'h41bb5231, 32'h413ff107, 32'hc2b618aa};
test_weights[1408:1415] = '{32'h428934bb, 32'h42a80c96, 32'h423921b0, 32'h41b50c59, 32'hc2bc5daa, 32'h427f62bf, 32'hc28365a0, 32'hc1e581e0};
test_bias[176:176] = '{32'h420d10d2};
test_output[176:176] = '{32'h46b90431};
test_input[1416:1423] = '{32'hc21d6c65, 32'h41992bb1, 32'hc24632d0, 32'hc2a2adca, 32'h41daf2aa, 32'hc209ee6e, 32'h412f1a15, 32'h41da784a};
test_weights[1416:1423] = '{32'h41ea015d, 32'h42418502, 32'hc2b23a06, 32'h426b3841, 32'hc19bb1e2, 32'hc2946d37, 32'hc1d9ea79, 32'h4274143b};
test_bias[177:177] = '{32'hc277eee3};
test_output[177:177] = '{32'h452b4366};
test_input[1424:1431] = '{32'hc1f1fd5a, 32'hc2be3034, 32'hc2b1374b, 32'hc19e7c68, 32'h42ad9859, 32'hc1c9fdb1, 32'h421ed874, 32'h423871cc};
test_weights[1424:1431] = '{32'h42422c29, 32'hc26ae111, 32'hc22d0c2e, 32'h4284202a, 32'h429f2b2f, 32'h41b9255f, 32'hc0beb037, 32'hc298dc5a};
test_bias[178:178] = '{32'hc2afcf61};
test_output[178:178] = '{32'h460e6ac0};
test_input[1432:1439] = '{32'h422b6360, 32'hbebf0664, 32'h429784c2, 32'hbf7c9f17, 32'h423f2f45, 32'h42bfe31d, 32'h42c37d41, 32'hc28a0ee9};
test_weights[1432:1439] = '{32'h420a015c, 32'hc22f638d, 32'hc2849378, 32'hc2878c73, 32'h4252ba2a, 32'hc026771b, 32'h4265c9f7, 32'hc2ab31e0};
test_bias[179:179] = '{32'hc09dd83b};
test_output[179:179] = '{32'h46215bda};
test_input[1440:1447] = '{32'h42091c15, 32'h4249203d, 32'h42a17fea, 32'h4227d427, 32'h40e109f1, 32'hc28d5d6f, 32'h42c6c324, 32'h4243c4c0};
test_weights[1440:1447] = '{32'h429ec57f, 32'h40e02712, 32'h41fc80e8, 32'hc282704c, 32'hc2a9e86d, 32'hc0b1e5a5, 32'h41e44285, 32'hc2935a16};
test_bias[180:180] = '{32'hc0f9d379};
test_output[180:180] = '{32'h44ede213};
test_input[1448:1455] = '{32'hc2b8fa39, 32'h4294512d, 32'hc2109184, 32'h42b980cb, 32'hc2bfcddf, 32'hc17468eb, 32'hc2a4c1b1, 32'hc172236a};
test_weights[1448:1455] = '{32'h3ff5d2be, 32'hc1f3bb2e, 32'hc264d888, 32'hc2b4e213, 32'h42bd0c54, 32'h42aac46d, 32'h4296627a, 32'hc22dfee6};
test_bias[181:181] = '{32'hc22451ec};
test_output[181:181] = '{32'hc6c10054};
test_input[1456:1463] = '{32'h418c2944, 32'h40c8c15d, 32'hc2817213, 32'hc25ebfb9, 32'hc263affc, 32'h42b0af70, 32'h420ed866, 32'hc291aa19};
test_weights[1456:1463] = '{32'h429761ac, 32'h41f921c7, 32'h42b5146e, 32'hc262be58, 32'h41b58aaa, 32'hc29af9fc, 32'hc2b99631, 32'hc2b6963f};
test_bias[182:182] = '{32'h419be968};
test_output[182:182] = '{32'hc5ba61f0};
test_input[1464:1471] = '{32'h420ee67f, 32'h416c741d, 32'hc079b9bc, 32'hc28638cd, 32'hc2b57a7f, 32'hc2123cff, 32'hc203e32a, 32'h412921ab};
test_weights[1464:1471] = '{32'h4206b942, 32'hc28fba82, 32'hc2a092e6, 32'h4287af4a, 32'hc26e07b5, 32'h42c4ab3c, 32'hc2c23e3e, 32'h425a2e96};
test_bias[183:183] = '{32'h428cdf1f};
test_output[183:183] = '{32'h44c26dd4};
test_input[1472:1479] = '{32'hc29993ac, 32'h4222d324, 32'h41e32703, 32'hc2079d64, 32'h405bd7c7, 32'h42b34c88, 32'h41b7a7c8, 32'hc2b2352d};
test_weights[1472:1479] = '{32'h40f766b1, 32'h42c46093, 32'h41147673, 32'h424d10b5, 32'hc0d0aa15, 32'hc23ddfac, 32'hc2673606, 32'h42bc4973};
test_bias[184:184] = '{32'hc2afa235};
test_output[184:184] = '{32'hc63de2c7};
test_input[1480:1487] = '{32'hc1cf8ffc, 32'hc29fa2b1, 32'hc26dd231, 32'h422070da, 32'h40ecee1c, 32'hc1701b6e, 32'h42b5a42f, 32'hc1bd59c1};
test_weights[1480:1487] = '{32'hc2a5a3e2, 32'hc1beb6c9, 32'h41c816a3, 32'hc1374b86, 32'hc20e8fe2, 32'h40e96b7e, 32'h419bc610, 32'h40cbd268};
test_bias[185:185] = '{32'h42995562};
test_output[185:185] = '{32'h455620b2};
test_input[1488:1495] = '{32'hc29840e2, 32'hc294bb50, 32'hc22844a8, 32'h41b42dc6, 32'h428dec2e, 32'h419c2d38, 32'h4237712a, 32'h428b59ce};
test_weights[1488:1495] = '{32'hc2a71143, 32'hc28f3395, 32'hc25e8d9b, 32'hc02608de, 32'hc2c40e4f, 32'h42aae5e9, 32'h40ac8128, 32'h41b515f4};
test_bias[186:186] = '{32'h41ffbc33};
test_output[186:186] = '{32'h462498d0};
test_input[1496:1503] = '{32'hc2ae6982, 32'hc2c2ffbb, 32'hc277210b, 32'h419796d4, 32'hc26ca32e, 32'h425a448e, 32'hc2a4755d, 32'h41f6f22c};
test_weights[1496:1503] = '{32'hc2bc6034, 32'hc1b96a63, 32'hc23d269f, 32'h42758218, 32'h429ddddb, 32'hc02b50e7, 32'h4211fbcf, 32'h42bd1617};
test_bias[187:187] = '{32'hc1a41025};
test_output[187:187] = '{32'h46169cbd};
test_input[1504:1511] = '{32'h4219a5db, 32'hc2358c6a, 32'h42c2d2e8, 32'h42bd225d, 32'hc2356439, 32'h419f4876, 32'h420f71ba, 32'h421770f1};
test_weights[1504:1511] = '{32'h41f35b87, 32'h41011016, 32'h415b7640, 32'h422aea98, 32'hc22eaa7f, 32'h419bdcc5, 32'hc2881957, 32'h428176f3};
test_bias[188:188] = '{32'h41d86fa0};
test_output[188:188] = '{32'h46062384};
test_input[1512:1519] = '{32'hc20b5c3a, 32'hc1a0f78b, 32'hc28d40f8, 32'h427b3d74, 32'h42779121, 32'hc22b1e32, 32'hc2375d21, 32'h4200103c};
test_weights[1512:1519] = '{32'hc24741d5, 32'h421a126d, 32'hc2896161, 32'h402a6c50, 32'h42bef879, 32'h4246e827, 32'h41e4dc9c, 32'h41912a3a};
test_bias[189:189] = '{32'hc12c219b};
test_output[189:189] = '{32'h460cf198};
test_input[1520:1527] = '{32'h42c59bbe, 32'hc2adc146, 32'hc28406c1, 32'h428770da, 32'h41318020, 32'hc19c22ca, 32'hc2027616, 32'hc2031168};
test_weights[1520:1527] = '{32'h42a1cc8d, 32'h424eaf97, 32'h423af0ee, 32'hc1a1b532, 32'hc216188c, 32'h41dd9060, 32'h41d169ca, 32'h428357cb};
test_bias[190:190] = '{32'h41095263};
test_output[190:190] = '{32'hc5993de6};
test_input[1528:1535] = '{32'hc1ebcc29, 32'h42a5c224, 32'h3fcada49, 32'h42a26a33, 32'hc2a3476c, 32'hc262eb25, 32'h4256ecbb, 32'h428af31f};
test_weights[1528:1535] = '{32'h42b7e3a4, 32'h4088d402, 32'hc1d7c2b0, 32'h42b65aa8, 32'h427f5d67, 32'hc1ea5b97, 32'h4259709d, 32'hc26c5182};
test_bias[191:191] = '{32'hc0fdb20c};
test_output[191:191] = '{32'h43840f7c};
test_input[1536:1543] = '{32'h421801ba, 32'h42b9edb9, 32'hc25fa90a, 32'h416de2df, 32'h422da84d, 32'hc213262b, 32'hc2b00e76, 32'hc2b260ba};
test_weights[1536:1543] = '{32'hc2b4023f, 32'h424ee205, 32'h4229edf3, 32'h42bee2e7, 32'hc2c050fb, 32'h41816e39, 32'hc2be1007, 32'hc211898a};
test_bias[192:192] = '{32'hc2b6923a};
test_output[192:192] = '{32'h45e06742};
test_input[1544:1551] = '{32'hc2566e31, 32'hc28cea17, 32'hc26badf2, 32'hc136dc5b, 32'hc10d960a, 32'hc2c6be0a, 32'h421743ac, 32'hc2319f74};
test_weights[1544:1551] = '{32'h4213e847, 32'hc2a4c347, 32'hc29dc214, 32'h4292ddc6, 32'h42a204f3, 32'h4225ea46, 32'hc2b25b13, 32'h412ce907};
test_bias[193:193] = '{32'h42a7cd61};
test_output[193:193] = '{32'hc47425bc};
test_input[1552:1559] = '{32'hc08da0c3, 32'hc2715ba3, 32'hc1c20df9, 32'h428e0154, 32'h41e16b9d, 32'hc1e3a978, 32'h4185a032, 32'h4246253b};
test_weights[1552:1559] = '{32'hc15fb2d4, 32'hc1c917d1, 32'hc1309e89, 32'h4280d8d2, 32'hc2292d2a, 32'hc24883eb, 32'hc22a41c0, 32'hc2a0921b};
test_bias[194:194] = '{32'hc0946c38};
test_output[194:194] = '{32'h44f558d3};
test_input[1560:1567] = '{32'h4292627c, 32'hc242ed65, 32'h417b5256, 32'h429ccc84, 32'hc21d5006, 32'hc2a4dcdd, 32'hc220f3f4, 32'h42bb4562};
test_weights[1560:1567] = '{32'h414903d8, 32'h413ed495, 32'h42b352c6, 32'hc2587ff6, 32'h427ca3d0, 32'h42bb936e, 32'h4207ed72, 32'h42bab0ce};
test_bias[195:195] = '{32'hc2a9d508};
test_output[195:195] = '{32'hc5a97c6d};
test_input[1568:1575] = '{32'hc2a3fb49, 32'h3fbf589d, 32'hc273bc33, 32'h40d1e9d8, 32'h41f5595c, 32'hc28eef83, 32'hc26dcc96, 32'h42ba8d86};
test_weights[1568:1575] = '{32'hc2247a48, 32'hc22d1183, 32'hc1e2496a, 32'h41b824ef, 32'h422b1ae5, 32'h424e77b7, 32'hc2098222, 32'hc1c6c6be};
test_bias[196:196] = '{32'hc1e3e173};
test_output[196:196] = '{32'h451c5d0e};
test_input[1576:1583] = '{32'hc26c7616, 32'h405ed403, 32'hc1e4dc1b, 32'h41d0e3c0, 32'h41bcc98f, 32'hc2939d8e, 32'hc2035ef2, 32'hc2a4f60c};
test_weights[1576:1583] = '{32'hc1a28f1f, 32'h4279512c, 32'hc2867095, 32'h42a7ee3b, 32'h4290cbc8, 32'h41f95cd2, 32'hc149aa6c, 32'hc235c999};
test_bias[197:197] = '{32'h421e2682};
test_output[197:197] = '{32'h460eddfc};
test_input[1584:1591] = '{32'h42020769, 32'h4243ccf2, 32'hc2bca639, 32'h41cb9c42, 32'h42817787, 32'hc29acd6a, 32'hc1e2db84, 32'hc21fc653};
test_weights[1584:1591] = '{32'h4261f0d9, 32'h4256444d, 32'hc2b03af6, 32'h428fb960, 32'hc2970dad, 32'h41e0b3d2, 32'hc1d64c82, 32'h4202d630};
test_bias[198:198] = '{32'hc2680ddc};
test_output[198:198] = '{32'h45d8950d};
test_input[1592:1599] = '{32'hc155916a, 32'h403f2518, 32'hc2017d92, 32'h42aaefb5, 32'hc2124aa9, 32'h426f6d10, 32'hc20bb37c, 32'h4232deb9};
test_weights[1592:1599] = '{32'hc10c2a7b, 32'hc2a05747, 32'h410275da, 32'h4209ffff, 32'h4168a1b8, 32'h428c3d7f, 32'hc124fbdc, 32'h40e1c0fe};
test_bias[199:199] = '{32'hc1daa4c3};
test_output[199:199] = '{32'h45d6ded5};
test_input[1600:1607] = '{32'h4231bc99, 32'h42aaf8b6, 32'hc237b1f8, 32'hc2864d2c, 32'hc244e78e, 32'h42c04039, 32'h42169edf, 32'h42916702};
test_weights[1600:1607] = '{32'h42c322b7, 32'hc27677c7, 32'h41db60e1, 32'h42465cd3, 32'hc2c12bd7, 32'h425236dd, 32'hc2bc5b6a, 32'h42998b60};
test_bias[200:200] = '{32'hc1de88af};
test_output[200:200] = '{32'h45c4a154};
test_input[1608:1615] = '{32'h42454691, 32'h40f35eba, 32'h411f4a08, 32'h4298bd9b, 32'hc232edaa, 32'hc1c0c081, 32'h429839bb, 32'h4232025b};
test_weights[1608:1615] = '{32'h42456b9b, 32'hc28b8468, 32'hc2c462cb, 32'hc1aaf881, 32'h4208d2e4, 32'hc213b6bc, 32'h41ce669f, 32'hc2288039};
test_bias[201:201] = '{32'h429c5f17};
test_output[201:201] = '{32'hc49366ea};
test_input[1616:1623] = '{32'hc2467f91, 32'hc2a75aed, 32'h41736e4d, 32'h4131311f, 32'h42271126, 32'h42a5e3ab, 32'h42aa11c1, 32'hc2230f64};
test_weights[1616:1623] = '{32'h42c2edeb, 32'h4277205e, 32'h42801aae, 32'h422cf2ed, 32'hc269c1b5, 32'hc1e1cce2, 32'hc1fb0a50, 32'h42add90a};
test_bias[202:202] = '{32'hc1e99684};
test_output[202:202] = '{32'hc698f005};
test_input[1624:1631] = '{32'hc29f8fe0, 32'h42bf22a7, 32'hc21f7583, 32'h42c6cbc7, 32'h42c69c25, 32'h41d8682d, 32'h4294e598, 32'h425b6918};
test_weights[1624:1631] = '{32'hc29fb771, 32'h427c445c, 32'hc20e16ec, 32'h3ff484c3, 32'hc2b1dcf3, 32'hc233378d, 32'hc1fb5291, 32'h42ab5e99};
test_bias[203:203] = '{32'hc2a1c88a};
test_output[203:203] = '{32'h45c30a2f};
test_input[1632:1639] = '{32'h424bc0cc, 32'hc290553b, 32'h40efae70, 32'h42adb8b5, 32'hc1b98ef1, 32'h42b1fc72, 32'hc1ac1ea0, 32'hc27e6f6e};
test_weights[1632:1639] = '{32'hc114b2fe, 32'h42ace815, 32'h41849453, 32'hc1041243, 32'h41b69bf9, 32'hc223806e, 32'hc24307a8, 32'hc281ec2f};
test_bias[204:204] = '{32'h42a04655};
test_output[204:204] = '{32'hc5c218da};
test_input[1640:1647] = '{32'h42a8ed63, 32'h42a04d88, 32'hc18b0e99, 32'hc273ed2b, 32'hc19fe308, 32'h418b896b, 32'hc1778936, 32'h42012603};
test_weights[1640:1647] = '{32'hc2b0f8f8, 32'h425db0fc, 32'h41da921b, 32'hc02459bd, 32'h42b20be3, 32'h41f47b06, 32'hc2b08f22, 32'hc14ab87f};
test_bias[205:205] = '{32'hc05da191};
test_output[205:205] = '{32'hc563ae64};
test_input[1648:1655] = '{32'hc24b229f, 32'hc17048e4, 32'h42b8b9c9, 32'hc29a575b, 32'h4208e0bb, 32'h422bbece, 32'hc20c9473, 32'hc2084899};
test_weights[1648:1655] = '{32'h41f95f86, 32'h4233991d, 32'hc1f12b8b, 32'hc27e5bdb, 32'h42bdacb7, 32'hc254edef, 32'hc29d651a, 32'h42673153};
test_bias[206:206] = '{32'h42895f22};
test_output[206:206] = '{32'h44d35032};
test_input[1656:1663] = '{32'h402a4843, 32'h426b396b, 32'h42502194, 32'hc2207019, 32'h419f1a58, 32'hc139f43d, 32'h4251e3f3, 32'hc1ae8357};
test_weights[1656:1663] = '{32'h41f36507, 32'h423c1c6f, 32'hc1bed01c, 32'h421fd225, 32'hc2afd8d7, 32'hc26cab59, 32'h42b5b32f, 32'h41e3dd69};
test_bias[207:207] = '{32'h4214d2d4};
test_output[207:207] = '{32'h45434dd2};
test_input[1664:1671] = '{32'h4272f5b1, 32'hc2bdf7df, 32'h41aab312, 32'hc25865cb, 32'h4212c2aa, 32'hc0be5ad7, 32'h42bc99fb, 32'hc0a6feb1};
test_weights[1664:1671] = '{32'hc244a4c1, 32'hc21c3ccf, 32'hc25d55a9, 32'hc2870910, 32'hc11f397f, 32'h42657007, 32'hc2b2811f, 32'h427371fa};
test_bias[208:208] = '{32'h425fbc00};
test_output[208:208] = '{32'hc5c16496};
test_input[1672:1679] = '{32'hc283e0dc, 32'hc10cf163, 32'hc0644b24, 32'hc29cd13d, 32'hc25b163d, 32'h424b61b2, 32'h42a88c27, 32'h418fcb65};
test_weights[1672:1679] = '{32'hc0a2aaaa, 32'hc27fd96c, 32'hc0f1d655, 32'h424f33d0, 32'h421d9837, 32'h4273a097, 32'hc271be7d, 32'h413f01dd};
test_bias[209:209] = '{32'hc180735b};
test_output[209:209] = '{32'hc5dd9e36};
test_input[1680:1687] = '{32'h423f06ec, 32'h419d0851, 32'h4245c740, 32'h412c6959, 32'h4278f6ee, 32'h4291d6d2, 32'hc26c2e12, 32'hc2662e86};
test_weights[1680:1687] = '{32'h422dd590, 32'h41669877, 32'hc25f187b, 32'hc29fefca, 32'h4295d7be, 32'hc25d90e9, 32'h42418d18, 32'hc22debea};
test_bias[210:210] = '{32'h40668f0e};
test_output[210:210] = '{32'hc47718b0};
test_input[1688:1695] = '{32'hc2b7c7f0, 32'h4295fd55, 32'hc180f916, 32'hc2c78809, 32'h428b29ea, 32'hc10fed7f, 32'h42477904, 32'h42b776bc};
test_weights[1688:1695] = '{32'hc2099a4f, 32'hc228de46, 32'hc2afc66e, 32'h42472bdc, 32'h409ffc16, 32'h41fc767d, 32'hc1e8ce94, 32'h40782e47};
test_bias[211:211] = '{32'hc2374a12};
test_output[211:211] = '{32'hc590c801};
test_input[1696:1703] = '{32'h4296afbf, 32'hc2a87134, 32'hc2c5e900, 32'h42207cd1, 32'h416e3878, 32'h428ca715, 32'hc2bd2785, 32'h42bbae67};
test_weights[1696:1703] = '{32'h41f3c41d, 32'h411aeab5, 32'h42c19c8f, 32'hc291576f, 32'hc1b67a14, 32'h42bb15c8, 32'hc2bb74e1, 32'h4264f365};
test_bias[212:212] = '{32'h42858fab};
test_output[212:212] = '{32'h4614daa0};
test_input[1704:1711] = '{32'hc2872768, 32'hc2ada733, 32'h4248a834, 32'hc29f7fd0, 32'hc2b7ff28, 32'hc1e7229e, 32'hc216a338, 32'h400d1bb9};
test_weights[1704:1711] = '{32'hc07b00de, 32'hc164103d, 32'h41e60bf2, 32'hc2a27c1b, 32'hc1e1c603, 32'h415108c1, 32'hc22dc1f2, 32'h428f6554};
test_bias[213:213] = '{32'h4221edf0};
test_output[213:213] = '{32'h46529649};
test_input[1712:1719] = '{32'h41aacee8, 32'hc1a08c2b, 32'hc03f404e, 32'h424e6078, 32'hc0e5edf7, 32'hc11c77bd, 32'h40a34748, 32'hc276f8a1};
test_weights[1712:1719] = '{32'hc2780268, 32'hc1983275, 32'h4229441b, 32'h42ba6c68, 32'hc281be8c, 32'h428edfb6, 32'hc2b77342, 32'hc1a97d02};
test_bias[214:214] = '{32'h4229dfcd};
test_output[214:214] = '{32'h45893629};
test_input[1720:1727] = '{32'hc146bb5e, 32'hc23a97e9, 32'hc16f86ee, 32'h42373840, 32'h42179e7b, 32'h429fe7e6, 32'h429f091c, 32'h42c7c444};
test_weights[1720:1727] = '{32'h4247eaad, 32'hc28202a7, 32'hc1683ce5, 32'hc2a338dc, 32'h427eadfc, 32'hc0c41fe6, 32'hc2b93bab, 32'hc270a5f7};
test_bias[215:215] = '{32'h41b7861a};
test_output[215:215] = '{32'hc643e352};
test_input[1728:1735] = '{32'hc23be356, 32'hc2a84861, 32'h42164344, 32'h4225fc31, 32'hc0755cfb, 32'hc28af74c, 32'hc29e259b, 32'hc2997adf};
test_weights[1728:1735] = '{32'hc08fd7a1, 32'h4229ec80, 32'h41b87ecd, 32'h4228a804, 32'h42bfa9aa, 32'h42bd8d06, 32'hc286fae0, 32'hc13764bb};
test_bias[216:216] = '{32'hc291e7b1};
test_output[216:216] = '{32'hc4c29475};
test_input[1736:1743] = '{32'h41c02de6, 32'h42a2d86c, 32'h403b7f9d, 32'h401ce9dc, 32'hc29022e5, 32'hc198a412, 32'h42b0b87f, 32'hc29a99c3};
test_weights[1736:1743] = '{32'h42663af3, 32'h42b836cf, 32'h42190e44, 32'h423647e2, 32'h4279ca5a, 32'h401f1ddc, 32'h42745f40, 32'hc2bd7b40};
test_bias[217:217] = '{32'hc2c34bf0};
test_output[217:217] = '{32'h46863c72};
test_input[1744:1751] = '{32'h422cd98b, 32'h408e86ff, 32'h42957d29, 32'hc125efdd, 32'h428ddfde, 32'hc294ddb5, 32'hc2bd8568, 32'h41a2ff6d};
test_weights[1744:1751] = '{32'h42b3edd3, 32'h410eaff3, 32'h41b9ea28, 32'h4225134f, 32'h41a72017, 32'h4257830d, 32'h41bc5439, 32'h4291da58};
test_bias[218:218] = '{32'h4187f925};
test_output[218:218] = '{32'h44f780c6};
test_input[1752:1759] = '{32'h42246ee4, 32'h428d5e27, 32'hc24b32a5, 32'hc19bdd30, 32'h420c8ddc, 32'hc24ef3b8, 32'h41976bd6, 32'h427c403b};
test_weights[1752:1759] = '{32'h42891873, 32'hc206b9d1, 32'hc25dd90c, 32'hc28fb420, 32'hc2adc7bb, 32'hc1c512c8, 32'h423101a2, 32'hc255cd2a};
test_bias[219:219] = '{32'h41eb8c68};
test_output[219:219] = '{32'h43ba0cc7};
test_input[1760:1767] = '{32'h418d89f1, 32'hc135abf1, 32'h40d2b7eb, 32'h42aef3d4, 32'hc0bc322f, 32'hc200835e, 32'h41ca41d6, 32'hc27c249f};
test_weights[1760:1767] = '{32'hc245d23d, 32'h427be951, 32'hc0a5ad0a, 32'hc18e0bcb, 32'h41bedd7f, 32'hc23bc38a, 32'h3e3b74b0, 32'h42168ab1};
test_bias[220:220] = '{32'hc1aee1c9};
test_output[220:220] = '{32'hc5833937};
test_input[1768:1775] = '{32'h423f3773, 32'h422690b1, 32'hbb90eaf9, 32'hc29c3b43, 32'h3fdecdb7, 32'h41ba8c1b, 32'hc183b8ac, 32'hc275f1f7};
test_weights[1768:1775] = '{32'hc1ac61c7, 32'hc1441a28, 32'hc04b14a8, 32'hc14368dc, 32'h4278663f, 32'hc199efac, 32'hc27a160e, 32'h42bd26a2};
test_bias[221:221] = '{32'h42777d10};
test_output[221:221] = '{32'hc5b0964c};
test_input[1776:1783] = '{32'hc2a42357, 32'h42bad52a, 32'hc2b0e8f8, 32'h417716ba, 32'h423a3ec8, 32'hc2ad2cd6, 32'h4222b0fb, 32'h425024b6};
test_weights[1776:1783] = '{32'h42b5bea6, 32'hc10eddf3, 32'h415e82e7, 32'h428ab750, 32'h40a0ffba, 32'h422eb9f0, 32'h4270e6d3, 32'h41bbaf68};
test_bias[222:222] = '{32'hc2a9f30f};
test_output[222:222] = '{32'hc6037691};
test_input[1784:1791] = '{32'h4212477a, 32'hc28c8c62, 32'h42144769, 32'h42b0495f, 32'hc1d65fb7, 32'hc13d60c6, 32'hc1a20d42, 32'h42186f4e};
test_weights[1784:1791] = '{32'h409591a0, 32'h424f3d8d, 32'h429b4f66, 32'h40043b08, 32'hc27c889e, 32'hc29d7d2b, 32'hbf96d0cb, 32'h42a6b666};
test_bias[223:223] = '{32'h42b300f9};
test_output[223:223] = '{32'h45ac0461};
test_input[1792:1799] = '{32'h42655a34, 32'hc216e2d0, 32'hc29c88ac, 32'hc146431d, 32'h41d941c0, 32'h4298e498, 32'hc2b7cd34, 32'h42c517c8};
test_weights[1792:1799] = '{32'h417004c3, 32'h40eb8886, 32'h42b3ffec, 32'hc0af83de, 32'hc282f029, 32'h421c8509, 32'hc27f98e1, 32'hbe603236};
test_bias[224:224] = '{32'h408fabc7};
test_output[224:224] = '{32'h4428c971};
test_input[1800:1807] = '{32'hc2a5e456, 32'hc29b0765, 32'h41dd3356, 32'hc12ae3d9, 32'hc2387ad4, 32'hc1f3ef6c, 32'hc13da562, 32'hc299d1c7};
test_weights[1800:1807] = '{32'h4152f86c, 32'h429c0301, 32'hc1b57daa, 32'h4198b8ab, 32'hc1add98d, 32'h4117bf23, 32'hc287604d, 32'h427bd330};
test_bias[225:225] = '{32'hc23f9246};
test_output[225:225] = '{32'hc63147c3};
test_input[1808:1815] = '{32'hc26950c5, 32'h42b057f5, 32'h427b82af, 32'h42b4b6e8, 32'h40375aad, 32'hc2b466f1, 32'h41f59bf5, 32'hc25627ba};
test_weights[1808:1815] = '{32'hc093f95e, 32'h424b692b, 32'h42662f55, 32'h42ae9562, 32'hc19f7b17, 32'h42511ea4, 32'hc13c6785, 32'hc28821dc};
test_bias[226:226] = '{32'h41b3bce2};
test_output[226:226] = '{32'h46671e80};
test_input[1816:1823] = '{32'h428d9fd4, 32'hc225ecba, 32'h428605d5, 32'h420807a4, 32'h41c8e227, 32'h429c4064, 32'hc23ca468, 32'hc2c0c7bd};
test_weights[1816:1823] = '{32'hc2bb9b76, 32'hc291175a, 32'hc295b8e2, 32'h42625a40, 32'hc2c7073e, 32'hc2457212, 32'h411f6b30, 32'h40c32344};
test_bias[227:227] = '{32'hc28439de};
test_output[227:227] = '{32'hc65df14e};
test_input[1824:1831] = '{32'h42587bed, 32'hc21f2548, 32'hc2a67026, 32'hc28c0539, 32'h401eaf67, 32'h42921207, 32'hc253f07a, 32'hc0d93d0c};
test_weights[1824:1831] = '{32'h3c44a3c2, 32'h42c5a00a, 32'hbfdea4cb, 32'h41e2ea67, 32'hc232a83b, 32'h428c203a, 32'hc207c146, 32'h421bff1a};
test_bias[228:228] = '{32'h4163c32f};
test_output[228:228] = '{32'h44438f77};
test_input[1832:1839] = '{32'h42b6ab45, 32'h41f79b36, 32'hc294a84a, 32'hc186b0d2, 32'h428b3bd4, 32'h42915e7d, 32'hc09441c2, 32'hc2b651a5};
test_weights[1832:1839] = '{32'hc25ca861, 32'h428c0c50, 32'h421ca70e, 32'hc247ba14, 32'h41f8b151, 32'hc1af7f88, 32'h42c10b86, 32'h41e4c9c6};
test_bias[229:229] = '{32'hc1d1de53};
test_output[229:229] = '{32'hc5e8e191};
test_input[1840:1847] = '{32'hc2847d1a, 32'hc1bd46d6, 32'hc21dc2b1, 32'h42b83e31, 32'h429a3afe, 32'hc2c458ca, 32'hc1d6bccf, 32'hc09b9094};
test_weights[1840:1847] = '{32'h3f12adfc, 32'h421d1c2b, 32'h42918b3e, 32'hc2c23d8e, 32'hc181e527, 32'h427a765f, 32'hc1eba003, 32'hc288e1ff};
test_bias[230:230] = '{32'hc28cb688};
test_output[230:230] = '{32'hc695752c};
test_input[1848:1855] = '{32'hc24d3a13, 32'hc25055ed, 32'hc25e1856, 32'hc21c54da, 32'hc2b64ebc, 32'hc1e79f25, 32'hc0fc580a, 32'h41778be5};
test_weights[1848:1855] = '{32'hc1dbf7bc, 32'h429982aa, 32'h409f912e, 32'hc1e55463, 32'h427114a5, 32'hc230272a, 32'h42bf7b02, 32'h421a4834};
test_bias[231:231] = '{32'hc156767c};
test_output[231:231] = '{32'hc5bfafaa};
test_input[1856:1863] = '{32'hc20c5c5f, 32'hc052d3af, 32'hc27704d3, 32'hc2971425, 32'h42c6df6a, 32'h4160c76f, 32'hc22ed52f, 32'h4183d8ee};
test_weights[1856:1863] = '{32'h4244f029, 32'h42bf47e4, 32'hc2ba01b0, 32'h425faa28, 32'h41f28c7a, 32'hc1a31f47, 32'h42a7733d, 32'hc1b257ab};
test_bias[232:232] = '{32'hc2511ce1};
test_output[232:232] = '{32'hc4ea40d9};
test_input[1864:1871] = '{32'h40ba76b0, 32'h41ec7ba1, 32'h42915a70, 32'h4046105c, 32'hc221e1a7, 32'h424a8a6e, 32'hc1b260c4, 32'h42592523};
test_weights[1864:1871] = '{32'h3f3bfc8c, 32'h41c60200, 32'h416760da, 32'h422f1863, 32'h4297f298, 32'hc1ba6fb8, 32'h4265f362, 32'hc2b1733b};
test_bias[233:233] = '{32'h4242f2cf};
test_output[233:233] = '{32'hc602f7de};
test_input[1872:1879] = '{32'hc2a01836, 32'h42a70668, 32'h42b31864, 32'h418bc976, 32'hc16d5f9e, 32'h42c26b8c, 32'hc25a10f7, 32'hc127e19a};
test_weights[1872:1879] = '{32'h41d11867, 32'h415a736f, 32'hc1755486, 32'hc1bac842, 32'h3e66ec45, 32'hc0c2d1aa, 32'hc16ee439, 32'h42872826};
test_bias[234:234] = '{32'h4196ba29};
test_output[234:234] = '{32'hc54846ad};
test_input[1880:1887] = '{32'hc1a2a7c3, 32'h42995456, 32'h42c291ae, 32'h41746b3b, 32'hc2a99b78, 32'hc1fb5dfd, 32'h42994cbe, 32'hc24589dd};
test_weights[1880:1887] = '{32'h42c45b21, 32'hc04d5ebf, 32'hc202eac2, 32'hc1885ab7, 32'hc1da43b4, 32'h42b923c9, 32'hc190a00b, 32'hc1871d6f};
test_bias[235:235] = '{32'hc20a1a72};
test_output[235:235] = '{32'hc5d69d24};
test_input[1888:1895] = '{32'h42893d3f, 32'h42ab97bb, 32'h42053a7f, 32'h422ad391, 32'h42a702a6, 32'h421c5b10, 32'hc27d7b0a, 32'h42886a01};
test_weights[1888:1895] = '{32'hbfc6eeec, 32'h4240a1de, 32'h419a90f7, 32'hc17d6a77, 32'h422ac3b9, 32'hc2b7e05c, 32'h42b13c0e, 32'hc228fa2c};
test_bias[236:236] = '{32'hc1fc7174};
test_output[236:236] = '{32'hc58ea984};
test_input[1896:1903] = '{32'hc2a6ad80, 32'hc29309af, 32'h42a3f6db, 32'h42a42148, 32'h4292e00e, 32'h41862801, 32'h410b6a14, 32'hc221e9b4};
test_weights[1896:1903] = '{32'h420c125c, 32'h419abd01, 32'h42358c99, 32'h42a16755, 32'hc1b114de, 32'hc295a6ce, 32'h41ce5e54, 32'h427c99d8};
test_bias[237:237] = '{32'h41154921};
test_output[237:237] = '{32'h44483a1f};
test_input[1904:1911] = '{32'hc2c41bc8, 32'hc13a5d6b, 32'h42a8b62c, 32'h427571cc, 32'hc2a1ec46, 32'hc036da4b, 32'hc266492a, 32'hc272bf99};
test_weights[1904:1911] = '{32'hc0e798ec, 32'hc240fe90, 32'hc1c86355, 32'hc107c87c, 32'hc2a2157a, 32'hc26681b5, 32'h423f667a, 32'hc1a171a9};
test_bias[238:238] = '{32'h4230069f};
test_output[238:238] = '{32'h45725bfb};
test_input[1912:1919] = '{32'hc285dd14, 32'hc188bc4a, 32'hc2c092eb, 32'h428e912a, 32'h425af2aa, 32'hc0e60615, 32'hc29b5e9e, 32'hc229d2f1};
test_weights[1912:1919] = '{32'hc0918d99, 32'h4259d133, 32'hc2384191, 32'h418e1ee2, 32'h41fd6d36, 32'hc1ce562d, 32'hc1f9a979, 32'h41630fb6};
test_bias[239:239] = '{32'hc164ab36};
test_output[239:239] = '{32'h46098984};
test_input[1920:1927] = '{32'hc20203ed, 32'h411b4c52, 32'hc2bfbc64, 32'hc2aa6d84, 32'h429e22c9, 32'h42b88a00, 32'hc2c718df, 32'h42b3723d};
test_weights[1920:1927] = '{32'h422309ee, 32'hc24f966f, 32'hc2ab0f52, 32'hc28e2657, 32'hc18f8ce5, 32'h413d7ac2, 32'hc211d486, 32'h41c8c513};
test_bias[240:240] = '{32'hc1936c34};
test_output[240:240] = '{32'h468c582a};
test_input[1928:1935] = '{32'hc22a0fa2, 32'h429d7ba0, 32'hc0246ad8, 32'h4276b701, 32'hc282abe2, 32'hc2a50791, 32'hc1483b6b, 32'hc1b66e47};
test_weights[1928:1935] = '{32'hc2a35f06, 32'h42c7af1f, 32'hc16bad0b, 32'hc21a2c8b, 32'hc29e7113, 32'hc2990d42, 32'h41c9826a, 32'h3fb7c461};
test_bias[241:241] = '{32'h3f9f8a13};
test_output[241:241] = '{32'h469d55bd};
test_input[1936:1943] = '{32'h3fb7c886, 32'hc0d96d24, 32'hc1de50c3, 32'hc2202a38, 32'hc1c76258, 32'hc1ad1532, 32'hc1c73f57, 32'h42359f96};
test_weights[1936:1943] = '{32'hc2813b83, 32'hc200a91c, 32'hc24364a9, 32'h4235777a, 32'h424f42e7, 32'hc24506f7, 32'h411fa02f, 32'hc2a880f8};
test_bias[242:242] = '{32'h4130b77f};
test_output[242:242] = '{32'hc5906fb9};
test_input[1944:1951] = '{32'hc21ecaa9, 32'hc1e12efc, 32'hc2a0eb2b, 32'hc1ec0944, 32'h42b1d916, 32'hc1f4c9ab, 32'hc2bc1daf, 32'hc26fcc1c};
test_weights[1944:1951] = '{32'h40280ce1, 32'h42936370, 32'h42663490, 32'h42abb853, 32'hc18d2b6c, 32'h4295a7b8, 32'hc2c5bb42, 32'h428acd3c};
test_bias[243:243] = '{32'h42c411eb};
test_output[243:243] = '{32'hc5f8e45d};
test_input[1952:1959] = '{32'h42b198fc, 32'h42b11aa2, 32'hc1d8d973, 32'h4187f7b4, 32'hc2b09ead, 32'h429bb6aa, 32'hc19f54c5, 32'hc2c5ef31};
test_weights[1952:1959] = '{32'hc2a6bcab, 32'hc1a52131, 32'hc1bacd90, 32'hc290853c, 32'hc27928f0, 32'hc1afa9f1, 32'hc29830fa, 32'h420069b9};
test_bias[244:244] = '{32'hc2553731};
test_output[244:244] = '{32'hc5f22dac};
test_input[1960:1967] = '{32'h421868b1, 32'hbed1b19b, 32'hc2c243c7, 32'hc2654d56, 32'h426f05f9, 32'h42ae7627, 32'hc2bd9bef, 32'h42c74b32};
test_weights[1960:1967] = '{32'hc28083f3, 32'h409229dc, 32'hc23cac21, 32'h42b384fb, 32'h41d93072, 32'h41e9e2cf, 32'h429cbf53, 32'h41d96339};
test_bias[245:245] = '{32'h428b32ed};
test_output[245:245] = '{32'hc55a67e7};
test_input[1968:1975] = '{32'hc1a16c7b, 32'h4299f134, 32'hbf0f2806, 32'hc23ceeda, 32'h419845b7, 32'h42be55f8, 32'hc127f9a8, 32'h41bc5aad};
test_weights[1968:1975] = '{32'h42459f43, 32'hc236ea45, 32'hc2c264d4, 32'h41cf6912, 32'hc2a9084f, 32'hc2384bc5, 32'h420dd47b, 32'hc27938a8};
test_bias[246:246] = '{32'hc268c827};
test_output[246:246] = '{32'hc6542708};
test_input[1976:1983] = '{32'h423e749d, 32'h41e69832, 32'hc2705773, 32'h40e03191, 32'hc1122dc0, 32'hc2c4f157, 32'hc27f0cd1, 32'h428420df};
test_weights[1976:1983] = '{32'hc0a93963, 32'h424448fa, 32'h414a82fb, 32'h42c4bc1e, 32'h41f0d781, 32'hc151844f, 32'h4261038d, 32'hc207b5d7};
test_bias[247:247] = '{32'h4275d135};
test_output[247:247] = '{32'hc564d125};
test_input[1984:1991] = '{32'h42477189, 32'hc2c5e5de, 32'h42c33b73, 32'h429843f1, 32'hc17469a6, 32'h421d68e5, 32'hc2abe4dd, 32'hc1b7f813};
test_weights[1984:1991] = '{32'h41c0fd8c, 32'h421445ed, 32'hc2ae75d6, 32'h4249e9bc, 32'hc20856f4, 32'hc25b9a35, 32'h42825835, 32'hc1cf7746};
test_bias[248:248] = '{32'hc2c25f82};
test_output[248:248] = '{32'hc658dc27};
test_input[1992:1999] = '{32'h42acea40, 32'h40b112c6, 32'hc2abd938, 32'hc2914c09, 32'h42a81af2, 32'h4271778d, 32'hc1ae35f1, 32'hc21c1b48};
test_weights[1992:1999] = '{32'hc27f615d, 32'h42a9e3ab, 32'hc2a0ee9d, 32'hc1b870ef, 32'hc1d37bbc, 32'hbfb26721, 32'h42ad4050, 32'hc202f1e8};
test_bias[249:249] = '{32'hc1977c89};
test_output[249:249] = '{32'h44174e24};
test_input[2000:2007] = '{32'h428eb731, 32'hc15cb226, 32'hc04d8b1a, 32'hc2ae80ce, 32'hc2306742, 32'h414692ce, 32'h425b0145, 32'h429a2925};
test_weights[2000:2007] = '{32'h42b720fd, 32'h4294ea2c, 32'h41ff659e, 32'hc1896311, 32'hc1f650bb, 32'h425ef1b6, 32'h4202114f, 32'h429c4752};
test_bias[250:250] = '{32'hc2af4db5};
test_output[250:250] = '{32'h468237e5};
test_input[2008:2015] = '{32'hc20aaa5b, 32'hc20fd16e, 32'hc2966ae9, 32'hc168a219, 32'hc28c2e86, 32'hc1182b53, 32'h416e09d9, 32'h424bcb6d};
test_weights[2008:2015] = '{32'hc0b2f4a7, 32'hc21a07fb, 32'h413094b8, 32'h427323f4, 32'hc2bb5913, 32'hc19f4ebb, 32'hc1eb6571, 32'h42ae5e8f};
test_bias[251:251] = '{32'hc1f29620};
test_output[251:251] = '{32'h46258610};
test_input[2016:2023] = '{32'h42bc5d46, 32'h428eb9d7, 32'hc2b036ac, 32'h42c12b3f, 32'hc250ecc4, 32'hc2a2ae52, 32'hc292d4e1, 32'hc2b1e974};
test_weights[2016:2023] = '{32'hc14cd397, 32'hc2074d66, 32'h42669f79, 32'hc2866698, 32'h42c2b423, 32'hc288316d, 32'h4184e5e2, 32'hc2511a25};
test_bias[252:252] = '{32'hc0ae7a47};
test_output[252:252] = '{32'hc630ba5c};
test_input[2024:2031] = '{32'hc20c3cf9, 32'h42ae7f54, 32'h42066b0b, 32'hc2ad6244, 32'hc1e04017, 32'h41d46ed0, 32'h428b1588, 32'hc2949b5f};
test_weights[2024:2031] = '{32'hc249d5f5, 32'hc0a21bc5, 32'h42b1662d, 32'h4281fdd9, 32'h42942fc6, 32'h402de642, 32'hc0501839, 32'hc1e94c84};
test_bias[253:253] = '{32'hc27cb9fa};
test_output[253:253] = '{32'hc4b5c13a};
test_input[2032:2039] = '{32'hc2a144fe, 32'h42c391ae, 32'hc2944840, 32'h429c5225, 32'h4299bf90, 32'h42a5c6fc, 32'hc06f2c23, 32'h4162a0ab};
test_weights[2032:2039] = '{32'hc02a1062, 32'hc28d5b6a, 32'hc12cbb92, 32'h41670253, 32'hbfbc63d3, 32'h4280ff9e, 32'h42472273, 32'hc2316613};
test_bias[254:254] = '{32'h42955d8a};
test_output[254:254] = '{32'hc3894433};
test_input[2040:2047] = '{32'hc2b0ad7c, 32'hc25c5cd1, 32'hc26786e4, 32'h425c42df, 32'h42669657, 32'h42471f1f, 32'hc1b61db3, 32'hc2167612};
test_weights[2040:2047] = '{32'hc1c5115e, 32'h410971b2, 32'hc293bbf0, 32'h42205f5d, 32'hc29e918c, 32'h41bf7952, 32'h412a184d, 32'h4180efcd};
test_bias[255:255] = '{32'hc18f3f03};
test_output[255:255] = '{32'h45764f39};
test_input[2048:2055] = '{32'hc1fb4e73, 32'h428078da, 32'h415bef5f, 32'h415a9386, 32'hc291c70b, 32'h42470a34, 32'h4235029d, 32'h41f45ef6};
test_weights[2048:2055] = '{32'h4205319f, 32'h4257ecf0, 32'h4200e1e3, 32'h42a85965, 32'hc24c0ca9, 32'h42af9d37, 32'h42c0b13a, 32'hc17c9227};
test_bias[256:256] = '{32'hc0920b2c};
test_output[256:256] = '{32'h46799c03};
test_input[2056:2063] = '{32'h4211ed68, 32'h41a3e466, 32'h41a2a1ad, 32'hc1ac438c, 32'hc125b10a, 32'hc277b90d, 32'h423f6656, 32'hc2951199};
test_weights[2056:2063] = '{32'hc140ca1b, 32'hc2429b2d, 32'hc143d6b5, 32'h42629359, 32'hc2b65b30, 32'hc2a03cfc, 32'hc27e16cd, 32'h42a14b3b};
test_bias[257:257] = '{32'h42469cb2};
test_output[257:257] = '{32'hc5bb7cfc};
test_input[2064:2071] = '{32'hc22cf658, 32'hc265d0a5, 32'hc2c36485, 32'h423f8c99, 32'hc29dffd2, 32'hc1ab0c01, 32'h42af751a, 32'hc0c18a4f};
test_weights[2064:2071] = '{32'hc2ae15fa, 32'hc2b2c526, 32'h42b8f8e0, 32'hc294742e, 32'h424bbe45, 32'hc2c0333c, 32'h42122c37, 32'h42b51561};
test_bias[258:258] = '{32'hc0ce6eea};
test_output[258:258] = '{32'hc53c02ad};
test_input[2072:2079] = '{32'hc29ee5ca, 32'hc1096772, 32'hc241d8f5, 32'h423c8ecb, 32'h4293c4bf, 32'h422fa51f, 32'h41462845, 32'hc2469414};
test_weights[2072:2079] = '{32'hc17d109d, 32'hc2059396, 32'h42bdd699, 32'hc260747e, 32'hc28230e9, 32'h4229253f, 32'h42b4a49e, 32'hc0267391};
test_bias[259:259] = '{32'h428056b8};
test_output[259:259] = '{32'hc5e5743d};
test_input[2080:2087] = '{32'h41ea56a7, 32'hc0ddd458, 32'h4290b912, 32'h42ab5e36, 32'h427cece4, 32'hc24ff242, 32'hc29a0e04, 32'h42930ccf};
test_weights[2080:2087] = '{32'hbfc1426f, 32'hc2c4e50f, 32'hc14c0bc0, 32'hc1a5ed6c, 32'h41ba48bf, 32'hc2843fd5, 32'hc2468750, 32'hc1f5a81f};
test_bias[260:260] = '{32'hc2adc60f};
test_output[260:260] = '{32'h458734fc};
test_input[2088:2095] = '{32'hc1b0074a, 32'h41e3476e, 32'h423bc723, 32'hc2ab5952, 32'hc0b310e1, 32'hc2c2414c, 32'hc13baaca, 32'hc2808986};
test_weights[2088:2095] = '{32'hc244f6f1, 32'hc1299367, 32'hc1f6e531, 32'hc2c5eb5a, 32'hc2a77a4b, 32'hc120ae9b, 32'h41bdaea9, 32'h418359ab};
test_bias[261:261] = '{32'h3e88148f};
test_output[261:261] = '{32'h45f796d1};
test_input[2096:2103] = '{32'hc2b160fa, 32'hc257254c, 32'h417b9635, 32'h42aa24a6, 32'hc21746af, 32'hc144e382, 32'h4217ff67, 32'hc20490f4};
test_weights[2096:2103] = '{32'h41cb927f, 32'hc2139ac6, 32'hc1251d8b, 32'h41d0ed14, 32'h41ae428c, 32'h414c1b11, 32'hc1332b2a, 32'h41e3b4cc};
test_bias[262:262] = '{32'h428f05fc};
test_output[262:262] = '{32'hc3f55b03};
test_input[2104:2111] = '{32'h42ae2070, 32'hc21dd5ae, 32'hc2b3082a, 32'h4294af9d, 32'h421c2f8f, 32'h42579dbe, 32'hbf5da38d, 32'h42830e03};
test_weights[2104:2111] = '{32'h429c55c5, 32'hc2673dee, 32'h4188faed, 32'h429b0435, 32'h41945320, 32'h42758ca4, 32'hc24520d4, 32'h429bc10b};
test_bias[263:263] = '{32'hc244febe};
test_output[263:263] = '{32'h46af5b25};
test_input[2112:2119] = '{32'hc009117b, 32'hc299f089, 32'h42b0af65, 32'hc2a85f57, 32'hc297f16c, 32'hc0e59e72, 32'hc16cad3a, 32'hc1f53dbb};
test_weights[2112:2119] = '{32'h4274c2a2, 32'hc20437b2, 32'h415aa773, 32'h423b2f6a, 32'hc25ff6e3, 32'hc28d4762, 32'h428f604f, 32'hc1c8ca91};
test_bias[264:264] = '{32'h4266178c};
test_output[264:264] = '{32'h45837f68};
test_input[2120:2127] = '{32'h422c59c0, 32'hc1e408ee, 32'h424bfd61, 32'h41a738f8, 32'hc2a01327, 32'hc1cf2950, 32'h40ee68e5, 32'h42880423};
test_weights[2120:2127] = '{32'h42b3e8f9, 32'h42a2ab21, 32'h412a522b, 32'h42c7d483, 32'hc26cbc26, 32'hc21c014c, 32'h42852ef7, 32'h422ca629};
test_bias[265:265] = '{32'h42893b74};
test_output[265:265] = '{32'h4651efba};
test_input[2128:2135] = '{32'h41387cf6, 32'h42b8fb84, 32'h4259ed77, 32'h42958bbf, 32'h42b2da71, 32'h426b43db, 32'hc27a2976, 32'h4287bed9};
test_weights[2128:2135] = '{32'h429d3d92, 32'h423ff3a3, 32'h42a4393b, 32'h41a70a78, 32'h4144a5be, 32'hc2a2a28b, 32'hc199e154, 32'hc13ca768};
test_bias[266:266] = '{32'hc13fda27};
test_output[266:266] = '{32'h45fcb6f7};
test_input[2136:2143] = '{32'hc1b0bc70, 32'h42335c08, 32'h42997cdb, 32'h427059a2, 32'h42291ad5, 32'hc1fa4c4b, 32'h4237cff4, 32'h42768f87};
test_weights[2136:2143] = '{32'h42c32056, 32'h42a3e6bd, 32'h419ed678, 32'hc282a5e2, 32'h402013eb, 32'h41d502b3, 32'h4230137c, 32'h42c49bc4};
test_bias[267:267] = '{32'hc26c318d};
test_output[267:267] = '{32'h45c86e51};
test_input[2144:2151] = '{32'hc279d7f8, 32'h41c9c91c, 32'hc2a2606a, 32'h41c52330, 32'hc297b8fc, 32'hc15b8138, 32'h42bcdf5d, 32'h42b64b11};
test_weights[2144:2151] = '{32'h42718998, 32'hc2407970, 32'hc2261f78, 32'hc210809f, 32'hc10da80d, 32'hc2b88533, 32'hc1ff83d0, 32'hc29a11d3};
test_bias[268:268] = '{32'h42902405};
test_output[268:268] = '{32'hc6249024};
test_input[2152:2159] = '{32'h4220044a, 32'hc2add8ce, 32'hc2b6094a, 32'h42354285, 32'h4244665c, 32'h42339226, 32'h40cbd926, 32'h421cab6d};
test_weights[2152:2159] = '{32'h42c3b0eb, 32'h42aaa774, 32'h416c1236, 32'h41f94f73, 32'hc2b1287c, 32'hc27558cd, 32'h41a0ca7b, 32'hc289141e};
test_bias[269:269] = '{32'hc2870c0d};
test_output[269:269] = '{32'hc64da0e5};
test_input[2160:2167] = '{32'hc2a8742e, 32'h41f1aef1, 32'hc2acf423, 32'h42b7a776, 32'h42130a65, 32'h425f2a80, 32'h42b9ef58, 32'hc2abc565};
test_weights[2160:2167] = '{32'h4288442a, 32'h42bc59a0, 32'h426a3f84, 32'hc184b7ea, 32'hc1f3970e, 32'h42a2dc37, 32'h421e2a8e, 32'hc267e834};
test_bias[270:270] = '{32'h40c4fc45};
test_output[270:270] = '{32'h4522c2e1};
test_input[2168:2175] = '{32'hc2970951, 32'hc1538638, 32'hc23a7358, 32'h4120a8a2, 32'h425b8fe0, 32'h41fb6c98, 32'h429e5b59, 32'hc0e6b00f};
test_weights[2168:2175] = '{32'h42b3262e, 32'h428d1902, 32'h423b334e, 32'h41fd3d87, 32'hc28885dd, 32'hc2c79181, 32'h42283c15, 32'h428e5e1b};
test_bias[271:271] = '{32'h41f40ee3};
test_output[271:271] = '{32'hc65470ff};
test_input[2176:2183] = '{32'hc20706be, 32'h4206612a, 32'h41ef625f, 32'h4293d064, 32'h427d470e, 32'h42452405, 32'h425851da, 32'h42839039};
test_weights[2176:2183] = '{32'hc26d4f6d, 32'hc1c795fd, 32'h42b28c48, 32'h42c112f9, 32'hc0925c1f, 32'hc0d66faf, 32'h411a7aff, 32'hc1e34cf8};
test_bias[272:272] = '{32'hc29b5f64};
test_output[272:272] = '{32'h460b78ee};
test_input[2184:2191] = '{32'h41b757aa, 32'h41d295b1, 32'h415aa442, 32'h3eacada3, 32'hc255fd0a, 32'hc2942191, 32'h4257b2fd, 32'hc27ad441};
test_weights[2184:2191] = '{32'hc2bbed48, 32'h42525cbf, 32'hc18297bc, 32'hc29794e2, 32'h4270297c, 32'h42809fd3, 32'h4273c48c, 32'hc29c618a};
test_bias[273:273] = '{32'hc21548b7};
test_output[273:273] = '{32'hc4523d38};
test_input[2192:2199] = '{32'hbff7a39b, 32'hc29136e6, 32'hc1951d9c, 32'h422bc067, 32'hc2bdb718, 32'h428cb7ef, 32'h42af75ff, 32'h416fc5a8};
test_weights[2192:2199] = '{32'h41bf6e22, 32'h41c1d354, 32'hc23b50f6, 32'h42685304, 32'h424578e0, 32'hc0e7d4b0, 32'h402bff5c, 32'hc1a70cae};
test_bias[274:274] = '{32'h41dcf87b};
test_output[274:274] = '{32'hc5660e1f};
test_input[2200:2207] = '{32'h3f8c20d1, 32'h416c0026, 32'h42b6c2de, 32'h42150d18, 32'h42ae2cc8, 32'h4252323e, 32'h4281909d, 32'h4203d88f};
test_weights[2200:2207] = '{32'h42b503fe, 32'hc23cf5b5, 32'h42868459, 32'hc284521e, 32'hc24697a2, 32'hc1d5114b, 32'h42a8d3b6, 32'h424472f4};
test_bias[275:275] = '{32'h4286ee62};
test_output[275:275] = '{32'h458d14c7};
test_input[2208:2215] = '{32'h42a5349a, 32'h42b215b4, 32'h41f98bbf, 32'hc2ac0b51, 32'hc245248e, 32'h41f1cccd, 32'hc26c613d, 32'h42989c04};
test_weights[2208:2215] = '{32'hc26cc115, 32'h41422c24, 32'hc206385d, 32'hc0d7c162, 32'h4294b807, 32'hc27d3fbb, 32'h40e90c3a, 32'hc29afffa};
test_bias[276:276] = '{32'hc1099336};
test_output[276:276] = '{32'hc67d3928};
test_input[2216:2223] = '{32'h429d5c2a, 32'hc2bb55bd, 32'h41ddb218, 32'h41005504, 32'hc282b81c, 32'hc284b26a, 32'hc2a9e119, 32'h4280bc4d};
test_weights[2216:2223] = '{32'hc2924b8d, 32'hc2b19952, 32'h42005cad, 32'hc14258da, 32'hc214e655, 32'hc2735905, 32'hc1c0ae57, 32'h42672aa3};
test_bias[277:277] = '{32'h3f5e98e4};
test_output[277:277] = '{32'h467398fd};
test_input[2224:2231] = '{32'h4281252a, 32'h42711402, 32'h42baa9bf, 32'hc11f1832, 32'hc239b5df, 32'hc19954ad, 32'hc19aa2a7, 32'h42898431};
test_weights[2224:2231] = '{32'h412fb1c5, 32'h41b7f9a9, 32'h4202ea83, 32'hbea7ff46, 32'h4263f7d6, 32'hc24ff1f1, 32'h425d94e0, 32'hc21bb165};
test_bias[278:278] = '{32'hc1746fa6};
test_output[278:278] = '{32'hc3817a60};
test_input[2232:2239] = '{32'h41c34b9f, 32'hc2967690, 32'hc2bd7e45, 32'h41bc78ca, 32'h41436e69, 32'hc185a038, 32'h426078be, 32'hc2b1c92c};
test_weights[2232:2239] = '{32'h41dbf000, 32'h4294f6e9, 32'h41cbc668, 32'hc29753de, 32'hc297fc4e, 32'hc1fab6f9, 32'hc29ab04d, 32'hc167caba};
test_bias[279:279] = '{32'h3f8078a3};
test_output[279:279] = '{32'hc644a242};
test_input[2240:2247] = '{32'hc238c178, 32'h4264238f, 32'hc23281c8, 32'h4102e1e2, 32'h415ea1bc, 32'hc29c065c, 32'hc2a7f2d4, 32'h421ee82e};
test_weights[2240:2247] = '{32'h41815704, 32'h416d5603, 32'h401eb37d, 32'hc2979bdd, 32'hc2883bcf, 32'h42381c68, 32'h4295a29e, 32'h412d919d};
test_bias[280:280] = '{32'hc21ac67f};
test_output[280:280] = '{32'hc62cd219};
test_input[2248:2255] = '{32'h4213fd17, 32'hc11e3acf, 32'h42b56fda, 32'h3fdf1aee, 32'hc270ac32, 32'hc1b0980b, 32'hc2526cd2, 32'h42a99e4d};
test_weights[2248:2255] = '{32'hc25ba355, 32'h42a2d716, 32'hc128a36e, 32'hc26b8d45, 32'hc2320c40, 32'h4057994b, 32'hc29da835, 32'hc2a40919};
test_bias[281:281] = '{32'h41ba34b5};
test_output[281:281] = '{32'hc57ed5cb};
test_input[2256:2263] = '{32'h4172abc0, 32'hc2b6f7a4, 32'h428bc431, 32'h41c1cec9, 32'h427115e6, 32'h4283127b, 32'hc219b277, 32'h4210621d};
test_weights[2256:2263] = '{32'h42399708, 32'hc09984d3, 32'h42aef648, 32'hc20bf2ff, 32'hc2a26657, 32'h41a354fc, 32'h41e075e9, 32'h41046130};
test_bias[282:282] = '{32'hc18ad865};
test_output[282:282] = '{32'h45007a2b};
test_input[2264:2271] = '{32'h420b7f65, 32'hc26e84dd, 32'hc29eb0a9, 32'hc2c2af1b, 32'h41823b4c, 32'hc20eac34, 32'hc240343f, 32'hc288385d};
test_weights[2264:2271] = '{32'hc1e59f4d, 32'hc21828b4, 32'hc1aa15af, 32'hc1bd4a5f, 32'h428d95e3, 32'hc1c3e741, 32'hc1e1bae7, 32'h42ae5a23};
test_bias[283:283] = '{32'h42771675};
test_output[283:283] = '{32'h452cb5d7};
test_input[2272:2279] = '{32'h427b4af5, 32'hc214758f, 32'hc28a8bae, 32'h4286feba, 32'h4264dede, 32'h41daafcc, 32'h41e419a1, 32'hc2b65fb0};
test_weights[2272:2279] = '{32'hc24314c6, 32'h422752fc, 32'hc2b5b40f, 32'hc2b5f483, 32'h41a473af, 32'h42570d29, 32'h424f4139, 32'hc1b747a5};
test_bias[284:284] = '{32'h42a4f59b};
test_output[284:284] = '{32'h44e4e2e1};
test_input[2280:2287] = '{32'h42b49f30, 32'h42b4c064, 32'h428b0740, 32'hc2a434af, 32'h40b31a20, 32'hc1ecca2a, 32'h428fbaaf, 32'h42556363};
test_weights[2280:2287] = '{32'h421b3204, 32'h420afd89, 32'hbf630377, 32'hc071913d, 32'h420fe305, 32'h412ad0d7, 32'h4285fa8b, 32'hc2a6fa3d};
test_bias[285:285] = '{32'hc2158b6f};
test_output[285:285] = '{32'h45dde64b};
test_input[2288:2295] = '{32'h421dbbba, 32'hc2c15ed8, 32'hc19114a3, 32'hc288a1a9, 32'h41db809f, 32'h41f0aa3b, 32'h4206a5ce, 32'h428b5f15};
test_weights[2288:2295] = '{32'h425a72e9, 32'hc14668d3, 32'hc120cf7b, 32'h4108b4a4, 32'hc138dae5, 32'hc21b7600, 32'hc1f90c2a, 32'h41da5cf6};
test_bias[286:286] = '{32'hc28350bd};
test_output[286:286] = '{32'h450cd64b};
test_input[2296:2303] = '{32'hc0e041e2, 32'hc1fdf578, 32'h40628a3c, 32'h421e8d06, 32'h42c607eb, 32'hc2bc9dc0, 32'h42b36eec, 32'hc16095cb};
test_weights[2296:2303] = '{32'hc2ba95cc, 32'h420c2faf, 32'h4256b194, 32'hc2790464, 32'hc1ac7cc3, 32'hc280f26a, 32'hc2b38bcd, 32'h420e1457};
test_bias[287:287] = '{32'h42009a35};
test_output[287:287] = '{32'hc5e47b81};
test_input[2304:2311] = '{32'h41899518, 32'hc18e45f2, 32'hc22ac5b9, 32'h42a6ae74, 32'hc128634f, 32'hc26ccc50, 32'hc2aae1d5, 32'hc25ceaa8};
test_weights[2304:2311] = '{32'hc1558ce5, 32'hc16b3c54, 32'h428d59eb, 32'hc1e2466f, 32'h41a2fce2, 32'hc2bdfc12, 32'h4297c4ef, 32'h42a9989a};
test_bias[288:288] = '{32'hc29ad14d};
test_output[288:288] = '{32'hc62ea7f3};
test_input[2312:2319] = '{32'hc2a53f20, 32'hc299ac53, 32'hc005f682, 32'hc235658a, 32'h429af7b7, 32'hc2847518, 32'h42b94821, 32'hc2376b47};
test_weights[2312:2319] = '{32'h4131bf54, 32'hc2355a36, 32'h42b6238c, 32'hc1fed8c4, 32'h42a52e5f, 32'hbe264a9b, 32'hc0792d15, 32'hc26f2e0d};
test_bias[289:289] = '{32'hc29df13d};
test_output[289:289] = '{32'h4643d0b0};
test_input[2320:2327] = '{32'h421aeb23, 32'h42a3718c, 32'h42801730, 32'hc1d83414, 32'hc0a09234, 32'hc28978e5, 32'hc22b66df, 32'hc256d936};
test_weights[2320:2327] = '{32'hc29eb046, 32'hc19ecfc5, 32'hc2010181, 32'hc20b08ed, 32'h42b65c14, 32'h4273e401, 32'h42180d55, 32'hc1c781b2};
test_bias[290:290] = '{32'h42be783c};
test_output[290:290] = '{32'hc626a0a0};
test_input[2328:2335] = '{32'h400fef1c, 32'hc2291711, 32'h42616740, 32'hc158c565, 32'h42a316a0, 32'hc2a5b7ba, 32'hc2756257, 32'h42adb283};
test_weights[2328:2335] = '{32'hc261a155, 32'hc2bb2ba8, 32'hc0face24, 32'h427d15bd, 32'hc1fecebf, 32'h412fdc77, 32'h4241866b, 32'hc28ed4e3};
test_bias[291:291] = '{32'hc16b073f};
test_output[291:291] = '{32'hc61ecabe};
test_input[2336:2343] = '{32'hc100d80b, 32'h41d1a16d, 32'hc1910c01, 32'h418b1b18, 32'hc1da1612, 32'h42c4868b, 32'h42a5d15b, 32'h42af38ab};
test_weights[2336:2343] = '{32'h42c30041, 32'hc1d9abea, 32'hc12d3f51, 32'hc20ec615, 32'hc22f1dc7, 32'hc221df8a, 32'hc25322a7, 32'h42971470};
test_bias[292:292] = '{32'hc2c60763};
test_output[292:292] = '{32'hc5202b01};
test_input[2344:2351] = '{32'hc2910c11, 32'hc2c2eda1, 32'hc229dd42, 32'hc2c3ce9a, 32'h422443e7, 32'hc2a70ab7, 32'hc20e548c, 32'h42a5bcfc};
test_weights[2344:2351] = '{32'hc1f047c4, 32'h42a6cf58, 32'hc1eeeb21, 32'h42759b12, 32'hc1a0cea5, 32'hc26e55c5, 32'hc20c9477, 32'hc26b6869};
test_bias[293:293] = '{32'hc23417aa};
test_output[293:293] = '{32'hc61f9988};
test_input[2352:2359] = '{32'hbfc4545a, 32'h3fbbc81c, 32'h425ec732, 32'h41ba2d17, 32'h42281be0, 32'hc2abdb83, 32'h42bd2993, 32'hc287a8c9};
test_weights[2352:2359] = '{32'hc164b75f, 32'hc2b1fe9f, 32'h41fdc36c, 32'hc2260249, 32'hc2b6b613, 32'h426bb6e4, 32'hc233180b, 32'h42665d5f};
test_bias[294:294] = '{32'hc2b60757};
test_output[294:294] = '{32'hc6807615};
test_input[2360:2367] = '{32'h42672d91, 32'h421f9e4d, 32'h4183913b, 32'hc2976aa7, 32'h42912939, 32'hc296de36, 32'h41e6c37e, 32'h411b2ca7};
test_weights[2360:2367] = '{32'h4134178f, 32'hc2793557, 32'h429c1f0f, 32'hc0492139, 32'h429c6b98, 32'hc2bbdaa0, 32'hc2b83233, 32'hc2949d6d};
test_bias[295:295] = '{32'hc238694f};
test_output[295:295] = '{32'h460d021f};
test_input[2368:2375] = '{32'h4239b87f, 32'hc27b30bd, 32'hbea1c9ae, 32'h3c29c7fb, 32'h41d04b0a, 32'h42026836, 32'h4229f621, 32'hc2bcf41e};
test_weights[2368:2375] = '{32'hc202a15a, 32'hc1e55cd8, 32'h4238e453, 32'h41a6d5f5, 32'h40e0fc51, 32'h42a347b7, 32'hc21c5e2c, 32'h41b18313};
test_bias[296:296] = '{32'h420e5c83};
test_output[296:296] = '{32'hc417d817};
test_input[2376:2383] = '{32'hc1c5de1f, 32'h418b7375, 32'hc2234279, 32'hc05f73b5, 32'h4292f20f, 32'h414382f0, 32'h4188c47a, 32'hc24f9738};
test_weights[2376:2383] = '{32'h42a53d89, 32'hc2144f22, 32'h428d8737, 32'h42c5d964, 32'hc1f345d3, 32'hc2bff1c1, 32'h42c48053, 32'h425526da};
test_bias[297:297] = '{32'hc2a59f4a};
test_output[297:297] = '{32'hc6240c19};
test_input[2384:2391] = '{32'h42481ca6, 32'hbcf26540, 32'h426f3076, 32'h41c9e4fc, 32'hc212b652, 32'hc29b1a72, 32'hc292e065, 32'h4263dcdd};
test_weights[2384:2391] = '{32'hc1e68ec9, 32'h420d4c7b, 32'h429bdc27, 32'hc28829bb, 32'h424b1dd4, 32'hc2c7fab1, 32'h42b91299, 32'h427ae9d1};
test_bias[298:298] = '{32'h4160bb1a};
test_output[298:298] = '{32'h4582b4b7};
test_input[2392:2399] = '{32'h42b29b63, 32'hc214fc8a, 32'hc2a78533, 32'hc29db8b9, 32'hc1e70e80, 32'hc2a8fb86, 32'h4265ded8, 32'h411defe1};
test_weights[2392:2399] = '{32'h42b5b963, 32'h41bf3fd3, 32'hc177fbe8, 32'h428af0cc, 32'h421b3039, 32'h424fd68e, 32'hc1c40664, 32'h42bbc5ed};
test_bias[299:299] = '{32'h42344901};
test_output[299:299] = '{32'hc535760c};
test_input[2400:2407] = '{32'hc24d2cbf, 32'h421e0317, 32'h4239efd6, 32'h428cff1a, 32'hc216483e, 32'hc28d7b50, 32'hc0ebf963, 32'h426ead42};
test_weights[2400:2407] = '{32'h424e6d0f, 32'hbfa39632, 32'hc1ec03e7, 32'h42c231ef, 32'hc2780d37, 32'hc20c1c34, 32'hc23ca628, 32'h42a3d495};
test_bias[300:300] = '{32'hc209ba2d};
test_output[300:300] = '{32'h4647c4a4};
test_input[2408:2415] = '{32'hc2986c69, 32'h42426720, 32'h4172853a, 32'h428c6ab3, 32'h42bb3304, 32'h405b4e59, 32'hc29a46be, 32'hc14c76c8};
test_weights[2408:2415] = '{32'h4242596a, 32'h429b024f, 32'h423f9a60, 32'h411d7bcf, 32'h4296ff12, 32'h42a96ac7, 32'h4201d835, 32'hc2c4b488};
test_bias[301:301] = '{32'hc2538479};
test_output[301:301] = '{32'h45eb8e5b};
test_input[2416:2423] = '{32'h42c5e297, 32'hc11e9b9f, 32'h412bea6b, 32'h428756fc, 32'hc138d659, 32'h42235a2d, 32'hc25e484a, 32'h42c48318};
test_weights[2416:2423] = '{32'hc28a9c7d, 32'hc1dadb2a, 32'hc1e8e5db, 32'hc1f5b115, 32'hc2708e8b, 32'hc1430f66, 32'h42715feb, 32'h428f1135};
test_bias[302:302] = '{32'h42ac44d6};
test_output[302:302] = '{32'hc59cd6bb};
test_input[2424:2431] = '{32'hc273bd7b, 32'hc2a12ba2, 32'h42621d03, 32'h426cac0c, 32'h423ce126, 32'hc1bf9df8, 32'h4219bce0, 32'h425fda0e};
test_weights[2424:2431] = '{32'h42879255, 32'hc25366b3, 32'h424910b5, 32'h42a1cc55, 32'hbc51d0e9, 32'h4021ce71, 32'hc2841de5, 32'h424469b1};
test_bias[303:303] = '{32'hbeb885cb};
test_output[303:303] = '{32'h45f7006c};
test_input[2432:2439] = '{32'h42bbe614, 32'h42bfcc78, 32'hc182a0f8, 32'hc244a2bb, 32'h42abb55f, 32'hc293cced, 32'hc16f3bf2, 32'h426bceed};
test_weights[2432:2439] = '{32'hc219e91b, 32'h4287cbf9, 32'h402464fb, 32'h423bd865, 32'hc1d229c8, 32'hc1ada712, 32'hc2825058, 32'hc2740235};
test_bias[304:304] = '{32'h424707df};
test_output[304:304] = '{32'hc5275906};
test_input[2440:2447] = '{32'hc18d9296, 32'hc1b83965, 32'h40d72342, 32'hc289b4f3, 32'h425b033d, 32'h42006261, 32'h41f23e16, 32'hc17a2e12};
test_weights[2440:2447] = '{32'hc2bddd80, 32'hc228065a, 32'h423276f1, 32'h419ce337, 32'h42963ae0, 32'hc1f3501d, 32'h4284a641, 32'hc2555585};
test_bias[305:305] = '{32'h42368370};
test_output[305:305] = '{32'h45ee2be2};
test_input[2448:2455] = '{32'hc12b2e73, 32'hc2bd3e87, 32'h420d2edc, 32'hc0f24b6a, 32'hc2224f18, 32'hc1b48229, 32'hc28d6232, 32'hc2b86e9c};
test_weights[2448:2455] = '{32'h429bd215, 32'hc291f3b1, 32'hc2883557, 32'hc1242607, 32'hc223c8bd, 32'h41cd9112, 32'hc29c496e, 32'hc2c7e9d1};
test_bias[306:306] = '{32'hc28ca28b};
test_output[306:306] = '{32'h4698551e};
test_input[2456:2463] = '{32'hc2aaf645, 32'hc2bbdb41, 32'h4047ab7e, 32'h411e7a18, 32'h426dd5ba, 32'h4211ee0f, 32'hc2a28ba1, 32'h41572844};
test_weights[2456:2463] = '{32'hc2483706, 32'hc2840fee, 32'h40688180, 32'hc27406eb, 32'hc2ad75b0, 32'h42b33a9b, 32'h41c996b1, 32'hc2a68fe1};
test_bias[307:307] = '{32'h41a20f38};
test_output[307:307] = '{32'h4597a676};
test_input[2464:2471] = '{32'hc248ecb6, 32'hc1ed3541, 32'h427af0e4, 32'h4227e0d9, 32'hc2926150, 32'hc27807c6, 32'hc0e74852, 32'hc2a9c2ac};
test_weights[2464:2471] = '{32'hc2a383ef, 32'h41883c77, 32'h40f5e12e, 32'h420dc2b4, 32'hc2617d37, 32'h4280cda4, 32'h42819f70, 32'hc27ad042};
test_bias[308:308] = '{32'hc2a08b04};
test_output[308:308] = '{32'h4623b576};
test_input[2472:2479] = '{32'h4277e7b4, 32'hc1befa55, 32'h4295ad43, 32'h428e7282, 32'hc275da64, 32'hc21a6ca4, 32'hc21d8969, 32'h429196e2};
test_weights[2472:2479] = '{32'h42b2fb6e, 32'h41d48322, 32'hc2b91bec, 32'h420e2c58, 32'h422702f5, 32'hc24be42b, 32'hc2a3ea83, 32'h41d58c95};
test_bias[309:309] = '{32'h423ceeaa};
test_output[309:309] = '{32'h45a08738};
test_input[2480:2487] = '{32'h4185eb0e, 32'hc0f7ee8e, 32'hc2c5047e, 32'hc2a008d0, 32'hc2c24941, 32'hc1f8fee0, 32'h416547e6, 32'h4250be7a};
test_weights[2480:2487] = '{32'hc1ae3d81, 32'h4179e061, 32'hc21a897c, 32'hc29671b0, 32'hc24449b4, 32'h42b72bfa, 32'h4151d0a9, 32'hc275b16d};
test_bias[310:310] = '{32'hc2b20698};
test_output[310:310] = '{32'h45fea982};
test_input[2488:2495] = '{32'h429ee6be, 32'h41be7028, 32'h427ded81, 32'h41e668d4, 32'hc2855e71, 32'h41956f58, 32'h40b1f111, 32'h4232ab7f};
test_weights[2488:2495] = '{32'hc1fb0a3e, 32'hc29b2eef, 32'hc1b22364, 32'h42940272, 32'hc1f9350e, 32'hc2173470, 32'h42b5fcab, 32'h426194ad};
test_bias[311:311] = '{32'h425ac739};
test_output[311:311] = '{32'h444f21ff};
test_input[2496:2503] = '{32'h4194d18d, 32'h404f8ff3, 32'h420e403c, 32'h41d69270, 32'hc207d121, 32'h41ad1d85, 32'hc289d907, 32'h421e78f4};
test_weights[2496:2503] = '{32'hc1be2ee0, 32'h42be89ed, 32'h4233db37, 32'h41dfc95c, 32'h424cb2d3, 32'h41d24790, 32'hc2c2a664, 32'hc2a30cb6};
test_bias[312:312] = '{32'hc25ec595};
test_output[312:312] = '{32'h458baddd};
test_input[2504:2511] = '{32'hc2145318, 32'h423ddf80, 32'h425c9992, 32'hc2a39826, 32'hc0c0e321, 32'h40c0ff8d, 32'hc0b889a7, 32'h42b7ddc8};
test_weights[2504:2511] = '{32'hc25a6cda, 32'hc262e2b8, 32'hc219322c, 32'hbf6c44fd, 32'h420da561, 32'hc214b364, 32'hc252b6d7, 32'hc1bbd870};
test_bias[313:313] = '{32'h42c066da};
test_output[313:313] = '{32'hc5992501};
test_input[2512:2519] = '{32'h411fdd71, 32'hc23acb3f, 32'h41cb1edc, 32'h418bff04, 32'hc2725946, 32'h42813cfa, 32'h41ac7335, 32'h42ade34c};
test_weights[2512:2519] = '{32'hc27f6441, 32'hc22ba903, 32'h421cd325, 32'h41eb544e, 32'h4203cd5a, 32'h42314306, 32'hc2392d52, 32'h42303628};
test_bias[314:314] = '{32'hc01c3fb1};
test_output[314:314] = '{32'h45cd6ac8};
test_input[2520:2527] = '{32'h42b9ec1f, 32'h428af768, 32'h42392f66, 32'h42be760e, 32'h42b26740, 32'hc0aadaa4, 32'hc2ae0963, 32'hc2a8d5a5};
test_weights[2520:2527] = '{32'h42a70b31, 32'h426e6668, 32'h41948c41, 32'h42c15a90, 32'h42504a27, 32'h4285f6a9, 32'hc2a43049, 32'hc2989f19};
test_bias[315:315] = '{32'hc25735d9};
test_output[315:315] = '{32'h471b6ee8};
test_input[2528:2535] = '{32'hc28a6b73, 32'h419fd2a3, 32'h41d37c22, 32'hc1ef55cd, 32'hc18d1242, 32'h421ae4a3, 32'hc2aa0a31, 32'h4287f961};
test_weights[2528:2535] = '{32'h41f1b343, 32'hc20ddbbf, 32'h4220385f, 32'hc1e0fb66, 32'hc236ed52, 32'h4258f035, 32'h424535fc, 32'hc2332e02};
test_bias[316:316] = '{32'h4245bbf4};
test_output[316:316] = '{32'hc5a1e3c4};
test_input[2536:2543] = '{32'h427023f8, 32'h4284f102, 32'h41ed7ceb, 32'hc21eacbf, 32'h4217aec9, 32'hc2469265, 32'h41779be5, 32'hc2a4f5b1};
test_weights[2536:2543] = '{32'h41d719f6, 32'h42c67850, 32'hc272a221, 32'hc2676394, 32'hbf844521, 32'hc2a2c7e7, 32'hc28f56ee, 32'hc297c18c};
test_bias[317:317] = '{32'h425f0828};
test_output[317:317] = '{32'h468bed86};
test_input[2544:2551] = '{32'h4292c5c9, 32'hc2c333f5, 32'hc2b5e54b, 32'hc24af5b0, 32'h42356856, 32'hc29a0270, 32'h41e05d90, 32'h420f5712};
test_weights[2544:2551] = '{32'h4159d2aa, 32'hc1054998, 32'h425e2150, 32'hc23da9f6, 32'h42b165aa, 32'hc235f432, 32'h4294da70, 32'hc2c3416a};
test_bias[318:318] = '{32'h413e08e4};
test_output[318:318] = '{32'h45a56d57};
test_input[2552:2559] = '{32'hc035a85e, 32'hc1a69dc6, 32'hc25718af, 32'hc250806d, 32'hc274ae34, 32'hc1e2f954, 32'hc20b5721, 32'h427fdf74};
test_weights[2552:2559] = '{32'hc29ac785, 32'h4096ca93, 32'h429b2b58, 32'h42b2358f, 32'hc033b7b5, 32'h427d46a1, 32'h4243574b, 32'hc205a2ff};
test_bias[319:319] = '{32'h426d692c};
test_output[319:319] = '{32'hc65c4b29};
test_input[2560:2567] = '{32'hc27e95fb, 32'h421cf400, 32'hc29e7e99, 32'h427a6cb6, 32'h425d0d29, 32'hc151a969, 32'h41e30cc1, 32'hc2b30ed8};
test_weights[2560:2567] = '{32'hc2bf44f7, 32'hc24c6003, 32'hc2b8a76f, 32'h4090d06b, 32'hc2beae72, 32'h429c227d, 32'h418c5e5a, 32'hc2be9390};
test_bias[320:320] = '{32'hc25661ca};
test_output[320:320] = '{32'h4660767b};
test_input[2568:2575] = '{32'h424e77d8, 32'h41668e15, 32'h4292b295, 32'h421d40a1, 32'hc18388b8, 32'hc17fed9c, 32'hc1982e0a, 32'hc1228ddc};
test_weights[2568:2575] = '{32'h42c5a031, 32'hc2b7e09c, 32'hc28e8bec, 32'h416cc750, 32'hc2a49bf1, 32'h42a9cb48, 32'hc1cebf91, 32'h42c3a7d4};
test_bias[321:321] = '{32'hc20b6098};
test_output[321:321] = '{32'hc4b088e9};
test_input[2576:2583] = '{32'h426c8b14, 32'hc220110b, 32'hc2b976fa, 32'hc1953c75, 32'hc2b509b1, 32'hc290481d, 32'hc2068145, 32'h410532ff};
test_weights[2576:2583] = '{32'hc1af6183, 32'hc2049ae1, 32'h426d48c4, 32'h42954055, 32'h41ca62a1, 32'h41379b9d, 32'hc280dcf4, 32'h42710dda};
test_bias[322:322] = '{32'hc2ae3219};
test_output[322:322] = '{32'hc5e73c3b};
test_input[2584:2591] = '{32'hc1adbcb5, 32'hc2bdbd40, 32'hc267b563, 32'hc26ee58c, 32'hc1e899f0, 32'h421946c2, 32'hc24aaed3, 32'hc29f8642};
test_weights[2584:2591] = '{32'hc1842e41, 32'h4286b5bb, 32'h42ad1881, 32'hc28ee0e9, 32'hc245a8fa, 32'hc2bb2e96, 32'hc2c18b38, 32'hc27d50eb};
test_bias[323:323] = '{32'h4177f7d1};
test_output[323:323] = '{32'h44825848};
test_input[2592:2599] = '{32'h416cc872, 32'h4282ecc9, 32'hc266874d, 32'hc2c13118, 32'h424a053b, 32'hc2c037fe, 32'h41e81654, 32'hc2bb19ae};
test_weights[2592:2599] = '{32'h4267348b, 32'h413e6f28, 32'hc213383a, 32'hc2a52cf0, 32'hc27912d5, 32'hc1a38755, 32'hc0a61946, 32'hc2900cc2};
test_bias[324:324] = '{32'h4287d6e5};
test_output[324:324] = '{32'h4686709f};
test_input[2600:2607] = '{32'h41c8258e, 32'hc1b1d7be, 32'hc2c4f50f, 32'hc28b3879, 32'hc07f281a, 32'h42982afe, 32'h42c0595b, 32'h42b3550a};
test_weights[2600:2607] = '{32'h42652372, 32'hc173c573, 32'hc2847166, 32'hc07442c0, 32'h414b4ebc, 32'h42a8ea4a, 32'h423500c0, 32'hc29a755a};
test_bias[325:325] = '{32'hc1da46cc};
test_output[325:325] = '{32'h4640b7f2};
test_input[2608:2615] = '{32'hc29782ed, 32'h41049108, 32'hc1f346ae, 32'hc257470f, 32'hc1164376, 32'hc16f2890, 32'h4264abc6, 32'hc1a18379};
test_weights[2608:2615] = '{32'h422c6e52, 32'h4231781b, 32'h41e93416, 32'h4266613c, 32'h4221b14c, 32'h42603df4, 32'h428fdada, 32'hc15a4649};
test_bias[326:326] = '{32'hc2a797c2};
test_output[326:326] = '{32'hc56d6441};
test_input[2616:2623] = '{32'hc27a2972, 32'h428019f1, 32'hc2c7fd6c, 32'h42a41acc, 32'h423eb46a, 32'h42c3f6f5, 32'h41916a3b, 32'h427a3923};
test_weights[2616:2623] = '{32'h42b8cbd7, 32'hc25e3385, 32'hc2b3f7a0, 32'hc1f2f408, 32'hc2b99cd0, 32'h423c763b, 32'h4291ae9a, 32'hc2b888e6};
test_bias[327:327] = '{32'h42933958};
test_output[327:327] = '{32'hc5db27fc};
test_input[2624:2631] = '{32'h42497c97, 32'h426fa879, 32'h40f15c72, 32'h4234ea58, 32'hc27ad9ba, 32'hc22c959e, 32'h4205c033, 32'hc2961036};
test_weights[2624:2631] = '{32'hc25a85d6, 32'h4258fce0, 32'h42c28971, 32'hc2b70a99, 32'hc2a6f5a4, 32'hc27d8539, 32'hc213067a, 32'hc11e04b5};
test_bias[328:328] = '{32'hc2618b07};
test_output[328:328] = '{32'h458d305f};
test_input[2632:2639] = '{32'h41214047, 32'hc087fc93, 32'h4293944d, 32'hc20525bb, 32'hc2b85f30, 32'h42b7bca3, 32'h424154dd, 32'hc1729bbb};
test_weights[2632:2639] = '{32'hc2784c53, 32'h4271f027, 32'h42a4ab10, 32'hc277f4dc, 32'hc1c231b4, 32'h40361df9, 32'h42c6c817, 32'h4216eb15};
test_bias[329:329] = '{32'h40623e62};
test_output[329:329] = '{32'h465a9a92};
test_input[2640:2647] = '{32'h427c2d16, 32'hc165c76a, 32'h428a6a66, 32'hc2251e8d, 32'hc0aa00ea, 32'hc1e96d44, 32'hc2c160c0, 32'hc2aefe65};
test_weights[2640:2647] = '{32'hc25ea7be, 32'hc180c1e9, 32'h4257bfa5, 32'hc2a42c9f, 32'hc22d7f6f, 32'hc2b526d3, 32'hc234af6e, 32'h428152c4};
test_bias[330:330] = '{32'h412d78e2};
test_output[330:330] = '{32'h45a9ea4d};
test_input[2648:2655] = '{32'hc2b4290a, 32'h42bd6f29, 32'h42c22005, 32'hc282b8ef, 32'h42c0c322, 32'hc27b6b06, 32'hc28b514c, 32'hc24f5543};
test_weights[2648:2655] = '{32'h408e20b8, 32'h42a3afe0, 32'hc0be2cec, 32'hc264a544, 32'hc12ca0f2, 32'h42bc3dfc, 32'h42b8a760, 32'h41f057e9};
test_bias[331:331] = '{32'hc0f7d07c};
test_output[331:331] = '{32'hc58ac7d5};
test_input[2656:2663] = '{32'h4232f5a2, 32'h4190cb78, 32'h41c7c2e9, 32'h42627a08, 32'h4116329c, 32'h42aa5c72, 32'hc1f38acb, 32'h42c6ba4c};
test_weights[2656:2663] = '{32'h427135ba, 32'h42616109, 32'hc237a07c, 32'hc2c5f8e9, 32'h41822ead, 32'hc0c938a4, 32'h420af027, 32'hc2716acf};
test_bias[332:332] = '{32'h42a1b6df};
test_output[332:332] = '{32'hc6225633};
test_input[2664:2671] = '{32'h42a99fd5, 32'h42890d2e, 32'h40c2343f, 32'h4179cc67, 32'h42bb2585, 32'h41e68c88, 32'h41d511b2, 32'h41b07eba};
test_weights[2664:2671] = '{32'hc199bbae, 32'h424c06f9, 32'h42365a44, 32'h4272b13c, 32'hc25b82a0, 32'h4287aad5, 32'hc29ab1f1, 32'hc1678814};
test_bias[333:333] = '{32'hc271024b};
test_output[333:333] = '{32'hc51e25b1};
test_input[2672:2679] = '{32'hc20cd949, 32'h421525cd, 32'hc1768db3, 32'h4208b849, 32'h42c6d04e, 32'h429b7ec8, 32'hc28bb708, 32'hc26e5c03};
test_weights[2672:2679] = '{32'h42c6bc55, 32'hc278e257, 32'h422e5bd5, 32'hc2b53ff6, 32'hc2a0b7d6, 32'h410b7103, 32'hc2379d38, 32'h428cc708};
test_bias[334:334] = '{32'h42adbbb8};
test_output[334:334] = '{32'hc68b0f95};
test_input[2680:2687] = '{32'h41c22d62, 32'hc202aac4, 32'hc0a45536, 32'h41e90826, 32'hc1e7ddc3, 32'h429c597d, 32'hc2c63361, 32'h42aa5d99};
test_weights[2680:2687] = '{32'hc18f100a, 32'hc2c5fce9, 32'hc1d20ff1, 32'hc22cef06, 32'h41c8be37, 32'hc21ee523, 32'h425789e8, 32'hc1de4e9d};
test_bias[335:335] = '{32'hc2271836};
test_output[335:335] = '{32'hc61ac915};
test_input[2688:2695] = '{32'hc27b0957, 32'h40900ddf, 32'h41d5c68c, 32'hc22720a5, 32'h406d8a6c, 32'hc2920a4a, 32'hc2a1078d, 32'h425fd1a3};
test_weights[2688:2695] = '{32'hc1b69ed3, 32'h4228b7a1, 32'h42b1f3cc, 32'hc2c74ca0, 32'hc251233b, 32'h42b26333, 32'h412cc32e, 32'hc271f605};
test_bias[336:336] = '{32'hc2a90c8f};
test_output[336:336] = '{32'hc5341ec0};
test_input[2696:2703] = '{32'h428fcbe1, 32'hbd684949, 32'h3f622333, 32'hc2a8a627, 32'h4211fb32, 32'hc22d7834, 32'h42b1fb2c, 32'hc1dafaa8};
test_weights[2696:2703] = '{32'hc2a242b9, 32'h41ef4048, 32'h3e043681, 32'h41f92cfd, 32'h428bbd12, 32'hc2bb6b24, 32'h425e4d42, 32'h41371a86};
test_bias[337:337] = '{32'h41300e07};
test_output[337:337] = '{32'h452ec1cd};
test_input[2704:2711] = '{32'hc25f19a0, 32'h411199d6, 32'h42a39861, 32'h42ad19a8, 32'hc1a74eba, 32'h413fbf26, 32'hc29506f6, 32'hc1e7e9e2};
test_weights[2704:2711] = '{32'hc21c4c83, 32'hc25ebae9, 32'h4248e87e, 32'h41af2cfc, 32'hc14e1dfd, 32'h401cbc8f, 32'h421f786f, 32'h41f472d2};
test_bias[338:338] = '{32'hc0a587f1};
test_output[338:338] = '{32'h45808b73};
test_input[2712:2719] = '{32'h416d569d, 32'hc1ab4d45, 32'hc2c48e54, 32'hc1a28d63, 32'h4229deec, 32'h429dde90, 32'hc2a87f46, 32'h4228936b};
test_weights[2712:2719] = '{32'hc1f7acb3, 32'hc22750f1, 32'h41a8bb52, 32'h42a1e8ea, 32'h3fd17d0e, 32'h429ddaa6, 32'hc281ec90, 32'h41146d81};
test_bias[339:339] = '{32'h4230687c};
test_output[339:339] = '{32'h460b7927};
test_input[2720:2727] = '{32'hc20de0d9, 32'h41a509d6, 32'hc1b82bd8, 32'h4282dbfa, 32'h42af5d03, 32'hc215dd47, 32'h4298177a, 32'hc20d8c38};
test_weights[2720:2727] = '{32'hc2829927, 32'h42c791a9, 32'hc2a09ddd, 32'h42780b5e, 32'h42af8b58, 32'h42bd3992, 32'h4238f90f, 32'h4215da06};
test_bias[340:340] = '{32'hc21e737b};
test_output[340:340] = '{32'h46818ec6};
test_input[2728:2735] = '{32'h41691c69, 32'hc2ac3225, 32'hc245d099, 32'h3f8c51c2, 32'h426685aa, 32'hc2a50ee5, 32'hc0547b34, 32'hc290c454};
test_weights[2728:2735] = '{32'hc1d5aa7e, 32'h429a2f0c, 32'hc224abcb, 32'hc2c7e8f5, 32'hc1d30177, 32'hc29f99a5, 32'h41f50959, 32'h428dfbc2};
test_bias[341:341] = '{32'hc175c302};
test_output[341:341] = '{32'hc5a5512f};
test_input[2736:2743] = '{32'h42771178, 32'hc29acd2f, 32'hc2168240, 32'hc2a2fa5a, 32'hc2a87e08, 32'hc2c1fb39, 32'hc23b64b9, 32'h40e13d11};
test_weights[2736:2743] = '{32'h42c4d18c, 32'h4289e917, 32'h42800409, 32'hc27350fa, 32'h417a7f7e, 32'hc27ca142, 32'h41bae328, 32'hc1a824b1};
test_bias[342:342] = '{32'hc1df0530};
test_output[342:342] = '{32'h45d551a3};
test_input[2744:2751] = '{32'h42513704, 32'h42bacb44, 32'hc2c42513, 32'h429727f3, 32'hc1bd2356, 32'hc28bb820, 32'hc186d9a6, 32'h418702d2};
test_weights[2744:2751] = '{32'h416101ec, 32'h40fa331d, 32'hc2aee6b1, 32'h4104e9f5, 32'hc1b571e0, 32'hc11d805c, 32'h42ab5046, 32'h42c1f3f2};
test_bias[343:343] = '{32'h421c258d};
test_output[343:343] = '{32'h463d7745};
test_input[2752:2759] = '{32'hc2b31c9e, 32'h42006ad5, 32'h4273e560, 32'h415c225f, 32'h42b45d94, 32'hc0a2c243, 32'h412ef2c4, 32'hc144f67e};
test_weights[2752:2759] = '{32'hc1baff84, 32'hc15cca92, 32'hc21518df, 32'h42a16c8e, 32'h42123666, 32'hc29b744e, 32'hc26c5425, 32'h427422fe};
test_bias[344:344] = '{32'h424527b3};
test_output[344:344] = '{32'h4530fc1b};
test_input[2760:2767] = '{32'h425b2a9c, 32'hc2b4005c, 32'hc22bacd5, 32'hc1a88308, 32'h40c79675, 32'h41f03135, 32'h42850ccb, 32'hc107d107};
test_weights[2760:2767] = '{32'h428c342d, 32'hc22580bf, 32'h41f9bde5, 32'hc2c73e7d, 32'hc240e341, 32'h40e76e9d, 32'h4291ca51, 32'h42087922};
test_bias[345:345] = '{32'hc181576f};
test_output[345:345] = '{32'h4647bd93};
test_input[2768:2775] = '{32'hc2aa4da2, 32'hc2bc1f29, 32'hc2765c2b, 32'h40a77a70, 32'h424f675e, 32'hc241bbe0, 32'hc2859987, 32'hc1e78c92};
test_weights[2768:2775] = '{32'hc21ff258, 32'h411ed50c, 32'hc164182d, 32'hc254e6ba, 32'h42c22294, 32'h3e4c0af9, 32'hc24ba0eb, 32'h42a104f0};
test_bias[346:346] = '{32'h42046204};
test_output[346:346] = '{32'h460fb5ea};
test_input[2776:2783] = '{32'h42c6103e, 32'hbe853c79, 32'hc2145071, 32'h4110eae8, 32'hc29f66ae, 32'h424f923a, 32'h42365f1b, 32'h418ed7c0};
test_weights[2776:2783] = '{32'hc28d43ef, 32'hc28093f0, 32'hc2a755dc, 32'hc2aa019c, 32'hc2a4751e, 32'hc18933fb, 32'hc2443bed, 32'hc21e5d37};
test_bias[347:347] = '{32'h410187c2};
test_output[347:347] = '{32'hc4efb3a3};
test_input[2784:2791] = '{32'h42be1d7e, 32'h3f6bb9e9, 32'hc1575281, 32'h425bd88a, 32'hc274341a, 32'h423bd6bb, 32'h42481544, 32'hc29b2135};
test_weights[2784:2791] = '{32'h422d7f76, 32'h4273a198, 32'h428656e3, 32'h42b333a6, 32'h42433fb2, 32'hc22f3ef0, 32'h40885870, 32'h42aefd77};
test_bias[348:348] = '{32'h4223e39e};
test_output[348:348] = '{32'hc552a08c};
test_input[2792:2799] = '{32'h42923289, 32'hc24397b1, 32'h41c99a43, 32'h416142bc, 32'h41221387, 32'h42812e86, 32'hc2b696b5, 32'hc14dd2e3};
test_weights[2792:2799] = '{32'hc29bf8e9, 32'hc1938887, 32'hc1acfcaa, 32'h41b34d33, 32'h428275bc, 32'h4297200a, 32'h41e063d3, 32'hc21acb49};
test_bias[349:349] = '{32'hc211f6fc};
test_output[349:349] = '{32'hc4c647d8};
test_input[2800:2807] = '{32'hc23dd734, 32'h4258a0de, 32'hc28f10d2, 32'hc2a0dfb0, 32'hc20d9757, 32'hc210319f, 32'h428b35d9, 32'hc2710904};
test_weights[2800:2807] = '{32'hc2496f21, 32'hc2451aa8, 32'h42ba458e, 32'h42a43927, 32'h42aa6b0d, 32'hbf2de605, 32'h42b9d8fc, 32'hc28904a4};
test_bias[350:350] = '{32'hc277972a};
test_output[350:350] = '{32'hc5bb9895};
test_input[2808:2815] = '{32'hc2a3ae61, 32'h419aa687, 32'hc2049f6a, 32'hc27e0c14, 32'h4276c797, 32'hc26d296b, 32'h41f095b1, 32'h426a5e5f};
test_weights[2808:2815] = '{32'h4294ee19, 32'hc2baf5ac, 32'hc2192d45, 32'h42b2e0c1, 32'hc2962cb0, 32'hc2a8b248, 32'h40eb6d3c, 32'hc1c202e1};
test_bias[351:351] = '{32'hc2c5acaf};
test_output[351:351] = '{32'hc64ee865};
test_input[2816:2823] = '{32'hc1525419, 32'hc235b6ce, 32'h423f6a40, 32'h429c8010, 32'h3fdbb87a, 32'hc28a027a, 32'hc166bc54, 32'hc2a9d14c};
test_weights[2816:2823] = '{32'hc0a1a29b, 32'h41ca12ca, 32'h41f0ee19, 32'hc2bd7caf, 32'hc2929651, 32'h428f53b4, 32'hc00b6e4f, 32'hc2ab810a};
test_bias[352:352] = '{32'h41822b69};
test_output[352:352] = '{32'hc595de09};
test_input[2824:2831] = '{32'h42695ba5, 32'hbfdba530, 32'h42b242d2, 32'h4284d55c, 32'hc26dae1d, 32'hc284e3d6, 32'h42aa8f6f, 32'h42c3eba6};
test_weights[2824:2831] = '{32'hc2450364, 32'hc2755404, 32'hc0c1dff0, 32'hc231b32d, 32'hc2566cd8, 32'hc23275b9, 32'h428721ac, 32'hc2b79638};
test_bias[353:353] = '{32'hc21e63d2};
test_output[353:353] = '{32'hc5532b08};
test_input[2832:2839] = '{32'hc2c05c2d, 32'hc287224e, 32'h3fdb3b69, 32'hc23f72cb, 32'h416841a6, 32'h4267d814, 32'hc23d928b, 32'hc295c995};
test_weights[2832:2839] = '{32'hc2150ff2, 32'hc2a18bc4, 32'hc2ad191c, 32'h429fb4a8, 32'h41d1fe11, 32'hc2ab2af0, 32'hc2442b49, 32'hc26a6c87};
test_bias[354:354] = '{32'h41493cc6};
test_output[354:354] = '{32'h45e19195};
test_input[2840:2847] = '{32'hc183df7a, 32'h429888de, 32'hc2989e49, 32'h42a15b01, 32'hc2949559, 32'h41da47ba, 32'hc296468e, 32'h4287a882};
test_weights[2840:2847] = '{32'h429ea014, 32'hc2c2f07b, 32'h420277f4, 32'hc205702d, 32'h42874c1b, 32'hc1b39b9a, 32'h410688ca, 32'hc2b4bfc3};
test_bias[355:355] = '{32'hc2401bde};
test_output[355:355] = '{32'hc6ce0351};
test_input[2848:2855] = '{32'hc22e51b1, 32'hc225c3e4, 32'hc292f02a, 32'hc2978416, 32'hc2b50ede, 32'hc24fcd27, 32'hc0c34399, 32'hc1967bbe};
test_weights[2848:2855] = '{32'hc21814e5, 32'hc1720a2d, 32'h42884255, 32'hc24143ca, 32'h42359649, 32'h42a323ae, 32'hc225b6dd, 32'h4234e774};
test_bias[356:356] = '{32'h41f89f95};
test_output[356:356] = '{32'hc5f93b2e};
test_input[2856:2863] = '{32'hc26afceb, 32'h42597853, 32'h427b5464, 32'h4223110a, 32'h428d701c, 32'hc267ad0a, 32'h428a61f2, 32'h4286b11e};
test_weights[2856:2863] = '{32'h428077d0, 32'h42c60c50, 32'hc2b8587a, 32'h3eab9845, 32'h423788c3, 32'h4207bb64, 32'h42c5951d, 32'hc2817a7f};
test_bias[357:357] = '{32'h426ed49d};
test_output[357:357] = '{32'hc3b07230};
test_input[2864:2871] = '{32'h42b81a91, 32'h4224e662, 32'h429ac5d6, 32'h425150d5, 32'h4220ea30, 32'h427c814b, 32'hc2b096bd, 32'hc24f9c5a};
test_weights[2864:2871] = '{32'hc2536f90, 32'h4210f2fe, 32'h41421e58, 32'h42bec759, 32'hc1b5a9de, 32'h42371698, 32'h410836e2, 32'hc2023f08};
test_bias[358:358] = '{32'h41fb30c4};
test_output[358:358] = '{32'h45ac0236};
test_input[2872:2879] = '{32'h41d29040, 32'h4253cb85, 32'hc2359533, 32'hc1ddb6a3, 32'hc2a27369, 32'hbf72dd5c, 32'h42b37cfc, 32'h41891e09};
test_weights[2872:2879] = '{32'hc1a5a81f, 32'hc191331d, 32'h42864f97, 32'hc1d68a81, 32'hc20c37e3, 32'h425abd2e, 32'hc2adb390, 32'hc2bfe784};
test_bias[359:359] = '{32'h4101aa06};
test_output[359:359] = '{32'hc6233b08};
test_input[2880:2887] = '{32'hc1dce348, 32'h42b54352, 32'hc2baa0de, 32'h41c7a534, 32'h4276a2dc, 32'h42c7a21d, 32'hc22af694, 32'hc2a29860};
test_weights[2880:2887] = '{32'h427024d0, 32'hc2105416, 32'hc2c4404c, 32'hc29a1b7e, 32'hc10c4e95, 32'h427027c5, 32'hc289b2ab, 32'h418b5a0f};
test_bias[360:360] = '{32'h4251dd1d};
test_output[360:360] = '{32'h4611e3be};
test_input[2888:2895] = '{32'hc03e2818, 32'h41df2af6, 32'hc1a2abd1, 32'hbfad6a43, 32'h42bcda9e, 32'h42097cda, 32'hc1cbf165, 32'h42c0401b};
test_weights[2888:2895] = '{32'hc1aebd20, 32'h42b2be6f, 32'hc1151d14, 32'hc210299e, 32'h42725620, 32'h4182a474, 32'h42b6866f, 32'h41f5d657};
test_bias[361:361] = '{32'hc25f0e39};
test_output[361:361] = '{32'h4616c80c};
test_input[2896:2903] = '{32'hc258105c, 32'hc26304f1, 32'hc199e5d7, 32'hc26773f2, 32'hc1dce077, 32'hc0cce93d, 32'h417a6dfb, 32'h41a53397};
test_weights[2896:2903] = '{32'hc21305b2, 32'h425e4dee, 32'h4271a1e6, 32'h42b3bcc0, 32'hc19e9fa6, 32'h42796961, 32'hc1a18fe4, 32'hc11dc72f};
test_bias[362:362] = '{32'h41df73a0};
test_output[362:362] = '{32'hc5f61507};
test_input[2904:2911] = '{32'h428e1a24, 32'h4225cd5d, 32'hc2ab053a, 32'hc223e2cb, 32'hc28911c5, 32'hc2a6ecdb, 32'h42a924e8, 32'hc0b42f4f};
test_weights[2904:2911] = '{32'h429bcfbd, 32'h4271aa0c, 32'h429c9d6b, 32'hbf311620, 32'hc21b7bc2, 32'h41b3c23b, 32'h42581df9, 32'hc2b7bafd};
test_bias[363:363] = '{32'hc05b3a96};
test_output[363:363] = '{32'h45e25d28};
test_input[2912:2919] = '{32'h404411ab, 32'h42b42810, 32'h423aa264, 32'hc1eb87b0, 32'hc211e08e, 32'h429ee2ee, 32'hc2839f1b, 32'h4219cb76};
test_weights[2912:2919] = '{32'h42a74d14, 32'hc20441c0, 32'hc1d72242, 32'hc2940e95, 32'hc2b6672f, 32'hc26801fa, 32'hc226361f, 32'hc21c328b};
test_bias[364:364] = '{32'hc2a2d0e2};
test_output[364:364] = '{32'hc4f0ea42};
test_input[2920:2927] = '{32'h420ef4bc, 32'h42b53504, 32'hc2887864, 32'h426db109, 32'h427b943f, 32'h3ee8a442, 32'hc27687f0, 32'h4239de9c};
test_weights[2920:2927] = '{32'h428c50e2, 32'hc1b2e895, 32'h42b5412e, 32'hc22109e4, 32'h41c0ecd7, 32'h42c522fe, 32'hc22cef37, 32'h4268d031};
test_bias[365:365] = '{32'hc27b12ab};
test_output[365:365] = '{32'hc4996732};
test_input[2928:2935] = '{32'hc19dcdee, 32'hc1f68f62, 32'hc210b35c, 32'h42933593, 32'hc15537b2, 32'hc2187b17, 32'hc2ab788e, 32'hc2c142c6};
test_weights[2928:2935] = '{32'hc24d7b55, 32'hc2b723e1, 32'h426e0fe3, 32'hc2882373, 32'hc2854738, 32'hc0aa7dfd, 32'h429c92f5, 32'h417f2dde};
test_bias[366:366] = '{32'hc0bd0310};
test_output[366:366] = '{32'hc623fe42};
test_input[2936:2943] = '{32'hc2b6de33, 32'h4272bd5b, 32'hc24b6dc5, 32'hc2b3c5d8, 32'hc150fa25, 32'hc2a87614, 32'hc1c66394, 32'hc137861f};
test_weights[2936:2943] = '{32'hc297c0c4, 32'hc2c1f4bb, 32'hc28469e0, 32'h42243649, 32'hc1e14c49, 32'h428493d6, 32'hc2067410, 32'h40729ca2};
test_bias[367:367] = '{32'hc2809541};
test_output[367:367] = '{32'hc56b0598};
test_input[2944:2951] = '{32'h42173848, 32'h428a2fe6, 32'hc2ad2461, 32'h4151682a, 32'hc0ccd332, 32'hc2639214, 32'h4288888d, 32'hc0ff6455};
test_weights[2944:2951] = '{32'hc15bf37d, 32'h41feb18f, 32'h428119d0, 32'h42a3293b, 32'h428b7302, 32'hc17fb2a8, 32'h40d6ac43, 32'h4217769a};
test_bias[368:368] = '{32'h41d9ddc6};
test_output[368:368] = '{32'hc50928ee};
test_input[2952:2959] = '{32'hc25f93ab, 32'h4157ee19, 32'hbcc45c94, 32'h427fbc1e, 32'h41ea84cb, 32'h40f60bac, 32'h42863103, 32'hc24122b0};
test_weights[2952:2959] = '{32'h422e4c2b, 32'h42659b95, 32'h422ca41f, 32'hc2300aa9, 32'h42809a7b, 32'hc281faed, 32'hc0bce356, 32'h411ed28a};
test_bias[369:369] = '{32'hc24795bc};
test_output[369:369] = '{32'hc57af9a8};
test_input[2960:2967] = '{32'h424fa9f5, 32'hc2c1dbda, 32'h421182d8, 32'hc16f14d2, 32'hc1e998e8, 32'h42bcd1f1, 32'hc2655f17, 32'h422b14eb};
test_weights[2960:2967] = '{32'hc210d1c2, 32'h420158fa, 32'h42b7a23e, 32'hc2115f12, 32'h41274ff4, 32'hc23c398b, 32'h425b96b8, 32'h41534791};
test_bias[370:370] = '{32'h424d795e};
test_output[370:370] = '{32'hc6036a57};
test_input[2968:2975] = '{32'hc256b924, 32'h4182debe, 32'hc25a28a3, 32'hc26e0ecf, 32'h42151d06, 32'hc16a46d1, 32'h40c4cc6c, 32'hc1b8d49c};
test_weights[2968:2975] = '{32'h4254fe32, 32'hc289ed7f, 32'hc2137f4f, 32'hc2a05d3d, 32'h42c408b2, 32'h428ed072, 32'hc1e9867c, 32'h423d215a};
test_bias[371:371] = '{32'hc289ac36};
test_output[371:371] = '{32'h457e01ea};
test_input[2976:2983] = '{32'h426cfdc3, 32'h3f86fb5b, 32'h40e1c44b, 32'hc2c09991, 32'hc13b8941, 32'hc22e02f1, 32'hc1c99d70, 32'hc28164e8};
test_weights[2976:2983] = '{32'h421202bb, 32'h419dda77, 32'h42054d4c, 32'hc2b2fce6, 32'h42b089e8, 32'hc2bd34dd, 32'hc1ebb496, 32'hc2aee220};
test_bias[372:372] = '{32'h42ad377d};
test_output[372:372] = '{32'h46a0f84e};
test_input[2984:2991] = '{32'h42968da9, 32'hc2b4b357, 32'h41a167b7, 32'hc2b9a35a, 32'hc22137c6, 32'h42bd293f, 32'hc296ad29, 32'h425e217d};
test_weights[2984:2991] = '{32'h422b0a7f, 32'h4298a758, 32'hc120fb31, 32'h42b49d41, 32'h429f30d8, 32'hc1ceabf4, 32'hc023b5cb, 32'h41eb7f97};
test_bias[373:373] = '{32'hc04b0a87};
test_output[373:373] = '{32'hc67b66bd};
test_input[2992:2999] = '{32'h4021a79c, 32'hc1777d93, 32'hc20da5db, 32'hc0ec3556, 32'h41c3203d, 32'hc237c19e, 32'hc1048a36, 32'hc292b559};
test_weights[2992:2999] = '{32'h41f6cb63, 32'hc1ec5e05, 32'h42a600c8, 32'hc23541e9, 32'h427ce480, 32'h41090c88, 32'hc25abaed, 32'h42220117};
test_bias[374:374] = '{32'h429a01c1};
test_output[374:374] = '{32'hc5522321};
test_input[3000:3007] = '{32'hc23e8804, 32'hc28b7a0a, 32'hc2012a65, 32'h42b15d37, 32'hc2bb98fd, 32'hc27e00c5, 32'h42b6cc29, 32'h41d76ee8};
test_weights[3000:3007] = '{32'hc18497c5, 32'h420de572, 32'h42960a84, 32'h4154825f, 32'hc160b5af, 32'hc24c39ce, 32'h42ad2f07, 32'h424c37ce};
test_bias[375:375] = '{32'h41d36eaa};
test_output[375:375] = '{32'h462b0831};
test_input[3008:3015] = '{32'hc16fa4c1, 32'h422b2ac4, 32'hc299ad07, 32'hc2926498, 32'h41de32d5, 32'hc2b8b3c9, 32'hc133114f, 32'hc23a1321};
test_weights[3008:3015] = '{32'hc275c363, 32'hc2547369, 32'h41e76685, 32'h3fa4fa81, 32'h4223a947, 32'hc23199fe, 32'h41bbd9c0, 32'h42030749};
test_bias[376:376] = '{32'h4213644f};
test_output[376:376] = '{32'hc3365a35};
test_input[3016:3023] = '{32'h4231bd21, 32'h41756e44, 32'h429d08da, 32'hc2ba7d24, 32'hc1d82579, 32'hc2287d98, 32'hc2a51f95, 32'hc278fd64};
test_weights[3016:3023] = '{32'hc09bfeb5, 32'h4266fd45, 32'hc209e6fd, 32'hc276af5f, 32'h4157840d, 32'h418f70cb, 32'hc061d9fa, 32'hc2132d3b};
test_bias[377:377] = '{32'h41ca8ba6};
test_output[377:377] = '{32'h45a284c2};
test_input[3024:3031] = '{32'hc19b2332, 32'hc1d8a765, 32'hc2a7ed1f, 32'h429c1a40, 32'hc28296b2, 32'hc054bcc5, 32'h41238f14, 32'hc2baa06b};
test_weights[3024:3031] = '{32'h42b0d5c8, 32'h4205544b, 32'h42811520, 32'h4238ecc2, 32'hc2c6b463, 32'hc2886701, 32'h3f943550, 32'h42a9bf94};
test_bias[378:378] = '{32'h4216c854};
test_output[378:378] = '{32'hc5ae8403};
test_input[3032:3039] = '{32'hc21a0252, 32'hc20af50f, 32'h42bc0eb9, 32'h4268ff1a, 32'h42be78bc, 32'h40e3e1f0, 32'hc00c04af, 32'h42a8da03};
test_weights[3032:3039] = '{32'hc2b8ab7e, 32'hc1469ea5, 32'hc20ff8c3, 32'hc2a68809, 32'h40079bd4, 32'h42043437, 32'h4187b516, 32'h426af7b0};
test_bias[379:379] = '{32'hc2180d48};
test_output[379:379] = '{32'h4486261f};
test_input[3040:3047] = '{32'h4281fbd9, 32'hc28fdb66, 32'h41c93261, 32'h42c069d1, 32'h42a4cf89, 32'h41e43d5c, 32'hc133f5cc, 32'h41c0b8ed};
test_weights[3040:3047] = '{32'h41b50bab, 32'hc2035119, 32'h41ba7dad, 32'h41de343d, 32'h42a0a606, 32'hc28969b4, 32'hc23e69f0, 32'hc222a70e};
test_bias[380:380] = '{32'hc17da95b};
test_output[380:380] = '{32'h46306641};
test_input[3048:3055] = '{32'h429562ef, 32'h4284ef75, 32'hc23a4b91, 32'hc1d3c593, 32'h411b53a8, 32'hc1b59bca, 32'hc2ad7788, 32'hc1419df9};
test_weights[3048:3055] = '{32'hc2bb1e49, 32'hc2167e9d, 32'hc2b7e559, 32'h42779279, 32'h4165cc29, 32'hc1f7438d, 32'hc240d618, 32'h4180a71c};
test_bias[381:381] = '{32'hc18aa8da};
test_output[381:381] = '{32'hc4fe51a0};
test_input[3056:3063] = '{32'h41df1657, 32'h42081cb9, 32'h42405064, 32'h420338ff, 32'h41c0aec0, 32'h42296e0d, 32'h42ab3629, 32'hc1e5d91d};
test_weights[3056:3063] = '{32'h42157d0d, 32'h4267a088, 32'hc09e0d3f, 32'h4131e428, 32'hc2b1f166, 32'hc22a792b, 32'hc271ac2c, 32'h4028f3e9};
test_bias[382:382] = '{32'h41944e43};
test_output[382:382] = '{32'hc5bcad6c};
test_input[3064:3071] = '{32'hc20b2871, 32'h42599e7d, 32'hc24c1083, 32'hc118dbab, 32'h4214935e, 32'h419d1f6f, 32'hc2587f78, 32'hc24cb58a};
test_weights[3064:3071] = '{32'hc2c77e30, 32'hc1164188, 32'h42a05692, 32'hc1de8387, 32'h41d48ae4, 32'hc252082d, 32'h41c7f15c, 32'hc27a9ab7};
test_bias[383:383] = '{32'hc2af0caa};
test_output[383:383] = '{32'h4456293f};
test_input[3072:3079] = '{32'hc2138af8, 32'h42a8d5b8, 32'h42592db9, 32'hc2a96753, 32'h428b9591, 32'h41ae3139, 32'h40882f21, 32'hc244b6fd};
test_weights[3072:3079] = '{32'hc2039cbb, 32'h42a32c45, 32'h428bd536, 32'h429798d2, 32'h41ab74c0, 32'h42b3127b, 32'h4218cfb5, 32'hc2791c94};
test_bias[384:384] = '{32'h42711bbd};
test_output[384:384] = '{32'h463ebefa};
test_input[3080:3087] = '{32'hc2c270f2, 32'h4154eb66, 32'h42bccc36, 32'hc18eb5fa, 32'h420eaee4, 32'hc2c5aeba, 32'hc045a5c7, 32'hbf8896ac};
test_weights[3080:3087] = '{32'hc29bf57a, 32'hc2797a86, 32'hc2b4b894, 32'hc25d7d6a, 32'h4118d4e7, 32'hc28aac2d, 32'h41380ea6, 32'h422f6579};
test_bias[385:385] = '{32'hc1855868};
test_output[385:385] = '{32'h45c500da};
test_input[3088:3095] = '{32'h3f4d9569, 32'h41e37ebc, 32'hc1d0afaa, 32'h429f6449, 32'h422246ba, 32'h4244d205, 32'hc2774dae, 32'hc2c45f70};
test_weights[3088:3095] = '{32'h413be2b5, 32'h429c7428, 32'hc2a53c84, 32'h403806b9, 32'hc2be2b5a, 32'hc2bb2dcc, 32'hc2a0bd75, 32'hc25027fe};
test_bias[386:386] = '{32'h42a4822a};
test_output[386:386] = '{32'h45c56370};
test_input[3096:3103] = '{32'hc2a798de, 32'h42188a33, 32'h41c3274d, 32'hc1ddf8a6, 32'hc2be1cab, 32'hc187a0e4, 32'h42bac4ca, 32'hc23e018e};
test_weights[3096:3103] = '{32'hc29fbc61, 32'h413dc778, 32'hc1cf9361, 32'hc2990b10, 32'hc2c24b63, 32'hc23bb098, 32'hc1de180f, 32'hc27872a1};
test_bias[387:387] = '{32'hc2877ec5};
test_output[387:387] = '{32'h469416f1};
test_input[3104:3111] = '{32'hc2c3164e, 32'h417f390a, 32'h41b9c57c, 32'h4239f8a5, 32'hc2981e34, 32'hc285e2d4, 32'h428e18fe, 32'hc29cf859};
test_weights[3104:3111] = '{32'h4254afb7, 32'h4243c7ad, 32'hc29785bd, 32'h42c645b8, 32'hc14fa639, 32'h40633488, 32'h40fbb484, 32'hc23f19a3};
test_bias[388:388] = '{32'hc2ad7cbd};
test_output[388:388] = '{32'h45557373};
test_input[3112:3119] = '{32'hc2bb0af8, 32'hc2bbc2d7, 32'h42783e1c, 32'hc2b88357, 32'hc2ba8f18, 32'hc29d0563, 32'hc1bf78f6, 32'h3ffdb1e5};
test_weights[3112:3119] = '{32'hc28f889e, 32'h42509c5f, 32'h421a0020, 32'h42b1891a, 32'h42528bc5, 32'hc244dd74, 32'hc195e531, 32'hc29af68f};
test_bias[389:389] = '{32'hc020640c};
test_output[389:389] = '{32'hc5940fe4};
test_input[3120:3127] = '{32'h42acbbd7, 32'hc0d9faff, 32'hc27cdb3e, 32'h41969bbb, 32'h4209e231, 32'h41e73930, 32'hc2652f4b, 32'hc2a68575};
test_weights[3120:3127] = '{32'h42c4d99c, 32'h4153d7ba, 32'hc2ba0a8e, 32'h4282e866, 32'hc20ba910, 32'h425edd0c, 32'hc29cf698, 32'hc2b5c179};
test_bias[390:390] = '{32'hc1cdfbae};
test_output[390:390] = '{32'h46da7e72};
test_input[3128:3135] = '{32'hc2c4ade2, 32'h42b126b6, 32'hc2271b6c, 32'hc29698d4, 32'h40834859, 32'hc290a09f, 32'hc25dc3c9, 32'h4288936e};
test_weights[3128:3135] = '{32'h422d36bc, 32'h4192d44e, 32'hc053843d, 32'h42ab1974, 32'h42a0bc4e, 32'hc10b6d36, 32'h41c6aae4, 32'hc28957ef};
test_bias[391:391] = '{32'h41999772};
test_output[391:391] = '{32'hc65b1e88};
test_input[3136:3143] = '{32'h42b154d5, 32'hc296639d, 32'h4190f7ed, 32'hc22e89fa, 32'h42befa8e, 32'hc16c3983, 32'h42b28cf1, 32'hc281cb94};
test_weights[3136:3143] = '{32'hc238abeb, 32'hc2624789, 32'h428d9e10, 32'h42be8f24, 32'h426be078, 32'hc243e57a, 32'h428ef96a, 32'h42430252};
test_bias[392:392] = '{32'hc1c98710};
test_output[392:392] = '{32'h45d58656};
test_input[3144:3151] = '{32'hc2938105, 32'h425e01ba, 32'hc29ec0e5, 32'hc2512038, 32'h4249a036, 32'hc264d02e, 32'hc20528ec, 32'h427e9e92};
test_weights[3144:3151] = '{32'hc28d3bc2, 32'h42c4ab9c, 32'hc2520aef, 32'h41cece48, 32'hc21bcd88, 32'hc295693c, 32'hc2328f9e, 32'hc1938669};
test_bias[393:393] = '{32'hc268f949};
test_output[393:393] = '{32'h467aba22};
test_input[3152:3159] = '{32'hc2c7335f, 32'hc1f112b2, 32'h41d6bd6a, 32'hc2bb52a7, 32'hc1f3fecc, 32'h418f3a48, 32'hc2a9f043, 32'h4259fd38};
test_weights[3152:3159] = '{32'hc2bee370, 32'hc2c6e32c, 32'h42981321, 32'hc1b4fd33, 32'h424d2f34, 32'hc24a54b7, 32'h41d194c0, 32'hc2a1146f};
test_bias[394:394] = '{32'h4214284a};
test_output[394:394] = '{32'h45edf536};
test_input[3160:3167] = '{32'h429f079a, 32'h429dcd2e, 32'h42b941c7, 32'hc13bf2b3, 32'h4225dd86, 32'h413beca6, 32'hc22e037a, 32'hc24ce00e};
test_weights[3160:3167] = '{32'h41b89cd3, 32'hc1b800d3, 32'h4271fa13, 32'hc0424f85, 32'h4243adff, 32'h4237efe4, 32'h42aa46f1, 32'h41d23874};
test_bias[395:395] = '{32'hc2510230};
test_output[395:395] = '{32'h45435fc6};
test_input[3168:3175] = '{32'h42a26e00, 32'h42b60842, 32'h42238e73, 32'h421b62ab, 32'h4190ac22, 32'h41e70b22, 32'hc2bc5ad7, 32'h427c5dc9};
test_weights[3168:3175] = '{32'hc1b5c8ab, 32'h406e55c4, 32'h429aac65, 32'hc28e3060, 32'h420988b4, 32'hc25162ea, 32'hc2b219ff, 32'hc2171a87};
test_bias[396:396] = '{32'h4217bd1a};
test_output[396:396] = '{32'h457cd21c};
test_input[3176:3183] = '{32'hc14a8783, 32'h42719d14, 32'h42af63e5, 32'h42215a68, 32'hc270d15b, 32'hc2995e91, 32'hc091db0b, 32'hc2b9776c};
test_weights[3176:3183] = '{32'h420fa554, 32'hc22603fb, 32'h42b650a3, 32'h41314424, 32'h42bbe2a3, 32'hc18c9d9a, 32'h422b6a9a, 32'h42c180f8};
test_bias[397:397] = '{32'hc138f39f};
test_output[397:397] = '{32'hc5fa3b9f};
test_input[3184:3191] = '{32'h42255a51, 32'h41e9b8f3, 32'hc29e4c63, 32'h420679fe, 32'h420fc9ee, 32'hc2c195ee, 32'hc2bf346c, 32'h410c3f91};
test_weights[3184:3191] = '{32'hc2024085, 32'h40e656b2, 32'hc1172fdb, 32'h42a48fd9, 32'hc1773dd3, 32'hc1e3a5cc, 32'hc2090bf1, 32'h42949a0c};
test_bias[398:398] = '{32'hc252e0f8};
test_output[398:398] = '{32'h46040ce7};
test_input[3192:3199] = '{32'hc25b9ba9, 32'hc283eac3, 32'h41e7a89d, 32'hc2364352, 32'hc1936685, 32'hc2b929b6, 32'hc26adf98, 32'h421cae4c};
test_weights[3192:3199] = '{32'h421ede75, 32'hc1a04914, 32'hc1a5fddd, 32'hc209c8eb, 32'h425e741f, 32'h423df739, 32'hc1861de3, 32'hc281d34f};
test_bias[399:399] = '{32'h41b4ca11};
test_output[399:399] = '{32'hc5d5fbb4};
test_input[3200:3207] = '{32'hc1034cc6, 32'h42a613e5, 32'hc2a11cca, 32'h423f2326, 32'h41abd100, 32'hc189d939, 32'hc2b946cb, 32'hc29b992a};
test_weights[3200:3207] = '{32'h3fe1f92a, 32'hc2990281, 32'h416f143b, 32'h422bb7c6, 32'hc2a7a791, 32'h42acf7c5, 32'h413d1aff, 32'h3eeacf06};
test_bias[400:400] = '{32'hc1e12a28};
test_output[400:400] = '{32'hc61bc410};
test_input[3208:3215] = '{32'hc2432e7c, 32'h3fc7ed31, 32'h42c5f85d, 32'hc21df9b4, 32'h42382821, 32'h4280bc0d, 32'hc2267ee3, 32'hc27e476b};
test_weights[3208:3215] = '{32'h42199319, 32'h429c03eb, 32'hc1bfbd21, 32'hc293542d, 32'h4095b47c, 32'h4286da5c, 32'hc234b02b, 32'h42406085};
test_bias[401:401] = '{32'hc0ada51b};
test_output[401:401] = '{32'h4506e346};
test_input[3216:3223] = '{32'h418810a5, 32'hc2a310ec, 32'h4293d6ae, 32'h41a68330, 32'h42ad9526, 32'h42a04255, 32'hc28e3975, 32'hc219855e};
test_weights[3216:3223] = '{32'h42ab36f8, 32'hc28e3cf9, 32'hc245aa8c, 32'hc26c50f5, 32'h40f0c1d1, 32'h41b4f606, 32'h42150f03, 32'hc28b5a8d};
test_bias[402:402] = '{32'hc225c96c};
test_output[402:402] = '{32'h4596a31d};
test_input[3224:3231] = '{32'h423d2358, 32'h4212f1c9, 32'hc2153b44, 32'hc285bdc1, 32'hc268b558, 32'hc2983aaa, 32'hc1a32ade, 32'h42528136};
test_weights[3224:3231] = '{32'hc2bbbc74, 32'hc2c247da, 32'h422ced1e, 32'hc29fbe4c, 32'h40c318ef, 32'hc2743a2b, 32'h429cda3c, 32'h428d8e6d};
test_bias[403:403] = '{32'hc18d1c88};
test_output[403:403] = '{32'h45049506};
test_input[3232:3239] = '{32'hc293ec84, 32'h423ab95c, 32'h415c2bf2, 32'hc255355b, 32'hc1f304a5, 32'hc1898e4e, 32'hc2bbd292, 32'hc2bc0e92};
test_weights[3232:3239] = '{32'hc2571f22, 32'hc214082d, 32'hc2648636, 32'hc2b2688f, 32'h41cc71c7, 32'h42b2b737, 32'hc26849b4, 32'hc2a09f3e};
test_bias[404:404] = '{32'hc2169028};
test_output[404:404] = '{32'h4683d2ee};
test_input[3240:3247] = '{32'h41c96cbd, 32'h42a42b13, 32'hc281f5cb, 32'hc2b5da26, 32'hc2b7119f, 32'h42c3f177, 32'h42303085, 32'hc13ae799};
test_weights[3240:3247] = '{32'hc29fe11b, 32'hc134febd, 32'h4266816a, 32'hc1995b95, 32'hc2187ed3, 32'hc2c188e3, 32'hc2950144, 32'h42bc36a4};
test_bias[405:405] = '{32'hc269a2e1};
test_output[405:405] = '{32'hc67033f3};
test_input[3248:3255] = '{32'hc29f376d, 32'h3fd9376e, 32'hc2b266d1, 32'h420f254e, 32'h42a0c95f, 32'h42bd1168, 32'h425db603, 32'h42bcbaf4};
test_weights[3248:3255] = '{32'hc2a5ce91, 32'hc2561c6e, 32'h4246c0e9, 32'h4271b28e, 32'h42033e21, 32'hc245f470, 32'h41301d18, 32'hc266569d};
test_bias[406:406] = '{32'hc1091491};
test_output[406:406] = '{32'hc5249f6b};
test_input[3256:3263] = '{32'hc2806503, 32'hc2320f26, 32'h429c0ffe, 32'h42b87566, 32'h429ac3f4, 32'hc281adf3, 32'hc225ba65, 32'h422ee3d4};
test_weights[3256:3263] = '{32'hc17e4970, 32'hc2bf85fe, 32'h40e00dd1, 32'hc2832acf, 32'h423b900b, 32'h42a0177b, 32'hc2105db9, 32'hc1c667dc};
test_bias[407:407] = '{32'hc28df482};
test_output[407:407] = '{32'hc4b41c88};
test_input[3264:3271] = '{32'hc24fecfe, 32'h4241d36f, 32'hc24ef8fa, 32'h41927c28, 32'hc1e57ce6, 32'hc002a56c, 32'hc28edd65, 32'h4287b721};
test_weights[3264:3271] = '{32'h42a764be, 32'h41ec0461, 32'hc2baf384, 32'hc252d22f, 32'h42051ce8, 32'h40f2c1f0, 32'h40194505, 32'h42ba167a};
test_bias[408:408] = '{32'h4195dc3f};
test_output[408:408] = '{32'h45bfeecb};
test_input[3272:3279] = '{32'hc1900f62, 32'hc20117cc, 32'h428a54c1, 32'hc1c7fa5a, 32'h40f4eaa5, 32'hc2adce88, 32'hc2a03727, 32'hc1ef33db};
test_weights[3272:3279] = '{32'h4277d90f, 32'hc1ac2451, 32'hc2170b18, 32'hc2702200, 32'h423422f2, 32'h428c9859, 32'hc19fd6ed, 32'h42afa3ca};
test_bias[409:409] = '{32'hc2c7be39};
test_output[409:409] = '{32'hc6039805};
test_input[3280:3287] = '{32'h41b01895, 32'h42c4e3db, 32'h40eb548b, 32'hc2872d1d, 32'hc144a34d, 32'hc1c14cc5, 32'h41186456, 32'h4285391e};
test_weights[3280:3287] = '{32'h429dd8a3, 32'hc0b113ea, 32'hc1f4e43c, 32'h42992437, 32'h42c78959, 32'hc2b88ea8, 32'h40bb026b, 32'hc21b01ac};
test_bias[410:410] = '{32'hc18462db};
test_output[410:410] = '{32'hc5b39462};
test_input[3288:3295] = '{32'hc2ac3469, 32'h42934585, 32'h4235942f, 32'h41098efd, 32'h41262a10, 32'h425a2c89, 32'h4211f446, 32'h42786355};
test_weights[3288:3295] = '{32'h412f6c39, 32'hc0dd5fc9, 32'hc13f8c86, 32'hbf5928bd, 32'hc2172ae7, 32'h427023b4, 32'h422d0cb5, 32'h42045ea5};
test_bias[411:411] = '{32'h3f9cf123};
test_output[411:411] = '{32'h458d04d5};
test_input[3296:3303] = '{32'hc2bd263b, 32'h4229c831, 32'hc21c1c5e, 32'hc1f5dea6, 32'hc0a76a08, 32'h426c7580, 32'h42ba7bd5, 32'h42b6cec7};
test_weights[3296:3303] = '{32'hc19566cf, 32'hc2b22212, 32'h41c402e1, 32'hc2c0a662, 32'hc2bb5132, 32'h42c05108, 32'h42be5f14, 32'hc2c0185d};
test_bias[412:412] = '{32'h42803a3f};
test_output[412:412] = '{32'h45c5a488};
test_input[3304:3311] = '{32'hc11b22ce, 32'hc2a227b9, 32'h41a08d7c, 32'h42c78cb9, 32'h42012b91, 32'hc281cc74, 32'h414fe6e9, 32'h42787d97};
test_weights[3304:3311] = '{32'hbfd1d0e6, 32'hc2c1e5ea, 32'h41c51eee, 32'h41ac3e5e, 32'hc21e1f94, 32'h42aa4330, 32'hc144c163, 32'hc2222dec};
test_bias[413:413] = '{32'h420e7cf4};
test_output[413:413] = '{32'h448651f4};
test_input[3312:3319] = '{32'h41bd4c96, 32'hc0d02cc1, 32'h4284f9ff, 32'h41bd2aee, 32'h4200845b, 32'h428d38c0, 32'hc2af3c0a, 32'h4296f4f6};
test_weights[3312:3319] = '{32'h42848ae8, 32'hc2b15df6, 32'h42c1ef46, 32'h42c64618, 32'hc29a5c5d, 32'h42937bca, 32'hc1c2c1ca, 32'h40184d4d};
test_bias[414:414] = '{32'h42c21b50};
test_output[414:414] = '{32'h467b2560};
test_input[3320:3327] = '{32'h41b89951, 32'hc2af5496, 32'hc27127b7, 32'h4246da11, 32'h4119be4a, 32'hc2891fa6, 32'h4264d5cb, 32'h41ffc4ec};
test_weights[3320:3327] = '{32'hc2a4922a, 32'h42802d92, 32'hc1f218e5, 32'hc271f542, 32'hc2b0e510, 32'h42c22c85, 32'h421203ed, 32'hc29554dd};
test_bias[415:415] = '{32'hc204e4c9};
test_output[415:415] = '{32'hc681343f};
test_input[3328:3335] = '{32'hc21ee6e8, 32'hc20a21a8, 32'h42b545f2, 32'h42a11177, 32'h42c1a07e, 32'h42c25116, 32'h40d81b2f, 32'h41eb57de};
test_weights[3328:3335] = '{32'h42035766, 32'h42bbc038, 32'hc2211fab, 32'h428a31be, 32'h42af5bd9, 32'hc252460d, 32'hc031cf5b, 32'hc18ae4d0};
test_bias[416:416] = '{32'hc1d6f521};
test_output[416:416] = '{32'h434044d7};
test_input[3336:3343] = '{32'h3fa878bf, 32'h41eabc0a, 32'hc2b3df99, 32'h41d312ed, 32'hc1272e9d, 32'hbfd9574f, 32'h40dddd8d, 32'hc2c53dae};
test_weights[3336:3343] = '{32'hc1de4c37, 32'h41ba32c7, 32'hc13dc2b1, 32'h42adbb12, 32'hc23849a0, 32'h42b358a0, 32'hc2981313, 32'hc280ff32};
test_bias[417:417] = '{32'hc024894e};
test_output[417:417] = '{32'h461ed47e};
test_input[3344:3351] = '{32'hc2b80ca5, 32'h417f5e97, 32'h3c764429, 32'hc25de69e, 32'h4205f300, 32'h42992e0d, 32'hc18aff52, 32'hc276d566};
test_weights[3344:3351] = '{32'hc137f6ba, 32'h429b1404, 32'hc13d3031, 32'h424f781e, 32'h42879669, 32'h40ae20b0, 32'h4035daad, 32'h42709927};
test_bias[418:418] = '{32'hc284df98};
test_output[418:418] = '{32'hc4d74da9};
test_input[3352:3359] = '{32'hc2bd9480, 32'hc2a88b2f, 32'hc2491e85, 32'h427599cc, 32'h427762a8, 32'h420998fd, 32'h429f6618, 32'hbfa4b3e4};
test_weights[3352:3359] = '{32'h41623345, 32'h4276f2ad, 32'h41f576ca, 32'h4272546e, 32'hc0011cd9, 32'h4178be71, 32'h412299b2, 32'hc2832d36};
test_bias[419:419] = '{32'hc21584ea};
test_output[419:419] = '{32'hc541ac31};
test_input[3360:3367] = '{32'h412b0c33, 32'h4218ff0f, 32'h4289a642, 32'hc272b8ac, 32'h42bab26d, 32'hc2b2cb88, 32'hc1b3430c, 32'hc222e351};
test_weights[3360:3367] = '{32'h42aa9dfd, 32'hc2455a57, 32'hc1a61b2f, 32'h424c223e, 32'hc13d90ea, 32'h429788db, 32'hc2bdd9f1, 32'hc29360c5};
test_bias[420:420] = '{32'hc2872d5e};
test_output[420:420] = '{32'hc6020035};
test_input[3368:3375] = '{32'h425dc8f3, 32'hc1437494, 32'hc2acbc3c, 32'hc1f07d3c, 32'hc22ad797, 32'h428bbc55, 32'hc090ddfb, 32'hc24cde04};
test_weights[3368:3375] = '{32'hc26ee584, 32'h425bb79a, 32'hc23943d2, 32'hbe8546ff, 32'h4191eaec, 32'hc235f540, 32'hc2bfc1d5, 32'hc0dc1df1};
test_bias[421:421] = '{32'hc187ff7b};
test_output[421:421] = '{32'hc545a5eb};
test_input[3376:3383] = '{32'hc29a240b, 32'h4116494a, 32'hc22dee30, 32'hc245a5cc, 32'h421358ff, 32'h42281b1b, 32'h42683ebd, 32'hc2becc85};
test_weights[3376:3383] = '{32'hc18ed6e8, 32'hc260df60, 32'h4290b4c1, 32'h4200cc00, 32'hc28eaa18, 32'hc175e793, 32'hc2bf29f3, 32'hc28191f6};
test_bias[422:422] = '{32'hbf821693};
test_output[422:422] = '{32'hc5cc2686};
test_input[3384:3391] = '{32'h41ac02b6, 32'h42bd8b3b, 32'h42045b74, 32'h426622f6, 32'hc28c29f2, 32'h42274f1a, 32'hc1736ca8, 32'hc0e77fcd};
test_weights[3384:3391] = '{32'hc289f415, 32'hc21e7406, 32'hc235093e, 32'hc1fd7a9e, 32'hc292f1d5, 32'hc25694dc, 32'hc1222663, 32'hc0d2d3c2};
test_bias[423:423] = '{32'hc0d5abc1};
test_output[423:423] = '{32'hc5aa8bab};
test_input[3392:3399] = '{32'hc25ea0c7, 32'h421cb202, 32'hc218ffd7, 32'h4231e806, 32'h425dd76b, 32'h41db0b37, 32'hc27ed60d, 32'hc18c5188};
test_weights[3392:3399] = '{32'h42aeb5be, 32'hc293965d, 32'hc20b4bba, 32'h42b0eb9b, 32'hc2af18e0, 32'h42c24903, 32'h4200b713, 32'h425f87e1};
test_bias[424:424] = '{32'hc252e963};
test_output[424:424] = '{32'hc5f2a769};
test_input[3400:3407] = '{32'hc2638860, 32'hbff3e9e0, 32'h4244cc5f, 32'h421e3250, 32'hc20510ef, 32'h425d3880, 32'hc184e117, 32'hc282417f};
test_weights[3400:3407] = '{32'h429e1f6f, 32'h4213480d, 32'hc28e01c0, 32'h410a0e13, 32'hbd4fe97b, 32'hc1bada1c, 32'h414b540a, 32'h4260bf75};
test_bias[425:425] = '{32'hc2b609c5};
test_output[425:425] = '{32'hc64aac04};
test_input[3408:3415] = '{32'h4291ab12, 32'hc1abbb34, 32'hc28f3f70, 32'h41de2734, 32'h42af267f, 32'h42a780a0, 32'hc2bea6d2, 32'h42a812f0};
test_weights[3408:3415] = '{32'h42918cd2, 32'h4257426d, 32'h41960a99, 32'h428ad20f, 32'h42c32b8d, 32'hc220fa5c, 32'h428ed8db, 32'h419ef5dc};
test_bias[426:426] = '{32'hc2345eab};
test_output[426:426] = '{32'h4593894c};
test_input[3416:3423] = '{32'h41b42d21, 32'h4229c63c, 32'h428c1f69, 32'hc2be3109, 32'h425fe72d, 32'hc1ecff35, 32'h42bfdc4a, 32'hc21276af};
test_weights[3416:3423] = '{32'hc2008876, 32'hc17cdbc0, 32'h42a4235f, 32'hc2898fcd, 32'h42b52a5e, 32'h41da90b7, 32'h42bbf6c5, 32'hc289aeea};
test_bias[427:427] = '{32'hc26437bb};
test_output[427:427] = '{32'h46d01935};
test_input[3424:3431] = '{32'hc2c60613, 32'h420dc439, 32'hc1ecc67a, 32'hc25730c7, 32'h41d60eec, 32'hc21953b8, 32'h42ac9c4d, 32'h41d6f2bc};
test_weights[3424:3431] = '{32'hc144fe5c, 32'h42748088, 32'hc2104d2b, 32'hc0b48e6d, 32'h41fb2ee6, 32'h421bb1b4, 32'h41af8d82, 32'h42bf19f9};
test_bias[428:428] = '{32'h42bc9455};
test_output[428:428] = '{32'h46075134};
test_input[3432:3439] = '{32'h40f5c80a, 32'hc299638b, 32'h401985ae, 32'hc2829a86, 32'h4222ef4a, 32'hc2b353b0, 32'hc294d998, 32'h424bf76d};
test_weights[3432:3439] = '{32'hc0e978ac, 32'hc22821ff, 32'h42b9ba47, 32'h428daaae, 32'hc2c26d9c, 32'hc27d3b64, 32'hc1c7b2da, 32'h428b5542};
test_bias[429:429] = '{32'h424b00b2};
test_output[429:429] = '{32'h45b9b329};
test_input[3440:3447] = '{32'h42160ed2, 32'hc17e45f3, 32'h41e35722, 32'h42c61533, 32'h41d0b8ef, 32'hc28f005e, 32'h4283e8f9, 32'h41b3e333};
test_weights[3440:3447] = '{32'hc25a9d83, 32'h4183ee35, 32'hc2086326, 32'hc1f71a49, 32'hc096864c, 32'hc2008cf8, 32'hc28f926f, 32'hc28c15c7};
test_bias[430:430] = '{32'h40f21cf7};
test_output[430:430] = '{32'hc6238db4};
test_input[3448:3455] = '{32'hc2752461, 32'hc2b5536a, 32'h41b99540, 32'h42207081, 32'h42bb6e41, 32'h409e3b6a, 32'h42c7bed0, 32'h4247a699};
test_weights[3448:3455] = '{32'h4187bf7c, 32'h41bce73e, 32'h425a9083, 32'hc2a35b01, 32'h425fda42, 32'h41ff7e67, 32'hc21107c6, 32'h41639f56};
test_bias[431:431] = '{32'hc2053d1e};
test_output[431:431] = '{32'hc52ab1d6};
test_input[3456:3463] = '{32'h40043b45, 32'hc27f75d5, 32'hc296f4e4, 32'hc03982cc, 32'h420f4e59, 32'hc194fdaa, 32'h42bb8eed, 32'h4176bc16};
test_weights[3456:3463] = '{32'hc2882cea, 32'h3fc5ced1, 32'h42c0c5a0, 32'hc28d986e, 32'hc2213bb3, 32'h4171f90f, 32'h4238a0f4, 32'h4292af9f};
test_bias[432:432] = '{32'h42bde8e7};
test_output[432:432] = '{32'hc55986a6};
test_input[3464:3471] = '{32'h4242b32e, 32'h42521b36, 32'h41abe36b, 32'h42496a14, 32'hc0c60c32, 32'hc29b63f2, 32'h42b0634d, 32'hc24a1153};
test_weights[3464:3471] = '{32'h42a75d7e, 32'hc17397d0, 32'h42924779, 32'hc2bf1aaa, 32'h42c58a47, 32'hc215eab3, 32'hc219dd77, 32'hc264ba76};
test_bias[433:433] = '{32'h4286627d};
test_output[433:433] = '{32'h44ed359c};
test_input[3472:3479] = '{32'hc22a753a, 32'hc00e1b99, 32'h417154a8, 32'hc2bb88e1, 32'h42231be5, 32'hc241b6a0, 32'h4265a7ab, 32'hc245279c};
test_weights[3472:3479] = '{32'h42b93416, 32'h42af166f, 32'h42573adf, 32'h410f3f02, 32'h42b9b7ae, 32'h4217b920, 32'h41cecc87, 32'hc245c881};
test_bias[434:434] = '{32'hc0faf6a2};
test_output[434:434] = '{32'h44d3d1a4};
test_input[3480:3487] = '{32'hc20bed73, 32'h40fd2ec5, 32'h428ee54e, 32'h423d7366, 32'hc1bd9710, 32'hc2852ddb, 32'h4222ced1, 32'hc24917ae};
test_weights[3480:3487] = '{32'hc1dc9f2a, 32'h42a31517, 32'h41aa3103, 32'hc11b56bc, 32'hc2af6399, 32'hc0856cef, 32'h421439e6, 32'h420ff229};
test_bias[435:435] = '{32'hc2af48d0};
test_output[435:435] = '{32'h4590eb2f};
test_input[3488:3495] = '{32'hc2bead49, 32'hc29c17a7, 32'h41c29cb6, 32'hc2148010, 32'h42b85506, 32'h4214bc31, 32'h42278715, 32'hc288f671};
test_weights[3488:3495] = '{32'h42361ad8, 32'hc23974e2, 32'hc25b44b2, 32'hc198b986, 32'hc18da200, 32'hc2adb7e0, 32'h42849f04, 32'h429d5c2a};
test_bias[436:436] = '{32'hc299ec05};
test_output[436:436] = '{32'hc60affcd};
test_input[3496:3503] = '{32'h42725df8, 32'hc28a7a2b, 32'h4235363b, 32'hc2bf331c, 32'h422aa2ff, 32'hc157c1e0, 32'hc29e2267, 32'hc1e404e8};
test_weights[3496:3503] = '{32'h42b5beb2, 32'h42c5b6e4, 32'h41908365, 32'h424190da, 32'hc1b07f47, 32'hc14b41c2, 32'hc147e842, 32'hc2afe653};
test_bias[437:437] = '{32'hc25d2f2a};
test_output[437:437] = '{32'hc51acf2e};
test_input[3504:3511] = '{32'hc240b121, 32'hbfd206cd, 32'hc21d3d6d, 32'h42acac25, 32'h41a9ebcf, 32'hc184fe03, 32'hc2c102f1, 32'hc2b2424c};
test_weights[3504:3511] = '{32'h429c862f, 32'h4246be56, 32'h41c08d87, 32'h4296ccae, 32'hc23e6f42, 32'hc28b7836, 32'h40330f4e, 32'h41d3f431};
test_bias[438:438] = '{32'hc23026e5};
test_output[438:438] = '{32'hc44bde1b};
test_input[3512:3519] = '{32'h42b09fdc, 32'h42577f92, 32'h42b2eb45, 32'hc267c9db, 32'h4203f611, 32'h408b36db, 32'hc277df87, 32'h42273be1};
test_weights[3512:3519] = '{32'hc2b13c04, 32'h42681e4e, 32'h42a2f428, 32'h4201d1d8, 32'hc285abd3, 32'hc2875a75, 32'hc1142b4c, 32'hc29e2258};
test_bias[439:439] = '{32'h42c61e71};
test_output[439:439] = '{32'hc58a3c71};
test_input[3520:3527] = '{32'hc0e74b79, 32'hc29ee907, 32'hc2b8c7f2, 32'h4297bc97, 32'hc28f4dac, 32'h416f93ba, 32'hc28960b2, 32'hc2825932};
test_weights[3520:3527] = '{32'hc1faa8d9, 32'hc2696f79, 32'h42950eda, 32'h42a737af, 32'h4268c43f, 32'hc243eed1, 32'hc124f539, 32'h414c9d33};
test_bias[440:440] = '{32'h425d99d5};
test_output[440:440] = '{32'hc423012b};
test_input[3528:3535] = '{32'hc287de92, 32'h424d5455, 32'h418e3946, 32'h426562bc, 32'h41e26aeb, 32'hc15d1d2a, 32'h426b3131, 32'hc2b91840};
test_weights[3528:3535] = '{32'h42355744, 32'hc29c947c, 32'hc225135a, 32'h41b44e7c, 32'hc2185393, 32'hc12e0931, 32'h416e9edb, 32'hc209d0dc};
test_bias[441:441] = '{32'h418a5ea8};
test_output[441:441] = '{32'hc55387bf};
test_input[3536:3543] = '{32'hc2445258, 32'hc2444110, 32'hc2823b5a, 32'hc28b12a4, 32'h40860940, 32'hc2035b58, 32'h41c90c26, 32'hc177048d};
test_weights[3536:3543] = '{32'h4291b026, 32'h42a9844c, 32'h419039a4, 32'h4273b87c, 32'h41f5409b, 32'h42983a66, 32'hbef77dcb, 32'hc2483737};
test_bias[442:442] = '{32'h41834a8d};
test_output[442:442] = '{32'hc6664a8a};
test_input[3544:3551] = '{32'h42c2c312, 32'hc21ea80c, 32'h4209666c, 32'hc10b8993, 32'h40d3586d, 32'hc16581b7, 32'h417186a4, 32'h428efee3};
test_weights[3544:3551] = '{32'hc257ffd3, 32'hc25ae40d, 32'h40a51c13, 32'hc2bf5155, 32'hc1b21473, 32'hc222fcda, 32'h420645b3, 32'hc2966761};
test_bias[443:443] = '{32'hc2ab1160};
test_output[443:443] = '{32'hc5ce1556};
test_input[3552:3559] = '{32'h42afa532, 32'h42600908, 32'h413190b0, 32'h427d0ec8, 32'hc28d4886, 32'h41c0a442, 32'h42af2922, 32'hc2b0474a};
test_weights[3552:3559] = '{32'hc2234dc9, 32'hc287f81d, 32'h4259a1f9, 32'h420452e3, 32'h4203be16, 32'h42bf60ad, 32'h42bbe525, 32'h42a031c1};
test_bias[444:444] = '{32'h42a362aa};
test_output[444:444] = '{32'hc558cfef};
test_input[3560:3567] = '{32'h4286a63a, 32'hc2c0930e, 32'h424892c3, 32'h41b8e2d4, 32'hc25caae1, 32'h4278b0f1, 32'h41dd15b1, 32'hc2b1b109};
test_weights[3560:3567] = '{32'h41da5c12, 32'hc21f28f0, 32'hc2bac861, 32'hc2622367, 32'h424a48d1, 32'h3f24d229, 32'h4204f5b6, 32'h42a70b60};
test_bias[445:445] = '{32'h41a64982};
test_output[445:445] = '{32'hc6153e96};
test_input[3568:3575] = '{32'hc292da1d, 32'h40b1d990, 32'h42b6ef36, 32'hc2c6d7ae, 32'hc2695595, 32'h42453c81, 32'h42175910, 32'h417658cc};
test_weights[3568:3575] = '{32'hc2b02fc8, 32'h420519f1, 32'hc2809740, 32'h42b42d0a, 32'h4277a92d, 32'h42967542, 32'hc247c155, 32'h41f0a61a};
test_bias[446:446] = '{32'hc1c220be};
test_output[446:446] = '{32'hc61504da};
test_input[3576:3583] = '{32'hc21c896d, 32'h42868702, 32'h419e05a2, 32'hc0f3190d, 32'hbf33a842, 32'hc2aae852, 32'hc2c19d93, 32'h424ca62d};
test_weights[3576:3583] = '{32'hc2075bb3, 32'h42b955c4, 32'h415ca3bc, 32'h42a3daa4, 32'h4204ae65, 32'h4160908b, 32'hc0fd0a8f, 32'hc21f8fed};
test_bias[447:447] = '{32'h411e6730};
test_output[447:447] = '{32'h45937a93};
test_input[3584:3591] = '{32'h42ac2846, 32'hc00d20f5, 32'h41e6cb71, 32'h42666db7, 32'hc2174728, 32'hbfb3662f, 32'hc27a4e81, 32'h4216610a};
test_weights[3584:3591] = '{32'h42c7768b, 32'hc29c8d42, 32'hc191735e, 32'h42b8f536, 32'hc21cc914, 32'hc29f49bb, 32'hc2ac9128, 32'hc2819924};
test_bias[448:448] = '{32'h404b1c3e};
test_output[448:448] = '{32'h468d9169};
test_input[3592:3599] = '{32'hc250b6a5, 32'hc1e2f1cf, 32'h4296faa9, 32'hc29ccd14, 32'h42512876, 32'h42a5388e, 32'h42a26882, 32'hc278de8f};
test_weights[3592:3599] = '{32'hc26f5cbd, 32'hc282c732, 32'h41e4ad59, 32'h4225d9fc, 32'h41e487d1, 32'hc26bdd0d, 32'h42963fb8, 32'h42c45de8};
test_bias[449:449] = '{32'h419883da};
test_output[449:449] = '{32'h440170ec};
test_input[3600:3607] = '{32'h422129b0, 32'h41ef248e, 32'h424287fc, 32'h42846dac, 32'h42baa48d, 32'hc21cd275, 32'hc256ac65, 32'h421874b7};
test_weights[3600:3607] = '{32'hc257fa02, 32'hc29c25b5, 32'h40d08267, 32'h413070d8, 32'h42b18c8b, 32'hbf9dd13f, 32'hc2ab1a76, 32'h423129ee};
test_bias[450:450] = '{32'h428b2377};
test_output[450:450] = '{32'h462f4f01};
test_input[3608:3615] = '{32'h42bca207, 32'hc139f8a7, 32'hc29baf27, 32'hc1b2b1f9, 32'hc228cea9, 32'hbef35b3d, 32'h41766f24, 32'hc01457d8};
test_weights[3608:3615] = '{32'h42a30c22, 32'h3fcf877a, 32'h41abbd3d, 32'h421313ed, 32'hc2c2cc41, 32'h42899c91, 32'hbff88c60, 32'hc2641e5b};
test_bias[451:451] = '{32'hc1b832e1};
test_output[451:451] = '{32'h4611db0b};
test_input[3616:3623] = '{32'hc14ccb83, 32'hc1b273a7, 32'hc2475a9d, 32'hc2637f07, 32'hc1866bb6, 32'h41a473b0, 32'h42942daf, 32'h42bf1e2d};
test_weights[3616:3623] = '{32'hbe897baa, 32'hc2a5ee76, 32'hc207770b, 32'h421479f1, 32'h42a12736, 32'hc0fe8e20, 32'hbeb8718b, 32'hc2a48efc};
test_bias[452:452] = '{32'hc225bd7d};
test_output[452:452] = '{32'hc5fa89ca};
test_input[3624:3631] = '{32'h42bf3e11, 32'hc2366d28, 32'h423baa51, 32'hc29415d4, 32'hc131333b, 32'hc0fd6a87, 32'hc099601b, 32'h42293f88};
test_weights[3624:3631] = '{32'h4213025a, 32'h41d0093e, 32'h425f8ac1, 32'hbfc1965e, 32'h412aec79, 32'hc2be8abc, 32'hc1c761a0, 32'h42b0e2dc};
test_bias[453:453] = '{32'hc210beb0};
test_output[453:453] = '{32'h4614cf8b};
test_input[3632:3639] = '{32'hc276f0c1, 32'hc22669f7, 32'h423e1252, 32'hc25f3c69, 32'h4299fbfb, 32'h42887e59, 32'hc051fa1f, 32'hbfa7530b};
test_weights[3632:3639] = '{32'hc287615a, 32'h42432563, 32'hc1e1f195, 32'h4218fed7, 32'h42935c5f, 32'hc2749321, 32'h41effab2, 32'hc1429e61};
test_bias[454:454] = '{32'hc188060d};
test_output[454:454] = '{32'h4291da64};
test_input[3640:3647] = '{32'hc1ca3681, 32'h4278b1ba, 32'h429dd8a6, 32'hc27d39ac, 32'h40096067, 32'hc24dec6a, 32'hc28638f5, 32'h421c7a74};
test_weights[3640:3647] = '{32'hc270bbd9, 32'h41ee2168, 32'hc267a1f3, 32'hc2b24b20, 32'h4232071e, 32'h414ac151, 32'hc1c0b472, 32'hc2c2e716};
test_bias[455:455] = '{32'hc2b2948f};
test_output[455:455] = '{32'h44c86bad};
test_input[3648:3655] = '{32'hc2c452e0, 32'h4226e795, 32'hc2ba6839, 32'hc2912cfa, 32'h4207c65d, 32'hc0dda9ad, 32'hc24c5118, 32'h428c0263};
test_weights[3648:3655] = '{32'h41f7da92, 32'h4213818f, 32'hc18b3e96, 32'h42036ca2, 32'hc2b198c4, 32'h41864978, 32'h4122087f, 32'h4249f035};
test_bias[456:456] = '{32'hc2bcc4e8};
test_output[456:456] = '{32'hc51a9225};
test_input[3656:3663] = '{32'hc0ef035e, 32'h41ca74f1, 32'h426c5a93, 32'h42632dcf, 32'h41d29e0a, 32'h42223e14, 32'h429d3940, 32'hc20634ec};
test_weights[3656:3663] = '{32'h42709101, 32'h4152f6c7, 32'hc29954a9, 32'h429536c5, 32'hc205e71b, 32'h4129423e, 32'h4050939a, 32'hc28922c3};
test_bias[457:457] = '{32'h41321c14};
test_output[457:457] = '{32'h44d56bf4};
test_input[3664:3671] = '{32'hc2896da6, 32'hc0d7554a, 32'hc1ab5f1c, 32'hc128e4e7, 32'hc2bbda2d, 32'h417536e2, 32'hc28186b6, 32'h42307e8f};
test_weights[3664:3671] = '{32'h4206fafb, 32'hc282325e, 32'hc087e192, 32'h41b755f4, 32'hc26e57c5, 32'hc2af2b88, 32'h420aca23, 32'hc26ba866};
test_bias[458:458] = '{32'h41084709};
test_output[458:458] = '{32'hc52376e7};
test_input[3672:3679] = '{32'h4201fe81, 32'h429b40af, 32'h427b2efc, 32'h42b97257, 32'h42b6872b, 32'h42884406, 32'h42915c40, 32'hc21454f6};
test_weights[3672:3679] = '{32'hc24ce6d9, 32'h412d2267, 32'h428f8a91, 32'hc21d751d, 32'hc20ff18b, 32'h41dba11d, 32'hc1a9438d, 32'hc2928c1b};
test_bias[459:459] = '{32'h42804b9c};
test_output[459:459] = '{32'hc309fdf7};
test_input[3680:3687] = '{32'hc269f688, 32'hc2114d90, 32'hc1b24020, 32'h41855d0b, 32'h4297a72c, 32'hc282d7b9, 32'h42685632, 32'hc245e6f6};
test_weights[3680:3687] = '{32'hc292aa23, 32'hc10d396d, 32'hc2a0e3cf, 32'hc2a067ee, 32'hc29ac67c, 32'hc2c35478, 32'hc1af1b07, 32'hc28167ed};
test_bias[460:460] = '{32'hc29addee};
test_output[460:460] = '{32'h45e87869};
test_input[3688:3695] = '{32'hc2b30660, 32'hc10ca6c6, 32'h4210c487, 32'hc2b695a5, 32'h409ca2b7, 32'hc01e3d93, 32'hc21976ee, 32'h41873be8};
test_weights[3688:3695] = '{32'hc2716e63, 32'hc2471373, 32'hc0019637, 32'h4263e08b, 32'hc2b907e9, 32'hc2745a8e, 32'hc21261ca, 32'hc2beb62d};
test_bias[461:461] = '{32'hc1d4b4c4};
test_output[461:461] = '{32'h41eed835};
test_input[3696:3703] = '{32'hc2b100c0, 32'h427887df, 32'h42b4e061, 32'h41a6ba29, 32'h409317a0, 32'h4209e2fb, 32'hc094bd56, 32'hc2a7ca5e};
test_weights[3696:3703] = '{32'hc27d260a, 32'h42be4d94, 32'hc13f9e07, 32'hc2353aaf, 32'hc29e498a, 32'h41e155ef, 32'hc2ac8116, 32'hc0f038b0};
test_bias[462:462] = '{32'hc28a03de};
test_output[462:462] = '{32'h462cba32};
test_input[3704:3711] = '{32'h401533ae, 32'h417eb71d, 32'hc2ae60ab, 32'hc1b072fd, 32'hc2111105, 32'h42c13e6a, 32'h4286c598, 32'h4137bd05};
test_weights[3704:3711] = '{32'h42998c87, 32'hc07cfd16, 32'h42c4baac, 32'h427bb1d7, 32'hc2095957, 32'hc1f97681, 32'hc2195490, 32'h4200c3b4};
test_bias[463:463] = '{32'hc17a64d4};
test_output[463:463] = '{32'hc6585332};
test_input[3712:3719] = '{32'h42b2d638, 32'h420c7948, 32'h421b5f92, 32'hc23a2213, 32'h42366cf2, 32'hc27cd549, 32'hc2251510, 32'hc244be54};
test_weights[3712:3719] = '{32'h4293b94e, 32'h423e05be, 32'h41d216a6, 32'hc13dbd20, 32'hc029c70b, 32'hc1e48847, 32'hc1814fa3, 32'hc0e39bf6};
test_bias[464:464] = '{32'hc19e389c};
test_output[464:464] = '{32'h4643ba9a};
test_input[3720:3727] = '{32'h419941d7, 32'hbfe58d8d, 32'hc17836d4, 32'h4258a4c0, 32'hc29a5848, 32'h4256b9a6, 32'h4276f296, 32'h4298d230};
test_weights[3720:3727] = '{32'h41acb766, 32'hc28449d7, 32'h422bd1d2, 32'h42a0b528, 32'h4251d01f, 32'hc28a9835, 32'h4255cdca, 32'hc1089bf4};
test_bias[465:465] = '{32'hc1c0cac0};
test_output[465:465] = '{32'hc467a8da};
test_input[3728:3735] = '{32'h426e19c5, 32'h42aadfae, 32'h4282e1ba, 32'hc14c8325, 32'hc296c450, 32'h40447dfc, 32'h42abf3ed, 32'h40d2f317};
test_weights[3728:3735] = '{32'h41bbe5b8, 32'hc252ea93, 32'h429d31a8, 32'h42b448d1, 32'h40ba4f7b, 32'hc28b1b52, 32'hc283e7fb, 32'hc16f0990};
test_bias[466:466] = '{32'h4212ed03};
test_output[466:466] = '{32'hc5abe239};
test_input[3736:3743] = '{32'hc26e25f3, 32'h418eb9b1, 32'h42289eee, 32'h428d45a8, 32'hc26b4a7d, 32'h426c4a8f, 32'hc263499d, 32'h4129e57f};
test_weights[3736:3743] = '{32'h41e231e2, 32'h40147974, 32'h424ddd9e, 32'hc137bd7a, 32'hc2035fd5, 32'h42ba893e, 32'h42935b5b, 32'hc2c3cc35};
test_bias[467:467] = '{32'hc1550f93};
test_output[467:467] = '{32'h44efd27b};
test_input[3744:3751] = '{32'hc2a75181, 32'h427f22f7, 32'h42c00c7c, 32'h418a5b46, 32'h40c1d80d, 32'h418d9ae9, 32'hc2a7fb60, 32'h4234f76e};
test_weights[3744:3751] = '{32'hc26796df, 32'h3fef140d, 32'h40a17b39, 32'hc2106998, 32'h4268fa24, 32'hc2232170, 32'hc2c5d657, 32'h42adcafb};
test_bias[468:468] = '{32'hc1e1bdd5};
test_output[468:468] = '{32'h46823296};
test_input[3752:3759] = '{32'h42372a96, 32'h42a001e9, 32'h41f5a28c, 32'hc21b90bb, 32'hc292c68d, 32'hc0deee9b, 32'hc1116f7a, 32'hc278abea};
test_weights[3752:3759] = '{32'hc15c2deb, 32'h4296ee6d, 32'h42356f3b, 32'h41fd6be2, 32'hc2a5c808, 32'hc2adfa56, 32'h423e9338, 32'hc28f668e};
test_bias[469:469] = '{32'hc25eb65f};
test_output[469:469] = '{32'h467d8802};
test_input[3760:3767] = '{32'hc2a7b1b4, 32'hc297ad5b, 32'hc2151011, 32'hc1f903cf, 32'hc2b98183, 32'h422b005f, 32'hc18a6f43, 32'hc2ba8ec6};
test_weights[3760:3767] = '{32'hc119463f, 32'h4006b0c5, 32'hc28f00ad, 32'h4278c015, 32'hc2ae6371, 32'hc2894f06, 32'hc1a27934, 32'hc2814bd6};
test_bias[470:470] = '{32'hc24284c8};
test_output[470:470] = '{32'h4648e862};
test_input[3768:3775] = '{32'h4203371b, 32'h42431fe6, 32'hc0f8d4bc, 32'hc1abea83, 32'h428ec06b, 32'hc2364774, 32'hc2199692, 32'hc244e57b};
test_weights[3768:3775] = '{32'hc22eb8c2, 32'h4269b2d2, 32'hc285b8cd, 32'h423b3594, 32'h42400f01, 32'hc010b591, 32'hc2950707, 32'hc2c39c83};
test_bias[471:471] = '{32'hc2c237f5};
test_output[471:471] = '{32'h463c1f35};
test_input[3776:3783] = '{32'h42ad18d5, 32'hc27097e4, 32'hc27fd68e, 32'h426fc36a, 32'h42a87270, 32'h40d6a015, 32'h42a39cd5, 32'hc1af954a};
test_weights[3776:3783] = '{32'h4244f852, 32'h4200ff89, 32'h42b0e00d, 32'hc24b56cf, 32'h4289bb58, 32'h427602fc, 32'hc2687062, 32'h424ddaeb};
test_bias[472:472] = '{32'hc1db4b91};
test_output[472:472] = '{32'hc5bdfb8f};
test_input[3784:3791] = '{32'hc215498c, 32'hc24b428c, 32'h42acb23b, 32'h40e5e409, 32'hc1185ddd, 32'hc21585dd, 32'hc2a86849, 32'h425ece56};
test_weights[3784:3791] = '{32'hc26d1f82, 32'hc283454a, 32'h41a319d6, 32'h42871449, 32'hc21ed59f, 32'hc25be509, 32'hc2c2dd5c, 32'hc2b16597};
test_bias[473:473] = '{32'hc2205209};
test_output[473:473] = '{32'h465227a6};
test_input[3792:3799] = '{32'hc1e4517a, 32'h4223b53f, 32'h42a0d212, 32'hc2bc9efc, 32'h40c4cefe, 32'h42b13ac1, 32'h3e154074, 32'h418a9394};
test_weights[3792:3799] = '{32'hc2c2f489, 32'hc2b62e06, 32'hc1e88a67, 32'hc1a239b7, 32'hc10c7ebd, 32'hc1deb653, 32'h41e3659d, 32'hc1ccf649};
test_bias[474:474] = '{32'hc1edc0c3};
test_output[474:474] = '{32'hc5884a10};
test_input[3800:3807] = '{32'h40ea7a26, 32'hc2b2068b, 32'hc22f7f7c, 32'hc04d8793, 32'hc05a7a03, 32'hc0e49340, 32'hc1385082, 32'hc281e9b3};
test_weights[3800:3807] = '{32'hc2031424, 32'h42075e02, 32'hc0d00aa8, 32'hc26cdd3e, 32'hc1a4446d, 32'h42385df9, 32'h42862718, 32'h42b5dca8};
test_bias[475:475] = '{32'hc2bff4ed};
test_output[475:475] = '{32'hc6194db5};
test_input[3808:3815] = '{32'h4226a851, 32'hc0edc8c6, 32'hc2703856, 32'hc21ede65, 32'hc2618cf7, 32'hc281a78f, 32'h428708a3, 32'hc18e0a6a};
test_weights[3808:3815] = '{32'h41945433, 32'hc24a5820, 32'h42bd3cc6, 32'h42ae95be, 32'h425d3f6e, 32'hc19a7f21, 32'hc2b829c1, 32'hc2b434f5};
test_bias[476:476] = '{32'h423fdeab};
test_output[476:476] = '{32'hc66194cd};
test_input[3816:3823] = '{32'h42763c07, 32'hc2411d93, 32'hc2556ef4, 32'h422164f2, 32'hc23b0597, 32'hc293bab1, 32'h416a198c, 32'hc2b322c7};
test_weights[3816:3823] = '{32'hc2a0c84b, 32'h4292448f, 32'hc25f53ba, 32'hc26cc2f4, 32'h41a434e6, 32'h41daf385, 32'hc296f704, 32'h42615412};
test_bias[477:477] = '{32'h41e2ee20};
test_output[477:477] = '{32'hc684bf40};
test_input[3824:3831] = '{32'hc2967e07, 32'hc25ad131, 32'hc246583f, 32'hc1889573, 32'h42a91834, 32'h424a853e, 32'h42a4a703, 32'h40c84771};
test_weights[3824:3831] = '{32'h42c0cd0a, 32'h41ced2ca, 32'hc1872c32, 32'h42246d06, 32'hc280a17b, 32'hc1e19fc0, 32'hc1a7cc2d, 32'hc2c2e4b8};
test_bias[478:478] = '{32'h4143fdbc};
test_output[478:478] = '{32'hc68a740c};
test_input[3832:3839] = '{32'h4283ed07, 32'hc235b4ec, 32'h4239d7b5, 32'hc238f068, 32'h4211082e, 32'h4281f0c6, 32'h423755ec, 32'hc032e1d5};
test_weights[3832:3839] = '{32'hc1da6a5c, 32'hc22a57ab, 32'h4257192f, 32'h42aa35c2, 32'h41870893, 32'h41fc7b5b, 32'hc21edc00, 32'hc1e6f276};
test_bias[479:479] = '{32'h411b9226};
test_output[479:479] = '{32'hc3b918c1};
test_input[3840:3847] = '{32'hc2b25fd3, 32'h42c4e39c, 32'h42c31946, 32'hc2a3f3ed, 32'h42607f44, 32'h41e33e35, 32'h42824013, 32'hc12bff93};
test_weights[3840:3847] = '{32'hc1745d65, 32'h4291996a, 32'hc2bdad13, 32'h417524e4, 32'h41d97882, 32'h42b9386c, 32'hc2bf6edb, 32'hc29d3b10};
test_bias[480:480] = '{32'hc20ec803};
test_output[480:480] = '{32'hc54ae5dd};
test_input[3848:3855] = '{32'hc1ada1cb, 32'hc0dde0c6, 32'h42bec613, 32'h426ef805, 32'hc1ec650e, 32'h408c95f2, 32'hc2bcea60, 32'h428297b0};
test_weights[3848:3855] = '{32'hc2ba2f85, 32'hc0ab4a90, 32'hc2a1d6ba, 32'h41fe8f7f, 32'h42473b66, 32'h42ac4aec, 32'hc2b47e8d, 32'h42c77c92};
test_bias[481:481] = '{32'hc2add563};
test_output[481:481] = '{32'h461dc47e};
test_input[3856:3863] = '{32'h429ccc0e, 32'hc1a04d7c, 32'hc2999266, 32'hc1f411f2, 32'hc2a2dc5b, 32'hc21383b4, 32'hc19f4657, 32'hc2969ca4};
test_weights[3856:3863] = '{32'h428e33d2, 32'hc2ba2091, 32'hc18a0f1c, 32'hc289b0c4, 32'h419635a3, 32'h421ecd24, 32'hc29982c0, 32'h42989a76};
test_bias[482:482] = '{32'h429f0fd9};
test_output[482:482] = '{32'h45695324};
test_input[3864:3871] = '{32'h41f3f682, 32'hc1ccfa02, 32'h42a5f1ff, 32'hc1937cea, 32'hc1a3dd39, 32'h425bc775, 32'hc28923f4, 32'h4294300e};
test_weights[3864:3871] = '{32'hc1c9c83b, 32'hc2abfab8, 32'h42af08f2, 32'hc27c398d, 32'h42a0cec6, 32'hc2c507d2, 32'hc2a3152d, 32'hc2bef72d};
test_bias[483:483] = '{32'hc2b7b9f9};
test_output[483:483] = '{32'h4498e1fb};
test_input[3872:3879] = '{32'hc2995637, 32'hc2287a18, 32'hc21a1524, 32'h422391e7, 32'h42bf37bd, 32'hc1bdf93d, 32'h42849cae, 32'h4284b0e2};
test_weights[3872:3879] = '{32'h42acea4a, 32'h42743afc, 32'h428c3231, 32'h42871d86, 32'h42922019, 32'hc24f91d3, 32'hc22ac17b, 32'hc1f9d7be};
test_bias[484:484] = '{32'h42b47f38};
test_output[484:484] = '{32'hc5b32395};
test_input[3880:3887] = '{32'hc126cca7, 32'hc00db9e1, 32'hc29e20b5, 32'hc065d70e, 32'h4243cfe8, 32'h41e81617, 32'hc0786a24, 32'h42133f42};
test_weights[3880:3887] = '{32'h40c0fc49, 32'hc13743f3, 32'hc09bcceb, 32'hc272b8da, 32'h419f026d, 32'h4283611f, 32'hc281d450, 32'h42644bd2};
test_bias[485:485] = '{32'h41f0b473};
test_output[485:485] = '{32'h45b618ec};
test_input[3888:3895] = '{32'h4259fb0e, 32'h424d7cdf, 32'h42c57b35, 32'h42b5df4c, 32'h42913728, 32'h417d4260, 32'h426b632e, 32'hc2213c98};
test_weights[3888:3895] = '{32'h42bef8f7, 32'h42832a78, 32'hc2995da4, 32'hc1cbba9c, 32'hc2248f70, 32'hc2695799, 32'hc2b56281, 32'h4201b4eb};
test_bias[486:486] = '{32'hc29abdd2};
test_output[486:486] = '{32'hc63aaaee};
test_input[3896:3903] = '{32'h42a4a0a7, 32'hc0a909a4, 32'hc27ba92f, 32'h40938937, 32'h422695f6, 32'hc290d6a4, 32'hc2130a7b, 32'h41996fe9};
test_weights[3896:3903] = '{32'h42202e8d, 32'hc1c1fac9, 32'hc2c0479c, 32'hc26942a2, 32'hc2028a09, 32'hc1a987c5, 32'h41e9e319, 32'h42b66af5};
test_bias[487:487] = '{32'hc1379943};
test_output[487:487] = '{32'h461ceb7d};
test_input[3904:3911] = '{32'h429829c7, 32'hc0bdd83c, 32'hc1fe2ca2, 32'h4208eb70, 32'hc2472d7b, 32'hc0829c79, 32'h42a3f451, 32'h42c12148};
test_weights[3904:3911] = '{32'h42bc0c88, 32'h4282f3cd, 32'h4075f3d6, 32'h4254e61d, 32'h42509007, 32'h4227463c, 32'h423fe51d, 32'hc20eb7fd};
test_bias[488:488] = '{32'hc27b2f05};
test_output[488:488] = '{32'h45bf534c};
test_input[3912:3919] = '{32'hc09e2f1f, 32'h4247947f, 32'h428e345e, 32'h4230463c, 32'hc0c648b7, 32'h4252e582, 32'hc28f5890, 32'h421d7d1c};
test_weights[3912:3919] = '{32'hc23e5183, 32'h423cba99, 32'h42c42284, 32'hc13e8220, 32'hc235fd18, 32'h4283452f, 32'h426cae41, 32'h423f8407};
test_bias[489:489] = '{32'hc1f9b1c6};
test_output[489:489] = '{32'h462263a8};
test_input[3920:3927] = '{32'h4265de15, 32'h42bb6fe6, 32'h424dd2e7, 32'hc2344977, 32'h42bbc044, 32'hc2b19652, 32'hc104dc6e, 32'h42b5f966};
test_weights[3920:3927] = '{32'hc224b323, 32'hc276eed8, 32'hc2c2dcde, 32'hc1cc434e, 32'h4270a29e, 32'h41e56f6e, 32'h41871675, 32'hc2329512};
test_bias[490:490] = '{32'hc077267d};
test_output[490:490] = '{32'hc64cfee1};
test_input[3928:3935] = '{32'hc2319a55, 32'h42a0d19e, 32'hc2a4b2e4, 32'h42a4d511, 32'hc06e8e8c, 32'h41da8230, 32'h4244f186, 32'h3fdd8412};
test_weights[3928:3935] = '{32'hc1da6443, 32'hc28fe1f3, 32'h4211ba0b, 32'hc2c66553, 32'h42086124, 32'hc1a8b93c, 32'hc284a116, 32'hc29c6c68};
test_bias[491:491] = '{32'hc081c2ec};
test_output[491:491] = '{32'hc69b1fd1};
test_input[3936:3943] = '{32'h422cd2c4, 32'hc1a79d56, 32'h42aa1696, 32'hc0d83692, 32'hc2b4ce93, 32'h4249cfef, 32'hc24fcbd4, 32'h421b77e5};
test_weights[3936:3943] = '{32'h422f1bab, 32'hc2a8c831, 32'hc28b4269, 32'h42a46b59, 32'h4291cd4b, 32'h418e0bc1, 32'hbfe22f21, 32'h4297dc53};
test_bias[492:492] = '{32'hc08020ed};
test_output[492:492] = '{32'hc5ab096a};
test_input[3944:3951] = '{32'hc23b0797, 32'h41b86f9c, 32'hc09dc280, 32'h4237cf38, 32'hc1c63a5e, 32'h427aaf29, 32'hc1f17a46, 32'hc2aea241};
test_weights[3944:3951] = '{32'hc2bccd66, 32'h421099cc, 32'hc177da10, 32'hc27c6090, 32'h42ba32fd, 32'h411335b5, 32'h4274ceb1, 32'h41abdd0b};
test_bias[493:493] = '{32'hc2005b4b};
test_output[493:493] = '{32'hc53f51ca};
test_input[3952:3959] = '{32'h42b329f7, 32'hc297f49f, 32'h42445dc1, 32'hc248a514, 32'h4124efe3, 32'h4280c571, 32'h40f827c3, 32'hc1cefee5};
test_weights[3952:3959] = '{32'hc1110d1d, 32'h4213b77c, 32'h4277cf17, 32'hc26612e1, 32'h427c6c79, 32'hc20c8555, 32'hc2b4d1bd, 32'hc1ad9424};
test_bias[494:494] = '{32'h413db709};
test_output[494:494] = '{32'h440e5a0c};
test_input[3960:3967] = '{32'h429aa3f1, 32'hc269db60, 32'h40501ddd, 32'hc2bfa4b2, 32'hc2008060, 32'h429d6546, 32'hc2929e7e, 32'h41e5aa96};
test_weights[3960:3967] = '{32'h420cad62, 32'h3f778f7a, 32'hc2187893, 32'hc0a56b85, 32'h41df6401, 32'h4267320a, 32'h4295b62e, 32'hc14d1a61};
test_bias[495:495] = '{32'hc28eaa11};
test_output[495:495] = '{32'h443daf53};
test_input[3968:3975] = '{32'hc1c3db35, 32'h41bd6be8, 32'h3f1c4695, 32'h42ab5c06, 32'h4259476f, 32'hc21f005a, 32'hc2408dba, 32'hc117d577};
test_weights[3968:3975] = '{32'h41fb2b38, 32'hc269f0ef, 32'h424c5d56, 32'h426c3bc6, 32'h4293fbeb, 32'hc26c5b82, 32'h41d41177, 32'h428593fb};
test_bias[496:496] = '{32'h42953f78};
test_output[496:496] = '{32'h45e97539};
test_input[3976:3983] = '{32'hc29a69c3, 32'h4265f992, 32'hc225da8c, 32'h4244f603, 32'h42a0f575, 32'h41c6005b, 32'hc1f976a5, 32'h42511998};
test_weights[3976:3983] = '{32'h40c41b1c, 32'hc28b3b4f, 32'hc2ab1d53, 32'h40f18039, 32'hc28df107, 32'h411ae368, 32'h42b30333, 32'hc260fe15};
test_bias[497:497] = '{32'hc17b0a7c};
test_output[497:497] = '{32'hc637fee9};
test_input[3984:3991] = '{32'hc1fbd1fe, 32'hc26109da, 32'h42a95c0f, 32'h424b8794, 32'h42753abb, 32'hc23d0ed9, 32'h42193be8, 32'hc2885934};
test_weights[3984:3991] = '{32'hc1cac68d, 32'hc0cb35e6, 32'hc1c69764, 32'hc2b20625, 32'h42444359, 32'h42123112, 32'h416a03dc, 32'hc2357166};
test_bias[498:498] = '{32'h410c42b8};
test_output[498:498] = '{32'hc4057b9e};
test_input[3992:3999] = '{32'h4186c1bd, 32'h41ab88e5, 32'hc26e80b8, 32'h422484fc, 32'hc2b4e536, 32'h41f6547c, 32'h42864688, 32'h42843414};
test_weights[3992:3999] = '{32'hc1e1a204, 32'hc2954661, 32'h428bb087, 32'hc2ac924d, 32'hc25a0947, 32'hc29fbda1, 32'h42997337, 32'hc2c5b9f6};
test_bias[499:499] = '{32'h4117f636};
test_output[499:499] = '{32'hc607d190};
test_input[4000:4007] = '{32'h42a680d2, 32'h422cbc21, 32'h41dae551, 32'hc2966500, 32'hc25f9432, 32'hc2803763, 32'h424e6e7b, 32'h42586d7c};
test_weights[4000:4007] = '{32'h4245405c, 32'h429621b9, 32'hc291ed9b, 32'h41a10d6b, 32'hc29ddb94, 32'hc27c1985, 32'h426a3e11, 32'hc2223245};
test_bias[500:500] = '{32'h42626eec};
test_output[500:500] = '{32'h464dd69a};
test_input[4008:4015] = '{32'h42869116, 32'h420987c6, 32'h427974c6, 32'hc29b2e8d, 32'h4080d599, 32'hc2030c81, 32'h41dc37b4, 32'hc28b477f};
test_weights[4008:4015] = '{32'hc245ff1e, 32'hc2807ce0, 32'h42386067, 32'hc18b7ec6, 32'h42a87d55, 32'hc2875746, 32'hc2c0187d, 32'hc1998ca9};
test_bias[501:501] = '{32'hc28a3239};
test_output[501:501] = '{32'hc303f439};
test_input[4016:4023] = '{32'hc173f059, 32'hc281b6d6, 32'hc016424c, 32'hc18f4f4b, 32'h42857bf5, 32'hc2be134b, 32'hc2c71666, 32'h41ac1c35};
test_weights[4016:4023] = '{32'h424982b7, 32'h42a3f8e5, 32'hc285eef1, 32'hc2b5d3ec, 32'h412f92b2, 32'h42b68247, 32'hc16bf3ec, 32'hc28716ae};
test_bias[502:502] = '{32'h4229e00e};
test_output[502:502] = '{32'hc63e5a24};
test_input[4024:4031] = '{32'hc21b6a9b, 32'hc20789cc, 32'hc2017e50, 32'hc292280b, 32'hc2518d9f, 32'h4084caee, 32'h420e54f8, 32'h42a157a0};
test_weights[4024:4031] = '{32'h42b717ea, 32'h429b045f, 32'h4272f339, 32'h420d12dd, 32'hc2688a32, 32'h4255dde0, 32'hc27366a6, 32'hc23e9138};
test_bias[503:503] = '{32'h3f6471ac};
test_output[503:503] = '{32'hc6526c88};
test_input[4032:4039] = '{32'hc2c4ec80, 32'hc1a394ee, 32'h419e950e, 32'h41dcf02f, 32'h41ad95b2, 32'hc104849f, 32'hc2b3e73a, 32'h4246165a};
test_weights[4032:4039] = '{32'hc1c5f1a7, 32'hc28a9a57, 32'h4283f821, 32'h422eeadb, 32'hc2649b5e, 32'h424e0426, 32'hc1608dd9, 32'h426dcca4};
test_bias[504:504] = '{32'h42b501da};
test_output[504:504] = '{32'h460c9d52};
test_input[4040:4047] = '{32'h429ae77c, 32'h42a0a136, 32'h40a44697, 32'hc2b071e4, 32'hc28f2b9d, 32'hc2200173, 32'hc2929d10, 32'h42b8d515};
test_weights[4040:4047] = '{32'hc2065f9b, 32'hc2ba647e, 32'h41e597ba, 32'hc280facc, 32'hc225c1bc, 32'h4289aad6, 32'h4226b6ea, 32'h407a0a29};
test_bias[505:505] = '{32'hc2234a5b};
test_output[505:505] = '{32'hc5d3a1f2};
test_input[4048:4055] = '{32'h423ad981, 32'hc153cf19, 32'hc22adda4, 32'hc1c9896c, 32'hc1fe57af, 32'h424921e2, 32'h4234bfac, 32'hc23c4f07};
test_weights[4048:4055] = '{32'hc2c55bd7, 32'hc1938a1d, 32'hc2a5ab46, 32'hc14f9a0a, 32'h424ae39f, 32'h420d2c9d, 32'h42b8680c, 32'h4268300f};
test_bias[506:506] = '{32'hc2193251};
test_output[506:506] = '{32'h44842aeb};
test_input[4056:4063] = '{32'hc23deeea, 32'hc226d347, 32'hc21b7e29, 32'hc2c31352, 32'hbf3c80c1, 32'h4298fae9, 32'hc2671a42, 32'h4246ef50};
test_weights[4056:4063] = '{32'h424c9644, 32'hc1c922a5, 32'h4290d9da, 32'hc119ddd8, 32'hc2916dfd, 32'hc27b5b8c, 32'hc2be3c43, 32'h425e3d5e};
test_bias[507:507] = '{32'h41799173};
test_output[507:507] = '{32'h4383e332};
test_input[4064:4071] = '{32'h427cce98, 32'hc188fa2d, 32'hc18f4083, 32'h4135d736, 32'h411a7e31, 32'h41a7d17c, 32'h4242cc31, 32'h42a5a19e};
test_weights[4064:4071] = '{32'h40c136d5, 32'h42b7f818, 32'h40e0c324, 32'hc1eaa8ae, 32'hc190f1b1, 32'hbf167c97, 32'h42934c57, 32'hc2b8caf1};
test_bias[508:508] = '{32'h4248195f};
test_output[508:508] = '{32'hc5b6f79a};
test_input[4072:4079] = '{32'hc1ba7f74, 32'h428f4c0d, 32'h42ad3fe9, 32'hc2b7b1ad, 32'hc1becf77, 32'hc212b08f, 32'h42acca3f, 32'h41afe0f9};
test_weights[4072:4079] = '{32'hc21fba69, 32'h42bd5111, 32'h41cc29b9, 32'hc2587542, 32'hc1b63714, 32'h412bb908, 32'hc1bf82a9, 32'h4180d566};
test_bias[509:509] = '{32'h42a4f900};
test_output[509:509] = '{32'h46518ffe};
test_input[4080:4087] = '{32'h4204c1e2, 32'h409361e4, 32'h42a3d84d, 32'hc2608c28, 32'hc23de653, 32'hc2474181, 32'hc2305032, 32'h420d94c1};
test_weights[4080:4087] = '{32'h42a1a065, 32'hc280b366, 32'h425c735c, 32'h42399f60, 32'h42827003, 32'h42bd45ad, 32'h4271d26d, 32'h429f9e08};
test_bias[510:510] = '{32'h4219adf7};
test_output[510:510] = '{32'hc54f44e6};
test_input[4088:4095] = '{32'h417ae77e, 32'hc1cc0b80, 32'h4106a7d5, 32'h4282d011, 32'hc20ebbb4, 32'h42be325c, 32'hc1f4cc80, 32'h42c77eda};
test_weights[4088:4095] = '{32'hc1e9c541, 32'hc2215cd9, 32'hc1f102ab, 32'hc219a404, 32'h4259a666, 32'hc2c089da, 32'hc29de19b, 32'hc214abea};
test_bias[511:511] = '{32'hc2c1dbcc};
test_output[511:511] = '{32'hc6656247};
test_input[4096:4103] = '{32'hc28487a1, 32'hc20cfb03, 32'h4204340b, 32'hc1c63c07, 32'hc204a695, 32'hc24e266c, 32'h4174ed31, 32'hc1acd5f6};
test_weights[4096:4103] = '{32'h425d3aae, 32'h42906394, 32'hc1bfeede, 32'h42b250d7, 32'h426f1952, 32'h42a6892f, 32'h42ba3c0e, 32'hc29cb405};
test_bias[512:512] = '{32'hc2aaff44};
test_output[512:512] = '{32'hc64292bf};
test_input[4104:4111] = '{32'hc0a90ff0, 32'hc23f958d, 32'hc18b0eb3, 32'h429c4fe1, 32'h4214bf39, 32'hc24b36aa, 32'h40d55151, 32'h42b24721};
test_weights[4104:4111] = '{32'h427352e9, 32'hc2b3e6b7, 32'hc215a394, 32'hc29ed75f, 32'h426411a5, 32'h41946b2a, 32'h427d6cb2, 32'hc28a8a2a};
test_bias[513:513] = '{32'hc016bd78};
test_output[513:513] = '{32'hc5c01770};
test_input[4112:4119] = '{32'hc229d778, 32'hc1c3bec1, 32'h4286c747, 32'h42afd5bb, 32'hc192c0ab, 32'h4254d7f0, 32'hc2037006, 32'h42ba36e8};
test_weights[4112:4119] = '{32'h422f322b, 32'hc163753f, 32'h423a7e53, 32'hc1e7fc3b, 32'h4277f306, 32'h42b8c38c, 32'h426485b6, 32'hc2b16778};
test_bias[514:514] = '{32'hc28081e1};
test_output[514:514] = '{32'hc5e56903};
test_input[4120:4127] = '{32'hc2b8c7f9, 32'h407b7f2a, 32'h42982d53, 32'h42a63c7d, 32'hc2bf18ec, 32'h4041bc40, 32'hc293e2a8, 32'hc1f5ad2a};
test_weights[4120:4127] = '{32'h41acb6ce, 32'h42a2e39e, 32'h415c808c, 32'h4178006a, 32'hc22e73b3, 32'h42b7abd4, 32'h42b05070, 32'hc238de43};
test_bias[515:515] = '{32'hc2c6b768};
test_output[515:515] = '{32'hc2b63c9b};
test_input[4128:4135] = '{32'h42c6d040, 32'hc2690e5c, 32'hc2458afa, 32'hc2c3b0d8, 32'hbf0d80f1, 32'h42bff16c, 32'hc278901a, 32'hc29b118b};
test_weights[4128:4135] = '{32'hc28056c4, 32'hc2403fe6, 32'h425bb5a7, 32'hc22ffb9f, 32'h429e3cac, 32'h42b94ea7, 32'h429bae21, 32'hc296af7d};
test_bias[516:516] = '{32'hc280d6f0};
test_output[516:516] = '{32'h45f3d125};
test_input[4136:4143] = '{32'h422c38ac, 32'h42a539fa, 32'h42aa64ac, 32'h41e70af8, 32'h428d562d, 32'hc292faf6, 32'hc1385da3, 32'hc2c68f74};
test_weights[4136:4143] = '{32'hc24872b7, 32'hc0730be4, 32'h424618a3, 32'hc20de5a4, 32'h3ec7eb12, 32'hc1810c93, 32'h42ad437b, 32'h41fce88c};
test_bias[517:517] = '{32'hc176b312};
test_output[517:517] = '{32'hc50a7bd4};
test_input[4144:4151] = '{32'hc1c7957b, 32'hc2c18e42, 32'h420dab6f, 32'h42c7ff7d, 32'hc1d25104, 32'h40f5906e, 32'h42b87be9, 32'h42a5e59b};
test_weights[4144:4151] = '{32'hc1df6e87, 32'hc28ed761, 32'h4258a0a2, 32'h4248201f, 32'hbf90ccb6, 32'h42203bcc, 32'h41b1433b, 32'h42ac67ef};
test_bias[518:518] = '{32'hc265b52e};
test_output[518:518] = '{32'h46bb87cb};
test_input[4152:4159] = '{32'h42744e74, 32'hc2870b0a, 32'hc2969c88, 32'h421db23c, 32'hc1f814db, 32'h42b94f06, 32'h41bc83dd, 32'hc239c6a3};
test_weights[4152:4159] = '{32'hc2363f3b, 32'h421eb5fc, 32'hc26c1488, 32'h42879caf, 32'hc1dd6488, 32'hc0d95b4b, 32'hc2ad9179, 32'h42588235};
test_bias[519:519] = '{32'hc265108b};
test_output[519:519] = '{32'hc52ab735};
test_input[4160:4167] = '{32'hc25bb647, 32'hbe58d0d8, 32'h41dabb09, 32'hc29331cd, 32'hc2211846, 32'hbf550557, 32'h42a68222, 32'h42976de5};
test_weights[4160:4167] = '{32'hc29f125b, 32'h4244bfc3, 32'h424b1aa8, 32'hc233a081, 32'h4252f7d0, 32'hc286b934, 32'h41e4644f, 32'h426ff75e};
test_bias[520:520] = '{32'hc14da221};
test_output[520:520] = '{32'h46590719};
test_input[4168:4175] = '{32'hc26c1aeb, 32'h41dc55a8, 32'h4184c79d, 32'hc29d87f2, 32'hc2898969, 32'h4265cf07, 32'hc10da58a, 32'hc2ad4418};
test_weights[4168:4175] = '{32'h424070d4, 32'hc2b1ecf0, 32'hc2b36b24, 32'h4197e435, 32'hc28b11a3, 32'hc183f2a3, 32'h419a9925, 32'h41c34197};
test_bias[521:521] = '{32'hc1e33177};
test_output[521:521] = '{32'hc5d31111};
test_input[4176:4183] = '{32'hc2b4a476, 32'hc294c1e9, 32'hc11aaa9b, 32'hc2b328bf, 32'h4293bb4a, 32'h407fc618, 32'h429c480f, 32'h4227ff2c};
test_weights[4176:4183] = '{32'h42c254f5, 32'h428f06d7, 32'hc196b112, 32'hc198127a, 32'hc234bf4f, 32'hc1daf922, 32'h42089c12, 32'hc2185566};
test_bias[522:522] = '{32'hc10a6952};
test_output[522:522] = '{32'hc6641390};
test_input[4184:4191] = '{32'h42935f73, 32'hc19c6bdd, 32'hc287b82b, 32'hc1dcbfac, 32'h42c261b4, 32'hc29e1282, 32'hc29ddd41, 32'hc2971960};
test_weights[4184:4191] = '{32'hc19c20b5, 32'h428f865f, 32'h42297cac, 32'hc1f5ac24, 32'hc1dc6e4a, 32'hc2719e9b, 32'h42b9ae62, 32'hc29b1eef};
test_bias[523:523] = '{32'hc2b18081};
test_output[523:523] = '{32'hc5875179};
test_input[4192:4199] = '{32'hc0f159a0, 32'hc28cb030, 32'h4285daf9, 32'h41d40919, 32'h407b231d, 32'hc2893e45, 32'h42424b25, 32'h4295a0fa};
test_weights[4192:4199] = '{32'hc1bb6e81, 32'h3fe4906b, 32'hc18f0658, 32'h424116af, 32'h424112ed, 32'hc283d40f, 32'hc28d9e20, 32'h42b2ff74};
test_bias[524:524] = '{32'h4268f497};
test_output[524:524] = '{32'h45ff0931};
test_input[4200:4207] = '{32'h40e25096, 32'hc2b5f0e6, 32'h42700117, 32'h41da57ac, 32'h4207616f, 32'hc29ea729, 32'h4288da4c, 32'h4291ed96};
test_weights[4200:4207] = '{32'hc266008e, 32'h41331296, 32'h3ff737a8, 32'h42831a37, 32'hc1a92d42, 32'hc298a58f, 32'h42badadd, 32'hc1032420};
test_bias[525:525] = '{32'hc26d6b88};
test_output[525:525] = '{32'h4634899a};
test_input[4208:4215] = '{32'hc2b265b1, 32'hc28c5989, 32'h42818d9b, 32'h42abc771, 32'hc24e8ea5, 32'h4283675a, 32'hc02f07f9, 32'h42bab60d};
test_weights[4208:4215] = '{32'h41d152f9, 32'hc0521cd0, 32'h42b387ff, 32'hc1d4b1d7, 32'h41a97511, 32'h421165e4, 32'h41b1d815, 32'h40c17bc2};
test_bias[526:526] = '{32'h42993dfa};
test_output[526:526] = '{32'h454e6516};
test_input[4216:4223] = '{32'hc26daa77, 32'hc1f9f26d, 32'hc202a97e, 32'hc02403e5, 32'hc1af63e3, 32'hc25ba9ad, 32'h3e886786, 32'h41084f48};
test_weights[4216:4223] = '{32'hc24a713f, 32'h4214a4be, 32'h41eb8131, 32'h3fc5b3bc, 32'hc1cda00a, 32'hc21df5d7, 32'hc251fb80, 32'hc1e99dd1};
test_bias[527:527] = '{32'h42c5740e};
test_output[527:527] = '{32'h4557898a};
test_input[4224:4231] = '{32'h42936780, 32'hc2b3b12f, 32'hc24fb026, 32'hc287c9b8, 32'hc2b8eeb8, 32'hc2022855, 32'h4296f0cf, 32'hc2a23e4b};
test_weights[4224:4231] = '{32'h41a44cda, 32'h4294a7a0, 32'hc27cdc06, 32'hc2c5c5b8, 32'hbf2082e3, 32'h425d0141, 32'hc29d4227, 32'h40630a14};
test_bias[528:528] = '{32'hc1afa21f};
test_output[528:528] = '{32'hc54501d1};
test_input[4232:4239] = '{32'h4295c182, 32'hc2a4cfc4, 32'hc2a16fc7, 32'h415c298a, 32'hc2a52df8, 32'h42b64290, 32'hc264d261, 32'hc273f6af};
test_weights[4232:4239] = '{32'h41071c38, 32'h4249ceab, 32'hc217f480, 32'hc27d46a5, 32'hc2bc2c11, 32'h4244d854, 32'hc1b71d92, 32'h417f3b9e};
test_bias[529:529] = '{32'h42961779};
test_output[529:529] = '{32'h4631224b};
test_input[4240:4247] = '{32'h41b1486d, 32'h41dfa149, 32'hc22f28d3, 32'hc2b71ea0, 32'h42a9b98c, 32'h4185c281, 32'hc04928ef, 32'h429d711f};
test_weights[4240:4247] = '{32'hc2239400, 32'h4251b8ba, 32'h423026e1, 32'h42c38a46, 32'hc194a32a, 32'hc168a2f2, 32'hc28a2b07, 32'hc276abe5};
test_bias[530:530] = '{32'h41b00f24};
test_output[530:530] = '{32'hc682e820};
test_input[4248:4255] = '{32'hc280d6a9, 32'hc1f29b97, 32'h4193621b, 32'hc22d7240, 32'h429f0892, 32'h421e4c18, 32'h42ba6f18, 32'hc2388977};
test_weights[4248:4255] = '{32'hc28f4f12, 32'hc2806ffd, 32'h42812c89, 32'hc1b32d3a, 32'h41a262a2, 32'h42411a4c, 32'h42c6e790, 32'hc25d0e06};
test_bias[531:531] = '{32'h42ab01b1};
test_output[531:531] = '{32'h46bcb55f};
test_input[4256:4263] = '{32'h423243e0, 32'hc2afce15, 32'h42a2c35b, 32'hc28a40ac, 32'hc276ba0d, 32'h42778554, 32'hc27ee0a7, 32'hc26afc9a};
test_weights[4256:4263] = '{32'hc186a06d, 32'hc21de8df, 32'h4207e2f5, 32'hc14e7925, 32'h419d6b90, 32'h428c35df, 32'hc2bc4bf9, 32'h42391706};
test_bias[532:532] = '{32'h42ad5264};
test_output[532:532] = '{32'h464912a7};
test_input[4264:4271] = '{32'h4240e539, 32'h422fdc34, 32'h42a6df97, 32'h41849062, 32'hc2825045, 32'h427d0079, 32'h3fbe9ef7, 32'hc2b04af4};
test_weights[4264:4271] = '{32'hc20e0c91, 32'hc298cd34, 32'h3f62444d, 32'h424b1b62, 32'hc2b35271, 32'h41ecca27, 32'hc23cbc78, 32'h428db146};
test_bias[533:533] = '{32'h424974b7};
test_output[533:533] = '{32'hc5292f31};
test_input[4272:4279] = '{32'hc25daa7d, 32'h42bd63e1, 32'h42700652, 32'h42392e08, 32'hc1da9417, 32'hc0f12cad, 32'h41b393ca, 32'h4285df0a};
test_weights[4272:4279] = '{32'h4272dfc5, 32'hc2a7dfd3, 32'h42a02ef0, 32'h42c6b260, 32'hc1e288ab, 32'h41f33bd7, 32'h41a0a79d, 32'hc194fe53};
test_bias[534:534] = '{32'hc241eec4};
test_output[534:534] = '{32'hc509fb65};
test_input[4280:4287] = '{32'h41ea9224, 32'hc293fbdb, 32'h420bda89, 32'h41a66d33, 32'hc29b970e, 32'h42858410, 32'h409c670f, 32'h418ef607};
test_weights[4280:4287] = '{32'hc18424f1, 32'h42bc04ac, 32'h41e6e216, 32'h425912c5, 32'hc28f7a63, 32'h40d86cec, 32'h422151b2, 32'h42c4b15d};
test_bias[535:535] = '{32'h428e95cd};
test_output[535:535] = '{32'h452c416b};
test_input[4288:4295] = '{32'hc1c60c4e, 32'h4284a9c6, 32'h42bb9af1, 32'h42c77aa6, 32'h428722ba, 32'h3fa4dc3d, 32'h40df58fa, 32'hc19c4cd6};
test_weights[4288:4295] = '{32'h42302142, 32'hc174e5b3, 32'hc29318ff, 32'h419045e6, 32'h40d18efc, 32'hc26d11d1, 32'h40ffecf1, 32'h416e780b};
test_bias[536:536] = '{32'hc170dc97};
test_output[536:536] = '{32'hc5dd8fd7};
test_input[4296:4303] = '{32'h426fb8d8, 32'h4219a00a, 32'h42aed38e, 32'h4200bbf3, 32'h42122abc, 32'h420f192a, 32'h41996eba, 32'hc1e50256};
test_weights[4296:4303] = '{32'h4208863e, 32'h417230d6, 32'h423201a4, 32'h42130fa7, 32'hc28740b6, 32'h42183574, 32'hc23b556d, 32'h4207e539};
test_bias[537:537] = '{32'hc2b1348e};
test_output[537:537] = '{32'h4590b6e8};
test_input[4304:4311] = '{32'h42b2bcc4, 32'hc2b7d0b5, 32'hc243d2b8, 32'hc205260b, 32'hc1f2cca4, 32'h41616d06, 32'hc11d2f1a, 32'h42ac11bb};
test_weights[4304:4311] = '{32'hc29d8d92, 32'hc180c995, 32'h3fc418ed, 32'hc25f468a, 32'h409338ca, 32'hc2b06b33, 32'hc28a29b5, 32'h41d3f8e0};
test_bias[538:538] = '{32'h42577349};
test_output[538:538] = '{32'hc5063d18};
test_input[4312:4319] = '{32'h42966cfa, 32'h4151a5bd, 32'h42a2f853, 32'h42548ef4, 32'hc1f7813d, 32'h4212c9cf, 32'hc29aeba9, 32'hc280ae79};
test_weights[4312:4319] = '{32'hc2295fb9, 32'hc2149427, 32'hc200687b, 32'h41f6d9b3, 32'hc26d68ad, 32'h428ca6f9, 32'hc1535b23, 32'hc18fe75e};
test_bias[539:539] = '{32'h41e2e165};
test_output[539:539] = '{32'h44f74acb};
test_input[4320:4327] = '{32'h42ae0744, 32'h4226fe7c, 32'hc222a1b4, 32'hc1403056, 32'h42c5e2a7, 32'h428640c2, 32'hc2c476ed, 32'h429941f5};
test_weights[4320:4327] = '{32'h42bc935f, 32'hc0afa678, 32'hc2845cfc, 32'h41e09777, 32'hc15d0e50, 32'hc2bc81b9, 32'hc2188b8d, 32'h428a3cfe};
test_bias[540:540] = '{32'hc09eb82a};
test_output[540:540] = '{32'h463662c2};
test_input[4328:4335] = '{32'h42823aff, 32'h42393e62, 32'h415dd15e, 32'h42ad5ee8, 32'hc1daec46, 32'hc265775a, 32'hc28b239e, 32'h42c2b28e};
test_weights[4328:4335] = '{32'h419cba7e, 32'h424e620e, 32'h421e573a, 32'hc298f543, 32'h41ad6ffa, 32'hc29721b4, 32'hc2a673b5, 32'hc288fb2d};
test_bias[541:541] = '{32'h42294ab5};
test_output[541:541] = '{32'h43f56a46};
test_input[4336:4343] = '{32'hc293bcea, 32'hc20688b9, 32'hc2328865, 32'h4200bc02, 32'hc2a28a01, 32'hc2ac8121, 32'h426dc832, 32'h422f63de};
test_weights[4336:4343] = '{32'hc224e882, 32'h42bf9b6a, 32'h420db252, 32'hc1fed5f3, 32'hc1d76221, 32'h42a69573, 32'hc263eb09, 32'hc2190eeb};
test_bias[542:542] = '{32'hc2ac640c};
test_output[542:542] = '{32'hc64a097a};
test_input[4344:4351] = '{32'hc1bc5d86, 32'hc292b686, 32'h428af79d, 32'hbefa83dd, 32'hc25a28bb, 32'h4245ce4d, 32'hc23ef721, 32'h403285ee};
test_weights[4344:4351] = '{32'hc299627f, 32'hc2b686ef, 32'h4270941e, 32'hc138270d, 32'h42c66e99, 32'hbfd6655a, 32'hc279cb6a, 32'hc1abb4d9};
test_bias[543:543] = '{32'hc2b3ab0a};
test_output[543:543] = '{32'h461c9b7f};
test_input[4352:4359] = '{32'hc2b572ca, 32'h4283f561, 32'hc2c5eecc, 32'h3fd2a28e, 32'h429e8d35, 32'hc149d5b9, 32'h42aa3ca4, 32'h41bdb8dd};
test_weights[4352:4359] = '{32'hc229d6b4, 32'hc24602ec, 32'h42b831ad, 32'hc1c0a53b, 32'hc0d01c2c, 32'h429f0ed7, 32'hc28b03d5, 32'h41912214};
test_bias[544:544] = '{32'hc2b419d8};
test_output[544:544] = '{32'hc674bca6};
test_input[4360:4367] = '{32'hc2106e1b, 32'hc02e8638, 32'h426dea91, 32'h4227fc58, 32'hc290f4d8, 32'h4280b645, 32'h420b073f, 32'h42bb862f};
test_weights[4360:4367] = '{32'hc17e1526, 32'hc27845d0, 32'hc2949a46, 32'h41c98b1d, 32'h42beefea, 32'hc2591052, 32'hc2384949, 32'h42532ff6};
test_bias[545:545] = '{32'hc1c00c29};
test_output[545:545] = '{32'hc617a5ad};
test_input[4368:4375] = '{32'h41b3100d, 32'hc26f7f37, 32'hc1e2e4b8, 32'h42c69063, 32'hc286c2c2, 32'h426227bd, 32'h42a86d74, 32'h42053698};
test_weights[4368:4375] = '{32'hc113f7c5, 32'h4220de23, 32'hc2b941d5, 32'h42973ca9, 32'hc18d7abd, 32'hc2b1a002, 32'hbfc4a813, 32'hc19240ab};
test_bias[546:546] = '{32'h4286d131};
test_output[546:546] = '{32'h453cb271};
test_input[4376:4383] = '{32'hc0e7d702, 32'h429d9840, 32'h418a21a0, 32'hc2c2e6d9, 32'h4285b912, 32'h42561bff, 32'h42113d68, 32'hc2178f30};
test_weights[4376:4383] = '{32'hc1d90484, 32'h41eda752, 32'hc2613905, 32'hc250d3b1, 32'h42c59e0f, 32'hc1b3a398, 32'hc22ccd43, 32'hc08cba07};
test_bias[547:547] = '{32'h42c55a5a};
test_output[547:547] = '{32'h462807ee};
test_input[4384:4391] = '{32'h41296ae8, 32'hc2a4c2a6, 32'h3fb10735, 32'hc2c0f4dc, 32'hc25dc7ce, 32'hc27a57b0, 32'hc284b0b7, 32'hc209b8ba};
test_weights[4384:4391] = '{32'hc2751ad1, 32'hc213aace, 32'h4228be80, 32'h42a1f8d5, 32'h426e18fe, 32'hc2a0f35d, 32'hc0d27e8c, 32'h42a1fd15};
test_bias[548:548] = '{32'hc299eb0e};
test_output[548:548] = '{32'hc5bd3cde};
test_input[4392:4399] = '{32'hc2c06c14, 32'h423c731c, 32'hc15da057, 32'h41ca5029, 32'h42249aea, 32'h42210cb3, 32'hc286d45e, 32'h428ca418};
test_weights[4392:4399] = '{32'h424eeb63, 32'h4260824e, 32'h41cb9064, 32'hc2bc8f07, 32'hc2a2766a, 32'hc1476b52, 32'hc2b8ab28, 32'h42a5c43f};
test_bias[549:549] = '{32'hc26286fb};
test_output[549:549] = '{32'h4540a773};
test_input[4400:4407] = '{32'hc2ade202, 32'hc20c2876, 32'h424ff3d8, 32'hc2a8bc46, 32'hc23a20ed, 32'hc0a3677b, 32'hc24eb3db, 32'hc231a61c};
test_weights[4400:4407] = '{32'hc240ad6c, 32'hc2423fba, 32'h401cbcb0, 32'hc28f6230, 32'h41cf391e, 32'h421931c5, 32'h421662e9, 32'h427007b3};
test_bias[550:550] = '{32'h41edc20b};
test_output[550:550] = '{32'h45be31ee};
test_input[4408:4415] = '{32'h41d8e51c, 32'h42c4c20f, 32'h42c182a8, 32'h4270baa0, 32'h425e7daa, 32'hc1a024c0, 32'h42a4ca0d, 32'h407861ac};
test_weights[4408:4415] = '{32'hc29bd0a4, 32'hc2c3714c, 32'h415539a0, 32'h41890408, 32'h42a82382, 32'hc2a98d66, 32'h4278a332, 32'h429d8848};
test_bias[551:551] = '{32'hc209460c};
test_output[551:551] = '{32'h45138640};
test_input[4416:4423] = '{32'h3fd5437e, 32'hc199b30a, 32'hc2a81140, 32'h419567da, 32'h4258de14, 32'hc1d066e7, 32'h4286d48c, 32'hc2abe179};
test_weights[4416:4423] = '{32'hc218e272, 32'hc2605734, 32'h421b6580, 32'hc1ba17aa, 32'h429004b9, 32'h41f77f07, 32'h420d7025, 32'hc208b71f};
test_bias[552:552] = '{32'hc1bca4c8};
test_output[552:552] = '{32'h45b2741f};
test_input[4424:4431] = '{32'hc28640ea, 32'h427c723a, 32'hc1ce8ea7, 32'hc188f8ef, 32'hc29c4c02, 32'h4120b8e5, 32'h4261c670, 32'hc24c5632};
test_weights[4424:4431] = '{32'h429d93bb, 32'h4182729e, 32'h4145e950, 32'h4235437f, 32'h426f964f, 32'hc29500d0, 32'hc1167426, 32'h4293faf9};
test_bias[553:553] = '{32'h42c4d5f3};
test_output[553:553] = '{32'hc66a5115};
test_input[4432:4439] = '{32'hc271de22, 32'hc13fbfc0, 32'hc19f5772, 32'h422e4ecc, 32'hc22d4c92, 32'h411fdbfe, 32'hc23b1e5d, 32'h4249fd2b};
test_weights[4432:4439] = '{32'h428e5b9f, 32'hc021c4e5, 32'hc10b8c39, 32'h4292caf0, 32'h423e4f76, 32'hc0a75ce5, 32'hc0deb2df, 32'hc2976f74};
test_bias[554:554] = '{32'h425c80fd};
test_output[554:554] = '{32'hc5c9cfc2};
test_input[4440:4447] = '{32'hc2991521, 32'h424570d3, 32'hc2b79718, 32'h4240f040, 32'h420d5744, 32'hc1fcf28c, 32'hc281b63f, 32'hc1e47e49};
test_weights[4440:4447] = '{32'hc2c64a96, 32'h418f6bca, 32'h42a5c89b, 32'hc2884ce7, 32'hc201b0af, 32'hc2c3cd30, 32'h42344488, 32'hc2bedfb4};
test_bias[555:555] = '{32'h42a420a5};
test_output[555:555] = '{32'hc412f0a8};
test_input[4448:4455] = '{32'hc1c1debf, 32'hc296b9a1, 32'hc198c3e6, 32'hc24a71b9, 32'h420198a2, 32'hc24c0878, 32'hc26b2ccb, 32'h42c2a843};
test_weights[4448:4455] = '{32'h4123c290, 32'h408398ea, 32'h427a323d, 32'hc21948e9, 32'hc2316932, 32'h42793066, 32'hbf95afcd, 32'hc2074cb0};
test_bias[556:556] = '{32'h429159a1};
test_output[556:556] = '{32'hc5ecd20d};
test_input[4456:4463] = '{32'h4003024f, 32'h429d9a2d, 32'hc29f9826, 32'hbffab201, 32'h427a79e5, 32'hc2a0b934, 32'hc25a674a, 32'hc29ee015};
test_weights[4456:4463] = '{32'h4298638b, 32'h428e40ae, 32'h42a39933, 32'hc1d9a718, 32'hc20289d5, 32'hc0974e74, 32'h411de4ca, 32'hc256c916};
test_bias[557:557] = '{32'hc28dbf08};
test_output[557:557] = '{32'h449fdfdd};
test_input[4464:4471] = '{32'hc1becd53, 32'h42c17e66, 32'h4214fedf, 32'h42ac429d, 32'h42bcc2db, 32'h426e40c9, 32'hc21c7f93, 32'h41f7c8f7};
test_weights[4464:4471] = '{32'hc1e88ed9, 32'hc25a8b2b, 32'h42b917cd, 32'h41e5bd12, 32'h427b6abb, 32'hc2151613, 32'hc2539d5a, 32'h427781b1};
test_bias[558:558] = '{32'h4295b85b};
test_output[558:558] = '{32'h460e363c};
test_input[4472:4479] = '{32'h42baca9f, 32'h41459098, 32'hc21bf75d, 32'hc246a906, 32'h429898a2, 32'hc2b471f0, 32'h421b7315, 32'h425b6b93};
test_weights[4472:4479] = '{32'h4171c324, 32'h429431fa, 32'hc255b6cd, 32'h41a3c217, 32'h41585c9a, 32'hc1c6662d, 32'h4257ba51, 32'hc27344b0};
test_bias[559:559] = '{32'hc24c86b7};
test_output[559:559] = '{32'h45a7d5c6};
test_input[4480:4487] = '{32'hc11c01c3, 32'hc22d2f2d, 32'h42b341f3, 32'hc2514b5a, 32'h428b2415, 32'h42b03b70, 32'hc171a47b, 32'hc281b76b};
test_weights[4480:4487] = '{32'h4260b3ac, 32'h41b43f23, 32'h41a5b5cd, 32'hc2acb33f, 32'h42bcb1c5, 32'hc230f98b, 32'h4244596a, 32'hc15c8b11};
test_bias[560:560] = '{32'hc21ef1d7};
test_output[560:560] = '{32'h45ee6ca7};
test_input[4488:4495] = '{32'hc194b2a5, 32'h429921d6, 32'hc2b0a955, 32'hc2afcc86, 32'h42b465a2, 32'h42145468, 32'hc25f0d2b, 32'hc1c065df};
test_weights[4488:4495] = '{32'hc2208955, 32'hc1fe1810, 32'hc0cea8bb, 32'hc1c94d42, 32'hc2088898, 32'hc286c6f9, 32'h408a9e0c, 32'h42b79ab4};
test_bias[561:561] = '{32'hc285271e};
test_output[561:561] = '{32'hc5daaa85};
test_input[4496:4503] = '{32'h423e7874, 32'h41a49ed2, 32'h42b78fb1, 32'hc1b86480, 32'hc207d8c0, 32'hc25f8707, 32'hc2aadd33, 32'hc2adb592};
test_weights[4496:4503] = '{32'hc1da4de7, 32'hc2274ce1, 32'h42b155d1, 32'h41ac4e58, 32'h426d95d1, 32'hc2a16e13, 32'hc21c5a98, 32'h4193edfa};
test_bias[562:562] = '{32'hc266fcc9};
test_output[562:562] = '{32'h4616c99f};
test_input[4504:4511] = '{32'hc2c464c1, 32'h421067d1, 32'h42a147d1, 32'h40cce212, 32'hc2454c46, 32'h423074c7, 32'hc29e655c, 32'h4293bee2};
test_weights[4504:4511] = '{32'h424beeab, 32'h41363864, 32'h423efbf5, 32'hc280d47e, 32'hc20cfe9a, 32'h4277239d, 32'h41de134f, 32'hc241428b};
test_bias[563:563] = '{32'hc1035bf2};
test_output[563:563] = '{32'hc51a50f9};
test_input[4512:4519] = '{32'hc142845e, 32'h42a5027f, 32'h41fbd9a2, 32'h42aa414f, 32'h4283baaf, 32'hc2be6212, 32'hc07de465, 32'h41aaa769};
test_weights[4512:4519] = '{32'hc2610219, 32'h41f163bf, 32'hc26903dc, 32'hc2a3936b, 32'h42992e2d, 32'hc2593f79, 32'h4161c789, 32'hc2772abb};
test_bias[564:564] = '{32'hc2ba6acd};
test_output[564:564] = '{32'h454345aa};
test_input[4520:4527] = '{32'h42c10c44, 32'hc18774da, 32'h421c994b, 32'hc21ddf19, 32'hc22d80da, 32'hc239b40a, 32'hc2b0afbd, 32'h40495d0e};
test_weights[4520:4527] = '{32'hc236c16a, 32'hc1b28cb1, 32'h41800164, 32'hc28dcc5e, 32'hc16003ef, 32'hc2ab2abc, 32'h42652667, 32'h42b060de};
test_bias[565:565] = '{32'h429209bb};
test_output[565:565] = '{32'hc4385980};
test_input[4528:4535] = '{32'h42b84241, 32'hc1b8ee52, 32'h419c879e, 32'hc22bb83e, 32'hc214ac4b, 32'hc2926e9e, 32'h419a8713, 32'h415d6989};
test_weights[4528:4535] = '{32'hc088658b, 32'hc0af9b0e, 32'h41e3ebd5, 32'h424322a4, 32'hc20d30d8, 32'hbf058018, 32'h4079b74e, 32'hc1e76594};
test_bias[566:566] = '{32'hc273f3a3};
test_output[566:566] = '{32'hc4519b88};
test_input[4536:4543] = '{32'h4205138e, 32'hc28322a9, 32'hc241f614, 32'hc2b887d8, 32'hc2a2c08e, 32'h42c3679b, 32'hc237e46e, 32'h42abf4f2};
test_weights[4536:4543] = '{32'hc0aab712, 32'h42abb422, 32'h428a1652, 32'h40ed0017, 32'hc2829dd8, 32'hc10e0e62, 32'hc1c6de31, 32'h42b090d9};
test_bias[567:567] = '{32'h42b5172c};
test_output[567:567] = '{32'h45568fe6};
test_input[4544:4551] = '{32'hc2469cc3, 32'hc2c1c0ef, 32'h429ea2b5, 32'h42b19eb9, 32'h410734f5, 32'hc28cac96, 32'hc2b9a56a, 32'hc28c6171};
test_weights[4544:4551] = '{32'hc1f672e5, 32'hc17b6a88, 32'hc2add808, 32'hc2b5c76d, 32'h4257487f, 32'hc28fcab0, 32'hc2a221da, 32'h40dc9565};
test_bias[568:568] = '{32'h427aea93};
test_output[568:568] = '{32'h442f3f72};
test_input[4552:4559] = '{32'hc1804fe1, 32'hc2210bb2, 32'hbeeeed67, 32'hc290c441, 32'hc29f1104, 32'h4232166c, 32'h42a2ed7c, 32'h40aae90f};
test_weights[4552:4559] = '{32'hc296d5cf, 32'h429e1d73, 32'h42567287, 32'hc235b925, 32'hc29ab8c0, 32'hc2bf456e, 32'h42b6de09, 32'hc28a27b9};
test_bias[569:569] = '{32'hc04d2a44};
test_output[569:569] = '{32'h4620555c};
test_input[4560:4567] = '{32'hc2bb58c6, 32'hc26099cc, 32'hc278bb4a, 32'h42a1e638, 32'hc2189b3c, 32'hc28e98c2, 32'h422587c5, 32'h42a40a87};
test_weights[4560:4567] = '{32'h410f5a5f, 32'h427e16b6, 32'hc2bc9e10, 32'hc2293cad, 32'h429d5fbb, 32'h424f7f23, 32'h428f3e19, 32'hc285e42b};
test_bias[570:570] = '{32'hc2bb7ad2};
test_output[570:570] = '{32'hc6305fc8};
test_input[4568:4575] = '{32'h41985ea1, 32'hc1138116, 32'h41a26ecf, 32'hc28fd69a, 32'h42a5bac6, 32'hc2a44a19, 32'hc19d3f32, 32'h415462c7};
test_weights[4568:4575] = '{32'hc275c04f, 32'h42b1749d, 32'hc1c94aec, 32'h41d80eb9, 32'hc295fa3b, 32'h42aa668d, 32'h41d604ec, 32'h429c7ab8};
test_bias[571:571] = '{32'h424859a5};
test_output[571:571] = '{32'hc6858675};
test_input[4576:4583] = '{32'h425bf215, 32'hc16e5a51, 32'h42b55de5, 32'h42a5c53a, 32'hc26fe6ed, 32'h42bc0415, 32'hc26c5a77, 32'hc231d0c6};
test_weights[4576:4583] = '{32'h42716ea3, 32'h42931c5f, 32'h423529aa, 32'hc23d45d3, 32'h420d8d1b, 32'hc0879797, 32'hc20c10e3, 32'h4277fc45};
test_bias[572:572] = '{32'hc2c3d2c7};
test_output[572:572] = '{32'hc4605400};
test_input[4584:4591] = '{32'hc2c791e1, 32'hc24d6416, 32'h426f975a, 32'hc25d6a0f, 32'hc2ba4ba5, 32'hc2877d57, 32'hc2be5c44, 32'hc268db34};
test_weights[4584:4591] = '{32'hc1a5e107, 32'h428d136a, 32'h42b7a2ba, 32'hc241ba5b, 32'hc251d2a1, 32'hc2c26b3e, 32'h4225839e, 32'h418585f2};
test_bias[573:573] = '{32'hc2385173};
test_output[573:573] = '{32'h464d5c59};
test_input[4592:4599] = '{32'h42c54e53, 32'hc286e0a9, 32'hc2b7d836, 32'h41078549, 32'hc2a8c447, 32'h4291e58d, 32'h41f11379, 32'h41491fdc};
test_weights[4592:4599] = '{32'h424f9f9c, 32'h41f5fc82, 32'h42b340bf, 32'h4259dca6, 32'hbfd53b84, 32'h428a4887, 32'h412f0c4e, 32'hc12f58b1};
test_bias[574:574] = '{32'hc1de638b};
test_output[574:574] = '{32'h441a8aad};
test_input[4600:4607] = '{32'hc1f63b7c, 32'hc2a0aa0e, 32'hc2a53515, 32'h42009723, 32'hc15e9749, 32'hc28bfe10, 32'hc267ff4c, 32'hc1ee4fa4};
test_weights[4600:4607] = '{32'hc28fe3eb, 32'hc0c2108b, 32'h41fb7d12, 32'h413d8b8e, 32'hc1e14a46, 32'h42a0f402, 32'h42c7b9d7, 32'hc2708ec6};
test_bias[575:575] = '{32'h42882c7f};
test_output[575:575] = '{32'hc607c006};
test_input[4608:4615] = '{32'h421a4dc1, 32'hbfcdae77, 32'hc2630920, 32'h421ea87e, 32'h422bac9b, 32'hc2c63276, 32'hc18ed94a, 32'h427dfe58};
test_weights[4608:4615] = '{32'hc2c56aea, 32'hc245c740, 32'h4271b44d, 32'hc2817a10, 32'h415b0597, 32'hc0db01f9, 32'h427e4aaa, 32'hc2b11a80};
test_bias[576:576] = '{32'h422a0e2b};
test_output[576:576] = '{32'hc66d1eb6};
test_input[4616:4623] = '{32'h423de0da, 32'hc2a95fbd, 32'hc12bfe25, 32'h42b344e2, 32'hc0b4769b, 32'hc200dbe6, 32'hc287a383, 32'h421df469};
test_weights[4616:4623] = '{32'hc1d0548d, 32'hc222370b, 32'h41b4b5f0, 32'h420ef65e, 32'h41917037, 32'h423c6139, 32'h42a2a93b, 32'h41b338db};
test_bias[577:577] = '{32'h429df157};
test_output[577:577] = '{32'hc47d36c1};
test_input[4624:4631] = '{32'h42c4894e, 32'h429b6ac9, 32'hc2c731ef, 32'h3fd7d46a, 32'hc28fc24e, 32'h42b0d526, 32'hc1d5bc21, 32'h3ffba796};
test_weights[4624:4631] = '{32'h429b33e7, 32'h422c15f4, 32'h422dc386, 32'hc2a66339, 32'h424e3cca, 32'h3f7f2639, 32'hc2a1e150, 32'h419d0038};
test_bias[578:578] = '{32'h426feb25};
test_output[578:578] = '{32'h45a0c8a2};
test_input[4632:4639] = '{32'h41acb5d6, 32'h41da8dca, 32'hc2515464, 32'h4231e8e5, 32'h417e28ca, 32'hbf89ad9c, 32'hc2012fed, 32'hc278e3e6};
test_weights[4632:4639] = '{32'hc2840f0d, 32'h4280714c, 32'h4274cb80, 32'hc207af59, 32'hc11ded1f, 32'hc233d68c, 32'h42c5f55d, 32'hc25bdea2};
test_bias[579:579] = '{32'hc199c22e};
test_output[579:579] = '{32'hc585f49c};
test_input[4640:4647] = '{32'hc1e7826c, 32'h414719d2, 32'h429bf4d9, 32'hc2034aec, 32'h426b6b30, 32'hc210ad6b, 32'hc2010208, 32'h40c94ea0};
test_weights[4640:4647] = '{32'h42bbc2a5, 32'h401cdeaa, 32'h418320dc, 32'hc2c61140, 32'hc256fb8f, 32'h42602637, 32'h41071237, 32'hc272dba9};
test_bias[580:580] = '{32'h41e5b43e};
test_output[580:580] = '{32'hc57850b0};
test_input[4648:4655] = '{32'h40fdcbbc, 32'h42a89037, 32'h42076ef3, 32'hc1254661, 32'h41a69892, 32'hc26a8ff0, 32'h40bf8b77, 32'h42c7f7ef};
test_weights[4648:4655] = '{32'h400de4d6, 32'h42131745, 32'hc2b64498, 32'hc1aff579, 32'h426bdb0b, 32'h3fd86697, 32'h428efba3, 32'h42489538};
test_bias[581:581] = '{32'hc1f9b37b};
test_output[581:581] = '{32'h45d46d48};
test_input[4656:4663] = '{32'h40febaae, 32'hc297ae1b, 32'h42a81817, 32'hc2b6f07f, 32'hc10e489e, 32'h42be4c79, 32'hc27ca6e8, 32'hc26d2ae9};
test_weights[4656:4663] = '{32'h426da13b, 32'hc17b89d5, 32'hc0be4ac7, 32'hc2b22637, 32'h42209b33, 32'hc2b2db94, 32'hc2b3442c, 32'hc2478431};
test_bias[582:582] = '{32'h429777b4};
test_output[582:582] = '{32'h460ed620};
test_input[4664:4671] = '{32'hc1aaed04, 32'hc29ca0b5, 32'h4299bb68, 32'h40f77ab3, 32'h4205ff70, 32'hc2828d9d, 32'h42ae1bca, 32'hc2c42970};
test_weights[4664:4671] = '{32'h422d40e3, 32'hc1416577, 32'h42ba7304, 32'hc29d0f69, 32'h41e85be3, 32'hc2308793, 32'hc21be240, 32'h419cfe10};
test_bias[583:583] = '{32'h42860d6f};
test_output[583:583] = '{32'h45a1f931};
test_input[4672:4679] = '{32'h41b63313, 32'hc2823af0, 32'h428887e5, 32'hc1d73ac4, 32'hc28e1f39, 32'h408dd2d1, 32'hc2766ff6, 32'hc231bb84};
test_weights[4672:4679] = '{32'hc20db2ab, 32'h428e514a, 32'hc1db39ac, 32'hc1ec7e6b, 32'hc29d289e, 32'hc253ae8a, 32'hc275c057, 32'h40ce188d};
test_bias[584:584] = '{32'hc2867021};
test_output[584:584] = '{32'h450d9775};
test_input[4680:4687] = '{32'hc2982ef7, 32'h423aab56, 32'h42465512, 32'hc1a6c6d3, 32'hc23cddd0, 32'hc27671cf, 32'hc2543b6a, 32'h42883d63};
test_weights[4680:4687] = '{32'hc205f82b, 32'h42b53974, 32'h42c5ac68, 32'hc27f157f, 32'hc2b6b0be, 32'hc27d3bd8, 32'h42b9019d, 32'hc21627bd};
test_bias[585:585] = '{32'h3ff71ce9};
test_output[585:585] = '{32'h4656f5d8};
test_input[4688:4695] = '{32'hc27b6ad0, 32'hc0f7287d, 32'h42822b2e, 32'hc003b0c8, 32'hc1b17fbe, 32'hc26f6df7, 32'hc2b7e122, 32'hc295349e};
test_weights[4688:4695] = '{32'hc1544fcd, 32'h4298be03, 32'hc21b942a, 32'h42a3b631, 32'hc20f437b, 32'h423f8109, 32'h41b30e79, 32'h4224061e};
test_bias[586:586] = '{32'hc0d8f547};
test_output[586:586] = '{32'hc616ca02};
test_input[4696:4703] = '{32'h3ef1e713, 32'hc2c02cdd, 32'hc23f129a, 32'h42a3f6d7, 32'hc1de7844, 32'hc2929206, 32'h41aee975, 32'h420253c7};
test_weights[4696:4703] = '{32'h40c434f5, 32'hc22044e8, 32'h401ccbc1, 32'h428c53be, 32'hc22df4df, 32'h4268a759, 32'hbf3ff430, 32'h4225d3bf};
test_bias[587:587] = '{32'h42384176};
test_output[587:587] = '{32'h45f43a16};
test_input[4704:4711] = '{32'h41ef6da0, 32'hc13b7d47, 32'h42711f9d, 32'h41895124, 32'hc2a1471b, 32'hc27445bc, 32'hc2a8c392, 32'h423a1663};
test_weights[4704:4711] = '{32'h422750e1, 32'hc199c8c1, 32'hc28eadfa, 32'hc1abbb9e, 32'h40f2271e, 32'hc24f8d18, 32'hc162d93d, 32'hc2025e40};
test_bias[588:588] = '{32'hc2acff98};
test_output[588:588] = '{32'hc481f4e7};
test_input[4712:4719] = '{32'h4160fe34, 32'hc202caad, 32'hc28f507e, 32'hc2ad5399, 32'hc1928d28, 32'hc2c0a73f, 32'hc24cb6f3, 32'hc29a3569};
test_weights[4712:4719] = '{32'hc2939197, 32'h428a049b, 32'hc288aa7d, 32'h4295146d, 32'h428e06c9, 32'hc1aedd50, 32'h41bde67f, 32'h42335f56};
test_bias[589:589] = '{32'h42c1b003};
test_output[589:589] = '{32'hc606d140};
test_input[4720:4727] = '{32'hc1c47054, 32'hc1fc9c16, 32'hc2273927, 32'h418795b0, 32'h418eadef, 32'h427b7063, 32'hc2381985, 32'h412ce2fe};
test_weights[4720:4727] = '{32'h429b55b9, 32'h421aa7e4, 32'hc28739b7, 32'h42a38b92, 32'h42415fcf, 32'hc2bc880a, 32'h42af4121, 32'hc2af14ae};
test_bias[590:590] = '{32'h42650a69};
test_output[590:590] = '{32'hc60b11eb};
test_input[4728:4735] = '{32'hc2b836fb, 32'h411279ff, 32'h41db4db4, 32'h4287ae07, 32'hc2ba61a9, 32'hc2a08721, 32'h42567ef8, 32'hc27af281};
test_weights[4728:4735] = '{32'h41bd2867, 32'h410461fb, 32'h3f84d26b, 32'hc0fba1ba, 32'hc264d256, 32'h422b7fed, 32'h4204b97d, 32'hc2a78b39};
test_bias[591:591] = '{32'h41febf8d};
test_output[591:591] = '{32'h45c66a88};
test_input[4736:4743] = '{32'hc1a07dcb, 32'hc1acab62, 32'hc1552e80, 32'h41f1e091, 32'h4275d3e0, 32'hc28d568b, 32'hc261e107, 32'hc21f4a7c};
test_weights[4736:4743] = '{32'hc27d2a9d, 32'hc085be46, 32'hc28153f5, 32'h42a86365, 32'h42911a3c, 32'h425c01ba, 32'hc1df162d, 32'hc2c536a0};
test_bias[592:592] = '{32'h41cb89b4};
test_output[592:592] = '{32'h4629c782};
test_input[4744:4751] = '{32'hc157b112, 32'hc1f57cdc, 32'hc2909ab3, 32'hc2b48c4b, 32'h429c5c06, 32'hc2853d91, 32'h42476dba, 32'hc1296bc7};
test_weights[4744:4751] = '{32'h4211527e, 32'h41df2c4d, 32'h42a7e1bc, 32'h3eeb54cf, 32'hc2ba08e1, 32'h42547964, 32'hc2a0cea7, 32'h428c5750};
test_bias[593:593] = '{32'h41273397};
test_output[593:593] = '{32'hc6b3c103};
test_input[4752:4759] = '{32'h42ac0ab4, 32'hc226d89b, 32'hc293c7c2, 32'h420b2a5e, 32'hc127ca31, 32'h42241fb3, 32'h41086b68, 32'h4112256c};
test_weights[4752:4759] = '{32'h42c1475f, 32'h4215c2fc, 32'hc2401ffc, 32'h4285da5a, 32'h427237bf, 32'h427fccc5, 32'hc186af20, 32'h42127df2};
test_bias[594:594] = '{32'hc175f498};
test_output[594:594] = '{32'h46672544};
test_input[4760:4767] = '{32'hc2a67c32, 32'hc2244564, 32'hc262c9cc, 32'hc1562beb, 32'hc2965bbc, 32'hc22c611c, 32'hc1c63253, 32'h41dcf684};
test_weights[4760:4767] = '{32'h41df3914, 32'h4185fd6c, 32'hc2c4c681, 32'hc21ba9eb, 32'h42551cf9, 32'hc25bbbd0, 32'hc2aaf4f5, 32'h42a9dd36};
test_bias[595:595] = '{32'hbf11df9d};
test_output[595:595] = '{32'h45b8cc9e};
test_input[4768:4775] = '{32'hc1dce88d, 32'h40bc71a6, 32'hc29058c3, 32'h3fa0811e, 32'hc2800a45, 32'hc2b6016c, 32'hc1a648fa, 32'hc1ce6ab9};
test_weights[4768:4775] = '{32'hc29edbed, 32'hc1000fe8, 32'h4286f8c8, 32'h4279cb56, 32'h423a7a89, 32'h404f0905, 32'hc2586cb1, 32'hc29cb142};
test_bias[596:596] = '{32'h420af218};
test_output[596:596] = '{32'hc52b84bc};
test_input[4776:4783] = '{32'h42a60cf7, 32'hc28f7491, 32'hc1660a46, 32'h41a8a18a, 32'h41836b2a, 32'h420ec88b, 32'h42c764b7, 32'h40dc3656};
test_weights[4776:4783] = '{32'h41d5c413, 32'h427761df, 32'hc251cca7, 32'hc1f6a0a1, 32'hc2aab56a, 32'hc2a2e3e9, 32'h42876c99, 32'h4166ef9b};
test_bias[597:597] = '{32'hc1dd7899};
test_output[597:597] = '{32'h43c7d2fe};
test_input[4784:4791] = '{32'h422bf6a1, 32'h4216e649, 32'h412d9ccf, 32'hc0adc484, 32'h4201b764, 32'h422b481d, 32'hc133107a, 32'h4201122b};
test_weights[4784:4791] = '{32'hc27ae63d, 32'hc2a04046, 32'hc2a5fe70, 32'hc2ad3f6f, 32'hc2b58571, 32'hc2812718, 32'h42a2f3b3, 32'h4275630f};
test_bias[598:598] = '{32'h4229a199};
test_output[598:598] = '{32'hc627ef97};
test_input[4792:4799] = '{32'h4296a101, 32'h418e4bed, 32'h42974436, 32'h41901500, 32'hc288b4a8, 32'hc28308bf, 32'h42b91075, 32'hc257e163};
test_weights[4792:4799] = '{32'hc20b541a, 32'h4276c644, 32'h3fa3a1aa, 32'hc0a68026, 32'hc2462e3f, 32'hc2bfd38b, 32'hc29fbf89, 32'h426cf460};
test_bias[599:599] = '{32'hc18a04eb};
test_output[599:599] = '{32'hc5199d27};
test_input[4800:4807] = '{32'hc1bc9cb3, 32'hc2ac9105, 32'hc2981d36, 32'hc160a01b, 32'h428b9b3e, 32'h424ff896, 32'hc2b1b60f, 32'h42b79d9e};
test_weights[4800:4807] = '{32'h42aef036, 32'hc2947895, 32'hc2b8a6f7, 32'h426c4795, 32'h429d6862, 32'hc28d4116, 32'hc2b71169, 32'h42adcdcd};
test_bias[600:600] = '{32'hc2bd022e};
test_output[600:600] = '{32'h46ddad30};
test_input[4808:4815] = '{32'h4209cf4d, 32'h424ad363, 32'hc2c6e914, 32'hc245e032, 32'hc2a0a4a0, 32'h4292369f, 32'hc26de561, 32'hc098aa50};
test_weights[4808:4815] = '{32'h42aff023, 32'hc24c0ea2, 32'hc24d5d5b, 32'h429bc220, 32'h42c53844, 32'hc2c596c2, 32'h42722556, 32'h411d4299};
test_bias[601:601] = '{32'h42625e5d};
test_output[601:601] = '{32'hc6851844};
test_input[4816:4823] = '{32'h40e01450, 32'hc2928e17, 32'hc147aaa1, 32'hc2a17956, 32'hc282548e, 32'h423a6f32, 32'h42b7a945, 32'h400a06c7};
test_weights[4816:4823] = '{32'h411ebdb9, 32'hc25b9fe0, 32'hc287e595, 32'hc1954235, 32'hc226c7f6, 32'h42839eb4, 32'h42ba378b, 32'h42c1e453};
test_bias[602:602] = '{32'hc0122cfd};
test_output[602:602] = '{32'h46a3f90e};
test_input[4824:4831] = '{32'hc288a4d5, 32'h41eac864, 32'h42c4ba06, 32'h413e11f7, 32'hc223b346, 32'hc241199e, 32'h4193877d, 32'hc2b4b8af};
test_weights[4824:4831] = '{32'h4193e824, 32'hc21ff8cd, 32'h41b9bdc6, 32'h4285403c, 32'hc2c41165, 32'hc2012218, 32'h4298ce6a, 32'h422a26d7};
test_bias[603:603] = '{32'h422129e2};
test_output[603:603] = '{32'h456e6637};
test_input[4832:4839] = '{32'hc2ad5253, 32'hc19f434f, 32'h408a936f, 32'h41ed2a22, 32'h429077eb, 32'h4225f5b7, 32'hc21c2a5a, 32'hc29fec24};
test_weights[4832:4839] = '{32'h416e2b2d, 32'hc21f0763, 32'hc2c5aaed, 32'h4236d582, 32'h4293cc5c, 32'h41afe386, 32'h42c49931, 32'hc1334e45};
test_bias[604:604] = '{32'hc263a1ef};
test_output[604:604] = '{32'h456603e5};
test_input[4840:4847] = '{32'hc2a1ba71, 32'hc2c7a772, 32'hc08a3d8c, 32'h428ca805, 32'h42567f68, 32'h4109ea08, 32'hc2aa620e, 32'h4215288c};
test_weights[4840:4847] = '{32'hc2946c4b, 32'h429b37c0, 32'hc2bb7094, 32'hc153e72e, 32'hc2b818ac, 32'h41f89ac8, 32'h4292ee56, 32'hc2b69c05};
test_bias[605:605] = '{32'h425417e4};
test_output[605:605] = '{32'hc6814eef};
test_input[4848:4855] = '{32'h41a7a156, 32'hc21342ac, 32'h4212642d, 32'hc20afbe8, 32'h42627e62, 32'hc026dfa1, 32'h427dffbf, 32'h3fb420e9};
test_weights[4848:4855] = '{32'hc28ad700, 32'hc246e86d, 32'h4036d324, 32'h42c0c47d, 32'h4127ba15, 32'hc1edb844, 32'hc24aeb7a, 32'hc0f7d842};
test_bias[606:606] = '{32'h42a5b247};
test_output[606:606] = '{32'hc5a71523};
test_input[4856:4863] = '{32'hc2a6617f, 32'h41f47e09, 32'h424dbf32, 32'h4241a428, 32'hc28cc92f, 32'h418e0f49, 32'h42a9bc0e, 32'h4291b288};
test_weights[4856:4863] = '{32'h42baca94, 32'hc208a44a, 32'hc29a9f35, 32'hc1d7fc5d, 32'h418f561a, 32'h4181c600, 32'hc1e5a18b, 32'h42020808};
test_bias[607:607] = '{32'h41ad1072};
test_output[607:607] = '{32'hc66c3295};
test_input[4864:4871] = '{32'h424cf0ac, 32'hc2213750, 32'h42ad098b, 32'h408bf628, 32'h412c799b, 32'hc2373f0f, 32'h40b25353, 32'hc2a4c15c};
test_weights[4864:4871] = '{32'h42b087bd, 32'hc2662aba, 32'hc2c138ee, 32'h429a4e2a, 32'hc27ee612, 32'hc2886634, 32'hc2a9101f, 32'h424e5118};
test_bias[608:608] = '{32'hc291df17};
test_output[608:608] = '{32'hc55cf5d8};
test_input[4872:4879] = '{32'h40c8e93f, 32'hc2197442, 32'hc26a88bb, 32'hc28abc5a, 32'hc16ea1f5, 32'h416ea2ff, 32'hc1f0b80a, 32'hc28b571c};
test_weights[4872:4879] = '{32'hc2631964, 32'hc1c4281b, 32'h4267c523, 32'h425d52eb, 32'h415dda3d, 32'h418f034f, 32'hc253ad69, 32'h41c24fae};
test_bias[609:609] = '{32'hc26d92e7};
test_output[609:609] = '{32'hc5d2f67f};
test_input[4880:4887] = '{32'h4100b7b0, 32'h40dc692f, 32'hc1a465bc, 32'h42568843, 32'hc2a6e25b, 32'h42548199, 32'h428950b7, 32'h41b629c7};
test_weights[4880:4887] = '{32'h41906778, 32'hc29e7601, 32'hc1f66c93, 32'h417ce65a, 32'hc27abd91, 32'hc2c65515, 32'h422b7086, 32'hc1ab3a92};
test_bias[610:610] = '{32'h41aa1c66};
test_output[610:610] = '{32'h455befd9};
test_input[4888:4895] = '{32'h40af3481, 32'hc28f3d1b, 32'hc12897e2, 32'hc29e968b, 32'h404a0887, 32'hbfa4efac, 32'h3f47b90d, 32'hc29d1228};
test_weights[4888:4895] = '{32'h41f5c63c, 32'h41691e26, 32'h4263d00a, 32'hc21c532e, 32'h4296d0fc, 32'h423b220c, 32'h4251fd85, 32'hc1d907d0};
test_bias[611:611] = '{32'h42c1349b};
test_output[611:611] = '{32'h457e5685};
test_input[4896:4903] = '{32'h411aa6c4, 32'hc1b802f4, 32'h4190f4c8, 32'h42a5ee69, 32'h42568024, 32'h419e6fa2, 32'hc23083b7, 32'h421662c6};
test_weights[4896:4903] = '{32'hc221a5aa, 32'h42aaca92, 32'hc20b8769, 32'h41aa3f5a, 32'h427af9c0, 32'h414ef4c5, 32'h42490c51, 32'h415f36fe};
test_bias[612:612] = '{32'h41c6e975};
test_output[612:612] = '{32'h4436b96b};
test_input[4904:4911] = '{32'hc2794258, 32'h4292b808, 32'h42789047, 32'h41ebc842, 32'hc2a62b9c, 32'h42b0d50c, 32'hc2b6f3d2, 32'hc21f3ad6};
test_weights[4904:4911] = '{32'hc25028ba, 32'hc297ee3d, 32'h4237aa61, 32'hc2c42cb9, 32'hc297b8b2, 32'h42965376, 32'h42085939, 32'h428b06f4};
test_bias[613:613] = '{32'hc2c34cf5};
test_output[613:613] = '{32'h458fb00b};
test_input[4912:4919] = '{32'hc2155d63, 32'h4288679f, 32'hc25213a6, 32'h42a165a6, 32'hbf05596a, 32'h42689dff, 32'h4261b468, 32'h42a4831c};
test_weights[4912:4919] = '{32'h42298ae2, 32'hc2b19ce9, 32'hc22062e7, 32'hc259ccd8, 32'hc2acf88c, 32'h41e7c642, 32'hc27185c1, 32'hc205a79a};
test_bias[614:614] = '{32'hbdffc8a1};
test_output[614:614] = '{32'hc6604607};
test_input[4920:4927] = '{32'hc2a29c7d, 32'hc260a371, 32'h42a9fb23, 32'hc1dceb5f, 32'h429f4bb5, 32'hc1a7d7a2, 32'h42980063, 32'h426cd279};
test_weights[4920:4927] = '{32'hc2c5960d, 32'hc1dea566, 32'hc263ac80, 32'hc20ebf69, 32'hc2a69e98, 32'h41b40dc2, 32'hc19f6d30, 32'hc2112805};
test_bias[615:615] = '{32'hc2c21e6a};
test_output[615:615] = '{32'hc5a0235d};
test_input[4928:4935] = '{32'h41ee4cc0, 32'hc2940a92, 32'h42acf6ec, 32'hc2698d33, 32'hc1d4a58f, 32'h41e3b456, 32'h41ab1380, 32'h42aa6798};
test_weights[4928:4935] = '{32'h42ab0ff3, 32'h4290f1b5, 32'h41277f42, 32'h42a48420, 32'h41d7769f, 32'h3f893e3b, 32'hc2a30e21, 32'h42631ce5};
test_bias[616:616] = '{32'hc2a56300};
test_output[616:616] = '{32'hc589208c};
test_input[4936:4943] = '{32'hc1549b87, 32'h428692d8, 32'h421349ef, 32'h42a981d1, 32'hc25f0164, 32'h3fe09829, 32'hc1304804, 32'h4120335e};
test_weights[4936:4943] = '{32'h4188f24e, 32'h42b6b3fd, 32'hc206829b, 32'hc1b26652, 32'hc119f4d1, 32'h41ccc371, 32'hc143ebc2, 32'hc20e71ed};
test_bias[617:617] = '{32'hc237317a};
test_output[617:617] = '{32'h45420f6c};
test_input[4944:4951] = '{32'hc22f7d33, 32'h420cb36e, 32'hc236dea1, 32'h42991b63, 32'hc2180071, 32'h4290ec2f, 32'hc1f554bb, 32'h42310bfb};
test_weights[4944:4951] = '{32'hc2a3343c, 32'hbf23e651, 32'h421c6e99, 32'h4266feeb, 32'h423f0d23, 32'h4291303b, 32'hc2ac3123, 32'h425a1015};
test_bias[618:618] = '{32'h4270296d};
test_output[618:618] = '{32'h46667416};
test_input[4952:4959] = '{32'h40ed07dc, 32'h425f9687, 32'h426d5be2, 32'hc2b09fe2, 32'h410445a2, 32'h412a779a, 32'h421c8f13, 32'hc26ee728};
test_weights[4952:4959] = '{32'h42847ebb, 32'h4280382a, 32'hc2896e0f, 32'hc23e15ba, 32'h42c5fa1e, 32'h42987d60, 32'hc1f4160e, 32'h429a3255};
test_bias[619:619] = '{32'h40468e1d};
test_output[619:619] = '{32'h41e21608};
test_input[4960:4967] = '{32'hc2551e40, 32'hc2764044, 32'h424c9f49, 32'hc21c75a2, 32'h4224119b, 32'hc2819f2b, 32'h416a3b7d, 32'hc2b6286e};
test_weights[4960:4967] = '{32'hc085d5a1, 32'hc22605ad, 32'hc2914138, 32'h412f0b0d, 32'h4219481a, 32'hc0a68de0, 32'h427bc1e4, 32'hc2b1e65d};
test_bias[620:620] = '{32'h41a82c02};
test_output[620:620] = '{32'h4615cf4d};
test_input[4968:4975] = '{32'h3f87d4ba, 32'h4291a6c0, 32'hc21c604c, 32'hc29d2dda, 32'hc0a0acef, 32'h422eba64, 32'h41ae4a99, 32'h42acfbc8};
test_weights[4968:4975] = '{32'hc0471d4d, 32'hc2c76f0c, 32'h42999713, 32'hc23d3bec, 32'hc2b7bd56, 32'h41ffc1fa, 32'h4295b718, 32'hc22d6a1d};
test_bias[621:621] = '{32'h428b0dbe};
test_output[621:621] = '{32'hc5d2a87e};
test_input[4976:4983] = '{32'hc0a43018, 32'h40b1a887, 32'h4221d0ea, 32'hc23183af, 32'hc1d80639, 32'hc1c5d9c5, 32'hc275c8b4, 32'h42aa0c47};
test_weights[4976:4983] = '{32'h42209591, 32'h42b2d4c9, 32'h425e9ed9, 32'hc2c127e6, 32'h4251a65c, 32'h42aafda5, 32'hc10c3713, 32'hc120cf5e};
test_bias[622:622] = '{32'hc1a89060};
test_output[622:622] = '{32'h453910e0};
test_input[4984:4991] = '{32'h424c45c4, 32'hc2a911b4, 32'h4160a0ff, 32'hc2574975, 32'hc21392ff, 32'hc29fd82c, 32'hc180aeb4, 32'h42a9be55};
test_weights[4984:4991] = '{32'hc1c47058, 32'h42bd8560, 32'h42119f30, 32'h422df262, 32'hc2995c01, 32'hc1f6af2a, 32'hc28a0463, 32'hc21bddac};
test_bias[623:623] = '{32'hc0e804f1};
test_output[623:623] = '{32'hc5fa270d};
test_input[4992:4999] = '{32'h42b4d01f, 32'hc1c3e138, 32'h427be147, 32'h42874d17, 32'hc2942279, 32'hc172a070, 32'hc2b741b5, 32'h42922e63};
test_weights[4992:4999] = '{32'h4289c78c, 32'hc2c2112b, 32'h424fb780, 32'hc2bfe1e6, 32'hc258eafe, 32'h40e0ce89, 32'h426c776d, 32'hc293f623};
test_bias[624:624] = '{32'hc1ad42af};
test_output[624:624] = '{32'hc4c20540};
test_input[5000:5007] = '{32'hc1d61571, 32'h4259cac8, 32'h420c7081, 32'h42a195cb, 32'h426cf61a, 32'h42739684, 32'h42c11fac, 32'hc23b802a};
test_weights[5000:5007] = '{32'h4289ac15, 32'hc242c0b6, 32'h42b19a12, 32'hc2407e1c, 32'hc2b57afc, 32'h427411a0, 32'h3f562fbf, 32'hc20a9ab1};
test_bias[625:625] = '{32'hc28176f9};
test_output[625:625] = '{32'hc5a51534};
test_input[5008:5015] = '{32'h429e6397, 32'h428e8bad, 32'hc2af8011, 32'hc22263cf, 32'hc0999e0d, 32'h4265a04e, 32'h42968c99, 32'hc21e649f};
test_weights[5008:5015] = '{32'hc082e9e6, 32'h428c0089, 32'hc25581bd, 32'hc2afbf90, 32'h3f2493f5, 32'h3fd03dcc, 32'h42996f1a, 32'h3febfbc9};
test_bias[626:626] = '{32'hc2ad230f};
test_output[626:626] = '{32'h46917c14};
test_input[5016:5023] = '{32'h420f2827, 32'h41b962c3, 32'h4295b7b8, 32'hc10da2c1, 32'h41a06d4e, 32'h4200b473, 32'h42ac74cd, 32'hc23f3d57};
test_weights[5016:5023] = '{32'hc25fda45, 32'h4268c034, 32'hc22a0b23, 32'h426bbaa2, 32'hc288bea6, 32'hc2c1ae94, 32'hc2438c48, 32'hc2c4a708};
test_bias[627:627] = '{32'h429aa722};
test_output[627:627] = '{32'hc6016ac2};
test_input[5024:5031] = '{32'hc20b7463, 32'h4186f008, 32'hc21ee738, 32'h42c35c1f, 32'hc2bf6a4b, 32'hc2839007, 32'h41f2cf94, 32'hc28973e0};
test_weights[5024:5031] = '{32'h4280cdf3, 32'hc299d6be, 32'h407cc16f, 32'hc1731e07, 32'hc20ac435, 32'h4270d8c6, 32'h41d9c9a9, 32'h420e9b5e};
test_bias[628:628] = '{32'hc29c9dd2};
test_output[628:628] = '{32'hc5eb3517};
test_input[5032:5039] = '{32'hc292757a, 32'hc180a53c, 32'h418e8727, 32'hc245def4, 32'hc25ce6ef, 32'h4261c8d4, 32'h429457bb, 32'h422c5f2c};
test_weights[5032:5039] = '{32'hc1880e4d, 32'hc1c48238, 32'h42244d9f, 32'h3fc456ea, 32'hc23bb773, 32'hc2bd06ce, 32'hc298c137, 32'h42aa196a};
test_bias[629:629] = '{32'hc2930381};
test_output[629:629] = '{32'hc51d85cf};
test_input[5040:5047] = '{32'h4145b8e0, 32'h41f660ab, 32'hc21f2de0, 32'hc279cba0, 32'h429e701c, 32'hc1a26904, 32'hc26840ed, 32'hc272d25c};
test_weights[5040:5047] = '{32'h424a4475, 32'hc226e93c, 32'hc2c6482c, 32'hc290b995, 32'hc01f2ee9, 32'hc222ce70, 32'hc0158799, 32'h41b94a0b};
test_bias[630:630] = '{32'hc1f898ab};
test_output[630:630] = '{32'h45dedef7};
test_input[5048:5055] = '{32'hc15dc5fa, 32'hc2bc4625, 32'hc10d4dfc, 32'hc1f58e6e, 32'hbfa2e6c6, 32'hc290e80b, 32'hc2189907, 32'hc290d2e5};
test_weights[5048:5055] = '{32'hc1617971, 32'h42af3a7e, 32'h4183c3d4, 32'hc12746dd, 32'hc29d090f, 32'hc24ba28c, 32'hc28e10a3, 32'h41a9b3f6};
test_bias[631:631] = '{32'h424d369f};
test_output[631:631] = '{32'hc532f738};
test_input[5056:5063] = '{32'h42bac61b, 32'h4233f402, 32'h4112ba4c, 32'hc14ee844, 32'h428dc33d, 32'hc2b2c630, 32'hc2492d83, 32'hc2b379b6};
test_weights[5056:5063] = '{32'hc2986fc7, 32'hc1fb2628, 32'h4292f5d5, 32'hc2b276e3, 32'h41357e49, 32'h42c42aa7, 32'h428800f1, 32'hc284c0ee};
test_bias[632:632] = '{32'h42270312};
test_output[632:632] = '{32'hc63cde4d};
test_input[5064:5071] = '{32'h42489683, 32'h427af991, 32'hc2a23a2f, 32'hc277b94f, 32'hc19fef3f, 32'h4194e41d, 32'hc249b216, 32'hc206d80e};
test_weights[5064:5071] = '{32'hc2ba651f, 32'h41d41de1, 32'hbfa08f7e, 32'h4216e2ba, 32'h419d73ea, 32'h4282220d, 32'hc267693d, 32'h42ac3e0a};
test_bias[633:633] = '{32'hc25a9e3e};
test_output[633:633] = '{32'hc58b9c54};
test_input[5072:5079] = '{32'h427c67c5, 32'hc20901f6, 32'h426bf238, 32'hc1b11eab, 32'h4255d011, 32'h41d473fb, 32'h4085a249, 32'h42167a3e};
test_weights[5072:5079] = '{32'hc20e8fd7, 32'hc206f019, 32'hc281c09f, 32'hc04c1601, 32'hc24fe845, 32'hc1790267, 32'h423a860b, 32'h426b04ac};
test_bias[634:634] = '{32'hc1a8fb25};
test_output[634:634] = '{32'hc5b0cb63};
test_input[5080:5087] = '{32'h4212d50b, 32'h42883192, 32'hc249a9f4, 32'hc2bfc83c, 32'h42437798, 32'h422b351f, 32'h4272fc9a, 32'h4216258e};
test_weights[5080:5087] = '{32'hc1bec1c5, 32'hc20dd5c7, 32'hc21d267f, 32'hc0b5fb36, 32'h42a8cf02, 32'hc29e28f7, 32'hc2332353, 32'hc27585c5};
test_bias[635:635] = '{32'hc211832c};
test_output[635:635] = '{32'hc59ee7ea};
test_input[5088:5095] = '{32'h42aa2d00, 32'hc2c6f9f3, 32'h418fa224, 32'h42b29642, 32'hc102aeae, 32'h42bdb0ea, 32'hc283f226, 32'hc2932d70};
test_weights[5088:5095] = '{32'hc203d18a, 32'hc299f74c, 32'hc2941049, 32'hc26322ca, 32'h42573950, 32'h420234a4, 32'h426d6a73, 32'hc25e7c8f};
test_bias[636:636] = '{32'h41e124fe};
test_output[636:636] = '{32'h44a3949a};
test_input[5096:5103] = '{32'hbe09b826, 32'hc285e4a8, 32'h4298ccd9, 32'h41bbc89e, 32'h427da155, 32'h42b2ab60, 32'h42b8fcc3, 32'h42b5c6d4};
test_weights[5096:5103] = '{32'hc2b1b38b, 32'h42658aec, 32'hc1ed3742, 32'h426b31f3, 32'hc1ab7e2a, 32'hc1162a8c, 32'h4130c305, 32'h42b28887};
test_bias[637:637] = '{32'h4122fb4b};
test_output[637:637] = '{32'h450b893c};
test_input[5104:5111] = '{32'hc24f9b47, 32'hc290c6ff, 32'h41470c0a, 32'h4283d9cd, 32'hc1b642db, 32'h4238dfdf, 32'h3f3f0a14, 32'hc196160b};
test_weights[5104:5111] = '{32'h42069298, 32'h4264d994, 32'h414b9122, 32'h40e71703, 32'hc25dc60e, 32'hc207183e, 32'h42c3aa84, 32'h4263cedb};
test_bias[638:638] = '{32'hc2b7b84f};
test_output[638:638] = '{32'hc5cf7395};
test_input[5112:5119] = '{32'h42b5c25e, 32'hc2a87769, 32'h3ff00c84, 32'h42bcfc48, 32'hc292e7d4, 32'hc287f7e0, 32'hc1d8dfb8, 32'hc1fe92a0};
test_weights[5112:5119] = '{32'h425df77f, 32'hc203fcb9, 32'hc2bb7c07, 32'h4238ea0b, 32'h41f7b1b3, 32'h4117fc87, 32'hc28b8823, 32'hc0905cd7};
test_bias[639:639] = '{32'hc085fa1a};
test_output[639:639] = '{32'h462dd66a};
test_input[5120:5127] = '{32'hc17b7cab, 32'h421c16ef, 32'hc2597a71, 32'h42aea7ca, 32'hc1c088e4, 32'hc244412b, 32'h421a3799, 32'hc21290e3};
test_weights[5120:5127] = '{32'hc1f9cb17, 32'h428d434c, 32'h4240f60f, 32'h41ca01c3, 32'hc293ded6, 32'h4232cfd6, 32'h4228faa8, 32'h425a24e7};
test_bias[640:640] = '{32'hc216b46f};
test_output[640:640] = '{32'h44fb0480};
test_input[5128:5135] = '{32'h429e5efc, 32'hc147a2b0, 32'h428e516b, 32'h4151d10c, 32'h4298ee09, 32'h42a7e4b1, 32'h4257f61c, 32'hc177c539};
test_weights[5128:5135] = '{32'h428f89f5, 32'hc0af8164, 32'h42982959, 32'h42a022e6, 32'hc25e3b0d, 32'h41c925a7, 32'h42a52d2e, 32'h42bbc547};
test_bias[641:641] = '{32'h428902c3};
test_output[641:641] = '{32'h464d7db9};
test_input[5136:5143] = '{32'hc2bc9124, 32'h420651be, 32'h42191d4c, 32'h4196bfeb, 32'hc169fb8e, 32'hbf0123f5, 32'h425f73c0, 32'hc288588e};
test_weights[5136:5143] = '{32'hc2a7bdb7, 32'hc234b9f8, 32'h41a6a5e7, 32'hc008d30d, 32'hc1aa4627, 32'hc293e28b, 32'hc25ba92a, 32'hc2764c18};
test_bias[642:642] = '{32'h41b76ad6};
test_output[642:642] = '{32'h460723e3};
test_input[5144:5151] = '{32'hc00d12c1, 32'h4279d9a9, 32'h4239bca8, 32'hc228c89a, 32'hc2181b1e, 32'h42bced16, 32'h42b288b1, 32'hc2163196};
test_weights[5144:5151] = '{32'h4293dd31, 32'hc277417c, 32'h4283ca4a, 32'h42293adb, 32'h4294b048, 32'hc1fb88e8, 32'hc2677fe5, 32'h4052ebd6};
test_bias[643:643] = '{32'hc2c3c7e5};
test_output[643:643] = '{32'hc659ba25};
test_input[5152:5159] = '{32'hc2864b3f, 32'hc281b2e9, 32'hc21f04fc, 32'h423f30b0, 32'hc25f5bc7, 32'hc231bac0, 32'h428587d3, 32'hc21ad3b5};
test_weights[5152:5159] = '{32'h40c7babc, 32'h4103e888, 32'h420b497e, 32'h4272894a, 32'h41d0ff51, 32'h41b69f79, 32'hc0aff337, 32'h429bbaa9};
test_bias[644:644] = '{32'h42558f61};
test_output[644:644] = '{32'hc5a3c4cb};
test_input[5160:5167] = '{32'h428047e9, 32'hc1b41d2c, 32'hc21fba88, 32'hc210d70b, 32'hbe24ea66, 32'h42b30359, 32'h4222ce89, 32'h423dd909};
test_weights[5160:5167] = '{32'h4012c967, 32'hc200d29e, 32'h42b730d5, 32'h426d5859, 32'hc2326235, 32'hc20586cf, 32'h4267593e, 32'hc26faf36};
test_bias[645:645] = '{32'hc20a5e7f};
test_output[645:645] = '{32'hc603dca5};
test_input[5168:5175] = '{32'h42c7df94, 32'hc1580ce5, 32'h42299155, 32'h42a01e4b, 32'hc194e382, 32'h4209ef9a, 32'h4294a938, 32'h421b21c4};
test_weights[5168:5175] = '{32'h427101e9, 32'hc2717ccf, 32'h42b656a7, 32'hc2303009, 32'hc293c7e7, 32'hc2b737d3, 32'hc0819529, 32'hc2aab9bb};
test_bias[646:646] = '{32'h419718ce};
test_output[646:646] = '{32'h44e0cef0};
test_input[5176:5183] = '{32'hc0a8dc75, 32'h4127ffbe, 32'hc2882657, 32'h4248352b, 32'h42a30cfd, 32'h42c3b773, 32'hc1751c27, 32'h421b2127};
test_weights[5176:5183] = '{32'h425313a1, 32'hc28ca518, 32'hc25426b3, 32'h42423b9c, 32'h41ecd440, 32'hc18afdef, 32'h4223c850, 32'hc2ac1a66};
test_bias[647:647] = '{32'hc2c1675d};
test_output[647:647] = '{32'h44d184a7};
test_input[5184:5191] = '{32'hc0519800, 32'hc203277d, 32'h4226533a, 32'hc24fd275, 32'h41b29c6b, 32'h41a9c6be, 32'h4173b418, 32'h422e80cb};
test_weights[5184:5191] = '{32'h41c5521e, 32'hc226d3db, 32'hc23f667a, 32'h428b3140, 32'h420c36e2, 32'h42bac255, 32'h3fdabaa4, 32'hc29e2d88};
test_bias[648:648] = '{32'hc2ac3269};
test_output[648:648] = '{32'hc59e4738};
test_input[5192:5199] = '{32'h42b5b688, 32'hc284b2ac, 32'h429cca16, 32'hc2c4201a, 32'h4218d9d0, 32'h425060d1, 32'hc0c0539d, 32'h4208f22f};
test_weights[5192:5199] = '{32'hc2c45ec7, 32'h41ac78e8, 32'hc23d72b6, 32'h42bdc22c, 32'h42982411, 32'h42555557, 32'hc278551e, 32'hc21c43c7};
test_bias[649:649] = '{32'hc2045d95};
test_output[649:649] = '{32'hc691f0e0};
test_input[5200:5207] = '{32'hc2769891, 32'hc22e8c86, 32'h4167dd86, 32'hc1eab2cc, 32'hc2b0c778, 32'hc1c34c0f, 32'hc298ffed, 32'h428067a0};
test_weights[5200:5207] = '{32'h41ca3889, 32'h42842aec, 32'hc238a778, 32'h42b685ab, 32'h42acc482, 32'h421e4cf2, 32'h42c0e99a, 32'hc2579b45};
test_bias[650:650] = '{32'h4297b387};
test_output[650:650] = '{32'hc6d4232c};
test_input[5208:5215] = '{32'hc2bb8d49, 32'hc24485cd, 32'h42555bbe, 32'h42a61000, 32'hc2b4526a, 32'hc1d6e29f, 32'h42c541e2, 32'hc2a94118};
test_weights[5208:5215] = '{32'h42900dfc, 32'hc27e6713, 32'hc222f8bd, 32'h42abe9dc, 32'h40ad2fec, 32'hc244734d, 32'hc230748a, 32'h41356d90};
test_bias[651:651] = '{32'h42469b0d};
test_output[651:651] = '{32'hc5417683};
test_input[5216:5223] = '{32'h4211d4b6, 32'h42a44bc1, 32'h4211e91e, 32'hc2482143, 32'h4218e141, 32'h41d29dfb, 32'hc1c11270, 32'h4297a8be};
test_weights[5216:5223] = '{32'h429ef2f9, 32'hc25d8d3c, 32'h42b1ed1a, 32'hc2454eab, 32'h4221c31d, 32'h42bfe1d1, 32'hc29ee511, 32'hc1cd0024};
test_bias[652:652] = '{32'hc0cddeed};
test_output[652:652] = '{32'h45fd1eee};
test_input[5224:5231] = '{32'h41ddc845, 32'hc1a05f74, 32'hc2837c49, 32'hc242439e, 32'h426c2cfd, 32'h426c2c01, 32'h427e7ac4, 32'h419ad408};
test_weights[5224:5231] = '{32'h42794d37, 32'hc2a935ad, 32'hc1dda295, 32'h411d1ee7, 32'hc2638037, 32'hc2734a64, 32'h42b57a51, 32'hc1028ea2};
test_bias[653:653] = '{32'h424ec423};
test_output[653:653] = '{32'h4559d992};
test_input[5232:5239] = '{32'h4214adec, 32'hc2ae6aa1, 32'h4204b8c6, 32'hc112a2a9, 32'hc257b7d5, 32'hc28acb6b, 32'h428677a3, 32'hc065d72b};
test_weights[5232:5239] = '{32'h425caf7f, 32'hc2956524, 32'h417a375b, 32'h41399f7d, 32'h42bbae98, 32'hc24e3b84, 32'hc24843dd, 32'hc1563b8c};
test_bias[654:654] = '{32'hc25a830a};
test_output[654:654] = '{32'h4580d049};
test_input[5240:5247] = '{32'h400e9270, 32'hc123c8f3, 32'hc2b71922, 32'h41d1cf77, 32'h429f64a0, 32'h42174ffe, 32'h41a3ddb1, 32'h4200daec};
test_weights[5240:5247] = '{32'hc1d2db72, 32'hc1d7e0ba, 32'hc27938ac, 32'hc21b9b8b, 32'hc24582e8, 32'hc2c43c92, 32'hc2bc1367, 32'hc2b745cf};
test_bias[655:655] = '{32'h41799e87};
test_output[655:655] = '{32'hc5edc158};
test_input[5248:5255] = '{32'h42331c76, 32'hc261ed36, 32'h42bf4adb, 32'hc2ad8908, 32'h4235030e, 32'hc2862f47, 32'h428b9e75, 32'h428d104b};
test_weights[5248:5255] = '{32'hc1d52770, 32'hc206e327, 32'hc22d2409, 32'h42998765, 32'hc2c651f4, 32'hc1186d8b, 32'h427a3b05, 32'h42233bdf};
test_bias[656:656] = '{32'hc2bc9742};
test_output[656:656] = '{32'hc5d41121};
test_input[5256:5263] = '{32'h420e8e8c, 32'h4285f6df, 32'hc22a93a9, 32'h425bb43d, 32'h428a6abc, 32'h4270cfc0, 32'h42c3dc4f, 32'h42a16d70};
test_weights[5256:5263] = '{32'hc2006655, 32'hc041a38c, 32'h42b21255, 32'h41b69c0a, 32'h4276ecd1, 32'h41a24b05, 32'hc21aa3b3, 32'hc24ad94c};
test_bias[657:657] = '{32'hc12e1d63};
test_output[657:657] = '{32'hc5c47161};
test_input[5264:5271] = '{32'hc11785bd, 32'hc28db4e0, 32'hc2b0ba59, 32'hc18fd90f, 32'hc2acebf5, 32'hc2c67e56, 32'h3fec8b51, 32'h41c8c721};
test_weights[5264:5271] = '{32'h4275dc74, 32'h425cbd2b, 32'h41f822b5, 32'hc1e777be, 32'hc19eb863, 32'hc243ffb7, 32'h42c2e0ce, 32'hc25f2b4f};
test_bias[658:658] = '{32'hc273adda};
test_output[658:658] = '{32'hc4b0e892};
test_input[5272:5279] = '{32'h41ff94b3, 32'hc28c3e72, 32'hc298b79f, 32'hc2bc672a, 32'h42406ef1, 32'hc2080d84, 32'h42010fc3, 32'h42afed5f};
test_weights[5272:5279] = '{32'hc1006346, 32'h429bafba, 32'h429172e0, 32'hc1b0df39, 32'h429bd5f9, 32'h41880239, 32'h424b582b, 32'hbfe76568};
test_bias[659:659] = '{32'hc28117cf};
test_output[659:659] = '{32'hc58fb315};
test_input[5280:5287] = '{32'hc159b03e, 32'hc2b9eee3, 32'h41e3d6ee, 32'h4240b180, 32'hc2c37da0, 32'h4293d180, 32'hc2b37f57, 32'h41e82d24};
test_weights[5280:5287] = '{32'hc10cd982, 32'hc2502197, 32'h426af50e, 32'hc1a00b21, 32'hc1fb6557, 32'h422a0a20, 32'h41a098b6, 32'h3f8c9f16};
test_bias[660:660] = '{32'hc2a6d16e};
test_output[660:660] = '{32'h461caa17};
test_input[5288:5295] = '{32'h429aa598, 32'hc226754e, 32'hc2b3d50b, 32'h4292d65c, 32'h42a7321b, 32'hc2a1d270, 32'hc29e11a5, 32'h42c15542};
test_weights[5288:5295] = '{32'h429cf2e9, 32'h41fd65dc, 32'h42bc8f77, 32'h424691e2, 32'h42704545, 32'hc121c983, 32'hc2053820, 32'hc27b3f79};
test_bias[661:661] = '{32'h42a29da7};
test_output[661:661] = '{32'h4515e8d1};
test_input[5296:5303] = '{32'hc2546808, 32'hc2b3c57b, 32'hc2c379d5, 32'hc27287bb, 32'h42a1f069, 32'h42b5b786, 32'h428eecc5, 32'h427b93df};
test_weights[5296:5303] = '{32'h42257b59, 32'hc0ab2d1b, 32'h4286e4f0, 32'h4268194b, 32'hc2135211, 32'hc1f4a5dd, 32'hc27d16cf, 32'hc24c3942};
test_bias[662:662] = '{32'hc27ce9c9};
test_output[662:662] = '{32'hc6c64deb};
test_input[5304:5311] = '{32'h42b15321, 32'hc2450d79, 32'h42b4d576, 32'hc27984d2, 32'h42b0e802, 32'hc258eae0, 32'hc0db2c90, 32'hc2bab7cd};
test_weights[5304:5311] = '{32'hc266e837, 32'hc28feb51, 32'h42678544, 32'h4212fae3, 32'hc0fc8f03, 32'hc2a7c4b7, 32'hc276b317, 32'hc2a7db2f};
test_bias[663:663] = '{32'hc2aa6318};
test_output[663:663] = '{32'h46513e0e};
test_input[5312:5319] = '{32'hc2a9194e, 32'hc26ddb6c, 32'h40010344, 32'h429f6510, 32'hc2b11002, 32'hc2a020c5, 32'hc23a2c01, 32'h42a14190};
test_weights[5312:5319] = '{32'hc28447fd, 32'hc23a6fe1, 32'h421437b9, 32'h42c14a2f, 32'hc2ba3259, 32'h42bf2313, 32'hc0c41a3a, 32'hc28d8d29};
test_bias[664:664] = '{32'h41d465fa};
test_output[664:664] = '{32'h4631223e};
test_input[5320:5327] = '{32'hc21631ab, 32'h4233b4e3, 32'hc11c19b5, 32'hc231f7cb, 32'h42c4846b, 32'hc2c0568d, 32'hc28743f9, 32'h41d60cd9};
test_weights[5320:5327] = '{32'h42547c70, 32'h4242ae1c, 32'hc1aea116, 32'h4239655b, 32'hc1f03165, 32'h41922434, 32'h40833105, 32'h41bed049};
test_bias[665:665] = '{32'h4201169d};
test_output[665:665] = '{32'hc5ba97d6};
test_input[5328:5335] = '{32'h4289435a, 32'hc17fe0df, 32'hc28c648a, 32'hc2bcd3f3, 32'hc2491750, 32'h4229feb5, 32'hc1a790cc, 32'h423f159a};
test_weights[5328:5335] = '{32'hc1d18a0b, 32'h41a18f8a, 32'hc2612f0e, 32'hc2a8e069, 32'hc284583e, 32'hc025d245, 32'hc28b405d, 32'h4193c977};
test_bias[666:666] = '{32'hc291807f};
test_output[666:666] = '{32'h466edff4};
test_input[5336:5343] = '{32'h4291c05c, 32'h42a87f4d, 32'hc2ba8c7f, 32'hc2327ce1, 32'h41d57eb5, 32'hc1b34aff, 32'hc1abe778, 32'h429980a5};
test_weights[5336:5343] = '{32'hc06cfa49, 32'h416623f6, 32'hc2b553d0, 32'hc1e3d3df, 32'hc2bef4a3, 32'hc28318fb, 32'h418478bc, 32'hc2b58fb5};
test_bias[667:667] = '{32'hc1fbb2b2};
test_output[667:667] = '{32'h450bb937};
test_input[5344:5351] = '{32'hc283e1e6, 32'h41b190d7, 32'hc2899a55, 32'hc1fe57bf, 32'hc2beef9e, 32'hc1e177a2, 32'h42233c39, 32'h4230ba47};
test_weights[5344:5351] = '{32'hc10673d3, 32'hc2bcbc75, 32'h425de0ac, 32'hc26487f0, 32'h40a575a4, 32'h425d8c28, 32'h424a7b82, 32'hc28642bc};
test_bias[668:668] = '{32'h425e7dee};
test_output[668:668] = '{32'hc5c93caa};
test_input[5352:5359] = '{32'hc0545770, 32'h414e5983, 32'h423e8b0d, 32'hc2797bec, 32'h429ae8b0, 32'h42add5ee, 32'hc2c533cc, 32'h42c14f8b};
test_weights[5352:5359] = '{32'hc1e3ce51, 32'hc285c032, 32'h42a0700f, 32'h41c47c7d, 32'h42c2a80c, 32'h42c0ce7f, 32'h41a26ab3, 32'hc2286445};
test_bias[669:669] = '{32'hc29cdf6f};
test_output[669:669] = '{32'h4630675c};
test_input[5360:5367] = '{32'h428b8baf, 32'hc1a691a9, 32'h421b2e7d, 32'h427da627, 32'h424389c7, 32'hc22334ca, 32'h4168ec26, 32'hc2807c9d};
test_weights[5360:5367] = '{32'h41b458fb, 32'h425ab8c4, 32'h424c9117, 32'hc2a02185, 32'hc1fc2dff, 32'hc1aa98b9, 32'h426fdf58, 32'h422b0593};
test_bias[670:670] = '{32'hc1e780ae};
test_output[670:670] = '{32'hc5a381ee};
test_input[5368:5375] = '{32'hc261af9d, 32'hc2945d49, 32'hc2c7c8ad, 32'h4273d975, 32'hc2a4aad6, 32'h4260adfc, 32'h429e5f49, 32'h42a8a41a};
test_weights[5368:5375] = '{32'hc23d0df5, 32'hc28a3c84, 32'hc25feeee, 32'h421e9f79, 32'h42ad0df1, 32'hc2a6275c, 32'hc0b19b2c, 32'h429f218c};
test_bias[671:671] = '{32'h418d999e};
test_output[671:671] = '{32'h4620f1fe};
test_input[5376:5383] = '{32'h427521c3, 32'h427ffd83, 32'h42049aed, 32'h420780e0, 32'hc2a74f49, 32'h429284c5, 32'h423454ba, 32'h427cae1d};
test_weights[5376:5383] = '{32'hc23361ce, 32'hc2903614, 32'h417f5f03, 32'h3fffdfcf, 32'hc27184f3, 32'h428dd495, 32'h4282b1da, 32'hc184a66b};
test_bias[672:672] = '{32'h424dac30};
test_output[672:672] = '{32'h45a9b225};
test_input[5384:5391] = '{32'hc1e2d1df, 32'h420e7009, 32'hc127fd95, 32'h41c77f67, 32'hc19258ce, 32'hc2480a82, 32'hc2b9c46f, 32'hc147eb47};
test_weights[5384:5391] = '{32'hc2b28156, 32'h4287cd59, 32'hc2c1a591, 32'hc0d8232e, 32'hc04b9700, 32'h41f747b9, 32'hbf28858e, 32'hc1f12ec0};
test_bias[673:673] = '{32'hc246cfe4};
test_output[673:673] = '{32'h4592c8ed};
test_input[5392:5399] = '{32'h4267ae06, 32'h42aeaabe, 32'h4252fb87, 32'h428e497e, 32'h42aa0a1a, 32'h42637b12, 32'hc29d4c2d, 32'h423d8456};
test_weights[5392:5399] = '{32'hc1e71b9a, 32'h42b886a9, 32'h40c11b7f, 32'h4207e76c, 32'h4287e628, 32'h428d63ae, 32'hbfb54028, 32'hc25baab4};
test_bias[674:674] = '{32'hc2371113};
test_output[674:674] = '{32'h467ff441};
test_input[5400:5407] = '{32'h420f15a0, 32'h429bb7a6, 32'hc24a557d, 32'h42b2d611, 32'hc2778012, 32'h42b2fdd1, 32'h42043ec6, 32'hc22fb9ea};
test_weights[5400:5407] = '{32'hc2c5b0d1, 32'hc27a2a70, 32'h42aa7594, 32'hc23d8bda, 32'h42c5d0ce, 32'h41a96795, 32'h4295f5e4, 32'h42754e4e};
test_bias[675:675] = '{32'h427deb15};
test_output[675:675] = '{32'hc6a6a45c};
test_input[5408:5415] = '{32'hc2add5dd, 32'h42ade3e8, 32'h42b95fc4, 32'h425a8e7b, 32'h42470110, 32'hc1bd31e5, 32'h40ff6592, 32'hc2149c33};
test_weights[5408:5415] = '{32'h4267a112, 32'hc26499b1, 32'hc23bbc31, 32'h41b56a67, 32'h420ce258, 32'h41e90ece, 32'hc2c4fd02, 32'hc24b6730};
test_bias[676:676] = '{32'hc102f8eb};
test_output[676:676] = '{32'hc62b2bab};
test_input[5416:5423] = '{32'h3ea6d5fa, 32'hc167cf09, 32'hc2627ae6, 32'hc258f018, 32'hc269e97f, 32'h42888b76, 32'h41eeff72, 32'hc297f1b9};
test_weights[5416:5423] = '{32'hc2175db6, 32'h42bf578f, 32'h4174f1b5, 32'hc2995368, 32'h4200f141, 32'h42a79a9e, 32'hc299c9e1, 32'h42970be5};
test_bias[677:677] = '{32'h404419b8};
test_output[677:677] = '{32'hc50fef22};
test_input[5424:5431] = '{32'h42895f72, 32'h42b6f540, 32'h42ac35d8, 32'h425cc4ce, 32'hc25c95a2, 32'hc294bfac, 32'hc0a4898c, 32'h41cf44d6};
test_weights[5424:5431] = '{32'h40cf16ce, 32'hc29063fe, 32'hc1e7af01, 32'h4248f810, 32'hc0cdc841, 32'hc2c21d31, 32'h41e48e86, 32'h4272203a};
test_bias[678:678] = '{32'h411824a8};
test_output[678:678] = '{32'h4543390f};
test_input[5432:5439] = '{32'hc22acb53, 32'h424b73d2, 32'h419807e9, 32'h428edc6e, 32'h422d62fc, 32'h41a321dd, 32'hc2c2b197, 32'hc2c3d3c7};
test_weights[5432:5439] = '{32'hc21765aa, 32'hc284588b, 32'hc2663a9b, 32'h42014f57, 32'h4115163f, 32'h419ce60c, 32'h41f71344, 32'hc247fd07};
test_bias[679:679] = '{32'h4231a85c};
test_output[679:679] = '{32'h4509ad8b};
test_input[5440:5447] = '{32'hc203a570, 32'hc2323ea2, 32'hc2b0c154, 32'h41dcf4d0, 32'hc2c22243, 32'h41fc7e3b, 32'hc138f203, 32'h4221bb66};
test_weights[5440:5447] = '{32'h42c09d8f, 32'hc2830e74, 32'h428c9075, 32'hbfb39fc6, 32'h421444f9, 32'h41a3a682, 32'h420ed419, 32'h41c5f9cd};
test_bias[680:680] = '{32'hc29b25ed};
test_output[680:680] = '{32'hc60bb766};
test_input[5448:5455] = '{32'hc23f830d, 32'h42a1f966, 32'h429b5b91, 32'h420ec271, 32'h42bec916, 32'hc2393078, 32'hc258c88a, 32'hc2b9b78a};
test_weights[5448:5455] = '{32'h42617d61, 32'h4095ce59, 32'hc2529e43, 32'h4250ca11, 32'hc1843aa8, 32'hc2bee52e, 32'hc22b5e07, 32'hc28c2b60};
test_bias[681:681] = '{32'hc2928d4c};
test_output[681:681] = '{32'h45dc5d9a};
test_input[5456:5463] = '{32'hc2ac34e0, 32'h40e02c5b, 32'hc2352e1c, 32'h42c40f3b, 32'h4092c00f, 32'hc28f2c62, 32'h4235bd46, 32'h42a59eaf};
test_weights[5456:5463] = '{32'hc23a8d4d, 32'h420219f5, 32'h41806900, 32'h42112890, 32'hc20f653e, 32'h42729a13, 32'h42254419, 32'h419000ab};
test_bias[682:682] = '{32'h4281674c};
test_output[682:682] = '{32'h45bb8271};
test_input[5464:5471] = '{32'h42a4310d, 32'hc25dc373, 32'h42877e28, 32'hc28e360d, 32'hc17faed0, 32'hc28cee73, 32'hc2be6ce2, 32'hc1f055c4};
test_weights[5464:5471] = '{32'h42b8580f, 32'h429f9311, 32'hc2b00446, 32'hc10f777e, 32'hc202ba59, 32'h42860ae5, 32'h3fbce33d, 32'h42293910};
test_bias[683:683] = '{32'h42851737};
test_output[683:683] = '{32'hc5f17464};
test_input[5472:5479] = '{32'h41f72cc0, 32'hbf292c6e, 32'hc29e317d, 32'h41af9bd0, 32'h40abf7cd, 32'hc1d6aa57, 32'h42a2e4f6, 32'hc1021a0a};
test_weights[5472:5479] = '{32'h42b39d5e, 32'hc294b927, 32'h4112117c, 32'hc271f6ce, 32'h409485be, 32'h413c760f, 32'h4237536e, 32'hc2b4ba87};
test_bias[684:684] = '{32'h42b54f5e};
test_output[684:684] = '{32'h459d890c};
test_input[5480:5487] = '{32'h4215f1ea, 32'hc21b7bdc, 32'h41a091aa, 32'h42b029e7, 32'h4229e448, 32'h428664ea, 32'hc2bbbc87, 32'hc1994606};
test_weights[5480:5487] = '{32'h40eb8b13, 32'hc2966569, 32'h411095b9, 32'hc2620d51, 32'hc2918dcb, 32'h42b0d5a6, 32'h423e4b22, 32'hbfef811d};
test_bias[685:685] = '{32'hc2a56a9b};
test_output[685:685] = '{32'hc54bb99d};
test_input[5488:5495] = '{32'h42062c4d, 32'hc2c72bd7, 32'hc2800b7c, 32'h42c12169, 32'h41b6db35, 32'hc090eb8b, 32'h40def684, 32'hc12b61a3};
test_weights[5488:5495] = '{32'hc24bb7eb, 32'hc1fe2ea7, 32'h42a22418, 32'h429b6073, 32'h4282b984, 32'hc23faf7e, 32'h4297c12f, 32'h428aab74};
test_bias[686:686] = '{32'hc237d7e0};
test_output[686:686] = '{32'h45a31401};
test_input[5496:5503] = '{32'hc158d24c, 32'h4299a177, 32'hc235f1f4, 32'h41f9a4d2, 32'hc28370ee, 32'hc1de5e44, 32'hc20a951f, 32'hc209cd7b};
test_weights[5496:5503] = '{32'h407914b0, 32'h4283efa7, 32'hc0e89d9f, 32'hc2935bbb, 32'hc2209b34, 32'h405fc43d, 32'hc27e7684, 32'h42a7017a};
test_bias[687:687] = '{32'hc1f61191};
test_output[687:687] = '{32'h4598a192};
test_input[5504:5511] = '{32'h42b7bf74, 32'hbf2cf631, 32'h42487791, 32'h4254f7a4, 32'h42a52390, 32'hc209978a, 32'hc14dd828, 32'hc17c29d4};
test_weights[5504:5511] = '{32'hc2a709b8, 32'hc1f84d21, 32'hc1879748, 32'hc21cd8db, 32'h4217ecfd, 32'h4045f454, 32'hc2415346, 32'hc1953010};
test_bias[688:688] = '{32'h42a16ecb};
test_output[688:688] = '{32'hc5cd19fd};
test_input[5512:5519] = '{32'h409a4811, 32'h411206d4, 32'h4282dbb0, 32'h42ab555a, 32'hc1acfa5f, 32'hc2a827b0, 32'h41f7f093, 32'hc284ab4f};
test_weights[5512:5519] = '{32'h40a9965e, 32'hc19bd20f, 32'h42876a8b, 32'h412d0264, 32'hc2655279, 32'hc2985d6f, 32'h416b0de3, 32'hc26acf0b};
test_bias[689:689] = '{32'hc2a56326};
test_output[689:689] = '{32'h4685b744};
test_input[5520:5527] = '{32'h3e8f315c, 32'h41a4c437, 32'hc2a23228, 32'h42161b40, 32'hc1a2ceea, 32'h420914d1, 32'hc1421aa2, 32'h424e9640};
test_weights[5520:5527] = '{32'hc24c1eae, 32'h413d876e, 32'h41aa1997, 32'hc26bae9c, 32'h4221317e, 32'h411dc913, 32'h41a9c735, 32'h41a4e76d};
test_bias[690:690] = '{32'h429491c8};
test_output[690:690] = '{32'hc54ea779};
test_input[5528:5535] = '{32'h4130472d, 32'hc24fddcc, 32'h42b68bba, 32'h41a44fcb, 32'h42869965, 32'hc1b9e9b1, 32'h42c64f31, 32'hc21f146f};
test_weights[5528:5535] = '{32'h417021fe, 32'hc2b0efce, 32'hc2846f7b, 32'h42499712, 32'hc2ae338f, 32'hc2a90ecf, 32'h424bad2d, 32'h4224e241};
test_bias[691:691] = '{32'hc2b772df};
test_output[691:691] = '{32'hc44e6c9c};
test_input[5536:5543] = '{32'hc287f909, 32'hc2bcc0d7, 32'h41f65632, 32'h4211020c, 32'h3fa13cde, 32'hc1427949, 32'h4290d68c, 32'h42b6cbea};
test_weights[5536:5543] = '{32'h418773c2, 32'h426dfa8e, 32'hc1a1f574, 32'h4249d0eb, 32'h42c4bcd9, 32'hc274b411, 32'hc2a82ec6, 32'h42b31e7d};
test_bias[692:692] = '{32'h428e4dc4};
test_output[692:692] = '{32'hc51ddf00};
test_input[5544:5551] = '{32'hc1fd5082, 32'hc27fb343, 32'h428e7cad, 32'h4199b903, 32'hc139c1bc, 32'h42c64b2d, 32'hc2954e2d, 32'hc29242be};
test_weights[5544:5551] = '{32'h4249d7b3, 32'hc2c46371, 32'hc2bb560b, 32'h411400d1, 32'hc28460d5, 32'h42a1ced4, 32'hc2c262a6, 32'h4196c71c};
test_bias[693:693] = '{32'h40a98285};
test_output[693:693] = '{32'h4648e11a};
test_input[5552:5559] = '{32'hc2b563e2, 32'hc2305211, 32'hc09b73f5, 32'hc2149304, 32'hc2151dd2, 32'hc2c18c18, 32'h42af2b33, 32'h41fc1626};
test_weights[5552:5559] = '{32'h420ffd7f, 32'h42b38fda, 32'h4251939d, 32'h42c1e9f1, 32'hc2210913, 32'hc0b6d541, 32'h428eadb6, 32'h42c1a378};
test_bias[694:694] = '{32'h4291135c};
test_output[694:694] = '{32'h43ad8f87};
test_input[5560:5567] = '{32'hc280b32c, 32'h42092f82, 32'hc0e7ed08, 32'hc20535e6, 32'h426acad3, 32'h42b7516e, 32'h42a17143, 32'hc2045155};
test_weights[5560:5567] = '{32'h42a484a2, 32'hc0711fb3, 32'h424fe560, 32'hc2bf2af7, 32'hc2b55719, 32'h428dbf41, 32'hc20bd5ba, 32'h429c4369};
test_bias[695:695] = '{32'hc2a5fdea};
test_output[695:695] = '{32'hc5d89bec};
test_input[5568:5575] = '{32'hc195c039, 32'hc28cbf4c, 32'hc1d63635, 32'h42c5777f, 32'hc2138079, 32'hc2c1bc72, 32'hc12f983a, 32'hc2589bfc};
test_weights[5568:5575] = '{32'hc28d18ce, 32'h42af350f, 32'hc17458ce, 32'hc29f7c93, 32'h42c2546c, 32'hc1abab9b, 32'h4281b7c3, 32'hc2261f75};
test_bias[696:696] = '{32'hc21f29bd};
test_output[696:696] = '{32'hc6406ef9};
test_input[5576:5583] = '{32'h42562a4f, 32'hc2adb8bb, 32'hc2a704c9, 32'h42c35cbb, 32'h42b1c18f, 32'hc23ad8a1, 32'hc22b9819, 32'hc212d4ef};
test_weights[5576:5583] = '{32'hc29afcc8, 32'hc2a094c4, 32'hc2735b68, 32'hc2400ca2, 32'hc2035381, 32'hc22ae763, 32'hc0f19f74, 32'hc2934022};
test_bias[697:697] = '{32'h423b23cf};
test_output[697:697] = '{32'h45a7b6df};
test_input[5584:5591] = '{32'h42c77b59, 32'hc22aba21, 32'h429f8f68, 32'h4210dd89, 32'hc1c6ba5c, 32'hc2c5b287, 32'h41828066, 32'hc28e6927};
test_weights[5584:5591] = '{32'hc29a626c, 32'hc2619ab0, 32'h41a95149, 32'hc1c29632, 32'h42bdaa82, 32'h412c3b90, 32'hc2c1d9f8, 32'hc150c8e8};
test_bias[698:698] = '{32'hc19a1a95};
test_output[698:698] = '{32'hc605fd58};
test_input[5592:5599] = '{32'hc2b90751, 32'hc287ae28, 32'h425f6a22, 32'hc2549e8a, 32'h42c5082e, 32'hc28b6a76, 32'h419bb983, 32'hc2488dde};
test_weights[5592:5599] = '{32'hc1a33b2c, 32'hc2c386ef, 32'hc1f88fa5, 32'hc1ea011d, 32'hc225db3a, 32'hc26251cb, 32'hc1c0004b, 32'h4233f031};
test_bias[699:699] = '{32'h42565235};
test_output[699:699] = '{32'h45accc0c};
test_input[5600:5607] = '{32'h42af4145, 32'hc246c0f3, 32'hc1e25d87, 32'hc1238021, 32'h3f214675, 32'hc27bf139, 32'hc29bad83, 32'hc2022b6d};
test_weights[5600:5607] = '{32'hc2355766, 32'hc2b69a60, 32'hc267418e, 32'h423d1afa, 32'hc20e38ec, 32'hc1cbe927, 32'h42a1beb0, 32'hc2890e88};
test_bias[700:700] = '{32'h40a55b75};
test_output[700:700] = '{32'hc43dfd62};
test_input[5608:5615] = '{32'h425e9f9b, 32'hc25b0f31, 32'hc265a97b, 32'hc1cf0b90, 32'h42a0d127, 32'h42c69c40, 32'h4259f516, 32'hc19749ff};
test_weights[5608:5615] = '{32'hbfac0e58, 32'h42aa58b9, 32'hc2b7f872, 32'h4164fb09, 32'h40692786, 32'h42109b8d, 32'hc2232d47, 32'hbeaaa1d0};
test_bias[701:701] = '{32'hc1c1ec4d};
test_output[701:701] = '{32'h44e2bcab};
test_input[5616:5623] = '{32'hc1983d65, 32'hc297c992, 32'h426a7cda, 32'hc2c268b3, 32'h429b4ce2, 32'hc238bd10, 32'h416dc012, 32'hc202a307};
test_weights[5616:5623] = '{32'h421fb09c, 32'h41424200, 32'hc22096f8, 32'hc0f5c2de, 32'h41554d27, 32'hc29d8c19, 32'hc18a6102, 32'h40a07a00};
test_bias[702:702] = '{32'hc2890d0b};
test_output[702:702] = '{32'h445ff53b};
test_input[5624:5631] = '{32'hc233b65a, 32'h419e3802, 32'hc29180cb, 32'h42a9b8e5, 32'hc2940a6f, 32'h4243e6fc, 32'h427bb36f, 32'hc2a21350};
test_weights[5624:5631] = '{32'hc214e5f3, 32'hc1568b75, 32'hc2803089, 32'h41f0cc38, 32'hc2c30fbf, 32'hc245d8ea, 32'hc1cbce7f, 32'hc271bd9d};
test_bias[703:703] = '{32'hc13d1642};
test_output[703:703] = '{32'h46828002};
test_input[5632:5639] = '{32'hc0b58842, 32'hc121bf5a, 32'h4208048f, 32'hc2b9a8a3, 32'h42b59d3e, 32'hc285193a, 32'h423fae54, 32'h4294ec04};
test_weights[5632:5639] = '{32'hc1e7d7cb, 32'h4267c1d0, 32'h429dab8d, 32'hc2872730, 32'h3f89383b, 32'hc2b685d1, 32'hc29f536f, 32'hc2c5b4ae};
test_bias[704:704] = '{32'h42c1806c};
test_output[704:704] = '{32'h45625d67};
test_input[5640:5647] = '{32'h4109b30b, 32'h42ae7748, 32'h4236f60c, 32'h3fe558c1, 32'hc27b3041, 32'h3faa22f3, 32'h424f1bb1, 32'h41b30fc9};
test_weights[5640:5647] = '{32'hc0c2a648, 32'hc2809aec, 32'h413a2dd1, 32'h42025eeb, 32'h4263ba94, 32'hc120ef41, 32'hc296f006, 32'h42940464};
test_bias[705:705] = '{32'hc284e7ed};
test_output[705:705] = '{32'hc62b8437};
test_input[5648:5655] = '{32'h41040278, 32'h427af4a0, 32'hc19ee80e, 32'hc236a242, 32'h42991e3c, 32'h41916965, 32'hc2379621, 32'h421a4d44};
test_weights[5648:5655] = '{32'hc2af0dff, 32'h4194aab2, 32'h428451aa, 32'h41a423a9, 32'hc2c564a8, 32'h425007ae, 32'hc2999ddd, 32'hc11e73af};
test_bias[706:706] = '{32'h421c40b0};
test_output[706:706] = '{32'hc5a39dbc};
test_input[5656:5663] = '{32'hc0e3af88, 32'hc111305e, 32'hc1bfdf7f, 32'h42aeaa57, 32'hc1c64e57, 32'h41fd0171, 32'h419a431d, 32'h42b963b8};
test_weights[5656:5663] = '{32'h3ec312ca, 32'hc1c9e75f, 32'h411bf9d9, 32'h4237b94e, 32'hc12073cb, 32'hc18dcbd4, 32'hc1347995, 32'hc1d976f1};
test_bias[707:707] = '{32'hc127d183};
test_output[707:707] = '{32'h446c0556};
test_input[5664:5671] = '{32'h426a7053, 32'h426f7741, 32'hc285bb4f, 32'hc2922fc9, 32'hbfef3de7, 32'hc1e1be21, 32'h42ae2a4e, 32'hc1d5e42c};
test_weights[5664:5671] = '{32'hc224e1c6, 32'hc1c70c97, 32'hc262a6a9, 32'hc2054083, 32'hc26d24a5, 32'hc2bfde32, 32'h42ba69b0, 32'h42589a8d};
test_bias[708:708] = '{32'hc2964131};
test_output[708:708] = '{32'h4637478a};
test_input[5672:5679] = '{32'hc26fa316, 32'hc27934b6, 32'hc0c5dcf6, 32'h42bbeab5, 32'hc2a0a2e6, 32'hc2af7b75, 32'hc232c968, 32'h42c14fed};
test_weights[5672:5679] = '{32'hc182d7b6, 32'h42b0304d, 32'hc29d3e8f, 32'h4219359b, 32'hc28faac9, 32'hc26dde1f, 32'hc26d1c39, 32'hc2a6ae1c};
test_bias[709:709] = '{32'hc1e56b84};
test_output[709:709] = '{32'h45a04917};
test_input[5680:5687] = '{32'h42862d0d, 32'hc1409e5d, 32'hc2a2da8f, 32'h422a57ff, 32'hc28d2ed3, 32'hc2c711ca, 32'h420a4d89, 32'h413c8cbc};
test_weights[5680:5687] = '{32'h41cce8fb, 32'h421bb8b9, 32'h429d09f5, 32'h4273e7b7, 32'hc1b97d3c, 32'h4263fa02, 32'hc26deb81, 32'h4282133a};
test_bias[710:710] = '{32'h426fbf43};
test_output[710:710] = '{32'hc5f42c15};
test_input[5688:5695] = '{32'hc19d8f91, 32'h429c7e5a, 32'hc2a5ae16, 32'h424c53dd, 32'hc2c7c7dc, 32'hc1998cee, 32'h42b9dd86, 32'h41b8d498};
test_weights[5688:5695] = '{32'hc26198d7, 32'h41355ebb, 32'hc25ea1be, 32'h41850926, 32'h4249c995, 32'h4282f01e, 32'hc1406b16, 32'hc2c52703};
test_bias[711:711] = '{32'h421a7ee8};
test_output[711:711] = '{32'hc50924d0};
test_input[5696:5703] = '{32'h41930563, 32'h42579ddb, 32'h429cbeab, 32'hc2a3f1ee, 32'h41097b80, 32'hc2799d02, 32'h4247a807, 32'hc2a61899};
test_weights[5696:5703] = '{32'h4254ddbd, 32'h42a5fa46, 32'h4288ba09, 32'hc22997cc, 32'h42179c6e, 32'hc2a3f210, 32'h42a7eb69, 32'h4159be4a};
test_bias[712:712] = '{32'hc2c07119};
test_output[712:712] = '{32'h46b1444a};
test_input[5704:5711] = '{32'hc0b1fbca, 32'hc2a7ab95, 32'h4272364a, 32'hc08578fe, 32'h41bd8179, 32'h41071fff, 32'hc297df5e, 32'hc183dbb8};
test_weights[5704:5711] = '{32'h42b2b270, 32'hc1a148eb, 32'h413a7a32, 32'hc2a54b7d, 32'hc2bf10ae, 32'h4279e1b3, 32'h41cd9b50, 32'hc29837b3};
test_bias[713:713] = '{32'h42bcb48e};
test_output[713:713] = '{32'hc2bd23b4};
test_input[5712:5719] = '{32'hc21e9d93, 32'hc1b573b3, 32'h4247eaa8, 32'h426291ce, 32'hc24a9e25, 32'h423b45a3, 32'h4216cf70, 32'h41dead0c};
test_weights[5712:5719] = '{32'h423b6134, 32'hc2b653dc, 32'h41aeb3ca, 32'h426cedea, 32'h42805952, 32'h42beaf3b, 32'h4158ddb1, 32'hc1f878c7};
test_bias[714:714] = '{32'hc294c4fe};
test_output[714:714] = '{32'h45aa0e49};
test_input[5720:5727] = '{32'h42acd5b5, 32'h429ebc91, 32'hc2b43400, 32'hc2c68bf4, 32'hc2a94768, 32'hc2baa60a, 32'h4206650a, 32'hc21f917e};
test_weights[5720:5727] = '{32'h42be3902, 32'hc19fa356, 32'hc08deb77, 32'h419a9e6f, 32'h42113bfc, 32'hc29aa40f, 32'hc2b94f37, 32'h42510a6f};
test_bias[715:715] = '{32'hc2815b8a};
test_output[715:715] = '{32'h4579c9f4};
test_input[5728:5735] = '{32'h421dd7fd, 32'hc2463a54, 32'h42171abb, 32'hc1a82d89, 32'h4223fadb, 32'hc28316ed, 32'h42c26be6, 32'hc28b3f5b};
test_weights[5728:5735] = '{32'hc1e4d523, 32'h423f4935, 32'h4195fea0, 32'h428608c7, 32'hc2b836b9, 32'h4245ccae, 32'h428766b9, 32'hc2798a7b};
test_bias[716:716] = '{32'h420e5cc5};
test_output[716:716] = '{32'hc37ffe43};
test_input[5736:5743] = '{32'hc1a5f63d, 32'h42c70e1a, 32'hc1d3bac0, 32'hc204b8c5, 32'h4130213c, 32'hc2a9766c, 32'hc135ac17, 32'h412a47d4};
test_weights[5736:5743] = '{32'h4237163f, 32'hc2846900, 32'h42b24ee5, 32'h429710d1, 32'h42acb7d3, 32'hc24f2bab, 32'h41e608a6, 32'h42bbcb89};
test_bias[717:717] = '{32'h427087c6};
test_output[717:717] = '{32'hc5c5e3fb};
test_input[5744:5751] = '{32'hc2927215, 32'hc2a151bf, 32'h4209875c, 32'h42a9c4eb, 32'hc16f52cb, 32'h40f68554, 32'hc22f55a0, 32'h41d2c75f};
test_weights[5744:5751] = '{32'h420b3729, 32'h421c7788, 32'h401ae94d, 32'h42a9f9e8, 32'hc03834f7, 32'h429b725f, 32'h42630824, 32'h4255101e};
test_bias[718:718] = '{32'h42480cf2};
test_output[718:718] = '{32'h44962503};
test_input[5752:5759] = '{32'h4285fad0, 32'h42c7a38c, 32'h4282ee08, 32'hc28318bf, 32'h417ac210, 32'h425dbc6b, 32'hc2a1e4a5, 32'hc2b6e2f9};
test_weights[5752:5759] = '{32'hc1f4b7ab, 32'hc284dc31, 32'h42c4b1b5, 32'hc2c528ce, 32'h429b4509, 32'h4201ff71, 32'hc2c76fb1, 32'h42afe7af};
test_bias[719:719] = '{32'h41feb039};
test_output[719:719] = '{32'h45e418ec};
test_input[5760:5767] = '{32'hc015886e, 32'h4297901a, 32'h422932bc, 32'h428e86f9, 32'hc281c901, 32'h40de7e5a, 32'h4299c657, 32'hc1afab0c};
test_weights[5760:5767] = '{32'hc1d988ef, 32'hc287950a, 32'hc2aa76ab, 32'hc226acef, 32'hc2281601, 32'hc26dc459, 32'hc297ea77, 32'hc20ee952};
test_bias[720:720] = '{32'hc296d347};
test_output[720:720] = '{32'hc662080f};
test_input[5768:5775] = '{32'hc2c73746, 32'h41f749c1, 32'h4225327c, 32'hc2ab8a5f, 32'hc2af6682, 32'h42a6e5ba, 32'h428b1708, 32'h4284bc68};
test_weights[5768:5775] = '{32'hc2a64f2d, 32'h424dc129, 32'hc1e0b752, 32'hc16f217d, 32'h4222ee4d, 32'h425905fa, 32'hc29a4063, 32'h422ca717};
test_bias[721:721] = '{32'hc201dce4};
test_output[721:721] = '{32'h460389f6};
test_input[5776:5783] = '{32'hc25c26f3, 32'hc29278dd, 32'h41fe3981, 32'hc2b6e450, 32'h428148c8, 32'hc2643d44, 32'h42a90e28, 32'hc2661cdb};
test_weights[5776:5783] = '{32'h4265c44e, 32'h4206950e, 32'hc238568b, 32'h42c32c95, 32'h424eab0e, 32'h4285bf80, 32'h420a5546, 32'hc2a7f33a};
test_bias[722:722] = '{32'h41b4054d};
test_output[722:722] = '{32'hc60824f4};
test_input[5784:5791] = '{32'hc2ac9fab, 32'hc2c57ca3, 32'hc2a6099b, 32'h423c51df, 32'h42152de9, 32'h4296cc3b, 32'hc0e55a48, 32'h4264a34d};
test_weights[5784:5791] = '{32'h4202a9c2, 32'h42312fd3, 32'hbea8d838, 32'h41ed87f6, 32'h408a0f04, 32'h428225e6, 32'h428d3f09, 32'h42b77092};
test_bias[723:723] = '{32'h41d3ba9c};
test_output[723:723] = '{32'h457de27f};
test_input[5792:5799] = '{32'h422f2222, 32'hc2b7eb7f, 32'hc2727bf7, 32'h427b8365, 32'h422fc747, 32'h428c1275, 32'hc2b47ef1, 32'hc258820f};
test_weights[5792:5799] = '{32'hc1a92c84, 32'h421fae22, 32'h3f1fdc67, 32'hc073b2cd, 32'h42bd38c5, 32'hc1d3cebe, 32'hc1e2ea3a, 32'hc299017b};
test_bias[724:724] = '{32'hc25f5865};
test_output[724:724] = '{32'h457ea06b};
test_input[5800:5807] = '{32'hc2a7d2db, 32'hc2c78704, 32'h4230843e, 32'hbfc39bb3, 32'hc2301510, 32'hc208d740, 32'hbf9cc463, 32'h42a739a1};
test_weights[5800:5807] = '{32'h41af48af, 32'h4096156d, 32'h428ff62b, 32'h4297ef27, 32'h421159e6, 32'h429b6369, 32'h42be61dc, 32'hc1f055f3};
test_bias[725:725] = '{32'hc231f5f1};
test_output[725:725] = '{32'hc5c104c9};
test_input[5808:5815] = '{32'hc26ce8e6, 32'hc2014ca6, 32'hc0d1dc44, 32'hc272a0ac, 32'h419b33ad, 32'hc03ace51, 32'h42aa6999, 32'h42b95422};
test_weights[5808:5815] = '{32'hc22f1b40, 32'hc2b2c66a, 32'hc20126c5, 32'hc2418175, 32'h40c8fd2b, 32'h41f53c17, 32'hc2112884, 32'hc272d571};
test_bias[726:726] = '{32'h42c5726a};
test_output[726:726] = '{32'h42274a0c};
test_input[5816:5823] = '{32'hc2b2855a, 32'h412bf4a1, 32'hc27ee6aa, 32'hc20c9dd6, 32'h4232de0d, 32'h4278bcb7, 32'h40928ea6, 32'hc197b42a};
test_weights[5816:5823] = '{32'h41f7358a, 32'h42a48148, 32'h42b11a0e, 32'h410ec658, 32'hc2b88a54, 32'h41fa2a9d, 32'hc1813bc9, 32'h42a04400};
test_bias[727:727] = '{32'hc252807b};
test_output[727:727] = '{32'hc6362a21};
test_input[5824:5831] = '{32'hc25dbeb2, 32'hc2b9ff7a, 32'h42750b6a, 32'hc28f4075, 32'hc2675091, 32'h42256df1, 32'h426ea0cb, 32'h40adaf7d};
test_weights[5824:5831] = '{32'hc2add81f, 32'hc24c96a6, 32'hc2aec333, 32'hc2c5c7c8, 32'h41f377ee, 32'hc18177b0, 32'h41f2b09b, 32'h4288a5db};
test_bias[728:728] = '{32'hc19b7f04};
test_output[728:728] = '{32'h462c74e4};
test_input[5832:5839] = '{32'h429996fa, 32'hc13a5a9e, 32'h418c6872, 32'hc20d7fb5, 32'hc1929e7f, 32'h428f7c20, 32'hc0ae36dc, 32'hc2063d93};
test_weights[5832:5839] = '{32'hc242acf1, 32'hc2459676, 32'h424ef471, 32'hc295cac9, 32'hc29e0978, 32'hc16f9985, 32'h42937fac, 32'hc0d2eb40};
test_bias[729:729] = '{32'hc1e8d680};
test_output[729:729] = '{32'h440bf06c};
test_input[5840:5847] = '{32'h427a3c66, 32'hc293242e, 32'h422718db, 32'hc28d56d6, 32'hc2946589, 32'h4101ecb3, 32'hc2652b65, 32'hc1c181e5};
test_weights[5840:5847] = '{32'h4194c958, 32'hc2a08ef7, 32'hc25d8364, 32'hc2b7d245, 32'h42aff048, 32'h424b1e8e, 32'h42939093, 32'hc0609511};
test_bias[730:730] = '{32'hc044edde};
test_output[730:730] = '{32'h4477d98e};
test_input[5848:5855] = '{32'hc2227329, 32'h401c87de, 32'hc1d1f207, 32'hc08514bd, 32'h4164de3e, 32'h4265bc15, 32'hc1da403a, 32'hc23dc121};
test_weights[5848:5855] = '{32'h4251bab6, 32'h426858bc, 32'h4252a2f1, 32'h4299a64f, 32'hc2bb8ed8, 32'hc0ca94a6, 32'h4285b6a8, 32'hc2bd7f5c};
test_bias[731:731] = '{32'h42203c60};
test_output[731:731] = '{32'hc527af21};
test_input[5856:5863] = '{32'h4220f4cd, 32'hc212ae30, 32'h4180e820, 32'hc1cd105e, 32'hc2b89c14, 32'h425809e1, 32'hc2996db7, 32'hc1e33262};
test_weights[5856:5863] = '{32'hc21fd111, 32'h42610ad8, 32'hc251d4e7, 32'hc289df1d, 32'hc2a30e64, 32'h4235a04c, 32'hc26d97a5, 32'hc2089706};
test_bias[732:732] = '{32'hc24962fa};
test_output[732:732] = '{32'h46468398};
test_input[5864:5871] = '{32'hc2a591d3, 32'h4242790c, 32'h41dc2db7, 32'h41ce7c04, 32'h42b3267e, 32'hc2aeb3c8, 32'hc25e02cd, 32'hc289babd};
test_weights[5864:5871] = '{32'hc29bedc3, 32'h41fe4e9c, 32'h4299471e, 32'hc2ba523c, 32'h429b1e65, 32'hc2478de5, 32'hc2718997, 32'hc29faf99};
test_bias[733:733] = '{32'hc191772a};
test_output[733:733] = '{32'h46d982d1};
test_input[5872:5879] = '{32'hc23b28dd, 32'h4218cab2, 32'h420aaa28, 32'hc00949d2, 32'h42c1713a, 32'h425430fb, 32'h42b640e3, 32'hc2227b8c};
test_weights[5872:5879] = '{32'hc2070da7, 32'h40efd760, 32'h42616ca2, 32'hc25b6310, 32'hc23d2154, 32'h40932a18, 32'h4032308e, 32'h3c1f2ac6};
test_bias[734:734] = '{32'hc2835a9e};
test_output[734:734] = '{32'hc34c3c2e};
test_input[5880:5887] = '{32'h42946ece, 32'hc2ab8cfd, 32'hc16d14c6, 32'hc1922328, 32'hc262539b, 32'h40e329b9, 32'hc281e76d, 32'hc29f96f7};
test_weights[5880:5887] = '{32'h41a67cc1, 32'hc2469d31, 32'h4287c919, 32'hc2a175f1, 32'hc28e3b06, 32'h41c1256d, 32'hc219f471, 32'h42b4122c};
test_bias[735:735] = '{32'hc1bebbb0};
test_output[735:735] = '{32'h45b3f97b};
test_input[5888:5895] = '{32'hc2718451, 32'hc2c6b6ed, 32'hc2bc017e, 32'hc0e8a08e, 32'h42011f8b, 32'h41a8c8cb, 32'h42620b06, 32'h421068db};
test_weights[5888:5895] = '{32'hc27e51dd, 32'hc252ace5, 32'h41bcb2ee, 32'hc278e5fe, 32'hc2909a2a, 32'h4249e223, 32'h42bd0fa4, 32'hc2ab973d};
test_bias[736:736] = '{32'h41c77347};
test_output[736:736] = '{32'h4601cda5};
test_input[5896:5903] = '{32'hc25d86e2, 32'h42a1ceb3, 32'hc286a6c6, 32'hc21e2c8a, 32'h4283cb0b, 32'h42a7faca, 32'hc237c9c9, 32'hc2b8b481};
test_weights[5896:5903] = '{32'hc1acd433, 32'hc1235914, 32'hc167c169, 32'hc2883bc6, 32'hc1de6348, 32'hc294aea6, 32'h422629b5, 32'hc0da7c4a};
test_bias[737:737] = '{32'h429f8bd2};
test_output[737:737] = '{32'hc5a39691};
test_input[5904:5911] = '{32'hc01fc05b, 32'h415a2b74, 32'hc26cdd1a, 32'hc174fc0c, 32'h424eb1b5, 32'hc2b4a12e, 32'hc28f0a0d, 32'hc29fe46d};
test_weights[5904:5911] = '{32'h42359dca, 32'hc2bbafeb, 32'hc238804e, 32'h41ee4bce, 32'h4222b7c7, 32'h42833cbb, 32'hc1d6c1ff, 32'h425ca151};
test_bias[738:738] = '{32'hbee4578e};
test_output[738:738] = '{32'hc5a9c0eb};
test_input[5912:5919] = '{32'hc266a105, 32'h420945f4, 32'h417164a9, 32'hc18e8f45, 32'h4233c8a0, 32'hc1cd4b1b, 32'h4198af1b, 32'h426fe06b};
test_weights[5912:5919] = '{32'hc25752ca, 32'h42c00cfe, 32'h42ac5bbe, 32'hc0d25564, 32'h4145f0a1, 32'h428a3426, 32'h4272c6aa, 32'h40880c1d};
test_bias[739:739] = '{32'hc1e24a1e};
test_output[739:739] = '{32'h45f9826d};
test_input[5920:5927] = '{32'h4227674b, 32'h40a84577, 32'hc2423857, 32'hc2240870, 32'hc1c3aa1a, 32'h42a871df, 32'h42acd8f3, 32'h42c0d269};
test_weights[5920:5927] = '{32'hc2570f55, 32'h423874fa, 32'hc00cc793, 32'hc2c36417, 32'h41a59f82, 32'hc29796f9, 32'h427b9326, 32'h4260a77d};
test_bias[740:740] = '{32'h41255c64};
test_output[740:740] = '{32'h45bde139};
test_input[5928:5935] = '{32'h3f98fac7, 32'hc2862639, 32'h40ee00da, 32'hc24dff61, 32'hc2a0c407, 32'h423fca14, 32'h4195d7fa, 32'hc2344fe4};
test_weights[5928:5935] = '{32'hc1654d55, 32'hc2380dc6, 32'hc2a3d90c, 32'hc2ac9fbe, 32'hc138bbf3, 32'h403d7995, 32'hc240bb80, 32'hc2b4e7d6};
test_bias[741:741] = '{32'h42bfef5b};
test_output[741:741] = '{32'h462fb76d};
test_input[5936:5943] = '{32'hc24b4d6f, 32'h42bce7a3, 32'hbf67b610, 32'h4251d268, 32'h42521660, 32'hc1e5d984, 32'h41df9d5c, 32'hc1464a80};
test_weights[5936:5943] = '{32'hc2891327, 32'hbf8845c3, 32'h428c6a78, 32'hc29b2b59, 32'hbfdf383e, 32'h42887323, 32'hc2a64901, 32'h42b2da62};
test_bias[742:742] = '{32'h420f254d};
test_output[742:742] = '{32'hc5c1b529};
test_input[5944:5951] = '{32'h42b26987, 32'hc2bc2eaa, 32'hc25a103e, 32'hc1ad0393, 32'hc2110c31, 32'h42ba28b1, 32'h4285eedd, 32'h42839ab6};
test_weights[5944:5951] = '{32'hc257dde5, 32'hc2aa0043, 32'hc2c67c48, 32'h42863f58, 32'h424913ba, 32'hc2b65d82, 32'h42a23a1d, 32'h423b4c0e};
test_bias[743:743] = '{32'h429a3957};
test_output[743:743] = '{32'h45a97294};
test_input[5952:5959] = '{32'hc2234c99, 32'h41e8d20a, 32'hc2b8bf40, 32'hc2007852, 32'h4229026e, 32'h42a52b76, 32'hc27b5d7e, 32'h41da7cab};
test_weights[5952:5959] = '{32'h4241f7fb, 32'h4285b7c3, 32'hc158e174, 32'h423e4fb0, 32'h4186bab5, 32'hc2544e83, 32'hc2a61ff9, 32'hc19ba091};
test_bias[744:744] = '{32'hc211abf6};
test_output[744:744] = '{32'h44279afa};
test_input[5960:5967] = '{32'hc2234bd2, 32'h420c597e, 32'h42c2dc76, 32'h419e7567, 32'h414a415b, 32'hc2a19e23, 32'hc2a7fc07, 32'hc2863bdc};
test_weights[5960:5967] = '{32'h42315c9e, 32'h41a487e6, 32'h423dc511, 32'h42896fc6, 32'h4262e43b, 32'h4214ceec, 32'hc2b8b76e, 32'hc2c1994c};
test_bias[745:745] = '{32'hc2bb2f26};
test_output[745:745] = '{32'h4682fcbe};
test_input[5968:5975] = '{32'h409ffc13, 32'hc11520fd, 32'h419a1f7f, 32'h41d98294, 32'hc232b6c8, 32'hc23a25b3, 32'h42c25ad7, 32'h42080ab2};
test_weights[5968:5975] = '{32'hc14439a4, 32'hc26a40d4, 32'hbf39f9cb, 32'hc1b63503, 32'h427de489, 32'hc2864fbc, 32'h41ae491b, 32'h4229213c};
test_bias[746:746] = '{32'h42a07a6f};
test_output[746:746] = '{32'h456bff96};
test_input[5976:5983] = '{32'h41c4a945, 32'h4299f267, 32'h416ff6ba, 32'hc2105ea4, 32'h42ab79f0, 32'hc2510df0, 32'hc2885875, 32'hc13216fd};
test_weights[5976:5983] = '{32'h421fbb9e, 32'h42410b19, 32'hc1c7978d, 32'hc21c1ff7, 32'h42196811, 32'hc2830c04, 32'h423f5998, 32'h425d2d77};
test_bias[747:747] = '{32'h42a65772};
test_output[747:747] = '{32'h460728d4};
test_input[5984:5991] = '{32'h413ae57b, 32'hc274ec65, 32'hc02be812, 32'hc1988a39, 32'hc2a326af, 32'h4295aedb, 32'hc0f392ec, 32'hc231723e};
test_weights[5984:5991] = '{32'hc2c1ab8b, 32'h40c9ffd7, 32'h42b57f7a, 32'h42c1b12c, 32'h42b9d35a, 32'h4138dba7, 32'hc2a2f80d, 32'hc231cf92};
test_bias[748:748] = '{32'hc2412098};
test_output[748:748] = '{32'hc5f3165e};
test_input[5992:5999] = '{32'hc2b86340, 32'h41d8deb7, 32'hc2bde002, 32'h415ab3ae, 32'hc2b3d358, 32'h41fd6fba, 32'h42c7bea7, 32'hc1902bb5};
test_weights[5992:5999] = '{32'h41a91703, 32'hc246a15a, 32'hc2b584cc, 32'h415b4bdf, 32'hc296da85, 32'hc26fbcc3, 32'h42b1b788, 32'h427907ad};
test_bias[749:749] = '{32'hc22ae321};
test_output[749:749] = '{32'h468d6bfa};
test_input[6000:6007] = '{32'h41e1bdaf, 32'h42076c38, 32'hc276bbbd, 32'hc116b1bc, 32'hc2b1307a, 32'h422db91e, 32'hc251db9d, 32'hc27d8426};
test_weights[6000:6007] = '{32'h420e4434, 32'hc2a6d8b7, 32'hc21343b1, 32'h4243d9a9, 32'h424cc87c, 32'h41b03781, 32'h418573ab, 32'h40d609af};
test_bias[750:750] = '{32'h428bb373};
test_output[750:750] = '{32'hc59699db};
test_input[6008:6015] = '{32'hc1a1a00f, 32'h4267ff30, 32'hc2bac877, 32'hc2523d2f, 32'h416da1f3, 32'h4204eb68, 32'hc29e89bc, 32'hc0971d97};
test_weights[6008:6015] = '{32'hc1e4013e, 32'h42b462be, 32'h41734cda, 32'hc22354cc, 32'hc182a749, 32'hc2940e4c, 32'hc2517abf, 32'h42bab83a};
test_bias[751:751] = '{32'h424e2e0d};
test_output[751:751] = '{32'h45ed4359};
test_input[6016:6023] = '{32'hc1b160f3, 32'hc2b5ffdd, 32'hc1968f5f, 32'hc2234957, 32'hc21d868a, 32'h42b6f37e, 32'h41c80867, 32'hc11cf9b1};
test_weights[6016:6023] = '{32'hc2445a9a, 32'hc1f4227d, 32'h4237ca8e, 32'h428e2f97, 32'h412dcd1b, 32'h42466ff1, 32'h42c6759a, 32'hc1393f0c};
test_bias[752:752] = '{32'h426974aa};
test_output[752:752] = '{32'h45d66f65};
test_input[6024:6031] = '{32'h42b36265, 32'hc19972cd, 32'h42413361, 32'h42bf06ab, 32'hc2163ca5, 32'hc1d04bfe, 32'hc205a90f, 32'hc2563d3b};
test_weights[6024:6031] = '{32'h423d8977, 32'hc0a34699, 32'h429794ae, 32'h40ff0492, 32'hc2500e12, 32'hc2b36d5f, 32'h41ddbd0b, 32'hc23adc5e};
test_bias[753:753] = '{32'h41f11f3a};
test_output[753:753] = '{32'h466524e7};
test_input[6032:6039] = '{32'h4227ad0c, 32'h40d41bd3, 32'hc14faf69, 32'hc0e22ae9, 32'h42bf7284, 32'hc283c636, 32'hc2c0756b, 32'h42a915ea};
test_weights[6032:6039] = '{32'h42a03274, 32'h422069cf, 32'h420842e1, 32'hbf2c9928, 32'hc1dcc5aa, 32'hc1604705, 32'hc2b15c9c, 32'hc28df46d};
test_bias[754:754] = '{32'hc2a9b1dc};
test_output[754:754] = '{32'h4574c351};
test_input[6040:6047] = '{32'h4280eb43, 32'hc2a45ea4, 32'hc290f542, 32'hc28f150f, 32'hc172a71d, 32'h42140c2c, 32'hc2a87498, 32'hc093732b};
test_weights[6040:6047] = '{32'h41c30b9d, 32'hbe9cd155, 32'hc1cbd09c, 32'h429baa96, 32'hc25a2b5b, 32'hc1bd04ad, 32'hc293fff2, 32'h429df879};
test_bias[755:755] = '{32'h420a474d};
test_output[755:755] = '{32'h45693272};
test_input[6048:6055] = '{32'h42152080, 32'hc2b2a5c1, 32'hc23ba709, 32'h41a3c61d, 32'h42696e03, 32'h4275c204, 32'hc0f450c2, 32'hc1e03cb7};
test_weights[6048:6055] = '{32'h41918419, 32'h42352394, 32'hc2bb3145, 32'hc2411ff7, 32'hc2b22533, 32'hc254f660, 32'hc2921a3e, 32'h425f18c8};
test_bias[756:756] = '{32'hc0a52478};
test_output[756:756] = '{32'hc6139107};
test_input[6056:6063] = '{32'h4231eb03, 32'hc23b114c, 32'hc273f0af, 32'h4246a918, 32'hc260f960, 32'hc27ab773, 32'h418bf867, 32'hc2a79e9a};
test_weights[6056:6063] = '{32'hc2aee4db, 32'hc1e8d5b0, 32'hc26dfc17, 32'h42ae9b96, 32'hc295d62f, 32'hc218cd3d, 32'hc23eebf0, 32'h42b124d6};
test_bias[757:757] = '{32'h4287fb38};
test_output[757:757] = '{32'h4570d970};
test_input[6064:6071] = '{32'hc2975490, 32'h41207952, 32'hbf88da4d, 32'hc2b8128b, 32'h4290ca90, 32'h42a9c9a9, 32'h41848c37, 32'hc211655a};
test_weights[6064:6071] = '{32'hc2b969a0, 32'hc1b48978, 32'hc2096e65, 32'hc1832ca1, 32'hc24cdcd2, 32'hc27cacad, 32'h4122e382, 32'h42c7894e};
test_bias[758:758] = '{32'h41370c62};
test_output[758:758] = '{32'hc582b523};
test_input[6072:6079] = '{32'h421ab8a5, 32'hc1ec7010, 32'hc0bf7b4c, 32'h42529949, 32'hc20107b4, 32'h422edddd, 32'hc1b50409, 32'h42c64559};
test_weights[6072:6079] = '{32'hbe6deae2, 32'hc293985f, 32'h4247fac5, 32'h424272ce, 32'h4288d4dc, 32'h4225fac7, 32'hc2b045ba, 32'h42176c7c};
test_bias[759:759] = '{32'hc2aaf01b};
test_output[759:759] = '{32'h46179453};
test_input[6080:6087] = '{32'hc08a713a, 32'hc1f2e609, 32'h427330af, 32'hc211f1b7, 32'hc2c7b91f, 32'hc2a8e865, 32'hc1463edb, 32'hc1c920ba};
test_weights[6080:6087] = '{32'hc1b8a362, 32'h42c2382d, 32'hc2141203, 32'h41b4bd42, 32'h42be5d6f, 32'h42c09db9, 32'hc22ed705, 32'hc261c589};
test_bias[760:760] = '{32'h424bd0f3};
test_output[760:760] = '{32'hc6a85d38};
test_input[6088:6095] = '{32'hc22454ce, 32'hc2979290, 32'hc2bdf567, 32'hc2b40c77, 32'h3d2b5a16, 32'hc2bed76a, 32'hc2258132, 32'h4130ed4e};
test_weights[6088:6095] = '{32'h4298448a, 32'hc1322b07, 32'hc293a43f, 32'hc225ff33, 32'h41be9303, 32'h42ad309c, 32'hc23e08f0, 32'h429f3036};
test_bias[761:761] = '{32'h4093d4c2};
test_output[761:761] = '{32'h453ec0d5};
test_input[6096:6103] = '{32'hc2af5432, 32'h41ba37a9, 32'h42906045, 32'hc225ec89, 32'h428b4ced, 32'h42850aa9, 32'h42bc4f70, 32'hc2c70299};
test_weights[6096:6103] = '{32'hc272122d, 32'hc2b43ffc, 32'h41824526, 32'h40e92f60, 32'h41d4cb01, 32'h42be9df9, 32'hc2c2818c, 32'h421e7fe3};
test_bias[762:762] = '{32'h423745a3};
test_output[762:762] = '{32'hc4432b37};
test_input[6104:6111] = '{32'h41b54aea, 32'hbf5b03d7, 32'h42401e5e, 32'h400ee938, 32'h4232751f, 32'h4156ace0, 32'h41b632c7, 32'h41658636};
test_weights[6104:6111] = '{32'h42001f72, 32'h42a4f545, 32'h426e08ff, 32'h420e4fb3, 32'hc005baf8, 32'hc2c6d695, 32'hc2a8395e, 32'hc1d61b7b};
test_bias[763:763] = '{32'hc28c2a96};
test_output[763:763] = '{32'hc34bdc8c};
test_input[6112:6119] = '{32'h428779e0, 32'h41cafc58, 32'hc267c1a0, 32'h42b89394, 32'h42b2ffc8, 32'hc187baee, 32'h423a9522, 32'hc25a9a97};
test_weights[6112:6119] = '{32'h41c3517f, 32'h422ff1d4, 32'hc208e0bb, 32'hc27fe8f9, 32'h4289f110, 32'h427c0efd, 32'hc2a6c221, 32'hc0efb287};
test_bias[764:764] = '{32'h422cc70a};
test_output[764:764] = '{32'h4400cb2b};
test_input[6120:6127] = '{32'h41bcbbc2, 32'hc2907c45, 32'hc1cee86c, 32'h40cf61b6, 32'hc24816e5, 32'h422134b0, 32'h4193ced5, 32'h41b3945e};
test_weights[6120:6127] = '{32'h3f7520b4, 32'hc1b53051, 32'h42b88dc1, 32'hc198ed66, 32'h41ab19e7, 32'hc1aa8eec, 32'hc21ccfc6, 32'h419eba70};
test_bias[765:765] = '{32'hc07c686b};
test_output[765:765] = '{32'hc53f7a7b};
test_input[6128:6135] = '{32'hc197ed21, 32'h40d7c4b4, 32'h42c68e55, 32'hc219077a, 32'hc28acac3, 32'hc252d6fd, 32'h4218079d, 32'hc255cab1};
test_weights[6128:6135] = '{32'h42b8f93e, 32'hc1ce9eb7, 32'h414c27a3, 32'h4226beed, 32'hc202533b, 32'hc24b5e8c, 32'hc1db9bb4, 32'hc282c82f};
test_bias[766:766] = '{32'h42a03891};
test_output[766:766] = '{32'h45a2f0b3};
test_input[6136:6143] = '{32'h428aadc5, 32'hc2708b7b, 32'h41f3821b, 32'hc22f1fc0, 32'hc2111e2d, 32'hc2c7d9a6, 32'h40decd4a, 32'h414860fc};
test_weights[6136:6143] = '{32'h42a2caf9, 32'hc0dc8cb5, 32'h4265fa96, 32'hc21bb707, 32'hc27771ed, 32'h42821f16, 32'hc1ed7dbf, 32'h42a9cb3f};
test_bias[767:767] = '{32'hc1e11eb2};
test_output[767:767] = '{32'h45be229c};
test_input[6144:6151] = '{32'hc2be82a0, 32'hc109d4d0, 32'hc29ad8d6, 32'hc1fde736, 32'h42943769, 32'h420cceb4, 32'hc1c54a36, 32'h40ee7d72};
test_weights[6144:6151] = '{32'h42c58b80, 32'hc2b067c0, 32'h40653c63, 32'h42487cd5, 32'h4284ee87, 32'h42856c83, 32'h42b74180, 32'h42c5a4da};
test_bias[768:768] = '{32'hc11857e4};
test_output[768:768] = '{32'hc5953bc6};
test_input[6152:6159] = '{32'hc28a36ad, 32'h42342d94, 32'hc2301315, 32'hc28229f6, 32'h42bfb831, 32'h4177c225, 32'h429d74b7, 32'h410dcea9};
test_weights[6152:6159] = '{32'h42a374cb, 32'hc2c1b08c, 32'hc2810add, 32'hc1e726df, 32'h42856f76, 32'hc2896823, 32'hc214ffaa, 32'h42c73f7c};
test_bias[769:769] = '{32'hc28c5dfb};
test_output[769:769] = '{32'hc501dd12};
test_input[6160:6167] = '{32'hc12a4908, 32'h41f8dbe8, 32'hc24f2fee, 32'hc20058f7, 32'h428ae12b, 32'h422e0a25, 32'hc2603af8, 32'hc2a5ee53};
test_weights[6160:6167] = '{32'h425e5f69, 32'h42b5e433, 32'h41b9c683, 32'hc2bc2a0c, 32'h42af20fd, 32'hc208287c, 32'h429a60ad, 32'h42c1f78d};
test_bias[770:770] = '{32'h42b1e1a4};
test_output[770:770] = '{32'hc562f91d};
test_input[6168:6175] = '{32'hc2b43c39, 32'h4274b115, 32'hc18d7952, 32'h41aea4cd, 32'h41b980c0, 32'hc112f0b0, 32'h420b7c90, 32'hc0a9be93};
test_weights[6168:6175] = '{32'h4174f37b, 32'hc2a15824, 32'h423e71a8, 32'hc24f4919, 32'hc0e4a781, 32'hc14665ff, 32'hc207468d, 32'h4292d6c4};
test_bias[771:771] = '{32'hc1474eef};
test_output[771:771] = '{32'hc61b0393};
test_input[6176:6183] = '{32'h4273a1e3, 32'h40caf7d2, 32'h41309cc3, 32'hc0344748, 32'h427cd82e, 32'h422d0b45, 32'hc23a192f, 32'hc2269f40};
test_weights[6176:6183] = '{32'hc22928d6, 32'h4124507f, 32'hc194a6ee, 32'h4206afaf, 32'hc1414676, 32'h42a351a0, 32'hc29cc425, 32'h422852b6};
test_bias[772:772] = '{32'h42a8aa48};
test_output[772:772] = '{32'h44f2152b};
test_input[6184:6191] = '{32'hc2771b45, 32'h4231f5cc, 32'h422de272, 32'hc0ef3aa8, 32'hc2846bd0, 32'hc2a5c6e0, 32'h42081248, 32'hc128e4ac};
test_weights[6184:6191] = '{32'hc1fb25fd, 32'h403c3489, 32'h422f4948, 32'h415a5508, 32'h41e002b4, 32'hc2974b54, 32'hc24096b1, 32'hc2b6bae9};
test_bias[773:773] = '{32'h42107d2d};
test_output[773:773] = '{32'h45ef2147};
test_input[6192:6199] = '{32'h429b10f0, 32'h41ce64a2, 32'hc2053290, 32'hc285060e, 32'hc2456107, 32'hc18f366b, 32'hc22fe7e1, 32'hbe2c1824};
test_weights[6192:6199] = '{32'hc2b986fb, 32'h41c26a85, 32'h411659ba, 32'h423b1254, 32'hc25c4f02, 32'hc1a0cec0, 32'h3ff09d00, 32'h41e27a12};
test_bias[774:774] = '{32'hc24bea3d};
test_output[774:774] = '{32'hc5dc4cd6};
test_input[6200:6207] = '{32'h42229fc7, 32'hc0c24949, 32'hc1c080d6, 32'h4201bdf4, 32'h40d97c15, 32'h41f51c3f, 32'h41393207, 32'hc1871db2};
test_weights[6200:6207] = '{32'h4274ff57, 32'h42bfa14f, 32'hc25cc548, 32'h427f5d28, 32'hc20770ca, 32'hc22c471e, 32'hc24176a5, 32'hc26fd5f7};
test_bias[775:775] = '{32'h42a38d28};
test_output[775:775] = '{32'h4586211a};
test_input[6208:6215] = '{32'hc226217a, 32'h422809f1, 32'h42bb8f6d, 32'hc0b13146, 32'hc24ff9af, 32'hc2340d72, 32'hc290bfe1, 32'h405278c7};
test_weights[6208:6215] = '{32'hc239154b, 32'h4294e9ae, 32'hc24a726f, 32'hc2804881, 32'h40c6bcd4, 32'h408f0ffc, 32'hbfa59349, 32'h42bc5373};
test_bias[776:776] = '{32'h413cf02d};
test_output[776:776] = '{32'h44095857};
test_input[6216:6223] = '{32'hc23b0e5c, 32'hc19d531a, 32'hc27201d6, 32'h429c0f6e, 32'hc1b7b948, 32'h427f2b95, 32'h4241d305, 32'h42004dee};
test_weights[6216:6223] = '{32'h42adb18b, 32'hc24abc82, 32'h419b1e00, 32'h422fdf67, 32'hc2b36eba, 32'h428b22ea, 32'h41ef1eb6, 32'hc19ebed9};
test_bias[777:777] = '{32'h42a9af8e};
test_output[777:777] = '{32'h45cde162};
test_input[6224:6231] = '{32'h42b54b19, 32'hc1609817, 32'hc2aa86cb, 32'hc2ad03b0, 32'h421cc14c, 32'hc113cd5d, 32'h4033dc49, 32'h42583286};
test_weights[6224:6231] = '{32'hc286afaf, 32'hc29135f6, 32'h42676d2c, 32'h429d1991, 32'hc2607cb8, 32'hc12c3ddc, 32'hc287d992, 32'h400b4ccd};
test_bias[778:778] = '{32'hc1d428df};
test_output[778:778] = '{32'hc6948a37};
test_input[6232:6239] = '{32'h41d5f066, 32'hc2b1ffdb, 32'hc182c55b, 32'h41c518ff, 32'hc273c606, 32'hc22686c4, 32'h422e4c64, 32'h42c36332};
test_weights[6232:6239] = '{32'h42b42933, 32'h428c8a55, 32'h42240e58, 32'h42c631cc, 32'h42818c2a, 32'hc296291c, 32'hc1a9d6cb, 32'h41c7f280};
test_bias[779:779] = '{32'hc21001b2};
test_output[779:779] = '{32'hc4b0e6de};
test_input[6240:6247] = '{32'hc27cb358, 32'h421a15d6, 32'hc2300a78, 32'h42440e43, 32'h42b925c4, 32'h429964d1, 32'h40c8e683, 32'h403e4ed7};
test_weights[6240:6247] = '{32'h41cc0120, 32'hc2b6e1f7, 32'h429efadb, 32'hc280d373, 32'h424a0120, 32'h42696a15, 32'hc29c6485, 32'h4021cffc};
test_bias[780:780] = '{32'h4259c634};
test_output[780:780] = '{32'hc53fb4b7};
test_input[6248:6255] = '{32'hc2b9095f, 32'h42b747d0, 32'h416728a4, 32'h428431c7, 32'h42a9b637, 32'h410bcdb6, 32'hc28a5ade, 32'h41e2df96};
test_weights[6248:6255] = '{32'hc22e1e11, 32'hc24d4b46, 32'h42293f17, 32'hc1c1e5fc, 32'hbf405694, 32'h42a3fd33, 32'h425abb80, 32'h42b7cbe3};
test_bias[781:781] = '{32'hc2520802};
test_output[781:781] = '{32'hc50c3425};
test_input[6256:6263] = '{32'hc1be86b2, 32'hc22cc808, 32'h425fc728, 32'hc1c54b14, 32'h4146e72a, 32'hc22e75bb, 32'hc20a9568, 32'hc1e82998};
test_weights[6256:6263] = '{32'hc229f110, 32'h41a4a8ee, 32'h414645ea, 32'h41f42747, 32'h413a5d10, 32'hc1da3226, 32'hc206884d, 32'hc28faae0};
test_bias[782:782] = '{32'h423fdad8};
test_output[782:782] = '{32'h4592bcc0};
test_input[6264:6271] = '{32'h4138467b, 32'h42c619f5, 32'h42a4619c, 32'h4239e489, 32'hc2949b3d, 32'h42a26711, 32'h4284e846, 32'h4221d2b2};
test_weights[6264:6271] = '{32'h4172995e, 32'h423d32f6, 32'h42913fef, 32'h41a11a95, 32'hc0d1b319, 32'h4203783d, 32'h427538c0, 32'h424f471c};
test_bias[783:783] = '{32'hc2867b63};
test_output[783:783] = '{32'h46a43f2a};
test_input[6272:6279] = '{32'hc251cc2e, 32'hc2812464, 32'hc2997ddc, 32'h41d452a5, 32'hc2875f4b, 32'h429d38e4, 32'hc2395cf8, 32'h42bec316};
test_weights[6272:6279] = '{32'h42b39ef9, 32'hc295023d, 32'hc1b8548c, 32'hc2b822a8, 32'hc1e2eb06, 32'h3f7338aa, 32'h42c2e488, 32'hc21f26cf};
test_bias[784:784] = '{32'h42614091};
test_output[784:784] = '{32'hc5d595bb};
test_input[6280:6287] = '{32'hc1da2e8f, 32'h42a4809b, 32'h429ac4ab, 32'h428dcc8a, 32'h428edd0b, 32'h4242f75f, 32'hc24835c6, 32'hc256dfe7};
test_weights[6280:6287] = '{32'h4163c8da, 32'hc2b0509f, 32'hc2a7899f, 32'hc0a44c01, 32'h42b7715d, 32'h42a840d3, 32'hc2595fb4, 32'h421ca220};
test_bias[785:785] = '{32'h423a1c2d};
test_output[785:785] = '{32'hc546269d};
test_input[6288:6295] = '{32'h428fc812, 32'h40990509, 32'h42baa88f, 32'h42047ed3, 32'h4285e80a, 32'h426593e5, 32'h429a5a6b, 32'h42acb2a6};
test_weights[6288:6295] = '{32'h41a430ed, 32'hc26853de, 32'hc26d836c, 32'hc29d6725, 32'hc1ab0c34, 32'h42adc920, 32'hc2b38fd6, 32'hc1e38ecc};
test_bias[786:786] = '{32'hc289973f};
test_output[786:786] = '{32'hc648c4d1};
test_input[6296:6303] = '{32'hc244d0da, 32'hc01041e2, 32'h428fed64, 32'hc2bb391f, 32'hc201cc51, 32'h42905670, 32'hc2b56b41, 32'hc151821e};
test_weights[6296:6303] = '{32'hc20fb60c, 32'hc232bcc3, 32'h423941b3, 32'h427a4b62, 32'h41e63d86, 32'hc2c6143e, 32'hc22111da, 32'h4209cb93};
test_bias[787:787] = '{32'h428ba166};
test_output[787:787] = '{32'hc5aad21c};
test_input[6304:6311] = '{32'h42ac7077, 32'h427acc0c, 32'hc2384c03, 32'h418dccf2, 32'hc2af5a57, 32'hc29697f6, 32'h41879227, 32'h42981d20};
test_weights[6304:6311] = '{32'hc2a9e0a3, 32'hc2828ef0, 32'hc2c1543b, 32'hc25a2724, 32'h40060b7e, 32'hc2779b91, 32'h4163a34f, 32'hc232f0ef};
test_bias[788:788] = '{32'h42a76c09};
test_output[788:788] = '{32'hc5cc0c38};
test_input[6312:6319] = '{32'h402f61ae, 32'hc2bf059a, 32'hc2096f00, 32'h4287b141, 32'hc29cf4fb, 32'h4132bbaf, 32'h42294495, 32'hc265c6b4};
test_weights[6312:6319] = '{32'hc13e9fee, 32'hc29b1460, 32'h42281c8c, 32'h41e27379, 32'hc2853dfb, 32'h428de6b3, 32'hc06c2abb, 32'hc2937b3e};
test_bias[789:789] = '{32'hc219a3dd};
test_output[789:789] = '{32'h468bf008};
test_input[6320:6327] = '{32'h42c518ca, 32'hc201abff, 32'h428e5cf3, 32'h42aeae62, 32'hc274d3a3, 32'hc0870c50, 32'hc2a04977, 32'h42361698};
test_weights[6320:6327] = '{32'h42bd4bbf, 32'h41283f7c, 32'h42039b94, 32'h3facc71a, 32'hc2a07d80, 32'hc2c2ae11, 32'hc1e9c818, 32'hc02e7b97};
test_bias[790:790] = '{32'h40aaec89};
test_output[790:790] = '{32'h46945fff};
test_input[6328:6335] = '{32'h42c2eff2, 32'hc120e9c3, 32'h4213a7c1, 32'h42a17d25, 32'hc118724c, 32'hc2579ce0, 32'hc29abf46, 32'h425445bc};
test_weights[6328:6335] = '{32'h4183a947, 32'h428f380d, 32'hc2b1317e, 32'hc2b5d97e, 32'hc14c5040, 32'hc2abee09, 32'hc1ff2004, 32'hc162d21a};
test_bias[791:791] = '{32'hc2083d09};
test_output[791:791] = '{32'hc54db9cc};
test_input[6336:6343] = '{32'hc2966b4e, 32'h42c312fc, 32'h42526a72, 32'h42946604, 32'hc279f91f, 32'hc244c7fb, 32'h41b67703, 32'h40aae29f};
test_weights[6336:6343] = '{32'hc278f5c9, 32'h421f7cc6, 32'hc20915ed, 32'hc25720c6, 32'hc1ff2401, 32'hc2ad7eb1, 32'h41dc9ee6, 32'hc05500b4};
test_bias[792:792] = '{32'hc152cc42};
test_output[792:792] = '{32'h46168d45};
test_input[6344:6351] = '{32'h425a37ef, 32'hbf37dbc8, 32'h411cd634, 32'hc2a02d5a, 32'h418a94ea, 32'hc2add1b9, 32'h427db7f1, 32'hc1a8cbdf};
test_weights[6344:6351] = '{32'hc23d917d, 32'hc266b327, 32'h42bc3bc1, 32'hc24aaa17, 32'h42c55a26, 32'h40edb7c4, 32'hc2b7e64d, 32'hc2abc492};
test_bias[793:793] = '{32'hc18b2e77};
test_output[793:793] = '{32'hc4066749};
test_input[6352:6359] = '{32'h422d5422, 32'hc2684b00, 32'hc1da4849, 32'h42919ac9, 32'hc2786d97, 32'h41dfcb99, 32'hc29b093f, 32'hc294c5ee};
test_weights[6352:6359] = '{32'hc2bb4aa9, 32'h4264e7bc, 32'hc28f590a, 32'hc1e00dbc, 32'hc2b7f15c, 32'hc1d9a223, 32'h427afe2f, 32'h4071cf14};
test_bias[794:794] = '{32'h42be42f9};
test_output[794:794] = '{32'hc5ec5bf5};
test_input[6360:6367] = '{32'hc2a5d9f9, 32'h420b273b, 32'h42714419, 32'hc1e8eab9, 32'h41c85fd5, 32'hc1ad6cea, 32'hc1fdf2f9, 32'hc0928dbe};
test_weights[6360:6367] = '{32'hc1f9ec3d, 32'h428bdaf5, 32'h4234eeb3, 32'h3f4f95b6, 32'hc285fcb2, 32'hc207360d, 32'h4291d87a, 32'h42c463f7};
test_bias[795:795] = '{32'hc25af4cc};
test_output[795:795] = '{32'h4577b822};
test_input[6368:6375] = '{32'h419fed84, 32'hc28c959b, 32'hc24227d0, 32'hc29d823b, 32'hc291ca2e, 32'hc2838320, 32'h42a00c86, 32'h42a32f5a};
test_weights[6368:6375] = '{32'h426a547d, 32'h4229db8b, 32'hc26b0cbd, 32'h423126ce, 32'hc2b7451a, 32'h42b868a2, 32'h42b5af39, 32'h427f04dc};
test_bias[796:796] = '{32'hc189dd8c};
test_output[796:796] = '{32'h4625f666};
test_input[6376:6383] = '{32'h4187373a, 32'h428530db, 32'hc17fdb92, 32'h42bf37c5, 32'h41e0b913, 32'h427dd2f9, 32'h429c5c49, 32'h424c8e34};
test_weights[6376:6383] = '{32'hc28ca0e4, 32'h425a1b6a, 32'hc2ba0475, 32'h42978f99, 32'hc2bdd70c, 32'h41ba56c9, 32'hc2972020, 32'h4298c4d5};
test_bias[797:797] = '{32'h42a339af};
test_output[797:797] = '{32'h45fc1b36};
test_input[6384:6391] = '{32'hc21428e9, 32'hc1fe63ac, 32'hc1bf051c, 32'hc2b4a46c, 32'h401b4df2, 32'h427973a3, 32'hc0ac69b5, 32'hc225cbd7};
test_weights[6384:6391] = '{32'hc2853bae, 32'hc10aa679, 32'h419a01a1, 32'h41e57797, 32'h4094d8ee, 32'hc1aecdda, 32'hc081d9ba, 32'h42804c90};
test_bias[798:798] = '{32'hc27f995d};
test_output[798:798] = '{32'hc5883d93};
test_input[6392:6399] = '{32'h421604b9, 32'hc29bb8f2, 32'h406dd590, 32'hc26d0c3d, 32'h42924a2b, 32'h42b15120, 32'h42bd6515, 32'h421a6522};
test_weights[6392:6399] = '{32'h42935153, 32'h426966e9, 32'h42bf028c, 32'h408475a5, 32'hc0a56a06, 32'hc25b3bad, 32'hc29159c0, 32'h42bb3a16};
test_bias[799:799] = '{32'hc222d743};
test_output[799:799] = '{32'hc61fa7ab};
test_input[6400:6407] = '{32'hc2be0e03, 32'h42889779, 32'hc29b4188, 32'h4094fb01, 32'hc29cadfa, 32'hc2bff2eb, 32'hc20d81ba, 32'hc249b661};
test_weights[6400:6407] = '{32'h40b95553, 32'h4295d8ce, 32'h428c9524, 32'h410b96c0, 32'h422555c0, 32'hc26103e8, 32'h42648f12, 32'hc2a27873};
test_bias[800:800] = '{32'h41b779f8};
test_output[800:800] = '{32'h455518d5};
test_input[6408:6415] = '{32'hc16463b1, 32'hc2c053b8, 32'hc19ea7a4, 32'hc2898905, 32'hc2a71eef, 32'h4200a548, 32'hc26e2c62, 32'hc2b7d3b1};
test_weights[6408:6415] = '{32'hc28928f9, 32'hc0c52f4f, 32'h417eb5c3, 32'h41b9c59f, 32'h41675650, 32'h425bcacb, 32'hc1a59a33, 32'h4130b2b3};
test_bias[801:801] = '{32'hc10eb93f};
test_output[801:801] = '{32'h43d5437a};
test_input[6416:6423] = '{32'hc1e77247, 32'hc2632cd6, 32'hc0e5c70f, 32'hc229915f, 32'hc21d09a1, 32'hc21d32ba, 32'h429107f4, 32'hc2be2937};
test_weights[6416:6423] = '{32'hc2992ac9, 32'h42c0acf8, 32'hc29638e1, 32'hc2b2c8a0, 32'h3fe29cf8, 32'hc2b0d485, 32'h424722eb, 32'hc22217c3};
test_bias[802:802] = '{32'h42bb6b44};
test_output[802:802] = '{32'h463c0c20};
test_input[6424:6431] = '{32'h427f2d9e, 32'h41e02b09, 32'h424f534e, 32'h418a1837, 32'h41a2ce3c, 32'h428dcd2f, 32'h4274b9f0, 32'hc122b02d};
test_weights[6424:6431] = '{32'hc2c62e49, 32'hc0dfe04c, 32'hc2240858, 32'hc2a5b934, 32'h42438947, 32'hc23340c7, 32'hc2a5d58e, 32'hc1e2ec5f};
test_bias[803:803] = '{32'hc2888a27};
test_output[803:803] = '{32'hc685a946};
test_input[6432:6439] = '{32'hc0279892, 32'hc28743d1, 32'h42aead6a, 32'h42a6803c, 32'hc2b8ec7a, 32'hc17c59b3, 32'hc2aa4db6, 32'hc2c3e484};
test_weights[6432:6439] = '{32'h4139b173, 32'h429555b1, 32'hc1e448da, 32'hc1e497ab, 32'hc2941200, 32'hc2b392ac, 32'h427b7008, 32'hc1c97492};
test_bias[804:804] = '{32'h4233c44b};
test_output[804:804] = '{32'hc58d9843};
test_input[6440:6447] = '{32'hc25ee8c2, 32'hc1928bf3, 32'h41b398e6, 32'h428f43cc, 32'h42c5a663, 32'h421b8e1d, 32'h427785b7, 32'h41b6cdfe};
test_weights[6440:6447] = '{32'hc2ad688a, 32'hc2c61794, 32'hc2380803, 32'h42461ba2, 32'hc2ab53cb, 32'hc1aa6704, 32'hc2b73835, 32'hc0de8c0d};
test_bias[805:805] = '{32'h412bde50};
test_output[805:805] = '{32'hc5b9f088};
test_input[6448:6455] = '{32'hc2a05ee8, 32'hc2b95ecc, 32'hc2c69f10, 32'hc1e140fd, 32'h42927f6d, 32'hc29e8909, 32'hc1fbcb24, 32'hc18d26ff};
test_weights[6448:6455] = '{32'h41b4b6e7, 32'h423a1b54, 32'h41d6b7a1, 32'hc26a6573, 32'hc2c2d7d0, 32'hc2a08d1c, 32'h41e4b4ae, 32'hc278a8f5};
test_bias[806:806] = '{32'hc228b2b8};
test_output[806:806] = '{32'hc5f2686d};
test_input[6456:6463] = '{32'hc29642e0, 32'h420a04d4, 32'h41e98bdf, 32'hc253e1a8, 32'hc2c4f3ea, 32'h4190d6b0, 32'hc2420730, 32'h41eb39c0};
test_weights[6456:6463] = '{32'h428910c7, 32'h407645d5, 32'h402c74b7, 32'h424cc02d, 32'hc2191557, 32'hc0c7e63f, 32'h42c35d6c, 32'h423981ab};
test_bias[807:807] = '{32'hc298ab6a};
test_output[807:807] = '{32'hc5e8a1c8};
test_input[6464:6471] = '{32'hc281ee9c, 32'h40f644df, 32'h424e8874, 32'h41a115bd, 32'hc1ef1705, 32'hc2412d02, 32'hc1cb6c34, 32'hc265fa67};
test_weights[6464:6471] = '{32'h42afacba, 32'hc18cb63d, 32'h41f9fa55, 32'h42a3aadd, 32'hc259e176, 32'h42159fd9, 32'h4239e674, 32'h42aeb485};
test_bias[808:808] = '{32'h418e8984};
test_output[808:808] = '{32'hc60bc5d5};
test_input[6472:6479] = '{32'h428d5a72, 32'hc2a22f6a, 32'h424ab7c6, 32'hc251916f, 32'h42c03b57, 32'hc25704fa, 32'hc10825f6, 32'hc09e80a8};
test_weights[6472:6479] = '{32'h425f5ba6, 32'hc2a8c937, 32'h4254f677, 32'h411f9ad1, 32'h4057cf69, 32'hc22cef66, 32'h416d51ec, 32'h42106c83};
test_bias[809:809] = '{32'h42771c52};
test_output[809:809] = '{32'h46702a8c};
test_input[6480:6487] = '{32'hc1cecf2b, 32'h4289ba02, 32'h42766cd7, 32'h42aeb83b, 32'h420aa264, 32'hc164de36, 32'h41dc41b2, 32'h42865eea};
test_weights[6480:6487] = '{32'hc29723b7, 32'h41195e4d, 32'h421c50a6, 32'h419bebf7, 32'h42040616, 32'h42ad1c4f, 32'h4246cdd5, 32'h41c813cf};
test_bias[810:810] = '{32'h40606e33};
test_output[810:810] = '{32'h4617473d};
test_input[6488:6495] = '{32'hc2843198, 32'h42817058, 32'h42808d51, 32'hc2921f4a, 32'h427ff8e5, 32'hc2a1a796, 32'h42556dcc, 32'hc1f05404};
test_weights[6488:6495] = '{32'h427ad0bb, 32'hc21bf4cf, 32'hc2add0c7, 32'h425e9d38, 32'h417e189c, 32'hc23dff2e, 32'h42993c5b, 32'h4145d4b8};
test_bias[811:811] = '{32'hc2bf2647};
test_output[811:811] = '{32'hc5f51baf};
test_input[6496:6503] = '{32'hc23682b5, 32'hc188c6bb, 32'hc2a00329, 32'h413e64c1, 32'h42831d3f, 32'hc1c169b9, 32'hc23c4666, 32'hc29b8ebc};
test_weights[6496:6503] = '{32'hc2b0fd3d, 32'h42bfcd5d, 32'h42570403, 32'h40fde047, 32'hc26cd795, 32'h4130b25a, 32'hc2c66937, 32'hc295afd5};
test_bias[812:812] = '{32'hc2a4014a};
test_output[812:812] = '{32'h458b1fcf};
test_input[6504:6511] = '{32'h4252d9d1, 32'hc196cc9c, 32'hc100f753, 32'hc1853904, 32'h418d880e, 32'hc2167c2f, 32'h42b88342, 32'hc19f02f6};
test_weights[6504:6511] = '{32'hc2c22336, 32'hc2bb2a19, 32'h428b5f31, 32'h42a821b5, 32'h41c1aaba, 32'hc2be73ac, 32'h4243c051, 32'h409438a4};
test_bias[813:813] = '{32'hc2127570};
test_output[813:813] = '{32'h4540a92c};
test_input[6512:6519] = '{32'h42327604, 32'h419ed1fe, 32'h42013784, 32'h420b4c1c, 32'hc2b3d1fe, 32'h421a2f06, 32'hc10443e3, 32'h42488bfb};
test_weights[6512:6519] = '{32'h422a502a, 32'h42b51d91, 32'h4071767c, 32'h42460ae6, 32'hc2b7c19c, 32'h42a46e39, 32'h42a03a1e, 32'hc2491e82};
test_bias[814:814] = '{32'hc213b60f};
test_output[814:814] = '{32'h4656e51f};
test_input[6520:6527] = '{32'hc2985c5f, 32'hc18f43fb, 32'h42a13ac6, 32'h42819d2a, 32'h41f85d86, 32'hc2adf781, 32'h423d9a74, 32'hc0a752ae};
test_weights[6520:6527] = '{32'h41832021, 32'hc0cd74ef, 32'hc1e213e1, 32'h425e9348, 32'hc10aacd9, 32'h42b4c368, 32'h42c7ca5f, 32'h424ae21a};
test_bias[815:815] = '{32'hc2ac0363};
test_output[815:815] = '{32'hc55e0983};
test_input[6528:6535] = '{32'hc19de036, 32'h3f9ea663, 32'h424d5259, 32'h4276d17b, 32'hc1a92838, 32'hc2854ce8, 32'h41a232dc, 32'hc2231d28};
test_weights[6528:6535] = '{32'h424ed312, 32'h420d8418, 32'hc2540ac9, 32'hc2a9b473, 32'h4287c95d, 32'h426685d7, 32'hc27e94b6, 32'hc143b1f5};
test_bias[816:816] = '{32'h41691f0e};
test_output[816:816] = '{32'hc66a2c7e};
test_input[6536:6543] = '{32'hc193d35b, 32'h41561dc0, 32'hc27caddf, 32'hc234e0aa, 32'h42c03ca6, 32'hc1fb9efc, 32'h42884036, 32'h42bf0eb1};
test_weights[6536:6543] = '{32'hc1e5832d, 32'hc0dbf294, 32'hc11808d5, 32'h42b34399, 32'hc1aff1ad, 32'hc0b97b05, 32'h42bfb5d2, 32'hc203c539};
test_bias[817:817] = '{32'hc2983304};
test_output[817:817] = '{32'hc4cce78a};
test_input[6544:6551] = '{32'hc2505b73, 32'hc0a60a37, 32'h42664694, 32'h426c3e5f, 32'hc18100ad, 32'hc2a62b9d, 32'h41f029d0, 32'hc24a7286};
test_weights[6544:6551] = '{32'hc018923f, 32'hc20217f7, 32'h42189bcc, 32'hc2ac8b3f, 32'h425bf21f, 32'h42159a9c, 32'h42b62881, 32'hbf2a23cf};
test_bias[818:818] = '{32'h429a3ada};
test_output[818:818] = '{32'hc56ab25b};
test_input[6552:6559] = '{32'h406b12cf, 32'hbf2492cd, 32'hc211c66e, 32'hc0e5d507, 32'hc22f69a9, 32'hc207fc56, 32'h42b2558e, 32'hbfe5742f};
test_weights[6552:6559] = '{32'h42b8a019, 32'h42c35778, 32'hc2a1ca1d, 32'h421ffedc, 32'h427d85ef, 32'h403e3f41, 32'hc1dbc71e, 32'h422cc1e6};
test_bias[819:819] = '{32'h4113f94b};
test_output[819:819] = '{32'hc519d319};
test_input[6560:6567] = '{32'h4288a0f9, 32'h425865a5, 32'h429c48d1, 32'h4228642e, 32'hc2b48cd5, 32'h42c16cfd, 32'hc0c87b15, 32'h428069d2};
test_weights[6560:6567] = '{32'h40660f62, 32'hc18e8654, 32'hc2901c80, 32'h421aa54c, 32'hc247b472, 32'h4297fda3, 32'hc2156cf1, 32'hc1dbfdf3};
test_bias[820:820] = '{32'hc1dfb477};
test_output[820:820] = '{32'h45ae4018};
test_input[6568:6575] = '{32'h41f735da, 32'hc1c48ab0, 32'h42aba820, 32'h407c72ac, 32'h3f3c5c95, 32'hc19e98d4, 32'h425d8109, 32'hc0ad5329};
test_weights[6568:6575] = '{32'h41cb6492, 32'h426f2c43, 32'hc12d185b, 32'hc28164ee, 32'h429a1932, 32'h41a73b07, 32'hc281b72a, 32'hc1bc45bc};
test_bias[821:821] = '{32'h418130ad};
test_output[821:821] = '{32'hc5b145e2};
test_input[6576:6583] = '{32'hc255248b, 32'h4287f524, 32'h418587b5, 32'hc193fc66, 32'h42bfa3cd, 32'h411fd962, 32'hc2a64173, 32'hc2c63e77};
test_weights[6576:6583] = '{32'h42a02dfe, 32'h407df577, 32'h429caad0, 32'h42c305b7, 32'hc1ddbf22, 32'hc2891c67, 32'hc0e09378, 32'hc215adc2};
test_bias[822:822] = '{32'hc2470fce};
test_output[822:822] = '{32'hc5608543};
test_input[6584:6591] = '{32'h429776f3, 32'hc2ac3726, 32'hc2bcf076, 32'h424f6efa, 32'hc292b088, 32'hc2b00a1e, 32'hc23f5a10, 32'hc24473f7};
test_weights[6584:6591] = '{32'h422a1d4f, 32'hc21ea1af, 32'h40de2328, 32'h42c669ce, 32'h3ea19ab7, 32'h429d9ce8, 32'h4213b472, 32'hc24687bf};
test_bias[823:823] = '{32'h41e5bfda};
test_output[823:823] = '{32'h459805e0};
test_input[6592:6599] = '{32'h420c95dc, 32'hc29d6854, 32'hc19f8a10, 32'h42482aa4, 32'hc2c0fd5a, 32'hc198733c, 32'h4207efdc, 32'hc23d12bf};
test_weights[6592:6599] = '{32'h42000dbe, 32'hc200e717, 32'hc27c6e53, 32'h41f27924, 32'h42a983d4, 32'hc229d343, 32'hc192201e, 32'h426543d9};
test_bias[824:824] = '{32'h424d8313};
test_output[824:824] = '{32'hc5839c42};
test_input[6600:6607] = '{32'hc2b8475d, 32'hc29f0dcf, 32'h4297adb3, 32'hc2253e56, 32'h42780893, 32'h421180aa, 32'hc20d7d59, 32'hc29254df};
test_weights[6600:6607] = '{32'hc286db44, 32'hc2a77fd4, 32'hc242a12b, 32'hc2a4fa1c, 32'hc220a2f5, 32'h413b6510, 32'h4204563a, 32'h42560adb};
test_bias[825:825] = '{32'h426672ce};
test_output[825:825] = '{32'h45abd5c5};
test_input[6608:6615] = '{32'hc20402fd, 32'hc1bd9dca, 32'h41a6d098, 32'hc232dac6, 32'h4110e09c, 32'hc29fb362, 32'h42286262, 32'hc1105c3b};
test_weights[6608:6615] = '{32'hc2b0bef7, 32'h421376c8, 32'h4211f2d2, 32'h42225d78, 32'hc272aeae, 32'hc25f7f92, 32'h42b1b0d4, 32'h42be78d5};
test_bias[826:826] = '{32'hbf3dc913};
test_output[826:826] = '{32'h45f3270c};
test_input[6616:6623] = '{32'h42946d5b, 32'hc0a1b174, 32'hc17eddf9, 32'hc2a41640, 32'h426099d0, 32'hc2c02de2, 32'hc19b23cf, 32'h425a9638};
test_weights[6616:6623] = '{32'h4237280c, 32'hc2954f33, 32'h42501cbe, 32'h42827819, 32'hc1f1f9ea, 32'hc2608815, 32'h422e0c93, 32'h425795fb};
test_bias[827:827] = '{32'hc2a7b3fd};
test_output[827:827] = '{32'h454eb935};
test_input[6624:6631] = '{32'hc14bb174, 32'h4290245f, 32'h42771765, 32'h429996fb, 32'h42a2f3c8, 32'h41c6a8c3, 32'hc187902c, 32'h42986a8f};
test_weights[6624:6631] = '{32'hc22050f2, 32'hc0f93a17, 32'h42968fed, 32'h40fc16b2, 32'hc2aa4f32, 32'hc246d862, 32'hc2246f6f, 32'hbfde05ab};
test_bias[828:828] = '{32'hc2c4d27c};
test_output[828:828] = '{32'hc51c64ad};
test_input[6632:6639] = '{32'h42810ee4, 32'hc0d3b70d, 32'hc2adcf5d, 32'h421a92f6, 32'hc2b4adf4, 32'hc2bd4540, 32'h4284cc8d, 32'hc2c29832};
test_weights[6632:6639] = '{32'hbf4a269e, 32'h4238efc3, 32'h42009650, 32'hc1221a93, 32'hc2a1b228, 32'h4266215e, 32'h421be76a, 32'h42ae7dbc};
test_bias[829:829] = '{32'hc21fb136};
test_output[829:829] = '{32'hc5ee3cc4};
test_input[6640:6647] = '{32'hc2439375, 32'hc25e3c82, 32'h426bf026, 32'h4093a45e, 32'hc28b032b, 32'hc24dbec5, 32'h42af27d2, 32'hc2b89851};
test_weights[6640:6647] = '{32'hc1794810, 32'hc1f8e8f1, 32'hc2bafd2a, 32'h425049d8, 32'h4293cb7d, 32'h423b8d5a, 32'h4258b211, 32'h423ee55c};
test_bias[830:830] = '{32'h4289dbeb};
test_output[830:830] = '{32'hc61b0e4a};
test_input[6648:6655] = '{32'h4100288f, 32'hc2c49871, 32'h42b10927, 32'h429492af, 32'hc239c1fe, 32'h41ef5a68, 32'hc07af9d7, 32'h424274cd};
test_weights[6648:6655] = '{32'hc293faa9, 32'hc25ed032, 32'h420bf653, 32'hc12b1add, 32'hc1b54d45, 32'h42a21e81, 32'hc283777d, 32'hc2279e82};
test_bias[831:831] = '{32'h40fc04c9};
test_output[831:831] = '{32'h460aef8f};
test_input[6656:6663] = '{32'hc085d133, 32'hc2749d03, 32'hc28281ca, 32'hc25c2190, 32'hc2451e32, 32'hc29977c6, 32'hc2b1ce92, 32'h4194350a};
test_weights[6656:6663] = '{32'hc289e767, 32'hc1da8528, 32'h42bd2f6c, 32'h4222b565, 32'h3f709daf, 32'hc2c5420f, 32'hc16cb372, 32'h425b4269};
test_bias[832:832] = '{32'h424e2690};
test_output[832:832] = '{32'h4557bcc7};
test_input[6664:6671] = '{32'h41e5ed57, 32'h429971d3, 32'h4268c174, 32'h41886de4, 32'h42729875, 32'h42a96305, 32'h42150597, 32'h41efe531};
test_weights[6664:6671] = '{32'h422afd5f, 32'hc27ec49f, 32'h4282a894, 32'h42bdb0b5, 32'hc229db0e, 32'h40bb3207, 32'hc1da361e, 32'h4275b6c1};
test_bias[833:833] = '{32'h429dd8ca};
test_output[833:833] = '{32'h44126ea2};
test_input[6672:6679] = '{32'hc02b8dd5, 32'h42743ec2, 32'hc24f019c, 32'h419f0fa4, 32'h42aca8c1, 32'hc2610d8a, 32'h404e45f4, 32'h4273ac7d};
test_weights[6672:6679] = '{32'h420a372f, 32'h425e2099, 32'hc2a979e0, 32'hc1291ac2, 32'hc289afbb, 32'hc1979ac3, 32'h428808c3, 32'h42ac8283};
test_bias[834:834] = '{32'hc235e325};
test_output[834:834] = '{32'h45fac57b};
test_input[6680:6687] = '{32'h42874f6c, 32'h41cecca3, 32'hc2673915, 32'hc18ac2a7, 32'h4149ea3d, 32'h4248a698, 32'hc205a67d, 32'h4236ffd4};
test_weights[6680:6687] = '{32'hc2726d5e, 32'h4126a533, 32'h42c25372, 32'h429b57b2, 32'h42134820, 32'hc09b7628, 32'h42b0e5f8, 32'hc25f5676};
test_bias[835:835] = '{32'h41c6c55e};
test_output[835:835] = '{32'hc67aeb58};
test_input[6688:6695] = '{32'hc02260d4, 32'h42045c06, 32'hc16c1dc7, 32'h421d9a09, 32'h4243e838, 32'h4210150f, 32'hc259e439, 32'h4077c248};
test_weights[6688:6695] = '{32'h416c7f59, 32'h411e7edf, 32'hc25e339e, 32'hc18298f5, 32'hc28542eb, 32'hc2b8ccc7, 32'hc2c24960, 32'hc24eb72f};
test_bias[836:836] = '{32'h422125b8};
test_output[836:836] = '{32'hc4783966};
test_input[6696:6703] = '{32'hc28f4d6d, 32'hc2b27e2d, 32'h4257957b, 32'hc11ce301, 32'h424ce87b, 32'h42999a9c, 32'hc29fbc55, 32'h419da01f};
test_weights[6696:6703] = '{32'hc11f86f9, 32'h3fa622eb, 32'h429eef0f, 32'hc2ba37c5, 32'h419fd48e, 32'hc2c1aad0, 32'hc29d554a, 32'hc280eac3};
test_bias[837:837] = '{32'hc2a67813};
test_output[837:837] = '{32'h4586b49c};
test_input[6704:6711] = '{32'h42a89f51, 32'hc292313d, 32'h429f6698, 32'hc1b935b3, 32'h420e6a54, 32'hc1ab9b57, 32'hc2136730, 32'hc248ce30};
test_weights[6704:6711] = '{32'h41843938, 32'h42b93d43, 32'h3eefc4c1, 32'h40f486e1, 32'h42929b23, 32'hc2bd2a67, 32'hc2a9230d, 32'h42b2991f};
test_bias[838:838] = '{32'h4174b3cc};
test_output[838:838] = '{32'hc50b4b73};
test_input[6712:6719] = '{32'hc29c1a61, 32'hc248227f, 32'hc14d08ae, 32'hc27fca8f, 32'hc1d84bc8, 32'h41c71c1a, 32'hc1c09e5c, 32'hc2906f35};
test_weights[6712:6719] = '{32'h41872130, 32'h412fe207, 32'hc18e2969, 32'hc26007bc, 32'h420cd1cf, 32'hc12ad2ba, 32'h41f5f478, 32'h42a78546};
test_bias[839:839] = '{32'hc293c66e};
test_output[839:839] = '{32'hc5bfddda};
test_input[6720:6727] = '{32'h42aaf6ec, 32'hc1632d24, 32'hc2be09d4, 32'h41aee9d2, 32'hc19af773, 32'h415becd4, 32'hc1c673ac, 32'hc1c98847};
test_weights[6720:6727] = '{32'h42a9abb9, 32'h41d36a71, 32'h4100ec01, 32'h428a8c00, 32'hc0e8cc5b, 32'h4277822f, 32'hc254b3cd, 32'h41fa30fa};
test_bias[840:840] = '{32'h42824af7};
test_output[840:840] = '{32'h460ff61b};
test_input[6728:6735] = '{32'h42b2033d, 32'h42393e8a, 32'h41c12451, 32'h429aa85a, 32'hc2c3f355, 32'hc0d994df, 32'h42b7ec3e, 32'h41214dde};
test_weights[6728:6735] = '{32'h418828b1, 32'hc28164f0, 32'hc20a3eb5, 32'hc2a30f1b, 32'h416ca841, 32'h40bf5a84, 32'hc29f737c, 32'hc22e8f30};
test_bias[841:841] = '{32'hc12d4f03};
test_output[841:841] = '{32'hc68bc92a};
test_input[6736:6743] = '{32'hc2a52a4d, 32'hc2ac634e, 32'h413a425c, 32'hc2b508c3, 32'hc29a7c05, 32'h42b5cf17, 32'h426749bf, 32'h42bdb8b9};
test_weights[6736:6743] = '{32'hc1a71ee9, 32'h4171446e, 32'hc2a374d8, 32'h4291603d, 32'h42b9ba6a, 32'h41acaa77, 32'h421b97a8, 32'hc1af0e37};
test_bias[842:842] = '{32'h42572854};
test_output[842:842] = '{32'hc63ce52f};
test_input[6744:6751] = '{32'hc235f4b5, 32'h423fa3b9, 32'hc285b7b8, 32'h41d8270f, 32'hc14105eb, 32'h422998f6, 32'h40e5d4ec, 32'h42bbb9ff};
test_weights[6744:6751] = '{32'hc228c7a1, 32'hc27424b8, 32'h425052b7, 32'h4169a02a, 32'h4149b272, 32'h420482d0, 32'h400386f1, 32'h40ee6f98};
test_bias[843:843] = '{32'hc2857bca};
test_output[843:843] = '{32'hc50906e8};
test_input[6752:6759] = '{32'h415e6bb1, 32'h41622c04, 32'hc2048b1d, 32'hc1885627, 32'hc2c15136, 32'h42873d1c, 32'hc28438c0, 32'h42987d5b};
test_weights[6752:6759] = '{32'h42484002, 32'hc2c54fc7, 32'hc1d1982d, 32'h42a6ab55, 32'h41bb3550, 32'h4283b6f0, 32'hc240d329, 32'hc18e5839};
test_bias[844:844] = '{32'h42bf37d2};
test_output[844:844] = '{32'h453328cd};
test_input[6760:6767] = '{32'hc27f35e6, 32'h4206f65b, 32'h42618238, 32'h42b17b56, 32'h423434ef, 32'hc259f732, 32'h418061b2, 32'hc112cbc3};
test_weights[6760:6767] = '{32'h4288d2c9, 32'hc21b3dc2, 32'hc286fe8c, 32'hc2330257, 32'hc218e657, 32'h427ab1d3, 32'hc290d5ba, 32'hc278b8be};
test_bias[845:845] = '{32'hc2bceb8c};
test_output[845:845] = '{32'hc69694ba};
test_input[6768:6775] = '{32'hc29a1abd, 32'hc181da4a, 32'h42a8b651, 32'h41a95c3e, 32'h424d8611, 32'h41fd57d1, 32'hc29ac6e0, 32'h42824042};
test_weights[6768:6775] = '{32'h42a1beca, 32'h42c78e47, 32'hc0267fbd, 32'h428bb871, 32'hc1d694d9, 32'h4174605e, 32'h42970b73, 32'hc0a74d09};
test_bias[846:846] = '{32'hc2c7e9b6};
test_output[846:846] = '{32'hc6572be7};
test_input[6776:6783] = '{32'h42692439, 32'h41fdeffe, 32'hc2572b5e, 32'hc2241a73, 32'hc286d1f6, 32'h42b12c63, 32'h42a8cef6, 32'hc2063daa};
test_weights[6776:6783] = '{32'hc285b0f1, 32'hc1cfbe22, 32'hc201c8d1, 32'h42c4fdc6, 32'hc232722f, 32'hc2879800, 32'hc29d58de, 32'hc1d152f9};
test_bias[847:847] = '{32'h41cd8214};
test_output[847:847] = '{32'hc6761c77};
test_input[6784:6791] = '{32'h41bee6af, 32'h41bcee4b, 32'hc28cb0f5, 32'h429a4c1e, 32'hc264b176, 32'h40ed47de, 32'hc1a39f8a, 32'h42bf3bef};
test_weights[6784:6791] = '{32'hc1df6a0e, 32'hc28ca05b, 32'hc1916b5c, 32'h41e8b9c2, 32'hc2bd0268, 32'h429e26a5, 32'h41b5fad0, 32'hc2bd0b07};
test_bias[848:848] = '{32'hc2b4c344};
test_output[848:848] = '{32'hc5167f2f};
test_input[6792:6799] = '{32'hc28adad6, 32'hc298dfbc, 32'hc10e802e, 32'h4170db38, 32'hc285e5d6, 32'h427233e9, 32'hc24abe7d, 32'h426b118d};
test_weights[6792:6799] = '{32'hc2b70d97, 32'h42b792bb, 32'h429bf021, 32'h42930f4c, 32'hc26b0c9e, 32'h42b934b7, 32'h40c7df30, 32'hc0cf1f9a};
test_bias[849:849] = '{32'hc29d882e};
test_output[849:849] = '{32'h46051233};
test_input[6800:6807] = '{32'h42769e23, 32'hc1f3baa0, 32'hc29017d8, 32'h4136218f, 32'hc2119d6c, 32'hc12ef50d, 32'hc0af0e01, 32'hc237fcf9};
test_weights[6800:6807] = '{32'hc1f70adc, 32'hc296e6b8, 32'h4173ae0d, 32'h4296e57c, 32'h42c39339, 32'hc293a8e4, 32'hc29ecc5b, 32'hc293d4b0};
test_bias[850:850] = '{32'h40da0790};
test_output[850:850] = '{32'h449b9c8c};
test_input[6808:6815] = '{32'h427e41b8, 32'h418fc865, 32'hc17f9ca0, 32'h400c806f, 32'h42500140, 32'h41aa20f5, 32'hc1d14411, 32'hc217e12e};
test_weights[6808:6815] = '{32'h421a49c4, 32'h42162ec5, 32'h41a71c4d, 32'h4272daa2, 32'h41bbf30a, 32'h425efcab, 32'hc0a39942, 32'hc25a9205};
test_bias[851:851] = '{32'h41b54285};
test_output[851:851] = '{32'h45ec646f};
test_input[6816:6823] = '{32'hc1ba5853, 32'h42a929ff, 32'h4211efa8, 32'hc2c000a1, 32'hc0993f05, 32'h42154232, 32'hc2839d78, 32'hc19d4262};
test_weights[6816:6823] = '{32'h42002c2a, 32'h416d157c, 32'hc28276b6, 32'h40db4a48, 32'h41c6edfd, 32'h42895960, 32'h41fad472, 32'h41545b38};
test_bias[852:852] = '{32'h42a34599};
test_output[852:852] = '{32'hc5119f62};
test_input[6824:6831] = '{32'hc283a26d, 32'h42c2675a, 32'hc133f0f4, 32'h42b5e9c7, 32'hc1bfbdb6, 32'h427019ae, 32'h3f93f975, 32'h42930282};
test_weights[6824:6831] = '{32'hc2c777c1, 32'h4186e1a1, 32'h410fd822, 32'hc0692067, 32'h41ef8449, 32'h42869507, 32'hc2ab0a8a, 32'h426e2cc8};
test_bias[853:853] = '{32'hc293d77f};
test_output[853:853] = '{32'h466f00a7};
test_input[6832:6839] = '{32'h42681346, 32'h4298fd6e, 32'hc2be59f4, 32'h42c69578, 32'h42a58efb, 32'hc28a8567, 32'hc211076d, 32'h41bcef62};
test_weights[6832:6839] = '{32'hc27d965c, 32'hc234951b, 32'hc2405c40, 32'hc19ab691, 32'h4217fa88, 32'hc19646dd, 32'h41f594d5, 32'h42bf40e2};
test_bias[854:854] = '{32'hc28f7794};
test_output[854:854] = '{32'h4482a0c9};
test_input[6840:6847] = '{32'hbfc7cf49, 32'h429b1236, 32'h3f9c7883, 32'h4089c547, 32'h40fc6088, 32'hc2af16bc, 32'hc1a88b32, 32'hc2807185};
test_weights[6840:6847] = '{32'h40b95d8c, 32'hc096b52a, 32'hc23641b3, 32'hc29d98be, 32'h41e14a01, 32'h42a119a5, 32'hc1ae630b, 32'hc1e36118};
test_bias[855:855] = '{32'hc28092cd};
test_output[855:855] = '{32'hc5a813c0};
test_input[6848:6855] = '{32'h42593ae4, 32'hc14e630a, 32'h40c20954, 32'hc22ca119, 32'h41892f08, 32'h42844e7b, 32'h423604c6, 32'h41e919cb};
test_weights[6848:6855] = '{32'hc285e7ff, 32'h428b709f, 32'hc25ff4cb, 32'hc259356a, 32'h42c55ec9, 32'h3f32a054, 32'hc1b6f8b0, 32'hc2630224};
test_bias[856:856] = '{32'hc2b4d61a};
test_output[856:856] = '{32'hc55f9bc2};
test_input[6856:6863] = '{32'h4134d221, 32'hc1ad1ba1, 32'hc2416205, 32'h429d2ab4, 32'hc20e23f0, 32'h4273048c, 32'hc2989463, 32'hc2ab6d2c};
test_weights[6856:6863] = '{32'h42b1877d, 32'hc1b7d9a3, 32'hc1bb6d7c, 32'hc252eb14, 32'hc28125d2, 32'h42969898, 32'hc2833846, 32'h41a4534e};
test_bias[857:857] = '{32'h423317c8};
test_output[857:857] = '{32'h4607212e};
test_input[6864:6871] = '{32'h41827495, 32'hc2adab69, 32'hc21b75a3, 32'hc28eb1a9, 32'h418240cb, 32'h42458c99, 32'h42b4fc90, 32'hc1384c47};
test_weights[6864:6871] = '{32'hc1258038, 32'h42998bda, 32'hc28ea251, 32'hc2a3fd97, 32'hc2c40a09, 32'hc232cbdb, 32'h4204487a, 32'hc1b0bbea};
test_bias[858:858] = '{32'hc2846f2c};
test_output[858:858] = '{32'h44918127};
test_input[6872:6879] = '{32'h42b923df, 32'h4298bc53, 32'hc2b322ab, 32'h419f2c28, 32'h4278e953, 32'h4016e043, 32'h42847aba, 32'h426d9bd9};
test_weights[6872:6879] = '{32'hc1e2827e, 32'hc1b75dfe, 32'hc2428634, 32'h41a64fb5, 32'h417ba1fc, 32'hc204134b, 32'h41a6d38a, 32'h4173b665};
test_bias[859:859] = '{32'hc1a82f33};
test_output[859:859] = '{32'h455ebe89};
test_input[6880:6887] = '{32'hc2584789, 32'h40be845d, 32'hc2af4c72, 32'h42c27426, 32'h42b05b45, 32'h42ae3e11, 32'hc2882700, 32'hc0d76f10};
test_weights[6880:6887] = '{32'h41ccd0d2, 32'hc0c250de, 32'h4166924c, 32'h426760b1, 32'h42a3180f, 32'hc267aa4b, 32'hc1bd8a6c, 32'h4234ed46};
test_bias[860:860] = '{32'hc1975660};
test_output[860:860] = '{32'h45c7372e};
test_input[6888:6895] = '{32'h42ac53dc, 32'h3efe4c3d, 32'hc2c26011, 32'hc19de966, 32'hc215752a, 32'h424a3c48, 32'hc1d3207c, 32'h3fafc501};
test_weights[6888:6895] = '{32'h3faf7cbf, 32'hc076c81c, 32'h41c08bc4, 32'hc282dc3f, 32'h419952e7, 32'hbf31c42a, 32'h420bdb29, 32'h4241c696};
test_bias[861:861] = '{32'h422b705a};
test_output[861:861] = '{32'hc51bff5c};
test_input[6896:6903] = '{32'hbe3cf615, 32'h3ff79a0f, 32'hc1b757eb, 32'hc269d06f, 32'hc273f517, 32'hc241caae, 32'h4270e731, 32'h42283a06};
test_weights[6896:6903] = '{32'h41f0df6a, 32'h42791de8, 32'h3febd957, 32'h4272aef9, 32'h42b2deb7, 32'hc26069f3, 32'h41dbaec6, 32'h41eadc3a};
test_bias[862:862] = '{32'h4295f787};
test_output[862:862] = '{32'hc54aebdb};
test_input[6904:6911] = '{32'h40e77fba, 32'h425389e9, 32'hc2b57c9c, 32'hc2adce1e, 32'hc2a49e05, 32'hc28dcab1, 32'h42bfc8cc, 32'hc1af79bf};
test_weights[6904:6911] = '{32'hc116b358, 32'h4184708f, 32'h41f90300, 32'h42afd1d1, 32'hc2bc806e, 32'hc2c6c7a4, 32'hc2b8cff3, 32'hc25abb0c};
test_bias[863:863] = '{32'hc20ff008};
test_output[863:863] = '{32'hc51f653e};
test_input[6912:6919] = '{32'h41e8661b, 32'hbfdda527, 32'h42326416, 32'hc20431bc, 32'hc2a9456c, 32'hc0c2388e, 32'hc2b55d04, 32'h41ea0d8e};
test_weights[6912:6919] = '{32'hc29649b1, 32'hc1f7117a, 32'h40a9160b, 32'hc24c8b42, 32'h41ebdf89, 32'hc2795b4d, 32'h42a2a6d7, 32'hc18b797f};
test_bias[864:864] = '{32'hc21ac7a4};
test_output[864:864] = '{32'hc6201195};
test_input[6920:6927] = '{32'h423c6f62, 32'h42ace196, 32'hc1e26857, 32'h41ed7348, 32'h4256fe4b, 32'h41e88763, 32'hc1a0a3d9, 32'hc16e8fcd};
test_weights[6920:6927] = '{32'hc2c4763c, 32'hc1a9f3e8, 32'h420cec29, 32'hc169bd33, 32'h429ac008, 32'hc288defe, 32'h4148ac06, 32'hc2b84bed};
test_bias[865:865] = '{32'h42c3500d};
test_output[865:865] = '{32'hc58cc967};
test_input[6928:6935] = '{32'h42b5ff68, 32'hc2ab0d92, 32'h4249f1be, 32'h428c2f7a, 32'h42796cd2, 32'hc177b3bb, 32'hc23c598f, 32'h4135fecd};
test_weights[6928:6935] = '{32'hc28dfd40, 32'hc28a8ad3, 32'hc14c5af5, 32'h42b6a51e, 32'h42120549, 32'h426d7e8e, 32'h427bc26c, 32'h404a3bd5};
test_bias[866:866] = '{32'h42a5f959};
test_output[866:866] = '{32'h45694b4d};
test_input[6936:6943] = '{32'h42c557b2, 32'h42476863, 32'hc0c76c02, 32'h4283506b, 32'h42091328, 32'hc28d5c5e, 32'hc2bbfc81, 32'h4252d929};
test_weights[6936:6943] = '{32'hc2a43e7f, 32'hc1e1ab83, 32'hc1813bd0, 32'h42bf1709, 32'h42a95ed5, 32'h4269ad97, 32'hc260c208, 32'hc1571257};
test_bias[867:867] = '{32'h42a34671};
test_output[867:867] = '{32'h4391fcbc};
test_input[6944:6951] = '{32'h40bff2be, 32'hc28e7575, 32'h427feb03, 32'hc276a694, 32'hc28862da, 32'hc2be0e6c, 32'h42943b42, 32'hc0fce53c};
test_weights[6944:6951] = '{32'h4215ed7e, 32'h42841586, 32'hc131edca, 32'h4039f930, 32'hc281dd55, 32'hc277321e, 32'h4281683e, 32'h428c8818};
test_bias[868:868] = '{32'h41111efb};
test_output[868:868] = '{32'h460f6fa8};
test_input[6952:6959] = '{32'h42c0da21, 32'h41618f36, 32'hc1dbe65b, 32'hc25408ee, 32'hbf86a73f, 32'hc21568e4, 32'h41f4de35, 32'h420e85f6};
test_weights[6952:6959] = '{32'hc24981b4, 32'h42449817, 32'h421549ac, 32'hc20c046e, 32'h427be11b, 32'h4107a5ce, 32'hc1d204db, 32'hc2989577};
test_bias[869:869] = '{32'hc27bc69d};
test_output[869:869] = '{32'hc5e436d3};
test_input[6960:6967] = '{32'hc18f8b57, 32'h4002107a, 32'hc2782286, 32'hc289307e, 32'h415264af, 32'hc27597e0, 32'h4266c4f8, 32'h424d85e7};
test_weights[6960:6967] = '{32'h42987fb5, 32'hc1721ab2, 32'h4216b7be, 32'h41ff5b6d, 32'hc2967b34, 32'hc1c98111, 32'hc0a1a864, 32'h3fb01906};
test_bias[870:870] = '{32'h4109e2e6};
test_output[870:870] = '{32'hc5ae66b2};
test_input[6968:6975] = '{32'h41951715, 32'hc1984cad, 32'h4249d4ee, 32'h4215407e, 32'hc250e814, 32'h3fe1dd42, 32'hc24074a5, 32'hc2abd3f2};
test_weights[6968:6975] = '{32'h428c6f3d, 32'hc20b90bc, 32'hc163ff12, 32'hc26e8af0, 32'hc2878c46, 32'h42214a43, 32'hc214d64b, 32'hc0b59f07};
test_bias[871:871] = '{32'h429aad38};
test_output[871:871] = '{32'h459c1509};
test_input[6976:6983] = '{32'hc1d264cd, 32'hc17ce1bf, 32'h428b81e5, 32'hc2aa184a, 32'hc22d335f, 32'hbec744ce, 32'hc25f9bfc, 32'hc2b5c4bc};
test_weights[6976:6983] = '{32'hbe2f1425, 32'hc1baf03b, 32'h42abe7b2, 32'h42a1b562, 32'hc1f9d67d, 32'h424b9134, 32'hc167d817, 32'hc106bbbe};
test_bias[872:872] = '{32'h41326d5b};
test_output[872:872] = '{32'h4516bd60};
test_input[6984:6991] = '{32'h4152705c, 32'h42c2b94c, 32'h4232fd41, 32'hc1dd732f, 32'hc1ad3d93, 32'hc089d03d, 32'h42b525f6, 32'h4225de29};
test_weights[6984:6991] = '{32'h428cb82d, 32'h42662746, 32'hc2248d41, 32'h42a1f4e3, 32'hc2a40264, 32'h423072bb, 32'h41219446, 32'hc12ea892};
test_bias[873:873] = '{32'hc134b37b};
test_output[873:873] = '{32'h458c0cf8};
test_input[6992:6999] = '{32'h4259cba2, 32'hc2c16f97, 32'h42ae20e4, 32'h42440880, 32'hc1867898, 32'h4160195e, 32'hc278f283, 32'hc25babb1};
test_weights[6992:6999] = '{32'hc2a17c53, 32'hc2504f6b, 32'hc172acf5, 32'h3fb457d0, 32'hc283f38f, 32'h41c2a6b6, 32'h42bc569d, 32'hc29ad630};
test_bias[874:874] = '{32'h42ba6030};
test_output[874:874] = '{32'hc4294c62};
test_input[7000:7007] = '{32'hc215cfc3, 32'hc2b48abf, 32'hc2c7e814, 32'h428c9f1d, 32'h420408e1, 32'hc211147b, 32'hc25b0909, 32'h4197d057};
test_weights[7000:7007] = '{32'hc1e5ef00, 32'hc2bd81e2, 32'h42217361, 32'h40e7d54a, 32'h42b82300, 32'hc228ec18, 32'hc2668ef0, 32'hc2613d31};
test_bias[875:875] = '{32'hc233179a};
test_output[875:875] = '{32'h4646baa1};
test_input[7008:7015] = '{32'hc221811b, 32'h4270918e, 32'hc23eda12, 32'h42ad5eaf, 32'hc218dae2, 32'hc24e3a98, 32'h42400682, 32'hc1eb89e7};
test_weights[7008:7015] = '{32'hc1df2bd8, 32'hc2948542, 32'hc29100c3, 32'h424969ba, 32'h420d0c61, 32'hc190ab6a, 32'hc1737e9c, 32'hc166539e};
test_bias[876:876] = '{32'h42c2f3d8};
test_output[876:876] = '{32'h45713e1f};
test_input[7016:7023] = '{32'h41920278, 32'h428596a1, 32'hc29e5bb2, 32'h3f157cde, 32'h429dcccd, 32'hc2b8ebb5, 32'hc0b84dcd, 32'hc1a78dcc};
test_weights[7016:7023] = '{32'h41ee11d8, 32'hc14158a1, 32'h4287284d, 32'h429aadef, 32'hc1ac5115, 32'hc189f5d1, 32'hc1f8dffd, 32'hc23731a4};
test_bias[877:877] = '{32'h42a5e1bd};
test_output[877:877] = '{32'hc58b2aba};
test_input[7024:7031] = '{32'hc2ac399c, 32'h423a5ac2, 32'h429a1961, 32'hc1fcb1cc, 32'h4229e235, 32'h42639d93, 32'hc2957cfb, 32'h4298b0d4};
test_weights[7024:7031] = '{32'h42c1fdc3, 32'h42852c06, 32'hc0c6d7e6, 32'hc209f01d, 32'hc1603402, 32'h42826095, 32'h42a43f4c, 32'hc2c693f9};
test_bias[878:878] = '{32'hc28baee4};
test_output[878:878] = '{32'hc66f47a1};
test_input[7032:7039] = '{32'hc22b1335, 32'h42078ee2, 32'h4295c521, 32'h4282f1e8, 32'hc2644072, 32'hc1ff9942, 32'hc20edb33, 32'h41c0b541};
test_weights[7032:7039] = '{32'h41c9aff2, 32'hbf9f0626, 32'hc1e6c37c, 32'h42adb3e6, 32'h42831a92, 32'hc236a640, 32'h4001918a, 32'hc26e8425};
test_bias[879:879] = '{32'h4138535c};
test_output[879:879] = '{32'hc4ab9cba};
test_input[7040:7047] = '{32'hc2075b0c, 32'hc276eca3, 32'hc28c5740, 32'h424ec2bb, 32'hc0a71918, 32'h4285d55a, 32'h4246e438, 32'hc1a016c2};
test_weights[7040:7047] = '{32'h42a73213, 32'hc1b05264, 32'hc254bd88, 32'h4207e951, 32'h42a4523c, 32'hc1c2ca6c, 32'hc2b5066f, 32'hc2bcf6a4};
test_bias[880:880] = '{32'hc2c24d95};
test_output[880:880] = '{32'hc43a5569};
test_input[7048:7055] = '{32'hc16f1fe2, 32'h421c6e74, 32'hc2b9b8dd, 32'h426d503c, 32'h3f78d3c5, 32'hc2a54f42, 32'h4299cd3b, 32'hc28f3eec};
test_weights[7048:7055] = '{32'hc28120db, 32'hc2a1c27b, 32'h42b3cc38, 32'h4267a036, 32'hc2258d15, 32'h42530155, 32'h424b58f2, 32'h3febc886};
test_bias[881:881] = '{32'h41b59210};
test_output[881:881] = '{32'hc5f0f778};
test_input[7056:7063] = '{32'h41cf908e, 32'h424ec310, 32'h4099788e, 32'hc21f98be, 32'h40e7df0b, 32'h429d1e37, 32'h429a9ae7, 32'hc1c7c546};
test_weights[7056:7063] = '{32'h423a05e7, 32'h42bc9844, 32'h41a80f1c, 32'hc28903ef, 32'h4283c67b, 32'hc1c13c32, 32'hbeead509, 32'hc02ccf7d};
test_bias[882:882] = '{32'h4254f177};
test_output[882:882] = '{32'h45ece10a};
test_input[7064:7071] = '{32'h41e6e68b, 32'h42636e5a, 32'h40823a1f, 32'h428920eb, 32'h410ef1ae, 32'hc21091b0, 32'h41efad8d, 32'h4267c34c};
test_weights[7064:7071] = '{32'hc289293a, 32'hc2c22e65, 32'h421d5a34, 32'h42929993, 32'h41f43376, 32'hc2043444, 32'h4291bd7e, 32'hc1b50952};
test_bias[883:883] = '{32'h41e132a3};
test_output[883:883] = '{32'h4255ed9d};
test_input[7072:7079] = '{32'hc29e9693, 32'hc2904846, 32'h4289d7a1, 32'h403302ad, 32'h426413c8, 32'hc2b486bd, 32'hc29196b5, 32'hc2bad8bd};
test_weights[7072:7079] = '{32'hc279b481, 32'h422a94b9, 32'h42b7cf11, 32'hc0ad5b57, 32'h42c18009, 32'h42a5468f, 32'hc2371c16, 32'hc1bcf7cd};
test_bias[884:884] = '{32'hc2c173ab};
test_output[884:884] = '{32'h4636b19b};
test_input[7080:7087] = '{32'h42b63770, 32'hc1af375a, 32'h428393c1, 32'hc25635a5, 32'h426771bc, 32'hc2641b06, 32'h41edde3e, 32'hc2a05e68};
test_weights[7080:7087] = '{32'h41ec8669, 32'h4259c196, 32'h41d95b41, 32'h417bebed, 32'hc15b6317, 32'h42332606, 32'h41b93720, 32'hc29b8524};
test_bias[885:885] = '{32'hc2bc8f70};
test_output[885:885] = '{32'h45b93b7a};
test_input[7088:7095] = '{32'h42a56b5f, 32'h41af45d7, 32'hc2b44b95, 32'hc2881dce, 32'h42ac6846, 32'h41556610, 32'h42a7b82f, 32'h41f21107};
test_weights[7088:7095] = '{32'h422cf157, 32'h42081a4c, 32'hc287d588, 32'hc19e7f77, 32'hc2853909, 32'hc2bfca9d, 32'h428a2daa, 32'h426701e9};
test_bias[886:886] = '{32'hc2749f5a};
test_output[886:886] = '{32'h463f6d9a};
test_input[7096:7103] = '{32'h426b3225, 32'hc1aa275e, 32'h428895fc, 32'h42b36802, 32'h41e37739, 32'hc2749b88, 32'hc26fd290, 32'h41afafb8};
test_weights[7096:7103] = '{32'h421a60d1, 32'hc2635e88, 32'h42bf03c7, 32'h42913b97, 32'h42abe27f, 32'hc29aa8e6, 32'h420b1376, 32'hc20e161d};
test_bias[887:887] = '{32'hc1519b4c};
test_output[887:887] = '{32'h46a292d4};
test_input[7104:7111] = '{32'h428cf9cd, 32'hc2b2168a, 32'hc2b3c7af, 32'h42844bd2, 32'hc0820a16, 32'hc21c43d3, 32'hc2892c98, 32'h42773275};
test_weights[7104:7111] = '{32'hc28af6cc, 32'h41b40b62, 32'hc16a57e5, 32'hc2a5608f, 32'hc1ee4df4, 32'hc211fe6e, 32'hc19b5af1, 32'hc21f7920};
test_bias[888:888] = '{32'h42201eb3};
test_output[888:888] = '{32'hc6259ee3};
test_input[7112:7119] = '{32'hc21c43a7, 32'hc18d9db2, 32'h41e87fb8, 32'h42817bb8, 32'h424c1ab5, 32'h42aac2a3, 32'hc16f4d49, 32'hc2c058ef};
test_weights[7112:7119] = '{32'hc1a74557, 32'h429a2802, 32'hc23941c3, 32'hc29149d6, 32'hc1943dc6, 32'hc2bbb99b, 32'h42b95eaf, 32'h40b9b1d9};
test_bias[889:889] = '{32'hc28753cf};
test_output[889:889] = '{32'hc6894070};
test_input[7120:7127] = '{32'h42a8f42c, 32'hc2527ac8, 32'hc2287993, 32'h3fdbe1b8, 32'hc2523226, 32'h4242e302, 32'h42108725, 32'h40e43240};
test_weights[7120:7127] = '{32'h423d8dd0, 32'h42c71618, 32'hc2275999, 32'h416d2061, 32'hc22a669e, 32'hc2010338, 32'hc28ec5ee, 32'hc2874a3a};
test_bias[890:890] = '{32'h42329c48};
test_output[890:890] = '{32'hc4e0a098};
test_input[7128:7135] = '{32'h410e615c, 32'h4209c20d, 32'hc23c45ac, 32'hc239900e, 32'h422c6049, 32'hc2b897ce, 32'h42a1aba8, 32'hc281b8a3};
test_weights[7128:7135] = '{32'h421bf855, 32'h41fd1ae2, 32'h419549cf, 32'h42c1f200, 32'h4201445d, 32'hc2abe5d4, 32'h424189fc, 32'h41797204};
test_bias[891:891] = '{32'hc2aa98fe};
test_output[891:891] = '{32'h46001f08};
test_input[7136:7143] = '{32'hc16aee4e, 32'hc29d36ed, 32'h42a269dc, 32'hc285f992, 32'hc285401b, 32'hc2c3522c, 32'h42a81cd3, 32'hc151d753};
test_weights[7136:7143] = '{32'hc0bad190, 32'hc2ba89e2, 32'h3fbf417f, 32'hc233c398, 32'h42c676c9, 32'h42331b85, 32'hc2c6325d, 32'h4169e638};
test_bias[892:892] = '{32'hc1a61f29};
test_output[892:892] = '{32'hc60c45b5};
test_input[7144:7151] = '{32'h42c33903, 32'h42374806, 32'h417dec34, 32'h42c2fc7e, 32'h42c558c5, 32'h4230b9fa, 32'hc2c1d663, 32'h42a1a13d};
test_weights[7144:7151] = '{32'hc137407f, 32'hc295a7da, 32'hc2a2d19f, 32'h4230d1f8, 32'hc02bb7dd, 32'h415e5888, 32'hc2ab6715, 32'hc2bf5ec9};
test_bias[893:893] = '{32'hc1f9d84a};
test_output[893:893] = '{32'hc41f67e9};
test_input[7152:7159] = '{32'h42a30e55, 32'h4289c82f, 32'h428afc00, 32'hc1d305d3, 32'hc02489ca, 32'h421d3e5c, 32'h421d3ebb, 32'hc2bee4fb};
test_weights[7152:7159] = '{32'hc2c53cff, 32'hc28635da, 32'hc299b89b, 32'hc291b853, 32'hc2619b25, 32'h42b6fb6b, 32'hc20d224f, 32'hc243e6a5};
test_bias[894:894] = '{32'h4271a833};
test_output[894:894] = '{32'hc60c83d2};
test_input[7160:7167] = '{32'hc24b6af6, 32'hc11bd0ff, 32'hc1fefdd8, 32'hc2518f89, 32'hc2a1fd79, 32'hc2121f16, 32'h42072e04, 32'hc27795f0};
test_weights[7160:7167] = '{32'h42a01904, 32'hc2179292, 32'hc0364504, 32'hc2c0fcb0, 32'hc19152e1, 32'hc29c73a4, 32'h4284214f, 32'h42a0a3a5};
test_bias[895:895] = '{32'h420234ca};
test_output[895:895] = '{32'h453faebd};
test_input[7168:7175] = '{32'hc00d3b16, 32'h4202869e, 32'hc2a50ea4, 32'h428b34e7, 32'hc21849c3, 32'h4210e90d, 32'hc18323bb, 32'h40de15a9};
test_weights[7168:7175] = '{32'hc205c7c1, 32'h429f38e0, 32'hc22545e9, 32'hc08710da, 32'hc21e7910, 32'h42c1f65b, 32'h42adb04f, 32'hc172e9f1};
test_bias[896:896] = '{32'h4282e102};
test_output[896:896] = '{32'h46120809};
test_input[7176:7183] = '{32'hc215a1cb, 32'hc27d2f38, 32'h424b98d8, 32'h421f2339, 32'h42abd840, 32'hc259b442, 32'hc25ce550, 32'hc2a61819};
test_weights[7176:7183] = '{32'hc2b2e0bb, 32'h40d0f937, 32'hc208ca50, 32'h42aca9d6, 32'hc1b64304, 32'h4215b125, 32'h42b16275, 32'hc28ea832};
test_bias[897:897] = '{32'h41d48756};
test_output[897:897] = '{32'h44d28a6f};
test_input[7184:7191] = '{32'hc2af971a, 32'hc2a559a4, 32'h41a7916d, 32'hc20491dd, 32'hbd240d68, 32'hc2bc0d98, 32'h42b4a3f1, 32'h41bcfed9};
test_weights[7184:7191] = '{32'hc1c0b6bf, 32'h426761b7, 32'hc24f27dd, 32'hc1f9fd3b, 32'hc21bfbab, 32'hc2b1e269, 32'hc259bb7d, 32'hc24038f1};
test_bias[898:898] = '{32'h428805e1};
test_output[898:898] = '{32'hc3a7e1ef};
test_input[7192:7199] = '{32'hc2a1cdd6, 32'hc29dec4d, 32'h42aac99c, 32'hc2276e9d, 32'h4124f8ae, 32'hc2a08175, 32'h42c002b5, 32'hc27a2879};
test_weights[7192:7199] = '{32'h421f923c, 32'hc0e8d487, 32'hc282c2ce, 32'hc23f1b7d, 32'h42c5f93e, 32'hc2250b19, 32'h42336ab0, 32'hc1701a9c};
test_bias[899:899] = '{32'h4281408e};
test_output[899:899] = '{32'h4554d289};
test_input[7200:7207] = '{32'h42a1a709, 32'hc2514b2d, 32'hc203cad0, 32'h422e753c, 32'hc2920f8d, 32'h42841450, 32'hc1cd403a, 32'h4254a9a4};
test_weights[7200:7207] = '{32'h42c3b05d, 32'hc299ca01, 32'h42aef514, 32'h41ac6f48, 32'hc230a03e, 32'h42919123, 32'h428b8e3a, 32'hc293e45a};
test_bias[900:900] = '{32'h429cbfe9};
test_output[900:900] = '{32'h464166dd};
test_input[7208:7215] = '{32'hc2760f04, 32'hc1b3821c, 32'h4280807d, 32'hc23b40cc, 32'h423bcd29, 32'hc245c04b, 32'hc20ad3b7, 32'h42a69374};
test_weights[7208:7215] = '{32'h423d945c, 32'h4282d3a2, 32'h42b6957e, 32'hc2682e5a, 32'h423d193a, 32'h40ca8973, 32'hc29e6a9c, 32'hc148cf3e};
test_bias[901:901] = '{32'hc11421e1};
test_output[901:901] = '{32'h45f3c628};
test_input[7216:7223] = '{32'h4215b296, 32'hc26175a4, 32'h42b3f393, 32'hc2bcdeb4, 32'hc2c1c6b3, 32'hc182aedd, 32'h421907a9, 32'h41ace53f};
test_weights[7216:7223] = '{32'hc1c43460, 32'hc08290a1, 32'h414d4bda, 32'hc2665a68, 32'hc285981b, 32'h415211c1, 32'h42284e15, 32'h42ad92eb};
test_bias[902:902] = '{32'hc0dcf0e7};
test_output[902:902] = '{32'h4674631f};
test_input[7224:7231] = '{32'hc2992006, 32'h42c0317e, 32'hc21187c9, 32'h422f038b, 32'h425be4d0, 32'hc275efc9, 32'hc2c0249b, 32'hc1b7e9ac};
test_weights[7224:7231] = '{32'h429ed335, 32'h42abf882, 32'hc1c86516, 32'h42b8b640, 32'hc1bb0423, 32'hc20bd398, 32'h42a5b56a, 32'h42a3d981};
test_bias[903:903] = '{32'hc255f102};
test_output[903:903] = '{32'hc4ed300a};
test_input[7232:7239] = '{32'h426d9a13, 32'hc23a9f1b, 32'hc281d697, 32'h408dba5e, 32'hc2adf7a7, 32'hc27f914c, 32'h42b3ee23, 32'h4209d31e};
test_weights[7232:7239] = '{32'hc2a554d0, 32'h42b60e6a, 32'h42b051ec, 32'hc29f9bc9, 32'h42b74721, 32'h4116d724, 32'h42c5ddb0, 32'h40b80d11};
test_bias[904:904] = '{32'h425b94be};
test_output[904:904] = '{32'hc664f799};
test_input[7240:7247] = '{32'hc24ab094, 32'hc1c86a82, 32'hc23722c3, 32'hc2c5aecc, 32'hc20d9dca, 32'h42c2901e, 32'hc22e9a78, 32'hc2874098};
test_weights[7240:7247] = '{32'hc2b87e16, 32'h419e316a, 32'hc265e41a, 32'hc275ebcc, 32'hc136a185, 32'hc2033f25, 32'h41f33e95, 32'h41d9da4e};
test_bias[905:905] = '{32'hc2c63187};
test_output[905:905] = '{32'h45d57ac2};
test_input[7248:7255] = '{32'hc120bff5, 32'hc062b41c, 32'h3f406323, 32'h42ad5671, 32'h427f1a18, 32'h4225b03c, 32'h4285cbca, 32'hc2b12135};
test_weights[7248:7255] = '{32'hc24aa9a5, 32'h41e4d030, 32'h42b0709b, 32'hc2230635, 32'hc2680a38, 32'hc2bef104, 32'h428f25bd, 32'hc1ee270e};
test_bias[906:906] = '{32'hc23a5db2};
test_output[906:906] = '{32'hc55066f8};
test_input[7256:7263] = '{32'h410153de, 32'hbfcc0dbd, 32'h42b66174, 32'hc1da95be, 32'h425aa05c, 32'h42a82338, 32'h4293928c, 32'h421e2ffd};
test_weights[7256:7263] = '{32'hc2c7b389, 32'hc1f7159d, 32'hc0da30ac, 32'h42bc5ad2, 32'hc27d4881, 32'hc2a89ca7, 32'hc2a01459, 32'hc2ac2216};
test_bias[907:907] = '{32'h40a2dab5};
test_output[907:907] = '{32'hc6b9fb4e};
test_input[7264:7271] = '{32'h3f75b704, 32'h41f59695, 32'h41e1a87a, 32'hc1086783, 32'h428af074, 32'h41179c6a, 32'hc200d305, 32'hc215cdfa};
test_weights[7264:7271] = '{32'hc20ddabb, 32'hc2c257ce, 32'h40dde5a6, 32'h4280af61, 32'hc19cd019, 32'h425a28bb, 32'hc29951c0, 32'hc2907427};
test_bias[908:908] = '{32'hc2a4493f};
test_output[908:908] = '{32'h445b34f3};
test_input[7272:7279] = '{32'hc1ee78e8, 32'h40907b28, 32'hc288aaae, 32'h421934ba, 32'hc2918225, 32'hc2bb63de, 32'hc1a466dd, 32'hc12ae7f9};
test_weights[7272:7279] = '{32'hc0da7600, 32'hc2b3cc0f, 32'h425bd9b3, 32'h419a7608, 32'hc21f8366, 32'h42056a10, 32'hc268f0fa, 32'hc26bb387};
test_bias[909:909] = '{32'h42bce69b};
test_output[909:909] = '{32'hc4be3951};
test_input[7280:7287] = '{32'h41341de2, 32'hc29c1420, 32'h42b0c0eb, 32'h404b75af, 32'h41bb68bd, 32'h42c3c599, 32'h4259daf8, 32'hc258647f};
test_weights[7280:7287] = '{32'h42b0955f, 32'h425a437a, 32'h41f8da5f, 32'h420d5122, 32'hc26802b4, 32'hc2c639b5, 32'hc1206df0, 32'hc1f604f4};
test_bias[910:910] = '{32'h42b686ea};
test_output[910:910] = '{32'hc6203a96};
test_input[7288:7295] = '{32'hc08dab1c, 32'hc26cb2b6, 32'hc16b573f, 32'hc291268e, 32'hc216790f, 32'h422d9e4b, 32'hc11c77e5, 32'hc2c5d630};
test_weights[7288:7295] = '{32'h427d4c1f, 32'h42950cfc, 32'hc2ae152b, 32'hc206a0e1, 32'h42bde759, 32'hc2a7f6d9, 32'h41d0d89e, 32'h42be8efc};
test_bias[911:911] = '{32'hc2bc0953};
test_output[911:911] = '{32'hc68c4d6b};
test_input[7296:7303] = '{32'hc2827e85, 32'hc13c50f8, 32'h41fe213a, 32'hc2b92e2a, 32'h40e0bd63, 32'h4295b7b1, 32'h429b9d92, 32'hc24aad00};
test_weights[7296:7303] = '{32'h41eac3d6, 32'h420d3972, 32'h417a0e33, 32'h42a5e5de, 32'h4228b2d6, 32'h42c31288, 32'h418f02be, 32'hc29558c2};
test_bias[912:912] = '{32'h424f5790};
test_output[912:912] = '{32'h454edf2c};
test_input[7304:7311] = '{32'hc2b6a290, 32'hc1fa9541, 32'hc2a5756b, 32'h429278ad, 32'hc288ede6, 32'h42afc671, 32'hc2666d63, 32'h42c7c274};
test_weights[7304:7311] = '{32'h42389593, 32'h42082e67, 32'hc08e57e9, 32'h416627ee, 32'h41fbd24a, 32'h427808a4, 32'h42241d01, 32'h41b2fefe};
test_bias[913:913] = '{32'hc22a5083};
test_output[913:913] = '{32'hc437e1f5};
test_input[7312:7319] = '{32'h41be2e6c, 32'h42c3da0b, 32'h42888640, 32'hc1cb93f0, 32'h42387fec, 32'h42ae0592, 32'h41c86c01, 32'h41e71ee3};
test_weights[7312:7319] = '{32'h4266a800, 32'h42aac0bd, 32'h423de44c, 32'h426f85b8, 32'hc25b4883, 32'hc1da8aa8, 32'hc27d54ed, 32'h42420e51};
test_bias[914:914] = '{32'hc295a7b8};
test_output[914:914] = '{32'h45c455ef};
test_input[7320:7327] = '{32'hc19aaf56, 32'hc26729a2, 32'h429825c5, 32'hc234b617, 32'h42c76272, 32'hc27ba498, 32'hc22036c8, 32'hc2b6fa0c};
test_weights[7320:7327] = '{32'h41d46b81, 32'h42ad7d64, 32'hc0fd0a15, 32'hc21d73a0, 32'h4105c107, 32'h42bb82bd, 32'hc219068f, 32'h42c7bda9};
test_bias[915:915] = '{32'hc1901c8a};
test_output[915:915] = '{32'hc6851a65};
test_input[7328:7335] = '{32'h42808ab2, 32'h42262f45, 32'h425c986e, 32'h42ae8b67, 32'hc2be98ed, 32'hc15d52ea, 32'h42453175, 32'hc158bc33};
test_weights[7328:7335] = '{32'h4203930c, 32'h42a88d48, 32'hc10b4c92, 32'h4211fd7a, 32'hc13886ca, 32'hc1e9b8c3, 32'h41b05ae7, 32'h41b3763d};
test_bias[916:916] = '{32'hc17195c7};
test_output[916:916] = '{32'h46257e05};
test_input[7336:7343] = '{32'h423fa6fb, 32'h41ea943e, 32'hc29b093d, 32'hc289e0fe, 32'hc25f06a2, 32'hc2b5da46, 32'h42b742f1, 32'h42a9fd94};
test_weights[7336:7343] = '{32'hc20b3d9f, 32'h42b9c956, 32'h40548e93, 32'h40a25821, 32'h4221f7c5, 32'hc22c6908, 32'hc1840508, 32'hc2841f18};
test_bias[917:917] = '{32'hc28050b4};
test_output[917:917] = '{32'hc59ec710};
test_input[7344:7351] = '{32'h415c487e, 32'hc221a237, 32'h4000edfb, 32'h424cfa6f, 32'hc2370a5b, 32'h41e69684, 32'h42908a1e, 32'hc2596727};
test_weights[7344:7351] = '{32'h4242c7b6, 32'hc1d3588b, 32'hc1859929, 32'h4287fbbe, 32'hc11b3b90, 32'hc11d2e97, 32'hc1c94819, 32'h41a50435};
test_bias[918:918] = '{32'hc20b8f3b};
test_output[918:918] = '{32'h45147001};
test_input[7352:7359] = '{32'hc29a789c, 32'hc23228c3, 32'hc2c77464, 32'hc290247a, 32'hc2718c1b, 32'hc1576b40, 32'h4280fcab, 32'h428713e3};
test_weights[7352:7359] = '{32'hc2043daf, 32'h42a2ccd5, 32'h41a72c57, 32'hc292e89e, 32'h4212bc84, 32'h41905e43, 32'hc2b1e167, 32'h41833ff8};
test_bias[919:919] = '{32'hc28afdd3};
test_output[919:919] = '{32'hc59ccec3};
test_input[7360:7367] = '{32'h3f59e1ea, 32'hc0db353e, 32'h416e4dcc, 32'h4203ef50, 32'hc20eee91, 32'h41b54adc, 32'hc1941e64, 32'h41b390d6};
test_weights[7360:7367] = '{32'h4288b06c, 32'hc23aebc7, 32'hc0972fe6, 32'hc21990bc, 32'h42bae484, 32'h42a6d5a1, 32'h401bb54e, 32'hc2567d8b};
test_bias[920:920] = '{32'h42ad6671};
test_output[920:920] = '{32'hc55f1118};
test_input[7368:7375] = '{32'h419aa19d, 32'h41d25366, 32'h41ff3774, 32'h42222fbb, 32'hc2210893, 32'hc2817200, 32'hc2b45810, 32'hc2ad456a};
test_weights[7368:7375] = '{32'h42856540, 32'h42697013, 32'hc2395130, 32'hc2a9daaa, 32'h41545b54, 32'hc2a11c97, 32'hc10f62e3, 32'h421ff648};
test_bias[921:921] = '{32'hc1332d0c};
test_output[921:921] = '{32'hc2ac7be5};
test_input[7376:7383] = '{32'hc1b8336a, 32'hc2064f33, 32'h427ee2d8, 32'hc2348e9f, 32'h42a9ca01, 32'h41897e02, 32'h42a0b8cd, 32'hc28b7721};
test_weights[7376:7383] = '{32'h42867ff0, 32'hc2628940, 32'h42ab1f7e, 32'h42270bdb, 32'hc2c5e348, 32'hc13f6064, 32'hc2b281a3, 32'hc2ac9eec};
test_bias[922:922] = '{32'h419bceca};
test_output[922:922] = '{32'hc5b5dc00};
test_input[7384:7391] = '{32'hc1e309cb, 32'hc1c5fd27, 32'h42710903, 32'hc1c2474f, 32'h41ca6cee, 32'hc285048f, 32'h42563787, 32'hc244be75};
test_weights[7384:7391] = '{32'h3f0c4f56, 32'hc1fed339, 32'h42a217ad, 32'hc2467f37, 32'h424c6e97, 32'h42bb4d8d, 32'h425b69c3, 32'hc2818c23};
test_bias[923:923] = '{32'hc2abdd92};
test_output[923:923] = '{32'h45f8de91};
test_input[7392:7399] = '{32'h3f5a375e, 32'hc1afa646, 32'hc295dbf0, 32'h3faa349a, 32'h4238442d, 32'h42a05259, 32'h4290f0c0, 32'hc2b84157};
test_weights[7392:7399] = '{32'h4266510f, 32'hc1df6b4a, 32'hc2644c65, 32'hc2575ba2, 32'h42b594fc, 32'h416c531c, 32'h419ce4b8, 32'h42aa05b1};
test_bias[924:924] = '{32'hc218292a};
test_output[924:924] = '{32'h456c905d};
test_input[7400:7407] = '{32'hc287b637, 32'h41996b27, 32'h40f7aadc, 32'h42a69080, 32'hc21bd1c5, 32'h42876ff8, 32'h425682a0, 32'h3f1fdf5a};
test_weights[7400:7407] = '{32'h425e6697, 32'hc2be294a, 32'h4223e17e, 32'h425490bc, 32'hc1c48d5e, 32'h4241451c, 32'hc282e9d9, 32'hc116e81b};
test_bias[925:925] = '{32'hc20222bb};
test_output[925:925] = '{32'hc32cffa7};
test_input[7408:7415] = '{32'h42aae122, 32'hc28a8346, 32'h3ee16875, 32'hc189f5aa, 32'h42208c4c, 32'hc1031e67, 32'hc2630365, 32'h42811cf2};
test_weights[7408:7415] = '{32'h42c2dee5, 32'hc2c14b31, 32'hc0853c3b, 32'hc1b90dfa, 32'hc1e71ec7, 32'hc1b142fc, 32'hc29211c6, 32'h429d876b};
test_bias[926:926] = '{32'hc20a17a6};
test_output[926:926] = '{32'h46b8a11d};
test_input[7416:7423] = '{32'hc2a70ad7, 32'hc202e3c8, 32'hc192ad3d, 32'hc2ba6e7b, 32'h428c4bb7, 32'h425e03c4, 32'hc230bdf8, 32'h40a0d8a6};
test_weights[7416:7423] = '{32'h40a82752, 32'hc2351446, 32'h42ae29ac, 32'h411095ba, 32'hc2132f42, 32'h4197293e, 32'h42618791, 32'hc28129fb};
test_bias[927:927] = '{32'h41545ccf};
test_output[927:927] = '{32'hc5b31c6b};
test_input[7424:7431] = '{32'h42379347, 32'h420553b5, 32'h42a168ed, 32'h42198898, 32'h42c5c289, 32'h42b60c69, 32'hc201b714, 32'hc248d712};
test_weights[7424:7431] = '{32'hc0bc531f, 32'h42595527, 32'hc24d8e93, 32'hc27581b3, 32'h42b18d22, 32'h42abad5a, 32'h425eaaa6, 32'hc2805587};
test_bias[928:928] = '{32'hc2a3331c};
test_output[928:928] = '{32'h464a9112};
test_input[7432:7439] = '{32'hc2b4a0ad, 32'h40fd4c8c, 32'hc290e8c0, 32'hc202e50f, 32'h40a325a6, 32'h428892d2, 32'hc24309ce, 32'h427d6e48};
test_weights[7432:7439] = '{32'h4180118d, 32'h42b930e6, 32'h421a30c5, 32'h421196cd, 32'h42a2e4e0, 32'hc20fe6f3, 32'h411b0055, 32'h40e4f040};
test_bias[929:929] = '{32'h42c2dfa6};
test_output[929:929] = '{32'hc5d01f3a};
test_input[7440:7447] = '{32'hc2a8e6f7, 32'h412cab2b, 32'h42887574, 32'h418f75a4, 32'h4291460b, 32'hc2228246, 32'h42a3512b, 32'hc244c17c};
test_weights[7440:7447] = '{32'hc2b3d79c, 32'h42ae974a, 32'h4197ac22, 32'hc250f669, 32'h42af73c8, 32'h42259df1, 32'hc18592d2, 32'hc1e556bd};
test_bias[930:930] = '{32'h42938c67};
test_output[930:930] = '{32'h46561cfa};
test_input[7448:7455] = '{32'h422990c1, 32'hc2029a89, 32'h4288c556, 32'hc1f65a7d, 32'hc2be6dc2, 32'hc226d238, 32'h41b14e40, 32'hc2753f52};
test_weights[7448:7455] = '{32'hc2b639c6, 32'h429c3ea6, 32'hc287288f, 32'hc1a5bced, 32'h4234c7b0, 32'hc22539de, 32'hc27e397d, 32'hc2bffff5};
test_bias[931:931] = '{32'hc2780773};
test_output[931:931] = '{32'hc605c74c};
test_input[7456:7463] = '{32'h41eba151, 32'h4212c0f9, 32'h42252e16, 32'hc1800fc2, 32'h418e50bf, 32'hc27182fb, 32'hc2c79161, 32'hc17cf3e5};
test_weights[7456:7463] = '{32'hc294165e, 32'h4246484c, 32'hc161a9c5, 32'hc2abc7b1, 32'hc2b9ae6d, 32'h41b7ebdb, 32'h417c4f89, 32'h420e0c57};
test_bias[932:932] = '{32'hc2515752};
test_output[932:932] = '{32'hc595e595};
test_input[7464:7471] = '{32'h408797c8, 32'h41cc0386, 32'hc253b4ae, 32'hc0d09895, 32'h4197a988, 32'h40a853ef, 32'hc1e560d8, 32'h41f594fb};
test_weights[7464:7471] = '{32'h420451f2, 32'h4285f514, 32'hc2363b62, 32'h429d940b, 32'h42b0a22f, 32'hc246ad97, 32'hc22804c2, 32'h41324c17};
test_bias[933:933] = '{32'hc2902d74};
test_output[933:933] = '{32'h45cf49f6};
test_input[7472:7479] = '{32'h42842c73, 32'h42bb9562, 32'hc2295d34, 32'h42239658, 32'hc24dfea3, 32'h4268f88e, 32'hc27ac363, 32'h424aba07};
test_weights[7472:7479] = '{32'hc2c1a27a, 32'h4202a7cc, 32'h3eb6dc9a, 32'h424f3a24, 32'h42b288b0, 32'hc2485463, 32'hc281403a, 32'h4299e4f7};
test_bias[934:934] = '{32'h41f3b5fe};
test_output[934:934] = '{32'hc43ee061};
test_input[7480:7487] = '{32'h41a28a4d, 32'h41b58fef, 32'h4220bb15, 32'hc0385f46, 32'h42821f8f, 32'hc2b34c77, 32'h3fe271b0, 32'h42bb9cee};
test_weights[7480:7487] = '{32'h4272d054, 32'h42bfb1c3, 32'h41183e40, 32'h4218f3ec, 32'hc2b20dd2, 32'hc2ac02b5, 32'hc290cad5, 32'hc25b43cb};
test_bias[935:935] = '{32'h40278ef2};
test_output[935:935] = '{32'h43a5a839};
test_input[7488:7495] = '{32'h42ac38f1, 32'hc2660fd3, 32'hc1d98a37, 32'hc2740832, 32'hc2447ca4, 32'hc1979492, 32'h42ba2c92, 32'h42b119be};
test_weights[7488:7495] = '{32'h409a8977, 32'hc2c519d9, 32'h416dae20, 32'h4244933f, 32'hc2ae443a, 32'hc26d6ac4, 32'h42c7fe5b, 32'h41146be2};
test_bias[936:936] = '{32'hc2a54ce0};
test_output[936:936] = '{32'h468dabb5};
test_input[7496:7503] = '{32'h42367871, 32'hc112483a, 32'h42b90a6d, 32'h42a67d3b, 32'h411306d9, 32'hc281ba53, 32'h4204376f, 32'h42a3fe60};
test_weights[7496:7503] = '{32'h42bc7fa4, 32'h429532e3, 32'h425b8256, 32'h42b0675f, 32'h4291747f, 32'hc281f40c, 32'h4235f0ed, 32'h4249380e};
test_bias[937:937] = '{32'h42aaf26e};
test_output[937:937] = '{32'h46d0136e};
test_input[7504:7511] = '{32'hc260b073, 32'hc25e73ec, 32'h420feeb2, 32'h426ddb5d, 32'h4279a267, 32'h4110c8c8, 32'hc181bdde, 32'h418ef347};
test_weights[7504:7511] = '{32'hc2c2f520, 32'hc2b2e657, 32'hc29e4185, 32'h40be0afc, 32'h423c4ec4, 32'h41d3a63e, 32'hc2549332, 32'h426e385a};
test_bias[938:938] = '{32'hc2209731};
test_output[938:938] = '{32'h464b6d8b};
test_input[7512:7519] = '{32'h420b9f33, 32'h41f01919, 32'hc1051a8e, 32'h3fa0e099, 32'hc25cd988, 32'hc285e2f3, 32'h42c394ef, 32'hc2948386};
test_weights[7512:7519] = '{32'hc2a8b4e9, 32'hc244022b, 32'h42912047, 32'h42854951, 32'hc24e68af, 32'hc2a77da0, 32'h4166890a, 32'hc2bdf8fe};
test_bias[939:939] = '{32'h42100f87};
test_output[939:939] = '{32'h463bcafa};
test_input[7520:7527] = '{32'hc1f3198d, 32'hc2c128de, 32'h4228abe7, 32'h4092d130, 32'h3e7c2cc6, 32'hc294adb9, 32'h423d6794, 32'h42b84a57};
test_weights[7520:7527] = '{32'h41b38972, 32'hc1977535, 32'h4193afbc, 32'hc254a25e, 32'hc2aea4b7, 32'hc10d202e, 32'hc0edbe65, 32'hc2bef154};
test_bias[940:940] = '{32'h421e866f};
test_output[940:940] = '{32'hc5d450fb};
test_input[7528:7535] = '{32'hc2a6ff17, 32'hc2ae3b7b, 32'h419eba7e, 32'h42487e64, 32'h407982e4, 32'h417fd8f8, 32'hc2934509, 32'hc28d6f48};
test_weights[7528:7535] = '{32'h422975fe, 32'hc25505a7, 32'hc2c21d46, 32'h4227d598, 32'hc1fb9c48, 32'hc0974ff0, 32'h4290a76c, 32'hc29eca74};
test_bias[941:941] = '{32'h41de7275};
test_output[941:941] = '{32'h44aeba03};
test_input[7536:7543] = '{32'h42868e70, 32'h41df12bb, 32'hc017a758, 32'h422f504a, 32'hc2b97fec, 32'h428bb3fb, 32'h417c4827, 32'hc25b7c9e};
test_weights[7536:7543] = '{32'h429fc076, 32'h41549bb1, 32'h4131b2d4, 32'hc2b6f918, 32'h418d6eec, 32'h41d2bc8a, 32'hc1c021f0, 32'hc2827a84};
test_bias[942:942] = '{32'hc2adbcf6};
test_output[942:942] = '{32'h459cf781};
test_input[7544:7551] = '{32'h42698670, 32'h42ba3d13, 32'h41351211, 32'hc2ad6cde, 32'hbfd87f2a, 32'h424cbbf5, 32'h42bd43c4, 32'h422e3b58};
test_weights[7544:7551] = '{32'hc2a2486e, 32'hc21f5f47, 32'hc294639c, 32'hc2241e1b, 32'h42351d7a, 32'hc25f69a6, 32'hc1ff8c32, 32'hc29555dd};
test_bias[943:943] = '{32'h4230c437};
test_output[943:943] = '{32'hc668be64};
test_input[7552:7559] = '{32'hc229d9e7, 32'h40462385, 32'h4289c23e, 32'h40e79b1f, 32'h41a897cf, 32'hc26282ec, 32'h41a674a3, 32'h41eb198e};
test_weights[7552:7559] = '{32'h42ae98d3, 32'h40cd980c, 32'hc2808fb7, 32'h41c63e3a, 32'hc208d3d2, 32'hc0f46a24, 32'h4297f4d3, 32'h41c894ce};
test_bias[944:944] = '{32'hc275fe2d};
test_output[944:944] = '{32'hc5ba7bc1};
test_input[7560:7567] = '{32'hc0c94de0, 32'hc264bf58, 32'h427e9718, 32'h40cc692e, 32'hc0015cc3, 32'hc1dd7820, 32'hc269311b, 32'h419aa80b};
test_weights[7560:7567] = '{32'h42b91109, 32'h42abac75, 32'h402a80de, 32'hc2725173, 32'hc22c0876, 32'h42b45ad8, 32'h41f6472b, 32'h417d039a};
test_bias[945:945] = '{32'hc2325557};
test_output[945:945] = '{32'hc616cd4e};
test_input[7568:7575] = '{32'hc2832e66, 32'hc2966fb7, 32'h4024538a, 32'h42aadb79, 32'hc2a2325a, 32'h4247697a, 32'h4201911f, 32'hc0389b5d};
test_weights[7568:7575] = '{32'h421b97f5, 32'hc0c7bd18, 32'hc1042feb, 32'h41c05f08, 32'h42b0bb0a, 32'h4279a03b, 32'hc244c8ae, 32'h41905fb7};
test_bias[946:946] = '{32'hc170511b};
test_output[946:946] = '{32'hc5b424a1};
test_input[7576:7583] = '{32'hc1d38678, 32'hc2906c25, 32'hc2993df3, 32'h425e0afd, 32'hc12355d4, 32'h42a26051, 32'hc2544237, 32'h42b02499};
test_weights[7576:7583] = '{32'hc24c0f62, 32'hc280e5d1, 32'hc1f1416f, 32'hc29f4631, 32'h4076a95f, 32'hc2860065, 32'hc1d40293, 32'h427b247c};
test_bias[947:947] = '{32'hc21bff07};
test_output[947:947] = '{32'h45a5f51b};
test_input[7584:7591] = '{32'h429beac5, 32'h421fc76b, 32'hc21afd9a, 32'h41827645, 32'h41e7e631, 32'h418017fd, 32'h42a982b2, 32'h41aa9ab3};
test_weights[7584:7591] = '{32'hc25971d6, 32'hc291ee24, 32'h42274bfd, 32'hc20821e1, 32'hc0b0a6e7, 32'hc23c4e70, 32'hc1e369d7, 32'hc29e8206};
test_bias[948:948] = '{32'h429517a5};
test_output[948:948] = '{32'hc65eeb1d};
test_input[7592:7599] = '{32'h41b5f65a, 32'hc28d2639, 32'hc2a23b43, 32'h4295c258, 32'hc2c659ef, 32'hc182a59b, 32'hc24afea4, 32'hc2c0a681};
test_weights[7592:7599] = '{32'h427dab50, 32'hc299a286, 32'h42a67a46, 32'h4299403d, 32'h42af6a53, 32'h40c16d43, 32'hc0ddc842, 32'h42953706};
test_bias[949:949] = '{32'h42b4fcaf};
test_output[949:949] = '{32'hc617701d};
test_input[7600:7607] = '{32'hc21d6e4c, 32'hc290808d, 32'hc2c29462, 32'hc2c54806, 32'hc1ac38c5, 32'hc2c42b21, 32'h428b0b10, 32'h4263988b};
test_weights[7600:7607] = '{32'h426b4dd9, 32'h41a69006, 32'hc2a244dd, 32'h42a307ee, 32'hc2995b3f, 32'hc2970725, 32'hc2ad4c30, 32'h42b0ec21};
test_bias[950:950] = '{32'hc2345d97};
test_output[950:950] = '{32'h457d6ffb};
test_input[7608:7615] = '{32'hc19a3574, 32'h42868bfc, 32'hc2a24e17, 32'hc2a57123, 32'h419ec4c4, 32'h42a4e5da, 32'h41d1c7e8, 32'hc28bd58c};
test_weights[7608:7615] = '{32'h4061f51b, 32'h40729378, 32'h40a9c89f, 32'h42b2711d, 32'h42c04884, 32'h4214618c, 32'h4243c3c1, 32'h42a15cfc};
test_bias[951:951] = '{32'h42142fb5};
test_output[951:951] = '{32'hc5da119b};
test_input[7616:7623] = '{32'hc2a21065, 32'h42922068, 32'hc2765047, 32'h42b17a24, 32'hc18b8bff, 32'hc22f4fa6, 32'hc20fe730, 32'h429c7141};
test_weights[7616:7623] = '{32'hc28f9798, 32'hc1ad51cb, 32'h42c6aca9, 32'hc22179f2, 32'hc23d0379, 32'h42b17f0e, 32'h42474fef, 32'h41ec53fc};
test_bias[952:952] = '{32'h42996769};
test_output[952:952] = '{32'hc5f7f7f7};
test_input[7624:7631] = '{32'hc20feb8a, 32'h420c4fe0, 32'hc26d4282, 32'h42a78cdb, 32'hc20e4484, 32'hc205b463, 32'hc2add49e, 32'hc2901122};
test_weights[7624:7631] = '{32'h42c7460b, 32'h42adb6bc, 32'h4281f505, 32'h41ca889f, 32'hc22e7ddd, 32'h423954a9, 32'hc21fb51d, 32'hc2838b6e};
test_bias[953:953] = '{32'h422b8623};
test_output[953:953] = '{32'h45baf25e};
test_input[7632:7639] = '{32'h4288159f, 32'h41b8d543, 32'h421a3d39, 32'hc2a8e31c, 32'h4227a161, 32'hc2c25afa, 32'h414b6a68, 32'hc2330eda};
test_weights[7632:7639] = '{32'hc1092c9e, 32'hc26f9489, 32'h404aa42f, 32'h40b82f6a, 32'hc2b9788f, 32'h42b4d54b, 32'h42b029bd, 32'hc2b7fd54};
test_bias[954:954] = '{32'h42b1a6a5};
test_output[954:954] = '{32'hc61734b0};
test_input[7640:7647] = '{32'hc2a8623b, 32'hc2c50dfc, 32'h4152efec, 32'h420648c8, 32'h422650fc, 32'hc293accd, 32'h41d88c95, 32'h42b8ca9a};
test_weights[7640:7647] = '{32'h4211a2db, 32'h42883a72, 32'hc18233bc, 32'h4064bee3, 32'hc2337f80, 32'hc283678e, 32'h41ef37a1, 32'hc2902cf5};
test_bias[955:955] = '{32'h42a6129f};
test_output[955:955] = '{32'hc645b6f0};
test_input[7648:7655] = '{32'h41f9b8bb, 32'h42840ba4, 32'h4235d5b0, 32'hc2a0df38, 32'h42091878, 32'h42961b05, 32'h423d78e7, 32'hc18ea8c5};
test_weights[7648:7655] = '{32'h426dbaea, 32'hc2c37f59, 32'hc2c2bc1a, 32'h4269df06, 32'hc13affdc, 32'hc14bc280, 32'h3e5b7935, 32'hc213d309};
test_bias[956:956] = '{32'hc2aeca09};
test_output[956:956] = '{32'hc6629893};
test_input[7656:7663] = '{32'h427903e7, 32'h422d9dfb, 32'h42aa50ab, 32'hc2668e55, 32'h415a6217, 32'h4184387c, 32'hc26b61b2, 32'h42b8123a};
test_weights[7656:7663] = '{32'hc27bddc3, 32'hc2846ebf, 32'hc150c06f, 32'hc1aeb1a4, 32'hc2114993, 32'hc2370486, 32'h422269d2, 32'hc263eec9};
test_bias[957:957] = '{32'h428b1dd5};
test_output[957:957] = '{32'hc6719a5b};
test_input[7664:7671] = '{32'h4200675f, 32'h41f08e8a, 32'h42c3c403, 32'hc299ff79, 32'hc2972742, 32'hc2a7e06d, 32'h428f3960, 32'hc241f40b};
test_weights[7664:7671] = '{32'h429e0c9d, 32'h4292968e, 32'h420e13f7, 32'h4231d344, 32'h415ff179, 32'h4211fa11, 32'hbe2f9797, 32'h42893a2b};
test_bias[958:958] = '{32'h4292c8b2};
test_output[958:958] = '{32'hc5220916};
test_input[7672:7679] = '{32'h42be2714, 32'hc2b59b74, 32'hc2859805, 32'hc2816a93, 32'h426ca87d, 32'h3eaf77a8, 32'hc2b24f77, 32'hc240a15f};
test_weights[7672:7679] = '{32'hc286c9cd, 32'h4204a8d2, 32'h42c5a21c, 32'h42852898, 32'hc295155a, 32'hc2acae5e, 32'hc22bc849, 32'h4270f32e};
test_bias[959:959] = '{32'h404d7f23};
test_output[959:959] = '{32'hc6ba393c};
test_input[7680:7687] = '{32'hbfc60263, 32'h42a3858c, 32'hc2c105a4, 32'hc1a95e94, 32'hc2097b5a, 32'hc20610c4, 32'h42428cc1, 32'h41c90ebf};
test_weights[7680:7687] = '{32'hc28c46ec, 32'h42ba462f, 32'h426ef567, 32'h421532f4, 32'h3fc58bbf, 32'hc2a4d28b, 32'h41e9ead0, 32'h41b06cd5};
test_bias[960:960] = '{32'h42adf22a};
test_output[960:960] = '{32'h45b9a587};
test_input[7688:7695] = '{32'hc089effc, 32'hc23b561f, 32'h42976a58, 32'hc287fced, 32'hc235e48a, 32'h4173a426, 32'h422b08d3, 32'hc210bb5c};
test_weights[7688:7695] = '{32'hc0267865, 32'h41d8b8de, 32'hc23871f6, 32'h4161453e, 32'hc28e2d52, 32'hc2b7fb21, 32'h429f0f80, 32'hc1ff05a3};
test_bias[961:961] = '{32'hc291a82a};
test_output[961:961] = '{32'h4417cd37};
test_input[7696:7703] = '{32'hc138edf5, 32'hc2382823, 32'h427323e7, 32'hc1afb005, 32'h427f8dc6, 32'hc22e1f14, 32'h42be7d76, 32'h42bc58f0};
test_weights[7696:7703] = '{32'h42ab06de, 32'hc2b339b3, 32'h41fd14db, 32'hc2c0343b, 32'h42b42109, 32'hc2c63e8c, 32'h41e28d56, 32'h42b7cc5a};
test_bias[962:962] = '{32'h423e2353};
test_output[962:962] = '{32'h46dfbddb};
test_input[7704:7711] = '{32'hc27f7c64, 32'h41d0a12a, 32'hc2a1f831, 32'h423c9c55, 32'h4205a304, 32'h42739501, 32'hc1e11d21, 32'hc226a256};
test_weights[7704:7711] = '{32'h41daca1f, 32'hc22fa94f, 32'hc2027e12, 32'h4239a453, 32'h4102a8a7, 32'hc173b869, 32'hc1d465b1, 32'hc28c548b};
test_bias[963:963] = '{32'hc1099e6d};
test_output[963:963] = '{32'h459a87ed};
test_input[7712:7719] = '{32'h42091352, 32'h429ceb16, 32'h41694ab4, 32'h41fc9f3f, 32'h4295c4b9, 32'hc2b61372, 32'h412f67d1, 32'h4288e61c};
test_weights[7712:7719] = '{32'hc26efb26, 32'h41507243, 32'hc20b37d7, 32'hc281c866, 32'hc2bbe34a, 32'h40ba4ce1, 32'hc20c051a, 32'hc2ae89b9};
test_bias[964:964] = '{32'h415dacbc};
test_output[964:964] = '{32'hc688a460};
test_input[7720:7727] = '{32'hc242f25d, 32'hc274c7fe, 32'h4107fe7a, 32'hbff5b294, 32'h42252341, 32'h4257c2e7, 32'hc28ccc31, 32'h422996e9};
test_weights[7720:7727] = '{32'hc2241934, 32'hc297ff8d, 32'hc287562b, 32'h4206fdf4, 32'h42ae12d9, 32'hc2c5d133, 32'h42a9d231, 32'hc2402aca};
test_bias[965:965] = '{32'hc0d2eb19};
test_output[965:965] = '{32'hc56a8ad3};
test_input[7728:7735] = '{32'hc2b6e433, 32'hc23d5921, 32'h428d141e, 32'h41f4c25c, 32'hc1fd4a21, 32'h4214d90d, 32'hc2182229, 32'hc29fecdc};
test_weights[7728:7735] = '{32'hc238f3c9, 32'hc0efac25, 32'h428373ab, 32'h42bf361e, 32'hc26746e5, 32'h42a29cd9, 32'hc2912d1f, 32'h418094af};
test_bias[966:966] = '{32'hc2150a84};
test_output[966:966] = '{32'h46900d3d};
test_input[7736:7743] = '{32'h3f9dcd08, 32'hc27c3bcc, 32'h4235b4f8, 32'h41fe5bd6, 32'hc1894f00, 32'hc25a5a05, 32'hc2366085, 32'hc14f2a93};
test_weights[7736:7743] = '{32'hc29a8eb1, 32'hc2c543ec, 32'h429d9e6f, 32'h4233eb79, 32'hc25b48f1, 32'hc1d215f1, 32'h419f222e, 32'hc2ba76fc};
test_bias[967:967] = '{32'hc0931ff5};
test_output[967:967] = '{32'h4657b263};
test_input[7744:7751] = '{32'hc2212209, 32'h421734d1, 32'h4296f73d, 32'h420c7dbd, 32'hc11e0a88, 32'h41f556b1, 32'h41b35806, 32'hc2c4416e};
test_weights[7744:7751] = '{32'h426a5f71, 32'hc0b65ea2, 32'h42979f24, 32'hc2c65961, 32'hc13efe26, 32'hc294a5ea, 32'hc12a65dd, 32'h42be2813};
test_bias[968:968] = '{32'h4238fd0b};
test_output[968:968] = '{32'hc63bd16f};
test_input[7752:7759] = '{32'hc1ac255f, 32'h411cc9e6, 32'hc2899dcd, 32'hc23ff0f4, 32'hc234d0c0, 32'h41c51cec, 32'hc0eaecca, 32'h425e4905};
test_weights[7752:7759] = '{32'h425d0a6c, 32'h413b5f4d, 32'h421030e8, 32'h4208619c, 32'h412fe43e, 32'hc239dcb2, 32'hc20d7c18, 32'hc181d795};
test_bias[969:969] = '{32'hc20d74ec};
test_output[969:969] = '{32'hc5eab1df};
test_input[7760:7767] = '{32'h422ddd6e, 32'h425341c7, 32'hc2349247, 32'h42bd9662, 32'hc290683b, 32'hc171ded1, 32'h42b8983e, 32'hc181d83e};
test_weights[7760:7767] = '{32'h421d4062, 32'hc1b027d2, 32'h40447596, 32'hc1e8d215, 32'h42c45690, 32'hc18b6839, 32'hc2a15434, 32'h42a0753c};
test_bias[970:970] = '{32'h4212e4da};
test_output[970:970] = '{32'hc68bbd85};
test_input[7768:7775] = '{32'hc2bb7740, 32'hc20b429e, 32'hc28053c7, 32'hc2bd09b5, 32'h42bbff23, 32'h4236e882, 32'hc267551d, 32'h42a3a305};
test_weights[7768:7775] = '{32'h4228699c, 32'h41818907, 32'h42b7aa92, 32'h4175b7cc, 32'hc25c3399, 32'hc22f892c, 32'h42a271b5, 32'hc2ae9725};
test_bias[971:971] = '{32'h4184d5a6};
test_output[971:971] = '{32'hc6f114f9};
test_input[7776:7783] = '{32'hc270b6b6, 32'hc1b19026, 32'hc0904094, 32'hc229279b, 32'hc1a0828c, 32'hc2af5a1e, 32'hc1e1ce19, 32'hc286823b};
test_weights[7776:7783] = '{32'hc29ebadc, 32'hc1f318b3, 32'hc2a21ca3, 32'h426b00a2, 32'h426b04a0, 32'hc0820bc4, 32'hc26d2597, 32'h4216044c};
test_bias[972:972] = '{32'hc082a766};
test_output[972:972] = '{32'h44cefc87};
test_input[7784:7791] = '{32'hc19a769d, 32'hc180297b, 32'h42c4be69, 32'hc1cbbe17, 32'h42a1fdc3, 32'hc1443d76, 32'h3e1ccd72, 32'h417edc39};
test_weights[7784:7791] = '{32'hc1d302f3, 32'h4290d60d, 32'h42389559, 32'hc298f9bb, 32'hc2939d41, 32'h428d16d0, 32'h4203746b, 32'hc0be7db4};
test_bias[973:973] = '{32'hc2422c89};
test_output[973:973] = '{32'hc48f2236};
test_input[7792:7799] = '{32'h429980b8, 32'hc2adcf67, 32'h41ff9b3c, 32'hc1edc040, 32'hc11bcdbc, 32'hc2b74dbd, 32'hc2a1cb15, 32'hc2b2ac52};
test_weights[7792:7799] = '{32'h42625d86, 32'hc19846ae, 32'hc24d0563, 32'h41666549, 32'hc20e2c3b, 32'h41a11ad7, 32'h4226c5d1, 32'hc222b1cc};
test_bias[974:974] = '{32'h41570c91};
test_output[974:974] = '{32'h45292bae};
test_input[7800:7807] = '{32'h4268f2e7, 32'hc291dcb7, 32'h4211c454, 32'hc296009a, 32'hc299a507, 32'hc11bfd2c, 32'hc2302072, 32'hc28d4f81};
test_weights[7800:7807] = '{32'h42a09430, 32'h42832209, 32'h42a5c4fc, 32'hc2c1f0bf, 32'hc28cc48f, 32'h42b5e11f, 32'hc2415b9f, 32'hc2b51176};
test_bias[975:975] = '{32'h41a74f02};
test_output[975:975] = '{32'h46b5abc8};
test_input[7808:7815] = '{32'hc2b071eb, 32'hc1ce3945, 32'hbe389030, 32'h41912a30, 32'h42300e9b, 32'h41c4af6e, 32'h4269bd1a, 32'hc2bb4fd9};
test_weights[7808:7815] = '{32'hc2a33fea, 32'hc27fa3db, 32'hc1fa8b45, 32'h42127621, 32'h4157e81e, 32'h428e2af9, 32'hc192620d, 32'hc1b759e1};
test_bias[976:976] = '{32'h4211a0e1};
test_output[976:976] = '{32'h464ab7ab};
test_input[7816:7823] = '{32'h4193ffc3, 32'h42aaf95c, 32'h421410b7, 32'hc22ec673, 32'hc1f6b41e, 32'hc1ad2ae5, 32'hc27cd72b, 32'h42a1a558};
test_weights[7816:7823] = '{32'hc0a1aa51, 32'hc2975b0d, 32'hc2c3bd04, 32'h4287c3e3, 32'hc2c13397, 32'h4255e97e, 32'h424bed9e, 32'hc211e75d};
test_bias[977:977] = '{32'h405876fe};
test_output[977:977] = '{32'hc688b34b};
test_input[7824:7831] = '{32'h41a7332a, 32'hc289f10e, 32'hc1a097c3, 32'hc2c15a40, 32'h429fa7fa, 32'hc297a1b9, 32'h42a73e11, 32'h429c007b};
test_weights[7824:7831] = '{32'h42a24368, 32'h42601e61, 32'hc2afa1dd, 32'hc28670d1, 32'hc2ac51b8, 32'h40daf54a, 32'h423f1081, 32'h42846d5c};
test_bias[978:978] = '{32'h41b56b1b};
test_output[978:978] = '{32'h45f62cf5};
test_input[7832:7839] = '{32'hc28e29c0, 32'hc18db37d, 32'hc16845de, 32'hc2c494f2, 32'hc1cfde7b, 32'hc2375a25, 32'hc12cb791, 32'h4280d621};
test_weights[7832:7839] = '{32'h4282e1de, 32'hc2afea8b, 32'h4191290f, 32'hc286acbb, 32'hc2829451, 32'h41a105dd, 32'h402dcb1d, 32'hc05edc01};
test_bias[979:979] = '{32'hc1da0763};
test_output[979:979] = '{32'h456aa826};
test_input[7840:7847] = '{32'hc19b5fa4, 32'hc293d997, 32'h42a9df28, 32'h415c3ffa, 32'hc2027066, 32'hc16b045c, 32'h41d5a2db, 32'h41866457};
test_weights[7840:7847] = '{32'hc28111f3, 32'h42a34fa2, 32'hc281e275, 32'hc2ab30f0, 32'h42033ab1, 32'hc2bb4841, 32'hc16a67c1, 32'hc09c4029};
test_bias[980:980] = '{32'h4277116f};
test_output[980:980] = '{32'hc634fc56};
test_input[7848:7855] = '{32'h42c6940b, 32'hc29ad819, 32'hc1f3e232, 32'h401ed888, 32'h42351092, 32'h41d8798b, 32'hc23b3543, 32'h428499d7};
test_weights[7848:7855] = '{32'h4118f882, 32'hc29b426e, 32'hc187881d, 32'h41a1d556, 32'h41f8f2f6, 32'hc2470ca4, 32'hc1cd0dd9, 32'h42108cd2};
test_bias[981:981] = '{32'hc266630f};
test_output[981:981] = '{32'h462dd8f9};
test_input[7856:7863] = '{32'hc2219ee4, 32'hc216fe7c, 32'hc2b95dae, 32'h42873cec, 32'hc2a3695c, 32'hc1fb24c8, 32'hc21b6092, 32'h41ce8a1c};
test_weights[7856:7863] = '{32'hc16723de, 32'hc1a7340d, 32'hc147fe2c, 32'hc230dc6a, 32'h41b167e2, 32'h429d3b57, 32'h422b8493, 32'hc2363bbc};
test_bias[982:982] = '{32'h4235e052};
test_output[982:982] = '{32'hc5eb76d9};
test_input[7864:7871] = '{32'h4207051f, 32'hc25d7adf, 32'h42a9c7d8, 32'hc2869937, 32'hc2984d0d, 32'h429721dd, 32'h41acb122, 32'hc29b452c};
test_weights[7864:7871] = '{32'hc2732918, 32'hc26b872a, 32'h422ea601, 32'hc1ab5950, 32'h426e5a11, 32'h42c3402d, 32'hc12da0a1, 32'h41694293};
test_bias[983:983] = '{32'hc1af48b7};
test_output[983:983] = '{32'h45f3fe74};
test_input[7872:7879] = '{32'hc2b0147d, 32'h429b2ac2, 32'h4283bd17, 32'h42835bb0, 32'h41cd4100, 32'hc22db91d, 32'hc114d47a, 32'hc285b4c0};
test_weights[7872:7879] = '{32'hc2ac337d, 32'h42ba960b, 32'hc256e9cc, 32'h4225a7ed, 32'hc1fd8f06, 32'h42a02cd5, 32'h424ba7d6, 32'hc2b071d0};
test_bias[984:984] = '{32'hc2923e67};
test_output[984:984] = '{32'h466b4c2b};
test_input[7880:7887] = '{32'h421bbb22, 32'h426d95fc, 32'h42ac9357, 32'hc233f9f9, 32'h42bedc4f, 32'hbd4086ba, 32'hc258ee92, 32'h42a83b4d};
test_weights[7880:7887] = '{32'hc00ffe4c, 32'h3e6b8e0d, 32'h426a2378, 32'h4284f55d, 32'hc29d3286, 32'hc2c5e1de, 32'hc1caf53e, 32'h428eadac};
test_bias[985:985] = '{32'hc29cbea5};
test_output[985:985] = '{32'h44df7de9};
test_input[7888:7895] = '{32'h41c88d1d, 32'h4200be95, 32'h41ae5037, 32'h401c1bc3, 32'hc2898b4e, 32'h425acd5f, 32'h422c9d40, 32'hc1de0e68};
test_weights[7888:7895] = '{32'hc1f0b25c, 32'h41d10d6c, 32'hc18d10cd, 32'h41eddd88, 32'h42a39a36, 32'h40a6c113, 32'hc2c7ca1f, 32'hc21c1763};
test_bias[986:986] = '{32'hc2a5cc6f};
test_output[986:986] = '{32'hc60ab00c};
test_input[7896:7903] = '{32'hc12699b7, 32'hc0e9d9ad, 32'h42990e8c, 32'hc1e5d49b, 32'hc2bfd977, 32'h420a7d4b, 32'h424bd42c, 32'h423336e6};
test_weights[7896:7903] = '{32'h4284e97e, 32'hc1738d9a, 32'h42113cb1, 32'h41fd10e1, 32'hc21d8349, 32'h412a7af7, 32'hc2501ace, 32'hc14b63ed};
test_bias[987:987] = '{32'hc2260bbf};
test_output[987:987] = '{32'h4507d41f};
test_input[7904:7911] = '{32'hc298e477, 32'hc24db648, 32'hc1a67d4f, 32'hc2961c1d, 32'h41d70abc, 32'h4136bb96, 32'hc202721d, 32'h425455f6};
test_weights[7904:7911] = '{32'h4281f302, 32'hc1c05468, 32'h4200cba8, 32'hc270e07b, 32'h429e1088, 32'hbfc1d28b, 32'h416e5f0b, 32'hc2a511ff};
test_bias[988:988] = '{32'h429e1a61};
test_output[988:988] = '{32'hc5202004};
test_input[7912:7919] = '{32'h42684011, 32'hc2756b60, 32'hc25976c5, 32'hc29aabc1, 32'h429ec683, 32'hc2bf4300, 32'hc2c3ceec, 32'hc26e91aa};
test_weights[7912:7919] = '{32'h417134b9, 32'hc265e61e, 32'hc29b7475, 32'hc29373eb, 32'hc20c36d1, 32'hc29e5662, 32'h42475201, 32'h42ba88c9};
test_bias[989:989] = '{32'h420c8474};
test_output[989:989] = '{32'h46081c70};
test_input[7920:7927] = '{32'h42c14fb8, 32'h428a1931, 32'h42afafaf, 32'hc296b5aa, 32'hc1ce84f0, 32'h42c1fb64, 32'h41f95382, 32'h420379a4};
test_weights[7920:7927] = '{32'hc205a443, 32'h42c0794d, 32'h414787be, 32'h4185beab, 32'h4217a3e2, 32'h42ada162, 32'hc26da111, 32'h4269d83b};
test_bias[990:990] = '{32'hc1fa21da};
test_output[990:990] = '{32'h4627af9b};
test_input[7928:7935] = '{32'hc20e81d3, 32'h4259e9f4, 32'hc07b9de3, 32'h42b949f7, 32'hc2b5447b, 32'h418fb6ab, 32'hc238f178, 32'hc1be4ca6};
test_weights[7928:7935] = '{32'hc2c76e08, 32'hc1c3d475, 32'hc1ba2521, 32'h42979ca4, 32'hc28f3d86, 32'h428042b3, 32'h42a8dfa8, 32'hc1bf04d6};
test_bias[991:991] = '{32'h42bf7c87};
test_output[991:991] = '{32'h4656a1a2};
test_input[7936:7943] = '{32'h4127c804, 32'h42c6f9f9, 32'h42594518, 32'hc20f171e, 32'hc2023fb4, 32'h4276838d, 32'hc28fefc9, 32'hc220e25b};
test_weights[7936:7943] = '{32'h3e1298ad, 32'h42697611, 32'hc26bb58b, 32'hc286a672, 32'hc2a03cf3, 32'h4063d369, 32'hc01c9148, 32'h426be0f8};
test_bias[992:992] = '{32'h41b1cf5d};
test_output[992:992] = '{32'h45b133c8};
test_input[7944:7951] = '{32'h42076f96, 32'h42a4a0ca, 32'hc1936e60, 32'hc12fba63, 32'h4212f1a4, 32'h42716446, 32'h428e06c8, 32'h42bc4813};
test_weights[7944:7951] = '{32'hc2863d66, 32'h426f19d3, 32'hc282b3f8, 32'h42b427c1, 32'hc1a51154, 32'hc2bb8ead, 32'h41dd6412, 32'hc284f61a};
test_bias[993:993] = '{32'h4277f928};
test_output[993:993] = '{32'hc5f34f52};
test_input[7952:7959] = '{32'hc0ec3d43, 32'h3f257300, 32'hc2afa55f, 32'hc2bb7d5d, 32'h41c95d79, 32'hc14b70e2, 32'hc2885b7d, 32'h423861fa};
test_weights[7952:7959] = '{32'hc1b2315a, 32'h4295d1c6, 32'h42c7600d, 32'hc2ba7ee0, 32'hc2888d3a, 32'hc1ef43be, 32'hc29d7948, 32'h404bc190};
test_bias[994:994] = '{32'hc284db46};
test_output[994:994] = '{32'h4586add4};
test_input[7960:7967] = '{32'hc2a95942, 32'h42bbc0d7, 32'hc26c0f34, 32'hc2c7beb4, 32'h4285dd34, 32'h425c43a6, 32'h4286c076, 32'h42869afb};
test_weights[7960:7967] = '{32'hc21e1b9a, 32'h42aae38c, 32'hc2bac678, 32'h42acd610, 32'h425084a9, 32'hc27b0580, 32'h41a95c34, 32'h42be4291};
test_bias[995:995] = '{32'hc0f59104};
test_output[995:995] = '{32'h467b9d00};
test_input[7968:7975] = '{32'hc11d2e44, 32'hc281a5ad, 32'hc23873e3, 32'hc2c6480b, 32'hc1abe6f6, 32'h428afd97, 32'h429ad15c, 32'hc2b65d49};
test_weights[7968:7975] = '{32'hc2c39202, 32'hc1f5b37c, 32'hc24a96e9, 32'hc2a5c605, 32'hc283b6fb, 32'hc20092c4, 32'hc1c8ca27, 32'h4251d464};
test_bias[996:996] = '{32'hc2a19b5f};
test_output[996:996] = '{32'h45b7b7a9};
test_input[7976:7983] = '{32'h4298bece, 32'h428a3c50, 32'hc1f67db1, 32'h42049ffa, 32'hc2090d13, 32'hc2add1db, 32'h4260e72f, 32'h42671144};
test_weights[7976:7983] = '{32'hc1df81ae, 32'hc2bdf00a, 32'h426aaaed, 32'h42aca4e1, 32'hc2603748, 32'h428db63f, 32'hc28562e6, 32'hc1dd525c};
test_bias[997:997] = '{32'h426abe9d};
test_output[997:997] = '{32'hc6862430};
test_input[7984:7991] = '{32'h3f9ca7e7, 32'h414bae60, 32'hc222609d, 32'h42572df9, 32'h424081c3, 32'h425a6861, 32'hc2b1280e, 32'h41c368e8};
test_weights[7984:7991] = '{32'hc187a867, 32'h40ec968a, 32'h429ab959, 32'h41f8e57f, 32'h420208f5, 32'h41421b36, 32'hc1bddb61, 32'hc1e8e987};
test_bias[998:998] = '{32'hc0c42bb3};
test_output[998:998] = '{32'h450aa65e};
test_input[7992:7999] = '{32'hc2a81ce9, 32'hc1fe8161, 32'hc0fc8674, 32'h42055b32, 32'hc1f20747, 32'hc296598f, 32'h422dec94, 32'h42a919e7};
test_weights[7992:7999] = '{32'h419997bc, 32'hc1e2ddfc, 32'hc2857b5d, 32'hc19eaa5a, 32'hc29954be, 32'h42b9c5f5, 32'h41b342f3, 32'h4208525d};
test_bias[999:999] = '{32'hc2a8fb6a};
test_output[999:999] = '{32'hc4d945b4};
test_input[8000:8007] = '{32'h42b8059b, 32'hc0da6aaf, 32'hc1ed2cee, 32'h428f4fcc, 32'h42a935a6, 32'hc2bc1c5f, 32'hbfd7de26, 32'h42b50064};
test_weights[8000:8007] = '{32'h420f0ac5, 32'hc28ecb98, 32'h426be276, 32'hc1df3e4b, 32'hc0f091f1, 32'hc0c30745, 32'h42821d27, 32'h425bd617};
test_bias[1000:1000] = '{32'h41337704};
test_output[1000:1000] = '{32'h45975282};
test_input[8008:8015] = '{32'h40cae321, 32'hc2b551a7, 32'h40f09a86, 32'hc0e51cb0, 32'hc260ccff, 32'h41359048, 32'hc221483a, 32'h42710ff6};
test_weights[8008:8015] = '{32'hc2c519d7, 32'hc206235a, 32'h41a54b5a, 32'hc13f9d05, 32'hc2a211a9, 32'hc17d1e0a, 32'h42b6ce52, 32'h427ebe10};
test_bias[1001:1001] = '{32'hc253c761};
test_output[1001:1001] = '{32'h45ded67e};
test_input[8016:8023] = '{32'hc2c0d16d, 32'hc19ed761, 32'hc269ffc3, 32'hc2ab2c35, 32'hc10f50b2, 32'hc0e843e2, 32'hc0fb765e, 32'hc27899e7};
test_weights[8016:8023] = '{32'hc215f743, 32'h4266ec49, 32'h4287a11b, 32'hbfd14e8c, 32'hc17475f9, 32'h41d2623d, 32'hc2bc2767, 32'h426a4f09};
test_bias[1002:1002] = '{32'hc12ce796};
test_output[1002:1002] = '{32'hc5872892};
test_input[8024:8031] = '{32'hc18d97e0, 32'h422c5cbf, 32'h429f5c01, 32'h4287d121, 32'hc1f87097, 32'h428ac4e1, 32'h42bbc2eb, 32'h42a91d18};
test_weights[8024:8031] = '{32'hc22eaf7b, 32'hc234e550, 32'hc189a55f, 32'hc2596b4e, 32'hc1b7f848, 32'h421d60cf, 32'h415fb5a2, 32'h40d11e11};
test_bias[1003:1003] = '{32'hc2c22fbe};
test_output[1003:1003] = '{32'hc4803726};
test_input[8032:8039] = '{32'hc2bc61e8, 32'h425b1c6a, 32'h42a8bf4d, 32'hc2c3f500, 32'h415a75e0, 32'h4278bcfe, 32'hc05945c7, 32'h421282bc};
test_weights[8032:8039] = '{32'hc2b5734e, 32'hc152aefb, 32'hc269ad77, 32'h42335130, 32'hc2ac4050, 32'h3fc295d4, 32'hc2ae22b0, 32'hc20371e7};
test_bias[1004:1004] = '{32'h4294f4da};
test_output[1004:1004] = '{32'hc55541e4};
test_input[8040:8047] = '{32'h41829719, 32'h3f47f92d, 32'h4233ce7d, 32'h41f85c86, 32'h4282cb02, 32'h42972809, 32'h41e933b7, 32'h4239f748};
test_weights[8040:8047] = '{32'h3f93f790, 32'hc2a88739, 32'hc2c630b3, 32'hc13c5c41, 32'h405517cc, 32'h42c79971, 32'h42c49676, 32'hc20693c5};
test_bias[1005:1005] = '{32'hbfa8d819};
test_output[1005:1005] = '{32'h45830a67};
test_input[8048:8055] = '{32'hc255e6a0, 32'hc27e66e5, 32'hc2ab3c73, 32'hc1baa482, 32'h42a53dc4, 32'hc1b60e62, 32'hc2634c1d, 32'h422a61f3};
test_weights[8048:8055] = '{32'hc2657906, 32'hc1ee8229, 32'h42584119, 32'h40645675, 32'hc2c195df, 32'h421f55cd, 32'hc2acacc6, 32'h42affaaf};
test_bias[1006:1006] = '{32'h41e5566f};
test_output[1006:1006] = '{32'h41f8191e};
test_input[8056:8063] = '{32'h410227ac, 32'h42c27fde, 32'h42446cfc, 32'h41233c7f, 32'h428e6b04, 32'hc2c6cbe0, 32'h4214f4e7, 32'h41ed9536};
test_weights[8056:8063] = '{32'hc289dc73, 32'hc291d0a4, 32'hc2a97047, 32'hc193e514, 32'hc291160b, 32'hc0ac4bb1, 32'hc2770a48, 32'hc1758451};
test_bias[1007:1007] = '{32'h42c19e7a};
test_output[1007:1007] = '{32'hc696b252};
test_input[8064:8071] = '{32'hc1db92eb, 32'hc287732b, 32'h42a862ae, 32'hc2ad5d70, 32'h427097c6, 32'hc20905d0, 32'hc258d659, 32'hc28b2123};
test_weights[8064:8071] = '{32'h424d824d, 32'h42b77333, 32'hc178d9a4, 32'h425361f3, 32'hc2a6f10e, 32'h42335425, 32'h422f1e82, 32'hc2be72d3};
test_bias[1008:1008] = '{32'hbe9611b8};
test_output[1008:1008] = '{32'hc677289f};
test_input[8072:8079] = '{32'hc1840bf1, 32'hc201a0c3, 32'h427dd591, 32'h40f0066f, 32'h4159fc2a, 32'h41a8a284, 32'hc1c3d95b, 32'hc25315f6};
test_weights[8072:8079] = '{32'h4102d83a, 32'hc276c24a, 32'h428c607e, 32'h42bcf0a9, 32'hc1b1527d, 32'hc23af010, 32'hc1d9f1cb, 32'hc249c638};
test_bias[1009:1009] = '{32'h429992b9};
test_output[1009:1009] = '{32'h460ee5ce};
test_input[8080:8087] = '{32'h425b4101, 32'hc296413f, 32'hc21fa4de, 32'h41a6fa3f, 32'h42a08a43, 32'hc23971ea, 32'h412dccb5, 32'h42a7c5c8};
test_weights[8080:8087] = '{32'hc1fcfeaa, 32'h420c08f0, 32'h4281c7b2, 32'h42aa2b4c, 32'h3fbb1596, 32'hc2558d61, 32'h42bfb35f, 32'h42c28664};
test_bias[1010:1010] = '{32'hc2af69df};
test_output[1010:1010] = '{32'h45cbfb76};
test_input[8088:8095] = '{32'hc240e85b, 32'hc28d47bf, 32'hc29f2e42, 32'hc2594667, 32'hc2539f98, 32'hc280cc41, 32'h42565c05, 32'h42866214};
test_weights[8088:8095] = '{32'h4102c51f, 32'hc2bb6aa9, 32'h418db15d, 32'h423b090a, 32'hc26e742d, 32'hc220985a, 32'hc2a69cf9, 32'h4225b07d};
test_bias[1011:1011] = '{32'hc2196e94};
test_output[1011:1011] = '{32'h45c4be31};
test_input[8096:8103] = '{32'hc0a8147d, 32'hc2bed5f5, 32'hc28b0ca9, 32'hc1d68e83, 32'h42a0d8c2, 32'hc244e61d, 32'hc2bda9c4, 32'h4265d28b};
test_weights[8096:8103] = '{32'h42bec722, 32'hc29a397c, 32'h3fc3d424, 32'h4143adcb, 32'hc29dd903, 32'h410e5476, 32'hc2914a45, 32'hc2817d40};
test_bias[1012:1012] = '{32'hc11741ad};
test_output[1012:1012] = '{32'h452ecefb};
test_input[8104:8111] = '{32'h42c06675, 32'h41b52e3a, 32'h42b92894, 32'h42658f2c, 32'hc2671b67, 32'h41feaeff, 32'hc2bfca7a, 32'hc28bc5e0};
test_weights[8104:8111] = '{32'hc1cd89fd, 32'hc186ebbb, 32'h41abb9ed, 32'h428ae4d1, 32'hc260de91, 32'hc26062d6, 32'h413bce3e, 32'h4288415a};
test_bias[1013:1013] = '{32'hc290f6cc};
test_output[1013:1013] = '{32'hc4ac3a51};
test_input[8112:8119] = '{32'hc2bece39, 32'hc121b41d, 32'hc250cdae, 32'h42870cfd, 32'h418269ea, 32'h409f6792, 32'hc269698e, 32'h42805374};
test_weights[8112:8119] = '{32'hc07ab7e5, 32'hc2968827, 32'hc269ce51, 32'hc111d9ba, 32'h40dffb32, 32'h42495587, 32'h4187acdf, 32'hc1b1f057};
test_bias[1014:1014] = '{32'hc2ac0733};
test_output[1014:1014] = '{32'h44b3047b};
test_input[8120:8127] = '{32'h42245477, 32'hc23a384b, 32'hc2773e89, 32'hc2ac1bea, 32'hc2ae8641, 32'hc28eccfc, 32'hc29db7ce, 32'h4238d1b5};
test_weights[8120:8127] = '{32'hc2aca538, 32'h42631d89, 32'h42b64c50, 32'h42a787bd, 32'hc21f6c9e, 32'hc25746d2, 32'h4202bc62, 32'h42b2d503};
test_bias[1015:1015] = '{32'hc23bb5d6};
test_output[1015:1015] = '{32'hc61f715e};
test_input[8128:8135] = '{32'hc129c878, 32'h4214d0b8, 32'hbf97a109, 32'h42436edc, 32'hc10be42c, 32'h421c2620, 32'hc1b16683, 32'h41b3ac6c};
test_weights[8128:8135] = '{32'hc2c51ac8, 32'h42418433, 32'hc2ae6159, 32'h42b10726, 32'hc190c27e, 32'h41357502, 32'hc2b35a77, 32'h42197035};
test_bias[1016:1016] = '{32'hc2aa52bd};
test_output[1016:1016] = '{32'h46263de6};
test_input[8136:8143] = '{32'hc28cc0f9, 32'hc132df84, 32'hc2b585e8, 32'h42b6c240, 32'hc21ecb39, 32'h42c71a70, 32'hc0b42990, 32'hc24e3345};
test_weights[8136:8143] = '{32'h42201732, 32'hc29902f2, 32'hc29d64ea, 32'h428f2bd9, 32'h429b77f0, 32'hc233caa7, 32'hc29b15bf, 32'h41e040c6};
test_bias[1017:1017] = '{32'h425ccbf7};
test_output[1017:1017] = '{32'h45488ec1};
test_input[8144:8151] = '{32'h4273d0a6, 32'h4218e0b5, 32'h417e4f50, 32'hc1e9ace9, 32'h422ad11d, 32'h42a4394d, 32'h4286564f, 32'h426e0662};
test_weights[8144:8151] = '{32'h422fd150, 32'hc23856e7, 32'h41b9b778, 32'hc25e9b4e, 32'h419e3f40, 32'hc20ca908, 32'h41f5ce98, 32'hc2a5f39b};
test_bias[1018:1018] = '{32'h42b777cf};
test_output[1018:1018] = '{32'hc4ef0c82};
test_input[8152:8159] = '{32'h42798d69, 32'hc29e5824, 32'h41adada8, 32'hc179e327, 32'hc2918d78, 32'h421af7e8, 32'hc19e175c, 32'h4292ea1f};
test_weights[8152:8159] = '{32'h414a86d4, 32'h428965c0, 32'hc10f9f4a, 32'hc1cd03f5, 32'h41b49202, 32'h424306cc, 32'h419e6f03, 32'h40df77f8};
test_bias[1019:1019] = '{32'h421bf4d5};
test_output[1019:1019] = '{32'hc57c5115};
test_input[8160:8167] = '{32'h424229bc, 32'hc26c842d, 32'h42b6138d, 32'hc192e748, 32'hc18c7726, 32'hc29c1259, 32'hc21d4282, 32'hbf6ef92f};
test_weights[8160:8167] = '{32'hc18c3d72, 32'h4133c0df, 32'h422ba80e, 32'h42b93e5d, 32'h4214b94f, 32'h422df331, 32'hc1de0c24, 32'h3f5e7b6a};
test_bias[1020:1020] = '{32'h4189076d};
test_output[1020:1020] = '{32'hc50c8113};
test_input[8168:8175] = '{32'hc1247d21, 32'hc2aaf48c, 32'h424267b3, 32'hc25f2486, 32'h41231f2b, 32'h4253762a, 32'h42a6558d, 32'hc236af4d};
test_weights[8168:8175] = '{32'hc1f5ee15, 32'hc26fc4b8, 32'h419c4369, 32'h42875083, 32'hc2a7b54f, 32'h42aef25b, 32'h41ac6990, 32'h424355b0};
test_bias[1021:1021] = '{32'h40fd970c};
test_output[1021:1021] = '{32'h45ba1184};
test_input[8176:8183] = '{32'h41bef793, 32'h424704ee, 32'h42a5bf94, 32'h429b681b, 32'hc072f277, 32'hc2186e5a, 32'h42a720c6, 32'h4245ddb9};
test_weights[8176:8183] = '{32'hc2839ec9, 32'h4037e3a9, 32'h412de555, 32'hc2bf715a, 32'h40fae33c, 32'h41b033d6, 32'hc29698fa, 32'h42a2c15a};
test_bias[1022:1022] = '{32'h42453ddb};
test_output[1022:1022] = '{32'hc62caee8};
test_input[8184:8191] = '{32'h42ae3570, 32'hc137e8b9, 32'hc23529ce, 32'h426dd373, 32'hc258da9a, 32'hc262c157, 32'hc0ba2d37, 32'hc2919c22};
test_weights[8184:8191] = '{32'hc25be468, 32'hc10c93af, 32'hc06621b8, 32'hc29a6acb, 32'h422c6475, 32'hc27c2d79, 32'hc28b91e3, 32'hc1dab9bf};
test_bias[1023:1023] = '{32'hc1bbb153};
test_output[1023:1023] = '{32'hc5ac04c7};
test_input[8192:8199] = '{32'hc2a38e4a, 32'h42ad61f0, 32'h42a73ae1, 32'hbe449f71, 32'h42253b6a, 32'hc27377c2, 32'hc1049c23, 32'hc29d946a};
test_weights[8192:8199] = '{32'h4226a67b, 32'h420046a6, 32'hc1f1da9f, 32'hc0f6b896, 32'h4189bf2d, 32'h427f0447, 32'h4229262d, 32'hc29c81ad};
test_bias[1024:1024] = '{32'hc2bd41d2};
test_output[1024:1024] = '{32'hc41688aa};
test_input[8200:8207] = '{32'hc2038381, 32'h429c6c2d, 32'hc17709ca, 32'hc25d934e, 32'h4281a60b, 32'hc2aefebf, 32'h42401789, 32'hc1a9397a};
test_weights[8200:8207] = '{32'h429c4944, 32'hc2a1ab43, 32'hc1ded289, 32'h421c84fd, 32'hc2b19159, 32'hc2133c76, 32'hc2bf922e, 32'hc21ea666};
test_bias[1025:1025] = '{32'h4190ee83};
test_output[1025:1025] = '{32'hc68414b8};
test_input[8208:8215] = '{32'hc2877e96, 32'hc296e5e1, 32'h419dff56, 32'hc289925a, 32'h42a7d050, 32'hc1be17f9, 32'hc281072d, 32'hc28cbc9e};
test_weights[8208:8215] = '{32'hc28b7d03, 32'h4231ed9b, 32'hc25ca475, 32'hc2094c8b, 32'hc2a39cd9, 32'h4285f413, 32'h41e14a05, 32'hc27c2a68};
test_bias[1026:1026] = '{32'h42855f4d};
test_output[1026:1026] = '{32'hc5439120};
test_input[8216:8223] = '{32'hc29271db, 32'h41ad1476, 32'h4147b6e0, 32'hc278b3a2, 32'h4251f7f3, 32'h428c3d03, 32'hc17cee55, 32'hc21824af};
test_weights[8216:8223] = '{32'hc18a8001, 32'hc2beed87, 32'hc1dd0a0c, 32'h420128c4, 32'hc28b3026, 32'h41d77036, 32'hc27570e6, 32'hc176b8f9};
test_bias[1027:1027] = '{32'hc2c1b018};
test_output[1027:1027] = '{32'hc557f638};
test_input[8224:8231] = '{32'hc1ab56e0, 32'hc2944f45, 32'h4286db88, 32'hc245fc10, 32'h42ba3b7f, 32'h42336b74, 32'hc0ad4b8d, 32'h4275932e};
test_weights[8224:8231] = '{32'h42329d55, 32'h420dca59, 32'h41df3964, 32'hc158edc1, 32'hc27ceb27, 32'h42931b08, 32'h425ed148, 32'h42890ff3};
test_bias[1028:1028] = '{32'h42268970};
test_output[1028:1028] = '{32'h43a33515};
test_input[8232:8239] = '{32'hc2415c81, 32'h4289a98d, 32'hc28e5f00, 32'h41e76677, 32'h3ed01c6b, 32'hc2bd15ea, 32'h4266c190, 32'h42889c3d};
test_weights[8232:8239] = '{32'h42b37a51, 32'h428ba80e, 32'h41ee9bdc, 32'h42b291d1, 32'hc29bae4a, 32'hc2762867, 32'h4137f0dd, 32'h422ad977};
test_bias[1029:1029] = '{32'h418ca001};
test_output[1029:1029] = '{32'h462121db};
test_input[8240:8247] = '{32'h42ae93ba, 32'h42a1e75e, 32'h429902ac, 32'hc2b96b4e, 32'hc19f2cd9, 32'h427391d5, 32'hc2219f7c, 32'h411b16d0};
test_weights[8240:8247] = '{32'h42953a3e, 32'hc26b8218, 32'hc28abf4e, 32'h426475ae, 32'hc18b92d4, 32'hc24fbc37, 32'h42bdd92a, 32'h42578762};
test_bias[1030:1030] = '{32'h42901801};
test_output[1030:1030] = '{32'hc66900e0};
test_input[8248:8255] = '{32'hc0e017a5, 32'hc2847062, 32'hc2b299ae, 32'hc17f5c7c, 32'hc293ba08, 32'h42af674e, 32'hc2882995, 32'h42b52398};
test_weights[8248:8255] = '{32'h422e811c, 32'hc2a02df5, 32'h41940ece, 32'h4241578f, 32'hc24b33e1, 32'hc01e20ec, 32'hc2a8d58c, 32'hc10460fd};
test_bias[1031:1031] = '{32'hc2554fb5};
test_output[1031:1031] = '{32'h462cb816};
test_input[8256:8263] = '{32'hc2c26928, 32'hc26c389b, 32'h428d8043, 32'hc2bfe513, 32'hc2c43803, 32'h41673b58, 32'h42652d61, 32'h42c08f4c};
test_weights[8256:8263] = '{32'hc2c2031d, 32'h42a8d9be, 32'hc2901e32, 32'h42c24830, 32'hc10c71fb, 32'hc0593263, 32'hc227286e, 32'h4288d5db};
test_bias[1032:1032] = '{32'h4256ef43};
test_output[1032:1032] = '{32'hc599a079};
test_input[8264:8271] = '{32'hc2ad21b4, 32'hc26eca22, 32'h42a99987, 32'hc18fe35e, 32'hc285f151, 32'h41c917d1, 32'h42a10375, 32'hc25fb79e};
test_weights[8264:8271] = '{32'h422a6d18, 32'hc28c65bd, 32'hc158b26c, 32'hc2ae3ca3, 32'hc2ac8091, 32'h4296e567, 32'h420bd070, 32'hc2b95936};
test_bias[1033:1033] = '{32'hc2713ece};
test_output[1033:1033] = '{32'h4681252b};
test_input[8272:8279] = '{32'h41221f54, 32'hc086836b, 32'h4151bfcc, 32'hc29a8686, 32'hc21b54a4, 32'hc18617b6, 32'h428a00bc, 32'hc2898d64};
test_weights[8272:8279] = '{32'h42526f2c, 32'h424790bb, 32'h42a18320, 32'h420bcf13, 32'hc2c76922, 32'h416d994f, 32'hc2963183, 32'h42405a48};
test_bias[1034:1034] = '{32'h42862109};
test_output[1034:1034] = '{32'hc5bf2cf9};
test_input[8280:8287] = '{32'hc24c36eb, 32'h4264571d, 32'hc1dd88e3, 32'hc2b28a24, 32'hc28534fb, 32'h41f67834, 32'h42627bda, 32'hc16ebe62};
test_weights[8280:8287] = '{32'hc28b78a2, 32'h42442035, 32'h4297a30c, 32'h4298c23c, 32'hc0cd3342, 32'hc17e9628, 32'hc28f4c24, 32'h42a9e045};
test_bias[1035:1035] = '{32'hc2a99dfe};
test_output[1035:1035] = '{32'hc5faf6d4};
test_input[8288:8295] = '{32'hc2c5c8d4, 32'h42b5bc16, 32'hc1fcfc15, 32'h42936cc5, 32'hc1f95e0f, 32'hc28782b0, 32'hc2b80e7c, 32'h4269b5a0};
test_weights[8288:8295] = '{32'h424d8c6f, 32'hbf15cbdd, 32'h428cc2eb, 32'hc29dace3, 32'hc0e92709, 32'hc2b0a7bc, 32'h423ff291, 32'hc26c11e5};
test_bias[1036:1036] = '{32'h42957cf8};
test_output[1036:1036] = '{32'hc6667736};
test_input[8296:8303] = '{32'hc2c56d5a, 32'hc260eb9c, 32'h4224e514, 32'hc2b0debd, 32'h415a057c, 32'h42461353, 32'hc22b367e, 32'h420fdd0a};
test_weights[8296:8303] = '{32'hc2737771, 32'hc1b7cef0, 32'hc22c9fb6, 32'hc2acc0bb, 32'h421f0c30, 32'h428aad8a, 32'hc04f0c98, 32'h41bcb738};
test_bias[1037:1037] = '{32'hc2a956ea};
test_output[1037:1037] = '{32'h468ceb28};
test_input[8304:8311] = '{32'h3f96fb4b, 32'hc28a42e7, 32'h4113106d, 32'hc2a8247c, 32'hc20a3ed1, 32'h41e7d64d, 32'hc2095caa, 32'hc14d3d64};
test_weights[8304:8311] = '{32'hc2947255, 32'hc22b8b35, 32'hc208883c, 32'hc29fa4cf, 32'hc28a4abe, 32'h422e1132, 32'hc296ac24, 32'hc22c573e};
test_bias[1038:1038] = '{32'hc2a51466};
test_output[1038:1038] = '{32'h4679b918};
test_input[8312:8319] = '{32'h41c3ca5a, 32'hc2b436e4, 32'h4280f397, 32'hc2a333a7, 32'h420fb01c, 32'h42728668, 32'hc00b94c8, 32'hc2734337};
test_weights[8312:8319] = '{32'hc2aa0431, 32'hc280a10e, 32'hc2811eb0, 32'h428bc7d4, 32'h429b5281, 32'hc2b122ed, 32'h42638708, 32'h41bba352};
test_bias[1039:1039] = '{32'hc2905a94};
test_output[1039:1039] = '{32'hc621c759};
test_input[8320:8327] = '{32'h40170d26, 32'h42538a93, 32'h42284940, 32'h42bf889c, 32'hc1aa0160, 32'h42a04030, 32'hc2ae4eed, 32'hc258517c};
test_weights[8320:8327] = '{32'h429af7fc, 32'hc131dd3a, 32'h4292c3ac, 32'h4277448c, 32'hc1b403af, 32'h429132a2, 32'h4265ecd4, 32'hc194c834};
test_bias[1040:1040] = '{32'h3ec2744d};
test_output[1040:1040] = '{32'h462a378b};
test_input[8328:8335] = '{32'hc1fded5c, 32'h4278f776, 32'h4279c345, 32'hc13af710, 32'hc27a70ef, 32'h428a5658, 32'h41e736fc, 32'hc21241c2};
test_weights[8328:8335] = '{32'h42b4ad0f, 32'hc1f31b93, 32'h4244e1d5, 32'hc0c091aa, 32'h42351196, 32'h41a147c2, 32'hc2844e2b, 32'h42943170};
test_bias[1041:1041] = '{32'h428ee5d0};
test_output[1041:1041] = '{32'hc5eda55c};
test_input[8336:8343] = '{32'h4219f09a, 32'hc29062ef, 32'h4252cbf1, 32'h4086705c, 32'h4288782f, 32'h42c5ba9d, 32'h42b1e757, 32'h41de9aa2};
test_weights[8336:8343] = '{32'h427e20ae, 32'hc120826f, 32'h3f8473a2, 32'h4236c177, 32'hc2981807, 32'h41dfb6d6, 32'h41f598ef, 32'h42a81c7f};
test_bias[1042:1042] = '{32'h4215581c};
test_output[1042:1042] = '{32'h45be9318};
test_input[8344:8351] = '{32'hc1b8a4bd, 32'hc0c88541, 32'hc24ad2a9, 32'hc21c08fc, 32'hc217b771, 32'hc1dd3b0b, 32'hc20dcb78, 32'hc2a40d3c};
test_weights[8344:8351] = '{32'h407b8731, 32'h4254dbb0, 32'hc2a2be74, 32'h42b51da4, 32'h41ff3d64, 32'h4295c49d, 32'h42712eec, 32'h42b7a075};
test_bias[1043:1043] = '{32'h42a554c0};
test_output[1043:1043] = '{32'hc64665dd};
test_input[8352:8359] = '{32'h410d4632, 32'hc27f7bd1, 32'h42b7d2b5, 32'h41ad65bc, 32'h42bb0c21, 32'h4265dc98, 32'h4223425f, 32'hc2ab1a99};
test_weights[8352:8359] = '{32'hc28f71ea, 32'hc261d775, 32'h41f8807b, 32'hc24d7ff3, 32'hc1c35288, 32'hbfe950b8, 32'hc204e79c, 32'hc23c3c6f};
test_bias[1044:1044] = '{32'hc19ed49b};
test_output[1044:1044] = '{32'h459b81f3};
test_input[8360:8367] = '{32'h4196eeb2, 32'hc21c2426, 32'h4171529d, 32'h41adf686, 32'h4287dadd, 32'h42c63480, 32'hc1e4dd2a, 32'hc2aa5138};
test_weights[8360:8367] = '{32'hc1565163, 32'h42bf338d, 32'hc160a9fb, 32'h42803189, 32'hc1bc1921, 32'h40d99815, 32'h41673aca, 32'hc2b35b2a};
test_bias[1045:1045] = '{32'hc2830f9b};
test_output[1045:1045] = '{32'h45568262};
test_input[8368:8375] = '{32'hc2ab5297, 32'hc218a059, 32'hc25b75cf, 32'hc22b3c6c, 32'h42b9b001, 32'h42bcb309, 32'h423fba4e, 32'h41a02e15};
test_weights[8368:8375] = '{32'hc2981e44, 32'hc1f36f68, 32'h4209b809, 32'h427a884f, 32'h41d0fa5a, 32'hc272fe62, 32'h42b57330, 32'h415ed4a3};
test_bias[1046:1046] = '{32'hc2a44f1c};
test_output[1046:1046] = '{32'h4587c95b};
test_input[8376:8383] = '{32'h426f75ff, 32'hc24fe1c7, 32'hc11b3d68, 32'h426640ee, 32'hc11b44f5, 32'h42a60a11, 32'h42c56c8d, 32'hc206e43c};
test_weights[8376:8383] = '{32'h425b6877, 32'hc122c22e, 32'hc236fba5, 32'h4231c77e, 32'h42b63638, 32'h42a27554, 32'hc2b2c324, 32'h41241796};
test_bias[1047:1047] = '{32'h3f52c881};
test_output[1047:1047] = '{32'h455b21c0};
test_input[8384:8391] = '{32'hc1f7e465, 32'hc1c70bee, 32'h423e9498, 32'hc28d3e47, 32'hc22e37f0, 32'hc21460be, 32'h422951c3, 32'h425d1af9};
test_weights[8384:8391] = '{32'hc28620db, 32'h403b283a, 32'hc2459fa3, 32'hc08bfe7f, 32'h41fb6050, 32'h42ad2c64, 32'h41ab66dd, 32'h424321b6};
test_bias[1048:1048] = '{32'h42c7fc58};
test_output[1048:1048] = '{32'hc4652ad7};
test_input[8392:8399] = '{32'hc211f214, 32'h42a3abbe, 32'h42913c50, 32'hc1a7969d, 32'h42866dff, 32'hc247b65e, 32'h4164d032, 32'h426b7ef9};
test_weights[8392:8399] = '{32'h42ae7d19, 32'h427182d6, 32'h42afef24, 32'hc28639a0, 32'h41b8dc08, 32'hc0f93cc8, 32'hc27e50e6, 32'h42c12374};
test_bias[1049:1049] = '{32'hc29d97ab};
test_output[1049:1049] = '{32'h467cfc79};
test_input[8400:8407] = '{32'h428b01e9, 32'hc08f5682, 32'hc12bc314, 32'h41aac33f, 32'hc258b75c, 32'h41b189b9, 32'h418bd3eb, 32'h428f5488};
test_weights[8400:8407] = '{32'h42ad001a, 32'hc280aa1e, 32'h401f325e, 32'h41ecaba0, 32'hc1d8cdb2, 32'hc2714d31, 32'hc2ada48a, 32'hc20fcce5};
test_bias[1050:1050] = '{32'h3f84a3a9};
test_output[1050:1050] = '{32'h4537db54};
test_input[8408:8415] = '{32'hc29f6513, 32'h40550edd, 32'h427a142d, 32'hc137e2a1, 32'h412afab1, 32'h4110931e, 32'h42a0005c, 32'h424146b5};
test_weights[8408:8415] = '{32'hc1780c12, 32'h41be015e, 32'hc25f95e7, 32'h421dfc25, 32'h4269ce11, 32'hc2718591, 32'hc20e9bf3, 32'h423f4c53};
test_bias[1051:1051] = '{32'hc1a5f351};
test_output[1051:1051] = '{32'hc542d064};
test_input[8416:8423] = '{32'h42b7d3f4, 32'h418bf7cf, 32'hc2108890, 32'h4215ffc1, 32'h416cf793, 32'hc1926a7f, 32'h422de1b6, 32'hc29e0fe7};
test_weights[8416:8423] = '{32'h42155aba, 32'hc210fd50, 32'hc2493194, 32'h41b649a4, 32'hc252dd45, 32'h4205fd79, 32'hc2c30fad, 32'hc20454e6};
test_bias[1052:1052] = '{32'h42aceecc};
test_output[1052:1052] = '{32'h451e9335};
test_input[8424:8431] = '{32'hc20e37f8, 32'hc22e68ad, 32'hc2bfd7d3, 32'hc2a72d31, 32'h3f56e7fc, 32'hc2c50f96, 32'h42b3e07d, 32'hc284ebb0};
test_weights[8424:8431] = '{32'h428500b7, 32'h42820751, 32'hc2bd0f9b, 32'hc2849af3, 32'h4272e0f3, 32'h41de4406, 32'hc2302d06, 32'h42c7efb8};
test_bias[1053:1053] = '{32'hc25a5cec};
test_output[1053:1053] = '{32'hc575fd8c};
test_input[8432:8439] = '{32'hc1ee7524, 32'h424785c8, 32'h41c7b893, 32'hc237ee1c, 32'h42ba8700, 32'hc2311dd1, 32'hc1ca5985, 32'hc2c09670};
test_weights[8432:8439] = '{32'h4047fa17, 32'h41993476, 32'h42a55ef0, 32'h426a0dcd, 32'h420ffe79, 32'h4262bfdb, 32'h408a3631, 32'hc26cbe1b};
test_bias[1054:1054] = '{32'h414764ba};
test_output[1054:1054] = '{32'h45d0ebd2};
test_input[8440:8447] = '{32'hc2272944, 32'h40cdb4f7, 32'h41d56080, 32'hc1461927, 32'h419bec66, 32'hc272b691, 32'h42c4fe50, 32'hc236d7df};
test_weights[8440:8447] = '{32'h4280b856, 32'hc26f6f48, 32'hc2684d50, 32'hc25efda8, 32'h421efb3b, 32'h42ae15db, 32'hc209cd14, 32'hc2116a9e};
test_bias[1055:1055] = '{32'h42890001};
test_output[1055:1055] = '{32'hc61ddc69};
test_input[8448:8455] = '{32'hc2ab528d, 32'h41f9fe74, 32'hc2c59a2a, 32'hc23c4188, 32'hc2965b3a, 32'hc0b10a02, 32'hc1d50902, 32'hc26391ca};
test_weights[8448:8455] = '{32'hc23c7c91, 32'h42b003fe, 32'h42a5b4ef, 32'h419c64e3, 32'h426d8de1, 32'h409eedd1, 32'hc289f9b3, 32'hc217a29e};
test_bias[1056:1056] = '{32'h42b9539e};
test_output[1056:1056] = '{32'hc52a51c8};
test_input[8456:8463] = '{32'hc2a3d982, 32'hc25074f4, 32'h42b503fb, 32'hc23e5cc9, 32'h428173a9, 32'hc296015c, 32'hc221c8c8, 32'h42b75221};
test_weights[8456:8463] = '{32'hc2aba0ed, 32'hc2c5701d, 32'hc28e6e62, 32'h4288fbb6, 32'hc2b2e24a, 32'h412897a5, 32'h42b903ca, 32'hc20d0b0a};
test_bias[1057:1057] = '{32'hc1fd9432};
test_output[1057:1057] = '{32'hc62dabbc};
test_input[8464:8471] = '{32'hc20039e8, 32'h425d53dc, 32'hc28a8f6d, 32'hc2a2b036, 32'h4221e69a, 32'h42c3ccca, 32'hc28cb782, 32'h412206ed};
test_weights[8464:8471] = '{32'h42c1efcb, 32'hc0ee77d3, 32'h4290be76, 32'hc2930f88, 32'hc1ff4a1c, 32'hc247f51f, 32'hc1bac37d, 32'hc2a2b38b};
test_bias[1058:1058] = '{32'h424d0d9e};
test_output[1058:1058] = '{32'hc5f5e87b};
test_input[8472:8479] = '{32'hc1f466fa, 32'hc15884fb, 32'hc1cb9686, 32'h427c2ca6, 32'hc27ec816, 32'h4269fb42, 32'hc113366e, 32'h42b53b96};
test_weights[8472:8479] = '{32'h410e5e6f, 32'hc1a537f3, 32'hc2b7704f, 32'h42a6642a, 32'hc2a5e522, 32'hc2674e9a, 32'h427944f8, 32'hc26c2dfc};
test_bias[1059:1059] = '{32'h418c9dfe};
test_output[1059:1059] = '{32'h455fd431};
test_input[8480:8487] = '{32'hc1a76de7, 32'h41f78cc0, 32'h42806162, 32'h427893d9, 32'hc24fd9cc, 32'h42aa548c, 32'h410c2212, 32'hc203cc24};
test_weights[8480:8487] = '{32'h40dc93f5, 32'hc2035d6e, 32'hc0f88267, 32'h428dd534, 32'h4224cd24, 32'h41c4919d, 32'hc1835712, 32'hc299f970};
test_bias[1060:1060] = '{32'hc25d9424};
test_output[1060:1060] = '{32'h459d6a42};
test_input[8488:8495] = '{32'h428b05a7, 32'hc2b4f710, 32'hc2c5f7b6, 32'hc233c382, 32'hc21edafb, 32'hc0e18287, 32'h428bc574, 32'hc28342db};
test_weights[8488:8495] = '{32'hc01a9f7a, 32'h4196224d, 32'h42b626ce, 32'h412cb1e3, 32'h41ea0b9a, 32'h3f7119d4, 32'h424dfa25, 32'h41f86d12};
test_bias[1061:1061] = '{32'h42396d53};
test_output[1061:1061] = '{32'hc62abe41};
test_input[8496:8503] = '{32'h41fdc14c, 32'hc2716fa7, 32'hc275d1d3, 32'h4246ff36, 32'hc2b76aef, 32'hc2a54be6, 32'hbe9d2637, 32'hc1f675c4};
test_weights[8496:8503] = '{32'hc29a1a3f, 32'h428d2bb7, 32'hc1d0177a, 32'hc13e10aa, 32'hc2c40273, 32'hc29178e4, 32'hc2179487, 32'h429e3ee4};
test_bias[1062:1062] = '{32'hc22df7a3};
test_output[1062:1062] = '{32'h45d5886f};
test_input[8504:8511] = '{32'h41eedde7, 32'hc28ba7e2, 32'hc1d1cb0f, 32'hc2b72f2d, 32'hc2a1b7e5, 32'h411ff4d7, 32'h42275432, 32'hc2bf68ac};
test_weights[8504:8511] = '{32'hc1f09d6c, 32'h422f03fe, 32'h42b2a53e, 32'hc26a3c88, 32'hc23e5145, 32'h42983b4c, 32'hc1bd3027, 32'h40666e36};
test_bias[1063:1063] = '{32'h41bd8cdd};
test_output[1063:1063] = '{32'h4513ddfb};
test_input[8512:8519] = '{32'hc2075b48, 32'h41e24ffd, 32'hc2bb4484, 32'h42bd455b, 32'hc2961ac7, 32'h412ec37c, 32'hc25ee27b, 32'h41f11270};
test_weights[8512:8519] = '{32'h4289ea40, 32'hc23372d3, 32'h42c41916, 32'h418d42f7, 32'h402812d7, 32'h4270f731, 32'hbfe87799, 32'hc21ca6a2};
test_bias[1064:1064] = '{32'h420a75ff};
test_output[1064:1064] = '{32'hc636be93};
test_input[8520:8527] = '{32'h41e1bc88, 32'h42bdd769, 32'h40d157b4, 32'hc17eba2e, 32'h429e5aa8, 32'h41e43686, 32'h429d6593, 32'hc2b16e40};
test_weights[8520:8527] = '{32'h4271174a, 32'hc0e2ff1e, 32'h42c4a222, 32'h4204b4ce, 32'hc185af7b, 32'h42c750c7, 32'hc29b52a6, 32'h42010386};
test_bias[1065:1065] = '{32'hc287cef6};
test_output[1065:1065] = '{32'hc5c7576b};
test_input[8528:8535] = '{32'h42360880, 32'h42361180, 32'hc269908c, 32'hc2afaec6, 32'hc2b922f6, 32'hc1c30b2d, 32'h42399ec4, 32'h41795313};
test_weights[8528:8535] = '{32'hc26c5423, 32'hc2b0ac96, 32'h422cecd9, 32'hc26490c7, 32'h426ea0a3, 32'hbff17592, 32'h429ebb52, 32'h40d9e42a};
test_bias[1066:1066] = '{32'hc292d436};
test_output[1066:1066] = '{32'hc5bab99a};
test_input[8536:8543] = '{32'h4133f7af, 32'h4139516b, 32'h4244aa73, 32'h42b9fa9d, 32'h428486d7, 32'h42505784, 32'hbfdf886f, 32'h41a06a96};
test_weights[8536:8543] = '{32'h41cc5e1f, 32'hc2b706d4, 32'h42459c24, 32'h42b4ab02, 32'h42c28978, 32'h40829ff7, 32'hc29ead63, 32'h41a6288d};
test_bias[1067:1067] = '{32'hc2897d46};
test_output[1067:1067] = '{32'h46866162};
test_input[8544:8551] = '{32'hc25e694a, 32'hc265ba3e, 32'h42a437a3, 32'h42b51e87, 32'h426314b5, 32'h428d80f1, 32'hc2a06dd8, 32'h41cbcb43};
test_weights[8544:8551] = '{32'h42892d83, 32'hc2b013fa, 32'hc2183fba, 32'hc2c5b466, 32'h41d43d5d, 32'h420e4326, 32'hc28547b0, 32'h42031dd4};
test_bias[1068:1068] = '{32'h42b54024};
test_output[1068:1068] = '{32'hc4074af5};
test_input[8552:8559] = '{32'hc155ffaa, 32'hc223ac88, 32'h41ba278f, 32'hc25d5ca5, 32'hc2b8c691, 32'hc238d2eb, 32'h4262c6ee, 32'h42ab0780};
test_weights[8552:8559] = '{32'hc273fbcb, 32'h42bec80a, 32'hc29418d1, 32'hc2899816, 32'hc18c1fdd, 32'hc14555ed, 32'h4220728a, 32'hc1d85a5a};
test_bias[1069:1069] = '{32'hc231a4a9};
test_output[1069:1069] = '{32'h4489bd3e};
test_input[8560:8567] = '{32'hc290a72d, 32'hc28e179f, 32'h40e6e194, 32'hc2c2200d, 32'hc1bd1711, 32'hc27fc858, 32'h4185a382, 32'hc29498fd};
test_weights[8560:8567] = '{32'hc2850880, 32'hc0f71b60, 32'hc2a0d686, 32'h42ab0626, 32'h418e1960, 32'hc1d453e6, 32'h42859ea4, 32'hc2b15c27};
test_bias[1070:1070] = '{32'h419aa55b};
test_output[1070:1070] = '{32'h45ab46aa};
test_input[8568:8575] = '{32'h4220a694, 32'hc197789a, 32'hc28600f6, 32'h42629c85, 32'h4178ce1e, 32'h40eb23a7, 32'hc2b6f772, 32'hc21aa99a};
test_weights[8568:8575] = '{32'h429eb148, 32'hc17e6af0, 32'hc2371a6b, 32'hc24d9fd6, 32'h42abb7bd, 32'h427778c1, 32'h428cbe99, 32'h41727fb6};
test_bias[1071:1071] = '{32'hc29e0916};
test_output[1071:1071] = '{32'hc4d0d2ee};
test_input[8576:8583] = '{32'h423cab4e, 32'h42a3b07b, 32'hc2ae48d8, 32'hc1b29b48, 32'hc290e160, 32'hc2575906, 32'hc18f2d9a, 32'h425c1281};
test_weights[8576:8583] = '{32'hc292cf06, 32'h4190df3d, 32'hc28091c1, 32'h420530d9, 32'h4278587f, 32'h426ae67f, 32'hc294ac64, 32'hc205c139};
test_bias[1072:1072] = '{32'hc29cf65a};
test_output[1072:1072] = '{32'hc5a7c483};
test_input[8584:8591] = '{32'hc2a3d787, 32'h41c36d56, 32'hc2247353, 32'hc2641b4f, 32'h419cc890, 32'hc27e7f38, 32'hc2217445, 32'h42c3f361};
test_weights[8584:8591] = '{32'h410556c3, 32'h42ba2f8c, 32'hc2532048, 32'hc1cfae00, 32'h414e1e1e, 32'hc28cf74d, 32'h423bc73a, 32'hc239b79e};
test_bias[1073:1073] = '{32'h4114aa91};
test_output[1073:1073] = '{32'h455d8365};
test_input[8592:8599] = '{32'hc223312a, 32'h421990a3, 32'hc292c50b, 32'h414c2004, 32'hc20f5473, 32'hc2005e56, 32'hc2be711a, 32'hc2a4ebe6};
test_weights[8592:8599] = '{32'hc22fcde4, 32'h424233fd, 32'h42a51800, 32'hc1d8f38e, 32'h41ffa80a, 32'h42a5cecf, 32'h40e1c291, 32'h40dae19e};
test_bias[1074:1074] = '{32'h4181d03b};
test_output[1074:1074] = '{32'hc5f2df11};
test_input[8600:8607] = '{32'hc1c843c8, 32'h4294c428, 32'hc29e69df, 32'h42b5800e, 32'h4293b3cf, 32'h422bac91, 32'h429c98b6, 32'hc203e91d};
test_weights[8600:8607] = '{32'hc20a7841, 32'hc23a844d, 32'h428b2baa, 32'h40095a9f, 32'h42899ad8, 32'h423c7b00, 32'hc2a46076, 32'h4268e31d};
test_bias[1075:1075] = '{32'h424528ce};
test_output[1075:1075] = '{32'hc60e84b4};
test_input[8608:8615] = '{32'hc1f129cb, 32'h420c4d57, 32'hc1b1dee6, 32'hc17fcb84, 32'hc1438073, 32'hbfbf9b49, 32'h42a4f529, 32'hc1cd5196};
test_weights[8608:8615] = '{32'h425b0e10, 32'h420abecd, 32'h42bb5cbe, 32'h4238275d, 32'h42baea14, 32'h423ed9c0, 32'h42425b72, 32'hc20452e7};
test_bias[1076:1076] = '{32'hc21321e9};
test_output[1076:1076] = '{32'h43b0a7c2};
test_input[8616:8623] = '{32'h41dba86d, 32'h40afd72e, 32'hc123353f, 32'h42921479, 32'h42be440a, 32'hc0b6c2e6, 32'h412ad77e, 32'hc1fcaf86};
test_weights[8616:8623] = '{32'h424e91b5, 32'hc29d9e1b, 32'hc2beb61f, 32'h419828a4, 32'hc2b23951, 32'hc12c64f2, 32'hc2b6d963, 32'hc293cecb};
test_bias[1077:1077] = '{32'hc28baf9c};
test_output[1077:1077] = '{32'hc56c4e37};
test_input[8624:8631] = '{32'h42658038, 32'hc12f8526, 32'hc2aeb317, 32'hc249cd1d, 32'h4261eeea, 32'hc26005c5, 32'hc21fc958, 32'h4181411a};
test_weights[8624:8631] = '{32'hc0a4bdf2, 32'h42973ab3, 32'hc20b3cf0, 32'hc2be0e84, 32'h42815e62, 32'h4293919c, 32'h4260823d, 32'hc212baf9};
test_bias[1078:1078] = '{32'h42323302};
test_output[1078:1078] = '{32'h45570f86};
test_input[8632:8639] = '{32'h4283fb09, 32'hc2a4bb6d, 32'hc2ad405c, 32'h407e54ed, 32'h4249e558, 32'h42067478, 32'h42276ac8, 32'hc2815266};
test_weights[8632:8639] = '{32'h42aaf272, 32'hc0d495a0, 32'hc1edb22e, 32'hc19346a6, 32'h42c0eaa2, 32'hc2b67e8a, 32'hc29e8aa6, 32'h4260346d};
test_bias[1079:1079] = '{32'hc2aff313};
test_output[1079:1079] = '{32'h455839f5};
test_input[8640:8647] = '{32'h419f8f84, 32'hc285ac4d, 32'hc222ef02, 32'h41ff06a2, 32'hc2827846, 32'h425f4374, 32'hc29493a6, 32'hc2b0026d};
test_weights[8640:8647] = '{32'hc20f13e3, 32'h40cc7918, 32'h4271a7a9, 32'h429a2ce9, 32'h424261e7, 32'h41edaf6a, 32'hc0d4a927, 32'h428439d8};
test_bias[1080:1080] = '{32'hc21f8539};
test_output[1080:1080] = '{32'hc5faa168};
test_input[8648:8655] = '{32'hc2591628, 32'hc2957d19, 32'hc280604e, 32'h41ada2d6, 32'hc26da614, 32'hc2a69689, 32'h425210d3, 32'hc1f87dcb};
test_weights[8648:8655] = '{32'hc297ca9f, 32'h4256852f, 32'h425d8489, 32'hc27a36ad, 32'h421ff478, 32'h4244fd74, 32'hc286ca5c, 32'hc16eab04};
test_bias[1081:1081] = '{32'h42a4d1e3};
test_output[1081:1081] = '{32'hc65f059a};
test_input[8656:8663] = '{32'h3fa1a7ac, 32'h42aa2b76, 32'h42a97188, 32'h40672b3b, 32'h42c39057, 32'h42518e47, 32'hc21c4545, 32'hc1d4cbd2};
test_weights[8656:8663] = '{32'h4259e713, 32'h4216fa67, 32'hc2b65900, 32'hc21eccde, 32'hc25d98cb, 32'hc2689bb1, 32'h42949128, 32'h4209851d};
test_bias[1082:1082] = '{32'h42390211};
test_output[1082:1082] = '{32'hc6836acd};
test_input[8664:8671] = '{32'h422a628c, 32'h4295f8fe, 32'hc296c234, 32'h41a91850, 32'hc22f3fdf, 32'h42510daa, 32'hc2a34ea8, 32'h42348a41};
test_weights[8664:8671] = '{32'hc286476d, 32'hc0f9e3be, 32'hc261668f, 32'h4231630b, 32'h41b0bc74, 32'h4195d029, 32'h412d117b, 32'hbe54b37e};
test_bias[1083:1083] = '{32'h42a79536};
test_output[1083:1083] = '{32'h446b619c};
test_input[8672:8679] = '{32'h418e9b4b, 32'hc1748bca, 32'h42a9cb48, 32'h41dbf39c, 32'h40ea1387, 32'h42b691b9, 32'h421715e1, 32'h41c755f1};
test_weights[8672:8679] = '{32'hc1553cc7, 32'h3f2bd04e, 32'hc229aa02, 32'h4285ee75, 32'h41f3e861, 32'hc2885ad9, 32'h3f519dbe, 32'hc2c0060d};
test_bias[1084:1084] = '{32'h42ba925e};
test_output[1084:1084] = '{32'hc620913e};
test_input[8680:8687] = '{32'h422022d7, 32'hc2af8791, 32'hc213b217, 32'h421ddbc7, 32'h41a96c5d, 32'h40b0db88, 32'h4253a0b1, 32'h42a33193};
test_weights[8680:8687] = '{32'hc2532826, 32'h42591f96, 32'hc2bfe452, 32'hc26b7705, 32'hc22c34cd, 32'hc2aa48a8, 32'h413da711, 32'h4230d1f3};
test_bias[1085:1085] = '{32'hc15cd00d};
test_output[1085:1085] = '{32'hc5303bd3};
test_input[8688:8695] = '{32'h429a8f88, 32'h424fef47, 32'hc21342ae, 32'h41bfc808, 32'hc2615343, 32'hc297d026, 32'hc1af88d0, 32'hc1ce5943};
test_weights[8688:8695] = '{32'h423ef7db, 32'hc26e4fd9, 32'h417d211b, 32'hc2a1a67b, 32'hc2aa5214, 32'hc2471685, 32'hc17b781e, 32'h425bc91b};
test_bias[1086:1086] = '{32'hc23a9a95};
test_output[1086:1086] = '{32'h45acc47b};
test_input[8696:8703] = '{32'h41e55d79, 32'h4214fc0a, 32'h423c4b54, 32'hc2a383bd, 32'hc200fff1, 32'h42913de3, 32'h41b96d08, 32'hc25e895e};
test_weights[8696:8703] = '{32'hc28e0eab, 32'hc221b377, 32'hc16e11c6, 32'hc22d133c, 32'h4242f0cb, 32'h417c59ea, 32'hc2b012f3, 32'hc17afed8};
test_bias[1087:1087] = '{32'hc1affdb4};
test_output[1087:1087] = '{32'hc511122a};
test_input[8704:8711] = '{32'hc13ae9b8, 32'hc1850806, 32'hc1af3446, 32'h422725d3, 32'h42b297c6, 32'hc1a2aff1, 32'h4284d017, 32'h4248c724};
test_weights[8704:8711] = '{32'hc258841d, 32'hc28f2ef5, 32'hc28b5c1c, 32'h42bd4735, 32'hc1f7688e, 32'hc24ddd54, 32'hc22def78, 32'h42bb4d79};
test_bias[1088:1088] = '{32'hc2237fbd};
test_output[1088:1088] = '{32'h45e606d7};
test_input[8712:8719] = '{32'hc26e8ab4, 32'h426fb0cf, 32'hc2c13d8d, 32'hc220f20f, 32'hc2480e43, 32'hc113df1d, 32'h4232bf5f, 32'h3f4fa1fb};
test_weights[8712:8719] = '{32'h428f53ef, 32'h429d59ff, 32'h42633c4f, 32'h42c1f0dc, 32'hc2096456, 32'hc20a012d, 32'hc2557f94, 32'hc1849e26};
test_bias[1089:1089] = '{32'hc25f35b2};
test_output[1089:1089] = '{32'hc6125e20};
test_input[8720:8727] = '{32'h421dda16, 32'h42afb634, 32'h423bb299, 32'hc269f777, 32'h429d83cc, 32'hc2399e5e, 32'hc2963c9a, 32'h41a43717};
test_weights[8720:8727] = '{32'hc25219f0, 32'h42a703fc, 32'h41618afe, 32'h415fdabe, 32'hc2a3fd83, 32'h4046630d, 32'h428caf96, 32'hc2c3ebb8};
test_bias[1090:1090] = '{32'hc261eea3};
test_output[1090:1090] = '{32'hc60a37db};
test_input[8728:8735] = '{32'h42b48a80, 32'h42a0e48f, 32'hc171d921, 32'h41b9924e, 32'hc1e334d5, 32'hc13a4b80, 32'h413eacd2, 32'h420a06c9};
test_weights[8728:8735] = '{32'h41fe4488, 32'h42993461, 32'h41b0bf50, 32'h41549150, 32'h418a8125, 32'h42c22837, 32'hc0978b49, 32'h42166f12};
test_bias[1091:1091] = '{32'h42671f46};
test_output[1091:1091] = '{32'h4607ab0f};
test_input[8736:8743] = '{32'hc2c37502, 32'hc0f89599, 32'hc1f4ea1f, 32'hc22cd05a, 32'hc2b20f50, 32'h4297a6e7, 32'h4280fc6a, 32'h4245df48};
test_weights[8736:8743] = '{32'hc2b8e6e5, 32'hc28be477, 32'hc2baaf1e, 32'h420b1301, 32'h41b9c9ec, 32'h4290218e, 32'hc2134714, 32'h4213728c};
test_bias[1092:1092] = '{32'h42807168};
test_output[1092:1092] = '{32'h46584f94};
test_input[8744:8751] = '{32'hc265cb45, 32'h41e93438, 32'hc07d0b2e, 32'hc299bf4f, 32'h4175c11d, 32'hc14241f0, 32'h4229d738, 32'hc2ad9e4e};
test_weights[8744:8751] = '{32'h41ab64ad, 32'h424c2090, 32'hc17e0b34, 32'hc20742c7, 32'h41db68c3, 32'hc2c28fd2, 32'h429225ce, 32'hc272616e};
test_bias[1093:1093] = '{32'hc009d0f3};
test_output[1093:1093] = '{32'h464948f2};
test_input[8752:8759] = '{32'h425252a8, 32'hc2a01ae5, 32'hc227a2e9, 32'h42830785, 32'h42c2d3c2, 32'hc18a88dd, 32'hc26a785d, 32'h42048796};
test_weights[8752:8759] = '{32'hc2c58818, 32'hc29b4302, 32'hc1a816b8, 32'h42159a2e, 32'h42829aef, 32'hc0f7d8fd, 32'h4214a581, 32'h42bbedea};
test_bias[1094:1094] = '{32'h42c0037d};
test_output[1094:1094] = '{32'h46399aa0};
test_input[8760:8767] = '{32'hc24e4e27, 32'hc29800f7, 32'h41df73ca, 32'h42c32b69, 32'hc29c8bdd, 32'hc28ec8f9, 32'h4285e50e, 32'hc2b3dbc1};
test_weights[8760:8767] = '{32'h411185ee, 32'hc2884f11, 32'h429cc73b, 32'h4294d160, 32'hc1ddb96a, 32'hc27ae54d, 32'hc1864d68, 32'hc2976869};
test_bias[1095:1095] = '{32'hc15ee8e2};
test_output[1095:1095] = '{32'h46cede16};
test_input[8768:8775] = '{32'h3f82a4a3, 32'hc24bb762, 32'h4111944c, 32'h420092f4, 32'hc1afe1d2, 32'hc2a61c84, 32'h41f19769, 32'hc2978dc9};
test_weights[8768:8775] = '{32'hc1ebd41c, 32'hc2aebbd9, 32'h4291b28a, 32'h42717e51, 32'hc03627d4, 32'hc0082d86, 32'h42b5c281, 32'h429b7521};
test_bias[1096:1096] = '{32'hc2315189};
test_output[1096:1096] = '{32'h457e8442};
test_input[8776:8783] = '{32'hc288aa48, 32'h41c5b4b4, 32'hc29288c5, 32'hc2affba3, 32'h41f76073, 32'hc29d6bfb, 32'hc2aa3faa, 32'hc2b433ce};
test_weights[8776:8783] = '{32'h42a40f3e, 32'h41f3a2f5, 32'h42369699, 32'h4233b8fe, 32'h4229cf6c, 32'h4196543c, 32'hc28bcf53, 32'h428f8fbf};
test_bias[1097:1097] = '{32'h418bc473};
test_output[1097:1097] = '{32'hc64841a6};
test_input[8784:8791] = '{32'h42526bfa, 32'hc1c06c57, 32'hc0d55e6c, 32'hc1890e1e, 32'hc2bbdd8b, 32'hc1393f10, 32'h42230b39, 32'h4295a809};
test_weights[8784:8791] = '{32'hc29fec5f, 32'hc1f22619, 32'h409ebe78, 32'hc2907e1c, 32'hc227c027, 32'h429feec8, 32'hc20ae399, 32'h42b1ab3f};
test_bias[1098:1098] = '{32'hc1ce250e};
test_output[1098:1098] = '{32'h45b9cfdf};
test_input[8792:8799] = '{32'hc20d2c2d, 32'h41fd4d7d, 32'hc253571c, 32'h4201bb51, 32'hc140098a, 32'h40531378, 32'h429a93f2, 32'h428b1d83};
test_weights[8792:8799] = '{32'h42b67234, 32'hc218c8fc, 32'h42876621, 32'hc08b85c3, 32'h424987c4, 32'hc1ab9fae, 32'hc2b54e93, 32'h42334eae};
test_bias[1099:1099] = '{32'hc2133c29};
test_output[1099:1099] = '{32'hc6473000};
test_input[8800:8807] = '{32'hc2acfaa5, 32'h41e4085e, 32'h41c5626a, 32'h4145a863, 32'hc14fd70a, 32'h42c6eba1, 32'hc29b6ed0, 32'hc1a54396};
test_weights[8800:8807] = '{32'h4281bb4a, 32'hc29b6fd1, 32'hc2823239, 32'h42ad9bdb, 32'h42a9d616, 32'h429cc578, 32'hc0b9a3ff, 32'h41fec55b};
test_bias[1100:1100] = '{32'hc288649c};
test_output[1100:1100] = '{32'hc4f2ac2e};
test_input[8808:8815] = '{32'hc2be211c, 32'h422926b5, 32'hc1e0dc94, 32'hc0a5ad70, 32'hc23b4e3d, 32'h42547563, 32'hc2a9e381, 32'hc1899992};
test_weights[8808:8815] = '{32'h42b31f5b, 32'hc27328de, 32'hc27d5d4a, 32'hc1aa3a1c, 32'hc1acae0b, 32'hc2b2b1d4, 32'hc2130cfa, 32'h42bc724d};
test_bias[1101:1101] = '{32'h421f56a5};
test_output[1101:1101] = '{32'hc631ecab};
test_input[8816:8823] = '{32'h419e4fe0, 32'h429f8127, 32'hc1d72280, 32'h42959f15, 32'h3faf5cbb, 32'h42a1f046, 32'h422e21a1, 32'h42b8dd28};
test_weights[8816:8823] = '{32'h42878ad2, 32'h420ccb48, 32'h42496ac3, 32'h41937431, 32'hc2b31783, 32'h42c3bb31, 32'h4243a4be, 32'hc09b19b1};
test_bias[1102:1102] = '{32'h41d6bb58};
test_output[1102:1102] = '{32'h4655ca32};
test_input[8824:8831] = '{32'hc2be4dac, 32'hc28b2c7c, 32'h42bdc835, 32'h424bd9ef, 32'hc2627ca6, 32'h42a9c213, 32'hc2a40686, 32'h420c6f7a};
test_weights[8824:8831] = '{32'hc29f80fb, 32'hc26fb102, 32'h42962033, 32'h423f877b, 32'h41eb8181, 32'h421f14e8, 32'hc1cbedae, 32'h424b7462};
test_bias[1103:1103] = '{32'h42077e27};
test_output[1103:1103] = '{32'h46d278e6};
test_input[8832:8839] = '{32'h42bc5cf6, 32'h42960524, 32'hc2710371, 32'hc20e5a94, 32'h4298c7f3, 32'h414ce3b2, 32'hc114c10e, 32'h4205c94b};
test_weights[8832:8839] = '{32'hc2b72991, 32'hbf970ed6, 32'hc20a2f73, 32'h40fcbc21, 32'hc170e0b2, 32'hc1395c24, 32'h42857baf, 32'h4114293c};
test_bias[1104:1104] = '{32'hc2c20a32};
test_output[1104:1104] = '{32'hc606ae22};
test_input[8840:8847] = '{32'hc19b2c5f, 32'hc29d23b9, 32'h4197b1ce, 32'hc1955776, 32'hc2a127b2, 32'h4186be60, 32'hc23f984d, 32'h413d29c5};
test_weights[8840:8847] = '{32'hc29825ef, 32'h427ef3a5, 32'hc22370bb, 32'hc2827797, 32'h42c1ec86, 32'h41b21b8a, 32'h42a65f83, 32'h410eb61a};
test_bias[1105:1105] = '{32'h42858e6c};
test_output[1105:1105] = '{32'hc6600e57};
test_input[8848:8855] = '{32'h40957268, 32'h42270d79, 32'hc2570bb4, 32'hc139e460, 32'h415d0248, 32'hc292dcbf, 32'h42aef13b, 32'hc1b80b02};
test_weights[8848:8855] = '{32'hc28e9ff6, 32'h42a0f441, 32'h4292743d, 32'h4097492e, 32'h423b65e9, 32'h406eddbf, 32'hc0cf393a, 32'h422a5ddb};
test_bias[1106:1106] = '{32'hc28a3bec};
test_output[1106:1106] = '{32'hc509e1c2};
test_input[8856:8863] = '{32'hc21e6b36, 32'h4278cf09, 32'hc1f26991, 32'hc2b77c93, 32'hc2776836, 32'hc2c4881c, 32'hc2415109, 32'h40cf7452};
test_weights[8856:8863] = '{32'hc1cc39f8, 32'hc194176c, 32'hc28637f9, 32'h428e3661, 32'hc2306bd1, 32'hc2a9e34d, 32'h40660aa5, 32'hc1c5fba7};
test_bias[1107:1107] = '{32'h42b6ef68};
test_output[1107:1107] = '{32'h45c1cfd5};
test_input[8864:8871] = '{32'hc1dd6533, 32'h42b410a6, 32'h42a4725a, 32'h41b19166, 32'h41fadce9, 32'hc252ac3a, 32'h420cd15c, 32'hc2457b28};
test_weights[8864:8871] = '{32'hc25b3287, 32'h4224693e, 32'hc2bf065d, 32'hc2ba3350, 32'hc1ef3874, 32'hc260800c, 32'hc0e71d5f, 32'h4248ddd0};
test_bias[1108:1108] = '{32'hc2a5fd94};
test_output[1108:1108] = '{32'hc5abe684};
test_input[8872:8879] = '{32'hc2a0bbbb, 32'hc22f04fe, 32'h429add15, 32'h4177fe7a, 32'hc18c4838, 32'h420c8056, 32'hc0e08764, 32'hc1e56c43};
test_weights[8872:8879] = '{32'h41a64221, 32'hc2731994, 32'hc261261e, 32'hc271e3e1, 32'h4024eec3, 32'h423d15ac, 32'hc29ca4ff, 32'h425ed737};
test_bias[1109:1109] = '{32'h42110b11};
test_output[1109:1109] = '{32'hc5677562};
test_input[8880:8887] = '{32'hc1a13e98, 32'h42775712, 32'h42b62e57, 32'hc2a12688, 32'h417a8021, 32'h429ae574, 32'h3fdc4ccb, 32'hc1fe6ee3};
test_weights[8880:8887] = '{32'hc1afc0e8, 32'h42b716cd, 32'hc2a6732a, 32'hc211d3ef, 32'hc2154d27, 32'hc285df7e, 32'hc2b42435, 32'h42429b12};
test_bias[1110:1110] = '{32'h42355a3a};
test_output[1110:1110] = '{32'hc5ba6bf6};
test_input[8888:8895] = '{32'hc241d0fc, 32'h42c2f04f, 32'hc095bed5, 32'hc12139bd, 32'h42946a56, 32'hc204d896, 32'h41f26b27, 32'h4283e800};
test_weights[8888:8895] = '{32'h407f580a, 32'hc2b74289, 32'hc27b2f48, 32'hc2a1673a, 32'h416f56de, 32'hc205bb7b, 32'h42a2d331, 32'h42597a74};
test_bias[1111:1111] = '{32'hc2aa415e};
test_output[1111:1111] = '{32'h432abdb9};
test_input[8896:8903] = '{32'hc29a9c7a, 32'hc1d4d18d, 32'h4213497f, 32'h429b7db9, 32'h412f826e, 32'h42a3602c, 32'h41d6b8e8, 32'hc1bf5d65};
test_weights[8896:8903] = '{32'hc1f31fcc, 32'h41c1e2ff, 32'hc23b324c, 32'h41055a98, 32'hc2c391f1, 32'hc2bd03e0, 32'hc2103e67, 32'h42972543};
test_bias[1112:1112] = '{32'h41d1f18f};
test_output[1112:1112] = '{32'hc62a830e};
test_input[8904:8911] = '{32'h42575607, 32'h42aaee4c, 32'hc18d845b, 32'h42a114ca, 32'h4283b8c7, 32'h3fba5873, 32'h42aa9253, 32'hc123b499};
test_weights[8904:8911] = '{32'hc06ab6f5, 32'h4241bad8, 32'hc1e5d016, 32'hc29531ef, 32'hc298e373, 32'h429d8f4f, 32'h42ae2d28, 32'hc14e572a};
test_bias[1113:1113] = '{32'hc20638b3};
test_output[1113:1113] = '{32'h4482f5ee};
test_input[8912:8919] = '{32'h4208af42, 32'hc1284952, 32'hc28c862e, 32'hc2614e42, 32'h4034babc, 32'hc242c001, 32'hc2552223, 32'hc21bb53f};
test_weights[8912:8919] = '{32'hc28d1909, 32'h42564b9b, 32'hc183f508, 32'hc2890660, 32'hc1c78007, 32'hc063ce4b, 32'hc21a833b, 32'hc27f044d};
test_bias[1114:1114] = '{32'h40a65ce4};
test_output[1114:1114] = '{32'h45d11eea};
test_input[8920:8927] = '{32'h428c31a7, 32'h4290edcb, 32'hc18b6f74, 32'h4182c2f7, 32'hc1282fbe, 32'hc1e66f30, 32'h421a556a, 32'hc27ca4e9};
test_weights[8920:8927] = '{32'hc2bc61f1, 32'hc2742db3, 32'h3e3f44d6, 32'hc0910a46, 32'hc1ff8828, 32'h429d22bc, 32'h42521696, 32'h41c1190c};
test_bias[1115:1115] = '{32'h4292ffdc};
test_output[1115:1115] = '{32'hc6429d43};
test_input[8928:8935] = '{32'hc2407fea, 32'hc2c4adcb, 32'hbf7f0d0f, 32'h425e3bbf, 32'hc20be3d1, 32'h4279e376, 32'hc2959689, 32'hc2077612};
test_weights[8928:8935] = '{32'hc29bdf43, 32'hc1e2f430, 32'hc2aa758f, 32'h42ac7607, 32'h4064762d, 32'hc2b47cf6, 32'h4295946f, 32'hc29df6e0};
test_bias[1116:1116] = '{32'hc23b2d1b};
test_output[1116:1116] = '{32'h4527fc33};
test_input[8936:8943] = '{32'h4277e830, 32'h41a0ab0f, 32'hc2bba9c6, 32'hc2b5e23a, 32'h4246d43b, 32'h41057ff4, 32'h4166701f, 32'hc08f8bfb};
test_weights[8936:8943] = '{32'hc155c009, 32'hc29161ee, 32'hc205ec24, 32'h4221b727, 32'h416915db, 32'hc2bfbcb1, 32'h41f86bb8, 32'h4291f81b};
test_bias[1117:1117] = '{32'hc286705e};
test_output[1117:1117] = '{32'hc531e2a3};
test_input[8944:8951] = '{32'h42ad091a, 32'hc1d89283, 32'hc18b3041, 32'h42903f97, 32'hc1cb4a1d, 32'hc1930ef6, 32'hc242b956, 32'hc1e36bfc};
test_weights[8944:8951] = '{32'h428482ae, 32'hc2c16cfe, 32'h42b33dc8, 32'h4220afcf, 32'hc291cf69, 32'hc26472b1, 32'hc158e5e6, 32'h421a01ae};
test_bias[1118:1118] = '{32'hc272d627};
test_output[1118:1118] = '{32'h463cfea4};
test_input[8952:8959] = '{32'h4215aebc, 32'h42b0ff13, 32'h42050291, 32'hbfd10365, 32'hc1f2edec, 32'hc1b630f1, 32'hc2b2ffa6, 32'hc23718e6};
test_weights[8952:8959] = '{32'h40d8bacd, 32'h42631af5, 32'hc1fe3a2b, 32'hc1efcd4a, 32'hc228d3ec, 32'hc24ec671, 32'hc28ecee8, 32'h428cf4d2};
test_bias[1119:1119] = '{32'hc2befb63};
test_output[1119:1119] = '{32'h46191901};
test_input[8960:8967] = '{32'hc1b8f686, 32'hc26fe94f, 32'hc127c024, 32'hc1b9b44a, 32'hc2bd14e7, 32'h4272fb9e, 32'h42c5896d, 32'hc1a96ee7};
test_weights[8960:8967] = '{32'h4275fe01, 32'hc12c34f3, 32'h4221e5f7, 32'h42b348c8, 32'h427cfb79, 32'h3fd97b91, 32'hc1e251e4, 32'h429bcabf};
test_bias[1120:1120] = '{32'h40bd3302};
test_output[1120:1120] = '{32'hc6546e87};
test_input[8968:8975] = '{32'h42689f73, 32'hc149bc6d, 32'hc1a1c823, 32'hc288464d, 32'hc2bf143b, 32'hc2ba0b09, 32'hc2b7f703, 32'hc1c0bf62};
test_weights[8968:8975] = '{32'h3ff248a6, 32'hc223a14e, 32'h42b7a89f, 32'h42b55cfc, 32'h42a38a8f, 32'hbfd6f564, 32'hc210f31e, 32'h42ba3c66};
test_bias[1121:1121] = '{32'h427c3c08};
test_output[1121:1121] = '{32'hc659656a};
test_input[8976:8983] = '{32'h41e1201e, 32'hc25962fc, 32'hc285d17b, 32'hc2c49ea7, 32'hc20ff5ca, 32'hc257182a, 32'hc2b5fb77, 32'h42744189};
test_weights[8976:8983] = '{32'h408bc6cb, 32'h41b8db17, 32'h42b25664, 32'hc28d9daa, 32'h40898ad0, 32'hc20a07b6, 32'h423a48e9, 32'hc283b5da};
test_bias[1122:1122] = '{32'hbf875c38};
test_output[1122:1122] = '{32'hc5d14871};
test_input[8984:8991] = '{32'hc235f072, 32'hc282293a, 32'h4268a78f, 32'hc28c86d7, 32'hc1923c51, 32'h4285be3d, 32'hc13601aa, 32'hc26b4177};
test_weights[8984:8991] = '{32'h4248e7e8, 32'h420f4284, 32'h3fa80255, 32'hbf2cee47, 32'hc2b73dc8, 32'h42baa4e0, 32'hc2c59847, 32'hc2c37ee5};
test_bias[1123:1123] = '{32'hc286badd};
test_output[1123:1123] = '{32'h461fd4d2};
test_input[8992:8999] = '{32'hc2afc1fe, 32'hc2914b2f, 32'h42c512d9, 32'h42ba00d7, 32'hc1b9c906, 32'h41c53fe8, 32'hc0444ad7, 32'h3fa9d965};
test_weights[8992:8999] = '{32'h427443ee, 32'hbe6cd4c1, 32'h421c3bc3, 32'h42aca38e, 32'hc1ffcbd9, 32'h40c15bbc, 32'hc1f6291b, 32'h428daf70};
test_bias[1124:1124] = '{32'h425cad25};
test_output[1124:1124] = '{32'h45ef6fd2};
test_input[9000:9007] = '{32'h4284ab6d, 32'hc2709614, 32'h42b31a28, 32'hc2ab5ffc, 32'hc2a42cb3, 32'hbf5e0966, 32'hc2a60dca, 32'hc2b30c8d};
test_weights[9000:9007] = '{32'hc13bb620, 32'hc2c1ff74, 32'hc2312141, 32'hc2847838, 32'h41849854, 32'h42a29d51, 32'h41c230dd, 32'hc15e2928};
test_bias[1125:1125] = '{32'hc1fe8abc};
test_output[1125:1125] = '{32'h458d952f};
test_input[9008:9015] = '{32'hc26af73f, 32'hc23124bd, 32'hc239d754, 32'hc2187fd5, 32'hc21b080c, 32'h4075ffdd, 32'h4208321e, 32'h429df9bf};
test_weights[9008:9015] = '{32'h427de3a3, 32'hc2434826, 32'hc19c7ab0, 32'h42b647bb, 32'hc2846ce7, 32'h41a10ea1, 32'hc2c0bed3, 32'h41ad0814};
test_bias[1126:1126] = '{32'h41d61c38};
test_output[1126:1126] = '{32'hc53dae5e};
test_input[9016:9023] = '{32'hc210e53e, 32'hc20c6765, 32'hc2495a5b, 32'h40a1b121, 32'hc18527da, 32'hc2c47396, 32'hc262c3a0, 32'h420c8e9c};
test_weights[9016:9023] = '{32'h426a1a83, 32'h4035c1f6, 32'hc2a1ca99, 32'hc29dcdc7, 32'hc1a9359f, 32'h4227b1a0, 32'h423a1234, 32'hc2c0da27};
test_bias[1127:1127] = '{32'h42480685};
test_output[1127:1127] = '{32'hc6017e93};
test_input[9024:9031] = '{32'hc1fd3865, 32'hc2bc4101, 32'h4184b9f5, 32'h40d05071, 32'hc28a7bf8, 32'hc27f8a32, 32'hc2aa4d7a, 32'h42a1fa76};
test_weights[9024:9031] = '{32'h411fa869, 32'hc1e1c0b1, 32'h4236bcb7, 32'hc29b68cb, 32'h42912e2c, 32'hc28592f9, 32'h421134cf, 32'hc291feed};
test_bias[1128:1128] = '{32'hc2594d2b};
test_output[1128:1128] = '{32'hc5e1c56e};
test_input[9032:9039] = '{32'h42427129, 32'h4200691c, 32'hc2bb7b46, 32'hc128135f, 32'hc24b1962, 32'h41e623db, 32'hc201896b, 32'hc21fec20};
test_weights[9032:9039] = '{32'h420d479e, 32'hc210cd43, 32'hc1dbff14, 32'h42a7c99d, 32'h41bf76bc, 32'hc2b1ba45, 32'hc1882a8c, 32'hc1373165};
test_bias[1129:1129] = '{32'hc19eea0f};
test_output[1129:1129] = '{32'hc404c942};
test_input[9040:9047] = '{32'hc2671c28, 32'hc282a19e, 32'hc29c111b, 32'hc292a931, 32'hc2a59c10, 32'hc24a4416, 32'h42b4d4be, 32'hc1b6bf81};
test_weights[9040:9047] = '{32'hc2c18701, 32'h420223df, 32'hc26992ea, 32'hc2b213c0, 32'h415d0253, 32'hc19a24dc, 32'hc028ba9a, 32'h429802b7};
test_bias[1130:1130] = '{32'h417cada2};
test_output[1130:1130] = '{32'h46421d45};
test_input[9048:9055] = '{32'hc205cb63, 32'hc285e85b, 32'hc2a84a01, 32'hc21b5591, 32'hc2863c99, 32'hc12a93c3, 32'h42698f0d, 32'hc1e7bba9};
test_weights[9048:9055] = '{32'hc24dd35c, 32'hc14ad9bf, 32'h412f745f, 32'hc28e00d1, 32'hc1baecfa, 32'h42317514, 32'hc2a1e3ab, 32'hbec6e026};
test_bias[1131:1131] = '{32'hc2145791};
test_output[1131:1131] = '{32'h443ae97d};
test_input[9056:9063] = '{32'h42a9b0fc, 32'hc281616e, 32'h42434c08, 32'h425d8d86, 32'hc0c0c8a2, 32'hc1e1ffe8, 32'h423c5cdb, 32'hc1ba318e};
test_weights[9056:9063] = '{32'hc2474952, 32'h41bed892, 32'h41bbf3a5, 32'h42ad459a, 32'h4249ed4b, 32'h411a6b8a, 32'hc2c04e14, 32'hc26159ea};
test_bias[1132:1132] = '{32'h41ae5537};
test_output[1132:1132] = '{32'hc560c598};
test_input[9064:9071] = '{32'hc284a29f, 32'h42bf9344, 32'h4149d514, 32'hc2ac8cad, 32'h42815c2a, 32'hc21597b6, 32'hc1763809, 32'hc176eee5};
test_weights[9064:9071] = '{32'hc23cf13c, 32'hc286bd5a, 32'h429f4fe5, 32'h41e227b2, 32'h427d18bc, 32'h4211e475, 32'hc2b8c72e, 32'h42105a5b};
test_bias[1133:1133] = '{32'h429e7638};
test_output[1133:1133] = '{32'hc4874641};
test_input[9072:9079] = '{32'hc0649aa3, 32'hc201b952, 32'hc13ab7ba, 32'h4204b4b7, 32'h41aa37b7, 32'h4246a886, 32'hc1161a23, 32'hc2a955b8};
test_weights[9072:9079] = '{32'h42684623, 32'hc2a34fcb, 32'h42b31492, 32'h427d74f1, 32'hc1ed8cea, 32'hc2b086ee, 32'hc297ddad, 32'hc20f07ad};
test_bias[1134:1134] = '{32'h42b0234d};
test_output[1134:1134] = '{32'h45106970};
test_input[9080:9087] = '{32'hc261b9ee, 32'hc1fae872, 32'hc2033785, 32'hc25b5812, 32'hc2b29d20, 32'h42bff88f, 32'h4190d025, 32'hc2ab7073};
test_weights[9080:9087] = '{32'h428693b7, 32'hc24f4ba9, 32'h429a82ff, 32'hc27eed36, 32'h4293940f, 32'hc278bd55, 32'hc05d8792, 32'h422bd02a};
test_bias[1135:1135] = '{32'hc22e4213};
test_output[1135:1135] = '{32'hc6892c78};
test_input[9088:9095] = '{32'h421009d1, 32'hc2c0bc42, 32'hc1fe7e31, 32'h41d654f1, 32'hc2946796, 32'h41a7bb24, 32'hc1f4e5a8, 32'h402d4a8a};
test_weights[9088:9095] = '{32'h42afa960, 32'h41e5ea85, 32'h421b4029, 32'hc24d4fec, 32'hc2be0101, 32'h42b59608, 32'h409fb0b0, 32'h429fb146};
test_bias[1136:1136] = '{32'h42a4d831};
test_output[1136:1136] = '{32'h45d71153};
test_input[9096:9103] = '{32'h428abbe9, 32'h426308fa, 32'h40df3892, 32'h42acc1c3, 32'hc29ad17e, 32'hc29f9def, 32'h411ea7e6, 32'hc218b340};
test_weights[9096:9103] = '{32'h40e9ada5, 32'h42724ec5, 32'hc2bab760, 32'h42836163, 32'h428f6a07, 32'h4293eaa8, 32'h428f1a41, 32'hc29f9dea};
test_bias[1137:1137] = '{32'hc2085780};
test_output[1137:1137] = '{32'h449a9404};
test_input[9104:9111] = '{32'hc17106a9, 32'h427ad4e0, 32'hc1e13cc5, 32'h422a36de, 32'hc29f41e4, 32'hc2b0c4b9, 32'h428f2c0e, 32'h40c56f75};
test_weights[9104:9111] = '{32'hc2090215, 32'h420a2426, 32'h41862b52, 32'hc27b6292, 32'hc27c5843, 32'h42af8ef4, 32'hc232ef8a, 32'h428ed27e};
test_bias[1138:1138] = '{32'h421be821};
test_output[1138:1138] = '{32'hc5b913df};
test_input[9112:9119] = '{32'h42bb6a00, 32'hc036579d, 32'h42c5cedc, 32'h4287a92e, 32'h41c561df, 32'h421386d5, 32'h4279d767, 32'h427fa6b2};
test_weights[9112:9119] = '{32'hc24d4d20, 32'h41ecb215, 32'h41adf59c, 32'hc2a1c47f, 32'hc2c2f6ad, 32'hbf3ac8ed, 32'hc1eaf68e, 32'h410bb15b};
test_bias[1139:1139] = '{32'hc14a18cb};
test_output[1139:1139] = '{32'hc63abae5};
test_input[9120:9127] = '{32'hc2665452, 32'h40ae4cd7, 32'h42725c9d, 32'hc26292ec, 32'h408dd654, 32'hc1af0ee4, 32'h423d2ad2, 32'h42376a06};
test_weights[9120:9127] = '{32'h42044dd0, 32'hc250119e, 32'h42bd4630, 32'hc202e7d5, 32'h42997d06, 32'h412dcccb, 32'h428ab68f, 32'h4152c34f};
test_bias[1140:1140] = '{32'hc2a0ce00};
test_output[1140:1140] = '{32'h461167f6};
test_input[9128:9135] = '{32'hc29492fc, 32'h42036af5, 32'hc108eaf0, 32'h428f280c, 32'h3f904124, 32'h40c30511, 32'hc226e2e3, 32'hc2b6f05d};
test_weights[9128:9135] = '{32'h4298781a, 32'h42b80878, 32'hc1a6933d, 32'h40edd225, 32'hc28567d4, 32'hbf620a07, 32'h42b67a01, 32'h4227849d};
test_bias[1141:1141] = '{32'hc2a2618e};
test_output[1141:1141] = '{32'hc61803fa};
test_input[9136:9143] = '{32'hc2b4639c, 32'hc2c5b2a3, 32'h42629991, 32'hc29f3939, 32'h4207fb2e, 32'h4298717d, 32'h42566f09, 32'h41c414cb};
test_weights[9136:9143] = '{32'hc2a7afdc, 32'hc06288dd, 32'h41a2b8e4, 32'hc113353f, 32'hc21da7a5, 32'h42915c48, 32'hc2c7b31a, 32'hc17a30f7};
test_bias[1142:1142] = '{32'hc263b69d};
test_output[1142:1142] = '{32'h46002f30};
test_input[9144:9151] = '{32'hc1e07d9b, 32'hc248e65b, 32'hc28e51cb, 32'hc209368d, 32'h41e4c310, 32'h426dfe7a, 32'hc2201cdc, 32'h41d50fe7};
test_weights[9144:9151] = '{32'h4128de4b, 32'hc2868bad, 32'h42ba8427, 32'h4297c131, 32'h428dd8ef, 32'h41d56bd9, 32'h42ae3207, 32'h429a7f5a};
test_bias[1143:1143] = '{32'h428de767};
test_output[1143:1143] = '{32'hc573b28f};
test_input[9152:9159] = '{32'h42c2f820, 32'h4142f9fc, 32'hc259091f, 32'hc2a62ffb, 32'hc214e545, 32'hc1a410b6, 32'hc2c36a39, 32'hc276f392};
test_weights[9152:9159] = '{32'hc28b0784, 32'hc2b60ed2, 32'hc1f3aa31, 32'h41889940, 32'hc2927ecc, 32'hc2ae5843, 32'h42ba1772, 32'hc23668c5};
test_bias[1144:1144] = '{32'hc10c60c9};
test_output[1144:1144] = '{32'hc61339b4};
test_input[9160:9167] = '{32'hc28830d0, 32'h4271743b, 32'h42131a04, 32'h4269173d, 32'hc2bbb7f6, 32'hc258829a, 32'h42658869, 32'h4210474e};
test_weights[9160:9167] = '{32'hc207b2f1, 32'h42905318, 32'h42b04824, 32'h428e7c90, 32'hc2450083, 32'hc230caa0, 32'hc200902d, 32'h41a95e95};
test_bias[1145:1145] = '{32'hc2b75829};
test_output[1145:1145] = '{32'h469b7b35};
test_input[9168:9175] = '{32'hc26861ae, 32'h42bbcade, 32'hc2b45843, 32'hc27259d0, 32'hc299830f, 32'h4181d32a, 32'h428c26cd, 32'h42b3338e};
test_weights[9168:9175] = '{32'hc29708dc, 32'hc262a306, 32'hc11c9059, 32'hc2937fa5, 32'hc25e7dd3, 32'hc1ce0829, 32'h42b60a54, 32'h4251c236};
test_bias[1146:1146] = '{32'hc27db05a};
test_output[1146:1146] = '{32'h4696a580};
test_input[9176:9183] = '{32'hc23ce00c, 32'h41d74df9, 32'hc0ac2c06, 32'hc1a9adea, 32'hc26d77a0, 32'hc0e3dc90, 32'h41f9b13b, 32'hc281b703};
test_weights[9176:9183] = '{32'h42874b35, 32'h4152283f, 32'h4274f334, 32'h42a3084a, 32'h426a3597, 32'hc1e64d68, 32'h3e3da8b4, 32'h41b87a75};
test_bias[1147:1147] = '{32'h420932c2};
test_output[1147:1147] = '{32'hc61666f0};
test_input[9184:9191] = '{32'h42af11d4, 32'hc2aca012, 32'hc299a454, 32'h42558b8f, 32'hc28824a7, 32'h40ce6e86, 32'hc2c084cf, 32'h42514590};
test_weights[9184:9191] = '{32'h420a598d, 32'h4135a426, 32'hc2c45f93, 32'h423aff31, 32'hc1e05e8e, 32'h410ef131, 32'h41bc71fb, 32'h4191251b};
test_bias[1148:1148] = '{32'hc2206b12};
test_output[1148:1148] = '{32'h46465aea};
test_input[9192:9199] = '{32'h42c72c6f, 32'h423b4035, 32'hc116f4cc, 32'hc2c7c5dc, 32'hc1b2f20c, 32'h422b82e4, 32'h42a2dba1, 32'hc2a43487};
test_weights[9192:9199] = '{32'h42a156bc, 32'h3ff8aea2, 32'hc1c51a78, 32'h429a4f8e, 32'hc27f5938, 32'hc06f041a, 32'hc2c6d46e, 32'h4201e77e};
test_bias[1149:1149] = '{32'h429403ac};
test_output[1149:1149] = '{32'hc6090661};
test_input[9200:9207] = '{32'hc2b062af, 32'hc2656a28, 32'hbff0ef01, 32'hc24908a2, 32'hc19144e5, 32'hc23f5dd7, 32'hc1d213c4, 32'h424bf0b5};
test_weights[9200:9207] = '{32'h42b73f7d, 32'h41ea4045, 32'h41b4a43c, 32'h4213afc0, 32'h41d096c6, 32'hc1fce4a4, 32'hc2c22709, 32'hc276351f};
test_bias[1150:1150] = '{32'hc2a9cbad};
test_output[1150:1150] = '{32'hc630748c};
test_input[9208:9215] = '{32'h42007ada, 32'h41dffc6c, 32'hc285dafa, 32'hc1a4c1c4, 32'h41e17156, 32'h422282c8, 32'h415916b4, 32'h41ee347c};
test_weights[9208:9215] = '{32'h4199af24, 32'hc0ed5349, 32'h42a196e7, 32'hc2185ac0, 32'hc2b6c52b, 32'hc237aa40, 32'hc2c76118, 32'hc2c47d64};
test_bias[1151:1151] = '{32'h42c2f62b};
test_output[1151:1151] = '{32'hc6488af7};
test_input[9216:9223] = '{32'h4244b9b2, 32'h41c2b112, 32'h42bbfcfb, 32'hc0c66a36, 32'hc14d7e19, 32'hc20d1605, 32'h41f2ca39, 32'hc1a421b9};
test_weights[9216:9223] = '{32'hc29992ed, 32'h4271896c, 32'hc2b09bd4, 32'h413fa5f3, 32'hc1f4c0fc, 32'hc2418bae, 32'h426258e0, 32'h42c549f9};
test_bias[1152:1152] = '{32'h425169a7};
test_output[1152:1152] = '{32'hc60a0f6f};
test_input[9224:9231] = '{32'hc2803d2e, 32'hc2c0c929, 32'h4135293c, 32'h428f034f, 32'h4207fbca, 32'hc1ce0173, 32'hc205d4c4, 32'hc1eb9510};
test_weights[9224:9231] = '{32'h42b1d584, 32'h42a51650, 32'hc259ae23, 32'h42868b26, 32'hc1f6c560, 32'h42505e3d, 32'h41eb8aa8, 32'hc2285ee3};
test_bias[1153:1153] = '{32'hc29d966e};
test_output[1153:1153] = '{32'hc636788e};
test_input[9232:9239] = '{32'hc29cf50d, 32'hc2ac9d2e, 32'hc2126c3d, 32'hc193f2ff, 32'hc293187d, 32'h4195223d, 32'h4295f27a, 32'hc25b1fa7};
test_weights[9232:9239] = '{32'h3ef93b95, 32'hc1bcf26d, 32'hc2b8c70f, 32'h425b5bc1, 32'hc225aa2d, 32'h3e01ef4c, 32'hc268f575, 32'h423affb6};
test_bias[1154:1154] = '{32'h42b1c2e5};
test_output[1154:1154] = '{32'h441078b5};
test_input[9240:9247] = '{32'h42b55fbf, 32'h42a10343, 32'h417a56dc, 32'h4196a6db, 32'h4156a5a0, 32'h42c0153d, 32'h42a9b787, 32'h42c5cdb5};
test_weights[9240:9247] = '{32'hc1fc115e, 32'hc028a197, 32'hc24aeba6, 32'h42b35c41, 32'hc10c1ecc, 32'h41f6c9cd, 32'h3fdf66a3, 32'h4188bc09};
test_bias[1155:1155] = '{32'hc2c1aae8};
test_output[1155:1155] = '{32'h4516c7a6};
test_input[9248:9255] = '{32'h42b23f97, 32'h42141f41, 32'hc1621315, 32'h40e10d83, 32'hc25176e7, 32'h41619276, 32'hc232dad9, 32'hc214f07a};
test_weights[9248:9255] = '{32'hbff91677, 32'h41ef8656, 32'h42b97e9a, 32'h428128f0, 32'h42069a78, 32'hc1b02f42, 32'h42a22d3b, 32'hc2b2a496};
test_bias[1156:1156] = '{32'h416ebbb2};
test_output[1156:1156] = '{32'hc50e6a4d};
test_input[9256:9263] = '{32'hc29b7c44, 32'hc1807c75, 32'h42a6fce5, 32'h42c3efbe, 32'hc07e07de, 32'h41fc886b, 32'h41440cd8, 32'h42c436cd};
test_weights[9256:9263] = '{32'h41feeae8, 32'h427b290c, 32'h42c63eca, 32'hbff9bc60, 32'h42938882, 32'hc29a28d9, 32'h3f2ebf65, 32'hc0f6c594};
test_bias[1157:1157] = '{32'h42809e07};
test_output[1157:1157] = '{32'h4494ae9b};
test_input[9264:9271] = '{32'hc2c35602, 32'hc20b03b3, 32'h41ccc3f7, 32'hc25efd09, 32'h42a1d11c, 32'hc1e30d60, 32'h42c529fb, 32'h429562a2};
test_weights[9264:9271] = '{32'h410bfa55, 32'h41819801, 32'hc1658f11, 32'h42981a13, 32'hc2bb8f24, 32'hc15e4e5c, 32'hc297e93d, 32'h41d669d4};
test_bias[1158:1158] = '{32'hc27e05d8};
test_output[1158:1158] = '{32'hc6929df5};
test_input[9272:9279] = '{32'h403758c9, 32'h4294781a, 32'hc0189afb, 32'h41ebe889, 32'hc13bbaa4, 32'h4278b11a, 32'hc1e06c71, 32'hc2c427bc};
test_weights[9272:9279] = '{32'h42642874, 32'h41a338dc, 32'hc2b0ca67, 32'h42c07b1b, 32'h4183139d, 32'hc2a37d2e, 32'hc108a3a6, 32'h42935e57};
test_bias[1159:1159] = '{32'h415d2fa0};
test_output[1159:1159] = '{32'hc5eb093f};
test_input[9280:9287] = '{32'h3fa45e6e, 32'h41ef25ac, 32'h3f5acfdb, 32'h42566f96, 32'h416d53ae, 32'hc2a05635, 32'hc236aa90, 32'hc1596cc7};
test_weights[9280:9287] = '{32'h40cabe29, 32'h4111fbb8, 32'hc2be202b, 32'hc220583d, 32'hc0daabc7, 32'hc2a38a35, 32'hc21cb5e8, 32'hc1666f62};
test_bias[1160:1160] = '{32'h428d0bd0};
test_output[1160:1160] = '{32'h45ccfff8};
test_input[9288:9295] = '{32'hc2b3d228, 32'hc11d0efb, 32'h4286f5fe, 32'h41d6563b, 32'hc1fdb9a9, 32'h4295be7b, 32'hc2b2cd3b, 32'h41d32134};
test_weights[9288:9295] = '{32'h41636d74, 32'hc2aab895, 32'hc1dfab86, 32'hc29c028d, 32'hc220080b, 32'hc2c7c84a, 32'hc1bee31c, 32'hc28e0813};
test_bias[1161:1161] = '{32'hc2c341d4};
test_output[1161:1161] = '{32'hc6238600};
test_input[9296:9303] = '{32'hc2b4c2d3, 32'hc1f989e3, 32'h420d668d, 32'h4214829f, 32'hc17945fd, 32'h42ad8a8d, 32'h42850dc0, 32'h41e5d7ee};
test_weights[9296:9303] = '{32'h429af3c4, 32'hc1b9fcbf, 32'h42a50d0a, 32'hc29e2877, 32'h4249ab4e, 32'hc29f9fcb, 32'hc1980fb6, 32'hc1c146ac};
test_bias[1162:1162] = '{32'h41a1dcfc};
test_output[1162:1162] = '{32'hc679246f};
test_input[9304:9311] = '{32'h41165e33, 32'hc175b204, 32'h425e574a, 32'hbf6fcbe9, 32'hc2304645, 32'hc09bcb3a, 32'hc2b3ab3b, 32'hc0fa70ef};
test_weights[9304:9311] = '{32'hc159ed62, 32'h42845796, 32'hc2a847be, 32'h42b487d4, 32'hc14b0217, 32'hc28d0f5b, 32'h42a6bf15, 32'h42018c3a};
test_bias[1163:1163] = '{32'hc2b05a4a};
test_output[1163:1163] = '{32'hc6488a24};
test_input[9312:9319] = '{32'hc0c21078, 32'h42764a25, 32'hc1503d57, 32'h42967fe1, 32'hc273dba2, 32'hc23308ee, 32'h41da7b78, 32'h41d707be};
test_weights[9312:9319] = '{32'hc18248d7, 32'hc1d6f09b, 32'h4132229d, 32'hc293cef6, 32'h429977d7, 32'hc08889e9, 32'h4259548d, 32'hc249ed07};
test_bias[1164:1164] = '{32'hc0c03db8};
test_output[1164:1164] = '{32'hc635af55};
test_input[9320:9327] = '{32'h41d4bd8d, 32'hc29bbaaf, 32'h4265bb6a, 32'hc165df98, 32'h42478bc9, 32'hc245c263, 32'hc2228c39, 32'h423c9a4e};
test_weights[9320:9327] = '{32'hc2b391c4, 32'hc22d4ec0, 32'hc262e642, 32'hc23a8cc3, 32'hc2c02b4f, 32'h41d8ecd8, 32'h41db60e3, 32'h4289a16e};
test_bias[1165:1165] = '{32'h412a5955};
test_output[1165:1165] = '{32'hc5aed5fc};
test_input[9328:9335] = '{32'hc1e9d60b, 32'hc26d7e8b, 32'hc29cabc2, 32'hc2c3042b, 32'h42bbbf31, 32'hc2c2c384, 32'h42388ea0, 32'hc29f7fc0};
test_weights[9328:9335] = '{32'h41fc9388, 32'h42917820, 32'h429e1a96, 32'h42a7e4b7, 32'h41ea4682, 32'hbfa99e5e, 32'hc2664620, 32'h4286bc35};
test_bias[1166:1166] = '{32'hc2183284};
test_output[1166:1166] = '{32'hc6c1d02b};
test_input[9336:9343] = '{32'h4297117f, 32'h42c43acf, 32'h41948fa1, 32'h42468d33, 32'hc02cc6b0, 32'h4236f8d5, 32'hc26d40c0, 32'h42ad1e64};
test_weights[9336:9343] = '{32'h42aa849b, 32'h427685de, 32'hc1c05beb, 32'h41d8d077, 32'h42b9e79f, 32'hc1b97a14, 32'hc2a7fec2, 32'hc1d5f326};
test_bias[1167:1167] = '{32'h42993dbf};
test_output[1167:1167] = '{32'h4667880f};
test_input[9344:9351] = '{32'h41f90669, 32'h424ac4be, 32'hc2978a62, 32'h41ff3540, 32'h42ac4377, 32'hc1f79316, 32'hc26eef9e, 32'hc15aa711};
test_weights[9344:9351] = '{32'h4217f872, 32'h41a44d88, 32'hc1debfa0, 32'h4132ff16, 32'hc233c438, 32'h3fc68e6e, 32'hc1f3117f, 32'h42a66227};
test_bias[1168:1168] = '{32'hbfa42095};
test_output[1168:1168] = '{32'h44b506ad};
test_input[9352:9359] = '{32'hc2b1561b, 32'h4238256f, 32'hc296c336, 32'h429fbc76, 32'h4212dd0e, 32'hc2368959, 32'hc1e199aa, 32'h41ead8a0};
test_weights[9352:9359] = '{32'h42b5f83d, 32'h42bfb444, 32'hc2031e2a, 32'h429d9b82, 32'hc24a34b8, 32'hc282a0e4, 32'hc22f800f, 32'hc29ff393};
test_bias[1169:1169] = '{32'h42b279d6};
test_output[1169:1169] = '{32'h45a2eb12};
test_input[9360:9367] = '{32'h420a70cc, 32'h42956e7c, 32'h4294f4aa, 32'h409e0245, 32'hc2426f72, 32'h4228cd62, 32'h420640f1, 32'hc195d5a0};
test_weights[9360:9367] = '{32'h429f6501, 32'hc28d52df, 32'h424fd18d, 32'h428b40ee, 32'h42bf4947, 32'h428dff25, 32'h4288fd24, 32'h42b40b99};
test_bias[1170:1170] = '{32'h424a663d};
test_output[1170:1170] = '{32'h442fa423};
test_input[9368:9375] = '{32'hc2afa26b, 32'h3fe02a81, 32'hc1f0c985, 32'hc1b3ca13, 32'hc2b3d5a7, 32'h4078176b, 32'hc17d19ac, 32'h41f87f66};
test_weights[9368:9375] = '{32'h42baf1c1, 32'h427878c0, 32'hc2bf2c40, 32'h4218723e, 32'hc267cfb1, 32'hc21beb47, 32'h41dbfcfb, 32'h42c12b3a};
test_bias[1171:1171] = '{32'h4224e214};
test_output[1171:1171] = '{32'h44c660c0};
test_input[9376:9383] = '{32'hc29c29a0, 32'hc1da7927, 32'h42a599d4, 32'h42bfe8e9, 32'hc2b7c633, 32'h420c4af2, 32'hc2285d4e, 32'hc2aa6e01};
test_weights[9376:9383] = '{32'h424d4832, 32'hc1fbf589, 32'hc25d6a48, 32'hc22f7671, 32'hc1b85fb7, 32'hc2baa966, 32'hc1f0c3db, 32'h42a548aa};
test_bias[1172:1172] = '{32'hc2078a17};
test_output[1172:1172] = '{32'hc693b15a};
test_input[9384:9391] = '{32'hc2766ca1, 32'h42aa8d99, 32'hc1548dd2, 32'hc29b4b15, 32'hc29d5bb8, 32'h410df519, 32'hc2a095bc, 32'h419f8374};
test_weights[9384:9391] = '{32'h4284ff4b, 32'h41c01460, 32'h42806770, 32'hc2bf71f3, 32'h40e34285, 32'h423973bb, 32'hc2af4d6d, 32'h4114ce81};
test_bias[1173:1173] = '{32'hc2aac11b};
test_output[1173:1173] = '{32'h4634031d};
test_input[9392:9399] = '{32'hc27ded61, 32'h41cb42e2, 32'hc16d6348, 32'h4289a3af, 32'h4221be57, 32'hc1b61b71, 32'h42c19b9f, 32'h421c02b9};
test_weights[9392:9399] = '{32'h42b4db3c, 32'h42339e78, 32'hc1b45233, 32'h41423946, 32'hc24f2fe0, 32'hc12cbbd5, 32'h42b2fccc, 32'hc270bcb0};
test_bias[1174:1174] = '{32'h42973dff};
test_output[1174:1174] = '{32'h448b2412};
test_input[9400:9407] = '{32'h42b2a6a0, 32'hc2135146, 32'h415faf8b, 32'hc29f7849, 32'h42a64cb8, 32'hc2ab2e12, 32'hc24686e3, 32'hc2437973};
test_weights[9400:9407] = '{32'hc196bb76, 32'h428070f2, 32'h4154ab47, 32'h41971b2c, 32'h427fc41c, 32'h4294865f, 32'hc2b2eea1, 32'h40c3fde3};
test_bias[1175:1175] = '{32'h42b79861};
test_output[1175:1175] = '{32'hc507f030};
test_input[9408:9415] = '{32'h42864a96, 32'hc2b8a4c4, 32'h426ec103, 32'hc22fcc98, 32'hc2a0486e, 32'hc291b4a9, 32'h42ad1051, 32'hc1d698df};
test_weights[9408:9415] = '{32'hc18105f9, 32'hc2221221, 32'hc1a3d584, 32'h426712bf, 32'h42252726, 32'h421a8762, 32'hc1b8a8fc, 32'hc18facc9};
test_bias[1176:1176] = '{32'h426c78a7};
test_output[1176:1176] = '{32'hc607ad9a};
test_input[9416:9423] = '{32'h42bdef94, 32'h40b35939, 32'hc1a57c87, 32'hc2197129, 32'h42c55aa6, 32'h42a4ef8e, 32'h41800595, 32'hc29d6c70};
test_weights[9416:9423] = '{32'h417b9970, 32'h4124d550, 32'hc2a3e81f, 32'hc1f7d7d7, 32'h41cfea55, 32'h422b6303, 32'h412f1ca2, 32'h42548db4};
test_bias[1177:1177] = '{32'h428a2ca8};
test_output[1177:1177] = '{32'h45ce1395};
test_input[9424:9431] = '{32'h42ac4274, 32'h4246da38, 32'hc035b15e, 32'hc2a4dc7a, 32'h42b73d17, 32'hc296ec05, 32'hc1d68693, 32'hbe7fa039};
test_weights[9424:9431] = '{32'hc2b2383a, 32'h42c58be4, 32'h41bdb747, 32'hc284fa1c, 32'hc267f8cf, 32'h425c02bf, 32'h426e3be4, 32'h41900592};
test_bias[1178:1178] = '{32'h42388756};
test_output[1178:1178] = '{32'hc602ca7b};
test_input[9432:9439] = '{32'hc28a05d4, 32'h4012deda, 32'h428de45b, 32'hc18ef90f, 32'hc2aa7d8d, 32'hc1d89b55, 32'h404f57d3, 32'hc1b37d68};
test_weights[9432:9439] = '{32'hc2038c60, 32'h42becdfe, 32'hc20e62e0, 32'h4238d517, 32'h42abfffb, 32'hc2007a2a, 32'hc0ea7797, 32'h41987504};
test_bias[1179:1179] = '{32'h42825c14};
test_output[1179:1179] = '{32'hc5f0f24a};
test_input[9440:9447] = '{32'h411a94bd, 32'hc28ba445, 32'h41b7e5d7, 32'h4241d957, 32'hc29264e2, 32'h41be66b8, 32'hc2740fe3, 32'h42a8d1f2};
test_weights[9440:9447] = '{32'h425f5faa, 32'hc24d1bc7, 32'hc29027d3, 32'h40ff5df1, 32'hc26024b9, 32'hc224e59e, 32'hc1b2683c, 32'h429e83e7};
test_bias[1180:1180] = '{32'hc2be992d};
test_output[1180:1180] = '{32'h465996a5};
test_input[9448:9455] = '{32'hc1f2a4ef, 32'hc24f8a01, 32'h41883acb, 32'h428844bd, 32'hc1ab29fd, 32'hc2631411, 32'hc2837b79, 32'h42b8cdc9};
test_weights[9448:9455] = '{32'h4253791c, 32'hc283e47c, 32'hc266f963, 32'hc20d4c02, 32'hc2b06077, 32'hc25d86d6, 32'h4216ec15, 32'hc2723a5d};
test_bias[1181:1181] = '{32'hbf562785};
test_output[1181:1181] = '{32'hc5905058};
test_input[9456:9463] = '{32'h423aad3f, 32'hc21396cf, 32'hc1a51c0f, 32'hc193360f, 32'h42a580e0, 32'hc2b7a8d2, 32'h424053df, 32'h41136697};
test_weights[9456:9463] = '{32'hc2576f6a, 32'h429cc97e, 32'hc1d969a9, 32'hc2bd63e4, 32'h42b8ccf2, 32'hc29d60dd, 32'hc2c3d484, 32'h42c56a22};
test_bias[1182:1182] = '{32'h4283e4df};
test_output[1182:1182] = '{32'h45fb27f5};
test_input[9464:9471] = '{32'h42b3426f, 32'hc16488bd, 32'hc2b97bd1, 32'hc2aca170, 32'hc2458445, 32'hc1bfe24e, 32'h4110e8f0, 32'hc206e79c};
test_weights[9464:9471] = '{32'h41ccaf57, 32'hc29c6e1c, 32'hc27bef9d, 32'hc1c33eeb, 32'h41542194, 32'hc28a7943, 32'h410ebe28, 32'hc22b738a};
test_bias[1183:1183] = '{32'hc1db2efe};
test_output[1183:1183] = '{32'h46589d00};
test_input[9472:9479] = '{32'h427d0fbf, 32'h41cb5313, 32'hc274b64c, 32'h42bc321f, 32'hc1fb9322, 32'hc1cb1385, 32'hc21f656b, 32'hc1c4e10a};
test_weights[9472:9479] = '{32'h419dacb9, 32'hc24f4b99, 32'hc22c0015, 32'hc20a92d8, 32'hc10ca84f, 32'hc2ac997b, 32'hc282e581, 32'hc13809ae};
test_bias[1184:1184] = '{32'hc29360dd};
test_output[1184:1184] = '{32'h458f491e};
test_input[9480:9487] = '{32'h40764af9, 32'hc2a1e24b, 32'h4274a227, 32'hc252db63, 32'h42c19709, 32'h428efc00, 32'hc07f9f6c, 32'hc20eff06};
test_weights[9480:9487] = '{32'h4249f576, 32'h42ab4300, 32'hc19c6020, 32'h41da3607, 32'h428fd7de, 32'h422e9103, 32'hc1f208ee, 32'h42b39dd6};
test_bias[1185:1185] = '{32'hc21402bb};
test_output[1185:1185] = '{32'hc516f2e2};
test_input[9488:9495] = '{32'h4011f67e, 32'h41d55d13, 32'hc2825432, 32'h42b70bf2, 32'hc237794a, 32'hc2c2c427, 32'h42c1c1ea, 32'hc13b2d6b};
test_weights[9488:9495] = '{32'h4228770c, 32'hc22ce263, 32'h423ff476, 32'h424def00, 32'hc27876c1, 32'h4231f35c, 32'hc2c24d08, 32'hc2978497};
test_bias[1186:1186] = '{32'hc2621a88};
test_output[1186:1186] = '{32'hc6150499};
test_input[9496:9503] = '{32'h41104113, 32'h42b7cc5f, 32'h4236fcf7, 32'hc28099d1, 32'hc2a044ad, 32'h41cda22b, 32'h42bf6fda, 32'hc26dbae9};
test_weights[9496:9503] = '{32'hc28ea64a, 32'h42252399, 32'hc230776f, 32'h42c36db7, 32'hc0a9176b, 32'h4285f222, 32'h420270f4, 32'hc2c1f4a8};
test_bias[1187:1187] = '{32'h42b8b03d};
test_output[1187:1187] = '{32'h45baa021};
test_input[9504:9511] = '{32'h42a35c81, 32'h42b3497c, 32'hc0beb08d, 32'h41038ce9, 32'h424a0dc8, 32'h4295eb53, 32'hc1941a51, 32'h41ac241d};
test_weights[9504:9511] = '{32'hc233a2ac, 32'h421f1828, 32'h42b70bbe, 32'hc20a2f9f, 32'h41006d6f, 32'hc2083705, 32'hc2b72124, 32'hc28cf515};
test_bias[1188:1188] = '{32'h427c78c3};
test_output[1188:1188] = '{32'hc5315a87};
test_input[9512:9519] = '{32'hc2ad36d1, 32'h42058304, 32'hc2624e82, 32'hc104b81e, 32'hc23ded08, 32'h4289aea4, 32'hc204f46e, 32'h428d3402};
test_weights[9512:9519] = '{32'hc26e49f9, 32'hc1dc70ef, 32'h4286e0a3, 32'h42afd397, 32'hc289c136, 32'h426d25e0, 32'hc2754c2b, 32'h42876e31};
test_bias[1189:1189] = '{32'hc226d78f};
test_output[1189:1189] = '{32'h465800a5};
test_input[9520:9527] = '{32'h42c531ff, 32'h42c6d62f, 32'hc24d172e, 32'hc1fe56f4, 32'hc2998876, 32'h4295e6c6, 32'hc2468528, 32'h4293426f};
test_weights[9520:9527] = '{32'h4204df5e, 32'h419ba329, 32'h424b5530, 32'h41c94751, 32'hc2a05225, 32'hc25a5e95, 32'hc1a6a5b6, 32'hc23395f6};
test_bias[1190:1190] = '{32'hc221f931};
test_output[1190:1190] = '{32'h44c2155f};
test_input[9528:9535] = '{32'h42a39987, 32'h420f11b6, 32'h410ca89d, 32'hc2b714bc, 32'h423f5e94, 32'h42b49e5c, 32'hc294c5d9, 32'hc2b18063};
test_weights[9528:9535] = '{32'h42aab6c9, 32'h416942b9, 32'hc292ed6b, 32'h424a6945, 32'h4298fe52, 32'h4288a65c, 32'hc1bb2055, 32'hc2b59c82};
test_bias[1191:1191] = '{32'h42a88fd0};
test_output[1191:1191] = '{32'h46ab6622};
test_input[9536:9543] = '{32'hc294c632, 32'hc244393d, 32'h42ad2f8d, 32'hc1d1cd56, 32'h4297e67a, 32'hc2390f31, 32'h42213ec8, 32'hc2a66c95};
test_weights[9536:9543] = '{32'h4078c4d0, 32'hc256a183, 32'hc246cfbc, 32'hc2616aec, 32'hc2a84121, 32'h4235556c, 32'hc1f949c1, 32'h41fbee76};
test_bias[1192:1192] = '{32'hc0cd5120};
test_output[1192:1192] = '{32'hc648d30d};
test_input[9544:9551] = '{32'hc2650732, 32'hc1846b07, 32'hc216b4cc, 32'h416e2ccc, 32'h42bda085, 32'h420e12aa, 32'hc1c89d4d, 32'h40b51e90};
test_weights[9544:9551] = '{32'h4173f125, 32'h41166baa, 32'h42901770, 32'h4192e026, 32'h41f80fa1, 32'h4286322d, 32'hc0c5db47, 32'h4291c50b};
test_bias[1193:1193] = '{32'h4293c766};
test_output[1193:1193] = '{32'h451bee5b};
test_input[9552:9559] = '{32'hc13832d4, 32'hc27deb92, 32'hc2b20e8d, 32'hc2331568, 32'h3fc0853a, 32'hc233608e, 32'hc206f472, 32'h4203753b};
test_weights[9552:9559] = '{32'h42162d8e, 32'hc23a880d, 32'hc2c289fd, 32'hc2c29559, 32'hc2a6b4e0, 32'hc05f3ea6, 32'h42a641cc, 32'hc29d0365};
test_bias[1194:1194] = '{32'hc246905d};
test_output[1194:1194] = '{32'h461e7137};
test_input[9560:9567] = '{32'hc29cc234, 32'h41d4856c, 32'hc2113f0c, 32'hc0afef4e, 32'h41a1ae4d, 32'h4204a5d4, 32'h426ea115, 32'h42b40ed4};
test_weights[9560:9567] = '{32'h41d5ec90, 32'h427636cd, 32'h42a00d13, 32'hc29b7c8e, 32'h42a0d744, 32'hbf48e9e5, 32'hc2c1257c, 32'hc22ad632};
test_bias[1195:1195] = '{32'h42c5ccbd};
test_output[1195:1195] = '{32'hc6297d50};
test_input[9568:9575] = '{32'h41254bd1, 32'h41c4aff0, 32'h42c46076, 32'h429bf4ff, 32'hc0758fcb, 32'h4132cc7a, 32'hc26adfb0, 32'h40bf25f0};
test_weights[9568:9575] = '{32'hc1e421a9, 32'h4219364b, 32'h428e2630, 32'hc202bafe, 32'h4216b62f, 32'h4286f209, 32'hc2153aa8, 32'hc2730d54};
test_bias[1196:1196] = '{32'hc2a86520};
test_output[1196:1196] = '{32'h45e83162};
test_input[9576:9583] = '{32'h41fb895f, 32'hc10d9374, 32'h42c3d933, 32'h42214771, 32'hc1198626, 32'hc1f9c2e5, 32'h4291aee5, 32'h42a68e69};
test_weights[9576:9583] = '{32'hc2c4203c, 32'hc106ed12, 32'h4247a56f, 32'h40cf3c8e, 32'hc1eb1995, 32'hc1927c89, 32'hc2bbb474, 32'h429b3462};
test_bias[1197:1197] = '{32'h420e8c50};
test_output[1197:1197] = '{32'h4525f7af};
test_input[9584:9591] = '{32'hc2299a94, 32'hbfb1941c, 32'hc24ae9a6, 32'hc2b7749c, 32'h40cd80fc, 32'h426cae77, 32'hc1bdb011, 32'hc1817d83};
test_weights[9584:9591] = '{32'h4229ae51, 32'h41410ee0, 32'hc2b07d64, 32'h417acc4a, 32'h42c385bf, 32'hc26a3ebb, 32'h42bbf1ae, 32'h42188f62};
test_bias[1198:1198] = '{32'h426e1d22};
test_output[1198:1198] = '{32'hc5897fc4};
test_input[9592:9599] = '{32'hc1e094c4, 32'hbfbf6d03, 32'hc282b983, 32'h41da134c, 32'hc111127d, 32'hc2c5f6a2, 32'hc0871a96, 32'h429899bc};
test_weights[9592:9599] = '{32'h41a5d630, 32'h421c747c, 32'h429b7bf5, 32'hc2264d95, 32'h42afcb66, 32'hc19b3ab3, 32'hc1cee9b7, 32'h42bc1bf7};
test_bias[1199:1199] = '{32'hc2872e5b};
test_output[1199:1199] = '{32'h44b9cf3d};
test_input[9600:9607] = '{32'hc1b45195, 32'h41c4cfb6, 32'hc2a9c177, 32'h42a84fe2, 32'h4028856f, 32'h42c3baee, 32'h41de3980, 32'h42356635};
test_weights[9600:9607] = '{32'hc2619931, 32'hc1624f77, 32'h42607443, 32'hc211da67, 32'hc28043b1, 32'hc2730000, 32'h429d1112, 32'hc196b191};
test_bias[1200:1200] = '{32'h42c30a65};
test_output[1200:1200] = '{32'hc635361a};
test_input[9608:9615] = '{32'hc206d560, 32'h42102d62, 32'h42b6ac95, 32'h41f30580, 32'hc296b069, 32'hc2432941, 32'hc182c207, 32'hc1f0ed2a};
test_weights[9608:9615] = '{32'hc29a8e76, 32'h42939cf8, 32'h41134e45, 32'hc2c7d313, 32'hc006fb27, 32'h4248c5d0, 32'hc283d4b8, 32'hc2a4e4d6};
test_bias[1201:1201] = '{32'h40b93495};
test_output[1201:1201] = '{32'h4587d8ef};
test_input[9616:9623] = '{32'h428f58c6, 32'h4222236f, 32'hc27a7fcb, 32'hc1d13775, 32'h428d7223, 32'hc18fc4b3, 32'h42895376, 32'h41ff0027};
test_weights[9616:9623] = '{32'h423faeef, 32'hc22735ce, 32'hc29727e1, 32'hc2a19746, 32'h41b8c7f4, 32'h4154831f, 32'h40dad9d2, 32'hc2a4ac49};
test_bias[1202:1202] = '{32'h4274fff6};
test_output[1202:1202] = '{32'h45f67b5a};
test_input[9624:9631] = '{32'hc1e3be0e, 32'hc18c7144, 32'h423c4747, 32'hc248750f, 32'hc269a801, 32'hc27a473e, 32'h40530c0c, 32'hc2203597};
test_weights[9624:9631] = '{32'h42239129, 32'h427336b1, 32'h4240925a, 32'hc2911bc0, 32'h41836bf3, 32'hc23255b1, 32'hc2ba38a0, 32'hc2160150};
test_bias[1203:1203] = '{32'hc253e0fb};
test_output[1203:1203] = '{32'h45cf9435};
test_input[9632:9639] = '{32'h41b420f9, 32'h41c6e2ba, 32'h40de1815, 32'hc1262185, 32'h41d5425d, 32'h424f9dfe, 32'hc21d69da, 32'h422fafcc};
test_weights[9632:9639] = '{32'h4267b58f, 32'hc1a0a9f1, 32'hc2a92c08, 32'hc27e0a75, 32'h429c184c, 32'h429ec8a5, 32'hc2c5729a, 32'hc28592f0};
test_bias[1204:1204] = '{32'h41fd6b58};
test_output[1204:1204] = '{32'h45fbf0e7};
test_input[9640:9647] = '{32'hc23d35d7, 32'hc2a713a8, 32'h42b1be2b, 32'h421520cf, 32'hc2a207a3, 32'hc1dc134b, 32'h414b8814, 32'hc1b4c3ff};
test_weights[9640:9647] = '{32'h42b892fc, 32'h4295901d, 32'h428de86c, 32'hc2a0c466, 32'hc2209780, 32'hc20b8518, 32'h4268593d, 32'h42463bb7};
test_bias[1205:1205] = '{32'h423b50a9};
test_output[1205:1205] = '{32'hc5561950};
test_input[9648:9655] = '{32'h42a35607, 32'h4168d076, 32'hc29a8792, 32'hc19a2632, 32'h4266ecf5, 32'h424ef739, 32'hc26faa5f, 32'h428f9556};
test_weights[9648:9655] = '{32'hc2a44b29, 32'h4161095e, 32'hc2ace6b9, 32'hbf9d1413, 32'h40b79403, 32'h42a7460c, 32'h4201a0e4, 32'hc287e60f};
test_bias[1206:1206] = '{32'h42200d63};
test_output[1206:1206] = '{32'hc4f042fd};
test_input[9656:9663] = '{32'h40d48f9d, 32'h42044027, 32'hc2af8261, 32'hc23ea608, 32'h42423367, 32'h42c4df69, 32'h427c94db, 32'hc29649dd};
test_weights[9656:9663] = '{32'h4225d225, 32'h42b8441c, 32'hc1eea8c9, 32'hc20c6590, 32'h4078c60e, 32'h425fff4b, 32'h426ec00d, 32'hc207eb57};
test_bias[1207:1207] = '{32'hc125a39e};
test_output[1207:1207] = '{32'h469952f5};
test_input[9664:9671] = '{32'h429666a5, 32'hc26b2faf, 32'hc20077eb, 32'h42ba1769, 32'hc1b33327, 32'h42b9093c, 32'h42844839, 32'h42684117};
test_weights[9664:9671] = '{32'h422bc543, 32'h42a1a32d, 32'h42990a6f, 32'h42c6d03a, 32'h42879129, 32'hc24c18f8, 32'h42c78b27, 32'hc291e60d};
test_bias[1208:1208] = '{32'hc27abb79};
test_output[1208:1208] = '{32'h44a659c3};
test_input[9672:9679] = '{32'hc2c11b3c, 32'hc1b55ce6, 32'h42837dea, 32'hc1ee6518, 32'h4253a8bc, 32'hc29bf4a3, 32'hc27cb2b0, 32'h411a71d7};
test_weights[9672:9679] = '{32'h418329db, 32'hc27abc14, 32'h42933da0, 32'h4044c506, 32'h424a1be7, 32'h423ff625, 32'hc1aabb42, 32'hc2c2b4cb};
test_bias[1209:1209] = '{32'h4196a59d};
test_output[1209:1209] = '{32'h45769709};
test_input[9680:9687] = '{32'hc20d620f, 32'hc16bd31b, 32'h428ba76e, 32'hc1953742, 32'h428f102b, 32'hc2c2cc54, 32'hc18e421b, 32'h42c0cfaa};
test_weights[9680:9687] = '{32'h42383493, 32'hc2c60d31, 32'hc28041a0, 32'hc20c2231, 32'hc1b3ed58, 32'h41c8c1fb, 32'hc2be4d2a, 32'hc2bc03b6};
test_bias[1210:1210] = '{32'hc2bc127a};
test_output[1210:1210] = '{32'hc67259f2};
test_input[9688:9695] = '{32'h42857319, 32'hc27a7847, 32'h42357cc1, 32'h41c3f5a3, 32'hc2b44a95, 32'h427c77b1, 32'h41056afa, 32'h412c76e0};
test_weights[9688:9695] = '{32'hc2165bbe, 32'hc28b84a9, 32'hc23cb60d, 32'hbf872016, 32'h4272f3d3, 32'hc23c6c7c, 32'h3f89a41a, 32'h41cd64ad};
test_bias[1211:1211] = '{32'hc0c6f10c};
test_output[1211:1211] = '{32'hc6046d8c};
test_input[9696:9703] = '{32'h42b1d86a, 32'h42aa9040, 32'hc21165f4, 32'h42b98813, 32'hc156f628, 32'h4250b06d, 32'hc05b2a16, 32'h42c7309e};
test_weights[9696:9703] = '{32'hc25ce2e5, 32'hc1ee8f8c, 32'h42b49f19, 32'hc2275a8e, 32'hc13f698d, 32'h414d3c51, 32'h4289351b, 32'h42079be3};
test_bias[1212:1212] = '{32'hc250f319};
test_output[1212:1212] = '{32'hc62728da};
test_input[9704:9711] = '{32'h40dfdd61, 32'h4249b9f4, 32'hc2468c19, 32'hc224d15e, 32'h42a19238, 32'h41ee8195, 32'hc24f526e, 32'hc2800f76};
test_weights[9704:9711] = '{32'h41eaa806, 32'h41acd507, 32'h40fdf3fe, 32'hc1d0f3d4, 32'hc2488927, 32'h428f7845, 32'hc1876bd6, 32'h42c43304};
test_bias[1213:1213] = '{32'hc2bcd9da};
test_output[1213:1213] = '{32'hc5a9c687};
test_input[9712:9719] = '{32'h42bbe5d1, 32'hc2689d36, 32'h4232b535, 32'h414e87b2, 32'hc27f9f58, 32'hc23aeb49, 32'hc1b5ad98, 32'hc2b4268c};
test_weights[9712:9719] = '{32'h413ae129, 32'h42be89f8, 32'h425b017a, 32'hc29506df, 32'h418ab49c, 32'h4226c8c5, 32'h4207d653, 32'hc1aaacaf};
test_bias[1214:1214] = '{32'h405a72da};
test_output[1214:1214] = '{32'hc597e987};
test_input[9720:9727] = '{32'h41de91ad, 32'h423723ad, 32'h41e7c227, 32'h42818426, 32'hc2b0e79f, 32'h4275e480, 32'hc0ae0c83, 32'h429988f0};
test_weights[9720:9727] = '{32'h417298fa, 32'hc1e1992e, 32'h41a70499, 32'hc2a88ed7, 32'h42615b6a, 32'hc2bae4bc, 32'h4231e4aa, 32'hc01734b8};
test_bias[1215:1215] = '{32'h42711129};
test_output[1215:1215] = '{32'hc6835a0f};
test_input[9728:9735] = '{32'h42b5bc12, 32'hc294d570, 32'hc16a859d, 32'h4282de86, 32'hc20d6be4, 32'hc10aba44, 32'h428c2c84, 32'hc1c0fb5c};
test_weights[9728:9735] = '{32'hc268d676, 32'h421ec743, 32'hc2156989, 32'hc1c79583, 32'hc203fb07, 32'hc0cff81a, 32'hc29d70ef, 32'hc2ba156b};
test_bias[1216:1216] = '{32'h429d74b6};
test_output[1216:1216] = '{32'hc6308dde};
test_input[9736:9743] = '{32'hc27b1a4b, 32'hc2985101, 32'h42b8cea3, 32'h426b9ba9, 32'hc211bfe3, 32'hc2b79d55, 32'h41833d2d, 32'h40d69f8c};
test_weights[9736:9743] = '{32'hc09f96c7, 32'hc1c9be04, 32'h4085cb24, 32'hc27f1bb9, 32'hc296a16f, 32'hc21c0d20, 32'hc2111433, 32'h42a41791};
test_bias[1217:1217] = '{32'h42895dad};
test_output[1217:1217] = '{32'h45a2ea37};
test_input[9744:9751] = '{32'hc28ae53d, 32'h429d26e5, 32'hc1f2bbd2, 32'hc2aac38f, 32'hc2b36161, 32'h40e1ffdd, 32'h423c6382, 32'h42a42ed8};
test_weights[9744:9751] = '{32'h423f940e, 32'h4292ae34, 32'h427d3f74, 32'h4280c0d8, 32'h416f9f75, 32'hc25ec993, 32'h412479dc, 32'hc2bc5846};
test_bias[1218:1218] = '{32'h429bacfe};
test_output[1218:1218] = '{32'hc658f969};
test_input[9752:9759] = '{32'h40c9542a, 32'h42b71223, 32'hc295cc7b, 32'hc27d672d, 32'h42b1e362, 32'h4277f8bb, 32'hc2870743, 32'hc29b4e62};
test_weights[9752:9759] = '{32'h41e6b2bf, 32'h42a9db87, 32'h420543cc, 32'h42b10405, 32'hc262a45d, 32'h411d073c, 32'h42b337c6, 32'h427d8799};
test_bias[1219:1219] = '{32'h4239c0c0};
test_output[1219:1219] = '{32'hc6723dda};
test_input[9760:9767] = '{32'hc28bb4bf, 32'hc2978761, 32'hc2654709, 32'hc2046305, 32'hc0969bae, 32'h405080b5, 32'hc22edc2c, 32'h3fc733c1};
test_weights[9760:9767] = '{32'h41f1d037, 32'hc184b610, 32'hc0a251f0, 32'h4234b6f2, 32'h4266ad96, 32'hc2b71fbc, 32'h4248f5c3, 32'h411a8056};
test_bias[1220:1220] = '{32'h42995aaf};
test_output[1220:1220] = '{32'hc593eabe};
test_input[9768:9775] = '{32'hc275692c, 32'hc20cd90d, 32'h411d7253, 32'hc2a10743, 32'h428601bd, 32'h4262a149, 32'hc2329514, 32'h4283f216};
test_weights[9768:9775] = '{32'hc20e9d65, 32'h413e6c0d, 32'hc1d7bb8a, 32'h4195783c, 32'h419cc1a2, 32'hc2638ed0, 32'hc1c18e29, 32'h42bbfd14};
test_bias[1221:1221] = '{32'hc208759c};
test_output[1221:1221] = '{32'h45a6bc3a};
test_input[9776:9783] = '{32'hc227f1cb, 32'hc26933f8, 32'h42a22988, 32'h42be532e, 32'hc2886ba4, 32'hc1444147, 32'h40fba500, 32'hc2754c7b};
test_weights[9776:9783] = '{32'h414a45fc, 32'hc2a3f43c, 32'hc23c6a4f, 32'hc22c4e6d, 32'hc1bd09eb, 32'h427f002f, 32'hc16dff4c, 32'hc284ed7c};
test_bias[1222:1222] = '{32'h42b3f602};
test_output[1222:1222] = '{32'h449717ec};
test_input[9784:9791] = '{32'hc2ad4cb9, 32'hbfcffafe, 32'hc2799ac5, 32'h420724c3, 32'h420e566b, 32'h40fc4b77, 32'hc1953739, 32'hc0c1ff60};
test_weights[9784:9791] = '{32'h42bf12ff, 32'h421349ee, 32'h423853b7, 32'hc192a176, 32'hc29f4c7d, 32'hc1b513b1, 32'hc2ad18ea, 32'h41afd56a};
test_bias[1223:1223] = '{32'hc25eb5c4};
test_output[1223:1223] = '{32'hc651b114};
test_input[9792:9799] = '{32'hc0ae15cf, 32'hc239d5c9, 32'hc190a656, 32'hc22ade02, 32'h4188c59e, 32'hc2c22450, 32'h41437f2a, 32'hc222e82a};
test_weights[9792:9799] = '{32'h41cdff1d, 32'h41ea953a, 32'hc2a11bbb, 32'h42aeb3c9, 32'hc120b7a4, 32'h415e938d, 32'h41e55930, 32'hc2c47ef5};
test_bias[1224:1224] = '{32'hc2bb8065};
test_output[1224:1224] = '{32'hc4822ed2};
test_input[9800:9807] = '{32'hc298d1f4, 32'hc28d8365, 32'hc2c39051, 32'hc29fb291, 32'h422618f4, 32'hc25b1aca, 32'h4182ee1b, 32'h41d1209a};
test_weights[9800:9807] = '{32'hc1d13fd7, 32'h40c025e3, 32'h40956ec8, 32'h41cc4829, 32'hc25f68f9, 32'hc2bc8921, 32'h4299a7e5, 32'h428889ba};
test_bias[1225:1225] = '{32'hc00725d7};
test_output[1225:1225] = '{32'h459b1370};
test_input[9808:9815] = '{32'h42525808, 32'h41745827, 32'h42316b45, 32'h419e07a5, 32'hc219dc60, 32'h41b53609, 32'hc2941733, 32'h42b6101e};
test_weights[9808:9815] = '{32'h41cda359, 32'h42330cc1, 32'hc1c8fa57, 32'hc1ddce71, 32'h42274f6a, 32'h42bb2a40, 32'hc2786878, 32'h42858e94};
test_bias[1226:1226] = '{32'hc2be7eeb};
test_output[1226:1226] = '{32'h463328fe};
test_input[9816:9823] = '{32'hc1694f3e, 32'hc2a56c73, 32'hc15f4918, 32'h41e08276, 32'h42c699d6, 32'hc29d92cf, 32'h4260291d, 32'h427a302d};
test_weights[9816:9823] = '{32'hc08da01a, 32'h41c8d461, 32'hc1093bd8, 32'hc2176c76, 32'h42c6220c, 32'h41cc16c4, 32'h42a30733, 32'hc2117835};
test_bias[1227:1227] = '{32'hc1f94862};
test_output[1227:1227] = '{32'h45def8f9};
test_input[9824:9831] = '{32'h428ba09e, 32'h420c510e, 32'hc1af80ca, 32'h427c7811, 32'hc2b5af67, 32'hc27b1242, 32'h3fc014fc, 32'hc26e9db9};
test_weights[9824:9831] = '{32'h41b6885b, 32'hc2713a2f, 32'h42afd241, 32'h428085d8, 32'h42c67e29, 32'h42c3f695, 32'h429fa531, 32'hc2bb332b};
test_bias[1228:1228] = '{32'h416c1197};
test_output[1228:1228] = '{32'hc5f5174b};
test_input[9832:9839] = '{32'hc247e8d7, 32'hc1c7d917, 32'h41655d22, 32'hc0ec6fb4, 32'h4283ad4c, 32'h42c76947, 32'h42bd72aa, 32'h42955c03};
test_weights[9832:9839] = '{32'h42a72926, 32'hc1eca0a5, 32'h41e4f1ed, 32'h42833945, 32'hc2a41901, 32'hc22f17a1, 32'hc2c6bad4, 32'h42c12db5};
test_bias[1229:1229] = '{32'h42bc9d84};
test_output[1229:1229] = '{32'hc6705f4b};
test_input[9840:9847] = '{32'h420fe4d6, 32'h424004da, 32'hc246bba2, 32'hc27c736b, 32'h41cfa30e, 32'h42a343b9, 32'h42096548, 32'hc18fb2fd};
test_weights[9840:9847] = '{32'h420a057c, 32'hc2175ebd, 32'hc21ee996, 32'h3f2ee114, 32'hc1ed82a4, 32'hc2bd9d44, 32'hc292cf0b, 32'h42baf72d};
test_bias[1230:1230] = '{32'h428ce26b};
test_output[1230:1230] = '{32'hc6305273};
test_input[9848:9855] = '{32'hc2c081f2, 32'hc2bb797b, 32'hc26754ae, 32'hc242b891, 32'hc1c8928e, 32'h429cbc3b, 32'hc1a05dc4, 32'hc244cdb2};
test_weights[9848:9855] = '{32'h3efab65a, 32'h3ff7febe, 32'hc2b5a682, 32'h41a42fa8, 32'h42019d0c, 32'hc0491d4f, 32'hc2c127be, 32'hc2a3296a};
test_bias[1231:1231] = '{32'hbfed1538};
test_output[1231:1231] = '{32'h460b489a};
test_input[9856:9863] = '{32'h3fbdfcb4, 32'h429a9972, 32'hc2a3b53b, 32'h405a6afe, 32'hc2bfe71f, 32'h42be9ac6, 32'h417eba24, 32'hc146df4a};
test_weights[9856:9863] = '{32'h421b8f66, 32'h424702e6, 32'hc295ed5a, 32'hc1d7e012, 32'hc0d9450f, 32'h41b86faa, 32'h42971524, 32'h41da8c88};
test_bias[1232:1232] = '{32'hc2724c0c};
test_output[1232:1232] = '{32'h46547ae6};
test_input[9864:9871] = '{32'h40fe27af, 32'hc02e3914, 32'h4182ebc4, 32'hc1ecccee, 32'h41be4eca, 32'h428fb02b, 32'hc1615f5d, 32'hc2bbca31};
test_weights[9864:9871] = '{32'hc2561786, 32'hc23b3a66, 32'h40041026, 32'hc1db8637, 32'hc2c057af, 32'h423faac2, 32'h4214ba5f, 32'hbf81dfbc};
test_bias[1233:1233] = '{32'hc26fdc1a};
test_output[1233:1233] = '{32'h4497d55b};
test_input[9872:9879] = '{32'hc2057282, 32'h4224479c, 32'h4109e277, 32'h42b49381, 32'hc15770d0, 32'h4202712e, 32'h4207f04d, 32'h422c8dfb};
test_weights[9872:9879] = '{32'hc126a4a4, 32'hc214ec49, 32'h427004df, 32'h42b7bac8, 32'h423be3fe, 32'hc1bf09e1, 32'hc296b37e, 32'h42873a7a};
test_bias[1234:1234] = '{32'h40ce3a7d};
test_output[1234:1234] = '{32'h45cda873};
test_input[9880:9887] = '{32'hc1e0141f, 32'hc196c986, 32'hc0aa8979, 32'hc1eccb8e, 32'hc29ca88c, 32'h408bde97, 32'hc2be312a, 32'hc0787246};
test_weights[9880:9887] = '{32'hc2c44fa8, 32'h420a2877, 32'h418ca7a9, 32'hc2ac94a4, 32'hc2265b68, 32'h41198e3f, 32'hc286af4e, 32'hc247df46};
test_bias[1235:1235] = '{32'hc1fafda1};
test_output[1235:1235] = '{32'h466163c7};
test_input[9888:9895] = '{32'h41fc68c0, 32'hc2098cc0, 32'hc2b0155e, 32'hc2270f8f, 32'h4239d097, 32'h42084ecb, 32'h4225a20a, 32'h4247e89c};
test_weights[9888:9895] = '{32'h42a2a823, 32'hc290eccf, 32'hc2180db5, 32'hc29bd7f0, 32'h42102483, 32'hc1600751, 32'hc0840f04, 32'h4292933a};
test_bias[1236:1236] = '{32'hc2832fa0};
test_output[1236:1236] = '{32'h467e6842};
test_input[9896:9903] = '{32'h41abd947, 32'hc28c6319, 32'h42b46116, 32'hc258fa73, 32'hc1f06703, 32'h40dc9bd6, 32'h42c6f836, 32'hc21721e0};
test_weights[9896:9903] = '{32'h4240affe, 32'hc0d7c12a, 32'hc289f849, 32'hc27948e4, 32'h4181dc2b, 32'h42bae5bd, 32'hbec92f34, 32'hc24a7bf4};
test_bias[1237:1237] = '{32'hc1b4d84d};
test_output[1237:1237] = '{32'h44289208};
test_input[9904:9911] = '{32'hc2314cff, 32'hc27ed978, 32'h42824695, 32'h41d5b190, 32'h4092ae74, 32'h4285f9a0, 32'h41892049, 32'hc238b784};
test_weights[9904:9911] = '{32'h41d19595, 32'hc2612ad8, 32'hc250c02c, 32'hc2b1e7b6, 32'h423a2fcb, 32'h401f2e26, 32'hc26489a1, 32'hc1c634fd};
test_bias[1238:1238] = '{32'hc23fa8c0};
test_output[1238:1238] = '{32'hc53255a9};
test_input[9912:9919] = '{32'h4110c8d3, 32'h42ac97de, 32'hc227bd72, 32'h4282c84b, 32'h41e8d9b2, 32'hc28dfe95, 32'hc186930a, 32'h42800040};
test_weights[9912:9919] = '{32'h4290c8c6, 32'h41b6567b, 32'hc19c8233, 32'hc29d1f85, 32'h4105cbc9, 32'hc2ae1cbb, 32'h429feac6, 32'hc29e75f5};
test_bias[1239:1239] = '{32'h411c533b};
test_output[1239:1239] = '{32'hc4d19935};
test_input[9920:9927] = '{32'h3fecd751, 32'h409c6268, 32'h42270179, 32'hc219f968, 32'hc2192d30, 32'hc17d30a6, 32'h42a133e6, 32'hc28382c8};
test_weights[9920:9927] = '{32'hc2735e9c, 32'h421599c1, 32'hc2c588ad, 32'h40c7e341, 32'h41907fef, 32'h42ae00e2, 32'h41dc1690, 32'h426e78d8};
test_bias[1240:1240] = '{32'hbf8cb0e6};
test_output[1240:1240] = '{32'hc5fc11d8};
test_input[9928:9935] = '{32'hc2b01f9b, 32'h42603b63, 32'h42139943, 32'hc2c1d096, 32'hc25f4f2f, 32'h4253f7f4, 32'h4208612c, 32'h42b8fb69};
test_weights[9928:9935] = '{32'h4294c03a, 32'hc2c0d676, 32'h426c2007, 32'hc286bf4e, 32'h4269f350, 32'h42a04982, 32'hc22a203d, 32'hc01116fd};
test_bias[1241:1241] = '{32'hc2a4caaf};
test_output[1241:1241] = '{32'hc57a7d98};
test_input[9936:9943] = '{32'h42919d2f, 32'hc22e5e25, 32'h419cbe60, 32'h412caed5, 32'hc29e0fb4, 32'hc29e4be4, 32'h42185cc3, 32'h41d30cf9};
test_weights[9936:9943] = '{32'hc29b6b57, 32'hc29ec69e, 32'h42c5e4fd, 32'hc28d9cfb, 32'h42ad60be, 32'hc1f0c852, 32'hc1a91b5f, 32'hc29381c7};
test_bias[1242:1242] = '{32'h41ff4b95};
test_output[1242:1242] = '{32'hc6004a1f};
test_input[9944:9951] = '{32'hc2b8f739, 32'h425fb150, 32'h42695ce5, 32'hc1c1e310, 32'h400cc436, 32'hc286c16d, 32'h41f77c26, 32'h42ad8697};
test_weights[9944:9951] = '{32'h41e575bd, 32'h42823435, 32'h428fbf3f, 32'h411ea933, 32'hc26b4ffc, 32'hc295dbc4, 32'hc1213367, 32'h42b6b579};
test_bias[1243:1243] = '{32'hc230e733};
test_output[1243:1243] = '{32'h46882cac};
test_input[9952:9959] = '{32'hc2c140d0, 32'h42a37689, 32'h41c97848, 32'h42c4e361, 32'hc2ba9543, 32'h41a379ca, 32'h426e4127, 32'h41a5e191};
test_weights[9952:9959] = '{32'h42a4ad1e, 32'h41784ea0, 32'hc26a5837, 32'h4291c831, 32'hc279d808, 32'hc2bbd92c, 32'h42b56941, 32'hc2b57766};
test_bias[1244:1244] = '{32'hc11671d4};
test_output[1244:1244] = '{32'h45c90333};
test_input[9960:9967] = '{32'h42ad48f8, 32'h427f7d56, 32'hc18ec23a, 32'h42380756, 32'hc1077be6, 32'h41093bc5, 32'h42aa472c, 32'h42b19c81};
test_weights[9960:9967] = '{32'hc2c68e70, 32'hbfa83aa3, 32'hc13d3f5d, 32'hc2a62c75, 32'h428cb02e, 32'h42519df4, 32'hc28afa53, 32'h42aaca0f};
test_bias[1245:1245] = '{32'hc20ba969};
test_output[1245:1245] = '{32'hc628ebdc};
test_input[9968:9975] = '{32'h42a4d9e8, 32'hc2bd6a42, 32'h42956cec, 32'hc2a97bc2, 32'hc23041b8, 32'hc2c7ac4a, 32'hc20f69fa, 32'h41d8c122};
test_weights[9968:9975] = '{32'hc10daf48, 32'hc280648b, 32'h425bb48e, 32'hc2bd5d44, 32'hc04c8813, 32'h4273e677, 32'hc1c13c20, 32'hc2a41a8a};
test_bias[1246:1246] = '{32'h42064f93};
test_output[1246:1246] = '{32'h461f7bc7};
test_input[9976:9983] = '{32'hc2bfb4c8, 32'h414f233c, 32'hc2bb759d, 32'hc2378988, 32'hc2af1a74, 32'h4224009b, 32'h4281fdd8, 32'h413b6b21};
test_weights[9976:9983] = '{32'hc1658c45, 32'hc2916515, 32'hc2719868, 32'hc1da4092, 32'hc2358f6b, 32'hc28b3231, 32'h420b029f, 32'h42551ab2};
test_bias[1247:1247] = '{32'h424c3d3b};
test_output[1247:1247] = '{32'h4632252c};
test_input[9984:9991] = '{32'h41278aaa, 32'h4222a25c, 32'h42059513, 32'h421bfdfe, 32'hc2980270, 32'h42c70628, 32'h42559875, 32'h42c41aae};
test_weights[9984:9991] = '{32'hc14f1add, 32'h42a0b25c, 32'hc2a085c5, 32'hc287fe3d, 32'hc23b458d, 32'hc2a2b305, 32'h3fd4831b, 32'hc2bc2954};
test_bias[1248:1248] = '{32'hc26c4c85};
test_output[1248:1248] = '{32'hc678f3a7};
test_input[9992:9999] = '{32'h42ab814f, 32'h41b3a778, 32'hc27fa91c, 32'h428ce30e, 32'h42be3e70, 32'h42c6aac6, 32'h410294cd, 32'hc039a971};
test_weights[9992:9999] = '{32'h418d2270, 32'h4216f4bc, 32'hc1acd12d, 32'h4174028c, 32'h42c3d055, 32'hc258eb71, 32'hc26a9e4f, 32'h4238b9d0};
test_bias[1249:1249] = '{32'h42aa24dd};
test_output[1249:1249] = '{32'h460057f0};
test_input[10000:10007] = '{32'hc2973747, 32'h421c00d6, 32'hc2b3dcea, 32'h3e5026ea, 32'hc1cf03aa, 32'h42a1521d, 32'hc16ee428, 32'hc2bebb76};
test_weights[10000:10007] = '{32'h3e96e37f, 32'hc285f26c, 32'hc127dd09, 32'h41db674c, 32'hc0c442f9, 32'h4259a9d2, 32'hc28b1b82, 32'h42b3826e};
test_bias[1250:1250] = '{32'hc1ac15e8};
test_output[1250:1250] = '{32'hc5923f25};
test_input[10008:10015] = '{32'h420ed48a, 32'h423b4fa3, 32'h42c13586, 32'h413c1842, 32'h41b9ac27, 32'h42673e14, 32'h414a2bf3, 32'hc231e12e};
test_weights[10008:10015] = '{32'hc2799fce, 32'hbe110f4f, 32'h4146e0ee, 32'h4295cb2b, 32'hc1dd5599, 32'h41ebba63, 32'h40e9bcad, 32'hc2c77942};
test_bias[1251:1251] = '{32'h41b46c96};
test_output[1251:1251] = '{32'h45aa8dd5};
test_input[10016:10023] = '{32'h42b1329f, 32'hc20e5f77, 32'h424d7db7, 32'h40dece27, 32'h42bbfebc, 32'hc1bb5ce6, 32'hc26dbbcd, 32'hc0f09e66};
test_weights[10016:10023] = '{32'h418fa149, 32'hc0962d98, 32'h42a163ab, 32'hc198eb73, 32'h4151303e, 32'hc2147ef5, 32'h4212e040, 32'h4192c860};
test_bias[1252:1252] = '{32'hc1a86ce2};
test_output[1252:1252] = '{32'h45acb992};
test_input[10024:10031] = '{32'h42875b4a, 32'hc211bc76, 32'h424cbdce, 32'h42606329, 32'hc2805f9b, 32'hc148b61a, 32'hc11e1c89, 32'hc1f5cdcb};
test_weights[10024:10031] = '{32'h42be5368, 32'h41a6e3bf, 32'hc2572266, 32'h42500515, 32'hc22df09d, 32'h40b4f034, 32'h421f953b, 32'hc285a244};
test_bias[1253:1253] = '{32'hc26c1c89};
test_output[1253:1253] = '{32'h461ed2e2};
test_input[10032:10039] = '{32'hc1b96bf8, 32'h4275189b, 32'hc28b8b75, 32'h429e90f4, 32'hc2b218d1, 32'hc2bdeec8, 32'h407eeba1, 32'h4164dc92};
test_weights[10032:10039] = '{32'h42563d60, 32'h413212ea, 32'hc20be5c4, 32'h421bf3e2, 32'hc23254a6, 32'h42415770, 32'hc2825692, 32'h4298d71f};
test_bias[1254:1254] = '{32'h41761821};
test_output[1254:1254] = '{32'h45a284c4};
test_input[10040:10047] = '{32'h4295f541, 32'hc28686c7, 32'h41af8951, 32'h428a4a2e, 32'hc29904d3, 32'hc29858e2, 32'hc2ba5faf, 32'h418b9964};
test_weights[10040:10047] = '{32'hc1507212, 32'h42019d13, 32'h413f02e4, 32'h41da2302, 32'h42c77686, 32'hc2aee19e, 32'hc19be84e, 32'h42913b0e};
test_bias[1255:1255] = '{32'h42c5e78c};
test_output[1255:1255] = '{32'h44966c07};
test_input[10048:10055] = '{32'hc276c674, 32'h41ca874e, 32'h423ffad8, 32'hc2a9de1c, 32'h41598af9, 32'h427d175d, 32'hc21aeaa6, 32'hc1022e49};
test_weights[10048:10055] = '{32'hc2a9d459, 32'h428abf97, 32'h42a6bda8, 32'hc2a1ba90, 32'h41eb8d99, 32'hc0ef624c, 32'h40be93db, 32'h4092f0b7};
test_bias[1256:1256] = '{32'hc2821fac};
test_output[1256:1256] = '{32'h468864d0};
test_input[10056:10063] = '{32'hc18cd1a3, 32'hc26c0fde, 32'h3f96c0ed, 32'h422fade4, 32'hc2a57b96, 32'hc194f413, 32'h421a9bd6, 32'h4205680a};
test_weights[10056:10063] = '{32'h424b08aa, 32'hbf47f786, 32'h41e8bece, 32'h42ac6eba, 32'hc1d70c73, 32'hc11b2736, 32'hc09ef14c, 32'hc1cc7262};
test_bias[1257:1257] = '{32'h422f5fc8};
test_output[1257:1257] = '{32'h4588ce0f};
test_input[10064:10071] = '{32'h414230c3, 32'h428063fe, 32'h3cd3a4d5, 32'h41b18c2f, 32'hc2aa7015, 32'h4243c625, 32'h409bad44, 32'h4240a296};
test_weights[10064:10071] = '{32'hc105ca31, 32'h429926da, 32'h4220f6be, 32'h41fe65d1, 32'h429ba372, 32'hc26a831d, 32'hc2736267, 32'h4293554c};
test_bias[1258:1258] = '{32'h42413e14};
test_output[1258:1258] = '{32'hc42a01d0};
test_input[10072:10079] = '{32'hc23c2529, 32'hc2516a7d, 32'h40b11e4c, 32'h42c3ce32, 32'hc2a95730, 32'h415e6f7c, 32'hc1616aa2, 32'h42bcc792};
test_weights[10072:10079] = '{32'h4288d0e1, 32'hc1efad83, 32'h42c27cc7, 32'hc187944a, 32'hc1695a83, 32'hc2903150, 32'h4281d2f2, 32'h41273053};
test_bias[1259:1259] = '{32'h4281eb0a};
test_output[1259:1259] = '{32'hc5160c51};
test_input[10080:10087] = '{32'hbf247061, 32'hc118fcf3, 32'h42b551d5, 32'h429de19d, 32'hc193e8ed, 32'hc0aaac42, 32'hc1b2b779, 32'h411769c0};
test_weights[10080:10087] = '{32'hc2c4f3bf, 32'h42c21bd0, 32'hc24f358c, 32'h42192b2f, 32'hc246894b, 32'h4246823a, 32'h4286f30d, 32'h42894690};
test_bias[1260:1260] = '{32'h42a5d606};
test_output[1260:1260] = '{32'hc52643f2};
test_input[10088:10095] = '{32'hc25a6f7f, 32'hc2599e73, 32'hc28d3684, 32'hc10706a7, 32'h4274ff92, 32'hc2840bab, 32'h42a33d0c, 32'hc2bc709a};
test_weights[10088:10095] = '{32'hc24614a4, 32'hc10c617d, 32'h41077fd0, 32'h424b6e97, 32'h424991fc, 32'hc27045a8, 32'h427871ca, 32'h42a75505};
test_bias[1261:1261] = '{32'hc2720b0f};
test_output[1261:1261] = '{32'h45c5e611};
test_input[10096:10103] = '{32'h427ae59d, 32'hc1f40aed, 32'h42310032, 32'h42bfeeb4, 32'h428dda19, 32'h41c42974, 32'hc224e8e3, 32'h428e1b85};
test_weights[10096:10103] = '{32'hc2a8ff54, 32'h4298a747, 32'hc2241ee2, 32'h42c1c147, 32'hc21f6bde, 32'hc2605cf3, 32'h40a45252, 32'hc2a2d25c};
test_bias[1262:1262] = '{32'h41453e7f};
test_output[1262:1262] = '{32'hc62174b3};
test_input[10104:10111] = '{32'h423bf5be, 32'h3f0e2fc1, 32'hc0271db4, 32'hc2b050e9, 32'hc2433722, 32'hc1a85b15, 32'hc19b8ebd, 32'hc1a51076};
test_weights[10104:10111] = '{32'h429bdf10, 32'hc1c6d7ee, 32'hc1c51876, 32'hc2714f87, 32'hc2bbf41d, 32'hc2af61b9, 32'h422701ca, 32'h42c0b4bd};
test_bias[1263:1263] = '{32'h411ac948};
test_output[1263:1263] = '{32'h464602c7};
test_input[10112:10119] = '{32'hc22386c0, 32'hc1a452d9, 32'h42042f5b, 32'hc26e8ca6, 32'hc290cdf3, 32'hc26ad001, 32'h42b013b5, 32'h41cad737};
test_weights[10112:10119] = '{32'h4226e65d, 32'h42b7e8d6, 32'hc29554d4, 32'h41b046a7, 32'h421b6093, 32'h4290eb19, 32'h414fcb91, 32'hc2267194};
test_bias[1264:1264] = '{32'hc1a56d17};
test_output[1264:1264] = '{32'hc66099b2};
test_input[10120:10127] = '{32'h424326d7, 32'h42729faf, 32'h42514c98, 32'hc2b59932, 32'hc0840179, 32'hc211289d, 32'hc217e182, 32'h42b47ff9};
test_weights[10120:10127] = '{32'h41e7fd54, 32'hc2b5cb19, 32'h4069bbfa, 32'h429a627b, 32'hc0d1d654, 32'hc28b004a, 32'hc271c10b, 32'h4202c148};
test_bias[1265:1265] = '{32'h4254c6fc};
test_output[1265:1265] = '{32'hc53fd207};
test_input[10128:10135] = '{32'hc2662273, 32'h42a44fe5, 32'hc29c2623, 32'hc22a4640, 32'h4252f89d, 32'h428c6454, 32'h4246501a, 32'hc045f085};
test_weights[10128:10135] = '{32'hc1aa23fd, 32'h42afc033, 32'hc25988a9, 32'h42a61693, 32'h42651cbb, 32'hc0fd99b3, 32'h4194a824, 32'h4203d2c1};
test_bias[1266:1266] = '{32'hc1ec0622};
test_output[1266:1266] = '{32'h4641e219};
test_input[10136:10143] = '{32'hc2b19bf6, 32'h42c6ebc2, 32'hc29de7d0, 32'h420eb536, 32'h42a26628, 32'h41ca39c1, 32'hc2a17351, 32'hc25fbf93};
test_weights[10136:10143] = '{32'hc2ab3d78, 32'h420ff43f, 32'h3eb10c23, 32'hc2bd5633, 32'hc1f84e82, 32'hc2663e5d, 32'h42a91106, 32'hc1f9740f};
test_bias[1267:1267] = '{32'h425c7d73};
test_output[1267:1267] = '{32'hc498bb5f};
test_input[10144:10151] = '{32'hc25394b0, 32'hc2952605, 32'h423577ab, 32'h4075f1c8, 32'hc166b1c4, 32'h40c70ce4, 32'hc2571571, 32'h4209034a};
test_weights[10144:10151] = '{32'hc2bd6321, 32'h4184bd66, 32'hc1825da8, 32'hc23b0329, 32'hc239f048, 32'h41f911e9, 32'h41efef2f, 32'hc1a3fab1};
test_bias[1268:1268] = '{32'hc0b07d99};
test_output[1268:1268] = '{32'h44ae835f};
test_input[10152:10159] = '{32'hc26f58ad, 32'h42a94154, 32'hc282c259, 32'h42c3b630, 32'hc17af8b1, 32'hc296be47, 32'h41f538d3, 32'hc284ab1e};
test_weights[10152:10159] = '{32'hc2a91823, 32'hbeba3b09, 32'hc2beb022, 32'hc22584ea, 32'h4239e28c, 32'h416e85ab, 32'hc2824c1c, 32'hc21bcc88};
test_bias[1269:1269] = '{32'hc19c26c1};
test_output[1269:1269] = '{32'h45b9396b};
test_input[10160:10167] = '{32'h424dbc68, 32'hc22e22a0, 32'h41ff0ba2, 32'hc29aa074, 32'h41c7009d, 32'hc23384ed, 32'hc2b22aac, 32'h41774054};
test_weights[10160:10167] = '{32'h42a639ad, 32'h42c57be4, 32'h3f9841bb, 32'hbfc2a47f, 32'hc11bda72, 32'hc2315428, 32'h420bc37d, 32'hc18449e2};
test_bias[1270:1270] = '{32'h4096b21c};
test_output[1270:1270] = '{32'hc4b98f3c};
test_input[10168:10175] = '{32'h42172165, 32'h3d6874e5, 32'hc2ba3472, 32'hc2b7c87a, 32'hc0b11899, 32'hc1824580, 32'h41d1646e, 32'hc2820e99};
test_weights[10168:10175] = '{32'hc0e92537, 32'h4296ba4f, 32'hc08082b3, 32'h421a9250, 32'h41482c26, 32'h42bd9ec0, 32'h42ba06de, 32'h42b6a113};
test_bias[1271:1271] = '{32'h42959684};
test_output[1271:1271] = '{32'hc604a799};
test_input[10176:10183] = '{32'h414ba3fd, 32'h425936b7, 32'h428cda02, 32'hc273aae3, 32'hc21a4927, 32'h422e04da, 32'hc2995fbc, 32'h42b81282};
test_weights[10176:10183] = '{32'hc29f7383, 32'hc299e893, 32'h426c5a92, 32'h42996f16, 32'h42ae68ac, 32'hc2077221, 32'hc2c52e1a, 32'hc2b2b6e2};
test_bias[1272:1272] = '{32'h418176b0};
test_output[1272:1272] = '{32'hc62ed6ad};
test_input[10184:10191] = '{32'hc281f067, 32'hc209f20f, 32'h41679c99, 32'hc298014c, 32'hc196e585, 32'hc1a4b40f, 32'hc2a6c235, 32'h42b4a6ee};
test_weights[10184:10191] = '{32'h4238dbcd, 32'h416a94d6, 32'hc293210d, 32'h42c0fb3b, 32'h429a39af, 32'h42252dc0, 32'hc29a5419, 32'hc2bfbda3};
test_bias[1273:1273] = '{32'hc2001ab9};
test_output[1273:1273] = '{32'hc680a9fa};
test_input[10192:10199] = '{32'h42681e36, 32'h42b58d17, 32'h42b8dc0d, 32'hc16440e5, 32'h41508dcb, 32'hc2b09fdb, 32'h40c24047, 32'hc180dd7b};
test_weights[10192:10199] = '{32'h4224e352, 32'hc2b386b8, 32'hc198c95b, 32'hc25f2d5c, 32'hc20559cf, 32'hc1b77812, 32'hc2b7a9cc, 32'hc0f2d179};
test_bias[1274:1274] = '{32'h420cebd8};
test_output[1274:1274] = '{32'hc5acf5c6};
test_input[10200:10207] = '{32'hc22f2da2, 32'h42c0f610, 32'hc282c157, 32'hc294ee5d, 32'hc1bca567, 32'hc297a62c, 32'hc1c5dac9, 32'h40a92816};
test_weights[10200:10207] = '{32'hc2963ad3, 32'hc2c78232, 32'h4104ef96, 32'h42c615e3, 32'h404be86a, 32'h42a29b6f, 32'hc2237e03, 32'hc2a88580};
test_bias[1275:1275] = '{32'hc1668d97};
test_output[1275:1275] = '{32'hc69bcc2d};
test_input[10208:10215] = '{32'h4298c2e1, 32'h410f61a8, 32'h41edd819, 32'hc1913db6, 32'hc2bfd0fa, 32'h42a5201d, 32'h4287de65, 32'h42afbc97};
test_weights[10208:10215] = '{32'h42b19179, 32'hc28e32fd, 32'h421994f5, 32'hc1b18d52, 32'h42ab1984, 32'h42abca43, 32'hc1a3351b, 32'h428b61ad};
test_bias[1276:1276] = '{32'hc1d006aa};
test_output[1276:1276] = '{32'h46305cb6};
test_input[10216:10223] = '{32'h42823d04, 32'hc22c67f3, 32'hc0e915c0, 32'hc2bca3ab, 32'hc2027631, 32'hc1d75db4, 32'hc2bc25e8, 32'h429ca7a5};
test_weights[10216:10223] = '{32'hc2b36427, 32'h42a1ff9f, 32'h42a62cd7, 32'h41c95607, 32'h42bbc00b, 32'h41dfa3ee, 32'hc186c0c8, 32'hc2595e35};
test_bias[1277:1277] = '{32'h42a498ed};
test_output[1277:1277] = '{32'hc69235ec};
test_input[10224:10231] = '{32'h41e618dc, 32'hc29f6c24, 32'hc2b1f6e8, 32'h4248c022, 32'h418fc36f, 32'hc2c35d4e, 32'hc2936b37, 32'hc2920145};
test_weights[10224:10231] = '{32'h42b4c81e, 32'hc29e4434, 32'hc28d99a7, 32'h4116ef24, 32'hc1e3f2a7, 32'h420a3b8f, 32'h42c101ba, 32'hc18dd495};
test_bias[1278:1278] = '{32'h428635d6};
test_output[1278:1278] = '{32'h45bccb54};
test_input[10232:10239] = '{32'h42a04cc7, 32'hc29d4902, 32'h41a6dca3, 32'h42adce04, 32'h41a84a7f, 32'h427c06b1, 32'hc107637b, 32'hc2a2e60b};
test_weights[10232:10239] = '{32'hc258ab2f, 32'h41cccefa, 32'hc2b7c357, 32'h42255556, 32'h4283af4f, 32'h4271da8b, 32'hc2944f14, 32'hc23eac5d};
test_bias[1279:1279] = '{32'hc2c1b5d1};
test_output[1279:1279] = '{32'h459a0460};
test_input[10240:10247] = '{32'h429cdcc8, 32'hc28c719e, 32'h417790b0, 32'hc2599e4a, 32'hc1bd2a9d, 32'h4297a099, 32'h4282771b, 32'hc2a155f3};
test_weights[10240:10247] = '{32'hc1e32930, 32'h429d759a, 32'h4277232f, 32'h422b63aa, 32'h4049e58d, 32'hc272dc66, 32'h42ba1187, 32'h427c89d9};
test_bias[1280:1280] = '{32'hc153d2d9};
test_output[1280:1280] = '{32'hc648b6ad};
test_input[10248:10255] = '{32'h4246813a, 32'hc25964f6, 32'hc27d38bb, 32'h4297c796, 32'h428c3db8, 32'hc2505ab9, 32'h42c63783, 32'h4134b7f8};
test_weights[10248:10255] = '{32'h42c102f6, 32'h41b3a41d, 32'h42c093f9, 32'h42a50945, 32'h426376d3, 32'h42b88573, 32'h41d049fa, 32'hc24a79b7};
test_bias[1281:1281] = '{32'h40c4733a};
test_output[1281:1281] = '{32'h459a2042};
test_input[10256:10263] = '{32'hc22bb487, 32'hc29f4680, 32'hc0be5143, 32'hc1c76095, 32'h42bc5365, 32'h41ac9122, 32'hc29c7f75, 32'h42a4695e};
test_weights[10256:10263] = '{32'h4207a011, 32'h4295ca78, 32'h428c0c84, 32'h41ba549d, 32'hc2be1a14, 32'h4116d87c, 32'hc224e24a, 32'h422c7b3c};
test_bias[1282:1282] = '{32'hc2a0d760};
test_output[1282:1282] = '{32'hc623a7f6};
test_input[10264:10271] = '{32'hc14df40c, 32'hc1eeef15, 32'hc2758bcb, 32'h42b5f455, 32'h422dc6d3, 32'hc29cad19, 32'hc1ca8455, 32'hc229dde3};
test_weights[10264:10271] = '{32'hc2b76ca1, 32'hc187d3e6, 32'hc11cf562, 32'hc2af9a5e, 32'hc1ba6269, 32'h42bf21ca, 32'hc0b1833a, 32'hc24d0897};
test_bias[1283:1283] = '{32'h4289f03a};
test_output[1283:1283] = '{32'hc6388a4a};
test_input[10272:10279] = '{32'h42b78972, 32'h428ebc7e, 32'h42068bba, 32'h428c100c, 32'h42a4ddbe, 32'hc24a18f5, 32'h423ff504, 32'hc14b818c};
test_weights[10272:10279] = '{32'hc285c286, 32'h42a70ff0, 32'hc250924d, 32'h41da6cae, 32'hc28f6913, 32'hbfce1234, 32'h42bfd1e8, 32'hc0003cee};
test_bias[1284:1284] = '{32'hc0ee7932};
test_output[1284:1284] = '{32'hc4995640};
test_input[10280:10287] = '{32'hc24961f2, 32'hc2820579, 32'hc2b6baf1, 32'h42092b22, 32'hc28e4e37, 32'hc2b077e9, 32'h41b44263, 32'h42ad967a};
test_weights[10280:10287] = '{32'h42143469, 32'h42340de4, 32'hc0dc9d94, 32'hc289c10d, 32'h428e8634, 32'h42aabe07, 32'h42b414ec, 32'hc20f7bb0};
test_bias[1285:1285] = '{32'h4294a0a5};
test_output[1285:1285] = '{32'hc69d5248};
test_input[10288:10295] = '{32'h41ac0303, 32'hc24eea10, 32'hc1f0c45c, 32'h4287e800, 32'h424c7e49, 32'h41a36031, 32'hc16b6b48, 32'hc21d7663};
test_weights[10288:10295] = '{32'h41609ef2, 32'h4294e0c5, 32'h41af8f55, 32'hc28d923c, 32'h42811360, 32'h40f3fef2, 32'hc2475d79, 32'h4264e361};
test_bias[1286:1286] = '{32'h4023309b};
test_output[1286:1286] = '{32'hc5dd473b};
test_input[10296:10303] = '{32'hc28e2638, 32'hc2c2d0ac, 32'h420429e3, 32'hc00d2683, 32'h41b4a72f, 32'h42830821, 32'h417925d8, 32'h42893c61};
test_weights[10296:10303] = '{32'hc2098a6a, 32'h4229e6e4, 32'hc21ce4b7, 32'h404b309c, 32'hc1056003, 32'hc206c394, 32'hc2b57b1d, 32'hc1ecc980};
test_bias[1287:1287] = '{32'h424fefaf};
test_output[1287:1287] = '{32'hc609400e};
test_input[10304:10311] = '{32'h41c568c7, 32'hc236162f, 32'h40aed4fd, 32'hc2845ec5, 32'hc02fed28, 32'h42a196f3, 32'h41ae8540, 32'hc2845c76};
test_weights[10304:10311] = '{32'hc2345498, 32'h421215d1, 32'hc05a8069, 32'h42b9238b, 32'h41cd5301, 32'hc1d0a1fd, 32'hc290a178, 32'h426933d6};
test_bias[1288:1288] = '{32'h42ba022f};
test_output[1288:1288] = '{32'hc68071c3};
test_input[10312:10319] = '{32'hc25b48b5, 32'hc12a02df, 32'h42ab0fe4, 32'hc296ca0d, 32'h42a28925, 32'h424f6f20, 32'h41380733, 32'h42a0c3c1};
test_weights[10312:10319] = '{32'hc2adacbb, 32'hc1c4e64c, 32'hc1e51307, 32'hc2b7bd3b, 32'hc08564f2, 32'hc29ef7fa, 32'h4265ff57, 32'hc2ab3d14};
test_bias[1289:1289] = '{32'hc296612f};
test_output[1289:1289] = '{32'hc49d2e42};
test_input[10320:10327] = '{32'h41ec3772, 32'hc28c5057, 32'h426ad81c, 32'hc2c6cef1, 32'h42195e92, 32'hc2c5646e, 32'h42c74428, 32'h42b040ed};
test_weights[10320:10327] = '{32'hc23e509b, 32'h4113a14b, 32'hc2b2a102, 32'h41d28086, 32'h424e31ea, 32'hc243ce4c, 32'h41a29c1f, 32'hc2339d01};
test_bias[1290:1290] = '{32'hc235f134};
test_output[1290:1290] = '{32'hc59ec9c0};
test_input[10328:10335] = '{32'hc29c356d, 32'hc1e65222, 32'hc21ec9d2, 32'hc0293596, 32'hc26bd6bb, 32'h4088d11d, 32'h423ac594, 32'hc1248043};
test_weights[10328:10335] = '{32'hc264463c, 32'hc2b29690, 32'h4293f42e, 32'h413226f8, 32'hc24bb6f4, 32'hc252b674, 32'h42bdb9a4, 32'h428b0798};
test_bias[1291:1291] = '{32'hc1bc38f4};
test_output[1291:1291] = '{32'h46248ab6};
test_input[10336:10343] = '{32'h417c1b0c, 32'h42874ed3, 32'h42b3a76b, 32'hc2a43ca2, 32'hc2463076, 32'hc29c6494, 32'hc28214d5, 32'h42452598};
test_weights[10336:10343] = '{32'h40521640, 32'h417dc690, 32'h420da3b7, 32'h42a61131, 32'hc29f8765, 32'h42a42f73, 32'h42b24592, 32'hc1da3f7a};
test_bias[1292:1292] = '{32'h42c51b9f};
test_output[1292:1292] = '{32'hc63bdf1d};
test_input[10344:10351] = '{32'h427c1675, 32'hc1f21a6a, 32'h42c45652, 32'h42b7b1f6, 32'hc2b103cc, 32'hc2012341, 32'h42944274, 32'h42118724};
test_weights[10344:10351] = '{32'hc2159872, 32'h42883182, 32'hc29e9b70, 32'h41d52652, 32'h41a53f2f, 32'hc297f720, 32'h42a9df54, 32'h428f7d8d};
test_bias[1293:1293] = '{32'h41a5e381};
test_output[1293:1293] = '{32'hc34b952f};
test_input[10352:10359] = '{32'hc1ac848e, 32'hc27e3263, 32'h40d9fa01, 32'h42be56cf, 32'hc2b87ad3, 32'h412fea28, 32'h41988ae7, 32'h427e16a8};
test_weights[10352:10359] = '{32'hc2bcb793, 32'hc1880081, 32'hc2c690ac, 32'hc2bd33e8, 32'hc2add371, 32'h40763ea8, 32'h42060252, 32'h421ba89b};
test_bias[1294:1294] = '{32'h411cc4c2};
test_output[1294:1294] = '{32'h45903b44};
test_input[10360:10367] = '{32'h40bc5c66, 32'h428ec4ca, 32'h41afba04, 32'hc1d7cd92, 32'hc2b72854, 32'hc14b8d07, 32'h429929fc, 32'hc228983b};
test_weights[10360:10367] = '{32'h4295665c, 32'h425734c2, 32'hc26b82c9, 32'hc2426295, 32'hc0abd6d1, 32'h42aab298, 32'h419da7b9, 32'h41396568};
test_bias[1295:1295] = '{32'h42a294e2};
test_output[1295:1295] = '{32'h45962fbc};
test_input[10368:10375] = '{32'h41fd71c6, 32'h4297a0c6, 32'hc2c50ce5, 32'h419b69a7, 32'h41fc42d7, 32'hc2ba2cf3, 32'hc2a69295, 32'h400450ce};
test_weights[10368:10375] = '{32'hc25871c7, 32'h423da2d5, 32'hc2af30d2, 32'h41a9897e, 32'hc1a7500c, 32'hc2b74ced, 32'hc1e1aa0e, 32'hc2604035};
test_bias[1296:1296] = '{32'h42325f9e};
test_output[1296:1296] = '{32'h46a4a038};
test_input[10376:10383] = '{32'hc1e88f6e, 32'hc188bfae, 32'hc1483be2, 32'h41e8d04d, 32'hc2948a9e, 32'hc244cbaf, 32'h425b6c39, 32'hc1f2b53b};
test_weights[10376:10383] = '{32'h41e31aa9, 32'h425733b0, 32'h4093a29e, 32'h404653f9, 32'h41c79fa6, 32'h42c09bb9, 32'h42a0ffa6, 32'h40b4e017};
test_bias[1297:1297] = '{32'hc2a2a2eb};
test_output[1297:1297] = '{32'hc58165d6};
test_input[10384:10391] = '{32'h40f58299, 32'h42830afb, 32'hc1a4d6eb, 32'hc2b073a5, 32'h426f75b7, 32'hc23badcf, 32'hc29c0624, 32'h42b6a650};
test_weights[10384:10391] = '{32'hc2aaea4b, 32'h42990687, 32'hc29d3224, 32'h4270c1aa, 32'h3f823dc4, 32'h42233a05, 32'h3f8c4fb3, 32'hc2986621};
test_bias[1298:1298] = '{32'h425baec4};
test_output[1298:1298] = '{32'hc5ff8302};
test_input[10392:10399] = '{32'h42a0b8a1, 32'h4156934d, 32'h424a8b47, 32'h41cafb4d, 32'h42ad4ec1, 32'hc25017f5, 32'hc07872f2, 32'hc239eee7};
test_weights[10392:10399] = '{32'hc17733a6, 32'h426167d7, 32'hc2bc8d64, 32'h42575fc8, 32'h42b978fe, 32'h42177cc2, 32'hc2545eda, 32'hc29e265f};
test_bias[1299:1299] = '{32'hc2688887};
test_output[1299:1299] = '{32'h45bb5f3f};
test_input[10400:10407] = '{32'h42246aef, 32'h42224548, 32'hc273a2d1, 32'h42b4b467, 32'h423a85f0, 32'h42915da7, 32'h42bf0232, 32'hc2b7f1e5};
test_weights[10400:10407] = '{32'hc1bb6bf2, 32'h42713eb3, 32'h4246735f, 32'h42789735, 32'hc1848714, 32'h40ccd1c1, 32'h42c2e7cb, 32'hc172c416};
test_bias[1300:1300] = '{32'hc1b78666};
test_output[1300:1300] = '{32'h4661c5d8};
test_input[10408:10415] = '{32'h4104b862, 32'hc248242d, 32'hc28c7792, 32'h428d6917, 32'h40145e41, 32'h410771f5, 32'h41ac23e1, 32'hc20660d0};
test_weights[10408:10415] = '{32'hc1469a68, 32'hc292828b, 32'hc1468519, 32'h42b1a5a0, 32'hc262bbb4, 32'h40b7e7cb, 32'h42c57358, 32'hc2a23cd6};
test_bias[1301:1301] = '{32'hc0aba3a5};
test_output[1301:1301] = '{32'h4671cdbe};
test_input[10416:10423] = '{32'hc21e0c42, 32'hc28e9274, 32'h422a3f0c, 32'h420bb7d7, 32'hc0758344, 32'h42651083, 32'hc138c952, 32'h4296f1cf};
test_weights[10416:10423] = '{32'hc27d7fdb, 32'h41a41239, 32'hc2b07f30, 32'h423f8f80, 32'hc22c1321, 32'hc2a4f114, 32'hc241f086, 32'hc1bbe26f};
test_bias[1302:1302] = '{32'hc2824c58};
test_output[1302:1302] = '{32'hc5d6e4d3};
test_input[10424:10431] = '{32'hc2106581, 32'hc2889b88, 32'h42be04c0, 32'hc2a10bfb, 32'hc1ed33fa, 32'h42357aa7, 32'h4139d7cc, 32'h42b352bc};
test_weights[10424:10431] = '{32'h4040c7bc, 32'hc2123a44, 32'h424f46b0, 32'hc22c5826, 32'h42072799, 32'hc2038fb3, 32'h413b02c1, 32'h418285a5};
test_bias[1303:1303] = '{32'hc1e9054e};
test_output[1303:1303] = '{32'h461a017e};
test_input[10432:10439] = '{32'h426f4a1c, 32'hbfd75ea3, 32'hc15c4c6c, 32'h425df9f6, 32'hc005d615, 32'hc004821c, 32'h428f930e, 32'hc1f97642};
test_weights[10432:10439] = '{32'hc22f1571, 32'h42b8620b, 32'h42aa9e37, 32'hc1d1bb3c, 32'hc284e6e0, 32'h42c2a954, 32'h41a8c763, 32'hc2c5b33e};
test_bias[1304:1304] = '{32'h42b07206};
test_output[1304:1304] = '{32'hc4431c68};
test_input[10440:10447] = '{32'h429310fc, 32'h41c16f15, 32'h42739051, 32'hc21af033, 32'hc2972b5f, 32'hc00394e2, 32'hc0bee2a8, 32'hc2051613};
test_weights[10440:10447] = '{32'hc233200b, 32'hc14362e5, 32'hc2abfaaf, 32'h42bdccd1, 32'hc2abbad5, 32'h42c1f610, 32'h428a797b, 32'h42a93532};
test_bias[1305:1305] = '{32'hc2a9a5bb};
test_output[1305:1305] = '{32'hc614c887};
test_input[10448:10455] = '{32'hc2b813ca, 32'h41bda513, 32'hc19fcc30, 32'h42012b03, 32'h421c5f42, 32'h429aac9d, 32'hc16eb44d, 32'hc20fe7bb};
test_weights[10448:10455] = '{32'hc234b621, 32'hc29e26eb, 32'hc26a62a6, 32'h42affadf, 32'h42538b63, 32'hc28c46ac, 32'h3fc96de6, 32'h41d58df6};
test_bias[1306:1306] = '{32'hc0933a71};
test_output[1306:1306] = '{32'h44f3c49c};
test_input[10456:10463] = '{32'h424c23b1, 32'hc20dae10, 32'hc262b015, 32'h42c2c509, 32'hc26154bd, 32'h429be22d, 32'hc22f90c6, 32'h41b260b6};
test_weights[10456:10463] = '{32'h40ada9d7, 32'h4243cda6, 32'h421c9fba, 32'hc2a994a6, 32'h42918a47, 32'h42a5c833, 32'h4280aabd, 32'h426f1cb0};
test_bias[1307:1307] = '{32'h41cfa22f};
test_output[1307:1307] = '{32'hc62c72e7};
test_input[10464:10471] = '{32'hc1a5d723, 32'hc290f79e, 32'h42b1a7e6, 32'hc275f858, 32'h42aa9530, 32'hc1fb391b, 32'hc282537c, 32'h426c6e39};
test_weights[10464:10471] = '{32'hc22ce322, 32'h4280b4b1, 32'h42af607f, 32'h42544439, 32'hc20bd0cd, 32'h41471a17, 32'h418ddd6c, 32'hc297b289};
test_bias[1308:1308] = '{32'hc2957595};
test_output[1308:1308] = '{32'hc6022070};
test_input[10472:10479] = '{32'hc27b3d48, 32'hc206adcb, 32'hc2ad6d38, 32'h42b3bdf0, 32'h429dd612, 32'h4288bd46, 32'h419e6e00, 32'h4298cac2};
test_weights[10472:10479] = '{32'hc29b7bc2, 32'hc26dc56e, 32'hc16e435f, 32'h423bf840, 32'h3fc98596, 32'hc28def02, 32'hc1f7d4bd, 32'hc2af0b23};
test_bias[1309:1309] = '{32'hc2c2b1e7};
test_output[1309:1309] = '{32'h438902e2};
test_input[10480:10487] = '{32'h425c9709, 32'h42b8362e, 32'hc2c4e288, 32'hc14978e9, 32'h4277afb0, 32'hc1fe18be, 32'h426afcf3, 32'hc29cf4d8};
test_weights[10480:10487] = '{32'h4298707d, 32'hc1eb3347, 32'hc29fcaed, 32'hc1d61c7b, 32'h416e36bb, 32'h422fad76, 32'h429ffb6d, 32'hc1b88db0};
test_bias[1310:1310] = '{32'h426b8a61};
test_output[1310:1310] = '{32'h4676c46a};
test_input[10488:10495] = '{32'hc23ae126, 32'hc1ddaf47, 32'h42c50931, 32'h41048b70, 32'h427e6da3, 32'h41d449b5, 32'h42c60622, 32'hc2af3dbb};
test_weights[10488:10495] = '{32'hc14d48d7, 32'h41c07411, 32'h425253c6, 32'hc2887fa4, 32'hc1d9514f, 32'h428c1bfc, 32'h41839c1c, 32'hc1bae4fe};
test_bias[1311:1311] = '{32'hc1ae6f4e};
test_output[1311:1311] = '{32'h46023346};
test_input[10496:10503] = '{32'hc2a4fbc8, 32'hc29f6438, 32'hc286ad03, 32'hc2bf35c3, 32'hc25f835f, 32'hbf100c82, 32'h4217e546, 32'h426c1f76};
test_weights[10496:10503] = '{32'h4216b3e3, 32'hc1862175, 32'h4282264b, 32'hc122199c, 32'hc2a0ebcc, 32'h427dbff9, 32'h42ad4525, 32'hc25ddf86};
test_bias[1312:1312] = '{32'hbffb09fa};
test_output[1312:1312] = '{32'hc431d014};
test_input[10504:10511] = '{32'hc06a219f, 32'hc0b91413, 32'h40ccf480, 32'h429db095, 32'h42320597, 32'h4289304f, 32'h409373af, 32'h4218fbcb};
test_weights[10504:10511] = '{32'hc23a0cdd, 32'h41289310, 32'hc21249af, 32'hc16506f1, 32'h42bc0d7e, 32'hc197828d, 32'h42509e7e, 32'h4198083c};
test_bias[1313:1313] = '{32'hc28d37e4};
test_output[1313:1313] = '{32'h451e083f};
test_input[10512:10519] = '{32'h42855f92, 32'h42bd6d5c, 32'hc25e59b6, 32'h42515cbb, 32'hc2423a0f, 32'h4193a40d, 32'h410cae2f, 32'h40d56fba};
test_weights[10512:10519] = '{32'h422de33c, 32'hc29dd62b, 32'h42c0e570, 32'hc2662308, 32'hc2164510, 32'h42c57f72, 32'h41bfb27c, 32'hc28bbb86};
test_bias[1314:1314] = '{32'h41b4aaef};
test_output[1314:1314] = '{32'hc614f9f4};
test_input[10520:10527] = '{32'h4271b55e, 32'hc22c0bea, 32'hc2670f4f, 32'hc25e63b9, 32'hc1e775ac, 32'hc15dc41d, 32'h4228f4bb, 32'hc27550f2};
test_weights[10520:10527] = '{32'h42b5107a, 32'h42b81ff3, 32'hc1d0e187, 32'h42488b50, 32'hc2c6e38d, 32'h425b7360, 32'h42889ce8, 32'hc2a27bda};
test_bias[1315:1315] = '{32'h42a8644e};
test_output[1315:1315] = '{32'h4620f12e};
test_input[10528:10535] = '{32'h4228d973, 32'hc2c3961e, 32'h42ac45ed, 32'h42a3cf00, 32'hc20b1f90, 32'h429b04ef, 32'h42b26515, 32'h41b6a109};
test_weights[10528:10535] = '{32'h40c89537, 32'h42ad1a62, 32'h42a412fd, 32'h42ad23e3, 32'hc1b7d4a3, 32'hc1381fd7, 32'hc2af75f1, 32'hc2620ac8};
test_bias[1316:1316] = '{32'hc255ae51};
test_output[1316:1316] = '{32'hc54e83d5};
test_input[10536:10543] = '{32'h41f64531, 32'h4289cbc5, 32'h4223bfc0, 32'hc2ac8651, 32'h42452cfe, 32'h4216af15, 32'hc0d09502, 32'h413f1212};
test_weights[10536:10543] = '{32'hc1b80ff8, 32'hc2a65aac, 32'h40fb6bef, 32'h41d208dd, 32'hc2bf20d8, 32'hc2787ac3, 32'h4260caaf, 32'hc2869351};
test_bias[1317:1317] = '{32'h42b6654b};
test_output[1317:1317] = '{32'hc680ff40};
test_input[10544:10551] = '{32'h429d9477, 32'h42bf570a, 32'hc1f61579, 32'hc209236e, 32'hc0fc6db6, 32'hc22dccba, 32'h410f15bd, 32'hc1855931};
test_weights[10544:10551] = '{32'h42c12cc0, 32'h428dfd3f, 32'h422ca7ee, 32'hc268a52b, 32'h42a525f9, 32'h4251b2b7, 32'hc2b0f230, 32'h42b428b8};
test_bias[1318:1318] = '{32'h41bb1c87};
test_output[1318:1318] = '{32'h461a37c5};
test_input[10552:10559] = '{32'h42489221, 32'h428480a5, 32'hc21aba2e, 32'h4222481e, 32'h41ed572d, 32'h42039c7e, 32'hc2a0f13d, 32'h42615009};
test_weights[10552:10559] = '{32'h3f8210da, 32'hc1d85919, 32'hc29da54c, 32'h428cecb4, 32'h41a12faf, 32'h42bc08d8, 32'hc2b7b9d7, 32'h42c0b67f};
test_bias[1319:1319] = '{32'hc140509d};
test_output[1319:1319] = '{32'h46a17419};
test_input[10560:10567] = '{32'h423e9c80, 32'h4278fb49, 32'hc2ab58b3, 32'h41068133, 32'hc195d5b9, 32'h42892d60, 32'h42920eea, 32'hc09f0c0c};
test_weights[10560:10567] = '{32'h40489b18, 32'h42c180ef, 32'h429d3ef8, 32'h429c6855, 32'h4045e273, 32'h417d7f52, 32'hc1d8321b, 32'h40d9a35b};
test_bias[1320:1320] = '{32'h419c0911};
test_output[1320:1320] = '{32'hc4587556};
test_input[10568:10575] = '{32'h429db406, 32'h4121d504, 32'h42bee35c, 32'hc20956a5, 32'h42c36cb8, 32'hc2939b45, 32'hc2b31a51, 32'hc1b77d62};
test_weights[10568:10575] = '{32'h42bfbe5b, 32'hc267d496, 32'hc1f63d99, 32'h4162604a, 32'h40e776f5, 32'hc29e1b3d, 32'hc2c79958, 32'hc1c0d11b};
test_bias[1321:1321] = '{32'hc2c670e8};
test_output[1321:1321] = '{32'h469833a0};
test_input[10576:10583] = '{32'h40f61feb, 32'hc2a1421b, 32'hc2359a99, 32'h41a655e3, 32'hc2026d9f, 32'h4203f853, 32'hc0fc8c9f, 32'h42497453};
test_weights[10576:10583] = '{32'hc0e2865c, 32'hc2992be6, 32'h42051e0c, 32'hc29b5412, 32'h4290569d, 32'hc2add2d0, 32'h4159c944, 32'hc25f7c2f};
test_bias[1322:1322] = '{32'h423b5472};
test_output[1322:1322] = '{32'hc59f61ef};
test_input[10584:10591] = '{32'h425e5eea, 32'hc2a50440, 32'hc05d3bc1, 32'h4299b69d, 32'hc1b4ebe4, 32'hc2c2ce9a, 32'h428a2c6b, 32'h420197e7};
test_weights[10584:10591] = '{32'hc266f2d1, 32'hc236dd70, 32'h42c71365, 32'hc29a323d, 32'hc1ba9046, 32'hc2327080, 32'h429f56ea, 32'h420c97e0};
test_bias[1323:1323] = '{32'h41bdb21e};
test_output[1323:1323] = '{32'h45b63e16};
test_input[10592:10599] = '{32'h42bca583, 32'hc2bfbcc1, 32'h42518621, 32'h42a2cad5, 32'h40b528c7, 32'hc16db0db, 32'h42b5b909, 32'hc2a518d2};
test_weights[10592:10599] = '{32'h4259528c, 32'h4230c23c, 32'h42c0b216, 32'hc28fd3d4, 32'h42298d1b, 32'h422751d6, 32'hc1b6189e, 32'h419833fc};
test_bias[1324:1324] = '{32'hc26bff85};
test_output[1324:1324] = '{32'hc579d9f0};
test_input[10600:10607] = '{32'h42578d29, 32'h424900fe, 32'h40b1d616, 32'h42c3932a, 32'hc2bc32d4, 32'h4204c52d, 32'hc21e90f0, 32'hc2639656};
test_weights[10600:10607] = '{32'h42c66c50, 32'hc2a635e4, 32'h423b9dcb, 32'h424a1ad4, 32'hc2043b94, 32'h427ec06f, 32'h42b9ad6d, 32'hc2bebfd5};
test_bias[1325:1325] = '{32'h42a7e80b};
test_output[1325:1325] = '{32'h4651ca55};
test_input[10608:10615] = '{32'h42440ce4, 32'h429fa9d4, 32'h428291bc, 32'hc2b3c689, 32'hc2170835, 32'h42528fa3, 32'h426c7d6e, 32'h41ebfb58};
test_weights[10608:10615] = '{32'h41f498bc, 32'hc2b5ac95, 32'h417299ad, 32'hc124d689, 32'h4297e747, 32'hc2423fda, 32'hc2769d78, 32'h408ef537};
test_bias[1326:1326] = '{32'hc16e759e};
test_output[1326:1326] = '{32'hc647d64a};
test_input[10616:10623] = '{32'h404e8f5e, 32'hc0ae964e, 32'hc24c14e0, 32'hc2c371a1, 32'h42076576, 32'h41e2a0a2, 32'h42c29d08, 32'h4285196d};
test_weights[10616:10623] = '{32'h42280cfb, 32'h42479e17, 32'hc1c445c0, 32'h42142997, 32'hc23fd3cf, 32'hc2c4f1a7, 32'h40a41f24, 32'hc16bd3b1};
test_bias[1327:1327] = '{32'h427ff44d};
test_output[1327:1327] = '{32'hc5e53a6c};
test_input[10624:10631] = '{32'h418fcb3a, 32'h42a3d8a6, 32'hc28b29a2, 32'h42a56fc8, 32'hc05a19e1, 32'hc26df644, 32'h42a28f1c, 32'h4257f173};
test_weights[10624:10631] = '{32'hc2807cc1, 32'hc1ec4918, 32'h42491f94, 32'h41b94fbf, 32'h420b21e5, 32'h4178adfa, 32'hc283da14, 32'h42348d57};
test_bias[1328:1328] = '{32'hc273acf7};
test_output[1328:1328] = '{32'hc60f7a71};
test_input[10632:10639] = '{32'hc2b6c96f, 32'hc1ce7f86, 32'h4212953e, 32'hc1a6482c, 32'h427ae35f, 32'h3f486569, 32'hc23a2d1b, 32'h42808b4d};
test_weights[10632:10639] = '{32'hc1ad56b3, 32'h40c5c1ca, 32'hc28519c3, 32'h42b699e0, 32'hc282879f, 32'hc29ec050, 32'hc1ce6c4e, 32'hc2ae0a13};
test_bias[1329:1329] = '{32'hc13d7c83};
test_output[1329:1329] = '{32'hc62d0cfa};
test_input[10640:10647] = '{32'h41dfe00a, 32'hc2a1ee0f, 32'hc20973cd, 32'h42c155d3, 32'hc216c885, 32'hc295481a, 32'hc2b26535, 32'h428b7274};
test_weights[10640:10647] = '{32'h3fd2404f, 32'h4247b637, 32'hc2522f18, 32'hc0a0258e, 32'hc2289597, 32'h412a55df, 32'hc23e5e5e, 32'h42ab7b5e};
test_bias[1330:1330] = '{32'hc23acff5};
test_output[1330:1330] = '{32'h4601a05d};
test_input[10648:10655] = '{32'hc245d4cb, 32'hc16e3372, 32'hc2912e11, 32'h421baa9a, 32'h4292d51e, 32'hc1ce05b8, 32'h4256437d, 32'hc2446173};
test_weights[10648:10655] = '{32'hc1e453ff, 32'h42aa491e, 32'h4181cf21, 32'hc2303bfe, 32'h425ebff0, 32'hc1a2aa49, 32'h4270c858, 32'h42a46029};
test_bias[1331:1331] = '{32'hc22da1e7};
test_output[1331:1331] = '{32'h447c62b0};
test_input[10656:10663] = '{32'hc28dfe26, 32'h428ef058, 32'h42b923c5, 32'h41fe25d5, 32'h42c35a04, 32'hc2af10c1, 32'h41a51b52, 32'hc29d2206};
test_weights[10656:10663] = '{32'hc1c00bd0, 32'hc259ac0a, 32'hc0feccf2, 32'h41cd2d4f, 32'h417e3ea0, 32'hc24fe301, 32'h416320ec, 32'h41a09010};
test_bias[1332:1332] = '{32'h411564e5};
test_output[1332:1332] = '{32'h4529f8dd};
test_input[10664:10671] = '{32'hc251da78, 32'hc195dcf6, 32'hc2034ad3, 32'hc2bbccae, 32'hc018a279, 32'h4224c875, 32'h421dc6d3, 32'hc1668ed7};
test_weights[10664:10671] = '{32'hc28916fa, 32'hc29528af, 32'hc0a34bd8, 32'h4291a0f0, 32'h420b31ab, 32'h402ae496, 32'h421bb11d, 32'h412f6744};
test_bias[1333:1333] = '{32'hc1a95fea};
test_output[1333:1333] = '{32'hc392b5a0};
test_input[10672:10679] = '{32'hc27afafa, 32'h4280da5e, 32'h420f1be0, 32'h42a4ab74, 32'hc29b783e, 32'hc29b8460, 32'hc2c6f4ac, 32'hc12ac224};
test_weights[10672:10679] = '{32'hc1dbc21e, 32'h42b32f2b, 32'hbfc97c5b, 32'h42c37e7d, 32'hc2c7514c, 32'h41c530b4, 32'h42bfc69e, 32'hc1e93663};
test_bias[1334:1334] = '{32'hc214b0e3};
test_output[1334:1334] = '{32'h463c5398};
test_input[10680:10687] = '{32'hc29a78d7, 32'h3ea5ee63, 32'h4238e62e, 32'h423cbce3, 32'h42422058, 32'h421c2b78, 32'hc2ba88c8, 32'hc29e17b4};
test_weights[10680:10687] = '{32'h422e45d8, 32'h42850c81, 32'hc184fe66, 32'hc0391512, 32'hc205da0f, 32'hc232f5ec, 32'hc1d7d0fe, 32'hc24d0056};
test_bias[1335:1335] = '{32'h4290f973};
test_output[1335:1335] = '{32'hc474dc9a};
test_input[10688:10695] = '{32'h41fdff5f, 32'h41314db7, 32'h414c614d, 32'hc2b05e27, 32'hc22422d8, 32'hc128050c, 32'hc292c6e2, 32'hc1ee3208};
test_weights[10688:10695] = '{32'h426d8c83, 32'hc2a77be2, 32'hc2034919, 32'h42993886, 32'h42413f2b, 32'h424c2116, 32'hc2c44269, 32'hc2089f9f};
test_bias[1336:1336] = '{32'hc29781c1};
test_output[1336:1336] = '{32'hc414422b};
test_input[10696:10703] = '{32'h3fdeb94c, 32'hc29ffda7, 32'hc291f7a2, 32'h42c301a1, 32'h4218b41a, 32'hc22dd8de, 32'hc158a8c0, 32'h41a16060};
test_weights[10696:10703] = '{32'hc11999d6, 32'h41cb4b9d, 32'hc23cea65, 32'hc22490d1, 32'hc2502f41, 32'h410e1795, 32'hc1204d5e, 32'hc1802172};
test_bias[1337:1337] = '{32'hc2709127};
test_output[1337:1337] = '{32'hc5a393af};
test_input[10704:10711] = '{32'hc1912058, 32'hc0dd4b03, 32'hc2af267f, 32'h42a6fdb5, 32'h429deb4c, 32'hc2b90165, 32'hc2be893f, 32'h41b6145e};
test_weights[10704:10711] = '{32'h41e049e4, 32'hc287e477, 32'h40c75d44, 32'h421ead97, 32'hc18dbe65, 32'h42a9f4ae, 32'hc2825f01, 32'hc2807d86};
test_bias[1338:1338] = '{32'hc1d44c69};
test_output[1338:1338] = '{32'hc4e24e19};
test_input[10712:10719] = '{32'hc28e96eb, 32'hc21f980c, 32'h4130df68, 32'h42905c7f, 32'h427d4f80, 32'hc26af526, 32'hc222f871, 32'hc271ac35};
test_weights[10712:10719] = '{32'h42b24fa4, 32'h4283fb7f, 32'h4236c8c4, 32'hc189b669, 32'hc2c65917, 32'hc2c55a9d, 32'hc2970417, 32'hc18cb710};
test_bias[1339:1339] = '{32'hc2af8a07};
test_output[1339:1339] = '{32'hc5c07c42};
test_input[10720:10727] = '{32'h42aafb70, 32'hc1b4e131, 32'hc255e754, 32'hc1940d3d, 32'hc1f450ca, 32'h41d10914, 32'hc28d4bba, 32'hc2b7642f};
test_weights[10720:10727] = '{32'hc2a123e2, 32'h3fcdc3da, 32'hc2b6da23, 32'h4246a3c2, 32'h42aa4a53, 32'h4285c3fa, 32'h40fcad7c, 32'h42266a77};
test_bias[1340:1340] = '{32'h400bdf24};
test_output[1340:1340] = '{32'hc5ff8c6f};
test_input[10728:10735] = '{32'hc22c99a7, 32'h42b05dd8, 32'h428a5c59, 32'hc2af76c4, 32'h42aa9c1b, 32'h425819ed, 32'h41808a77, 32'h42b560f0};
test_weights[10728:10735] = '{32'h42599960, 32'h42b75b18, 32'h4216c8ee, 32'h424efd10, 32'hc212a21a, 32'h42073a75, 32'hc25b8460, 32'hc2c72f7e};
test_bias[1341:1341] = '{32'h415b0b5f};
test_output[1341:1341] = '{32'hc5e71db9};
test_input[10736:10743] = '{32'h4299c79e, 32'hc2a3b140, 32'h4241f6aa, 32'hc271f593, 32'hc179cfe0, 32'hc0c4c2b9, 32'hc2c0def6, 32'hc1995d9c};
test_weights[10736:10743] = '{32'hc229ebaa, 32'h42bf04c6, 32'h4118d13d, 32'h42ac42ab, 32'hc2c7619b, 32'hc0aa509e, 32'h423117cf, 32'hc227861b};
test_bias[1342:1342] = '{32'h41ecaa27};
test_output[1342:1342] = '{32'hc68a1c18};
test_input[10744:10751] = '{32'h429ffcb1, 32'h421cc16a, 32'hc26de8c1, 32'h42c1de2b, 32'hc1b3848c, 32'h424dfe9d, 32'hc179f4b4, 32'hc29e50a1};
test_weights[10744:10751] = '{32'h424ae1e5, 32'h42997606, 32'h41f6c1c3, 32'h429872c2, 32'hc2834f23, 32'h42143c26, 32'hc0a6b76b, 32'hc2be6a8a};
test_bias[1343:1343] = '{32'hc25904f8};
test_output[1343:1343] = '{32'h46b81788};
test_input[10752:10759] = '{32'hc297f92f, 32'h4295b1dc, 32'hc1546385, 32'h4215771f, 32'hc2924ea0, 32'hc2c1c44e, 32'h41b70ee1, 32'h4117ec70};
test_weights[10752:10759] = '{32'hc274b781, 32'h42ba3e02, 32'hc209e570, 32'h42966d9f, 32'h42b2ec06, 32'hc26032cf, 32'hc21aecfe, 32'h4255ec63};
test_bias[1344:1344] = '{32'hc2445789};
test_output[1344:1344] = '{32'h4650847d};
test_input[10760:10767] = '{32'hc1a230ff, 32'h41680080, 32'hc28ece9c, 32'h41d9c75c, 32'h4098498b, 32'h4263efe8, 32'h42a4eaeb, 32'h4230e50a};
test_weights[10760:10767] = '{32'hc2a7daa2, 32'h41dc1d31, 32'hc2aecb4b, 32'h4228a1f8, 32'h426e1162, 32'hc281751b, 32'hc26adf86, 32'h4217d743};
test_bias[1345:1345] = '{32'hc1fa7ddb};
test_output[1345:1345] = '{32'h45348e69};
test_input[10768:10775] = '{32'hc1546ae4, 32'h42ae3780, 32'h426ca1cf, 32'h41c44333, 32'h42c5baf7, 32'hc28a8def, 32'hc2b82fb6, 32'hc2425f85};
test_weights[10768:10775] = '{32'hc264386f, 32'h425d1969, 32'hc2a72bfd, 32'hc2afb84e, 32'h42c6277e, 32'hc0b3eaab, 32'hc17be084, 32'hc293d7f1};
test_bias[1346:1346] = '{32'hc2b7dfbf};
test_output[1346:1346] = '{32'h46549b62};
test_input[10776:10783] = '{32'h426ca0a4, 32'h4249d012, 32'h429c6dc6, 32'hc2475852, 32'h41e86d75, 32'h428aa496, 32'hc2807da3, 32'h42651f23};
test_weights[10776:10783] = '{32'hc2ab1463, 32'h4279ee68, 32'h4251ea04, 32'h3dca12b2, 32'hc1e9f315, 32'hc1cd7c2c, 32'hc2aa3f04, 32'h429a54e6};
test_bias[1347:1347] = '{32'hc2839fe6};
test_output[1347:1347] = '{32'h4612a2c9};
test_input[10784:10791] = '{32'h3f25b8fd, 32'h407cab20, 32'hc0442720, 32'hc2b9cf69, 32'hc2ab3010, 32'h4280da7d, 32'hc1547a7b, 32'hc0f6149d};
test_weights[10784:10791] = '{32'hc20a10b8, 32'hc212092e, 32'h4196feed, 32'h417f96ef, 32'h42a06d51, 32'hc03abab8, 32'hc1eea9f5, 32'hc13256ad};
test_bias[1348:1348] = '{32'hc2845a87};
test_output[1348:1348] = '{32'hc60269e0};
test_input[10792:10799] = '{32'h42b8d9e5, 32'h41e0492e, 32'hc260a252, 32'h422fe2dc, 32'hc21a2b4d, 32'h41a343d7, 32'hc21d0469, 32'hc2789146};
test_weights[10792:10799] = '{32'h42025e94, 32'hc2a95c41, 32'hc297f01b, 32'hc239999e, 32'hc2c538db, 32'hc0b0dbd0, 32'hc07a6188, 32'h4132b574};
test_bias[1349:1349] = '{32'hc28d4e40};
test_output[1349:1349] = '{32'h45b9a87b};
test_input[10800:10807] = '{32'hc295be8a, 32'hc139064d, 32'h409e887c, 32'hc1a269ed, 32'hc03068c5, 32'h4185a071, 32'h4290184e, 32'hc1fbdf7c};
test_weights[10800:10807] = '{32'hc2c15ec2, 32'hc290fc1a, 32'h42166fcc, 32'hc0ec9e2e, 32'hc28b9ad5, 32'h425b84cf, 32'h42c71ae5, 32'h42aaaa46};
test_bias[1350:1350] = '{32'h4270e168};
test_output[1350:1350] = '{32'h465bd3ca};
test_input[10808:10815] = '{32'h42892094, 32'hc229d03f, 32'h41adc137, 32'hc2c14f62, 32'h42c10275, 32'h429686bc, 32'h42183fbc, 32'h429e01a7};
test_weights[10808:10815] = '{32'hc03b6980, 32'hc1bab86e, 32'hc2a85c56, 32'hc2a93f56, 32'hc2a525db, 32'h42161480, 32'h42a5473b, 32'h417fcd3c};
test_bias[1351:1351] = '{32'hc0a8c575};
test_output[1351:1351] = '{32'h45c7fb03};
test_input[10816:10823] = '{32'hc18c974f, 32'h40f41052, 32'h411a8300, 32'hbfbdbf68, 32'h4223e477, 32'h3f8870ce, 32'h42871804, 32'h4292c0ae};
test_weights[10816:10823] = '{32'h4279a2ce, 32'h428876c5, 32'hc298489e, 32'hc16dc6f7, 32'h4293092a, 32'h4235549e, 32'hc2bad0ff, 32'h416d4399};
test_bias[1352:1352] = '{32'hc1408d80};
test_output[1352:1352] = '{32'hc55866d2};
test_input[10824:10831] = '{32'h42c48935, 32'hc2106cd6, 32'hc26c7435, 32'hc24560d1, 32'hc2475b74, 32'h4235f566, 32'hc1332c67, 32'hc27ac04f};
test_weights[10824:10831] = '{32'hc28c733e, 32'h42a9809b, 32'h4288f53f, 32'hc18a4a44, 32'hc124b1b7, 32'h3f983f19, 32'hbf025012, 32'h418fa570};
test_bias[1353:1353] = '{32'hc18ef14e};
test_output[1353:1353] = '{32'hc6567a86};
test_input[10832:10839] = '{32'h42521007, 32'h429d3c65, 32'h4248cda4, 32'h4210dd76, 32'h42907724, 32'hc2b7b3ba, 32'hc1b4bb7c, 32'hc197730c};
test_weights[10832:10839] = '{32'hc253918a, 32'hc1a385a6, 32'hc2b438c1, 32'h41d5f9d3, 32'hc1dfb243, 32'hc1b8acd9, 32'h41d950e3, 32'hc2609e6d};
test_bias[1354:1354] = '{32'hc1fab44f};
test_output[1354:1354] = '{32'hc5e7e7fa};
test_input[10840:10847] = '{32'h40f1e013, 32'h41d09d87, 32'h42ae98e7, 32'h428716b7, 32'h41de5010, 32'hc298e59b, 32'h42717c2e, 32'hc265db2d};
test_weights[10840:10847] = '{32'h42b58a0e, 32'hc25b26b7, 32'h40a7a60b, 32'hc0cf43ea, 32'hc1e0b32e, 32'h427e32c2, 32'h42194b7b, 32'hc1a33644};
test_bias[1355:1355] = '{32'h42a3247e};
test_output[1355:1355] = '{32'hc52e9f36};
test_input[10848:10855] = '{32'hc1aec929, 32'h426533d7, 32'h4230b3ed, 32'h418d4e42, 32'h42bd7bfe, 32'h410362aa, 32'h425eb584, 32'h4162520c};
test_weights[10848:10855] = '{32'h4282a5df, 32'h40a8a88b, 32'h4221aafa, 32'hc1c0456f, 32'h429b6c99, 32'h41358470, 32'h4239172e, 32'h4218d1bb};
test_bias[1356:1356] = '{32'h42972430};
test_output[1356:1356] = '{32'h462a0f40};
test_input[10856:10863] = '{32'h42793fde, 32'h4291c659, 32'h4297db37, 32'hc1070f69, 32'h42be22c4, 32'h3e58a2f8, 32'h40ad25aa, 32'h42b2e750};
test_weights[10856:10863] = '{32'h40d55766, 32'h41d2f364, 32'h42515e57, 32'h4280cab9, 32'hc27b1bc6, 32'hc28b0354, 32'h42b2e155, 32'h417ee4ba};
test_bias[1357:1357] = '{32'h4223c4cc};
test_output[1357:1357] = '{32'h44d8e5dd};
test_input[10864:10871] = '{32'h418446ae, 32'hc2b9556d, 32'h42b80826, 32'h415ad9ed, 32'h42a357e3, 32'hc24086fb, 32'h41e471ae, 32'h41d0b034};
test_weights[10864:10871] = '{32'hc12abc83, 32'hc206a093, 32'hc1e28e39, 32'hc28e9047, 32'h42a9673d, 32'h3f7bac47, 32'h4122b9d6, 32'h4290fe8a};
test_bias[1358:1358] = '{32'h3fdd409b};
test_output[1358:1358] = '{32'h46037d33};
test_input[10872:10879] = '{32'hc2460b9a, 32'hc1ae60a9, 32'hc254a4ff, 32'hc15bff82, 32'hc29e3ebf, 32'hc11130cf, 32'hc2c51481, 32'h3fff7992};
test_weights[10872:10879] = '{32'h4210e8d4, 32'h429931e2, 32'h42481421, 32'hc2aa2247, 32'h42b41ae8, 32'hc2887cd0, 32'h42b7a4ef, 32'hc2c394fe};
test_bias[1359:1359] = '{32'hc1810d9a};
test_output[1359:1359] = '{32'hc6a1dc34};
test_input[10880:10887] = '{32'h423b8a27, 32'h425bcdcd, 32'hc22c0ea2, 32'h42c5d8ec, 32'hc2737051, 32'h428e2187, 32'hc2182dea, 32'h42ab629f};
test_weights[10880:10887] = '{32'h41ed8b12, 32'h408993dd, 32'hc28e3b0c, 32'hc2b7e919, 32'h4245680a, 32'h4220b14e, 32'h42a21a20, 32'h42b6b21b};
test_bias[1360:1360] = '{32'h4234a746};
test_output[1360:1360] = '{32'h4367a69c};
test_input[10888:10895] = '{32'hc162484e, 32'h3f99b425, 32'hc2121628, 32'h4236f889, 32'h42afef6e, 32'hc246ba7f, 32'hc2b8c64e, 32'hc246f664};
test_weights[10888:10895] = '{32'hc24034e2, 32'hc21f8470, 32'hc16a7583, 32'hc218a230, 32'hc09b2dea, 32'h423466d7, 32'h4287f9ab, 32'h41d65ab9};
test_bias[1361:1361] = '{32'h42a78190};
test_output[1361:1361] = '{32'hc6286051};
test_input[10896:10903] = '{32'h412afaa8, 32'hc2c23bfe, 32'hc1fc019c, 32'hc2920a27, 32'hc22d2800, 32'h4197d886, 32'h42838273, 32'h42c36959};
test_weights[10896:10903] = '{32'h423b800c, 32'hc2490289, 32'hc2458017, 32'hc292eddc, 32'h41813cc9, 32'h4241c470, 32'hc0cfe05c, 32'hc209aa8f};
test_bias[1362:1362] = '{32'hc2abebd7};
test_output[1362:1362] = '{32'h46071566};
test_input[10904:10911] = '{32'h415c032a, 32'hc2915f37, 32'h42b4bee8, 32'h413e87ee, 32'hc130ddab, 32'h42747b8b, 32'h42ab5c52, 32'hc2c07749};
test_weights[10904:10911] = '{32'hc20d4583, 32'hc09044cd, 32'hc26f16cf, 32'h410f2597, 32'h42a27db4, 32'hc2c7b6be, 32'h4278d8fb, 32'h42a781da};
test_bias[1363:1363] = '{32'hc28f34ca};
test_output[1363:1363] = '{32'hc66e5eff};
test_input[10912:10919] = '{32'h41808b0a, 32'hc162ab3f, 32'hc29ca54e, 32'h42798119, 32'hc22cff5a, 32'h42b6bf6b, 32'hc195614f, 32'hc1cfab97};
test_weights[10912:10919] = '{32'hc224aed7, 32'hc282f563, 32'hc14e1883, 32'hc223e559, 32'hc2ad9a32, 32'h42c21437, 32'hc1e53494, 32'hc120da87};
test_bias[1364:1364] = '{32'hc1898c3c};
test_output[1364:1364] = '{32'h463d5ba7};
test_input[10920:10927] = '{32'h422b649c, 32'h41399921, 32'h4120044c, 32'h42ba1bd9, 32'h421a9af1, 32'hbf1b674b, 32'hc2a7edc5, 32'hc1ba1106};
test_weights[10920:10927] = '{32'hc295cf13, 32'h41daa645, 32'hc1c0c7bd, 32'h42b81515, 32'hc18e024e, 32'hc1301ad0, 32'hc2ab17d8, 32'h41a775dc};
test_bias[1365:1365] = '{32'hc280a681};
test_output[1365:1365] = '{32'h4631de71};
test_input[10928:10935] = '{32'hc04f7314, 32'hc1bdad13, 32'hc1e54448, 32'h416c6241, 32'h420d597b, 32'h42c4aa69, 32'h3ea7d39c, 32'hc1f3d800};
test_weights[10928:10935] = '{32'h41e97d1d, 32'hc2c54783, 32'hc2427660, 32'hbf589878, 32'h42aacd97, 32'hc2a801a9, 32'h419cccd5, 32'hc26aaee2};
test_bias[1366:1366] = '{32'h4295e5f3};
test_output[1366:1366] = '{32'h437c1d3c};
test_input[10936:10943] = '{32'h41ad6cd1, 32'h42ae0c36, 32'h42b63f34, 32'h4244eb50, 32'h42432a0f, 32'hc2125df4, 32'h42612c69, 32'h429ab840};
test_weights[10936:10943] = '{32'hc2818bac, 32'h42af8d45, 32'h40b34a9c, 32'hc25f53ed, 32'h42b64342, 32'h4288a397, 32'h428d3583, 32'hc0eb8c32};
test_bias[1367:1367] = '{32'hc282635f};
test_output[1367:1367] = '{32'h46110b37};
test_input[10944:10951] = '{32'hc11854d5, 32'hc19f26d3, 32'hc0bb2de6, 32'h42921a4e, 32'hc2b79f4c, 32'h41c23b69, 32'h422b10b0, 32'h42855140};
test_weights[10944:10951] = '{32'hc0d6e428, 32'h42879103, 32'h41f8dd13, 32'h411f1c8d, 32'h42b2affc, 32'hc2767906, 32'h42bad5c4, 32'h428e3217};
test_bias[1368:1368] = '{32'h421110a0};
test_output[1368:1368] = '{32'hc4d084b0};
test_input[10952:10959] = '{32'h41ef89e4, 32'h42c19176, 32'h4131593a, 32'h4102680f, 32'hc1b6e672, 32'hc16e306e, 32'hc110aebd, 32'h429ba672};
test_weights[10952:10959] = '{32'hbebb9a00, 32'h42a296c5, 32'h426da6c4, 32'h427847d6, 32'hc1f3698d, 32'hc282a54d, 32'hc27fab7b, 32'hc27ebe0b};
test_bias[1369:1369] = '{32'h4269f794};
test_output[1369:1369] = '{32'h45c70da1};
test_input[10960:10967] = '{32'h413cdcce, 32'h41b77a40, 32'h429e10be, 32'hc1b2505b, 32'hc0ab32d2, 32'hc25208f8, 32'hc21bf8c8, 32'hc296e491};
test_weights[10960:10967] = '{32'hc1e45654, 32'h4260f175, 32'hc2b5ee52, 32'hc2884244, 32'hc18397f1, 32'hc005b28e, 32'h410f0bd9, 32'hc28f4c96};
test_bias[1370:1370] = '{32'h4179e0b0};
test_output[1370:1370] = '{32'h440a2351};
test_input[10968:10975] = '{32'hc2722062, 32'h40841979, 32'h3f1ddc8b, 32'hc07c8da3, 32'h424bc303, 32'hc29c708c, 32'hc1efe9fc, 32'h4210304d};
test_weights[10968:10975] = '{32'hc1c8b4ba, 32'hc27f83a8, 32'h42761c5c, 32'hc294647a, 32'hc2a918c7, 32'h426c0818, 32'h42affb5e, 32'hc216b2f6};
test_bias[1371:1371] = '{32'h42a3c61d};
test_output[1371:1371] = '{32'hc62fcf48};
test_input[10976:10983] = '{32'h42784f34, 32'hc291fb9f, 32'h421f3e48, 32'hc2b661f6, 32'h41b9ba9f, 32'h41697b38, 32'h4299368b, 32'hc2b3d1e7};
test_weights[10976:10983] = '{32'hc28aa757, 32'h40a0cc9c, 32'hc29daab0, 32'hc269b669, 32'h427a5eeb, 32'h40997c9b, 32'h4261fbc8, 32'hc0b62e1d};
test_bias[1372:1372] = '{32'hc28a2479};
test_output[1372:1372] = '{32'h456e5370};
test_input[10984:10991] = '{32'h41ac4831, 32'h4284e2ef, 32'h424d46d4, 32'hc2989e02, 32'h41436b57, 32'hc2b3fc6d, 32'hc267f3b1, 32'h425eed1b};
test_weights[10984:10991] = '{32'h408fc856, 32'h42097fe0, 32'h420c689a, 32'h427f994c, 32'h42b3d935, 32'hc2494f21, 32'hc1f8e166, 32'hc28e7235};
test_bias[1373:1373] = '{32'h41797aa2};
test_output[1373:1373] = '{32'h452dfb2a};
test_input[10992:10999] = '{32'hc26b6091, 32'hc2584a41, 32'h423be6c2, 32'h428508fc, 32'hc2aef85e, 32'hc22a92ad, 32'h42914de4, 32'hc24fd901};
test_weights[10992:10999] = '{32'h418b8c90, 32'hc0946c32, 32'h4249925f, 32'hc26da78c, 32'hc1e31baf, 32'h42093c45, 32'hc1b4734f, 32'h413f0006};
test_bias[1374:1374] = '{32'hc29db089};
test_output[1374:1374] = '{32'hc565ddaa};
test_input[11000:11007] = '{32'hc28bda1f, 32'h4280e211, 32'hc24eef67, 32'h429fab4b, 32'hc2910cb8, 32'hc274a114, 32'h4190d87d, 32'hc28fef84};
test_weights[11000:11007] = '{32'h429a3963, 32'hc264b52a, 32'hc18d9e9a, 32'hc21d1e26, 32'h41de16c3, 32'h423dc73f, 32'h42aa60fb, 32'h423625ac};
test_bias[1375:1375] = '{32'h41a42d91};
test_output[1375:1375] = '{32'hc68c0be7};
test_input[11008:11015] = '{32'h42ade561, 32'h418d4f51, 32'hc1b99d2e, 32'hc2bcdce0, 32'hc1c6e615, 32'h3c5a992f, 32'hc2a736ea, 32'hc2a6a703};
test_weights[11008:11015] = '{32'h42936d1e, 32'hc26a6a79, 32'hc22aae1d, 32'h4180a14b, 32'h41fe9e35, 32'h42ad0136, 32'h423a5a5c, 32'hc2261e8e};
test_bias[1376:1376] = '{32'h42811c38};
test_output[1376:1376] = '{32'h456658ab};
test_input[11016:11023] = '{32'h41641609, 32'hc27177be, 32'h429fcba7, 32'h418e1530, 32'h425a179b, 32'hc2159209, 32'h423ce349, 32'h420457a6};
test_weights[11016:11023] = '{32'h41db0cf2, 32'hc18d6695, 32'hc0fa871a, 32'hc1c6caf7, 32'h41fd580e, 32'hc24c23ea, 32'h4001c404, 32'hc297c35c};
test_bias[1377:1377] = '{32'h41389372};
test_output[1377:1377] = '{32'h44cac484};
test_input[11024:11031] = '{32'hc1cf80f5, 32'h424b76e0, 32'h4231a1b4, 32'hc26f25e9, 32'hc0cb4caf, 32'h41d64a33, 32'hc1f75c9d, 32'h41799ea8};
test_weights[11024:11031] = '{32'h4178d02a, 32'hc2bcc2b6, 32'hc19b978c, 32'h429b94cc, 32'h4232e67a, 32'h426729b5, 32'h422f441a, 32'hc2bf628f};
test_bias[1378:1378] = '{32'h42a1a0af};
test_output[1378:1378] = '{32'hc63ef6f9};
test_input[11032:11039] = '{32'hc298e19b, 32'h42286c09, 32'hc1d59ed7, 32'h4239a013, 32'h4194626b, 32'h415e6031, 32'h41a00e3d, 32'h422ee5a9};
test_weights[11032:11039] = '{32'h42b1ab9a, 32'h4298cdf5, 32'h42b9d93a, 32'hc2c2f48f, 32'h42bcc435, 32'hc273f0d3, 32'h420c37de, 32'hc2b5dded};
test_bias[1379:1379] = '{32'hc2929e27};
test_output[1379:1379] = '{32'hc64b7e05};
test_input[11040:11047] = '{32'hc204cb89, 32'h42aa0f95, 32'h423fd443, 32'hc18271ee, 32'hc24c2e00, 32'h428930c7, 32'hc2c295ef, 32'hc283a9c5};
test_weights[11040:11047] = '{32'h419c5ea3, 32'hc113254c, 32'hc2aa8ccd, 32'hbf51a48c, 32'h41e880b8, 32'h41386aea, 32'h42b2a496, 32'h41ed0d69};
test_bias[1380:1380] = '{32'h41e0969c};
test_output[1380:1380] = '{32'hc68359e0};
test_input[11048:11055] = '{32'hc18f962e, 32'hc0dc87c3, 32'h416016be, 32'h40888d5a, 32'hbfc69d46, 32'hc1f66cd5, 32'h40d9faae, 32'h428fa61a};
test_weights[11048:11055] = '{32'hc1dddc8f, 32'hc28b81c9, 32'h4296fcdd, 32'h4228991a, 32'h4284f94e, 32'h429c1101, 32'hc2ac1a91, 32'h42aecc46};
test_bias[1381:1381] = '{32'hbdba5efa};
test_output[1381:1381] = '{32'h45a8bf91};
test_input[11056:11063] = '{32'hc1194012, 32'hc2b6e252, 32'hc2aaa131, 32'hc2709fd5, 32'hc2200af4, 32'hc1320273, 32'h42b402c0, 32'hc2396527};
test_weights[11056:11063] = '{32'hc008f8ff, 32'hc1f64753, 32'h42b91474, 32'h41e879a2, 32'hc283fcab, 32'hc1ae6ab7, 32'h4191ed71, 32'hc1444a24};
test_bias[1382:1382] = '{32'h42ab702f};
test_output[1382:1382] = '{32'hc4cb8f74};
test_input[11064:11071] = '{32'h42af7c3f, 32'h42573463, 32'h419dc645, 32'h4227caa8, 32'hc2c146b3, 32'h423539e0, 32'hc0a160dd, 32'hc29e9374};
test_weights[11064:11071] = '{32'hc0c90310, 32'h42b31d6f, 32'hc2a552ab, 32'hc1ad9681, 32'hc2b643cf, 32'h4193e521, 32'h40a2e412, 32'hbf8a6104};
test_bias[1383:1383] = '{32'hc236aea6};
test_output[1383:1383] = '{32'h4631e607};
test_input[11072:11079] = '{32'hc03c21a4, 32'hc2adbb60, 32'hc2c6fcb8, 32'h421d7ba8, 32'hc2a02b09, 32'hbf4449c8, 32'hc27ec567, 32'h423f9b73};
test_weights[11072:11079] = '{32'h42046350, 32'h42be4aa9, 32'hc2b135b5, 32'h41971ade, 32'hc28f2645, 32'h42c7c061, 32'hc2a42346, 32'h42c1b858};
test_bias[1384:1384] = '{32'hc2921848};
test_output[1384:1384] = '{32'h46820cbe};
test_input[11080:11087] = '{32'hc0f48f11, 32'hc28f972c, 32'h427e260a, 32'hc19f4df8, 32'hc2c5b978, 32'h42120ff1, 32'hc2b9bb46, 32'hc2a6b4c4};
test_weights[11080:11087] = '{32'hc2c42345, 32'hc27c08b6, 32'hc1a2def7, 32'hc179725d, 32'hc265b2ac, 32'h411111d9, 32'h4223f39b, 32'hc14a1ffc};
test_bias[1385:1385] = '{32'h4218138d};
test_output[1385:1385] = '{32'h45ecf777};
test_input[11088:11095] = '{32'hc2a7a4b7, 32'hc209c2ad, 32'hc1fd7ff2, 32'h42b25683, 32'hc256943e, 32'hc24d0f47, 32'h42550b7f, 32'h41c36285};
test_weights[11088:11095] = '{32'h42563018, 32'hc21bede9, 32'hc26d61f7, 32'hc1a6cf6a, 32'hc24aa2d3, 32'hc1e66a00, 32'hc2a8427b, 32'hc2290d73};
test_bias[1386:1386] = '{32'h41905ab7};
test_output[1386:1386] = '{32'hc58a4c20};
test_input[11096:11103] = '{32'hc1f8019c, 32'hc2824025, 32'hc276b4e2, 32'h4220b337, 32'hc2260950, 32'hc1a273f9, 32'h4162872a, 32'h42718cf1};
test_weights[11096:11103] = '{32'hc1b6ad53, 32'h41764a17, 32'h4237e783, 32'h41572bc1, 32'h40f9e338, 32'h420fbdae, 32'h41cebb20, 32'h42c228eb};
test_bias[1387:1387] = '{32'h404c4d5d};
test_output[1387:1387] = '{32'h4521ba80};
test_input[11104:11111] = '{32'hc21d0876, 32'h4286ffaa, 32'h424fe642, 32'hc237c71c, 32'h423499ba, 32'hc29b8fbf, 32'hc22e1b73, 32'h41be69c0};
test_weights[11104:11111] = '{32'h428b6644, 32'h427e1f8d, 32'hc2674666, 32'hc19b57b7, 32'hc2896040, 32'hc29c5495, 32'h4227ac4f, 32'h41f31b2e};
test_bias[1388:1388] = '{32'hc258e4d4};
test_output[1388:1388] = '{32'h449dbfca};
test_input[11112:11119] = '{32'h428519ce, 32'hc2b33040, 32'hc2c143ff, 32'h429286f5, 32'h4294ad5c, 32'hc1d496f2, 32'h41f84faf, 32'hc2b4e01a};
test_weights[11112:11119] = '{32'h42419044, 32'hc19c0b48, 32'hc2a8074e, 32'h42bad887, 32'h400eef0b, 32'h426a5040, 32'hc27aed36, 32'h4218ad24};
test_bias[1389:1389] = '{32'h40e3c274};
test_output[1389:1389] = '{32'h464d71fc};
test_input[11120:11127] = '{32'hc2bcfc1c, 32'h429fb889, 32'h41b30214, 32'h41aeb294, 32'hc23655d7, 32'h4171e938, 32'hc2bdd3f2, 32'h40eeaa5d};
test_weights[11120:11127] = '{32'h4298d7f3, 32'h423e5874, 32'h429d64fa, 32'h4159e913, 32'hc215461b, 32'hc240e4da, 32'h413d9ad3, 32'hc293edff};
test_bias[1390:1390] = '{32'h428a491a};
test_output[1390:1390] = '{32'hc4f9bdc3};
test_input[11128:11135] = '{32'hc2b040e6, 32'h425f815e, 32'hc2c7f23c, 32'h428b9277, 32'hc22f4f3d, 32'hc15e89f7, 32'h423ba807, 32'hc2aef47e};
test_weights[11128:11135] = '{32'hc2048aad, 32'h41807cc3, 32'hc21bce13, 32'h40bcc2db, 32'hc21cba3b, 32'hc2be9c74, 32'hc1aeb1ed, 32'h42c60b1e};
test_bias[1391:1391] = '{32'h42a44aa0};
test_output[1391:1391] = '{32'h44c3333a};
test_input[11136:11143] = '{32'h429c3fed, 32'hc28658b0, 32'hc1800d82, 32'h4279a96c, 32'h41771b2a, 32'h41d3fb2e, 32'hc21bc4ed, 32'h41d1b61a};
test_weights[11136:11143] = '{32'h42a0dbc1, 32'hc1e754ed, 32'hc2bec212, 32'h42829975, 32'h4282ead1, 32'hc0acce9e, 32'hc2630fce, 32'h42906783};
test_bias[1392:1392] = '{32'h42553400};
test_output[1392:1392] = '{32'h4693498d};
test_input[11144:11151] = '{32'hc22a9aaa, 32'hc09be1f5, 32'h42a60e40, 32'hc29c7ed3, 32'hc2a15003, 32'hc2819f05, 32'h4293576c, 32'h41e79034};
test_weights[11144:11151] = '{32'h42b5b5bb, 32'h4206a0d4, 32'hc252b7ee, 32'h4222edc6, 32'hc249069a, 32'hc1a98d9f, 32'h424cb1a0, 32'hc1a6f24e};
test_bias[1393:1393] = '{32'h4261e649};
test_output[1393:1393] = '{32'hc538690d};
test_input[11152:11159] = '{32'h42bac359, 32'h420e76f2, 32'hc21b0d98, 32'h428ec316, 32'hc294655d, 32'h415384b3, 32'h4249b0d1, 32'h41b25196};
test_weights[11152:11159] = '{32'h42154bed, 32'h42c0fed4, 32'h4211eb9c, 32'hc289cd10, 32'hc23ee0b3, 32'hc2b44613, 32'h42c7b21c, 32'hc24029c8};
test_bias[1394:1394] = '{32'h4269f875};
test_output[1394:1394] = '{32'h45d98ab8};
test_input[11160:11167] = '{32'h42bf0215, 32'hc2798719, 32'h42450a9b, 32'h4200438d, 32'hc1ce6222, 32'h4259aa06, 32'h41046688, 32'hc0449097};
test_weights[11160:11167] = '{32'h4217b8f1, 32'h420c9c32, 32'hc2978eb2, 32'h401174a6, 32'hc218c790, 32'hc2a4ae99, 32'hc282ab43, 32'h42a656ee};
test_bias[1395:1395] = '{32'hc24a651a};
test_output[1395:1395] = '{32'hc5cd62fa};
test_input[11168:11175] = '{32'h42912249, 32'hc20abaa8, 32'hc2b3f438, 32'h42bf576b, 32'hc262cde0, 32'hc2696737, 32'h42a10e3e, 32'hc1a57bbd};
test_weights[11168:11175] = '{32'hc2ae71bb, 32'hc200a9c6, 32'hc14c3bc1, 32'hc29e5b75, 32'h42981fd3, 32'hc20fdd26, 32'hc18f3cf8, 32'h422e1877};
test_bias[1396:1396] = '{32'hc15463c4};
test_output[1396:1396] = '{32'hc67d47fe};
test_input[11176:11183] = '{32'h428f72da, 32'hc250e45e, 32'hc2902db3, 32'h429ae93e, 32'hc286b8f1, 32'hc264be0d, 32'h41d36112, 32'hc1106008};
test_weights[11176:11183] = '{32'hc21c20af, 32'h42ac476a, 32'hc29c0d0e, 32'h40b9d730, 32'hc2b7db3a, 32'hc23d4d47, 32'h428dd9d9, 32'h41931e5b};
test_bias[1397:1397] = '{32'hc2a19b29};
test_output[1397:1397] = '{32'h46115a86};
test_input[11184:11191] = '{32'h4283cceb, 32'h428bffb5, 32'hc27ba3a2, 32'h42c38478, 32'hc2916650, 32'h428de4e4, 32'h4281b7bb, 32'hc2806183};
test_weights[11184:11191] = '{32'hc1c1e92f, 32'h420030eb, 32'h42980571, 32'h4266d06a, 32'h426d287c, 32'hc2c3111f, 32'h4204c85c, 32'h42859ef3};
test_bias[1398:1398] = '{32'hc2b2a3b3};
test_output[1398:1398] = '{32'hc63ab6f5};
test_input[11192:11199] = '{32'h42b6f3fc, 32'h42b7e0aa, 32'hc2aafd73, 32'h4235fa5b, 32'hc035e929, 32'hc296f4b4, 32'hc22135c3, 32'hc1d82594};
test_weights[11192:11199] = '{32'hc2419e91, 32'hc12ba099, 32'hc1c99fce, 32'hc2417aaa, 32'h4284fdad, 32'h4273f80c, 32'h420e214a, 32'h41fafee4};
test_bias[1399:1399] = '{32'h418f238c};
test_output[1399:1399] = '{32'hc6438965};
test_input[11200:11207] = '{32'h42a56ebd, 32'h410b1878, 32'h427e26ac, 32'h42a7f304, 32'hc2702b80, 32'h429e2a89, 32'hc2c300fc, 32'h42a7c88c};
test_weights[11200:11207] = '{32'hc1d0ed0b, 32'hc204324b, 32'hc1b5a08e, 32'hc2567a5b, 32'hc2126611, 32'h427cacb8, 32'h42a3a155, 32'hc115256c};
test_bias[1400:1400] = '{32'h41b48c07};
test_output[1400:1400] = '{32'hc61b40af};
test_input[11208:11215] = '{32'h422c609f, 32'hc2bf97de, 32'hc2308228, 32'hc1b99d8d, 32'h429bb27d, 32'hc293ad01, 32'h42c69f72, 32'hc2291eb2};
test_weights[11208:11215] = '{32'hc1ff3617, 32'hc1debd3a, 32'hc274d404, 32'h42c1a386, 32'hc2430912, 32'h428bd506, 32'h423c60cc, 32'hc0ad088e};
test_bias[1401:1401] = '{32'h42391024};
test_output[1401:1401] = '{32'hc50d36c8};
test_input[11216:11223] = '{32'h42b47b77, 32'hc2c67733, 32'h42015aa6, 32'h42c71c81, 32'hc2905e54, 32'h41a1eb0b, 32'h423b3282, 32'h427b871a};
test_weights[11216:11223] = '{32'hc28eedb9, 32'h3ef575b0, 32'h40e7387f, 32'h42403ff9, 32'hc2963ed2, 32'h42bc0575, 32'h414494a0, 32'hc21ee897};
test_bias[1402:1402] = '{32'hc270846c};
test_output[1402:1402] = '{32'h45718222};
test_input[11224:11231] = '{32'hc287ae2b, 32'h41c53fea, 32'hc28e1588, 32'hc2bec025, 32'hc2066fe0, 32'hc24c3b4c, 32'hc2677152, 32'hc0ae8379};
test_weights[11224:11231] = '{32'hc239bbf2, 32'h4286b81d, 32'h4276d0ef, 32'h40f777cb, 32'h42a57718, 32'hc2696856, 32'h42b0a15d, 32'h42883700};
test_bias[1403:1403] = '{32'hc2519be5};
test_output[1403:1403] = '{32'hc5b06a94};
test_input[11232:11239] = '{32'hc23a9515, 32'h429ffa13, 32'h41f053fd, 32'h428eb54c, 32'h42283be3, 32'hc2ac00e1, 32'h4219ba8c, 32'h40f02d3a};
test_weights[11232:11239] = '{32'hc1c4c768, 32'hc1eeaded, 32'h42bb043a, 32'h418c40c1, 32'hc2229931, 32'hc119355c, 32'h4071c538, 32'h4142f902};
test_bias[1404:1404] = '{32'h4206cc56};
test_output[1404:1404] = '{32'h4509d23e};
test_input[11240:11247] = '{32'hc25efd7b, 32'h420bd637, 32'h404670bc, 32'hc254b184, 32'h421d55cc, 32'h42b04d88, 32'hc2bcdb82, 32'hc2140956};
test_weights[11240:11247] = '{32'h427fe7f9, 32'hc1607765, 32'hc23e5e69, 32'h429152c4, 32'h42b8747a, 32'h4273977e, 32'hc2b4f5b1, 32'h42a6a195};
test_bias[1405:1405] = '{32'hc26deb90};
test_output[1405:1405] = '{32'h45c5c557};
test_input[11248:11255] = '{32'hc2774025, 32'h419bc1b0, 32'h417df022, 32'h4207843a, 32'hc2925933, 32'hc2bda928, 32'hc02e08c7, 32'h411aa5ec};
test_weights[11248:11255] = '{32'h424a7303, 32'hc2743f95, 32'h426d1c5f, 32'hc1d67f4e, 32'hc23a5c93, 32'h429b622c, 32'hc1e24cd1, 32'h4267bb96};
test_bias[1406:1406] = '{32'hc0cbfe54};
test_output[1406:1406] = '{32'hc5ede5c8};
test_input[11256:11263] = '{32'hc0f256f2, 32'h4238d37e, 32'hc2bdbe0d, 32'hc24c5e0c, 32'hc23a4350, 32'hc2bca995, 32'h42b4a3fd, 32'hc2a288eb};
test_weights[11256:11263] = '{32'h4293824a, 32'h421aeb6a, 32'hc28dca5d, 32'hbd8ce456, 32'h41ebf402, 32'h4294a8de, 32'hc231f877, 32'hc115207d};
test_bias[1407:1407] = '{32'hc287d0a3};
test_output[1407:1407] = '{32'hc56a9a21};
test_input[11264:11271] = '{32'hc1fd1bdc, 32'hc2c261b8, 32'h415845a1, 32'h425b8eac, 32'h3f3253fd, 32'hc28b12c1, 32'hc24eb626, 32'hc263a217};
test_weights[11264:11271] = '{32'h428a0ab1, 32'h41a29cdd, 32'h42c22ac8, 32'h41a93151, 32'h421d4bff, 32'hc2c51f48, 32'h41ba7039, 32'hc2afd9c4};
test_bias[1408:1408] = '{32'hc2962caa};
test_output[1408:1408] = '{32'h460b5c6a};
test_input[11272:11279] = '{32'h428b4e0f, 32'h42923134, 32'hc181dd2d, 32'hc27480a2, 32'h42be33c0, 32'hc28750ff, 32'h41fed82d, 32'h41d3a09c};
test_weights[11272:11279] = '{32'hc294cd08, 32'hc27c5181, 32'h422b7342, 32'hc29604bc, 32'h423d9ffd, 32'hc24a119d, 32'hc28d4c2f, 32'hc2c6e409};
test_bias[1409:1409] = '{32'h4235d5cf};
test_output[1409:1409] = '{32'hc52fd544};
test_input[11280:11287] = '{32'h429fd17a, 32'hc0db3780, 32'h42b46820, 32'hc2c33100, 32'hc286ffa1, 32'h4284f2f0, 32'hc10aff98, 32'hc288cffb};
test_weights[11280:11287] = '{32'hc2056541, 32'h42b088b3, 32'hc2a41fda, 32'hc2104a41, 32'hc2992b95, 32'hc0afd26b, 32'h427fc870, 32'hc18ecade};
test_bias[1410:1410] = '{32'hc27441fb};
test_output[1410:1410] = '{32'hc4d9d711};
test_input[11288:11295] = '{32'h41d93787, 32'hc24db6bf, 32'hc28e1936, 32'h42bc3439, 32'h425ac271, 32'h429156af, 32'h419c62f7, 32'hc247bb29};
test_weights[11288:11295] = '{32'hc2b59125, 32'hc0d56b4d, 32'hc2c7d395, 32'hc2084896, 32'h42c3aee2, 32'h4132d920, 32'h42358976, 32'hc241b36e};
test_bias[1411:1411] = '{32'hbf70e3e1};
test_output[1411:1411] = '{32'h462f9896};
test_input[11296:11303] = '{32'h41fdc3f2, 32'hc18f4e93, 32'hc23a0908, 32'h42947c31, 32'h428be8a6, 32'h426a7f0b, 32'hc2c14d88, 32'h4253afcc};
test_weights[11296:11303] = '{32'hc2a76109, 32'h4260d969, 32'h41e914cf, 32'hc21d172a, 32'hc163c27f, 32'h4241f7c7, 32'hc2ac0cbd, 32'hc1d46e32};
test_bias[1412:1412] = '{32'h42796f82};
test_output[1412:1412] = '{32'h445d8847};
test_input[11304:11311] = '{32'hc2a5228e, 32'h42965cb0, 32'h428c57ba, 32'hc2558413, 32'hc0a88591, 32'hc28c9a3f, 32'hc25a1fd8, 32'hc20dc989};
test_weights[11304:11311] = '{32'hc22d34c5, 32'h4293f52d, 32'h42b5de1a, 32'h422e2739, 32'hc28e91d3, 32'hc102dc17, 32'hc29c2360, 32'hc2994018};
test_bias[1413:1413] = '{32'hc2a42193};
test_output[1413:1413] = '{32'h46a4574d};
test_input[11312:11319] = '{32'hc22aacec, 32'hc155e68a, 32'hc221c98c, 32'h42c7d2e8, 32'hc2555f29, 32'hc23e8137, 32'h41cae6c7, 32'h4211c006};
test_weights[11312:11319] = '{32'h429172c9, 32'h42b428e3, 32'h4290d6d9, 32'hc2430c3d, 32'h421598d0, 32'h42834cd8, 32'h400cb097, 32'h429a9738};
test_bias[1414:1414] = '{32'h41e88ec5};
test_output[1414:1414] = '{32'hc65fe2ef};
test_input[11320:11327] = '{32'hc299e616, 32'hc26683fd, 32'hc2aa1a13, 32'hc2264bb7, 32'hc2624bee, 32'h42944bb7, 32'hc2577473, 32'hc1a3a82a};
test_weights[11320:11327] = '{32'h42921115, 32'h4218fb46, 32'hc2b231aa, 32'hc24743e2, 32'hc2bbfdfe, 32'hc289974f, 32'h4212e457, 32'hc252ec83};
test_bias[1415:1415] = '{32'h4048486e};
test_output[1415:1415] = '{32'h448f2e76};
test_input[11328:11335] = '{32'hc13ab031, 32'hc28d0617, 32'hc18eebca, 32'h4169c33f, 32'hc1c9027a, 32'h40f8af11, 32'h42044b52, 32'hc18ca326};
test_weights[11328:11335] = '{32'hc18f1382, 32'h42b549ad, 32'hc289dd72, 32'h42b977a1, 32'hc1692612, 32'hc2b5249a, 32'h42acc92d, 32'hc2bda500};
test_bias[1416:1416] = '{32'h42973f6e};
test_output[1416:1416] = '{32'h44266d10};
test_input[11336:11343] = '{32'hc2409a8c, 32'hc27b34e3, 32'h413b1919, 32'h418ae055, 32'h424b4c42, 32'h42b6d6b5, 32'hc1927c6d, 32'hc2ba6b6a};
test_weights[11336:11343] = '{32'hc1ee766c, 32'hc2ad83df, 32'h42c3dee0, 32'h418a2cca, 32'h414e5660, 32'hc290d3b5, 32'h4207d2b4, 32'hc2acfdd5};
test_bias[1417:1417] = '{32'h428ba73a};
test_output[1417:1417] = '{32'h461a4a6e};
test_input[11344:11351] = '{32'hc2881e8b, 32'h424a6b20, 32'h401acf04, 32'hc24669eb, 32'h4006d9ee, 32'hc2aa7652, 32'h4223fe1f, 32'h42a3bf33};
test_weights[11344:11351] = '{32'h422c176a, 32'h42546615, 32'h42a3fd79, 32'hc2c46801, 32'h41a47cec, 32'hc28b2f88, 32'hc22c81e5, 32'hc29cc2fe};
test_bias[1418:1418] = '{32'h42abd840};
test_output[1418:1418] = '{32'h4528fce6};
test_input[11352:11359] = '{32'hc1a19e58, 32'h42be04a5, 32'hc26bf23a, 32'hc207f62c, 32'h409fa184, 32'h42825d04, 32'h4203a81a, 32'hc2a858b8};
test_weights[11352:11359] = '{32'h410fe423, 32'hc094b36f, 32'hc29209e0, 32'hc2c21bb6, 32'h42a35980, 32'h41f2ffb5, 32'hc23ab9f7, 32'hc053298d};
test_bias[1419:1419] = '{32'h428cfab0};
test_output[1419:1419] = '{32'h45ffaf66};
test_input[11360:11367] = '{32'h42b90475, 32'h42c22a02, 32'hc1d59bad, 32'hc1a95389, 32'hc1706b2e, 32'hc2c0e3c2, 32'hc26d51dd, 32'hc1c97f39};
test_weights[11360:11367] = '{32'hc2607322, 32'h4289c7ba, 32'h429f4076, 32'hc1bd488a, 32'h42a8c714, 32'hc22ce2b5, 32'h40f63310, 32'h428b7ded};
test_bias[1420:1420] = '{32'h4202449d};
test_output[1420:1420] = '{32'h4413e8f9};
test_input[11368:11375] = '{32'hc1838355, 32'hc09bf204, 32'h42b4218c, 32'h42bcbcd3, 32'hc0783a60, 32'h410c7f61, 32'hc192d732, 32'h4295b89d};
test_weights[11368:11375] = '{32'hc1883c12, 32'h3fa0880c, 32'h41a11568, 32'hc2721f8a, 32'h4202e7ef, 32'h41dbc270, 32'hc27eaa42, 32'hc292eb88};
test_bias[1421:1421] = '{32'hc2bf554a};
test_output[1421:1421] = '{32'hc5f80753};
test_input[11376:11383] = '{32'h41be6b7e, 32'hc1fa63b1, 32'hc21b0581, 32'h42041646, 32'hc0d8f0fd, 32'h4234092a, 32'hc20080c8, 32'hc115947e};
test_weights[11376:11383] = '{32'h427b8dfa, 32'hc2a1d7fa, 32'hc2a2f337, 32'h42c4f7cf, 32'hc1a765a7, 32'hc21db843, 32'h4285fa06, 32'hc24a75c5};
test_bias[1422:1422] = '{32'h42275a66};
test_output[1422:1422] = '{32'h45e00bf1};
test_input[11384:11391] = '{32'hc1c0232b, 32'h411827c6, 32'hc1ac81e0, 32'hc23a7b87, 32'hc09468e7, 32'hc1e1525f, 32'h4135597f, 32'h42bc8a78};
test_weights[11384:11391] = '{32'hc19c70c1, 32'hc25d6f4a, 32'h42bb4ecc, 32'hc28e4173, 32'hbf88d1f5, 32'hc27fb243, 32'hc1c9d0fd, 32'h42921f1a};
test_bias[1423:1423] = '{32'hc223d103};
test_output[1423:1423] = '{32'h461616dc};
test_input[11392:11399] = '{32'hc1354b1d, 32'h42a12ab7, 32'h429e27a1, 32'h42b23a2a, 32'hc2665b4b, 32'hc2a3e0f3, 32'hc293c9c3, 32'h41d70760};
test_weights[11392:11399] = '{32'hc1137a44, 32'hc22f859b, 32'hc2be62d2, 32'h425d503d, 32'hc22cf328, 32'h3fd15a10, 32'hc150f610, 32'hc28c2aed};
test_bias[1424:1424] = '{32'hc230fd0d};
test_output[1424:1424] = '{32'hc590dd3b};
test_input[11400:11407] = '{32'h42c2d3dd, 32'hc2affefb, 32'h42c74557, 32'h425d83b4, 32'h41fafdcc, 32'h3fb2bbfa, 32'hc25bd214, 32'h427d9cb0};
test_weights[11400:11407] = '{32'hc0e0e65c, 32'hc2aef366, 32'h4264050e, 32'hc2b624dd, 32'hc2390601, 32'h4202880b, 32'h42425e83, 32'h42328653};
test_bias[1425:1425] = '{32'h40a976bb};
test_output[1425:1425] = '{32'h45c84245};
test_input[11408:11415] = '{32'hc243673f, 32'h425ab072, 32'hc2b2da27, 32'hc0596bda, 32'hc2c134ca, 32'h428c8122, 32'hc2686f22, 32'h42648b89};
test_weights[11408:11415] = '{32'h4258b054, 32'h41d31700, 32'hc2a2680c, 32'h41a26232, 32'h42a7031e, 32'hc14bcae7, 32'h424df7c2, 32'hc2477f9e};
test_bias[1426:1426] = '{32'hc21d1524};
test_output[1426:1426] = '{32'hc60a574e};
test_input[11416:11423] = '{32'h4208b91a, 32'hc266c51e, 32'h4214d545, 32'hc2a3b212, 32'hc24f9da8, 32'hc213b3b9, 32'h41c4388f, 32'h42a9bef0};
test_weights[11416:11423] = '{32'h4290d7bb, 32'h4295b540, 32'hc2a4d7bc, 32'hc2199e12, 32'hc1cf7f93, 32'h427dc65a, 32'hc14be597, 32'hc1e7494c};
test_bias[1427:1427] = '{32'h42b9bb8a};
test_output[1427:1427] = '{32'hc5a9e371};
test_input[11424:11431] = '{32'hc24de9f7, 32'hc1c3eef6, 32'hc2a6fd8b, 32'h417ae2b9, 32'hc2c5b5e3, 32'h42925552, 32'h42be0fb6, 32'h429e54d1};
test_weights[11424:11431] = '{32'hc2a21923, 32'hc2b6da6d, 32'hc281908e, 32'hc25b8ec1, 32'h42ab1719, 32'hc2c2b834, 32'h411d1837, 32'hc2b882d4};
test_bias[1428:1428] = '{32'hc2abf87e};
test_output[1428:1428] = '{32'hc62d12ae};
test_input[11432:11439] = '{32'hc2ad1d49, 32'h42502d21, 32'h422c6df0, 32'hc2a9033a, 32'hc175018b, 32'h42708068, 32'hc1fd3706, 32'hc1536dec};
test_weights[11432:11439] = '{32'h42ab0d80, 32'h4160507e, 32'h42b10b0b, 32'h42a06308, 32'hc269bb22, 32'h42a390a4, 32'hc092ffde, 32'hc25c5805};
test_bias[1429:1429] = '{32'h412453ea};
test_output[1429:1429] = '{32'hc537aa0b};
test_input[11440:11447] = '{32'hc21b05eb, 32'h42073172, 32'hc2bc1f31, 32'hc0e23b91, 32'hc206d132, 32'h42b0ef38, 32'hc2a8de77, 32'h42961ab1};
test_weights[11440:11447] = '{32'hc229375c, 32'hc2885bb7, 32'hc1bb2581, 32'h41242645, 32'h422108da, 32'h42a05c2a, 32'hc22222d3, 32'hc28f431f};
test_bias[1430:1430] = '{32'h429c871f};
test_output[1430:1430] = '{32'h45a66113};
test_input[11448:11455] = '{32'h429f7e8c, 32'hc27c7ae1, 32'hc27196ac, 32'hc243e47b, 32'h41b09e59, 32'hc1a59618, 32'h42aee53e, 32'h426e8d2d};
test_weights[11448:11455] = '{32'h4254425f, 32'h422b3d68, 32'hc10987a7, 32'hc277741c, 32'hc281f8e9, 32'h427cdfad, 32'hc251eada, 32'h4249ec46};
test_bias[1431:1431] = '{32'hc291cf35};
test_output[1431:1431] = '{32'h442ae7d7};
test_input[11456:11463] = '{32'hc276b838, 32'h42ae3ada, 32'h3f5c1a4c, 32'h426063bc, 32'hc19380e2, 32'h410d7423, 32'h419b3d87, 32'h42afcb23};
test_weights[11456:11463] = '{32'hc203a320, 32'hc2bbdc6f, 32'hc2b02410, 32'h41e044fd, 32'hc2849575, 32'h410aa29a, 32'hc01e47f7, 32'hc2b3c68e};
test_bias[1432:1432] = '{32'hc23c08d6};
test_output[1432:1432] = '{32'hc63163e4};
test_input[11464:11471] = '{32'h42a45a2b, 32'h42b63b56, 32'hc2ae99f8, 32'hc288a3c2, 32'h41aade12, 32'h42451e4f, 32'hc2957520, 32'h42311ae7};
test_weights[11464:11471] = '{32'h42c10486, 32'h3f94fa06, 32'h42144312, 32'hc0d772c3, 32'h42484cbf, 32'hc2b25cd1, 32'hc1ba769a, 32'h4288eddd};
test_bias[1433:1433] = '{32'h4241c1b0};
test_output[1433:1433] = '{32'h45d32969};
test_input[11472:11479] = '{32'hc2c37290, 32'hc044a1d3, 32'h40d17b17, 32'hc2a2fb8d, 32'h40f7ec90, 32'h42c0978b, 32'h420910f5, 32'h411b4e10};
test_weights[11472:11479] = '{32'h41bdcd2c, 32'hc2c7de45, 32'hc0b7b4be, 32'h4295bb74, 32'h4013c476, 32'hc277622e, 32'h42066e1a, 32'hc2b7a12c};
test_bias[1434:1434] = '{32'hc287e9e0};
test_output[1434:1434] = '{32'hc6591cab};
test_input[11480:11487] = '{32'h42b92de5, 32'hc1e8219f, 32'hc2a61610, 32'hc1f3e24d, 32'hc2c625a9, 32'hc2c18dc8, 32'hc24c778e, 32'hc29bfef8};
test_weights[11480:11487] = '{32'hc1ff5065, 32'hc2868792, 32'hc2a31d6e, 32'hc26d1d10, 32'hc10217b5, 32'h41a2e73b, 32'h404ea1cc, 32'h4110fed8};
test_bias[1435:1435] = '{32'h41df45aa};
test_output[1435:1435] = '{32'h45adfd8d};
test_input[11488:11495] = '{32'h4229643d, 32'h40dbca93, 32'hc15793fd, 32'h42c669ba, 32'h42844382, 32'hc282ad2d, 32'hc22df899, 32'hc1c8b439};
test_weights[11488:11495] = '{32'h409bc15a, 32'h42c69531, 32'hc12a46c5, 32'h4221f33f, 32'h4095d82a, 32'hc2bea90f, 32'hc2b35f5e, 32'h4292fe66};
test_bias[1436:1436] = '{32'hc241dbbe};
test_output[1436:1436] = '{32'h46546b65};
test_input[11496:11503] = '{32'h4240a3f1, 32'hc245f514, 32'h41a748a3, 32'h423f5be6, 32'hc261aad6, 32'h40078bcc, 32'h417645ea, 32'h426dc733};
test_weights[11496:11503] = '{32'hc2a9498c, 32'h42b18cba, 32'hc1f5a31d, 32'hc2b0f910, 32'h42728164, 32'hc1b734c4, 32'hc23cf2b2, 32'hc1446099};
test_bias[1437:1437] = '{32'h426887f4};
test_output[1437:1437] = '{32'hc68e48ec};
test_input[11504:11511] = '{32'hc11ee276, 32'h3f447a05, 32'h42924dfc, 32'h41e3449c, 32'hc22f95a0, 32'hc283b9f6, 32'hc02b2da1, 32'h42bb274c};
test_weights[11504:11511] = '{32'h42707f0e, 32'h415bc32e, 32'hc230e2f9, 32'h422fcf0e, 32'hc1d82d6f, 32'h41e40919, 32'h418c8013, 32'hc2b6cce4};
test_bias[1438:1438] = '{32'hc243f492};
test_output[1438:1438] = '{32'hc63a23b5};
test_input[11512:11519] = '{32'hc2b35d6c, 32'h4140215b, 32'h42a4fcd0, 32'hc20135d5, 32'h41dd9d08, 32'hc20f7518, 32'h420f1dd8, 32'hc258f693};
test_weights[11512:11519] = '{32'h4269fc2e, 32'h41b653f8, 32'h4247fad0, 32'hc21bfb05, 32'hc22a9376, 32'h424e6a75, 32'h42c47f0c, 32'hc29c4467};
test_bias[1439:1439] = '{32'hc1c0e1dc};
test_output[1439:1439] = '{32'h459fa4d1};
test_input[11520:11527] = '{32'hc291c39c, 32'hc276006e, 32'hc2ab6f37, 32'h4131a914, 32'h42b3c5cb, 32'h42b41cd8, 32'hc1976a52, 32'hc10580bd};
test_weights[11520:11527] = '{32'hc1aad90b, 32'h42030096, 32'h41ea367e, 32'hc284bf62, 32'h42735a83, 32'h4283b6e3, 32'hc1dedf74, 32'hc1b48c91};
test_bias[1440:1440] = '{32'h42aa6acd};
test_output[1440:1440] = '{32'h4604bff4};
test_input[11528:11535] = '{32'h42486280, 32'h42343718, 32'hbff2059f, 32'hc2432bd4, 32'hc2b59488, 32'h429b0469, 32'hc27716b5, 32'hc1895eff};
test_weights[11528:11535] = '{32'hc28f205b, 32'hc1bad05c, 32'h408409b0, 32'h4188e5c3, 32'hc21f91ab, 32'hc151579d, 32'h42a0fe67, 32'h424487b9};
test_bias[1441:1441] = '{32'h421c84ed};
test_output[1441:1441] = '{32'hc60724be};
test_input[11536:11543] = '{32'h421187c8, 32'h4291ab7d, 32'hc2827cab, 32'h429b652d, 32'hc2214815, 32'hc26494b9, 32'h3fa4b009, 32'hc2a089d7};
test_weights[11536:11543] = '{32'h4289a721, 32'h424321dd, 32'hc29a5edf, 32'h41c298e7, 32'h41af0b02, 32'h42a2a250, 32'h41c535dc, 32'hc28c5676};
test_bias[1442:1442] = '{32'hc0b8deb4};
test_output[1442:1442] = '{32'h464ce0f2};
test_input[11544:11551] = '{32'hc283ffa2, 32'hc21218b0, 32'h41f139e4, 32'h420d7944, 32'hc28d5741, 32'h42b55ccb, 32'h42993f1c, 32'h42985b86};
test_weights[11544:11551] = '{32'h418ea3cd, 32'h419fa48e, 32'h4297cb9c, 32'hc283243e, 32'h421c313d, 32'h41d752a8, 32'h42110ef0, 32'h42a401d1};
test_bias[1443:1443] = '{32'hc1b03e1e};
test_output[1443:1443] = '{32'h45d2e4bf};
test_input[11552:11559] = '{32'hc0c1d941, 32'h41c6e93d, 32'h41ec336d, 32'hc1f8f61f, 32'hc2ac2108, 32'hc2b71c92, 32'hc28832bb, 32'h42132de4};
test_weights[11552:11559] = '{32'hc1ef0564, 32'hc29b8e44, 32'hc1065721, 32'h41834d36, 32'h42ba7c4f, 32'h4086bbc1, 32'hc2be09bc, 32'hc2a1f1c4};
test_bias[1444:1444] = '{32'hc20a4352};
test_output[1444:1444] = '{32'hc5e94912};
test_input[11560:11567] = '{32'h4244b316, 32'h4284219c, 32'h42824754, 32'hc29fd85b, 32'h42b9c2c1, 32'h3e12b663, 32'h4223abcc, 32'hc2bf4ef1};
test_weights[11560:11567] = '{32'h429129e4, 32'h40e9a668, 32'h40f7623b, 32'hc2ae90b2, 32'hc09fe969, 32'h420f6ff1, 32'h4141cb65, 32'h4296b822};
test_bias[1445:1445] = '{32'hc2158af6};
test_output[1445:1445] = '{32'h45870e0b};
test_input[11568:11575] = '{32'h416d330d, 32'h429ea297, 32'h428a8484, 32'hc1b876c3, 32'hc2474c17, 32'hc1920cad, 32'h42c14d00, 32'hc292b66d};
test_weights[11568:11575] = '{32'h42a4bdea, 32'h41b97467, 32'hc21edf31, 32'hc25a5943, 32'hc28b34ce, 32'h425d992f, 32'hc2a35391, 32'hc2c12881};
test_bias[1446:1446] = '{32'hc200c5d8};
test_output[1446:1446] = '{32'h4546ffa5};
test_input[11576:11583] = '{32'hc29bcefe, 32'hc1eb67b0, 32'h4281b1d6, 32'hc24aa401, 32'h42a5029a, 32'h3f25946f, 32'h4241f428, 32'h4012f71f};
test_weights[11576:11583] = '{32'h42303f6b, 32'hc29d175e, 32'h41ed00b3, 32'hc2c411c1, 32'h421c184a, 32'h4251efd2, 32'hc28d9dac, 32'h41b6373a};
test_bias[1447:1447] = '{32'hc1fbad1a};
test_output[1447:1447] = '{32'h45af3a61};
test_input[11584:11591] = '{32'h42a8de3c, 32'hc29c9553, 32'h42a4b7d6, 32'hc2a0cbeb, 32'hc180fb01, 32'hc29dc828, 32'hc18a2227, 32'hc194b47b};
test_weights[11584:11591] = '{32'hc2bdc2cd, 32'hc19e6133, 32'h42bf48c2, 32'hc2a3b129, 32'h42bedcd7, 32'hc190f434, 32'hc2ad91c9, 32'hc28bbe1e};
test_bias[1448:1448] = '{32'h427e26e9};
test_output[1448:1448] = '{32'h4627ef01};
test_input[11592:11599] = '{32'hc2b3a0d1, 32'hc24428ca, 32'hc24d85f3, 32'hc225b915, 32'hc2c6d61f, 32'h427b0f89, 32'h42b26149, 32'hc1b52173};
test_weights[11592:11599] = '{32'hc1854140, 32'h42843b93, 32'hc1a86320, 32'h42765f78, 32'hc2a714ef, 32'hc210928d, 32'hc21cba19, 32'h42b53849};
test_bias[1449:1449] = '{32'hc2a8c820};
test_output[1449:1449] = '{32'hc52fa449};
test_input[11600:11607] = '{32'hc21d8ee4, 32'h41f50d76, 32'h427be450, 32'hc27d20a7, 32'h42ad43db, 32'hc21a5a14, 32'hc27a94a1, 32'hc16685c2};
test_weights[11600:11607] = '{32'hc285577c, 32'hc2261351, 32'hc2007170, 32'h423ac906, 32'hc19e39b1, 32'h3eac4d00, 32'h42271999, 32'hc28aef9e};
test_bias[1450:1450] = '{32'h427723ce};
test_output[1450:1450] = '{32'hc5d7bc77};
test_input[11608:11615] = '{32'hc2bc9185, 32'h4214fd47, 32'h42210932, 32'hc23057d6, 32'h424ba5da, 32'hc101ff21, 32'hc28abb54, 32'h424304fd};
test_weights[11608:11615] = '{32'h41b88dd6, 32'hc27a2001, 32'h42a2a79d, 32'h42a222a6, 32'hc18de1a5, 32'h425a87ca, 32'h4293958a, 32'h425fd458};
test_bias[1451:1451] = '{32'h42766222};
test_output[1451:1451] = '{32'hc6047e8b};
test_input[11616:11623] = '{32'h422d3376, 32'hc2af3a59, 32'hc0088ec9, 32'hc217ab56, 32'hc130ce71, 32'hc1a60cba, 32'hc29b7e93, 32'hc2272b6f};
test_weights[11616:11623] = '{32'h40ae9685, 32'h41a83e29, 32'hc2c67544, 32'hc24bec68, 32'hc2065118, 32'hc277cec1, 32'hc2b36a2c, 32'h4269bc2c};
test_bias[1452:1452] = '{32'h42adcff9};
test_output[1452:1452] = '{32'h45d4f5e9};
test_input[11624:11631] = '{32'hc28dda82, 32'h426fad43, 32'h4246178b, 32'h41d23c3d, 32'hc281750b, 32'hc0284711, 32'hc2024f05, 32'hc294011d};
test_weights[11624:11631] = '{32'h42ab8ae1, 32'hc2b67005, 32'h42c23af7, 32'hc26fd37d, 32'hc2c6a32b, 32'h41fd77c6, 32'hc2ad63b7, 32'hc11e74cf};
test_bias[1453:1453] = '{32'hc248f4c0};
test_output[1453:1453] = '{32'h44c01e26};
test_input[11632:11639] = '{32'hc25f8c1e, 32'h3fef1a84, 32'h42c70074, 32'hc0a6e6e5, 32'hc0b8ddfc, 32'h42a9723c, 32'h429cc0db, 32'h429106b8};
test_weights[11632:11639] = '{32'h428fc5c7, 32'hc2773f18, 32'hc28108c3, 32'h410472a4, 32'h40ffc545, 32'hc25e1d44, 32'h413c4d8f, 32'hc1b6d8bc};
test_bias[1454:1454] = '{32'h421f6a57};
test_output[1454:1454] = '{32'hc67aa5d6};
test_input[11640:11647] = '{32'hc0db2b7c, 32'hc24b6083, 32'hc27e7142, 32'hc1dbc514, 32'h42c79443, 32'hc1e021e0, 32'h42940511, 32'h41b7b38d};
test_weights[11640:11647] = '{32'hc29eccee, 32'hc1b7061d, 32'hc1b155c5, 32'hc239d4cb, 32'hc1b7a6f0, 32'hc2802d06, 32'h421f8671, 32'hc26229f3};
test_bias[1455:1455] = '{32'h42049e9f};
test_output[1455:1455] = '{32'h45ae83bd};
test_input[11648:11655] = '{32'hc25899c7, 32'hc181544a, 32'hc28b290d, 32'h42528ef6, 32'h421edbbb, 32'hc203117b, 32'hc137fdff, 32'hc29c7bf9};
test_weights[11648:11655] = '{32'hc1571a57, 32'h42345fc5, 32'hc2966cc5, 32'hc28aa281, 32'h419bdc85, 32'hc24a70ad, 32'h4267fbc3, 32'h422c0ea8};
test_bias[1456:1456] = '{32'hc157f867};
test_output[1456:1456] = '{32'hc1f34507};
test_input[11656:11663] = '{32'hc1f84342, 32'hc0b16899, 32'h4273fd8c, 32'h4180cdbb, 32'h42990f4a, 32'hc2c493f0, 32'hc29623df, 32'h4159bf56};
test_weights[11656:11663] = '{32'h42ba0800, 32'h429fb4c2, 32'h411ec87a, 32'hc292caed, 32'h41b2759c, 32'h4257945b, 32'hc2b6b24f, 32'hc23d3233};
test_bias[1457:1457] = '{32'hc256e940};
test_output[1457:1457] = '{32'hc4a6f3d9};
test_input[11664:11671] = '{32'hc1902781, 32'h42c520fb, 32'h41d2b347, 32'hc1df06e3, 32'h4228e2b4, 32'h4291f7fd, 32'h41abe009, 32'h418c337a};
test_weights[11664:11671] = '{32'h429ef7a9, 32'h4189ed52, 32'hc2a337db, 32'hc1321b3f, 32'h42066c4d, 32'hc2af5c5b, 32'h416dd938, 32'h42c22eec};
test_bias[1458:1458] = '{32'h41c8f40f};
test_output[1458:1458] = '{32'hc58cd29d};
test_input[11672:11679] = '{32'hc2c23dde, 32'hc28a548b, 32'hc20e5777, 32'hc2c7a3e3, 32'h40585cfa, 32'h41a5ed34, 32'h429140e5, 32'hc2ad9828};
test_weights[11672:11679] = '{32'h4294e91b, 32'h42307845, 32'h40f35d68, 32'h42549a2e, 32'hc2b424c7, 32'h4235e169, 32'h41ac1b79, 32'hc297c6ac};
test_bias[1459:1459] = '{32'hc2500814};
test_output[1459:1459] = '{32'hc5de9643};
test_input[11680:11687] = '{32'h427699b4, 32'h42842bc4, 32'h4272be43, 32'hc22035d5, 32'hc23a668d, 32'hc2b7f3cb, 32'h40184497, 32'hc0bd4cdd};
test_weights[11680:11687] = '{32'hc295531a, 32'hc298ad5c, 32'hbf50985f, 32'h4170b1ee, 32'h42b9e138, 32'hc1de0ea2, 32'h411aae08, 32'h41cb1ce4};
test_bias[1460:1460] = '{32'hc262e98b};
test_output[1460:1460] = '{32'hc63f96e6};
test_input[11688:11695] = '{32'hc108a2fa, 32'hc2abc802, 32'hc2a890b4, 32'hc1b2fde4, 32'h40335051, 32'hc299427f, 32'hc210e702, 32'h42810c36};
test_weights[11688:11695] = '{32'h42c69c6b, 32'h422e3759, 32'hc2c02cf9, 32'h42b710e1, 32'h42862a26, 32'hc2b40e49, 32'h40a29873, 32'hc19507de};
test_bias[1461:1461] = '{32'hc23364f2};
test_output[1461:1461] = '{32'h45de6c07};
test_input[11696:11703] = '{32'h41807e60, 32'h429cf3c7, 32'h429d1876, 32'h41de122b, 32'hc2c1d6e9, 32'h4265b4ea, 32'h42b05549, 32'hc289338b};
test_weights[11696:11703] = '{32'hc2265e1c, 32'hc267495d, 32'hc2b05dc1, 32'h423d3c00, 32'h415861f7, 32'hc2904844, 32'hc1c3df36, 32'h4217a54d};
test_bias[1462:1462] = '{32'hc0befb84};
test_output[1462:1462] = '{32'hc6a45bea};
test_input[11704:11711] = '{32'h41e94f5b, 32'hc26434e7, 32'h427b019d, 32'h42884144, 32'h4181a85a, 32'hc24c9e00, 32'hc25b7920, 32'hc183a19b};
test_weights[11704:11711] = '{32'hc19149e8, 32'hc1382d17, 32'h42212470, 32'h42270886, 32'hc2c7781c, 32'h420d0292, 32'h42875421, 32'h425e8f77};
test_bias[1463:1463] = '{32'hc20c20e6};
test_output[1463:1463] = '{32'hc5216f0c};
test_input[11712:11719] = '{32'h426c152a, 32'h42686cae, 32'h404ae538, 32'h418c96fb, 32'h4082ab4a, 32'h42ae003b, 32'hc2c16345, 32'h4297dc64};
test_weights[11712:11719] = '{32'hc2b4c94b, 32'hc28bb33d, 32'hc21a2cd0, 32'h41369f9f, 32'h42b3b3c2, 32'hc2c7dd8c, 32'hc2beb3f0, 32'h42806896};
test_bias[1464:1464] = '{32'hc2ba07e2};
test_output[1464:1464] = '{32'hc5638bc4};
test_input[11720:11727] = '{32'h41ab33aa, 32'h423463a8, 32'h421abdc3, 32'hc2a55ea9, 32'hc08c83bc, 32'hc206ca4c, 32'hc22510d5, 32'h42a0fdaf};
test_weights[11720:11727] = '{32'hc234a44e, 32'hc1d5a7e0, 32'h42429681, 32'h41851fe4, 32'h4276c572, 32'h428b6808, 32'hc2251943, 32'hc2ac0a0e};
test_bias[1465:1465] = '{32'hc2b6f3ee};
test_output[1465:1465] = '{32'hc615f3f8};
test_input[11728:11735] = '{32'hc20502b9, 32'h42acb0c1, 32'hc190c15e, 32'h425aa55e, 32'hc2665ba1, 32'hc28309ca, 32'hc2216cc2, 32'h41be332e};
test_weights[11728:11735] = '{32'h428b9554, 32'hc2b07eca, 32'h4286c294, 32'h42bb1925, 32'hc2355cca, 32'hc2692b75, 32'hc1c0f3b5, 32'h417aa792};
test_bias[1466:1466] = '{32'h3f81e559};
test_output[1466:1466] = '{32'h44d8617b};
test_input[11736:11743] = '{32'h4286d38c, 32'h4212c87d, 32'hc0fe5dd4, 32'h41498b9d, 32'h4216c895, 32'h428c00f5, 32'h3f95847a, 32'h42c54739};
test_weights[11736:11743] = '{32'hc19fe1be, 32'h425f032a, 32'hc1a462b7, 32'hc2807cf4, 32'hc287cbcc, 32'hc28b5298, 32'hc1f135d1, 32'h41787b0b};
test_bias[1467:1467] = '{32'h41da3f0b};
test_output[1467:1467] = '{32'hc5b71a04};
test_input[11744:11751] = '{32'hc2316b37, 32'h41561a8d, 32'hc21cf2ea, 32'h4192c3eb, 32'hc24a7407, 32'hc1baf933, 32'hc2bec5f4, 32'hc1ea3715};
test_weights[11744:11751] = '{32'hc1139c79, 32'h429c166c, 32'h42356312, 32'hc22694be, 32'h42a54e2b, 32'h429d03be, 32'h416174a2, 32'h41073a4e};
test_bias[1468:1468] = '{32'h428d5093};
test_output[1468:1468] = '{32'hc606d32b};
test_input[11752:11759] = '{32'hc2bff3cd, 32'h4284803d, 32'hc2a2ce47, 32'hc229a3ed, 32'hc1ccbecf, 32'h42078f1e, 32'hc1eb9fb4, 32'hc245d96f};
test_weights[11752:11759] = '{32'hc1c12cdb, 32'hc16c1680, 32'hc219ca09, 32'hc21633a5, 32'hc2b76475, 32'h42548557, 32'hc2abdd7a, 32'h425cb73c};
test_bias[1469:1469] = '{32'h4298a99f};
test_output[1469:1469] = '{32'h461d9e62};
test_input[11760:11767] = '{32'h4239587b, 32'hc26a89bd, 32'hc051772f, 32'hc17a0fe1, 32'hc2ae7194, 32'hc299469d, 32'h4211cc2b, 32'hc2874f69};
test_weights[11760:11767] = '{32'h4200f9a3, 32'hbfae0adc, 32'hc2518f46, 32'hc20c5bff, 32'hc28286ad, 32'h427e5df2, 32'hc0a01249, 32'h4262f679};
test_bias[1470:1470] = '{32'hc21f456b};
test_output[1470:1470] = '{32'hc46d1ce5};
test_input[11768:11775] = '{32'h4291c46d, 32'h42335d76, 32'h40411601, 32'hc1d947d1, 32'h4297971f, 32'h3ffa996a, 32'hc22126ac, 32'h42b1a0a9};
test_weights[11768:11775] = '{32'hc02948fb, 32'h42a65aad, 32'hc2bce289, 32'hc2976dff, 32'hc2c333b5, 32'h41f3f9c7, 32'hc218508d, 32'h42c09400};
test_bias[1471:1471] = '{32'h3ffc64d5};
test_output[1471:1471] = '{32'h45fbd2f7};
test_input[11776:11783] = '{32'h42618c08, 32'hc1acca82, 32'hc0987128, 32'h42be790b, 32'hc28da225, 32'hc2467b7f, 32'hc1fd4d50, 32'h408926b4};
test_weights[11776:11783] = '{32'h3f558901, 32'h42b1dfc6, 32'hc27febcd, 32'h4284decc, 32'h420779d8, 32'hc1ae62d9, 32'h42280f64, 32'hc284d56f};
test_bias[1472:1472] = '{32'h425c21b0};
test_output[1472:1472] = '{32'h44eb248c};
test_input[11784:11791] = '{32'h42c52c72, 32'hc2c6f1ad, 32'h42974206, 32'hc2bacaa7, 32'h428c3cea, 32'h4230d43b, 32'hc25a5b4d, 32'hc243db77};
test_weights[11784:11791] = '{32'h42538f22, 32'h422bfd83, 32'h42553d8c, 32'h41b1c1f2, 32'hc1cfeab8, 32'h42855367, 32'hc1858ed1, 32'hc010936e};
test_bias[1473:1473] = '{32'hc2a07228};
test_output[1473:1473] = '{32'h459b00c8};
test_input[11792:11799] = '{32'hc01761ad, 32'hc2855c7a, 32'hc277eaa0, 32'hc03f194f, 32'hc1fe4383, 32'h427af355, 32'h425e139c, 32'hc278a19a};
test_weights[11792:11799] = '{32'hc2b081e1, 32'h4250c49d, 32'hc1ede6b3, 32'h42843dea, 32'hc1a95102, 32'h4296c365, 32'h425861e3, 32'hc201021e};
test_bias[1474:1474] = '{32'h41ad8b65};
test_output[1474:1474] = '{32'h460997b3};
test_input[11800:11807] = '{32'hc18c4af2, 32'h41b37af8, 32'hc2394069, 32'h4299f562, 32'h42c63e8a, 32'h40b5ad82, 32'h40dd271c, 32'h42844cd1};
test_weights[11800:11807] = '{32'h42a00c3e, 32'h42465612, 32'h42b987e9, 32'h429182c2, 32'h42a64dd6, 32'h42991acc, 32'h42803e98, 32'hc1778590};
test_bias[1475:1475] = '{32'h424a5341};
test_output[1475:1475] = '{32'h460f22d1};
test_input[11808:11815] = '{32'hc29e091e, 32'h4295db0a, 32'h420e7154, 32'hc2a7b952, 32'h42a2bf0e, 32'hc28c2b7f, 32'h41b7f837, 32'hc289f0af};
test_weights[11808:11815] = '{32'hc29ab5a8, 32'hc23dfe85, 32'hc2796ce2, 32'h41bcc03a, 32'hc28f839b, 32'h42a7170f, 32'hc268fef5, 32'h40196e5d};
test_bias[1476:1476] = '{32'h417de19f};
test_output[1476:1476] = '{32'hc667b443};
test_input[11816:11823] = '{32'hc1ef14d9, 32'h42b997aa, 32'h42993c9c, 32'hc28fb833, 32'hc21ea924, 32'h40d1a9cb, 32'hc299b492, 32'hc27c2845};
test_weights[11816:11823] = '{32'hc28fa775, 32'h426f4430, 32'h41b20dc7, 32'h42c20e1b, 32'hc2aa8174, 32'h42bccfc8, 32'hc26f80fc, 32'h4281d85d};
test_bias[1477:1477] = '{32'hc29d9e72};
test_output[1477:1477] = '{32'h45d663c7};
test_input[11824:11831] = '{32'hc2b50047, 32'h42be0aa8, 32'hc2b63e9f, 32'hc28893b8, 32'h4243adab, 32'hc2960091, 32'h42aa02e6, 32'hc2c6d999};
test_weights[11824:11831] = '{32'h420b8efc, 32'hc2b374b1, 32'hc19b7056, 32'hc096b9a3, 32'h425261e6, 32'h40c36949, 32'hc15b7541, 32'h42406502};
test_bias[1478:1478] = '{32'hc236685d};
test_output[1478:1478] = '{32'hc65278d8};
test_input[11832:11839] = '{32'hc20d42f9, 32'h42bcd644, 32'hc2c5f95c, 32'hc19343e2, 32'hc2828e4f, 32'h41c53038, 32'h4295f794, 32'h429760fa};
test_weights[11832:11839] = '{32'hc29e3421, 32'h400c67f7, 32'hc2303596, 32'hc10d6b37, 32'hc0d96a3c, 32'hc28b8f2e, 32'h41ea4ff8, 32'h40b297ef};
test_bias[1479:1479] = '{32'h42733f72};
test_output[1479:1479] = '{32'h460b7bc9};
test_input[11840:11847] = '{32'h429a8c93, 32'h428c2be4, 32'hc2b2e971, 32'hc0930b19, 32'hc0de874b, 32'hc0ed97e7, 32'h42a2f760, 32'h41493fbd};
test_weights[11840:11847] = '{32'hc27b3694, 32'hc2943cd7, 32'h3f9cba0a, 32'hc2c6b870, 32'hc29f8b06, 32'h42b48341, 32'hc2979d2c, 32'hc2643c08};
test_bias[1480:1480] = '{32'h42231c43};
test_output[1480:1480] = '{32'hc6823c11};
test_input[11848:11855] = '{32'hc20d5dd0, 32'hc28f8ff2, 32'h42a7fe23, 32'h428556da, 32'h428f6437, 32'h42a1b88f, 32'hc248ee67, 32'h41eb359c};
test_weights[11848:11855] = '{32'h412c34b7, 32'hc23f730a, 32'h42afa1eb, 32'h40da0137, 32'h418677df, 32'hc2bd21c4, 32'hc25e9f63, 32'h41929dce};
test_bias[1481:1481] = '{32'hc1b580c8};
test_output[1481:1481] = '{32'h45f2602a};
test_input[11856:11863] = '{32'h42be7e47, 32'h42a4de87, 32'hc284545f, 32'h421f78bf, 32'hc1178b8e, 32'h428088c5, 32'hc2b05af9, 32'hc2b78463};
test_weights[11856:11863] = '{32'h42bc6d72, 32'h4217ef51, 32'hc18dc5f0, 32'hc21cef63, 32'hc2952687, 32'h4293b527, 32'hc199bb95, 32'h421b2a61};
test_bias[1482:1482] = '{32'hc2aa76dd};
test_output[1482:1482] = '{32'h466dbe75};
test_input[11864:11871] = '{32'hc23e8fd5, 32'hc203396b, 32'h40f0c9d3, 32'h423914eb, 32'hc28f5398, 32'hc2216332, 32'h421cc73e, 32'h42b496a0};
test_weights[11864:11871] = '{32'h40cc2ddd, 32'hc2b96e34, 32'h417cb77a, 32'h413c062b, 32'hc2c57b9c, 32'hc092757d, 32'h42639ea0, 32'hc2b068ae};
test_bias[1483:1483] = '{32'hc1b98c0f};
test_output[1483:1483] = '{32'h45993ee3};
test_input[11872:11879] = '{32'hc2bf8aea, 32'h41cc436a, 32'h429d8c02, 32'hc24e532f, 32'hc249a900, 32'h42117fc5, 32'hc1a79fb3, 32'h42347e95};
test_weights[11872:11879] = '{32'hc1ce9f1a, 32'h3f7c0f05, 32'hc25cc2db, 32'hc29ee896, 32'hc2381e1e, 32'hc279a96f, 32'h3ed5a274, 32'hbfbb4e7c};
test_bias[1484:1484] = '{32'hc1a6aa98};
test_output[1484:1484] = '{32'h4509c217};
test_input[11880:11887] = '{32'hc234f884, 32'hc280581a, 32'h418048b2, 32'hc1df08c3, 32'h429b19e4, 32'hc2bf6363, 32'h42256487, 32'hc2b09f1b};
test_weights[11880:11887] = '{32'h41211277, 32'h40174ecf, 32'h42a1d841, 32'hc1ebe9db, 32'h41d77dcc, 32'h42090bd0, 32'h41a45d62, 32'hc2b506bf};
test_bias[1485:1485] = '{32'h428fa881};
test_output[1485:1485] = '{32'h4610562a};
test_input[11888:11895] = '{32'hc277bd1c, 32'hbfaa5bcf, 32'hc22f9db3, 32'h42bc0057, 32'hc261923e, 32'hc28401cd, 32'hc2441640, 32'h41882d2c};
test_weights[11888:11895] = '{32'h42180b44, 32'hc1a12dc3, 32'hc2ab8be0, 32'h4241fe41, 32'h428f8a32, 32'hc1d2eecc, 32'hc2818263, 32'h4265cd13};
test_bias[1486:1486] = '{32'h420fda61};
test_output[1486:1486] = '{32'h45f63434};
test_input[11896:11903] = '{32'hc2aedf74, 32'h4146fb67, 32'h4253569b, 32'hc1e73237, 32'hc218601c, 32'h422781ac, 32'h41d38ffa, 32'hc2bf13fc};
test_weights[11896:11903] = '{32'hc29ef4cf, 32'h4145fdbc, 32'hc1eef5e0, 32'hc28dc47a, 32'hc224eb06, 32'hc2c57094, 32'h4282c9c1, 32'hc151e5b0};
test_bias[1487:1487] = '{32'hc2413a77};
test_output[1487:1487] = '{32'h45f8438a};
test_input[11904:11911] = '{32'hc17c8b7b, 32'hc2c10ec2, 32'h412ac844, 32'hc09c5dee, 32'h415e5b3d, 32'hc22a0bf5, 32'h42948e24, 32'hc2b555a3};
test_weights[11904:11911] = '{32'hc2c3892b, 32'h42bfc8eb, 32'h4189f607, 32'hc2902fdc, 32'h425d8b66, 32'hc0dbbeab, 32'hc205e129, 32'h422cdbfc};
test_bias[1488:1488] = '{32'hc10a555d};
test_output[1488:1488] = '{32'hc643c05a};
test_input[11912:11919] = '{32'h4246efb9, 32'h423b410a, 32'h427f5816, 32'hc25f6dda, 32'hc2c0eab8, 32'hc24e65d9, 32'hc0b87d90, 32'hc256e784};
test_weights[11912:11919] = '{32'hc0b6a65f, 32'hc2a97359, 32'hc2b0ceb1, 32'hc0990263, 32'h41e1b96e, 32'hc27e539a, 32'h40f49d62, 32'h42a15aa4};
test_bias[1489:1489] = '{32'hc29dce06};
test_output[1489:1489] = '{32'hc65352ce};
test_input[11920:11927] = '{32'h42050682, 32'h420cc6f9, 32'h427fdb09, 32'h40d5ecb0, 32'h42bd3b4e, 32'hc1d21f80, 32'hc1042acf, 32'hc1b30ec2};
test_weights[11920:11927] = '{32'hc1a5a908, 32'hc2a07bdb, 32'h42501130, 32'hc1c27c9b, 32'hc2840315, 32'h40fc8d99, 32'hc1732589, 32'h418bc261};
test_bias[1490:1490] = '{32'hc0c4954a};
test_output[1490:1490] = '{32'hc5dd0168};
test_input[11928:11935] = '{32'h41b3ecca, 32'h4222209f, 32'h40443102, 32'hc14d691e, 32'h4245f0f7, 32'hc181f5a6, 32'h41389a35, 32'hc1e36f6f};
test_weights[11928:11935] = '{32'hc26a9b07, 32'hc2c71639, 32'h427b810e, 32'h42c22dae, 32'h426db41d, 32'hc1f4af38, 32'h4279a50d, 32'hc2a234c5};
test_bias[1491:1491] = '{32'h421c0776};
test_output[1491:1491] = '{32'h42bdc329};
test_input[11936:11943] = '{32'hc21f1157, 32'hc26a62a3, 32'hc2bf160f, 32'hc24161a3, 32'hc26fee8d, 32'hc2b4e861, 32'hc2c70d25, 32'h4084f8e6};
test_weights[11936:11943] = '{32'hc21762fa, 32'h42c25f0e, 32'hc202fb7b, 32'hc2b811f0, 32'h4207a421, 32'hc07114a4, 32'h42b3bb4b, 32'hc25583be};
test_bias[1492:1492] = '{32'h4286bdb2};
test_output[1492:1492] = '{32'hc5e75a65};
test_input[11944:11951] = '{32'h41e2f7e9, 32'hc20a9114, 32'hc1b591a7, 32'h42baf14b, 32'hc258f001, 32'hc189f42c, 32'h42ae6304, 32'hc24dd043};
test_weights[11944:11951] = '{32'h4220bdeb, 32'hc085d165, 32'hc2b0fb8a, 32'h41cacfc0, 32'h42ac98a5, 32'hc224715f, 32'h42bc63cf, 32'h41a2930d};
test_bias[1493:1493] = '{32'h42609ac2};
test_output[1493:1493] = '{32'h460b4d3a};
test_input[11952:11959] = '{32'h4276a4d2, 32'hc0e2277e, 32'h40d59627, 32'hc100769c, 32'h4273e0f0, 32'hc260cc70, 32'h42427884, 32'h42513af9};
test_weights[11952:11959] = '{32'hc2316084, 32'h41b6d6d2, 32'hc2b97112, 32'hc2566f62, 32'h41bc48df, 32'h42bb3729, 32'h406cc0c3, 32'h41d3bed5};
test_bias[1494:1494] = '{32'h4258fd62};
test_output[1494:1494] = '{32'hc5a55bb5};
test_input[11960:11967] = '{32'hc1d5568b, 32'h429015c2, 32'h427f1f19, 32'h40601ba2, 32'hc205c228, 32'h41fd0484, 32'hc280878d, 32'hc1a99087};
test_weights[11960:11967] = '{32'h426e4c7e, 32'h41dcde6d, 32'hc2a4a9d9, 32'h42b4e62c, 32'hc288eac4, 32'h426eb6d6, 32'h419256fa, 32'hc2527919};
test_bias[1495:1495] = '{32'hc1fc1881};
test_output[1495:1495] = '{32'hc3e09d8d};
test_input[11968:11975] = '{32'h41a77015, 32'hc22d141f, 32'h421bbcce, 32'h3faae472, 32'h4298c425, 32'h42c63966, 32'hc2a9db56, 32'hc2ae4d7f};
test_weights[11968:11975] = '{32'h42945198, 32'hc28731ac, 32'hc114cc05, 32'hc1cd988f, 32'h4193c0ca, 32'hc15103ef, 32'h428f71be, 32'h419e97db};
test_bias[1496:1496] = '{32'h42943e58};
test_output[1496:1496] = '{32'hc55dc342};
test_input[11976:11983] = '{32'hbf5e2269, 32'h42ac5ffe, 32'h42a30d2c, 32'h42803142, 32'h41e4ba6c, 32'hc262d071, 32'hc27c45b6, 32'hc1c7a446};
test_weights[11976:11983] = '{32'hc2b74de8, 32'h42a0ef63, 32'hc2094306, 32'h4241aad2, 32'hc28d2f5e, 32'hc29a3aee, 32'hc2b7e6cf, 32'h41c9bb35};
test_bias[1497:1497] = '{32'hc292adfb};
test_output[1497:1497] = '{32'h4666cdf9};
test_input[11984:11991] = '{32'hc1c3af35, 32'hc19d156e, 32'hc23836a7, 32'h425a9a8d, 32'hc19df030, 32'hbe740c06, 32'hc24481c1, 32'h4209cb5f};
test_weights[11984:11991] = '{32'h42634dc5, 32'h4284f672, 32'hc2a00d11, 32'hc25ad7a2, 32'h42c556ab, 32'hc2b43f07, 32'hc2766f84, 32'hc1f3154b};
test_bias[1498:1498] = '{32'h429b73b6};
test_output[1498:1498] = '{32'hc4e99896};
test_input[11992:11999] = '{32'h4299edf1, 32'hc2879de8, 32'h418f134d, 32'hc2a6f49e, 32'hc202302e, 32'h414f3fa6, 32'hc20acaf3, 32'h3f4cc910};
test_weights[11992:11999] = '{32'hc2851d39, 32'hc06b6aa8, 32'h42ad68a7, 32'h428c2e1b, 32'h42ba7c25, 32'h41fcceee, 32'h42b99739, 32'h41d538f7};
test_bias[1499:1499] = '{32'h422c0054};
test_output[1499:1499] = '{32'hc669a97d};
test_input[12000:12007] = '{32'h421a8a07, 32'h422969d0, 32'hc2a6b594, 32'h42b5c21e, 32'h42b2cc79, 32'h42c373e5, 32'hc2a639ee, 32'hc102d2a4};
test_weights[12000:12007] = '{32'h428de7c3, 32'hc17ce224, 32'h41dc8948, 32'hc2521023, 32'hc15bd74b, 32'h42ac1d13, 32'h415f60f6, 32'hc264c9ca};
test_bias[1500:1500] = '{32'h42313f20};
test_output[1500:1500] = '{32'h44bfd64b};
test_input[12008:12015] = '{32'hc1ca7cd5, 32'hc1a80f1f, 32'hc28ba5e8, 32'hc22e62ca, 32'hc2866b57, 32'hbf99bcef, 32'h429b1ab8, 32'hc2079d54};
test_weights[12008:12015] = '{32'h42663519, 32'h42809075, 32'hc16b2406, 32'h41c33fa1, 32'h41c03cfe, 32'hc29bfbca, 32'hc28f01be, 32'h4204319e};
test_bias[1501:1501] = '{32'hc1f5c2a3};
test_output[1501:1501] = '{32'hc62cdaf9};
test_input[12016:12023] = '{32'h40eae12e, 32'hc18e98ef, 32'hc2b9256f, 32'h42aeb8ab, 32'h4099b23b, 32'h4299ce99, 32'h42b4f599, 32'hc2c04033};
test_weights[12016:12023] = '{32'h42aa671a, 32'hc2c32327, 32'hc1b737b9, 32'hc20e87f8, 32'hc297ab84, 32'hc208caf6, 32'hc2c240e9, 32'hc278df2b};
test_bias[1502:1502] = '{32'h402d510d};
test_output[1502:1502] = '{32'hc58a5849};
test_input[12024:12031] = '{32'h42bb04ba, 32'hc203bac5, 32'hc1e77ae0, 32'h4138a1d2, 32'h4294636f, 32'h4272eda0, 32'hc2512bb9, 32'h42b57676};
test_weights[12024:12031] = '{32'hc2c129bd, 32'h41d116e5, 32'h4220bae7, 32'hc2961a57, 32'hc2956f85, 32'hc294354a, 32'h42aa65a3, 32'hc2bec3d1};
test_bias[1503:1503] = '{32'hc2251818};
test_output[1503:1503] = '{32'hc7092b91};
test_input[12032:12039] = '{32'h4299c171, 32'h42982d9c, 32'h42934ccd, 32'hc284f9a7, 32'hc037c8e6, 32'h423e210f, 32'h42c01867, 32'h4266f5bf};
test_weights[12032:12039] = '{32'h4190d996, 32'h4205241e, 32'h429379b5, 32'h42a59979, 32'hc1cf88d4, 32'hc2c54040, 32'hc21146b5, 32'h420a9905};
test_bias[1504:1504] = '{32'h419a60ca};
test_output[1504:1504] = '{32'hc50b7907};
test_input[12040:12047] = '{32'h40820173, 32'h4116ee9c, 32'hc1f44136, 32'h4294c891, 32'hc18edf52, 32'h41cb71e0, 32'h4177ec8e, 32'hc12eabcb};
test_weights[12040:12047] = '{32'hc24c1b03, 32'hbef3d46f, 32'hc2951206, 32'h41b4e905, 32'hc1470e10, 32'hc28b79a0, 32'h42676e39, 32'h41b4d1fd};
test_bias[1505:1505] = '{32'hc2346a83};
test_output[1505:1505] = '{32'h452ef8ef};
test_input[12048:12055] = '{32'h42c14539, 32'h42b94a52, 32'hc28dc817, 32'hc16e970a, 32'hc16066ca, 32'h410bc795, 32'h429ba2b6, 32'h41ffebfe};
test_weights[12048:12055] = '{32'hc2839332, 32'h425a849e, 32'h41378ebc, 32'h428b6714, 32'h42b59709, 32'h410301ca, 32'h429b0d8b, 32'h42aea1f5};
test_bias[1506:1506] = '{32'h42a6015f};
test_output[1506:1506] = '{32'h458e738b};
test_input[12056:12063] = '{32'h42854c66, 32'hc26637f8, 32'hc10be1c2, 32'h42afef7d, 32'hc244c247, 32'hbf598224, 32'h429e751c, 32'hc1c8ab29};
test_weights[12056:12063] = '{32'hc1385a4a, 32'h4277c684, 32'hc24c9df6, 32'h416a6f67, 32'hc22da51a, 32'h41b79d66, 32'h429a423a, 32'hc292cc73};
test_bias[1507:1507] = '{32'hc220510f};
test_output[1507:1507] = '{32'h45e836ad};
test_input[12064:12071] = '{32'h42a5a03d, 32'hc2a78b0b, 32'hc2c4df1a, 32'hc285d7a6, 32'hc20e8882, 32'h42c4c741, 32'h40aa37a7, 32'hc2667ee8};
test_weights[12064:12071] = '{32'hc22b3e5e, 32'hc298f53b, 32'h4293256d, 32'h41e3b6d2, 32'h4204fa3a, 32'h4288f34e, 32'hc24990b8, 32'hc28aa1c1};
test_bias[1508:1508] = '{32'hc2877aaf};
test_output[1508:1508] = '{32'h4536d760};
test_input[12072:12079] = '{32'h3fa325e2, 32'h42194398, 32'hc1c44501, 32'hc2a6a848, 32'hc29505ab, 32'h409149d0, 32'hc1cdad64, 32'hc13b93e8};
test_weights[12072:12079] = '{32'hc2111fb6, 32'hc2b6aafb, 32'h41972e67, 32'h428bb511, 32'hc247e1b6, 32'hc21860d1, 32'hc268767a, 32'hc2242450};
test_bias[1509:1509] = '{32'h427163ec};
test_output[1509:1509] = '{32'hc584a23e};
test_input[12080:12087] = '{32'hc2a37a3d, 32'hc28e5755, 32'hc217815a, 32'hc29e4774, 32'hc20f5b5b, 32'hc2bbc427, 32'h41005a30, 32'hc2a6c71f};
test_weights[12080:12087] = '{32'hc215c962, 32'h4259065b, 32'hc29a746a, 32'hc23368e5, 32'h42a02f3f, 32'hc27e9a15, 32'hc2c3aee3, 32'h41aff284};
test_bias[1510:1510] = '{32'hc24842a3};
test_output[1510:1510] = '{32'h45bef31d};
test_input[12088:12095] = '{32'h41cc10c8, 32'hc2ac1919, 32'h42abba23, 32'h42410516, 32'h413e67d9, 32'hc1727f29, 32'h42b3b85c, 32'h41fa923e};
test_weights[12088:12095] = '{32'hc209d633, 32'hc2a6dfcd, 32'h4188668b, 32'h429128df, 32'h4190f6d5, 32'hc28ccfb3, 32'hc27f728e, 32'hc1b376a3};
test_bias[1511:1511] = '{32'h429bbee1};
test_output[1511:1511] = '{32'h45c152a0};
test_input[12096:12103] = '{32'hc23348a9, 32'hc25c9e1a, 32'hc29171ba, 32'h429814b5, 32'h421fb844, 32'h41a06eb1, 32'h420a64e9, 32'h42094a4a};
test_weights[12096:12103] = '{32'hc2186a8e, 32'h423c133d, 32'h4297db95, 32'h42c16dcb, 32'hc08330b4, 32'h41bf93ca, 32'hc29cc124, 32'hc2a8bfb0};
test_bias[1512:1512] = '{32'h42bf9b0d};
test_output[1512:1512] = '{32'hc584c233};
test_input[12104:12111] = '{32'h4269175f, 32'hc2a0375e, 32'h418118b6, 32'h42b83a20, 32'h420ee002, 32'hc14b71df, 32'hc2889b69, 32'hc2be03ce};
test_weights[12104:12111] = '{32'hc1b7b44e, 32'hc1e73fee, 32'hc1a6561e, 32'hc0ca6a3f, 32'h4293d7c2, 32'hc293b6a1, 32'hc1260003, 32'hc28abef3};
test_bias[1513:1513] = '{32'hc2bf2862};
test_output[1513:1513] = '{32'h46296b4d};
test_input[12112:12119] = '{32'h42b0baf7, 32'hc227343c, 32'h4211a2a9, 32'hc078e6cc, 32'h42b2ce58, 32'hc20defbe, 32'h4242218a, 32'hc223d24f};
test_weights[12112:12119] = '{32'hc2a11665, 32'hc209762c, 32'hc28bf134, 32'h41ee5d39, 32'hc131424e, 32'hc2a1484c, 32'hc2b0089b, 32'hc21e6e98};
test_bias[1514:1514] = '{32'hc278cd12};
test_output[1514:1514] = '{32'hc60f83ae};
test_input[12120:12127] = '{32'h41d11252, 32'hc1c67e73, 32'h4223113b, 32'h4104ffff, 32'hc1958b6b, 32'hc2bc3a35, 32'hc235b97b, 32'h42a2497d};
test_weights[12120:12127] = '{32'h40a2ec1a, 32'hc20acd91, 32'hc2127385, 32'h409a663e, 32'h41d56d58, 32'h42bd78eb, 32'h428444b7, 32'hc26fbed0};
test_bias[1515:1515] = '{32'hc2bfc29b};
test_output[1515:1515] = '{32'hc68b59fa};
test_input[12128:12135] = '{32'hc2b97068, 32'hc22a7f79, 32'hc2b249a6, 32'h42715815, 32'h40dee542, 32'h427ba5fc, 32'hc2b354f2, 32'h40ece9dd};
test_weights[12128:12135] = '{32'h4291bdff, 32'hc289c384, 32'hc1e9cbcf, 32'hc23fe437, 32'hc0877ca4, 32'h426929eb, 32'h41d6b190, 32'hc227f9ec};
test_bias[1516:1516] = '{32'h426517fa};
test_output[1516:1516] = '{32'hc543c14d};
test_input[12136:12143] = '{32'h422e4971, 32'hc2a3ecc2, 32'hc20f6243, 32'hc2b9a03c, 32'h40f9a5aa, 32'h423f862d, 32'hc2b35e05, 32'hc29bd9d8};
test_weights[12136:12143] = '{32'hc286f4e1, 32'hc2a22ef9, 32'h41081afd, 32'h428574c7, 32'h428f9e16, 32'h42b6af3e, 32'h42543ceb, 32'hc13300dd};
test_bias[1517:1517] = '{32'h41aae503};
test_output[1517:1517] = '{32'hc4d76e53};
test_input[12144:12151] = '{32'hc2c680c0, 32'h429a8d54, 32'h416634f6, 32'hc1b2c770, 32'h42896704, 32'h4228d7a9, 32'hc2bb359c, 32'hc2139aa4};
test_weights[12144:12151] = '{32'h41b98dbd, 32'hc2952e12, 32'hc2c63162, 32'hc26eb34c, 32'h4229fd1d, 32'hc0eb9427, 32'hc296750b, 32'hc2a1c9b1};
test_bias[1518:1518] = '{32'hc262a5c0};
test_output[1518:1518] = '{32'h458a25d6};
test_input[12152:12159] = '{32'hc216ed78, 32'hc2b6f906, 32'hc2ac7191, 32'h404f2ac9, 32'hc1b9ce0e, 32'h417114a4, 32'h413ef2d2, 32'hc242aecd};
test_weights[12152:12159] = '{32'hc2908cf1, 32'h41cd912b, 32'h416a0ac4, 32'hc2a44d4b, 32'h42c09804, 32'h42835003, 32'h40f8e81e, 32'h420be6d6};
test_bias[1519:1519] = '{32'hc2663dc2};
test_output[1519:1519] = '{32'hc57e12ae};
test_input[12160:12167] = '{32'h42a9ecba, 32'h428e5920, 32'h42a4d21f, 32'hc265c9ff, 32'hc1b2560d, 32'h42542838, 32'h417a71b6, 32'h42a50199};
test_weights[12160:12167] = '{32'h42b1d09e, 32'hc2878ba6, 32'h42036ff3, 32'hc1469cbf, 32'h4282c6f5, 32'h4211ad6d, 32'h42ab2cb1, 32'h4280292e};
test_bias[1520:1520] = '{32'hc0d1469d};
test_output[1520:1520] = '{32'h464ef4ac};
test_input[12168:12175] = '{32'h42b9b7b3, 32'h41811e45, 32'h4274a7de, 32'hc22ab2c8, 32'h42ba6e20, 32'hc2a25d70, 32'h40a17dbf, 32'h420adc51};
test_weights[12168:12175] = '{32'hc2499f36, 32'hc23a14ae, 32'hc2a7c673, 32'hc2c1b2dc, 32'h4251f945, 32'hc2742b3d, 32'hc240dfa7, 32'hc1b6efde};
test_bias[1521:1521] = '{32'h422527c8};
test_output[1521:1521] = '{32'h451778bf};
test_input[12176:12183] = '{32'h42099e0c, 32'hc2bfb188, 32'h42120349, 32'hc19a4f88, 32'h42810ac5, 32'hc1683b12, 32'h426bfb25, 32'hc1a7305f};
test_weights[12176:12183] = '{32'h42c6b451, 32'hc2881e32, 32'h427463de, 32'hc281ff65, 32'hc1b270c9, 32'h429db9fb, 32'hc186d5a5, 32'hc230abb3};
test_bias[1522:1522] = '{32'h41d52614};
test_output[1522:1522] = '{32'h4628b3c8};
test_input[12184:12191] = '{32'hc1cb98b9, 32'h428d4f9b, 32'h4279666f, 32'h42aba919, 32'hc29494fd, 32'h427f0f62, 32'h428b2793, 32'hc2202948};
test_weights[12184:12191] = '{32'hc2b0cd14, 32'h42983592, 32'hc204da83, 32'h42b1a60b, 32'hc29f5b3d, 32'h42926509, 32'h42a11994, 32'hc2159fa6};
test_bias[1523:1523] = '{32'hc288f0d3};
test_output[1523:1523] = '{32'h46f0a0e5};
test_input[12192:12199] = '{32'h4201f5ca, 32'hc06dbfb7, 32'h41d860a6, 32'hc2b60e4a, 32'hc28946c0, 32'hc2b3950b, 32'hc10daf43, 32'hc242fd33};
test_weights[12192:12199] = '{32'hc29a188f, 32'h429bc144, 32'hc228d020, 32'h421af3bf, 32'h429274a4, 32'h417eb6b9, 32'h41196cea, 32'hc1a781ca};
test_bias[1524:1524] = '{32'h3f88d37d};
test_output[1524:1524] = '{32'hc64acc89};
test_input[12200:12207] = '{32'h4219e191, 32'h42731bab, 32'hc23c9fd8, 32'h4296a93c, 32'hc20da352, 32'h424a4d40, 32'hc271cacf, 32'hc278b382};
test_weights[12200:12207] = '{32'hc244cdf1, 32'hc2c3420a, 32'hc22a51b8, 32'h42910cb4, 32'hc0b963c3, 32'h428dd9a4, 32'hc24d60d4, 32'h3f13ba5e};
test_bias[1525:1525] = '{32'h4298fe42};
test_output[1525:1525] = '{32'h45cdaada};
test_input[12208:12215] = '{32'h4281e64f, 32'hc1791ad9, 32'hc0314b36, 32'hc235a546, 32'h42638ff2, 32'h4162d727, 32'hc28425e9, 32'hc2c38dac};
test_weights[12208:12215] = '{32'hc22eaf3f, 32'h42c4f2d4, 32'hc25230e1, 32'hc2aea700, 32'hc29842d1, 32'h426de08c, 32'hc29f1e94, 32'hc23461a9};
test_bias[1526:1526] = '{32'h42a0fa17};
test_output[1526:1526] = '{32'h45bb81a6};
test_input[12216:12223] = '{32'hc1b0226a, 32'hc289f710, 32'hc20b4b5b, 32'hc26d9655, 32'hc04578bc, 32'hc03b7fd5, 32'hc297f5df, 32'hc2b67315};
test_weights[12216:12223] = '{32'hc1c963ce, 32'hc03976b5, 32'h426e0718, 32'hc2279142, 32'h421a4285, 32'h418345db, 32'hc1c18b06, 32'h428b5422};
test_bias[1527:1527] = '{32'hc2b42f7c};
test_output[1527:1527] = '{32'hc5613f1d};
test_input[12224:12231] = '{32'h4283ae2b, 32'hc1a1c211, 32'hc1b34e11, 32'hc2b48c8b, 32'hc2b796f0, 32'hc2a5d8ba, 32'hc1f9297d, 32'hc1ed58e8};
test_weights[12224:12231] = '{32'hc1eddde5, 32'hc1163b96, 32'hc0d91643, 32'h424d25e7, 32'hc28adaf5, 32'hc2a609df, 32'hc233adab, 32'h416acb3d};
test_bias[1528:1528] = '{32'h428a7049};
test_output[1528:1528] = '{32'h45fb6470};
test_input[12232:12239] = '{32'h422ba5b1, 32'h423b6d60, 32'h4289ed9b, 32'h41ea0e82, 32'h41f0d2a1, 32'h42453ab0, 32'hc2c6e378, 32'h40c05c90};
test_weights[12232:12239] = '{32'h4250c7a0, 32'h42abc45c, 32'hc0453c0d, 32'h422972b6, 32'hc296ad2a, 32'hc22771d0, 32'h42aecc9a, 32'h422b8b6f};
test_bias[1529:1529] = '{32'hc29e240e};
test_output[1529:1529] = '{32'hc5ad8e02};
test_input[12240:12247] = '{32'h42427add, 32'hc297ec9e, 32'h423ec56a, 32'h427ba675, 32'hc2b2ec69, 32'hc2bdf1e7, 32'h41cbc186, 32'hc1e7c688};
test_weights[12240:12247] = '{32'hc2b2bf36, 32'h41ba636a, 32'h4213314b, 32'hc2800b83, 32'hc201b35c, 32'h42b630b7, 32'h421c4746, 32'hc2bd03f7};
test_bias[1530:1530] = '{32'h3f39d972};
test_output[1530:1530] = '{32'hc622932d};
test_input[12248:12255] = '{32'h425f01a0, 32'h42b73044, 32'hc2802a8c, 32'hc26f6ea7, 32'h41f0a765, 32'h42b6ea3c, 32'h42546235, 32'h41e98be5};
test_weights[12248:12255] = '{32'h4290512b, 32'hc2a73d6b, 32'h4273766c, 32'hc2989d0f, 32'h41d69238, 32'h42228c9f, 32'hc112db31, 32'h423710e3};
test_bias[1531:1531] = '{32'h41314632};
test_output[1531:1531] = '{32'h4516e319};
test_input[12256:12263] = '{32'hc11555ee, 32'hc25ea12f, 32'h42bbf431, 32'hc2bcbe87, 32'h4280ceff, 32'h42a6be62, 32'hc229162d, 32'h41b24d87};
test_weights[12256:12263] = '{32'h4218db15, 32'hc0a577fb, 32'hc0cd93b0, 32'hc2a9b5c0, 32'h41f13747, 32'hc16b208a, 32'h4219c485, 32'h429d3119};
test_bias[1532:1532] = '{32'hc165e764};
test_output[1532:1532] = '{32'h45ff2377};
test_input[12264:12271] = '{32'h428a57ae, 32'h428780ad, 32'h4161bba3, 32'hc1a46444, 32'hc2a0cf54, 32'h42801697, 32'h429dbca2, 32'h42bf3a7c};
test_weights[12264:12271] = '{32'hc2b32acf, 32'hc208d3f9, 32'hc2bbfcdd, 32'h42431bf1, 32'hc2874f49, 32'hc2571220, 32'hc29ff9e0, 32'h42bd37ae};
test_bias[1533:1533] = '{32'h42c666a4};
test_output[1533:1533] = '{32'hc5bbcda2};
test_input[12272:12279] = '{32'h4293ca51, 32'hc21b9564, 32'hc1caad9d, 32'hc1cf163f, 32'hc2138280, 32'h42956fcf, 32'h4221cc0f, 32'hc2802db9};
test_weights[12272:12279] = '{32'hc19d486a, 32'hc29cdf43, 32'h41dc79fa, 32'h41de7849, 32'h4227f9bd, 32'h42416b3c, 32'hc29ca735, 32'h4256da68};
test_bias[1534:1534] = '{32'hc12bada0};
test_output[1534:1534] = '{32'hc588c8d5};
test_input[12280:12287] = '{32'hc29d400a, 32'hc2428126, 32'h41affd12, 32'h429fce98, 32'hc1cafdb5, 32'hc2c3b16c, 32'h418b252f, 32'hc1b6f2d9};
test_weights[12280:12287] = '{32'hc2393cd7, 32'hc21fcf01, 32'hc19a9de3, 32'h420c862f, 32'h4245f1fc, 32'hc08f139c, 32'h424442c9, 32'hc215aeae};
test_bias[1535:1535] = '{32'h42397dd5};
test_output[1535:1535] = '{32'h460b1c4f};
test_input[12288:12295] = '{32'h40225fc5, 32'hc09e0e64, 32'h40d04f68, 32'h421ea85b, 32'hc29cdcc6, 32'h42b498f4, 32'h421b9b08, 32'h426c62a4};
test_weights[12288:12295] = '{32'hc25a7126, 32'hc06560dd, 32'hc106d9c5, 32'hc2b4860e, 32'hbc558687, 32'hc1d31cd4, 32'h422a3107, 32'hc1d91fcd};
test_bias[1536:1536] = '{32'hc24f2bcf};
test_output[1536:1536] = '{32'hc5bfd268};
test_input[12296:12303] = '{32'hc21db84d, 32'h41873683, 32'hc22a514f, 32'hc2b5b5e9, 32'h41daefd9, 32'h42a34c9e, 32'hc2b3a5cc, 32'hc2c3f88c};
test_weights[12296:12303] = '{32'hc228a7b4, 32'hc29c8b41, 32'hc267a033, 32'h41c5468e, 32'h422ab2f7, 32'hc26d6582, 32'h3faa746e, 32'h41b65099};
test_bias[1537:1537] = '{32'hc1c21eaf};
test_output[1537:1537] = '{32'hc5ab90a8};
test_input[12304:12311] = '{32'h41c7e21e, 32'hc2a18fdf, 32'h416e3821, 32'h41bf749e, 32'h428bf437, 32'hc2b94622, 32'h42b946ca, 32'hc292f342};
test_weights[12304:12311] = '{32'hc24fc740, 32'h428eff73, 32'h42a42996, 32'h4299d186, 32'h426d43e0, 32'hc0562fab, 32'h42b3cd49, 32'h428e61fc};
test_bias[1538:1538] = '{32'h428f9ba5};
test_output[1538:1538] = '{32'h45623225};
test_input[12312:12319] = '{32'h4124548b, 32'hc2a21ccf, 32'hc190e48c, 32'hc296ef0d, 32'h41b5ac21, 32'hc1f938bf, 32'h4289344b, 32'hc20bd2df};
test_weights[12312:12319] = '{32'h425ed822, 32'hc2b45778, 32'hc2640ac4, 32'h422ab2ec, 32'hc282a62d, 32'h428e14c2, 32'h4200e59b, 32'h4282cb8a};
test_bias[1539:1539] = '{32'hbfe6848a};
test_output[1539:1539] = '{32'h44efec06};
test_input[12320:12327] = '{32'h429abad8, 32'h410fab0e, 32'hc2c39ff6, 32'hc2c05f81, 32'h42b65bbb, 32'hc1c908e7, 32'h425d4203, 32'hc1ff1dcd};
test_weights[12320:12327] = '{32'h4242f8c6, 32'h3fdddb06, 32'hc2b4d525, 32'hbfaf44e8, 32'hc2201193, 32'h42899e76, 32'h42ad266a, 32'hc258e9d3};
test_bias[1540:1540] = '{32'hc1c8ded6};
test_output[1540:1540] = '{32'h4658d52c};
test_input[12328:12335] = '{32'h41536636, 32'h421b6c30, 32'h421448e4, 32'h42894225, 32'h42b0ec5c, 32'hc2c46b08, 32'hc2b87284, 32'h4085ac0e};
test_weights[12328:12335] = '{32'h419c0baa, 32'h42984fe6, 32'h42916462, 32'h42c44f41, 32'hc2c64a66, 32'hc2bb4434, 32'h4293c140, 32'h42b1fba1};
test_bias[1541:1541] = '{32'h4287690b};
test_output[1541:1541] = '{32'h45d15a57};
test_input[12336:12343] = '{32'hc2741725, 32'h42b692e1, 32'h42a94b4a, 32'h41605c66, 32'h42820720, 32'h41abd839, 32'hc2387ae8, 32'hc212ee53};
test_weights[12336:12343] = '{32'hc24439c7, 32'hc2637f87, 32'h42120b9b, 32'h4237ae1b, 32'h40cfd6e8, 32'h419d77cc, 32'hc20558dd, 32'hc18f2715};
test_bias[1542:1542] = '{32'h429d991f};
test_output[1542:1542] = '{32'h45917681};
test_input[12344:12351] = '{32'hc1949886, 32'hc11320d8, 32'hc2256d10, 32'h428825bd, 32'h40a3f5c3, 32'hc21ffb47, 32'h41d544b6, 32'hc038b832};
test_weights[12344:12351] = '{32'h41af6970, 32'h42bb81a7, 32'hc27574ce, 32'hc15adc1d, 32'hc2279fc3, 32'h427c5cbd, 32'hc05a1894, 32'hc28324ad};
test_bias[1543:1543] = '{32'h418b74db};
test_output[1543:1543] = '{32'hc50ecf27};
test_input[12352:12359] = '{32'h429f6bd4, 32'h429e96cb, 32'h4209d9e3, 32'hc0bf1603, 32'hc190752b, 32'hc2970fbf, 32'hc2980f3c, 32'h42b75d4b};
test_weights[12352:12359] = '{32'hc1fbc9c4, 32'hc200278a, 32'hc2b7dff1, 32'hc2032af3, 32'hc2a5b7dc, 32'hc2b4951e, 32'hc16398a6, 32'hc2941deb};
test_bias[1544:1544] = '{32'h42b9beb3};
test_output[1544:1544] = '{32'hc5a64ad8};
test_input[12360:12367] = '{32'hc20246a1, 32'h42463f5d, 32'hc22f4955, 32'h3fff1685, 32'h428a95d3, 32'hc2c2d764, 32'hc2bd86dc, 32'hc1494061};
test_weights[12360:12367] = '{32'h428fad90, 32'hc19f5455, 32'hc238e00f, 32'hc231b67d, 32'hc1b9c77a, 32'hc218236a, 32'h41d401c6, 32'h41ca7597};
test_bias[1545:1545] = '{32'h42c31108};
test_output[1545:1545] = '{32'hc4fd3b30};
test_input[12368:12375] = '{32'hc114513e, 32'h424cd928, 32'h413d0f1d, 32'h41e9ffa2, 32'hc235b485, 32'hc131ac64, 32'hc17940c0, 32'hc2a0e215};
test_weights[12368:12375] = '{32'hc10bd44f, 32'h42724418, 32'h4213375a, 32'hc2997c51, 32'hc2ab33f0, 32'hc19110ef, 32'h4228dd5c, 32'hc24d70be};
test_bias[1546:1546] = '{32'h425a5631};
test_output[1546:1546] = '{32'h460c7d00};
test_input[12376:12383] = '{32'hc186c52f, 32'h41943f7a, 32'hc2aac08a, 32'hc28c596a, 32'hc19f0b26, 32'hc29dd831, 32'hc2b81eea, 32'hc26c17c0};
test_weights[12376:12383] = '{32'h422cb79f, 32'h4282b342, 32'hc29d3559, 32'hc2621f81, 32'h424f3116, 32'h42ae43b0, 32'h429a2a0f, 32'hc21757e2};
test_bias[1547:1547] = '{32'hc2993d78};
test_output[1547:1547] = '{32'hc4d2915c};
test_input[12384:12391] = '{32'hc2a1ce6d, 32'hc29addc5, 32'h415eec3f, 32'hc1844a08, 32'h422423f2, 32'hc11221ec, 32'h42634f3b, 32'h427255c5};
test_weights[12384:12391] = '{32'hc2a2e2f3, 32'h429bca85, 32'hc2aa3ede, 32'h423c4043, 32'hc2661d08, 32'h42c5cc70, 32'hc2af9b39, 32'hc2c28b93};
test_bias[1548:1548] = '{32'hc2811ad9};
test_output[1548:1548] = '{32'hc67408b5};
test_input[12392:12399] = '{32'hc236f7bc, 32'hc2b27a47, 32'hc2acb942, 32'h428c68e8, 32'h4272259e, 32'h42454f93, 32'h415e43f3, 32'hc1322b0b};
test_weights[12392:12399] = '{32'hc1499408, 32'h427d3faa, 32'hc206e215, 32'hc2520565, 32'h429b2147, 32'h42793f34, 32'hc24426a9, 32'h428fb5a7};
test_bias[1549:1549] = '{32'hc10e18ef};
test_output[1549:1549] = '{32'h43d7b7f4};
test_input[12400:12407] = '{32'h413a8f38, 32'h40e3b4b8, 32'h4276a493, 32'hc29e8105, 32'h428196b6, 32'hc2a7da39, 32'h421e12ad, 32'hc2a8fad5};
test_weights[12400:12407] = '{32'h42b9e16a, 32'hc002538a, 32'h424a7118, 32'hc2b643f7, 32'hc0c08f9a, 32'h42c79312, 32'hc182abbb, 32'h4165f93e};
test_bias[1550:1550] = '{32'hc22e468b};
test_output[1550:1550] = '{32'h443a0c57};
test_input[12408:12415] = '{32'h4275d6cc, 32'h419371c1, 32'hc242d982, 32'h420035e6, 32'h427a832e, 32'hc2bfc605, 32'h4220ea8d, 32'h4288c3de};
test_weights[12408:12415] = '{32'h3e059e72, 32'hc0f1d51c, 32'hc1ea557a, 32'h42c6285d, 32'h3fe1381d, 32'h42b29277, 32'h42461963, 32'hc1f7ee2d};
test_bias[1551:1551] = '{32'hc20b428e};
test_output[1551:1551] = '{32'hc5816c71};
test_input[12416:12423] = '{32'hc1eeb6f7, 32'hc29b7952, 32'hc28cef26, 32'h42c47e9d, 32'h41919996, 32'hc1862616, 32'hc2c01e19, 32'h4281a207};
test_weights[12416:12423] = '{32'hc2afff46, 32'h41f592c2, 32'hc1ffe74e, 32'hc2162195, 32'hc2863154, 32'hc29f97e5, 32'hc27021a5, 32'hc1f31595};
test_bias[1552:1552] = '{32'hc1c7ffcf};
test_output[1552:1552] = '{32'h45287482};
test_input[12424:12431] = '{32'h429a7750, 32'h41e0f60b, 32'hc165053f, 32'h42b27a05, 32'hc20f2286, 32'h42b39494, 32'hc28a5a66, 32'h4262802f};
test_weights[12424:12431] = '{32'hc08e5824, 32'hc1851c14, 32'hc2aed985, 32'h413eb0ff, 32'hc2a63539, 32'h421ac417, 32'hc2a4ab7a, 32'hc28848e3};
test_bias[1553:1553] = '{32'hc2262ade};
test_output[1553:1553] = '{32'h46184bb0};
test_input[12432:12439] = '{32'hc28791be, 32'hc230bb13, 32'hc2b6367e, 32'hc2af1018, 32'hc2ba5e3a, 32'hc1c0a362, 32'hc214ae4e, 32'h421127dc};
test_weights[12432:12439] = '{32'hc0f9e325, 32'hc288bf61, 32'h40329a14, 32'hc247fc0a, 32'h4299094d, 32'h41ca17eb, 32'h4291343c, 32'hc2a8d864};
test_bias[1554:1554] = '{32'h425b26e9};
test_output[1554:1554] = '{32'hc5b46e22};
test_input[12440:12447] = '{32'h426b3146, 32'hc1622449, 32'hc2be4866, 32'hc22984af, 32'hc29e03da, 32'hc284f355, 32'h42b59d8f, 32'h425a7221};
test_weights[12440:12447] = '{32'hc0b9e91e, 32'hc133c2f6, 32'hc26f5a76, 32'hc23f5713, 32'hc231e2c7, 32'h428aed76, 32'hc29816ac, 32'hc137ec59};
test_bias[1555:1555] = '{32'hc0b28b66};
test_output[1555:1555] = '{32'hc48a28c4};
test_input[12448:12455] = '{32'h429c3ebc, 32'hc17a36e2, 32'h429a0f2b, 32'h421de5fc, 32'h42babd31, 32'h42a7a478, 32'h41b0f00f, 32'h428d6efb};
test_weights[12448:12455] = '{32'h40432b66, 32'hc1420bb5, 32'h42994735, 32'hc22b30ca, 32'hc292f690, 32'hc08ac022, 32'hc2b88294, 32'h42a0fc21};
test_bias[1556:1556] = '{32'hc2630c32};
test_output[1556:1556] = '{32'h447d2346};
test_input[12456:12463] = '{32'h4116d420, 32'h426cd01b, 32'h420beead, 32'h41d02857, 32'h418c98b8, 32'hc1443c02, 32'hc139b050, 32'hc2b38338};
test_weights[12456:12463] = '{32'hc2ad15f5, 32'hc26efee3, 32'h41a70a16, 32'h42bb40ca, 32'hc291f310, 32'hc23a0989, 32'hc2a779bc, 32'hc1955f31};
test_bias[1557:1557] = '{32'hc25f35aa};
test_output[1557:1557] = '{32'h442d5023};
test_input[12464:12471] = '{32'hc24a0dac, 32'hc2be2318, 32'h42b907cf, 32'hc11f778b, 32'h4174dcec, 32'h42b8711b, 32'h4222b1f1, 32'h42782917};
test_weights[12464:12471] = '{32'hc2199083, 32'hc22f7905, 32'h411612b8, 32'hc1f534f9, 32'h4237c760, 32'h4248d686, 32'hc2bc8a3f, 32'h42c0e656};
test_bias[1558:1558] = '{32'hc1fdd773};
test_output[1558:1558] = '{32'h466638d2};
test_input[12472:12479] = '{32'hc2753fcb, 32'hc101d21c, 32'h42117ce6, 32'hc2b0bc28, 32'hc20afdfd, 32'h42c193d6, 32'h42be189f, 32'hc1d53f0e};
test_weights[12472:12479] = '{32'hc24d7233, 32'hc2763cfc, 32'h42c78ca8, 32'h426353f1, 32'hc1fa36a9, 32'h42a05732, 32'hc1d4a7cc, 32'h428ebce4};
test_bias[1559:1559] = '{32'hc259fb42};
test_output[1559:1559] = '{32'h45ced34e};
test_input[12480:12487] = '{32'h4219005b, 32'h425c1afc, 32'h42b0b4ca, 32'h401b3205, 32'h4262f404, 32'h4256e165, 32'h429d01b1, 32'h422bc465};
test_weights[12480:12487] = '{32'hc296060f, 32'hc13e28db, 32'h413baeeb, 32'h4204706d, 32'h42ab0a4a, 32'h41a53c40, 32'h4254acaa, 32'hc2aeadb2};
test_bias[1560:1560] = '{32'hc2898474};
test_output[1560:1560] = '{32'h45745f1f};
test_input[12488:12495] = '{32'hc1f4583c, 32'hc2ad69b2, 32'h42934659, 32'h4284ef8f, 32'hc290e7e9, 32'hc267edda, 32'hc2204122, 32'h4282759d};
test_weights[12488:12495] = '{32'hc29dfe64, 32'h42aa6631, 32'h429866cd, 32'hc254676f, 32'h427df448, 32'h4280e2e0, 32'h42b318f4, 32'h42a707e5};
test_bias[1561:1561] = '{32'hc185e74a};
test_output[1561:1561] = '{32'hc612a813};
test_input[12496:12503] = '{32'hc2909e60, 32'h4208aa5b, 32'hc284d30f, 32'hc252384e, 32'h41371572, 32'h42574f24, 32'h429a933c, 32'h42ba8214};
test_weights[12496:12503] = '{32'hc27c6416, 32'hc1206e84, 32'h42a85d8f, 32'h42aa5468, 32'h420d2199, 32'h41be7077, 32'hc25d3f04, 32'hc1ec4de3};
test_bias[1562:1562] = '{32'hc23357f9};
test_output[1562:1562] = '{32'hc62f8f43};
test_input[12504:12511] = '{32'hc20c72fd, 32'hc234b1e5, 32'h40800c85, 32'h417a7b8b, 32'h42443261, 32'h40740f3d, 32'h41b23fde, 32'hc2646519};
test_weights[12504:12511] = '{32'hc2a17f8d, 32'hc2be778a, 32'hc1c1463c, 32'h423caab1, 32'h411eeb63, 32'h41e4d4a2, 32'hc215745a, 32'h4243f639};
test_bias[1563:1563] = '{32'hc1889ada};
test_output[1563:1563] = '{32'h4593c39a};
test_input[12512:12519] = '{32'hc20900dc, 32'hc0e75f68, 32'hc281274a, 32'hc29f91c8, 32'hc25f733c, 32'h41baa790, 32'h426dc692, 32'hc276f761};
test_weights[12512:12519] = '{32'hc2c4e9cb, 32'h429dcc6f, 32'h40b8e79a, 32'hbfbcc9a2, 32'h4288240f, 32'h418924cf, 32'h42aa7e61, 32'h41a90a59};
test_bias[1564:1564] = '{32'hc25325e4};
test_output[1564:1564] = '{32'h45325b02};
test_input[12520:12527] = '{32'hc20322fd, 32'hc0d009af, 32'hc2a6f3b7, 32'hc2883358, 32'h413ef062, 32'hc0a01c74, 32'hc2b83ae3, 32'h41eaaffa};
test_weights[12520:12527] = '{32'h41edc0d1, 32'h41aff60a, 32'hc096a751, 32'h42abca77, 32'hc2bd1661, 32'hc20c5def, 32'h42225603, 32'hc2c52199};
test_bias[1565:1565] = '{32'hc2afba0c};
test_output[1565:1565] = '{32'hc65e910e};
test_input[12528:12535] = '{32'hc29c75b9, 32'hc1019160, 32'hc2a3fc85, 32'hc09b10a3, 32'hc0889c7d, 32'hc202e14c, 32'hc1e3cae5, 32'hc209a01b};
test_weights[12528:12535] = '{32'h429b4935, 32'hc1383d41, 32'hc21e6706, 32'h42ace95f, 32'h41e6e9ab, 32'hc2b0b016, 32'hc09e47c1, 32'h421a6633};
test_bias[1566:1566] = '{32'h40271a8f};
test_output[1566:1566] = '{32'hc4c43ead};
test_input[12536:12543] = '{32'hc1e5d997, 32'hc1501c68, 32'hc28c6438, 32'hc15bf5c5, 32'h408a0935, 32'hc27be77c, 32'h421c4341, 32'h414ba146};
test_weights[12536:12543] = '{32'h420d4355, 32'h429d3f56, 32'h42740395, 32'h42a3ccf6, 32'h42263ad1, 32'hc2a38cf7, 32'h42858211, 32'h424b79cd};
test_bias[1567:1567] = '{32'hc243412d};
test_output[1567:1567] = '{32'h44884344};
test_input[12544:12551] = '{32'hc1901edb, 32'hc2a5091c, 32'h42c2ba2d, 32'hc1a06ab0, 32'h4266a5b1, 32'h422098cf, 32'h411ee452, 32'h42b3ef86};
test_weights[12544:12551] = '{32'hbfcbdc80, 32'h42ae574d, 32'hbfbb9dbb, 32'hc0bf1067, 32'h4299bb03, 32'h41ca10cf, 32'h41af9127, 32'hc28e7813};
test_bias[1568:1568] = '{32'h42c38e99};
test_output[1568:1568] = '{32'hc5f4d1c4};
test_input[12552:12559] = '{32'hc2886806, 32'hc21d633d, 32'h42302aa9, 32'h41e84694, 32'hc19929a0, 32'hc2b96cb8, 32'h42c0ae29, 32'h41ce1776};
test_weights[12552:12559] = '{32'hc292fa8e, 32'h4160e22b, 32'h4251bdba, 32'hc244f6e6, 32'h40e10b53, 32'hc245be7d, 32'h426f114b, 32'h411e23d6};
test_bias[1569:1569] = '{32'h3f2b3498};
test_output[1569:1569] = '{32'h4676e303};
test_input[12560:12567] = '{32'h41b19687, 32'hc232d94d, 32'hc29fd8c8, 32'h410a33d1, 32'hc28de7da, 32'h425f9c55, 32'h421b60cf, 32'h41bcfe6a};
test_weights[12560:12567] = '{32'hc291bf95, 32'hc1fb124e, 32'hc2b0119c, 32'hc030485a, 32'hc2bab9fa, 32'h428e4d53, 32'hc2c266a3, 32'h429e4219};
test_bias[1570:1570] = '{32'h4287fef4};
test_output[1570:1570] = '{32'h46732559};
test_input[12568:12575] = '{32'h4255aea7, 32'h42959125, 32'hc22dec5e, 32'hc1290461, 32'h3f740e47, 32'h4263cbb6, 32'h420fcafe, 32'hc180aa8a};
test_weights[12568:12575] = '{32'hc16aac0d, 32'h4278f76a, 32'h42878d9a, 32'hc1e6cf09, 32'h40f65caa, 32'hc2beaab1, 32'h414076c3, 32'h41326036};
test_bias[1571:1571] = '{32'h42636948};
test_output[1571:1571] = '{32'hc572ae92};
test_input[12576:12583] = '{32'h421363c6, 32'hc2b80fd7, 32'hc24283cb, 32'h420301f4, 32'h428ea430, 32'hc2689b76, 32'h42251afb, 32'hc1516664};
test_weights[12576:12583] = '{32'hc256f4b1, 32'hc1cbcc90, 32'h42b60595, 32'hc198af18, 32'h4262d920, 32'h423e6aea, 32'h4294fc36, 32'h4290faa9};
test_bias[1572:1572] = '{32'hc2b43a44};
test_output[1572:1572] = '{32'hc4abc262};
test_input[12584:12591] = '{32'h408bfad0, 32'hc2902930, 32'h42478e7a, 32'h40a854dc, 32'h4277662c, 32'hc190b58c, 32'h40fbdf82, 32'hc232056e};
test_weights[12584:12591] = '{32'h40a341e4, 32'h41faca9a, 32'hc1122cd2, 32'hc1fc3e49, 32'hc1d11328, 32'h420117fe, 32'hc24141b8, 32'hc1f05bf7};
test_bias[1573:1573] = '{32'h4279ffe1};
test_output[1573:1573] = '{32'hc57c7c8e};
test_input[12592:12599] = '{32'hc2404244, 32'h42c2a1c0, 32'h4225cec7, 32'hc2c3ffb0, 32'h42421d0b, 32'h42a20b3e, 32'h428d9617, 32'h41927e6b};
test_weights[12592:12599] = '{32'hc1d90131, 32'hc2a89bdc, 32'h40eba19d, 32'h4287f75e, 32'hc2bfc0eb, 32'h41a08342, 32'h42a0bad2, 32'h42c55072};
test_bias[1574:1574] = '{32'h42614283};
test_output[1574:1574] = '{32'hc608718b};
test_input[12600:12607] = '{32'hc1e51d26, 32'hc255fa22, 32'hbea6e56b, 32'h41c9642b, 32'hc13cf518, 32'h427878ae, 32'h419ec4b8, 32'h42a8ff8e};
test_weights[12600:12607] = '{32'h4136e69a, 32'hc2b42795, 32'hc242967b, 32'h42083617, 32'h42357215, 32'hc29ab9ff, 32'h41ccc467, 32'h40e663b6};
test_bias[1575:1575] = '{32'h41ed22f1};
test_output[1575:1575] = '{32'h44921f10};
test_input[12608:12615] = '{32'h4264a709, 32'h4263c66d, 32'h42767bb3, 32'h426404c9, 32'hc1513f43, 32'h4221c291, 32'h3fae3dbc, 32'h428503d9};
test_weights[12608:12615] = '{32'hc14b28d7, 32'h42aefb34, 32'hc2679c63, 32'hc1c884aa, 32'h4128f03b, 32'hc294f375, 32'h4201d9ee, 32'h42bef62e};
test_bias[1576:1576] = '{32'hc1d5eeae};
test_output[1576:1576] = '{32'h451ad29e};
test_input[12616:12623] = '{32'hc2ae2e59, 32'h42a58a0e, 32'hc1e8d112, 32'h41aab6d0, 32'hc1157358, 32'h42aa72d3, 32'h42bf9314, 32'h415ebaf0};
test_weights[12616:12623] = '{32'h42513c88, 32'h41cd800d, 32'hc28ee9fa, 32'hc12cd3c6, 32'h4272b4e7, 32'h418bddd4, 32'hc15d2b2a, 32'h4257cced};
test_bias[1577:1577] = '{32'hc2a43b5f};
test_output[1577:1577] = '{32'hc39c2dc8};
test_input[12624:12631] = '{32'h4299b881, 32'hc26e7c4b, 32'hc2c42ac7, 32'h41dc0754, 32'hc1c86ea5, 32'h427844fd, 32'h428a9483, 32'h40302f2e};
test_weights[12624:12631] = '{32'h41cf1aab, 32'hc27b2bce, 32'h421355f9, 32'h42337813, 32'hc2836f01, 32'hc0fa134d, 32'h4198eac6, 32'h42596264};
test_bias[1578:1578] = '{32'hc29173a6};
test_output[1578:1578] = '{32'h45b8ec27};
test_input[12632:12639] = '{32'h42b5889c, 32'hc228fc7d, 32'hc2833215, 32'hc2c2a2b7, 32'h42876094, 32'hc29496cf, 32'h42370676, 32'hc2118b40};
test_weights[12632:12639] = '{32'h41b7856b, 32'hc1b37b30, 32'h42907955, 32'h42933346, 32'h4254fc52, 32'hc1a0318d, 32'hc27eb66a, 32'hc28a7372};
test_bias[1579:1579] = '{32'hc26cd76f};
test_output[1579:1579] = '{32'hc5844aeb};
test_input[12640:12647] = '{32'hc28bff3c, 32'hc03bd153, 32'h42a054d5, 32'h4151a2af, 32'h41f615ec, 32'h428e911f, 32'h42bdd209, 32'hc16fbaab};
test_weights[12640:12647] = '{32'h421a4348, 32'h424c773c, 32'hc25062d0, 32'h424fd8cb, 32'hc2a6da19, 32'h41d29855, 32'hc2485009, 32'h40cc4b38};
test_bias[1580:1580] = '{32'h4224ef32};
test_output[1580:1580] = '{32'hc63908c0};
test_input[12648:12655] = '{32'hc2aaa8ab, 32'h40a3b348, 32'hc2c10884, 32'hc271de2c, 32'hc1a4f962, 32'hc147f9b0, 32'h4292ad3f, 32'hc1873f1f};
test_weights[12648:12655] = '{32'h42588960, 32'hc2c3d36f, 32'hc28ac56f, 32'hc29aeda9, 32'hc176a8e1, 32'h4293d88e, 32'hc23af6fb, 32'hc2c71f9d};
test_bias[1581:1581] = '{32'h4280cb9e};
test_output[1581:1581] = '{32'h4578666c};
test_input[12656:12663] = '{32'h41abd294, 32'hc2846a45, 32'h421d5bd3, 32'h41c20ed6, 32'hc2a023b2, 32'h4283c51b, 32'hc2b9495e, 32'h42bf6da5};
test_weights[12656:12663] = '{32'hc1a9df62, 32'hc21e1bba, 32'hc228ed30, 32'hc1f9b7da, 32'h42a6b8dc, 32'hc143a735, 32'hc155d5f8, 32'h4281ff25};
test_bias[1582:1582] = '{32'hc296d4e1};
test_output[1582:1582] = '{32'hc3b0ff3f};
test_input[12664:12671] = '{32'h429f6394, 32'h41bbe2d1, 32'hc214b54d, 32'hc23f728d, 32'h427e05f4, 32'h40edacb4, 32'h4271f585, 32'h426c5f46};
test_weights[12664:12671] = '{32'hc23f987f, 32'hc2a7ae74, 32'h41c844e2, 32'h427d08a2, 32'h42b43c63, 32'h4116fb0a, 32'h41eb6790, 32'h42518829};
test_bias[1583:1583] = '{32'h42a94b6b};
test_output[1583:1583] = '{32'h447c1e76};
test_input[12672:12679] = '{32'hc2471d63, 32'hc19efaae, 32'hc2b7b2c7, 32'h42a9bdad, 32'h41fb5d65, 32'hc1e62aef, 32'hc21c59d4, 32'h42560451};
test_weights[12672:12679] = '{32'hc2931925, 32'h414f8571, 32'hc2830614, 32'h42b952dc, 32'h4257237f, 32'h4201c808, 32'h42a66ea4, 32'h3ff26a0b};
test_bias[1584:1584] = '{32'h4245587d};
test_output[1584:1584] = '{32'h46696d30};
test_input[12680:12687] = '{32'hc25af1a2, 32'h41d61275, 32'h42a41a20, 32'h4253bcf0, 32'h428e753d, 32'h41e8fb8c, 32'h42182427, 32'h41a348fb};
test_weights[12680:12687] = '{32'h41a002af, 32'h428cae33, 32'hc0af40df, 32'hc2af5514, 32'h42251a30, 32'h426af785, 32'hc297d812, 32'hc2baa2ba};
test_bias[1585:1585] = '{32'hc270f18e};
test_output[1585:1585] = '{32'hc58cc300};
test_input[12688:12695] = '{32'h429fc3c9, 32'h42c06499, 32'hc1c232f8, 32'h42b778be, 32'hc2c653d3, 32'hc2425993, 32'h426714bb, 32'h426a155f};
test_weights[12688:12695] = '{32'h42c6ff35, 32'hc0b78a92, 32'h41d95d6b, 32'h420a80eb, 32'h42863589, 32'h40367cc7, 32'h419e737c, 32'h42086b80};
test_bias[1586:1586] = '{32'hc1c25db0};
test_output[1586:1586] = '{32'h45c2e18e};
test_input[12696:12703] = '{32'hc0832022, 32'h40ae7a3d, 32'h423fb83c, 32'h42c36240, 32'hc2b406c4, 32'hc2b6b57a, 32'hc2939a6c, 32'h428c0ca2};
test_weights[12696:12703] = '{32'h42572174, 32'hc280fdfe, 32'h419b1f5f, 32'hc29bccc9, 32'h42b7d65c, 32'hc2041b9c, 32'h4224821a, 32'hc2ad43cf};
test_bias[1587:1587] = '{32'hc2302e2f};
test_output[1587:1587] = '{32'hc6a92e97};
test_input[12704:12711] = '{32'hc2431086, 32'hc28828c0, 32'hc261cd18, 32'h415df308, 32'h41373b12, 32'hc0a732c3, 32'h422ac9a7, 32'hc2c62fb9};
test_weights[12704:12711] = '{32'hc16e4edb, 32'hc26d2fc2, 32'hc2c40a87, 32'hc2a47c52, 32'h40a528f5, 32'h4282bde5, 32'h42afd01a, 32'hc286cc29};
test_bias[1588:1588] = '{32'h42c34f22};
test_output[1588:1588] = '{32'h469795e7};
test_input[12712:12719] = '{32'h427f7ac2, 32'hc2064eff, 32'h42365f0d, 32'h42ba46f0, 32'h40dcf1dd, 32'h422fd709, 32'h4285fcd4, 32'hc0c790aa};
test_weights[12712:12719] = '{32'h42c399cf, 32'h429be6f4, 32'h427d9ca3, 32'h42808293, 32'h41ca958f, 32'h42b079eb, 32'h4235a8fb, 32'h42b76d5a};
test_bias[1589:1589] = '{32'hc275cb79};
test_output[1589:1589] = '{32'h46942ebd};
test_input[12720:12727] = '{32'h42b004c0, 32'h41d034d0, 32'h42874203, 32'h40946553, 32'hc083ef7b, 32'hc2122850, 32'h42892b54, 32'h421c825d};
test_weights[12720:12727] = '{32'hc0382937, 32'h428da723, 32'hc29f0442, 32'h421899da, 32'h40f9e37e, 32'h41d457ad, 32'hc1f75d22, 32'hc26779f8};
test_bias[1590:1590] = '{32'h4269a2c5};
test_output[1590:1590] = '{32'hc60baaa0};
test_input[12728:12735] = '{32'h4229fa47, 32'hc264553e, 32'hc23eade3, 32'hc2522d03, 32'h4269681a, 32'hc218dc10, 32'hc2843431, 32'h42155123};
test_weights[12728:12735] = '{32'hc2b4c68e, 32'h41ffb6a8, 32'hc24f4b68, 32'h42a656e0, 32'h41c42316, 32'hc2b845da, 32'hc2a9b72d, 32'hc1b8a087};
test_bias[1591:1591] = '{32'h428eb5b5};
test_output[1591:1591] = '{32'h4509d7b8};
test_input[12736:12743] = '{32'h41348611, 32'h42399683, 32'hc2a21c80, 32'h420340ad, 32'hc21f6224, 32'hc2106080, 32'hc0e67235, 32'hc2bc2e96};
test_weights[12736:12743] = '{32'hc014c234, 32'h429d8f59, 32'hc2899034, 32'hc29b9884, 32'h40b151e6, 32'hc2035cc1, 32'hc1e49262, 32'h42369a7b};
test_bias[1592:1592] = '{32'h420177af};
test_output[1592:1592] = '{32'h455e69fe};
test_input[12744:12751] = '{32'h4220f25f, 32'hc282eff9, 32'hc1c36971, 32'hc041adc4, 32'h4166e563, 32'hc27ab413, 32'h4224d724, 32'h42bbf4af};
test_weights[12744:12751] = '{32'hc293b051, 32'hc2036f53, 32'hc29b8f4c, 32'hc1c901e3, 32'hc2bc3f8b, 32'h42aa5826, 32'hc186a2d6, 32'hc1eb677d};
test_bias[1593:1593] = '{32'h4295a4e6};
test_output[1593:1593] = '{32'hc60b72e8};
test_input[12752:12759] = '{32'h425586d8, 32'h4249d8a0, 32'hc2969114, 32'h42a45d63, 32'h415f41cf, 32'hc2be4ae6, 32'h42842833, 32'h41dd3284};
test_weights[12752:12759] = '{32'hc1832eb3, 32'hc26e38ce, 32'h424de8ff, 32'h427d6b51, 32'h429a578a, 32'hc03900c4, 32'hc278eb11, 32'h409a7c5f};
test_bias[1594:1594] = '{32'hc18d5006};
test_output[1594:1594] = '{32'hc5a24dce};
test_input[12760:12767] = '{32'hc085cb44, 32'hc2c0ccd2, 32'hc104681f, 32'h4264e3bc, 32'hc1f41f00, 32'h4209de91, 32'hc20e3194, 32'hc092654f};
test_weights[12760:12767] = '{32'h42086210, 32'hc2778165, 32'hc27d04c5, 32'hc2af396b, 32'h40105952, 32'h42a06881, 32'h42417dcf, 32'h40f77eb8};
test_bias[1595:1595] = '{32'hc2ba7619};
test_output[1595:1595] = '{32'h45083d08};
test_input[12768:12775] = '{32'hc211f475, 32'h4268a8a3, 32'h42b8084e, 32'h424c4c10, 32'h41dd43a7, 32'hc29426fd, 32'hc25a8630, 32'hc12e7e47};
test_weights[12768:12775] = '{32'h41ab14e1, 32'hc228b00d, 32'h4225357b, 32'h420fa9d7, 32'h428aadf7, 32'hc2c337ba, 32'h42c71e8c, 32'hc28a9b26};
test_bias[1596:1596] = '{32'h423662f0};
test_output[1596:1596] = '{32'h45d80215};
test_input[12776:12783] = '{32'h428a3bb7, 32'h4041d020, 32'h41dc72dd, 32'hc2a7765a, 32'hc2389bda, 32'h415259a7, 32'hc27d091d, 32'hc02ed15d};
test_weights[12776:12783] = '{32'h41db24fa, 32'hc2abc54b, 32'h41862436, 32'hc1d2c15a, 32'h4239df1b, 32'h41a813ff, 32'h4292b448, 32'h428058f1};
test_bias[1597:1597] = '{32'h426ac169};
test_output[1597:1597] = '{32'hc5114086};
test_input[12784:12791] = '{32'h402cf67c, 32'h4295e6da, 32'h4292821f, 32'h42be8dd5, 32'h425fb35f, 32'hc14b9bc4, 32'h416455b7, 32'hc0e0ab11};
test_weights[12784:12791] = '{32'hc25df26b, 32'h42995153, 32'hc2973e71, 32'h423c7261, 32'h42b6cbde, 32'hc12999ce, 32'hc24af4ed, 32'hc1a842c1};
test_bias[1598:1598] = '{32'hc24cc954};
test_output[1598:1598] = '{32'h460f2dd5};
test_input[12792:12799] = '{32'h4231b5cd, 32'hc2a5cce7, 32'hc22f0c35, 32'hc2631b73, 32'hc27e6a05, 32'hc2163bdf, 32'h42b768d0, 32'hc2a1a6ae};
test_weights[12792:12799] = '{32'hc2c7a2d5, 32'h41edd526, 32'hc2abf55c, 32'hc2a33aec, 32'h42b5ec23, 32'hc2b666b2, 32'hc25750a3, 32'hc1e796f7};
test_bias[1599:1599] = '{32'hc29b902b};
test_output[1599:1599] = '{32'hc55d1312};
test_input[12800:12807] = '{32'h4237277f, 32'hc2b0874f, 32'hc1b92566, 32'hc2bf96ec, 32'hc2939950, 32'h4195c31f, 32'hc1797d91, 32'hc22795db};
test_weights[12800:12807] = '{32'hc24b956e, 32'h421a53bc, 32'hc2b38b82, 32'hc21079a8, 32'h428a2581, 32'hc29ea587, 32'h41de4ddc, 32'hc2b1b0ee};
test_bias[1600:1600] = '{32'hc1b68507};
test_output[1600:1600] = '{32'hc55ba8eb};
test_input[12808:12815] = '{32'hc29aaf7b, 32'hc2c008b8, 32'hc158b2e1, 32'hc19c56e5, 32'hc2a8c558, 32'h42b93e62, 32'h41963612, 32'h413c8d59};
test_weights[12808:12815] = '{32'h405ba66c, 32'hc2bfe91e, 32'hc2bbaad7, 32'hc290bad9, 32'hc1987639, 32'h42b57c83, 32'h42c7692f, 32'hc23d90f7};
test_bias[1601:1601] = '{32'hc27fd4c8};
test_output[1601:1601] = '{32'h46b2df33};
test_input[12816:12823] = '{32'h41d6a0f0, 32'hc29a88a5, 32'hc2aea535, 32'h41eb8a0d, 32'h42430f91, 32'hc14da08c, 32'hc27b443d, 32'hc2b06e19};
test_weights[12816:12823] = '{32'h422529d1, 32'h42aa20ba, 32'hc28808c7, 32'h429b031d, 32'hc19e1ec9, 32'hc1d99bfc, 32'h41a79503, 32'hc25fa472};
test_bias[1602:1602] = '{32'hc2c08182};
test_output[1602:1602] = '{32'h45b0f297};
test_input[12824:12831] = '{32'h42148060, 32'h4228686a, 32'h42544a4d, 32'h425cca61, 32'h426aa680, 32'hc26ef1f5, 32'h4143582c, 32'h42885395};
test_weights[12824:12831] = '{32'h429528bb, 32'h424db127, 32'hc2ba0175, 32'h408b2c3e, 32'hc2c0d0e2, 32'hc2b77061, 32'h414f328a, 32'hc2bab4b1};
test_bias[1603:1603] = '{32'hc217e9f9};
test_output[1603:1603] = '{32'hc5c12da3};
test_input[12832:12839] = '{32'h41d67152, 32'h4260b629, 32'h4198331b, 32'h428afb61, 32'h428256c0, 32'hc2266bde, 32'h4211c4e9, 32'hc1d3ca75};
test_weights[12832:12839] = '{32'hc24ef7b0, 32'h429c450f, 32'hc2a3d58a, 32'h416e9e00, 32'h42b65bd7, 32'h402f7685, 32'h4290ded4, 32'h4197c95e};
test_bias[1604:1604] = '{32'hc1c31b26};
test_output[1604:1604] = '{32'h4622d5ca};
test_input[12840:12847] = '{32'h40490869, 32'hc23f4174, 32'hc1152003, 32'h423ba2d4, 32'hc1593908, 32'h4225f44f, 32'h429d5d16, 32'hc27f245f};
test_weights[12840:12847] = '{32'h42ac97be, 32'h428822e1, 32'hc28ca74f, 32'hc204ea0b, 32'hc0f8c746, 32'hc2a568a7, 32'hc1443974, 32'hc12050fe};
test_bias[1605:1605] = '{32'hc2c16650};
test_output[1605:1605] = '{32'hc5ee9887};
test_input[12848:12855] = '{32'h4147aa2e, 32'h429fa1da, 32'h413fcb15, 32'hc25649b4, 32'h4105205a, 32'h420df8d7, 32'h4280f54b, 32'hc23c95d2};
test_weights[12848:12855] = '{32'h417b3c76, 32'hc1f4f6f5, 32'hc05997dc, 32'h42978066, 32'h421856ab, 32'hc2a57d57, 32'hc25dde89, 32'h41a54e4c};
test_bias[1606:1606] = '{32'hc291b263};
test_output[1606:1606] = '{32'hc65459cb};
test_input[12856:12863] = '{32'h42b05026, 32'hc1b8d0d3, 32'hc2be2318, 32'hc2bd338a, 32'h3fa3ca05, 32'h4190e1f9, 32'h423c4ecf, 32'h41e65fa2};
test_weights[12856:12863] = '{32'hc234f082, 32'hc15b9c09, 32'hc268f942, 32'h41467893, 32'hc0fd3f94, 32'h428a04ce, 32'hc240dcf8, 32'h4184d729};
test_bias[1607:1607] = '{32'hc2c6c522};
test_output[1607:1607] = '{32'h42264e59};
test_input[12864:12871] = '{32'h42bafe83, 32'hc29fb4e2, 32'hc2b870e3, 32'h41bf78fb, 32'h41773965, 32'h41a35568, 32'hc292c226, 32'hc2abe2c7};
test_weights[12864:12871] = '{32'h41a09dce, 32'hc2286c5e, 32'hc24ae63f, 32'hc114c5c2, 32'hc2a1a48d, 32'h42218d2b, 32'h421d7205, 32'h425e4797};
test_bias[1608:1608] = '{32'hc26fc44a};
test_output[1608:1608] = '{32'h44c14e4e};
test_input[12872:12879] = '{32'hc2329b2b, 32'h42abb922, 32'hc1e0d28e, 32'h4260e0f6, 32'hc16c8f80, 32'hc20ae17e, 32'hc115e0a8, 32'hc2903657};
test_weights[12872:12879] = '{32'hc2389a7a, 32'h41da307a, 32'hc0abf502, 32'hc29c0fa9, 32'h40ba0748, 32'hc275bb78, 32'h4281c0c2, 32'h428d0fe8};
test_bias[1609:1609] = '{32'hc2966bd2};
test_output[1609:1609] = '{32'hc55e3024};
test_input[12880:12887] = '{32'hc1aec716, 32'h41295824, 32'hc2771b8d, 32'hbfcd443f, 32'h4297e2a6, 32'hc194cdf0, 32'hc294c308, 32'hc27560c2};
test_weights[12880:12887] = '{32'h42ab676b, 32'hc2a799c2, 32'hc068d261, 32'hc1a4620e, 32'h41bdbd0c, 32'h4272f318, 32'hc24364a1, 32'hc0ebfd6b};
test_bias[1610:1610] = '{32'hc1b2917c};
test_output[1610:1610] = '{32'h450b940e};
test_input[12888:12895] = '{32'h426b9ec9, 32'h425a6f90, 32'hc2590e09, 32'hc2c77e6c, 32'hc28c9663, 32'h41f4eab4, 32'hc00f4863, 32'hc1e8a02f};
test_weights[12888:12895] = '{32'h425571a2, 32'h42b60603, 32'h428e692d, 32'hc2069ef4, 32'h42c7447c, 32'h41ce0510, 32'h42150236, 32'hc1fb3bfc};
test_bias[1611:1611] = '{32'h424cb886};
test_output[1611:1611] = '{32'h450e0281};
test_input[12896:12903] = '{32'h42289382, 32'hc1b75019, 32'hbeffdee2, 32'h429b6aae, 32'hc1e979c8, 32'hc26df56e, 32'hc189531c, 32'h4281e41f};
test_weights[12896:12903] = '{32'h42a72570, 32'hc27258ec, 32'h42ab7f85, 32'h42968e6e, 32'h41a95e66, 32'hc2b30f7a, 32'h41e24274, 32'hc0c1b197};
test_bias[1612:1612] = '{32'hc2161268};
test_output[1612:1612] = '{32'h4662b5c1};
test_input[12904:12911] = '{32'h428037b2, 32'hc232e707, 32'h42a491ba, 32'hc2021636, 32'h42c4bb24, 32'h41c4a87b, 32'hc2b5e0fa, 32'hc1df001b};
test_weights[12904:12911] = '{32'h420437b8, 32'h41c5f1bb, 32'hc287c574, 32'h42c6a7fa, 32'h42a81b06, 32'h422d7f4f, 32'h4208a34a, 32'hc277bf40};
test_bias[1613:1613] = '{32'h42b79516};
test_output[1613:1613] = '{32'h4372249e};
test_input[12912:12919] = '{32'hc2a17f7b, 32'hc207f745, 32'h421f0a55, 32'h4283da4e, 32'h413850e6, 32'h427cac73, 32'hc2165a0b, 32'hc20b185a};
test_weights[12912:12919] = '{32'h4292065c, 32'hc25224d8, 32'h4283bdc8, 32'hc29846a9, 32'h412cb0ca, 32'hc2bf00c7, 32'h426f9db8, 32'h40f99590};
test_bias[1614:1614] = '{32'h41320616};
test_output[1614:1614] = '{32'hc66949f3};
test_input[12920:12927] = '{32'h427fac1c, 32'hc24569e0, 32'h41bb83b8, 32'hc290c846, 32'h423785dc, 32'hc296de1e, 32'h41cda8e0, 32'hc2148d49};
test_weights[12920:12927] = '{32'h4295e290, 32'hc2ba8fa7, 32'hc22b816f, 32'hc23fba7a, 32'hc2923cac, 32'hc1bbd70b, 32'hc28948ac, 32'h42ba5260};
test_bias[1615:1615] = '{32'hc2379c22};
test_output[1615:1615] = '{32'h459c672f};
test_input[12928:12935] = '{32'h419cc2ba, 32'h424af38f, 32'h428083a7, 32'hc22cf776, 32'h420b9b7c, 32'hc2785064, 32'h428e0ce4, 32'hc21e971d};
test_weights[12928:12935] = '{32'hc28b87c8, 32'hc2bc590c, 32'h415f6993, 32'h428d7b90, 32'h42c535ce, 32'h42372bad, 32'h41cfe6fc, 32'hc28ac61a};
test_bias[1616:1616] = '{32'hc2ae986a};
test_output[1616:1616] = '{32'hc547eb2b};
test_input[12936:12943] = '{32'hc1dafcba, 32'h42537866, 32'hc283f08a, 32'hc2368228, 32'hc2b3bde4, 32'hc287198b, 32'h42c0bc90, 32'h40c775a3};
test_weights[12936:12943] = '{32'hc217118f, 32'h4285dcb3, 32'h42029231, 32'hc1fc20c5, 32'hc22339b7, 32'hc2340381, 32'h3f4bf138, 32'hc1ee038f};
test_bias[1617:1617] = '{32'h42770d41};
test_output[1617:1617] = '{32'h462454db};
test_input[12944:12951] = '{32'h408b8765, 32'hbf8a8b5b, 32'h429bb613, 32'hc16f89a3, 32'hc10c61da, 32'h4262d9e9, 32'hc26c0eac, 32'h4139464f};
test_weights[12944:12951] = '{32'hc26fe3a7, 32'hc24b073d, 32'hc2bb6265, 32'hc2944257, 32'hc2c53e7c, 32'hc23ea80f, 32'hc214a7ee, 32'hc29da2e3};
test_bias[1618:1618] = '{32'h4211c371};
test_output[1618:1618] = '{32'hc5d800fd};
test_input[12952:12959] = '{32'h3ff839a2, 32'hc264acd6, 32'hc126376d, 32'h4136c4db, 32'h4210e4cf, 32'h41198643, 32'h428fd453, 32'h427ab9d6};
test_weights[12952:12959] = '{32'h4081e49c, 32'h429f51f6, 32'h42a54ce8, 32'h4061e40c, 32'hc0709263, 32'h4036469c, 32'hc22d00f6, 32'h4209edfe};
test_bias[1619:1619] = '{32'h41e56800};
test_output[1619:1619] = '{32'hc5c7ccf8};
test_input[12960:12967] = '{32'h428d09f7, 32'hc2894996, 32'hc19420d1, 32'hc2915c4c, 32'hc231d737, 32'h428f1c04, 32'hc26d034e, 32'h41b0552d};
test_weights[12960:12967] = '{32'hc2c0050c, 32'h41922f8c, 32'h42355abe, 32'h4296427a, 32'h4205e111, 32'hc29e53e1, 32'hc181be7d, 32'h42bd5ebe};
test_bias[1620:1620] = '{32'h42bcb20e};
test_output[1620:1620] = '{32'hc68f3e4a};
test_input[12968:12975] = '{32'h41ba273d, 32'h42874f8f, 32'h42877f56, 32'hc2945e7a, 32'hc2115ceb, 32'hc207afac, 32'hc255b69c, 32'hc297a0b3};
test_weights[12968:12975] = '{32'hc225e44a, 32'h41f8ed58, 32'h41efa65a, 32'hc2847ab5, 32'h42c2d739, 32'h41f254b3, 32'hc271c0e5, 32'hc2b09e06};
test_bias[1621:1621] = '{32'hc1dcd2a5};
test_output[1621:1621] = '{32'h46519100};
test_input[12976:12983] = '{32'hbe05e5fd, 32'h419043a4, 32'hc259f35d, 32'h4172e0c0, 32'h4244aad6, 32'h4272e31c, 32'h429c7c24, 32'h4280095c};
test_weights[12976:12983] = '{32'h42aa564d, 32'hc27e906c, 32'h426f2cae, 32'h4286c326, 32'h415bc0ca, 32'h41e9e521, 32'hc22f2e50, 32'hc129f352};
test_bias[1622:1622] = '{32'h426bcfe9};
test_output[1622:1622] = '{32'hc59bf85a};
test_input[12984:12991] = '{32'h4266c7ba, 32'hc1c95794, 32'h42a25531, 32'h4145a662, 32'h400c26e2, 32'hc1dc1f9e, 32'hc2358d82, 32'h4228fcb8};
test_weights[12984:12991] = '{32'h42a25a37, 32'hc2ae4fdb, 32'h42574679, 32'hc2bb9395, 32'h4281b962, 32'hc1b4f465, 32'hc22aee4d, 32'hc2935a20};
test_bias[1623:1623] = '{32'hc2554c55};
test_output[1623:1623] = '{32'h46166313};
test_input[12992:12999] = '{32'hbfbfd848, 32'hc0a37517, 32'h42a4fd27, 32'h42b2bb51, 32'hc2911a4f, 32'hc2bf989d, 32'h4269cd03, 32'h424d9564};
test_weights[12992:12999] = '{32'h4286a72e, 32'h41af4b5b, 32'h42a9ab8d, 32'h3f645a53, 32'hc2bd0865, 32'hc214d379, 32'hc1803f12, 32'h423435d0};
test_bias[1624:1624] = '{32'hc0809b9f};
test_output[1624:1624] = '{32'h4691cace};
test_input[13000:13007] = '{32'hc292b024, 32'h42688d3a, 32'h4188d306, 32'hc187f58e, 32'hc2acf4d6, 32'hc27c7786, 32'h42a7d3c8, 32'h4292105b};
test_weights[13000:13007] = '{32'h427749c0, 32'h4295bdc7, 32'h42161ca7, 32'h42291c21, 32'h41dbf15f, 32'hc28d1a8f, 32'hc1d3542e, 32'h41cd73ee};
test_bias[1625:1625] = '{32'hc1d55572};
test_output[1625:1625] = '{32'h44b5332d};
test_input[13008:13015] = '{32'h42a66c57, 32'h41cc8caf, 32'hc17a1720, 32'hc2980a0c, 32'hc2a27a4a, 32'hc2b1f86f, 32'hc22dc9df, 32'hc2a798b9};
test_weights[13008:13015] = '{32'hc2486080, 32'h421085e9, 32'hc2b81033, 32'hc2a6388e, 32'h4198b4e1, 32'h418598e2, 32'hc29c5f9d, 32'h42487a85};
test_bias[1626:1626] = '{32'h42b2c78c};
test_output[1626:1626] = '{32'h443e68de};
test_input[13016:13023] = '{32'h42a67531, 32'hc1a45aaf, 32'hc2362c70, 32'hc1aa1e31, 32'h41b3e87e, 32'hc21805a5, 32'hc13c2b17, 32'h422e02db};
test_weights[13016:13023] = '{32'h42af16a7, 32'hbf2d56e1, 32'hc22b40e7, 32'hc2c11860, 32'h42a37475, 32'hc2662e21, 32'hc07727af, 32'h428eab2a};
test_bias[1627:1627] = '{32'hc1038e44};
test_output[1627:1627] = '{32'h469048e2};
test_input[13024:13031] = '{32'hc29a8902, 32'h421e1484, 32'hc29c8426, 32'h41a7b1dd, 32'h41acd9da, 32'hc2a93246, 32'hc288192d, 32'hc2990c57};
test_weights[13024:13031] = '{32'hbfdb186d, 32'hc23bc12b, 32'h41abc0f6, 32'h42b0441d, 32'h4245ab56, 32'hc1f83a7a, 32'hc12cbd52, 32'hc2a09f7d};
test_bias[1628:1628] = '{32'h422b3fef};
test_output[1628:1628] = '{32'h460d91e3};
test_input[13032:13039] = '{32'h421aa25e, 32'h427e6fc9, 32'h424bfb35, 32'h41ca721b, 32'h41a0a6b6, 32'hc2010153, 32'hc2095ea2, 32'hc2a24102};
test_weights[13032:13039] = '{32'h403499f6, 32'hc14a2434, 32'h42ab7507, 32'hc18312b2, 32'h421d38a7, 32'hc27859ae, 32'h41ddea6f, 32'hc2b0eb30};
test_bias[1629:1629] = '{32'hc296a212};
test_output[1629:1629] = '{32'h463eab33};
test_input[13040:13047] = '{32'h40b67c03, 32'hc1be1709, 32'h41f9da12, 32'hc1c3b8ce, 32'hc2a526bf, 32'h428b9294, 32'h416616b3, 32'hc2348f4c};
test_weights[13040:13047] = '{32'hc2b26951, 32'hc252830b, 32'hc11f3dd4, 32'hc25b5f5e, 32'hc178dcd1, 32'h40e84ca3, 32'hc21732ba, 32'hc27dfdc6};
test_bias[1630:1630] = '{32'h41c6710e};
test_output[1630:1630] = '{32'h45b8b9aa};
test_input[13048:13055] = '{32'h41ec3ca5, 32'hc24194be, 32'h41952bc5, 32'h429eedc9, 32'hc2a1e168, 32'hc2463b8c, 32'hc28ef54b, 32'hc298d524};
test_weights[13048:13055] = '{32'hc2266296, 32'h426abdfc, 32'hc27187b6, 32'hc2ad7e12, 32'hc1f366ba, 32'hc1eba638, 32'hc2c76a93, 32'hc2a8008e};
test_bias[1631:1631] = '{32'h428a5d85};
test_output[1631:1631] = '{32'h45aa50ef};
test_input[13056:13063] = '{32'hc1a469ab, 32'h428c15b9, 32'hc2026ad7, 32'hc2a8f44b, 32'hc21c2b2d, 32'hc0a5077f, 32'hc28be791, 32'hc23c7bc6};
test_weights[13056:13063] = '{32'hc1dca59e, 32'hc29677a3, 32'hc29c4486, 32'hc286e648, 32'h419c7229, 32'h4288cfd8, 32'hc263ce2d, 32'h41968ab9};
test_bias[1632:1632] = '{32'h420505db};
test_output[1632:1632] = '{32'h45ada723};
test_input[13064:13071] = '{32'hc1dc2db2, 32'h419bbe06, 32'hc2024be1, 32'hc1c68d5a, 32'hc2bc97c8, 32'hc2afd7b0, 32'h42068409, 32'h41b95bc0};
test_weights[13064:13071] = '{32'h42084337, 32'hc28b35d4, 32'hc26ef5e6, 32'h420a879c, 32'hc2aab1d0, 32'hc25963ff, 32'h42bd594f, 32'hc22620e5};
test_bias[1633:1633] = '{32'hc19f9ffb};
test_output[1633:1633] = '{32'h4657f688};
test_input[13072:13079] = '{32'hc29725c8, 32'h4286e10a, 32'hc28c5f24, 32'h41bab219, 32'hc2a91c0b, 32'hc20d23d1, 32'h429137a8, 32'hc2a4b738};
test_weights[13072:13079] = '{32'hc29b365f, 32'h4295c204, 32'h42040a18, 32'hc28da17f, 32'hc257689e, 32'h409fac90, 32'h41d4162c, 32'hc1a1372e};
test_bias[1634:1634] = '{32'h4043a8fd};
test_output[1634:1634] = '{32'h4668f98f};
test_input[13080:13087] = '{32'hc279d110, 32'hc29907c3, 32'hc28fc991, 32'hc22142e9, 32'hc28f8a02, 32'h3fca0ea8, 32'h3f4030ee, 32'hc2b6a6e9};
test_weights[13080:13087] = '{32'h42b5a9d4, 32'h42c38a0e, 32'hc234d551, 32'h4196275d, 32'hc1f3c63a, 32'h429f5f38, 32'h421f1f84, 32'h423cf84c};
test_bias[1635:1635] = '{32'h404cbcb6};
test_output[1635:1635] = '{32'hc6455359};
test_input[13088:13095] = '{32'h4210099c, 32'h42c0747c, 32'hc1cf259e, 32'h41be963b, 32'hc18ce0c4, 32'hc26c99f0, 32'h42927feb, 32'h4283f1b9};
test_weights[13088:13095] = '{32'h41ac3c4e, 32'h42bb7aaf, 32'h42834f1b, 32'hc1c284ae, 32'h42a6f733, 32'h42999828, 32'h428bf14b, 32'h3f38969b};
test_bias[1636:1636] = '{32'h40ad016d};
test_output[1636:1636] = '{32'h45d0cfe2};
test_input[13096:13103] = '{32'hc2a07245, 32'h429b2cae, 32'hc2283edd, 32'hc2adf95b, 32'h42c6d435, 32'hc2a69301, 32'h4124f043, 32'h429dac15};
test_weights[13096:13103] = '{32'hc2219e08, 32'hc233afb0, 32'hc20efa65, 32'hc23f641a, 32'h4298cc4b, 32'h4221916d, 32'hc288a28d, 32'hc29ef85e};
test_bias[1637:1637] = '{32'h42212c29};
test_output[1637:1637] = '{32'h452a2639};
test_input[13104:13111] = '{32'h41e1fe70, 32'hc2157dc3, 32'h404ff2e9, 32'h41b05d38, 32'hc1db2cdb, 32'hc255ee22, 32'hc222e8c2, 32'hc20db23a};
test_weights[13104:13111] = '{32'hc24bd3bc, 32'hc29267c6, 32'h42b3ce6e, 32'h420b2862, 32'h40a7a91e, 32'h426a44b4, 32'h42b8d39e, 32'h41f92792};
test_bias[1638:1638] = '{32'h428560f9};
test_output[1638:1638] = '{32'hc5b2c67a};
test_input[13112:13119] = '{32'hc20fa54a, 32'h429aa60a, 32'h41d87285, 32'hc2a6c3bb, 32'hc1b08bc3, 32'h42003745, 32'hc2b7402a, 32'hc23ff531};
test_weights[13112:13119] = '{32'h42a6ba13, 32'hc1a37132, 32'h42bcb605, 32'h42b140db, 32'hc2677681, 32'h421a95f1, 32'hc2b8e01c, 32'hc229afac};
test_bias[1639:1639] = '{32'h41d2abb9};
test_output[1639:1639] = '{32'h456350c4};
test_input[13120:13127] = '{32'h41cbb07b, 32'hc21e1575, 32'hc2a75744, 32'hc281a0ab, 32'hc2ac31c0, 32'hc1a6385e, 32'hc25e1fb7, 32'h4235bca5};
test_weights[13120:13127] = '{32'h41f53fc8, 32'h418389f2, 32'h429222b9, 32'hc2b9243d, 32'hc28942de, 32'h42a37915, 32'h4276b448, 32'hc1e7b4fc};
test_bias[1640:1640] = '{32'h41addfd1};
test_output[1640:1640] = '{32'hc3f5c472};
test_input[13128:13135] = '{32'h416f0ef1, 32'h3f4b71bd, 32'hc2236f66, 32'h42bfc27c, 32'h42905b81, 32'h429f57a3, 32'h420a5a8e, 32'hc0267043};
test_weights[13128:13135] = '{32'hc291735f, 32'hc28927cf, 32'hc20f31af, 32'h428cb88b, 32'hc2b7ef31, 32'h41533207, 32'hc2b2e8a8, 32'h41f5c8b8};
test_bias[1641:1641] = '{32'h427a4235};
test_output[1641:1641] = '{32'hc4cbc3fb};
test_input[13136:13143] = '{32'h42283029, 32'hc1ccf107, 32'h423b5dcb, 32'h413fdd02, 32'hc280a3eb, 32'h429438c0, 32'hc1cdb0d3, 32'hc2ad3245};
test_weights[13136:13143] = '{32'hc1df6e2f, 32'hc1caca59, 32'h429aed58, 32'hc2aa93a2, 32'hc1c5c01c, 32'hc12c7ca7, 32'hc21d9634, 32'h42b48619};
test_bias[1642:1642] = '{32'h42ac26d4};
test_output[1642:1642] = '{32'hc5705b07};
test_input[13144:13151] = '{32'hc14a5a28, 32'hc264b7bb, 32'hc11f3b37, 32'h42312b6c, 32'h4292db9d, 32'hbfc766f9, 32'hc295a49b, 32'h427bee10};
test_weights[13144:13151] = '{32'h42aebfe1, 32'h423904a8, 32'h42417370, 32'hc22b7694, 32'hc16cf4ae, 32'h41139cf3, 32'hc1f40aa6, 32'h4249df4c};
test_bias[1643:1643] = '{32'hc1e141c4};
test_output[1643:1643] = '{32'hc4e0d6df};
test_input[13152:13159] = '{32'h426f4be0, 32'h42a4e77f, 32'h42921967, 32'hc1f6cec2, 32'h41182fe1, 32'hc2b1e7cc, 32'hc148e723, 32'h41ba6551};
test_weights[13152:13159] = '{32'hc24c39c3, 32'hc1905d1e, 32'hc21c7e4c, 32'hc105bf51, 32'h429be97d, 32'h4264b1b3, 32'hc21f958a, 32'h42708056};
test_bias[1644:1644] = '{32'h42028b86};
test_output[1644:1644] = '{32'hc6154079};
test_input[13160:13167] = '{32'h424a1280, 32'hc2a28118, 32'h4205ae08, 32'h419e1f2c, 32'hc27e7065, 32'h42b6b52d, 32'hc2618e66, 32'hc24b4381};
test_weights[13160:13167] = '{32'hc2590894, 32'hc1a7933a, 32'hc2798023, 32'h41c8a8d1, 32'hc20188b5, 32'h42b55154, 32'h41e6baef, 32'hc29f7ca8};
test_bias[1645:1645] = '{32'hc297a34d};
test_output[1645:1645] = '{32'h461d40a8};
test_input[13168:13175] = '{32'hc1206ab4, 32'h41caae71, 32'hc229526b, 32'hc1ca7c9b, 32'h42897184, 32'h42837e33, 32'h41e629d5, 32'hc284de3a};
test_weights[13168:13175] = '{32'h4204beda, 32'hc2054537, 32'h429f3d96, 32'hc2803e8c, 32'hc13eb36e, 32'h42c118b2, 32'h42128e57, 32'h428da833};
test_bias[1646:1646] = '{32'hc1a9b930};
test_output[1646:1646] = '{32'hc4858376};
test_input[13176:13183] = '{32'hc1904ef8, 32'h410fe426, 32'hc20c2179, 32'h4263c513, 32'hc2c0a493, 32'h41d8c164, 32'hc290ca53, 32'hc24b59df};
test_weights[13176:13183] = '{32'hc2a0fe67, 32'h4088d8e7, 32'h41d5f2cc, 32'hc2297d8c, 32'h3f814943, 32'hc186693c, 32'h42bc1624, 32'hc1c1f214};
test_bias[1647:1647] = '{32'hc2a1f515};
test_output[1647:1647] = '{32'hc5fc23eb};
test_input[13184:13191] = '{32'h4219ef20, 32'h429d1edc, 32'h40a6c7b7, 32'h42a2ea33, 32'hc2066ce0, 32'h42414a96, 32'hc29ad728, 32'hc1e8344d};
test_weights[13184:13191] = '{32'h40f98d28, 32'h41fd53a8, 32'h42773c31, 32'h4246939d, 32'h429caf52, 32'h42bd19b5, 32'hbfb61a7d, 32'hc2551f60};
test_bias[1648:1648] = '{32'h419ee9ce};
test_output[1648:1648] = '{32'h462839d4};
test_input[13192:13199] = '{32'hc1b43676, 32'h413e1625, 32'hc15ae350, 32'hc2845e93, 32'h4232891a, 32'hc217a3ba, 32'hc245915d, 32'hc2b66a54};
test_weights[13192:13199] = '{32'hc265d5e4, 32'h3f8870a1, 32'hc23452cc, 32'h41c599da, 32'hc2b7c1d9, 32'hc280b6b5, 32'h4180bfd0, 32'h42ae27a1};
test_bias[1649:1649] = '{32'h42605bb4};
test_output[1649:1649] = '{32'hc61d1465};
test_input[13200:13207] = '{32'h42b070ec, 32'hc022843c, 32'hc23dd872, 32'hc260c439, 32'hc23a5b1b, 32'h3f29dae4, 32'h4196c804, 32'h42a6d78b};
test_weights[13200:13207] = '{32'h412fd47a, 32'hc0bad40f, 32'h428a72eb, 32'h40aa0754, 32'hc1ce6f61, 32'h42ade62b, 32'hc1a2c263, 32'hc0e38b10};
test_bias[1650:1650] = '{32'hc0aaf28c};
test_output[1650:1650] = '{32'hc5111d4b};
test_input[13208:13215] = '{32'hc2a97557, 32'h428387dd, 32'h420f0bb8, 32'h41f7f858, 32'h418fab34, 32'hc21cef0f, 32'hc2939c5e, 32'hbfe73260};
test_weights[13208:13215] = '{32'h421ad923, 32'hc2b01257, 32'hc1d1e87b, 32'h42a544c5, 32'h4236c27e, 32'hc23e3639, 32'h42c305fc, 32'hc2aa2a4d};
test_bias[1651:1651] = '{32'hc20f7c55};
test_output[1651:1651] = '{32'hc638fe6f};
test_input[13216:13223] = '{32'h426cfba5, 32'hc28aed2c, 32'h42790eb6, 32'hc29de794, 32'h42c031bd, 32'h418799ef, 32'hc22b5bfd, 32'h42a29eac};
test_weights[13216:13223] = '{32'h41a11e2b, 32'h42c67961, 32'h4242c61e, 32'h42250ad8, 32'h41adfae4, 32'hc1c697b4, 32'hc2bdc081, 32'hc2622036};
test_bias[1652:1652] = '{32'hc2acf78f};
test_output[1652:1652] = '{32'hc5985ae5};
test_input[13224:13231] = '{32'hc1ffbe96, 32'h4228dc07, 32'h429931e3, 32'h42ade58e, 32'hc272d21d, 32'hc2b912e7, 32'hc10a65c1, 32'hc0aa47cc};
test_weights[13224:13231] = '{32'h4197d66b, 32'hc2018e42, 32'h424d7a8b, 32'hc2aeb60a, 32'hc19ae76f, 32'hc284da7e, 32'hc2163ebb, 32'h424eb4a2};
test_bias[1653:1653] = '{32'hc2c2146a};
test_output[1653:1653] = '{32'h44cd11fa};
test_input[13232:13239] = '{32'h41c4161a, 32'h3f3e6174, 32'h42a95256, 32'h422bf684, 32'hc181fc85, 32'h42a37772, 32'hc2c7381d, 32'h4185b592};
test_weights[13232:13239] = '{32'hc0f0965a, 32'hc15e872f, 32'h428fd34c, 32'h42934474, 32'h425a1664, 32'hc2819385, 32'h42573bf7, 32'hc1c1ee3e};
test_bias[1654:1654] = '{32'h42a5c6d3};
test_output[1654:1654] = '{32'hc52f439f};
test_input[13240:13247] = '{32'hc199d611, 32'h42a268f9, 32'h41f2175e, 32'hc25af53a, 32'hc293a8c7, 32'h4286cdbd, 32'hc28ed5c7, 32'h42c66670};
test_weights[13240:13247] = '{32'hc00c97a2, 32'h40c2869d, 32'hc139c46e, 32'h410efd93, 32'hc21f5a40, 32'h410a41f0, 32'h42ba14b2, 32'hc1e795a8};
test_bias[1655:1655] = '{32'h4198d9d6};
test_output[1655:1655] = '{32'hc5c43227};
test_input[13248:13255] = '{32'h420b9db0, 32'h427d65b6, 32'hc28268e1, 32'hc1b95250, 32'hc24fae42, 32'h429134a4, 32'hc241b0e4, 32'hc232001d};
test_weights[13248:13255] = '{32'h42c75e7c, 32'hc27d701a, 32'hc1a675ee, 32'h42842ccc, 32'h4278c819, 32'h42be9551, 32'h42a32514, 32'h42a18aec};
test_bias[1656:1656] = '{32'hc299e159};
test_output[1656:1656] = '{32'hc5910470};
test_input[13256:13263] = '{32'hc275844e, 32'hc2560a4f, 32'h42a51386, 32'h42754392, 32'h41eb84f7, 32'h42b0bf84, 32'h426de8a3, 32'hc2887d8a};
test_weights[13256:13263] = '{32'hc2861271, 32'hc2b1d094, 32'h429c57b2, 32'h41f5eeaf, 32'h4297e64c, 32'h41f7b6fa, 32'h40bc4c55, 32'h4292f093};
test_bias[1657:1657] = '{32'h40cb598d};
test_output[1657:1657] = '{32'h4688e7c7};
test_input[13264:13271] = '{32'h42608e51, 32'h4099a7cc, 32'h41fdf6c2, 32'hc29bdd09, 32'h42816f42, 32'h421ae00a, 32'hc2246e56, 32'hc245f4bd};
test_weights[13264:13271] = '{32'h4270e960, 32'h4253b0b8, 32'h4226d55c, 32'hc1dcdb5b, 32'h42017054, 32'h42a326de, 32'hc2409473, 32'h4281c670};
test_bias[1658:1658] = '{32'hc202ae3d};
test_output[1658:1658] = '{32'h462d6b12};
test_input[13272:13279] = '{32'h4290b2ac, 32'hc2816313, 32'hc1c5ed21, 32'h414966c2, 32'hc22001d6, 32'h417bdf27, 32'hc2945cc4, 32'hc1e73860};
test_weights[13272:13279] = '{32'h41ba8187, 32'h42342895, 32'h425c9fc9, 32'hc29ae43c, 32'h42bdb7c7, 32'hc29ef42b, 32'h4219f923, 32'hc22a93b0};
test_bias[1659:1659] = '{32'h42b2e9a8};
test_output[1659:1659] = '{32'hc61e86c1};
test_input[13280:13287] = '{32'h427b6c69, 32'h4241a3ef, 32'hc15bcab0, 32'h4095e3e7, 32'h41e66dc1, 32'h3fba73a1, 32'hc05fecc6, 32'h40e0745b};
test_weights[13280:13287] = '{32'h42b13a58, 32'h42665d0a, 32'h42a6b53d, 32'h41c67c6c, 32'h416194da, 32'hc2033ed6, 32'hc2b780d1, 32'hc20721e6};
test_bias[1660:1660] = '{32'hc197d7d0};
test_output[1660:1660] = '{32'h45f2439e};
test_input[13288:13295] = '{32'h421416fe, 32'h4139d255, 32'hc153455c, 32'h42a60d8b, 32'hc29826ab, 32'hc27fe72f, 32'h428fe7c5, 32'hc2abadf7};
test_weights[13288:13295] = '{32'hc227dcbc, 32'h41ca5bb5, 32'h425b557c, 32'hc28e985a, 32'hc23b3ef8, 32'hc1a962c7, 32'hc23430c2, 32'h42c5b018};
test_bias[1661:1661] = '{32'hc21ef720};
test_output[1661:1661] = '{32'hc6668617};
test_input[13296:13303] = '{32'hc265a537, 32'h429242cc, 32'h4205a59f, 32'hc22f12e4, 32'hc24ffd79, 32'h425622c0, 32'hc2acdea7, 32'hc2bb7928};
test_weights[13296:13303] = '{32'h41b6892c, 32'hc2b2ef04, 32'h41bd554a, 32'hc287acc3, 32'hc2af8042, 32'hc2543ecb, 32'hc190feb8, 32'hc26ba3e3};
test_bias[1662:1662] = '{32'h418a8737};
test_output[1662:1662] = '{32'h4593faa4};
test_input[13304:13311] = '{32'h41d4deea, 32'h429a015f, 32'hc27b065b, 32'hc1ff55ef, 32'hc29277ca, 32'hc2255967, 32'hc17c3a55, 32'h42969a0d};
test_weights[13304:13311] = '{32'h42b3d07e, 32'h425613fb, 32'hc1157db2, 32'h42aba7af, 32'h4211f4fc, 32'hc16eeccd, 32'hc284ca31, 32'h427f6f90};
test_bias[1663:1663] = '{32'hc21b8a79};
test_output[1663:1663] = '{32'h45fdcf45};
test_input[13312:13319] = '{32'h4258b64f, 32'hc2abebf5, 32'hc29206a9, 32'hc2c2510a, 32'h42a158f6, 32'h40409587, 32'h423a14ee, 32'h42c2c1ea};
test_weights[13312:13319] = '{32'h42c4660e, 32'h42acf48f, 32'hc1129e64, 32'hc2560c9d, 32'hc2155bb8, 32'hc2371cce, 32'h41cc2eae, 32'h4292634a};
test_bias[1664:1664] = '{32'hc280d83a};
test_output[1664:1664] = '{32'h460a5c9b};
test_input[13320:13327] = '{32'hc2084cad, 32'h4244511f, 32'hc286ae5c, 32'hc20c2840, 32'h4298b179, 32'h428fb585, 32'h424d5df8, 32'h4194f3b5};
test_weights[13320:13327] = '{32'hc26cc64b, 32'h41ccff29, 32'h41e517cd, 32'hc2aa7010, 32'h42558d08, 32'hc1a7c5df, 32'hc1745e01, 32'h42858b26};
test_bias[1665:1665] = '{32'h41c7b72f};
test_output[1665:1665] = '{32'h45e6caf7};
test_input[13328:13335] = '{32'hc183fe28, 32'h4231291b, 32'hc26eb541, 32'hc2878980, 32'hc14f94d2, 32'h42424174, 32'h405791f2, 32'h42a7fe18};
test_weights[13328:13335] = '{32'hc2206849, 32'h41e3c2fd, 32'hc1c3bcdf, 32'h42763a6f, 32'h410ed722, 32'hc28c20bc, 32'h424c6b8e, 32'hc1cc3e7a};
test_bias[1666:1666] = '{32'hc18c131c};
test_output[1666:1666] = '{32'hc5c4c938};
test_input[13336:13343] = '{32'h424884c9, 32'h427127b9, 32'hc2c07c1e, 32'hc0ed21e2, 32'h42b988c6, 32'h42521c5d, 32'hc289b567, 32'h41fe1a8e};
test_weights[13336:13343] = '{32'hc21c0032, 32'hc2623467, 32'h428a7728, 32'hc28b8ccb, 32'hc185865c, 32'hc28ad819, 32'hc276a125, 32'h429b56de};
test_bias[1667:1667] = '{32'h41bd65ed};
test_output[1667:1667] = '{32'hc61bc58c};
test_input[13344:13351] = '{32'hc22a603a, 32'hc1cb7820, 32'hc20780c2, 32'hc2a996b4, 32'hc2bd9f09, 32'hc20e130a, 32'h42a094d6, 32'hbf2ee825};
test_weights[13344:13351] = '{32'hc22fdb55, 32'h428d1385, 32'h422e096c, 32'h42a51a09, 32'h41e6e972, 32'hc255047f, 32'h409065fb, 32'hc2593e18};
test_bias[1668:1668] = '{32'h41a42ab2};
test_output[1668:1668] = '{32'hc609d15d};
test_input[13352:13359] = '{32'h429629b3, 32'h426f8a80, 32'h4136fcc7, 32'h40d251b9, 32'hc1ed9e97, 32'hc22b022a, 32'h41db28d6, 32'hc0cf4ea5};
test_weights[13352:13359] = '{32'hc214a478, 32'h41d73c8b, 32'h420ff26d, 32'hc270ca98, 32'hc1b9ae0c, 32'h428a9d94, 32'h428c4f84, 32'hc2533d9a};
test_bias[1669:1669] = '{32'hc2922166};
test_output[1669:1669] = '{32'hc49bb561};
test_input[13360:13367] = '{32'h3f097ff1, 32'hc26d6861, 32'h412f6d6c, 32'h42b7aadb, 32'h42b8edbb, 32'h4257cc5a, 32'hc29d4e85, 32'h40af358a};
test_weights[13360:13367] = '{32'h42707400, 32'hc28193b0, 32'h42b8247e, 32'h41ea5886, 32'h41f36737, 32'h4267328c, 32'h423343b8, 32'hc2bc3076};
test_bias[1670:1670] = '{32'hc1351b31};
test_output[1670:1670] = '{32'h4613c50c};
test_input[13368:13375] = '{32'hc2c1d09c, 32'h42abb32e, 32'h42a8ddf9, 32'h422ebecc, 32'hc2a0cdeb, 32'h409cef39, 32'h41e9bbed, 32'hc27f4062};
test_weights[13368:13375] = '{32'hc1932350, 32'hc2b7b125, 32'h4213c18f, 32'hc185fcaf, 32'h421c28b4, 32'h41e0a36f, 32'hc0aa23ff, 32'h42101945};
test_bias[1671:1671] = '{32'h425d7fc5};
test_output[1671:1671] = '{32'hc60e6d8f};
test_input[13376:13383] = '{32'h40f7bd26, 32'hc1e803ed, 32'h4218c177, 32'h42400254, 32'hc0a3f1df, 32'h4203fc8b, 32'hc23c8ac4, 32'hc2a6069a};
test_weights[13376:13383] = '{32'h421f64f7, 32'hc0847d34, 32'h42af893f, 32'h42a32081, 32'hc25b634d, 32'hc2c3e6f6, 32'h42696d13, 32'h42b86bf5};
test_bias[1672:1672] = '{32'h42affee4};
test_output[1672:1672] = '{32'hc5ae26b2};
test_input[13384:13391] = '{32'hc224fe91, 32'h419ad47d, 32'hc1a1225a, 32'hc22c4398, 32'hc2881e95, 32'hc1cfa749, 32'hc26c901c, 32'h42545cc4};
test_weights[13384:13391] = '{32'h42b49ec8, 32'hc1ec67b0, 32'hc174e7a7, 32'h4284ec22, 32'h42c31642, 32'h429465ca, 32'h423c2da6, 32'hc292f5f0};
test_bias[1673:1673] = '{32'h42c0bcf1};
test_output[1673:1673] = '{32'hc6abe577};
test_input[13392:13399] = '{32'hc201b50b, 32'h41672d1e, 32'hc281be61, 32'h415099d7, 32'hc11a62e4, 32'hc11b2619, 32'h42c7e707, 32'hc18486c8};
test_weights[13392:13399] = '{32'h408bcb27, 32'h42bd5407, 32'h412c5907, 32'hc1ec7f81, 32'hc214b1a4, 32'h41e60fe7, 32'hc2a6fe52, 32'h4294cf9d};
test_bias[1674:1674] = '{32'h428e9645};
test_output[1674:1674] = '{32'hc61114a7};
test_input[13400:13407] = '{32'h42bf6eba, 32'hc2350d05, 32'hc27fd50e, 32'h41f5984a, 32'h42b6192b, 32'h423d4c3b, 32'hc26efb5f, 32'h424264a9};
test_weights[13400:13407] = '{32'hc1c339c3, 32'h4237e243, 32'h41f4a873, 32'h4117860a, 32'h42174a88, 32'h41c7f48b, 32'h42b74adc, 32'hc21d53cb};
test_bias[1675:1675] = '{32'hc14a5265};
test_output[1675:1675] = '{32'hc60a5b1d};
test_input[13408:13415] = '{32'hc2c01679, 32'hc2ba2176, 32'hc24841f7, 32'hc164a2d8, 32'h413ad0b0, 32'hc1cca534, 32'h42c42ff4, 32'hc29d41e2};
test_weights[13408:13415] = '{32'h429f8f8d, 32'h42076d16, 32'hc0cbeaab, 32'h420f5d34, 32'h427d4ef7, 32'hc10a98e6, 32'hc28f47f1, 32'h42b8d38f};
test_bias[1676:1676] = '{32'h4114ad50};
test_output[1676:1676] = '{32'hc6be13e1};
test_input[13416:13423] = '{32'hc21702f9, 32'hc2a5e30e, 32'h41debedc, 32'hc19d29c2, 32'h423a1565, 32'h423ceee9, 32'hc26fb1d7, 32'hc242c80f};
test_weights[13416:13423] = '{32'h428f2466, 32'hc1c1b6c2, 32'h425f3338, 32'hc19c828b, 32'hc2826558, 32'h4185600d, 32'h4231e268, 32'hc2222fa0};
test_bias[1677:1677] = '{32'h4203b815};
test_output[1677:1677] = '{32'hc4cf5747};
test_input[13424:13431] = '{32'h425e524b, 32'h42c46970, 32'h4286237c, 32'h42b1b014, 32'hc2a7efd5, 32'hc2b0c0e7, 32'h4191a277, 32'h425b54c4};
test_weights[13424:13431] = '{32'hc1d476e7, 32'hc1bd131a, 32'hc187e9cd, 32'hc29d8756, 32'hc25cff3a, 32'hc2728ace, 32'h424d105e, 32'h424e3830};
test_bias[1678:1678] = '{32'h42c7563f};
test_output[1678:1678] = '{32'h44f06f33};
test_input[13432:13439] = '{32'h42a885c3, 32'hc206f388, 32'h414b4867, 32'hc1f4dcc6, 32'hc2432b4e, 32'h421caddf, 32'hc24f2973, 32'hc2a92c83};
test_weights[13432:13439] = '{32'hc183facb, 32'h424f2620, 32'h4286aa65, 32'hc2aa0dc9, 32'hc273080d, 32'hc20cfeb9, 32'h42c6f064, 32'hc22c76ce};
test_bias[1679:1679] = '{32'h4146d7fb};
test_output[1679:1679] = '{32'h43ce34d3};
test_input[13440:13447] = '{32'h409105f9, 32'h4107f980, 32'h4222ff14, 32'hc290ff6b, 32'h4237a4b8, 32'h4211a484, 32'h42469224, 32'hc2994302};
test_weights[13440:13447] = '{32'h42224094, 32'hc2863d1a, 32'hc2ab1bd3, 32'h428a84ab, 32'h42af0a41, 32'hc2814986, 32'hc29c13bf, 32'hc218b372};
test_bias[1680:1680] = '{32'hc2019be1};
test_output[1680:1680] = '{32'hc6004ac2};
test_input[13448:13455] = '{32'h42b42183, 32'h42545620, 32'h427cb392, 32'h425df084, 32'h42249b72, 32'hc23d540d, 32'h42b17fe2, 32'h428cf308};
test_weights[13448:13455] = '{32'hc28a6d36, 32'h423de7c0, 32'hc295a6fb, 32'hc225b30c, 32'h40e9b671, 32'hc0da277d, 32'h42a86136, 32'hc2886909};
test_bias[1681:1681] = '{32'h4297a766};
test_output[1681:1681] = '{32'hc5e677a5};
test_input[13456:13463] = '{32'h417f340f, 32'hc1ea8d5d, 32'hc11e951b, 32'h422dd0a4, 32'hc25c8f0e, 32'h428fdb64, 32'h41a2cb97, 32'hc2b33029};
test_weights[13456:13463] = '{32'hc24f2c7c, 32'hc17388b3, 32'hc13e8560, 32'hc13b05c5, 32'hc2c0f320, 32'h42bdbcbe, 32'hc2bf65b8, 32'h420fd8a2};
test_bias[1682:1682] = '{32'h42b321e9};
test_output[1682:1682] = '{32'h45c4ae71};
test_input[13464:13471] = '{32'hc285d07b, 32'hc2430f73, 32'hc2b78b05, 32'hc11020d7, 32'hc235769d, 32'h4153a31d, 32'hc21764c4, 32'hc1620760};
test_weights[13464:13471] = '{32'hc1f71cab, 32'hc2c59bfa, 32'hc207e9a5, 32'h42990c59, 32'h41110868, 32'h42050743, 32'hc0c245bb, 32'h42bcc561};
test_bias[1683:1683] = '{32'hc2133e85};
test_output[1683:1683] = '{32'h46002860};
test_input[13472:13479] = '{32'hc2255ef6, 32'h42524749, 32'hc2025119, 32'h41598aa6, 32'h425cfed1, 32'h429ea3d4, 32'hc287e0df, 32'hc2c21370};
test_weights[13472:13479] = '{32'h4225216b, 32'h40eaad25, 32'h40e33408, 32'hc292f414, 32'hc2c3fa7a, 32'h42708a83, 32'h41764970, 32'hc1887a67};
test_bias[1684:1684] = '{32'h42025880};
test_output[1684:1684] = '{32'hc51f9280};
test_input[13480:13487] = '{32'hc23cb867, 32'hc10a2554, 32'h42974ba0, 32'hc294e828, 32'hc21fc61d, 32'hc006ff1e, 32'hc16fa64b, 32'hc1d000ca};
test_weights[13480:13487] = '{32'hc2234524, 32'h421a8843, 32'h41a8b296, 32'h42ba3de2, 32'hc24fee69, 32'hc27991a3, 32'hc18929d6, 32'h429ada37};
test_bias[1685:1685] = '{32'hbff5cb97};
test_output[1685:1685] = '{32'hc54e000e};
test_input[13488:13495] = '{32'hbf586653, 32'hc1f20c49, 32'hc2a2b057, 32'h427baaa5, 32'hc29ea769, 32'hc20dc48e, 32'h4212c33a, 32'hc1bc20b6};
test_weights[13488:13495] = '{32'hc2629137, 32'hc221bd38, 32'hc26743fe, 32'h3fb36046, 32'hc29fe60e, 32'hc2b72e31, 32'hc2a9df24, 32'h4021b99f};
test_bias[1686:1686] = '{32'h41944ef4};
test_output[1686:1686] = '{32'h46433618};
test_input[13496:13503] = '{32'h4087f1b4, 32'hc1a3a63b, 32'hc2b58608, 32'hc284ef21, 32'hc279a814, 32'hc2bc359d, 32'h4287ad65, 32'hc202b367};
test_weights[13496:13503] = '{32'h421fc314, 32'h42880712, 32'h42289b51, 32'h414ac3c0, 32'h42838051, 32'h3ffd43d2, 32'hc2927755, 32'hc283f59d};
test_bias[1687:1687] = '{32'hc2a2c8c1};
test_output[1687:1687] = '{32'hc64c44cd};
test_input[13504:13511] = '{32'hc2c78661, 32'h425ab3c4, 32'h4247c19f, 32'h428f2e3c, 32'h408725fb, 32'h428bcf92, 32'h42a34582, 32'h429f2149};
test_weights[13504:13511] = '{32'hc2c12207, 32'h42b8fd71, 32'h4205172c, 32'h40b61e21, 32'hc05e7e46, 32'h428483d9, 32'hc28613f6, 32'hc07e8171};
test_bias[1688:1688] = '{32'hc270f1f3};
test_output[1688:1688] = '{32'h46729e7a};
test_input[13512:13519] = '{32'hc237961b, 32'h4287e5bd, 32'h426a3ed1, 32'hbfb6fccd, 32'h4286f78d, 32'h42c3e67c, 32'h423f3532, 32'h41d1a6c1};
test_weights[13512:13519] = '{32'hc26a7b85, 32'hc1a50f67, 32'hc2863b26, 32'h422cf8f2, 32'h424fdf43, 32'h429ba553, 32'hc21fdce8, 32'h41a2b6ed};
test_bias[1689:1689] = '{32'hc1e0f4ba};
test_output[1689:1689] = '{32'h45db6467};
test_input[13520:13527] = '{32'hbc4949ee, 32'hc20a69ab, 32'hc2445ad7, 32'h426e7be0, 32'hc268a918, 32'hc2290157, 32'hc23d55e1, 32'h4299cee5};
test_weights[13520:13527] = '{32'h427f7ce7, 32'h4280a96f, 32'hc28c0ba0, 32'hc1edba13, 32'hc2940a62, 32'h4262bb09, 32'h42c2f4e4, 32'h42a11a89};
test_bias[1690:1690] = '{32'hc25a2bda};
test_output[1690:1690] = '{32'h4533b79e};
test_input[13528:13535] = '{32'hbfc276fe, 32'h421039cb, 32'h420592a1, 32'hc2b3c2a2, 32'h42561cc7, 32'hc2b33e8e, 32'h41cfe543, 32'h42214ed0};
test_weights[13528:13535] = '{32'h42864a14, 32'hc24771c0, 32'hc2a0e4ac, 32'hc1c3c62f, 32'hc28c214d, 32'hc2842aee, 32'hc2955e98, 32'h42c50910};
test_bias[1691:1691] = '{32'h4228fb81};
test_output[1691:1691] = '{32'h44e8799d};
test_input[13536:13543] = '{32'hc28800e6, 32'hc29e3627, 32'h426f9112, 32'hc2b3d7c9, 32'h42914837, 32'hc28f85dc, 32'h422c0fe2, 32'hc0d4bff1};
test_weights[13536:13543] = '{32'h42189d4e, 32'hc06e6115, 32'hc1b1007b, 32'h42a2b42b, 32'h40c1dc53, 32'h42b00454, 32'h41f8084d, 32'h419d2020};
test_bias[1692:1692] = '{32'h42aeb909};
test_output[1692:1692] = '{32'hc672957e};
test_input[13544:13551] = '{32'h425fde1f, 32'hc1bc526d, 32'h42b66b21, 32'h42b919ce, 32'h4276b7e5, 32'hc1b30ed1, 32'h42b5e3c0, 32'h4280ef87};
test_weights[13544:13551] = '{32'h420d2d77, 32'h415fbd53, 32'hc2c76ba3, 32'hc24423f1, 32'hc0ac209b, 32'hc2888eea, 32'h42ac34a8, 32'hc274fe55};
test_bias[1693:1693] = '{32'h41d653fc};
test_output[1693:1693] = '{32'hc5d70a0e};
test_input[13552:13559] = '{32'h42c48e25, 32'h42b5965b, 32'hc21c632f, 32'hc223ce63, 32'hc24070e7, 32'hc27b11b6, 32'h42c6dcdc, 32'hc2727044};
test_weights[13552:13559] = '{32'hc25c8b99, 32'h42a3dc4b, 32'h41f269d1, 32'hc22bffe9, 32'hc254bba6, 32'hc2437d46, 32'hc2869403, 32'h42bd78ac};
test_bias[1694:1694] = '{32'h4123a33c};
test_output[1694:1694] = '{32'hc5833e35};
test_input[13560:13567] = '{32'hc27c7c55, 32'hc142a009, 32'hc2989e99, 32'hc23a807e, 32'hc28f018b, 32'h42489003, 32'h3ef8c1bf, 32'hc2877b03};
test_weights[13560:13567] = '{32'hc1cb04e1, 32'hc2855aff, 32'hc22b71f1, 32'h42266f14, 32'h40d9b403, 32'hc2c20993, 32'h41c711ac, 32'hc21fc074};
test_bias[1695:1695] = '{32'hc2b00241};
test_output[1695:1695] = '{32'h447f86f3};
test_input[13568:13575] = '{32'h41683877, 32'h42582a22, 32'h403efd0c, 32'hc2290576, 32'h42c42da2, 32'h42882d8c, 32'hc2846170, 32'h42a2e6dd};
test_weights[13568:13575] = '{32'h42b51312, 32'hc249df63, 32'hc27d11d8, 32'h42382f6d, 32'hc1bb412f, 32'h41fa9a16, 32'hc29c14cd, 32'hc1f3b8a2};
test_bias[1696:1696] = '{32'hc28a98ca};
test_output[1696:1696] = '{32'hc48901c5};
test_input[13576:13583] = '{32'h41d4dfed, 32'hc2b9971f, 32'hc2aa59ad, 32'hc0e5f08a, 32'h42ae7b62, 32'h42af96e4, 32'hc2646db7, 32'hc0765714};
test_weights[13576:13583] = '{32'hc23271be, 32'hc2390240, 32'h42803289, 32'hc2bdecf1, 32'h42c28c83, 32'hc2c0d6a6, 32'h427080b8, 32'hc2a5af29};
test_bias[1697:1697] = '{32'h424cffc8};
test_output[1697:1697] = '{32'hc59354ed};
test_input[13584:13591] = '{32'hc2a23cff, 32'h42aee256, 32'hc2828353, 32'h42439ccb, 32'h427c92ec, 32'hc2787482, 32'h428f2e74, 32'hc1b2d3fa};
test_weights[13584:13591] = '{32'h4163aa3e, 32'h4287c758, 32'h42a8b7f8, 32'h428d9988, 32'hc0549e58, 32'h42304ab8, 32'h4127b1b8, 32'hc216dbd7};
test_bias[1698:1698] = '{32'hc2698e05};
test_output[1698:1698] = '{32'h44a5e552};
test_input[13592:13599] = '{32'h3d7b7c0b, 32'hc2b067aa, 32'h429023b9, 32'h428bb7a1, 32'hc2109c51, 32'h420cfdb3, 32'h425aafc5, 32'h42667666};
test_weights[13592:13599] = '{32'hc2bfb2e2, 32'hc17b8cfb, 32'hc18c27c8, 32'h42b68ecc, 32'h424c3591, 32'hc298e938, 32'h417cca20, 32'h42206cfa};
test_bias[1699:1699] = '{32'hc2b4fbf5};
test_output[1699:1699] = '{32'h459d7273};
test_input[13600:13607] = '{32'hc28491db, 32'h42421402, 32'h426beca2, 32'h428c6722, 32'hc25f2c3b, 32'h42c7689e, 32'h424ce1ee, 32'h422428fc};
test_weights[13600:13607] = '{32'h42a35caa, 32'hc2c65222, 32'h413245a4, 32'h3f833763, 32'hc23e5c18, 32'h42ab4daa, 32'hc218a5d4, 32'hc0e1841f};
test_bias[1700:1700] = '{32'hc28cdfd8};
test_output[1700:1700] = '{32'hc419e666};
test_input[13608:13615] = '{32'hc25105cc, 32'hc213110d, 32'h427e92d0, 32'h42b9a5ff, 32'h422b1966, 32'hc2353d1b, 32'hc289d7e7, 32'hc2891968};
test_weights[13608:13615] = '{32'hc12ea0ac, 32'h4293870e, 32'hbfdc11cf, 32'hc162f41f, 32'hc279ac4c, 32'h42464828, 32'h42983bbb, 32'h42a428c2};
test_bias[1701:1701] = '{32'h41c9afcf};
test_output[1701:1701] = '{32'hc6970655};
test_input[13616:13623] = '{32'h4236b2ac, 32'h42b1224c, 32'hc2444270, 32'h4215c2e1, 32'h41a3127a, 32'hc2760b3b, 32'h4257b7e3, 32'h42b7ddda};
test_weights[13616:13623] = '{32'hc2b0e883, 32'hc24480fc, 32'h425ade29, 32'h42828138, 32'hc2b1a05c, 32'h417e211b, 32'hc1ac6903, 32'hc294667e};
test_bias[1702:1702] = '{32'h42b69a00};
test_output[1702:1702] = '{32'hc696e0d6};
test_input[13624:13631] = '{32'h424c42c4, 32'hc2af2b1c, 32'h40e21a07, 32'h4292f5c4, 32'hc2b5b453, 32'h40be6c59, 32'h4222aa77, 32'hc1f3e721};
test_weights[13624:13631] = '{32'hc210d2c4, 32'h426bd36d, 32'hc2944fe7, 32'hc297e9cc, 32'h42457725, 32'hc1caada8, 32'hc2b2e014, 32'hc265a096};
test_bias[1703:1703] = '{32'hc2855494};
test_output[1703:1703] = '{32'hc699f647};
test_input[13632:13639] = '{32'h4158d42f, 32'hc1296e27, 32'hc2aa2219, 32'hc0c5097b, 32'hc1b189d2, 32'hc19cd520, 32'hc28f546f, 32'h40ad63cb};
test_weights[13632:13639] = '{32'h42035a16, 32'hc27ef372, 32'h42487f0d, 32'hc266f13a, 32'hc2ae203a, 32'hc1e93858, 32'h41135494, 32'hc28e90b7};
test_bias[1704:1704] = '{32'h42c4b6eb};
test_output[1704:1704] = '{32'hc49a1266};
test_input[13640:13647] = '{32'hc21af752, 32'h421de1ee, 32'h424c270d, 32'hc21a04fe, 32'h425335a2, 32'hc22b8cad, 32'h425bbe12, 32'h4275d9ca};
test_weights[13640:13647] = '{32'hc169ec27, 32'h4290e462, 32'h42b734c8, 32'h4180ceb8, 32'hc1502e64, 32'h41de97be, 32'hc2c74f8a, 32'hc2340702};
test_bias[1705:1705] = '{32'h42935f82};
test_output[1705:1705] = '{32'hc5206542};
test_input[13648:13655] = '{32'h41d2f341, 32'hc1d4ff72, 32'h42b0cf6c, 32'h42b2b3a3, 32'h41967a09, 32'h41badb12, 32'hc1d46a39, 32'hbe8ada82};
test_weights[13648:13655] = '{32'h4206e003, 32'hc12cf4f6, 32'h4273dcf4, 32'hc2c5460d, 32'h415dccad, 32'hc2119a1b, 32'hc189bd9c, 32'h419f87a9};
test_bias[1706:1706] = '{32'hc1357c14};
test_output[1706:1706] = '{32'hc515bb76};
test_input[13656:13663] = '{32'hc229dacd, 32'h41e37e38, 32'hc1da1cad, 32'h429f5cb6, 32'h42ba0257, 32'h41da7a41, 32'h4263a484, 32'h4276215f};
test_weights[13656:13663] = '{32'hc209382a, 32'h42195090, 32'h41b00a7e, 32'h427e97cd, 32'hc2bac46d, 32'hc26f1814, 32'hc154cb7c, 32'hc23078a3};
test_bias[1707:1707] = '{32'hc1fb8871};
test_output[1707:1707] = '{32'hc5d49212};
test_input[13664:13671] = '{32'h427f738e, 32'hc18b6863, 32'hc25dfa5f, 32'h41be5a8d, 32'h424401fb, 32'h424b0b7d, 32'h4285f88c, 32'h427f70b8};
test_weights[13664:13671] = '{32'h4242fc96, 32'hc2208e7d, 32'h42a11648, 32'hc2a06a57, 32'hc2c647d1, 32'h42a71bdc, 32'h42c3ab3c, 32'h4286cf53};
test_bias[1708:1708] = '{32'h42344f66};
test_output[1708:1708] = '{32'h45f14556};
test_input[13672:13679] = '{32'h421e4902, 32'h419277a1, 32'h41e69719, 32'hc02267c7, 32'h427d9759, 32'h41d5dbe9, 32'h4207e46e, 32'h4193bddf};
test_weights[13672:13679] = '{32'h422a42fe, 32'h42a761a3, 32'hc1cf5afe, 32'h420afc04, 32'h411cc122, 32'hc1f319fe, 32'h40d0074d, 32'h420a2c61};
test_bias[1709:1709] = '{32'h42109c7c};
test_output[1709:1709] = '{32'h4540d12a};
test_input[13680:13687] = '{32'hc1f14f86, 32'hc281bbe3, 32'h429a15cb, 32'h42b549f7, 32'hc27cdd2b, 32'hc27e0275, 32'h41b7f64b, 32'hc22ea251};
test_weights[13680:13687] = '{32'h41873342, 32'hc0f20e51, 32'hc221c428, 32'h4257c750, 32'hc28df1a4, 32'hc2681448, 32'h42b9fd9b, 32'h4278f579};
test_bias[1710:1710] = '{32'hc1098f36};
test_output[1710:1710] = '{32'h4611e9ed};
test_input[13688:13695] = '{32'hc0d9bded, 32'hc18b1b0b, 32'hc1f14b8c, 32'hc21dc5da, 32'h3fec3fad, 32'h41a8f583, 32'hc0b1bbc9, 32'h415c8589};
test_weights[13688:13695] = '{32'hc201aabe, 32'h41b295b6, 32'hc29f19e0, 32'h42b3f838, 32'h42ac4ea6, 32'h41f424c0, 32'hc20b594d, 32'hc20a0fec};
test_bias[1711:1711] = '{32'hc2a249c4};
test_output[1711:1711] = '{32'hc45b52d6};
test_input[13696:13703] = '{32'hc252e390, 32'h4227271a, 32'h424d2e53, 32'hc23f466d, 32'hc206dc60, 32'h41c19961, 32'hbf1941fc, 32'h425c148b};
test_weights[13696:13703] = '{32'hc015cd30, 32'h42ad71e4, 32'h3faf6867, 32'hc193c6cb, 32'hc2670cbe, 32'hc17366c3, 32'h421eb850, 32'hc0b49d32};
test_bias[1712:1712] = '{32'h4295958e};
test_output[1712:1712] = '{32'h45bc2673};
test_input[13704:13711] = '{32'hc27675cd, 32'h42c25850, 32'h4151e948, 32'hc25507bc, 32'hc184125f, 32'hc232133d, 32'hc2163fda, 32'hc108a9d8};
test_weights[13704:13711] = '{32'hc292b3a7, 32'hc27b267c, 32'hc1b1c06b, 32'h42ae851f, 32'h4193db2d, 32'h41831179, 32'h4202b052, 32'h41695703};
test_bias[1713:1713] = '{32'h42affbbb};
test_output[1713:1713] = '{32'hc609cb1b};
test_input[13712:13719] = '{32'hc282a07c, 32'hc2a357e8, 32'h41cc7017, 32'hc2985c34, 32'hc22597e8, 32'h41a632fc, 32'hc2796573, 32'hc27b11ec};
test_weights[13712:13719] = '{32'hc1991db8, 32'hc252170c, 32'hc1d15f7c, 32'hc2b2f418, 32'hc0ee296a, 32'hc297abc2, 32'h41b09a06, 32'hc25c93dc};
test_bias[1714:1714] = '{32'h426d88d3};
test_output[1714:1714] = '{32'h46445089};
test_input[13720:13727] = '{32'h41e482e2, 32'h42558ac0, 32'h425ce36d, 32'hc2774759, 32'h4249474e, 32'hc2ba2512, 32'hc0b4d463, 32'h42a05b42};
test_weights[13720:13727] = '{32'h42a4dbcb, 32'h421b4fb3, 32'hc293e283, 32'hc288b49c, 32'hc189096d, 32'h420e676e, 32'hc1a740c9, 32'h4190380a};
test_bias[1715:1715] = '{32'hc10bc1c9};
test_output[1715:1715] = '{32'h44f3a098};
test_input[13728:13735] = '{32'h41f1ff3f, 32'hc20463cc, 32'h42837b10, 32'h4012a72f, 32'h42a624f6, 32'hc212f724, 32'hc29a4e8e, 32'hc1c9f50f};
test_weights[13728:13735] = '{32'hc186680b, 32'hc1e66f35, 32'h426d7b1d, 32'hc2b46909, 32'h42931052, 32'hc2843028, 32'hc2a67ae3, 32'h416a3545};
test_bias[1716:1716] = '{32'h426b000c};
test_output[1716:1716] = '{32'h4692cb85};
test_input[13736:13743] = '{32'h41cb4f8c, 32'hc1c7ab4b, 32'hc29384fe, 32'h4214bcfa, 32'hc1f4b1a6, 32'h429ef66c, 32'h4230856b, 32'h4114253d};
test_weights[13736:13743] = '{32'hc225990e, 32'hc1488395, 32'h42987209, 32'hc2551ff0, 32'hc21a6c56, 32'h41db1c40, 32'h4140bdbf, 32'h423d08be};
test_bias[1717:1717] = '{32'hc1c16855};
test_output[1717:1717] = '{32'hc57c8040};
test_input[13744:13751] = '{32'hc178c9fc, 32'h41810782, 32'hc21e355e, 32'hc21cc820, 32'hc2a63882, 32'hc227e183, 32'h41cf0722, 32'hc29bc61f};
test_weights[13744:13751] = '{32'hc2b31d11, 32'hc28e79bd, 32'h42371a30, 32'hc2b446b4, 32'h41bfb8e5, 32'h424582ab, 32'hc1690cc4, 32'hc1e02ebb};
test_bias[1718:1718] = '{32'hc196697a};
test_output[1718:1718] = '{32'hc39b9c51};
test_input[13752:13759] = '{32'hc1e32d5f, 32'h42877214, 32'hc1d33780, 32'hc2b4b48e, 32'h4165a414, 32'hc1d856bd, 32'h4249fdb4, 32'hc28f438b};
test_weights[13752:13759] = '{32'hc2a9debd, 32'h4270e37d, 32'hc29ba30a, 32'h42c1ada0, 32'hc2644394, 32'h42a2fb30, 32'hc28ec1ee, 32'hc24ffb34};
test_bias[1719:1719] = '{32'h40d53bc7};
test_output[1719:1719] = '{32'hc541ccb0};
test_input[13760:13767] = '{32'h42027eb4, 32'hc2661077, 32'hc1de4247, 32'hc2a695ff, 32'hc0894f3c, 32'h422c6062, 32'hc2ab28a4, 32'h42874dc7};
test_weights[13760:13767] = '{32'h41b3cd9b, 32'hc2c08ad3, 32'h3fe16cea, 32'h42b9821f, 32'h4112df2a, 32'hc0c7d3d0, 32'hc19a2a3e, 32'h42673bee};
test_bias[1720:1720] = '{32'h421b9682};
test_output[1720:1720] = '{32'h456ca1a0};
test_input[13768:13775] = '{32'hc1d70acf, 32'h42916c29, 32'h42adbe8e, 32'hc2919b29, 32'hc2785315, 32'hc0596371, 32'h426cc90e, 32'h4280938b};
test_weights[13768:13775] = '{32'h42870475, 32'h4200232d, 32'hc2ad1a40, 32'h422a92fc, 32'h42ba9dc2, 32'hc226cf9d, 32'h40189a67, 32'hc28aa69e};
test_bias[1721:1721] = '{32'hbf2ff741};
test_output[1721:1721] = '{32'hc69cd87a};
test_input[13776:13783] = '{32'h41c45289, 32'hc2987f2e, 32'hc2c3487e, 32'h41903469, 32'hc2596191, 32'hc2789d26, 32'hc2ac7e75, 32'hc111da70};
test_weights[13776:13783] = '{32'h42881144, 32'hc1d8c476, 32'h42c23c5f, 32'hc2901691, 32'h42ab3792, 32'h42a29dfd, 32'hc214e28e, 32'h3fbf9b89};
test_bias[1722:1722] = '{32'h42863963};
test_output[1722:1722] = '{32'hc652c08d};
test_input[13784:13791] = '{32'hc0bb1488, 32'h42926890, 32'hc2968dfb, 32'h416a6894, 32'hc1166ae4, 32'hc2b55d7d, 32'hc19d4574, 32'h42b230c9};
test_weights[13784:13791] = '{32'h4276e8b2, 32'hc2c7fae7, 32'hc2282382, 32'h42c1141a, 32'hc1e4f797, 32'h4239db3c, 32'hc2623c77, 32'h42afd91d};
test_bias[1723:1723] = '{32'h41a15496};
test_output[1723:1723] = '{32'h44efe98e};
test_input[13792:13799] = '{32'hc2077f06, 32'hc1a3bc94, 32'hc208264c, 32'hc19558f5, 32'h406177c5, 32'hc11166ec, 32'hc2752356, 32'h412d2e99};
test_weights[13792:13799] = '{32'hc2845116, 32'hc2181251, 32'hc28f3af5, 32'hc283f71d, 32'hc2937c96, 32'hc1b3beae, 32'h42082407, 32'h42c02743};
test_bias[1724:1724] = '{32'hc238911c};
test_output[1724:1724] = '{32'h45ad2724};
test_input[13800:13807] = '{32'h4297f249, 32'hc2389e7e, 32'hc24dbb7b, 32'hc297add6, 32'h42c7b9a8, 32'hc17df999, 32'h42895f0b, 32'hc23d844b};
test_weights[13800:13807] = '{32'h414ad90d, 32'h403b6e52, 32'h422814d8, 32'h41298ad2, 32'h42306e3d, 32'hc2a9a674, 32'hc256775f, 32'hc0852a5b};
test_bias[1725:1725] = '{32'hc220cab1};
test_output[1725:1725] = '{32'h42b136b1};
test_input[13808:13815] = '{32'hc02d115e, 32'hc2b7a882, 32'h42b45046, 32'hc0589a62, 32'hc2120edd, 32'h4253f47e, 32'hc2b31e4a, 32'h423019da};
test_weights[13808:13815] = '{32'hc27466ff, 32'h402a8555, 32'hc24663b0, 32'h41d07bed, 32'hc1f82a86, 32'h42b1ac58, 32'hc1d52059, 32'h41209d3b};
test_bias[1726:1726] = '{32'hc240792e};
test_output[1726:1726] = '{32'h4578c9f7};
test_input[13816:13823] = '{32'h40e66afc, 32'hc2213722, 32'hc206d678, 32'h4057377c, 32'hc23a6667, 32'h428a43a8, 32'hc05cc905, 32'h426af193};
test_weights[13816:13823] = '{32'h412fd396, 32'h42b82ac1, 32'h4170c1cd, 32'hc2360918, 32'h41f007d2, 32'hc2499ced, 32'h4235d75b, 32'hc2c6852e};
test_bias[1727:1727] = '{32'h41afccb5};
test_output[1727:1727] = '{32'hc66c9072};
test_input[13824:13831] = '{32'hc257d73e, 32'hc1320a3a, 32'h427cf3df, 32'h42b2a9cb, 32'hc28d4dc3, 32'hc26a9ad0, 32'hc245b02c, 32'hc1203024};
test_weights[13824:13831] = '{32'hc114a4d8, 32'hc1698376, 32'h42bb0679, 32'h428755ab, 32'h421ee89e, 32'h41cdc94c, 32'h42b0abc8, 32'h429d2939};
test_bias[1728:1728] = '{32'h42900b39};
test_output[1728:1728] = '{32'h4549a2ce};
test_input[13832:13839] = '{32'hc2b70be4, 32'hc2749952, 32'hc20937dc, 32'hc2815aae, 32'hc246acbd, 32'hc293f40f, 32'h40b7cfd1, 32'hc0e847fd};
test_weights[13832:13839] = '{32'h42ac8181, 32'h426d0e6c, 32'h42b947ee, 32'h429a4977, 32'hc2227fd9, 32'h42891f0d, 32'h419123b4, 32'hc1bac860};
test_bias[1729:1729] = '{32'h3ec30879};
test_output[1729:1729] = '{32'hc6af8325};
test_input[13840:13847] = '{32'hc26d6a2f, 32'h4162e2bd, 32'hc23477fa, 32'hc2b1acf2, 32'hc2b2d5e6, 32'hc28e1da1, 32'hc231217c, 32'h42424de5};
test_weights[13840:13847] = '{32'h424c7d86, 32'h426b4e47, 32'hc2ab8adf, 32'hc2a62f08, 32'h40524617, 32'hc29c7a1a, 32'hc2c2891e, 32'hc1868450};
test_bias[1730:1730] = '{32'h42587c37};
test_output[1730:1730] = '{32'h468b8b37};
test_input[13848:13855] = '{32'hc26d60f6, 32'h42b530d4, 32'hc2669ef3, 32'h4254e4c5, 32'hc228b3eb, 32'h425888d3, 32'hc244470e, 32'hc2ac902b};
test_weights[13848:13855] = '{32'hc2a8d15f, 32'hc2655230, 32'h412422da, 32'h3fe4d7ab, 32'h4262dcf1, 32'hc2586524, 32'h41b82691, 32'hc1463248};
test_bias[1731:1731] = '{32'hc2816366};
test_output[1731:1731] = '{32'hc5bf7792};
test_input[13856:13863] = '{32'h3f825d88, 32'h419feb41, 32'hc21dd5d4, 32'hc2b55ee5, 32'h4285c556, 32'hc26771ea, 32'hc26ed919, 32'hc1fcd9be};
test_weights[13856:13863] = '{32'hc2834074, 32'h42000ef8, 32'h42171abb, 32'hc23b4898, 32'hc2c31568, 32'h4199915d, 32'h420520f5, 32'h410d5a7c};
test_bias[1732:1732] = '{32'h42a89643};
test_output[1732:1732] = '{32'hc5cac4e7};
test_input[13864:13871] = '{32'hc2968d31, 32'h42c56686, 32'h416f1ccb, 32'h42bd15a4, 32'h41b0062c, 32'hc29be0c7, 32'hc2ad0546, 32'h42496caf};
test_weights[13864:13871] = '{32'hc08448ba, 32'hc1bdb0b6, 32'hc2a2d1ae, 32'hc0be5085, 32'hc25c9659, 32'hc233d0ee, 32'hc2150d9e, 32'hc22e6f1f};
test_bias[1733:1733] = '{32'h429f59ac};
test_output[1733:1733] = '{32'hc3cd300e};
test_input[13872:13879] = '{32'h428bcb11, 32'h41a465f3, 32'h429e8104, 32'h4258bb1e, 32'hc229282f, 32'hc0940a96, 32'hc1c935e3, 32'h424d87f3};
test_weights[13872:13879] = '{32'hc22a6818, 32'h42a3abcc, 32'hc296d3e1, 32'hc275bd25, 32'hc18752ff, 32'h41cedb1c, 32'hc213b36a, 32'hbe87de70};
test_bias[1734:1734] = '{32'hc2a72498};
test_output[1734:1734] = '{32'hc60f58b0};
test_input[13880:13887] = '{32'hc21c31f4, 32'h42b0f387, 32'hc2088ddc, 32'hc2a7e277, 32'hc1d0769b, 32'h42a39e0b, 32'h42b23648, 32'h4281916b};
test_weights[13880:13887] = '{32'hc283576a, 32'h42b40935, 32'hc209a35e, 32'h426e15ba, 32'hc278eaec, 32'hc1952376, 32'h426e74a3, 32'h41a0d5b0};
test_bias[1735:1735] = '{32'hc2b9d629};
test_output[1735:1735] = '{32'h46503431};
test_input[13888:13895] = '{32'hc127206b, 32'hc2567bb8, 32'hc29ac18a, 32'h42544cd7, 32'hc2b9550f, 32'h42abc65b, 32'hc26517ad, 32'h42223846};
test_weights[13888:13895] = '{32'hc29b0815, 32'hc27832f2, 32'h4185628a, 32'hc296df09, 32'h428eb205, 32'h4126c2ae, 32'h40a7caeb, 32'hc2ac8cbb};
test_bias[1736:1736] = '{32'hc2347c5a};
test_output[1736:1736] = '{32'hc62776c8};
test_input[13896:13903] = '{32'hc17c4327, 32'hc182510b, 32'hc1c05c03, 32'hc0f7f9b6, 32'hc27655a4, 32'h429f9af5, 32'hc0dd0882, 32'hc282759c};
test_weights[13896:13903] = '{32'h41a338a9, 32'h42b49726, 32'h42591610, 32'h422d97cb, 32'hc24f0ecf, 32'h42a61f4e, 32'h40ccae3f, 32'h428bb394};
test_bias[1737:1737] = '{32'h42bb715f};
test_output[1737:1737] = '{32'h44ea7782};
test_input[13904:13911] = '{32'h415b79ab, 32'hc1f95001, 32'hc2bc426e, 32'hc1dae463, 32'hc2b3cf5c, 32'h42bdf61e, 32'h42b2840e, 32'h41a442ec};
test_weights[13904:13911] = '{32'h419170b5, 32'hc27d3328, 32'hc2aafe7a, 32'h402a22cb, 32'hc2376241, 32'h424e3a69, 32'h41836c27, 32'hc286818a};
test_bias[1738:1738] = '{32'hc216fa98};
test_output[1738:1738] = '{32'h46967f0d};
test_input[13912:13919] = '{32'hc18399a1, 32'h4231cb15, 32'h41308b9b, 32'h41877862, 32'h427a4143, 32'hc1f4ed8a, 32'hc219694f, 32'h4289cc1b};
test_weights[13912:13919] = '{32'h42a47590, 32'hc2241cb9, 32'hc21431a8, 32'h418fada1, 32'h41d48134, 32'hc28a012b, 32'hc1666085, 32'hc221d57f};
test_bias[1739:1739] = '{32'hc21b8cc3};
test_output[1739:1739] = '{32'hc4de96d5};
test_input[13920:13927] = '{32'h3f82552c, 32'h4138a571, 32'h424a30cd, 32'hc261cf2c, 32'hc2566ea3, 32'h4262c564, 32'hc1e40afa, 32'hc1a91de4};
test_weights[13920:13927] = '{32'hc2b9a73d, 32'hc23f08ca, 32'hc2bef7c9, 32'h41ecddba, 32'h427fae5d, 32'h40857bc4, 32'hc0a7e3ef, 32'h42c2117c};
test_bias[1740:1740] = '{32'hc11cb38a};
test_output[1740:1740] = '{32'hc63f5517};
test_input[13928:13935] = '{32'h424f234d, 32'hc28d2561, 32'h42b91f00, 32'h42028139, 32'hc25e886e, 32'h429f3d69, 32'hc1b48d6c, 32'h429cac5b};
test_weights[13928:13935] = '{32'h42c01429, 32'h42972ef9, 32'h42b74292, 32'hc19d89ed, 32'hc16a9144, 32'h42401483, 32'h4279b397, 32'h423da96d};
test_bias[1741:1741] = '{32'hc2ae9e88};
test_output[1741:1741] = '{32'h465ffa59};
test_input[13936:13943] = '{32'h4172fcb4, 32'hc2b1a581, 32'hc10e8b92, 32'h41e7291a, 32'hc2a723d6, 32'hc19d788e, 32'hc26b4918, 32'hc1b82212};
test_weights[13936:13943] = '{32'hc21c8653, 32'h4287701b, 32'h40b98f18, 32'hc226acfa, 32'h421ae245, 32'hc2759000, 32'h41d237bf, 32'h422e5056};
test_bias[1742:1742] = '{32'hc2b463da};
test_output[1742:1742] = '{32'hc643cd7d};
test_input[13944:13951] = '{32'h42b30b74, 32'hc1d23879, 32'hc2a4580d, 32'h42740cda, 32'h427cf9f5, 32'hc29fc000, 32'hc1f675ee, 32'h42466948};
test_weights[13944:13951] = '{32'h425088f1, 32'h42676ee6, 32'h3ffe19b9, 32'hc1a862f6, 32'h40051f30, 32'h41ba0250, 32'hc18b7e7b, 32'h426dca5b};
test_bias[1743:1743] = '{32'hc2621cd1};
test_output[1743:1743] = '{32'h4554b36c};
test_input[13952:13959] = '{32'hc0382e13, 32'h4255a269, 32'h41bc3a1d, 32'h42c784ff, 32'h42ad6616, 32'h42a0fffe, 32'h40a7184f, 32'hc1d8b4bf};
test_weights[13952:13959] = '{32'h4259add2, 32'h4297ffa6, 32'hc1f43600, 32'hc27a94fe, 32'h429776ed, 32'h40e836c3, 32'hc28c141c, 32'hc25d899f};
test_bias[1744:1744] = '{32'hc1e71696};
test_output[1744:1744] = '{32'h45a23375};
test_input[13960:13967] = '{32'hc2a16892, 32'hc1d886c9, 32'hc0e2bd54, 32'h4282b7d7, 32'hc1a061a4, 32'h41d09ff7, 32'hc213f27a, 32'hc26d21c6};
test_weights[13960:13967] = '{32'hc1971e4b, 32'hc2718137, 32'hc2aa778b, 32'h4251cd9e, 32'hc2b7ba97, 32'hc2590355, 32'hc19c4538, 32'hc2aa7f5f};
test_bias[1745:1745] = '{32'hc29a8ffe};
test_output[1745:1745] = '{32'h4650122b};
test_input[13968:13975] = '{32'hc264c1f8, 32'hc2709449, 32'hc28ef931, 32'hc27dc5d7, 32'hc2bdba18, 32'hc29a61c9, 32'h42ae3fe5, 32'h41d94ee7};
test_weights[13968:13975] = '{32'hc2942eca, 32'hc13f6806, 32'hc170b708, 32'hc239d47f, 32'hc2a02394, 32'hc105e262, 32'h423a1f0c, 32'hc29fb247};
test_bias[1746:1746] = '{32'hc224bd2c};
test_output[1746:1746] = '{32'h4694f217};
test_input[13976:13983] = '{32'hc230ac57, 32'hc186df6f, 32'hc00f960d, 32'h4171bec0, 32'hc22bccde, 32'hc133bca0, 32'h42c208b5, 32'h422ae015};
test_weights[13976:13983] = '{32'h4063c42d, 32'hc177e301, 32'h42be12fb, 32'h41eb0b49, 32'h42786573, 32'hbe5cdc13, 32'hc21190a1, 32'hc1da46ea};
test_bias[1747:1747] = '{32'hc2c2a739};
test_output[1747:1747] = '{32'hc5de9bfc};
test_input[13984:13991] = '{32'h4201f00e, 32'h428cbb3f, 32'hc28cb423, 32'h42ac55c1, 32'hc123367c, 32'hc20a72c5, 32'h428bfab8, 32'hc27400d5};
test_weights[13984:13991] = '{32'h4294ef4b, 32'hc1ed89dc, 32'h4272bcfb, 32'hc2c4e420, 32'hc0e10191, 32'hc2549fb3, 32'h41ed190d, 32'h41d9bbd7};
test_bias[1748:1748] = '{32'h41b4cbe9};
test_output[1748:1748] = '{32'hc61d6894};
test_input[13992:13999] = '{32'h41b14a78, 32'h42a5e16e, 32'hc2998840, 32'hc2945895, 32'hc2133bb0, 32'h4269c080, 32'h42b6cc23, 32'h429b4516};
test_weights[13992:13999] = '{32'h422194d1, 32'hc058ccc7, 32'h42382562, 32'h42ba389c, 32'h4298cee9, 32'hc137cfde, 32'h4291aa90, 32'h41225355};
test_bias[1749:1749] = '{32'h42704557};
test_output[1749:1749] = '{32'hc5b56970};
test_input[14000:14007] = '{32'hc220f97b, 32'h42aa368c, 32'h4221ed49, 32'h42638a1d, 32'hc1c731c8, 32'h421264fc, 32'hc29083b6, 32'h42b5c966};
test_weights[14000:14007] = '{32'hc2a3d7ce, 32'h42ad8745, 32'h41a9d8ae, 32'hc1ee4629, 32'h427e53d6, 32'h4233f298, 32'h42c05fcf, 32'hc22b11d4};
test_bias[1750:1750] = '{32'hc288465b};
test_output[1750:1750] = '{32'hc47906fc};
test_input[14008:14015] = '{32'hc1826b4e, 32'hbf2ad654, 32'h4158e7d7, 32'hc23db273, 32'hc2a8d4f0, 32'hc2adda34, 32'hc27c3206, 32'hc1b788e1};
test_weights[14008:14015] = '{32'hc239276c, 32'h4222632b, 32'h4189f353, 32'hc25ab1e1, 32'h419e67cb, 32'hc26daac2, 32'hc2ab8e79, 32'h427b4229};
test_bias[1751:1751] = '{32'h423a5ab9};
test_output[1751:1751] = '{32'h462cd507};
test_input[14016:14023] = '{32'hc19df959, 32'h42346b58, 32'hc2673c09, 32'h429a6ec9, 32'h422686cf, 32'hc0ca2fa3, 32'h41f1e767, 32'h421e54c3};
test_weights[14016:14023] = '{32'hc29378f0, 32'hc28a45c3, 32'hc2bec401, 32'hc21193c5, 32'hc2b3ac35, 32'hc1ce4c96, 32'h40414cb1, 32'h4177fd4e};
test_bias[1752:1752] = '{32'hc2b013ff};
test_output[1752:1752] = '{32'hc4efdd76};
test_input[14024:14031] = '{32'hc2aaf695, 32'h428f8779, 32'h4290923e, 32'h42700e38, 32'h426cb4ac, 32'h423aa1a0, 32'hc14bb93c, 32'h418981e7};
test_weights[14024:14031] = '{32'h429314d9, 32'h4159038f, 32'hc135caa7, 32'h41b09c3b, 32'h410f3dc2, 32'h4240c606, 32'h423af37c, 32'h421a3ede};
test_bias[1753:1753] = '{32'h424d08b8};
test_output[1753:1753] = '{32'hc4ef02ab};
test_input[14032:14039] = '{32'hc1ce3197, 32'h4272a80e, 32'hc20cbaa1, 32'hc2adf705, 32'h41a85667, 32'hbe98c742, 32'h41d33576, 32'h425d7335};
test_weights[14032:14039] = '{32'h42b4da5f, 32'h41dbbedb, 32'hc2a4f523, 32'h417360cf, 32'h41a1f490, 32'h4298d348, 32'hc279ac48, 32'h4282796e};
test_bias[1754:1754] = '{32'hc29a237c};
test_output[1754:1754] = '{32'h454843f7};
test_input[14040:14047] = '{32'hc25b671a, 32'h42895244, 32'h4100fa4a, 32'h40e0c6c6, 32'hc23ac429, 32'h421b7568, 32'h4233bc14, 32'hc23e863a};
test_weights[14040:14047] = '{32'h41691567, 32'hc297e8db, 32'hc15f3fcd, 32'hc2a1395d, 32'hc2533bce, 32'h42193030, 32'hc1edfba6, 32'h4200bd9e};
test_bias[1755:1755] = '{32'h4200b735};
test_output[1755:1755] = '{32'hc5ae4243};
test_input[14048:14055] = '{32'h42bbe9e7, 32'h42482f92, 32'hc2451e26, 32'hc25b8d59, 32'h42b92f79, 32'h4151b15a, 32'hc2a16bf2, 32'hc2074b34};
test_weights[14048:14055] = '{32'hc29050cd, 32'hc192c731, 32'hc25642c0, 32'h42956038, 32'hc25c83cf, 32'hc1bd9515, 32'hc26d85a8, 32'h428798cb};
test_bias[1756:1756] = '{32'hbfd1d219};
test_output[1756:1756] = '{32'hc63cac07};
test_input[14056:14063] = '{32'h3eab7f95, 32'hc126a4d9, 32'hc27878cd, 32'h4255f5a0, 32'h41e84bf8, 32'h42891aee, 32'hc2535d03, 32'hc2b7403e};
test_weights[14056:14063] = '{32'hc03aef96, 32'h425042b1, 32'h424ab75c, 32'h427b2e8a, 32'hc23975a6, 32'hc22f0979, 32'hc25af264, 32'hc26a1eee};
test_bias[1757:1757] = '{32'h42913f45};
test_output[1757:1757] = '{32'h456414b0};
test_input[14064:14071] = '{32'hc238aede, 32'h42a36102, 32'hc288e564, 32'hc2aa1d78, 32'h42987076, 32'h428310ea, 32'h42bbe83b, 32'hc2bc4449};
test_weights[14064:14071] = '{32'h42319dae, 32'hc217cfaa, 32'hc0fd07a7, 32'h4275f913, 32'hc244be62, 32'h4163e3ed, 32'hc2637bb7, 32'hc2780157};
test_bias[1758:1758] = '{32'h4146a390};
test_output[1758:1758] = '{32'hc63dd6c2};
test_input[14072:14079] = '{32'h42634764, 32'hc27e4c04, 32'hc18277af, 32'hc2c4c028, 32'h4277b1d4, 32'h42c00295, 32'h41b863b0, 32'h424e2bda};
test_weights[14072:14079] = '{32'h425c222b, 32'h42bfcc51, 32'hc1f837d7, 32'hc20e560b, 32'h4258a03c, 32'h42194bb6, 32'h41ee686a, 32'hc2aa2bd3};
test_bias[1759:1759] = '{32'hc202bcf7};
test_output[1759:1759] = '{32'h458792e6};
test_input[14080:14087] = '{32'hc12789df, 32'h424e4041, 32'hc28599bb, 32'hc1241070, 32'hbfd159e0, 32'h41c18e48, 32'h42098e10, 32'hc26becd8};
test_weights[14080:14087] = '{32'hc2358340, 32'hc287d0ca, 32'hc2b18464, 32'hc2b05703, 32'hc25adc6a, 32'h4142b35d, 32'h428817dc, 32'h42c3617f};
test_bias[1760:1760] = '{32'hc0d68be9};
test_output[1760:1760] = '{32'h443e8b03};
test_input[14088:14095] = '{32'hc15004b7, 32'hc06e912f, 32'h40faf95b, 32'hc1460aeb, 32'hc1217625, 32'h42aa89f3, 32'hc2a542d0, 32'h42247395};
test_weights[14088:14095] = '{32'hc28ef2f1, 32'hc28a6684, 32'h41d80606, 32'hc27b9741, 32'h42943991, 32'hc29845f9, 32'h427d323f, 32'h4290083e};
test_bias[1761:1761] = '{32'h41e08576};
test_output[1761:1761] = '{32'hc5e440bc};
test_input[14096:14103] = '{32'hbf552a23, 32'h41ec8ef3, 32'hc104aca4, 32'h429cea46, 32'hc105d4c5, 32'hc28e9ccb, 32'h42912b4e, 32'h41a7734c};
test_weights[14096:14103] = '{32'h40ba30a2, 32'h426b8f6c, 32'hc162a879, 32'h422b9e68, 32'hc1bf9c46, 32'hc2869650, 32'hbf633da0, 32'hc1e49fda};
test_bias[1762:1762] = '{32'h42808258};
test_output[1762:1762] = '{32'h46165283};
test_input[14104:14111] = '{32'h42971015, 32'hc2a7cfcb, 32'hc2662e2a, 32'hc2abcc0d, 32'hc21673e3, 32'h42c119c0, 32'hc2a754c6, 32'hc1ef1b8d};
test_weights[14104:14111] = '{32'hc21e05f5, 32'hc11899e3, 32'h4227962b, 32'h425b8bca, 32'hc259aaf8, 32'hc297e37f, 32'h4287c1d6, 32'hc29f4b8b};
test_bias[1763:1763] = '{32'h41b021fa};
test_output[1763:1763] = '{32'hc68b9ef8};
test_input[14112:14119] = '{32'hc1908803, 32'h42b1019b, 32'h41d25618, 32'h41eeb812, 32'hc24ef796, 32'hc203406b, 32'hc2b1d2ae, 32'h41b77790};
test_weights[14112:14119] = '{32'hbe9ecfca, 32'hbf98cb68, 32'h42349ff2, 32'hc23149d9, 32'h4232182a, 32'hc2b66f66, 32'hc1e1c53c, 32'hc19f44f0};
test_bias[1764:1764] = '{32'hc1fe599b};
test_output[1764:1764] = '{32'h451aadaa};
test_input[14120:14127] = '{32'h42c238f5, 32'h419bb507, 32'h427ceaf3, 32'hc180ec8e, 32'h42788c3a, 32'hc1c76985, 32'hc22a698b, 32'h421493a7};
test_weights[14120:14127] = '{32'h407714d1, 32'hc21df80e, 32'h426ac367, 32'h42288bcb, 32'hc1ff7770, 32'hc2a30ff3, 32'hc2522857, 32'h4214c8d4};
test_bias[1765:1765] = '{32'h42295f61};
test_output[1765:1765] = '{32'h45c66462};
test_input[14128:14135] = '{32'hc1a60ea1, 32'hc2651f8e, 32'h3fe06bee, 32'h42ad72df, 32'hc211e63c, 32'h41be8d0f, 32'hc27bdd5c, 32'hc19b230f};
test_weights[14128:14135] = '{32'hc2848ca9, 32'h4273f14f, 32'h42b60de8, 32'h422f64c5, 32'hc2a29ba9, 32'h426ca557, 32'h4181a167, 32'h425856fe};
test_bias[1766:1766] = '{32'h42a093bd};
test_output[1766:1766] = '{32'h45843497};
test_input[14136:14143] = '{32'hc23d9fb4, 32'h42c16a24, 32'h419c2992, 32'hc216e47e, 32'hc2ac15f7, 32'hc2b75124, 32'hc25b63a0, 32'h4254ccf1};
test_weights[14136:14143] = '{32'hc072a2d8, 32'h3f949fdb, 32'hc224b394, 32'h41c97554, 32'h42775d55, 32'hc2b5e1cf, 32'h424eeb0b, 32'hc214b3d6};
test_bias[1767:1767] = '{32'h423cfb26};
test_output[1767:1767] = '{32'hc548ee5f};
test_input[14144:14151] = '{32'h41e56b92, 32'hc270b715, 32'h42992c24, 32'hc28a30d5, 32'h42229d3b, 32'h42a53477, 32'hc2996b8e, 32'h4026750d};
test_weights[14144:14151] = '{32'h3f66def3, 32'hc28ffe2c, 32'h429a2400, 32'hc2bb0587, 32'hc2801d51, 32'h413c9139, 32'hbfb3b3fb, 32'hc2a57790};
test_bias[1768:1768] = '{32'hc1c24c01};
test_output[1768:1768] = '{32'h4669bf26};
test_input[14152:14159] = '{32'h4283fbf7, 32'h423bef38, 32'hc0516034, 32'hc275f58e, 32'h42c79f0a, 32'h42879383, 32'h422e6fd4, 32'hc242861b};
test_weights[14152:14159] = '{32'hc298ab43, 32'h41e78b46, 32'h42978b05, 32'hc08991bc, 32'h4226bd59, 32'h42a0b069, 32'h419420fe, 32'h42c2c52e};
test_bias[1769:1769] = '{32'hc2ada336};
test_output[1769:1769] = '{32'h44f151d3};
test_input[14160:14167] = '{32'hc22a8122, 32'h4051cdd7, 32'h42849b50, 32'hc2848144, 32'h3f6871ae, 32'hc2825aa0, 32'h420dd183, 32'hc225ce78};
test_weights[14160:14167] = '{32'hc234a9a2, 32'hc29685bc, 32'hc2612a0e, 32'h426cbc76, 32'h4285d04d, 32'h40e54806, 32'hc2bada98, 32'hc27cdda2};
test_bias[1770:1770] = '{32'h4214a9f4};
test_output[1770:1770] = '{32'hc5dbdf71};
test_input[14168:14175] = '{32'h42a46f66, 32'hc2700fc6, 32'hc28ca65d, 32'hc29e4b7c, 32'h425b68af, 32'h42ab8778, 32'h42b7576d, 32'h42c2fe4f};
test_weights[14168:14175] = '{32'h42c452c4, 32'hc284c16f, 32'h41bf0fe8, 32'h4283ad08, 32'h41e99d3c, 32'hc27ce3fe, 32'hc18cbf01, 32'h420add55};
test_bias[1771:1771] = '{32'h418fa71f};
test_output[1771:1771] = '{32'h4543d3d8};
test_input[14176:14183] = '{32'h422bc68a, 32'h423e0a86, 32'h42895ada, 32'h4185e753, 32'hc2834bf1, 32'h4095cf90, 32'h428f0bb0, 32'hc1ec9109};
test_weights[14176:14183] = '{32'hc0eafc10, 32'hc0abc5e8, 32'hc0be93db, 32'h42a8b950, 32'hc2c3a2c9, 32'h42899168, 32'hc1b95c83, 32'h41ecb5f7};
test_bias[1772:1772] = '{32'hc2453834};
test_output[1772:1772] = '{32'h458f9650};
test_input[14184:14191] = '{32'h4220f599, 32'h425ad3f0, 32'hc2101e9a, 32'h42af8627, 32'h41621675, 32'hc2c3dd8d, 32'h42a0264e, 32'hc1402a29};
test_weights[14184:14191] = '{32'h41c2272a, 32'hc2c4eaab, 32'h42b4dbb1, 32'h42182b64, 32'hc19a94aa, 32'h420941d8, 32'hc0aa6804, 32'h405a4379};
test_bias[1773:1773] = '{32'hc21bea65};
test_output[1773:1773] = '{32'hc6045484};
test_input[14192:14199] = '{32'hc121ecd7, 32'hc2984385, 32'hc2254b35, 32'hc2bd30b0, 32'h4288a5ce, 32'hc294ba52, 32'h42ab8067, 32'hc12be508};
test_weights[14192:14199] = '{32'h42c1d84e, 32'hc2654096, 32'h41ca5a1d, 32'h42a51dd3, 32'hc26bb03a, 32'hc0820d4a, 32'hc24c7bb6, 32'hc1f65f26};
test_bias[1774:1774] = '{32'h42a78273};
test_output[1774:1774] = '{32'hc64db3e2};
test_input[14200:14207] = '{32'hc24cec74, 32'h3f546af8, 32'hc2b88e4c, 32'hc238f27e, 32'h41ca22c7, 32'hc26bbf44, 32'hc28fa6a4, 32'h42b603fa};
test_weights[14200:14207] = '{32'hc28f508b, 32'h42271899, 32'h4112a6fa, 32'h4285a632, 32'hc279283c, 32'h420b8f07, 32'hc29d68bb, 32'h412909a9};
test_bias[1775:1775] = '{32'h41c0b4da};
test_output[1775:1775] = '{32'h452da981};
test_input[14208:14215] = '{32'hc28611bf, 32'h42ba7201, 32'h423abffe, 32'hc19fd844, 32'hc1f818e3, 32'h423697a5, 32'hc1896823, 32'hc2398acb};
test_weights[14208:14215] = '{32'h426f5231, 32'hc06351ba, 32'hc18e89a8, 32'hc26c3cfe, 32'h42bc691e, 32'hc2a4cab8, 32'hc28ceccc, 32'h42bc4fbf};
test_bias[1776:1776] = '{32'h42866baa};
test_output[1776:1776] = '{32'hc657195c};
test_input[14216:14223] = '{32'hc017110a, 32'h429fb884, 32'hc2be7a4b, 32'h422b278a, 32'hc2ba4799, 32'hc21de515, 32'hc20eeac0, 32'h420ae5ee};
test_weights[14216:14223] = '{32'hc209f962, 32'hc2753cf3, 32'hc2b73d07, 32'h428b106b, 32'h4253b7f8, 32'hc0a1125c, 32'hc1abe99d, 32'hc0d1cfa9};
test_bias[1777:1777] = '{32'h426ee1c5};
test_output[1777:1777] = '{32'h452c2c51};
test_input[14224:14231] = '{32'h420f04e2, 32'h42afb0e2, 32'h418af247, 32'h41e8f9b3, 32'h4124aab3, 32'h4155aabb, 32'hc29ce988, 32'h40e9cc87};
test_weights[14224:14231] = '{32'hc261b37b, 32'hc207bddb, 32'h429bf525, 32'hc01f9b00, 32'hc2919d4a, 32'hc2b8a21e, 32'h402475aa, 32'h40819b7d};
test_bias[1778:1778] = '{32'h4242b1ed};
test_output[1778:1778] = '{32'hc5b5f230};
test_input[14232:14239] = '{32'hc12fbc06, 32'h4135a453, 32'hc23e247d, 32'hc29ca532, 32'h419b5265, 32'hc2ac46a6, 32'h424916df, 32'hc127cb5a};
test_weights[14232:14239] = '{32'h423fbd0a, 32'hc28b0b21, 32'hc133032b, 32'h4293873c, 32'h4295b38d, 32'hc20a163e, 32'h427d6c90, 32'hc27377fa};
test_bias[1779:1779] = '{32'h42afadaf};
test_output[1779:1779] = '{32'h44de1961};
test_input[14240:14247] = '{32'hc2bed418, 32'h42c23c05, 32'h41cfe787, 32'h422a24d1, 32'h42b8ab68, 32'h42b3375c, 32'hc2356fb6, 32'h4298d623};
test_weights[14240:14247] = '{32'h41ed2b85, 32'hc2b1bfc8, 32'hc230ce7e, 32'hc29baffe, 32'hc2c1f5e6, 32'hc25d6cd9, 32'h42966c35, 32'h427d9939};
test_bias[1780:1780] = '{32'hc1958001};
test_output[1780:1780] = '{32'hc6de0849};
test_input[14248:14255] = '{32'hc2bbeb56, 32'hc28277f9, 32'h410c5298, 32'hc1abc9a1, 32'h42a2cb4f, 32'h41f1157e, 32'hc20d9a97, 32'hc1c456bb};
test_weights[14248:14255] = '{32'hc278986b, 32'hc1bf73a2, 32'h429d4089, 32'h422f5250, 32'hc1a443bf, 32'h41b5e2ae, 32'hc2a49842, 32'hc2869cea};
test_bias[1781:1781] = '{32'hc1d53c55};
test_output[1781:1781] = '{32'h462735c1};
test_input[14256:14263] = '{32'hc29f87f0, 32'hbc1b1cdb, 32'hc1cfa983, 32'h41f9c5bc, 32'hc29fbff0, 32'hc1a8a9db, 32'h42a67d69, 32'h428eb53c};
test_weights[14256:14263] = '{32'h424ba468, 32'hc1f675f7, 32'h41897140, 32'h429ad72f, 32'h42936896, 32'h424e7f10, 32'h3e6d3ff3, 32'h422179dd};
test_bias[1782:1782] = '{32'h42552a9c};
test_output[1782:1782] = '{32'hc5befeac};
test_input[14264:14271] = '{32'hc2994169, 32'h3fa340a5, 32'hc299b9da, 32'h4165f784, 32'hc24c56b1, 32'h3e8edf76, 32'h42a05eb5, 32'h4262c727};
test_weights[14264:14271] = '{32'hc24087a9, 32'h4121f6b9, 32'h42bf98cb, 32'hc1a301fb, 32'h428c9ebf, 32'hc1dfd863, 32'h41ba4de6, 32'hc2bb8ea3};
test_bias[1783:1783] = '{32'hc19cc9e0};
test_output[1783:1783] = '{32'hc62c3e49};
test_input[14272:14279] = '{32'h4219ae8e, 32'hc2bed9e5, 32'h42066a4d, 32'h42beeec8, 32'hc1fa1b8b, 32'h419d3bf2, 32'hc076d101, 32'hc21d4e57};
test_weights[14272:14279] = '{32'hc116191e, 32'h40063f1f, 32'hc0ba7703, 32'hc28e8ca9, 32'hc26ebc62, 32'h40ca2941, 32'h3e726520, 32'hc19401d9};
test_bias[1784:1784] = '{32'h42b0a185};
test_output[1784:1784] = '{32'hc5949d5e};
test_input[14280:14287] = '{32'hc21ac91d, 32'h41f2d5e5, 32'h4193e3c3, 32'hbd436d35, 32'h426d28d2, 32'h42b5f175, 32'hc28cc003, 32'h3f0fffd6};
test_weights[14280:14287] = '{32'hc2b2b1ca, 32'h416bd68f, 32'hc203230e, 32'hc2af2939, 32'hc2a1fb29, 32'h41e0c391, 32'h41f24c58, 32'hc14685f9};
test_bias[1785:1785] = '{32'h41684f09};
test_output[1785:1785] = '{32'hc4855fd5};
test_input[14288:14295] = '{32'h4233bff1, 32'h42449fca, 32'hc0b98630, 32'hc2b12a03, 32'h41b2b56e, 32'hc2c06324, 32'hc2703e68, 32'h41c89c80};
test_weights[14288:14295] = '{32'hc28b71a3, 32'h42832785, 32'h42283291, 32'h42a8146f, 32'hc290aff6, 32'hc2455710, 32'hc1b2d2ab, 32'hbfafa396};
test_bias[1786:1786] = '{32'hc2bd08ea};
test_output[1786:1786] = '{32'hc54b68ef};
test_input[14296:14303] = '{32'hc2c4aaf0, 32'h429efa1a, 32'h421ff6c0, 32'hc108e7f7, 32'hc26ec569, 32'h42acc94b, 32'hc1d64a0c, 32'h42215c54};
test_weights[14296:14303] = '{32'h4298dc4e, 32'hc2b5eae2, 32'h42982d00, 32'h4105fc31, 32'h42b0cbd6, 32'hc25ea246, 32'hc22b71e2, 32'hc28ebe27};
test_bias[1787:1787] = '{32'h42140395};
test_output[1787:1787] = '{32'hc6b803ef};
test_input[14304:14311] = '{32'h424e4cfd, 32'hc2556113, 32'hc21c91ce, 32'hc2649fda, 32'h42c4fd20, 32'h42a88f17, 32'hc2a1145e, 32'h4268916e};
test_weights[14304:14311] = '{32'hc2a57cbd, 32'h42b3114c, 32'hc28df80b, 32'h41df1638, 32'h42be019d, 32'h42baf6c2, 32'h423b1fc9, 32'h41775866};
test_bias[1788:1788] = '{32'h42a3e59a};
test_output[1788:1788] = '{32'h45cdef2e};
test_input[14312:14319] = '{32'hc20b7b5c, 32'hc2bb967b, 32'hc2c1552f, 32'h421d8aee, 32'h428c1898, 32'h425f796f, 32'h428185aa, 32'h42820591};
test_weights[14312:14319] = '{32'h41cc6ad9, 32'h42b03435, 32'h428e441d, 32'hc20553c2, 32'hc2c10d19, 32'hc28b69bf, 32'hc2b512a4, 32'hc2a8db43};
test_bias[1789:1789] = '{32'h40b84b92};
test_output[1789:1789] = '{32'hc719b179};
test_input[14320:14327] = '{32'hc20d252b, 32'hc232d1e5, 32'h404ebbca, 32'hc2bb5d2e, 32'h41c3c5a6, 32'hc188d2b2, 32'h41d0b785, 32'h4209e3b9};
test_weights[14320:14327] = '{32'hc2243d68, 32'hc2490c1a, 32'hc2a35296, 32'hc1d56d62, 32'h42666ee2, 32'hc102ec9b, 32'hc27106d9, 32'hc113d34a};
test_bias[1790:1790] = '{32'h42b9d714};
test_output[1790:1790] = '{32'h45b19afe};
test_input[14328:14335] = '{32'h419e6606, 32'h42bb48e2, 32'hc247fd87, 32'hc1f66704, 32'hc15bc674, 32'hc2a8af03, 32'h4215aa7f, 32'hc1c40861};
test_weights[14328:14335] = '{32'hc2878d5a, 32'h40062ec9, 32'h42a044a5, 32'h429a9060, 32'hc202c27f, 32'hc245ea73, 32'h4254270f, 32'hc2b7944f};
test_bias[1791:1791] = '{32'hc28cee22};
test_output[1791:1791] = '{32'h449c9fad};
test_input[14336:14343] = '{32'hc1f7c192, 32'h427c1a07, 32'hc2740888, 32'h41b8cd7c, 32'hc28fc39e, 32'h42362264, 32'h42b92d48, 32'h428b5b07};
test_weights[14336:14343] = '{32'hc19efd55, 32'h42887e96, 32'h4095d259, 32'h400576b1, 32'hc2423ca8, 32'hc2a55109, 32'hc1d4556c, 32'hc0bb060a};
test_bias[1792:1792] = '{32'h423c276d};
test_output[1792:1792] = '{32'h44c68f9e};
test_input[14344:14351] = '{32'h42794e82, 32'hc1b40550, 32'h3fc58097, 32'hc2b67ab3, 32'h42ab3ff6, 32'h416f8a3a, 32'hc2357ebe, 32'h4287c934};
test_weights[14344:14351] = '{32'hc2ba7a60, 32'h40bdea3c, 32'h4162d36f, 32'h415c2d70, 32'h429fc925, 32'hc2b8d71c, 32'hc2adb02d, 32'h424375e4};
test_bias[1793:1793] = '{32'hc10e1fca};
test_output[1793:1793] = '{32'h45acbe9c};
test_input[14352:14359] = '{32'hc1408b73, 32'hc25a2f62, 32'h4248f97b, 32'hc28dc412, 32'h42217660, 32'hc2445c86, 32'h42a05459, 32'h420cc8d4};
test_weights[14352:14359] = '{32'h4216b05d, 32'h40aefc34, 32'hc25e51bc, 32'h4295e5ac, 32'hc2793a30, 32'h4252a315, 32'hc22d5906, 32'hc2c4f99a};
test_bias[1794:1794] = '{32'hbf6b6d75};
test_output[1794:1794] = '{32'hc6a3447a};
test_input[14360:14367] = '{32'hc2b2ddbf, 32'h41bdf782, 32'hc18bd71f, 32'hc20a7b21, 32'h41f0554c, 32'h42a8c4e5, 32'h4297815c, 32'hc201a49e};
test_weights[14360:14367] = '{32'h42c40006, 32'h413b2738, 32'hc2c55640, 32'h41ed176c, 32'hc192e7ff, 32'hc25e1852, 32'h4248e840, 32'hc213269c};
test_bias[1795:1795] = '{32'h4153a34f};
test_output[1795:1795] = '{32'hc5fa7514};
test_input[14368:14375] = '{32'h40b7fa83, 32'h421397c0, 32'hc279caaa, 32'hc2b91a27, 32'h42a1d100, 32'hbfa15184, 32'h41379231, 32'hc2af53b3};
test_weights[14368:14375] = '{32'hc2b5661f, 32'h42818bfd, 32'h424e70ba, 32'h41f8a8a0, 32'h421f0b37, 32'hc29a3a29, 32'hc2abb9ab, 32'hc02c481e};
test_bias[1796:1796] = '{32'hc19a54fd};
test_output[1796:1796] = '{32'hc4d2aae4};
test_input[14376:14383] = '{32'hc2c35f47, 32'h4232eba4, 32'hc2a38ea4, 32'hc0b29058, 32'hc1007760, 32'h42b3be1b, 32'h4284c99a, 32'hc2b88b23};
test_weights[14376:14383] = '{32'h4136f730, 32'h425f6292, 32'h42241708, 32'h42c7fe5e, 32'h42130b07, 32'hc2c3cae0, 32'h4207dbc9, 32'h422f68f8};
test_bias[1797:1797] = '{32'h40f5ebac};
test_output[1797:1797] = '{32'hc65182a8};
test_input[14384:14391] = '{32'hc1fc1f9a, 32'h4206fd4a, 32'h4209eaba, 32'h419e1531, 32'h42811159, 32'hc293e43e, 32'h42341274, 32'h42942215};
test_weights[14384:14391] = '{32'hc1c60ff5, 32'h429fa9c4, 32'hc1d279ae, 32'h42273b3c, 32'hc1f6990f, 32'hc2a6900d, 32'h42988fd4, 32'h3fff0a22};
test_bias[1798:1798] = '{32'hc23b3e42};
test_output[1798:1798] = '{32'h462d64db};
test_input[14392:14399] = '{32'h429b74eb, 32'h424a107f, 32'h41b59a2e, 32'hc2aeed50, 32'h42824c09, 32'h41c8ef0f, 32'h417454a4, 32'hbf2017f0};
test_weights[14392:14399] = '{32'hc0bb61a0, 32'h42307181, 32'hbe610d6a, 32'hc204c406, 32'h413f1f26, 32'h42a0f36e, 32'hc21cd154, 32'h40f0b6ed};
test_bias[1799:1799] = '{32'hc031da67};
test_output[1799:1799] = '{32'h45d68440};
test_input[14400:14407] = '{32'hc2b70a76, 32'h4210cbfd, 32'h42c1d377, 32'h42ba7da0, 32'h428783dd, 32'hc2a07082, 32'h42c00795, 32'h4274fc54};
test_weights[14400:14407] = '{32'h4098da85, 32'h429ff74b, 32'h4207b067, 32'hc27d0384, 32'h421e84dd, 32'h426c7ac0, 32'h41a09747, 32'hc1ebdc3b};
test_bias[1800:1800] = '{32'hc2aa4978};
test_output[1800:1800] = '{32'hc507d3e6};
test_input[14408:14415] = '{32'h42abd6ba, 32'hc12b35df, 32'h4190e82f, 32'hc19e804a, 32'h425e2348, 32'hc27e5e9c, 32'h42801a0a, 32'hc20f2f34};
test_weights[14408:14415] = '{32'hc25ab41e, 32'h428c8817, 32'hc09612e6, 32'h41835c05, 32'hc1831ff9, 32'h41b09da6, 32'hc297d38d, 32'hc12d7bc3};
test_bias[1801:1801] = '{32'hc1f911c5};
test_output[1801:1801] = '{32'hc6461d73};
test_input[14416:14423] = '{32'h4281d734, 32'h41623192, 32'h40241884, 32'hc29542df, 32'h42b0068d, 32'h40a3c693, 32'h42b63898, 32'h4228bf6f};
test_weights[14416:14423] = '{32'h42a1d631, 32'h4060282a, 32'hc2af6809, 32'h42a5d483, 32'hc1cb0694, 32'h4296b5df, 32'hc2ba9a68, 32'hc2b0729c};
test_bias[1802:1802] = '{32'h42c67959};
test_output[1802:1802] = '{32'hc66ba5df};
test_input[14424:14431] = '{32'h42c31926, 32'hbe087207, 32'hc15c16bf, 32'h425de41d, 32'hc1b15b6a, 32'h41a156e1, 32'h42a8c5ea, 32'hc293cf03};
test_weights[14424:14431] = '{32'h42a8e98b, 32'hc26e972f, 32'h421aeb0a, 32'h42bff015, 32'hc1b8b188, 32'hbf38e33b, 32'h4232d50e, 32'h428eaad4};
test_bias[1803:1803] = '{32'hc2508b0e};
test_output[1803:1803] = '{32'h463b3e01};
test_input[14432:14439] = '{32'h42bd8734, 32'hc26c4357, 32'hc1fa1be9, 32'hc1132a8b, 32'h426b8b6d, 32'h41d7145d, 32'hc2327edc, 32'h42bf7db7};
test_weights[14432:14439] = '{32'h42a2a14a, 32'h42ba281d, 32'h42bc633a, 32'hc1022886, 32'h421070c8, 32'h42b52f13, 32'h40145f69, 32'hc26fe3db};
test_bias[1804:1804] = '{32'h429d9f33};
test_output[1804:1804] = '{32'hc4e95a0d};
test_input[14440:14447] = '{32'h42221e16, 32'hc0bf00a0, 32'hc2a3ff80, 32'hc2368500, 32'h42b7df50, 32'hc2815256, 32'h423eac56, 32'hc0753afb};
test_weights[14440:14447] = '{32'h41af3a7d, 32'h41d736fb, 32'hc0c1e334, 32'h4288a7f1, 32'h4127f294, 32'hc180db14, 32'h429ec54c, 32'hc249304f};
test_bias[1805:1805] = '{32'hc2298426};
test_output[1805:1805] = '{32'h457cf39b};
test_input[14448:14455] = '{32'h40df0ffe, 32'h428721e2, 32'hc13ee2d4, 32'hc20ee680, 32'h4268513a, 32'hc2381c15, 32'hc23b1b1d, 32'h42b93aa1};
test_weights[14448:14455] = '{32'hc265bbff, 32'hc0f1b8f2, 32'h414664ec, 32'h42a00871, 32'h4178e714, 32'hc2c2e2e0, 32'h42a88764, 32'h42a17f08};
test_bias[1806:1806] = '{32'h4299d7a9};
test_output[1806:1806] = '{32'h459ee891};
test_input[14456:14463] = '{32'hc279975f, 32'h4270f787, 32'h4299c5db, 32'h42b141e6, 32'hc2a4d34b, 32'h42151ee6, 32'hc25a8f1a, 32'h42908e06};
test_weights[14456:14463] = '{32'hc1f7cb83, 32'hc2c3bc6d, 32'h420c4bf9, 32'hc245be4e, 32'h4209cba3, 32'h42ae33ea, 32'hc2c3290f, 32'hc25db63a};
test_bias[1807:1807] = '{32'h4246ffad};
test_output[1807:1807] = '{32'hc5718427};
test_input[14464:14471] = '{32'h4190148f, 32'hc2835348, 32'hc1556af4, 32'hc1f48b03, 32'h4247dac3, 32'h41c231f1, 32'h421eff45, 32'h4289005b};
test_weights[14464:14471] = '{32'hc29af788, 32'h424dca00, 32'hc2872226, 32'h4286a9f1, 32'h4262ee5c, 32'hc165fc51, 32'hc244c0dd, 32'h4225f8e0};
test_bias[1808:1808] = '{32'h42a98ef7};
test_output[1808:1808] = '{32'hc51a90f1};
test_input[14472:14479] = '{32'h41f1b417, 32'hc2b7787c, 32'h3fd6fe39, 32'hc183a62d, 32'hc25c3292, 32'h42877f7a, 32'h4265146c, 32'h41d1b4d4};
test_weights[14472:14479] = '{32'hc214a3e2, 32'hc229a74d, 32'hc23afc36, 32'h42b89b8d, 32'h42ba836e, 32'h4287b105, 32'hc2901428, 32'hc2aebfc4};
test_bias[1809:1809] = '{32'hc2c6370b};
test_output[1809:1809] = '{32'hc5b7ce75};
test_input[14480:14487] = '{32'h42311978, 32'hc241681b, 32'h418a0f7a, 32'hc282a146, 32'hc0eff54a, 32'h423cda77, 32'h420ae228, 32'h42c33ab7};
test_weights[14480:14487] = '{32'hc2b8cc24, 32'h4228dd39, 32'hc285c7df, 32'hc2ae3bdd, 32'h413a43db, 32'h427f6eb5, 32'hc01b6738, 32'h422d5947};
test_bias[1810:1810] = '{32'hc20100e9};
test_output[1810:1810] = '{32'h45aa27b7};
test_input[14488:14495] = '{32'hc2a47e32, 32'hc0490593, 32'h42bc3488, 32'hc2a61569, 32'hc2a876be, 32'hc2b4c759, 32'hbfe7feb1, 32'h42a453a6};
test_weights[14488:14495] = '{32'hc167f391, 32'hc2b75957, 32'hc1fdcc30, 32'hc2b9628e, 32'h41b9a5ce, 32'hc20b9f6b, 32'h42851522, 32'hc2bc8fbd};
test_bias[1811:1811] = '{32'hc22fe0da};
test_output[1811:1811] = '{32'hc4019527};
test_input[14496:14503] = '{32'hbf835921, 32'hc2666c05, 32'hc22e0c28, 32'hc13c1016, 32'h41a49165, 32'h422aaf0d, 32'h42805e2b, 32'hc1ed5f26};
test_weights[14496:14503] = '{32'h42767cc6, 32'hc2b575c0, 32'hc1814169, 32'hc283cd47, 32'hc1a810f4, 32'h42538fbe, 32'hc2c37e61, 32'hc2b391ed};
test_bias[1812:1812] = '{32'h42047782};
test_output[1812:1812] = '{32'h4598c850};
test_input[14504:14511] = '{32'h419a1463, 32'h40f4e33c, 32'hc2b3203a, 32'h428433df, 32'hc23216b1, 32'hc1bf98dc, 32'h4076f32b, 32'h41c8d1aa};
test_weights[14504:14511] = '{32'h42b748df, 32'h42916f6c, 32'hc214366c, 32'h41df4e58, 32'h4191b11a, 32'hc0f51d23, 32'hc2ad3184, 32'hc22bfd9e};
test_bias[1813:1813] = '{32'hc2768b49};
test_output[1813:1813] = '{32'h45a835c6};
test_input[14512:14519] = '{32'h41005a08, 32'hc2834aa7, 32'hc2b251d7, 32'h42003cfa, 32'h40f7b740, 32'hc2933849, 32'h42401ebe, 32'h4286f5c0};
test_weights[14512:14519] = '{32'hc2858ab4, 32'h420f769e, 32'hc197a307, 32'h42c2564d, 32'h427a6ab0, 32'h4293d35b, 32'h4296e0bc, 32'h42a601fd};
test_bias[1814:1814] = '{32'hc27f1b85};
test_output[1814:1814] = '{32'h45bf3d48};
test_input[14520:14527] = '{32'hc1d55386, 32'h42944953, 32'h42b7a7b0, 32'hc181d21a, 32'hc2460331, 32'hc25167e3, 32'h42b5ea9e, 32'hc268ff2f};
test_weights[14520:14527] = '{32'hc2160d24, 32'h42725622, 32'h428526c0, 32'hc248430b, 32'h4171e255, 32'h3ff42039, 32'hc25854c1, 32'h427a5168};
test_bias[1815:1815] = '{32'h41cff75a};
test_output[1815:1815] = '{32'h453d76cf};
test_input[14528:14535] = '{32'h41ae9aeb, 32'h42a4f194, 32'hc2aebc3d, 32'hc290bc77, 32'h42b7603d, 32'h42553e88, 32'hc27bf654, 32'hc2af4214};
test_weights[14528:14535] = '{32'h42a9c2be, 32'hc2597026, 32'h422e4d75, 32'hc18818bc, 32'h425829ad, 32'h4209eb46, 32'h4262b5b2, 32'h422f949c};
test_bias[1816:1816] = '{32'h423ca792};
test_output[1816:1816] = '{32'hc5b4b7b8};
test_input[14536:14543] = '{32'h4242c3cd, 32'h42691f71, 32'hc239f890, 32'hc2a2644c, 32'hc2bf1472, 32'hc06d5d42, 32'hc2b71bb3, 32'h41d2a222};
test_weights[14536:14543] = '{32'hc1f7e671, 32'hc19a155f, 32'h41bfbaf9, 32'hc2b01017, 32'h4244fdf4, 32'h42170046, 32'h429506b7, 32'hc19df6c0};
test_bias[1817:1817] = '{32'hc25ef72a};
test_output[1817:1817] = '{32'hc60a2241};
test_input[14544:14551] = '{32'h42060bcb, 32'hc1b28080, 32'hc28a41ac, 32'hc2b2c662, 32'h4290d71a, 32'hc233b57d, 32'h42534b84, 32'hc290186c};
test_weights[14544:14551] = '{32'h420f354d, 32'hc18f229f, 32'hc29ffad9, 32'hc259fcdb, 32'h422d0d17, 32'hc2873182, 32'hc20e717f, 32'h42af03ab};
test_bias[1818:1818] = '{32'h42283bfd};
test_output[1818:1818] = '{32'h461ca8d3};
test_input[14552:14559] = '{32'h424e4ef3, 32'h4288a171, 32'hc16d3aee, 32'hc246fc0c, 32'hc28a3bfe, 32'h423fbfcb, 32'hc223173c, 32'h426ec92c};
test_weights[14552:14559] = '{32'hc21b4a69, 32'h41aaa3b4, 32'h41b2c5e8, 32'hc1ad8547, 32'hc1040f34, 32'hc2b220cd, 32'h42aff788, 32'hc1f190bd};
test_bias[1819:1819] = '{32'h425692c9};
test_output[1819:1819] = '{32'hc60a0338};
test_input[14560:14567] = '{32'hc0b11ade, 32'hc2900ba5, 32'hc281f8bd, 32'h42a5c794, 32'h428a0873, 32'h42ab6e07, 32'h4215d911, 32'h42b832d0};
test_weights[14560:14567] = '{32'h41237025, 32'hc1e58207, 32'hc2644033, 32'h421b736a, 32'h42b4738c, 32'hc0a32514, 32'h42ad4f2c, 32'h422f2676};
test_bias[1820:1820] = '{32'hc20f25af};
test_output[1820:1820] = '{32'h46aba937};
test_input[14568:14575] = '{32'hc1dadbc6, 32'h428aa042, 32'h40e1e139, 32'h42910192, 32'h4201370f, 32'hc1369538, 32'h420d1b13, 32'hc259b43f};
test_weights[14568:14575] = '{32'h41ea4654, 32'h4256b6bd, 32'hc27ee566, 32'h41dee25d, 32'h41f93171, 32'h42b4b792, 32'h41f6c904, 32'hc2bd555c};
test_bias[1821:1821] = '{32'hc2574398};
test_output[1821:1821] = '{32'h46266dec};
test_input[14576:14583] = '{32'h42629add, 32'h40309bfb, 32'hc1c62f2b, 32'hc1360e1e, 32'h421c8ab6, 32'hc249008b, 32'hc17bc3b2, 32'hc28b54d4};
test_weights[14576:14583] = '{32'h420e4ea9, 32'h422e63f1, 32'hbee16345, 32'h42a84a55, 32'h429426cb, 32'h414710d5, 32'hc15b7ea2, 32'h42b13c3f};
test_bias[1822:1822] = '{32'h4298c90b};
test_output[1822:1822] = '{32'hc517251d};
test_input[14584:14591] = '{32'h40a58fb5, 32'hc09934f8, 32'h4236cc54, 32'h42850f0a, 32'h41cbdd25, 32'h419113aa, 32'hc251f02b, 32'h42b56f2c};
test_weights[14584:14591] = '{32'h42031587, 32'h41b05a59, 32'hc1449875, 32'hc19c95e5, 32'h426ba7f1, 32'hc2770e8b, 32'h425ddd47, 32'h4180961d};
test_bias[1823:1823] = '{32'h428228b2};
test_output[1823:1823] = '{32'hc52f6607};
test_input[14592:14599] = '{32'hc2ae1c56, 32'hc276deaa, 32'h414fef13, 32'h42c3c1dd, 32'hc1959576, 32'hc2a4a720, 32'hc1a7be6d, 32'hc16ff180};
test_weights[14592:14599] = '{32'h4290ac1f, 32'h41e85139, 32'hc26368b7, 32'h4213bd47, 32'h428db315, 32'hc14d92e4, 32'hc29ba30a, 32'hc2c3af79};
test_bias[1824:1824] = '{32'hc2392af4};
test_output[1824:1824] = '{32'hc517b81b};
test_input[14600:14607] = '{32'hc2639813, 32'h4295cc11, 32'h42a35d32, 32'hc20d7386, 32'h42ab08d6, 32'hc295587d, 32'h41a3f31b, 32'h425cf8a5};
test_weights[14600:14607] = '{32'hc170bbdf, 32'hc2642887, 32'hc2b789f5, 32'hc2905b95, 32'h4119fd9d, 32'hc1801370, 32'hc267df68, 32'h4005707c};
test_bias[1825:1825] = '{32'hc1a873c8};
test_output[1825:1825] = '{32'hc5e85724};
test_input[14608:14615] = '{32'h425f5754, 32'h429e5a62, 32'h41f4dd3f, 32'h42c3ef38, 32'hbf1d26c5, 32'hc2b10dfa, 32'hc1fa067d, 32'h41171486};
test_weights[14608:14615] = '{32'hc04e7afd, 32'hc2380cfd, 32'hc25c500c, 32'hc2813512, 32'hc24ce275, 32'hc209d165, 32'h429ce48d, 32'hc145adb3};
test_bias[1826:1826] = '{32'h429a8694};
test_output[1826:1826] = '{32'hc62fbe85};
test_input[14616:14623] = '{32'hc165c9ff, 32'hc2148268, 32'h423dfd5d, 32'h42c2feed, 32'h425bf086, 32'hbfc6ca68, 32'h429659ac, 32'hc1c52279};
test_weights[14616:14623] = '{32'hc2432d9d, 32'hc256923f, 32'hc256906d, 32'hc1d0ca04, 32'hc19eda14, 32'h42716fa2, 32'h428cd94d, 32'hc2b0d089};
test_bias[1827:1827] = '{32'hc1cc8860};
test_output[1827:1827] = '{32'h4571596c};
test_input[14624:14631] = '{32'h4244cf1c, 32'hc1ce2355, 32'h429eba4f, 32'h41ba5a49, 32'h42a4b018, 32'h412454ca, 32'hc297627b, 32'hc29121a9};
test_weights[14624:14631] = '{32'hc2c3067a, 32'hc28c5b3e, 32'h427ab003, 32'h42c3ad3e, 32'h42445315, 32'h426a406f, 32'h42ba00e3, 32'hc243823b};
test_bias[1828:1828] = '{32'hc2c1eaf9};
test_output[1828:1828] = '{32'h45a625f2};
test_input[14632:14639] = '{32'hbf9ba4f1, 32'hc2246a1c, 32'h42c57094, 32'h40e4b87c, 32'h426573e5, 32'h4288be4a, 32'hc13546e4, 32'hc2aa450d};
test_weights[14632:14639] = '{32'h42853c41, 32'h42b00c94, 32'h41bf5825, 32'h42ac5187, 32'h429dc351, 32'hc107920d, 32'h42a2837e, 32'h41f41a25};
test_bias[1829:1829] = '{32'hc1cf330f};
test_output[1829:1829] = '{32'hc3a063ae};
test_input[14640:14647] = '{32'h42bb9ff8, 32'hc2b4165f, 32'h418f6d33, 32'hc06ae465, 32'h41ca3a65, 32'h42ae53c3, 32'hc1a9d55f, 32'h4254e427};
test_weights[14640:14647] = '{32'h429e8806, 32'hc25ee539, 32'hc2351dea, 32'hc208ef4f, 32'h40c5ac35, 32'h42b81ba3, 32'hc28dd4f9, 32'h4237cb84};
test_bias[1830:1830] = '{32'hc21916e9};
test_output[1830:1830] = '{32'h46ba6864};
test_input[14648:14655] = '{32'h42bf0e21, 32'hc2a9235e, 32'hc299f9b3, 32'hc29a1492, 32'h4277edd7, 32'hc26c1836, 32'h42670f28, 32'h42c26d50};
test_weights[14648:14655] = '{32'hbfa52f87, 32'h42193301, 32'h42374801, 32'h4288d9dd, 32'hc232a293, 32'hc15c0ea3, 32'hc29ea022, 32'hc16b5ab5};
test_bias[1831:1831] = '{32'h426363c4};
test_output[1831:1831] = '{32'hc69cd082};
test_input[14656:14663] = '{32'h429aa887, 32'h4236018b, 32'h42b3c9b7, 32'hc2556758, 32'h4246476f, 32'hc00c0e17, 32'hc0411d03, 32'hc2b6d7b3};
test_weights[14656:14663] = '{32'hc176211c, 32'hc26a84eb, 32'h40626f0e, 32'h4281e75b, 32'hc1d6e386, 32'hc2702014, 32'h41d2aa52, 32'hc2c4cb61};
test_bias[1832:1832] = '{32'h420ab1a5};
test_output[1832:1832] = '{32'h443a8c22};
test_input[14664:14671] = '{32'hc206f3d6, 32'hc2c53d21, 32'h4214a286, 32'hc29e94fd, 32'hc21fd03b, 32'h4299a237, 32'h42a7f773, 32'hc2105b3b};
test_weights[14664:14671] = '{32'hc05ccb87, 32'hc127b32a, 32'h42898568, 32'hc194a270, 32'hc2a29349, 32'h41583870, 32'h42448008, 32'h42831cb5};
test_bias[1833:1833] = '{32'hc139ee4d};
test_output[1833:1833] = '{32'h462f311b};
test_input[14672:14679] = '{32'h41b5a0b6, 32'hc2807e79, 32'h4254812b, 32'h424b0a48, 32'h4271bbc6, 32'h42ab9e49, 32'hc261f7df, 32'hc256a11d};
test_weights[14672:14679] = '{32'hc2b779e3, 32'h428608c7, 32'hc279cfa9, 32'h428826c9, 32'h3fefd539, 32'h426a68aa, 32'hc2a648a7, 32'hc278dc2b};
test_bias[1834:1834] = '{32'h42a87959};
test_output[1834:1834] = '{32'h45db13a0};
test_input[14680:14687] = '{32'hc24e30da, 32'hc1704d56, 32'h4239a657, 32'hc1eb3804, 32'hc2098c9e, 32'h400ebb73, 32'h41fae066, 32'hc2964a78};
test_weights[14680:14687] = '{32'h416d2997, 32'hc2ae21df, 32'h416a3386, 32'hc200d9fa, 32'hc1f036f7, 32'hc2a35ce4, 32'hc290c207, 32'h405094ba};
test_bias[1835:1835] = '{32'hc184f98d};
test_output[1835:1835] = '{32'h43f491e8};
test_input[14688:14695] = '{32'h428c2bbe, 32'h416bec71, 32'hc13cf79a, 32'h42667f19, 32'h422db9c7, 32'h42686a55, 32'hc20798a3, 32'h42381228};
test_weights[14688:14695] = '{32'hc223dbc9, 32'hc1c0f17d, 32'hc2c7ca96, 32'h426ec95e, 32'hc20d6b5f, 32'hc287fda7, 32'h411e6ccd, 32'h41bcff5b};
test_bias[1836:1836] = '{32'h41610222};
test_output[1836:1836] = '{32'hc54ff9c9};
test_input[14696:14703] = '{32'h42126f69, 32'h422525e3, 32'hc1bb041e, 32'h423faf35, 32'h42b1fa8e, 32'hc2142111, 32'h42b99a74, 32'hc1c0e88b};
test_weights[14696:14703] = '{32'h422d9ff6, 32'h42b49953, 32'h41ecfdc5, 32'h4113f831, 32'hc28776e1, 32'h42a4e12a, 32'hc2644525, 32'hbffa569d};
test_bias[1837:1837] = '{32'h42690ae9};
test_output[1837:1837] = '{32'hc60fcc0f};
test_input[14704:14711] = '{32'hc210386e, 32'h42bf2299, 32'h4170b2e5, 32'h42c0c958, 32'h423ff336, 32'h42b4663c, 32'hc19e3286, 32'hc26331d9};
test_weights[14704:14711] = '{32'h4223fe94, 32'h428519c6, 32'h425e46aa, 32'hc228e75a, 32'h414448c6, 32'h3fb828f1, 32'h42918f22, 32'h41680360};
test_bias[1838:1838] = '{32'h41b2e99d};
test_output[1838:1838] = '{32'h42fb1058};
test_input[14712:14719] = '{32'h428eb3ba, 32'h41ee2c33, 32'h42a25b8e, 32'h4288bd4c, 32'hc2a19b4d, 32'hc2c4e94c, 32'hc1261d35, 32'hc156bf00};
test_weights[14712:14719] = '{32'hc207d594, 32'hc297dcc0, 32'hc187ae88, 32'hc29f3745, 32'h427660fb, 32'hc236f141, 32'h424c15ea, 32'h428b926e};
test_bias[1839:1839] = '{32'hc1b116e3};
test_output[1839:1839] = '{32'hc6526716};
test_input[14720:14727] = '{32'h42451f2a, 32'hc247885e, 32'hc278ef1e, 32'h42776331, 32'h42bfa559, 32'h420f6b5d, 32'hc252d91b, 32'h413b0846};
test_weights[14720:14727] = '{32'hc1f1afe9, 32'hc08c921a, 32'hc1a1d26a, 32'h422df19b, 32'h41ef63e2, 32'hc2049c02, 32'h42566049, 32'h42ac6179};
test_bias[1840:1840] = '{32'h409ad37b};
test_output[1840:1840] = '{32'h451f0a8f};
test_input[14728:14735] = '{32'hc1756b4a, 32'h42614220, 32'h4268c9b2, 32'h418cd3c3, 32'hc2b8b421, 32'h41a159c4, 32'hc299ab62, 32'h429b4c8b};
test_weights[14728:14735] = '{32'h42b8c032, 32'hc19282e7, 32'hc200dee6, 32'hc2a338a5, 32'hc19d278d, 32'h428f667d, 32'hc0bfe02f, 32'hc280b423};
test_bias[1841:1841] = '{32'h4295344e};
test_output[1841:1841] = '{32'hc5d9890f};
test_input[14736:14743] = '{32'h42b3a920, 32'h41ff905b, 32'hc297d433, 32'h41a5e366, 32'hc2086e77, 32'hc2901242, 32'hc24f212c, 32'h41a7ad44};
test_weights[14736:14743] = '{32'h42c0de70, 32'h427f94b9, 32'h42c165ca, 32'h4245e39a, 32'hc27aa1d6, 32'h422f8466, 32'hc228e154, 32'h418ff9b1};
test_bias[1842:1842] = '{32'h42138fd8};
test_output[1842:1842] = '{32'h45ba6c49};
test_input[14744:14751] = '{32'h423ebef2, 32'hbf36e374, 32'h423742d4, 32'h41bb67aa, 32'h40e901eb, 32'hc2617bc8, 32'hc2229c27, 32'h416fd1b6};
test_weights[14744:14751] = '{32'h41a3145a, 32'h42958bb2, 32'h4253d7cc, 32'h411ad001, 32'h42c070a6, 32'hc08e56f5, 32'hc15e30ee, 32'hc0916a98};
test_bias[1843:1843] = '{32'h4184c155};
test_output[1843:1843] = '{32'h459d6107};
test_input[14752:14759] = '{32'h4295768b, 32'h426be617, 32'h42b14a39, 32'hc091770e, 32'h415b9f94, 32'h42087a2e, 32'hc23f545e, 32'hc22ca441};
test_weights[14752:14759] = '{32'h4254f1d8, 32'hc18066b3, 32'hc0733385, 32'h40e8cd58, 32'h41856b7e, 32'hc2905585, 32'hc211aaa3, 32'h425a9b58};
test_bias[1844:1844] = '{32'h4163eceb};
test_output[1844:1844] = '{32'hc32e125b};
test_input[14760:14767] = '{32'hc2b22ecf, 32'h4206d0b9, 32'h4212ee6a, 32'hc2bfc410, 32'h401e09cd, 32'h42c5e964, 32'h429c67cf, 32'hc027319f};
test_weights[14760:14767] = '{32'hc1e6e244, 32'hc2abc589, 32'h42835e8e, 32'h41388d13, 32'h429291d9, 32'hc2c6c507, 32'hc294f47d, 32'hc1d7bc3c};
test_bias[1845:1845] = '{32'hc284a8cc};
test_output[1845:1845] = '{32'hc6626a69};
test_input[14768:14775] = '{32'hc1f741eb, 32'h42c1f7c9, 32'h412caf0e, 32'hc128cb3c, 32'h42c27c05, 32'h406f8fbd, 32'hc2666197, 32'hc2bb61cf};
test_weights[14768:14775] = '{32'hc2008a30, 32'hc1d1c73c, 32'hc2ae9ac9, 32'h41f0c89a, 32'hc210e4e1, 32'hc2b429a5, 32'h428efcbc, 32'hc2b8089a};
test_bias[1846:1846] = '{32'hc2c5d69d};
test_output[1846:1846] = '{32'hc50d8cd8};
test_input[14776:14783] = '{32'hc2148e7f, 32'h42131b82, 32'h42a7be4a, 32'hc2b9cbc7, 32'h41492809, 32'h40a0e70e, 32'h429d97d7, 32'hbfde73e9};
test_weights[14776:14783] = '{32'h417b335e, 32'h42a0fb87, 32'hc25d1f6b, 32'h41eb4d2c, 32'h40a2bdb0, 32'hc1c3a2e5, 32'h4229900d, 32'h42a81314};
test_bias[1847:1847] = '{32'hc1c18a05};
test_output[1847:1847] = '{32'hc4eb1842};
test_input[14784:14791] = '{32'hc1026ef1, 32'hc05f5f87, 32'h42aacf45, 32'h419e0b32, 32'h4298d963, 32'hc2948df4, 32'hc2a54a02, 32'h4106ae0d};
test_weights[14784:14791] = '{32'h41fc7fff, 32'hc29de3a7, 32'hc2a57cf4, 32'h423d6e4e, 32'h4216e460, 32'h41f8b916, 32'h407c4222, 32'hc06eb3b5};
test_bias[1848:1848] = '{32'h42ad2ead};
test_output[1848:1848] = '{32'hc5b58e9c};
test_input[14792:14799] = '{32'h410db8cb, 32'hc1ea8a2b, 32'hc2854d31, 32'h428fa3e7, 32'hc2a7de44, 32'hc2608330, 32'h4111ab06, 32'hc29c06ed};
test_weights[14792:14799] = '{32'hc1446316, 32'hc20152a1, 32'hc2c0b897, 32'h42414441, 32'hc28e15a4, 32'h41bd57ff, 32'hc2522e55, 32'h42aefab4};
test_bias[1849:1849] = '{32'hc2bedb7e};
test_output[1849:1849] = '{32'h45f8f7e2};
test_input[14800:14807] = '{32'hc2a08672, 32'hc261c733, 32'h4008e9af, 32'hc19130e2, 32'h4224a3fb, 32'hc23682d7, 32'h41c26c07, 32'hc257cd32};
test_weights[14800:14807] = '{32'hc19eee6a, 32'hc2bd73df, 32'h40a24370, 32'h421a7f07, 32'hc2bcb6d5, 32'hc0f96a8a, 32'h4245036b, 32'hc1df105d};
test_bias[1850:1850] = '{32'h42c74efe};
test_output[1850:1850] = '{32'h45aca008};
test_input[14808:14815] = '{32'hc1c37ce1, 32'hc103498b, 32'h42853e88, 32'hc2c05910, 32'h4273091f, 32'hc2c259ee, 32'h42bd4f6e, 32'hc0ff71af};
test_weights[14808:14815] = '{32'hc2a764a4, 32'h42715fb3, 32'hc2a68355, 32'hc2b208e7, 32'hc1a8fe8d, 32'h415f63d4, 32'h42427a05, 32'hc291db90};
test_bias[1851:1851] = '{32'h424751d2};
test_output[1851:1851] = '{32'h45dfb25a};
test_input[14816:14823] = '{32'h4180daa0, 32'hc1e7bc1a, 32'h42a6d445, 32'h428973e3, 32'hc20a89cf, 32'hc2c6ce06, 32'hc25c73a8, 32'hc2abe115};
test_weights[14816:14823] = '{32'h42afe4bc, 32'hc22c47b6, 32'hc23b454c, 32'hc29e97ac, 32'hc23586b2, 32'h41922e33, 32'h423ccff6, 32'h42bfc761};
test_bias[1852:1852] = '{32'h42bda6ae};
test_output[1852:1852] = '{32'hc68a25a2};
test_input[14824:14831] = '{32'hc2a54944, 32'hc2256cf2, 32'h421ab437, 32'h42c2bea0, 32'h423d9398, 32'h41572db9, 32'h42645f08, 32'h41efb0a6};
test_weights[14824:14831] = '{32'hc2a35dc4, 32'h422e693c, 32'hc11100a2, 32'hc2a1c7fd, 32'hc18f7328, 32'hc2953216, 32'h41cc1348, 32'h41e98e97};
test_bias[1853:1853] = '{32'h415e02f6};
test_output[1853:1853] = '{32'hc52e3ce9};
test_input[14832:14839] = '{32'hc1a93897, 32'h4247afac, 32'h421ee896, 32'h41b44829, 32'hc2622097, 32'h4275b5b8, 32'hc1fbaf9c, 32'h42ab872b};
test_weights[14832:14839] = '{32'h41ac4ce0, 32'h42c25da7, 32'h410135e3, 32'hc1c1e52f, 32'hc25ebb06, 32'hc18331b4, 32'hc19a09db, 32'h42ac7722};
test_bias[1854:1854] = '{32'hc1531a1d};
test_output[1854:1854] = '{32'h465f6d30};
test_input[14840:14847] = '{32'h427990db, 32'h422632fd, 32'hc202d6ea, 32'hc2bfafeb, 32'h426d30c1, 32'hc1c8bc59, 32'hc1c0bce5, 32'hc1b4fe92};
test_weights[14840:14847] = '{32'h415992d8, 32'h42040109, 32'h42b95aca, 32'hc1e07a16, 32'h42873649, 32'hc1fcb89d, 32'h4283caa6, 32'hc2b8525a};
test_bias[1855:1855] = '{32'h42ad6fae};
test_output[1855:1855] = '{32'h45e2f9d1};
test_input[14848:14855] = '{32'h41d02d82, 32'h41eecbd7, 32'h419a1843, 32'h40c5a646, 32'hc1c7bc06, 32'h42855913, 32'hc2c313ad, 32'h4239130d};
test_weights[14848:14855] = '{32'hc20b0000, 32'h428544dd, 32'hc1010be4, 32'h42b54a45, 32'h42520b00, 32'h422c31c5, 32'hc2a6ff7f, 32'h4245dd3f};
test_bias[1856:1856] = '{32'h417089aa};
test_output[1856:1856] = '{32'h4652e24b};
test_input[14856:14863] = '{32'hc292d7a1, 32'hc2a5fe7e, 32'hc132cf49, 32'hc221dc60, 32'hbd412305, 32'h42bff780, 32'hc2000c92, 32'h4197cbcf};
test_weights[14856:14863] = '{32'hc1448990, 32'h41f7f653, 32'h42724a8a, 32'h400fb8ed, 32'h4010c260, 32'h42b20c18, 32'hc1536a24, 32'hc2849022};
test_bias[1857:1857] = '{32'h41b14d55};
test_output[1857:1857] = '{32'h45a56dd1};
test_input[14864:14871] = '{32'hc2802ebd, 32'h4235fd54, 32'hc1ac2854, 32'hc167ec06, 32'hc1933a90, 32'h42a63264, 32'h42994c9a, 32'h3ffb2253};
test_weights[14864:14871] = '{32'h423db295, 32'h42baf4a1, 32'hc0ea6649, 32'hc2c12dfa, 32'hc0cc0c01, 32'hc1dd636f, 32'hc263aeac, 32'h42c570dd};
test_bias[1858:1858] = '{32'hbf485ed6};
test_output[1858:1858] = '{32'hc55fd189};
test_input[14872:14879] = '{32'hc29b2056, 32'hc2a97938, 32'hc0aa75a1, 32'hc2a71267, 32'hc1ba53f0, 32'h42af2924, 32'h4153a3c7, 32'h42a4774b};
test_weights[14872:14879] = '{32'hc2bb0e92, 32'hc214c068, 32'hc15584b2, 32'h41e85838, 32'h423d9828, 32'hc29d9953, 32'hc286e9c2, 32'hc1814031};
test_bias[1859:1859] = '{32'h42a02990};
test_output[1859:1859] = '{32'hc502f89d};
test_input[14880:14887] = '{32'h415dd0f6, 32'hc1ab2b9b, 32'hc27964e4, 32'h4278fd88, 32'hc28db1d0, 32'h40bd9c81, 32'hc23ddae4, 32'hc18d1084};
test_weights[14880:14887] = '{32'h4134da14, 32'h425b945e, 32'h418ba6d0, 32'hc2bef669, 32'hc2bd6d26, 32'h41951b34, 32'h4055c45c, 32'h41a051fc};
test_bias[1860:1860] = '{32'hc27dfe02};
test_output[1860:1860] = '{32'hc4e18fde};
test_input[14888:14895] = '{32'hc2a9cdc3, 32'h419d27b7, 32'h42810e05, 32'hc27cef6c, 32'h428d3d44, 32'h42be22de, 32'h418eb24c, 32'hc0e013e4};
test_weights[14888:14895] = '{32'hc29eadbf, 32'h41fe176c, 32'hc0cf2f1f, 32'h4254dff2, 32'h3fd1fd18, 32'hc2351082, 32'hc1ddd773, 32'hc0c3e607};
test_bias[1861:1861] = '{32'hc03cae07};
test_output[1861:1861] = '{32'hc4852735};
test_input[14896:14903] = '{32'h42835003, 32'hc2193833, 32'h42bfe453, 32'hc29dce98, 32'h42414a4f, 32'h42c7d7fb, 32'hc18823eb, 32'h403f0b93};
test_weights[14896:14903] = '{32'h42b6ab1d, 32'h41c47149, 32'hc298381f, 32'h42816c0d, 32'h4110bfac, 32'hbf8150e8, 32'hc2aeb33e, 32'h427c75aa};
test_bias[1862:1862] = '{32'h42088854};
test_output[1862:1862] = '{32'hc5a5d836};
test_input[14904:14911] = '{32'h41d0b7cf, 32'h429efbf9, 32'hc2c112c6, 32'h427ffef5, 32'hc28e33ba, 32'hc138331c, 32'h42bace46, 32'hc2a03228};
test_weights[14904:14911] = '{32'hc2955e3f, 32'hc2ae626c, 32'h422dc711, 32'h410c129b, 32'h40849e44, 32'hc1c5c185, 32'h40c658b2, 32'h42850c23};
test_bias[1863:1863] = '{32'hc126e551};
test_output[1863:1863] = '{32'hc6870689};
test_input[14912:14919] = '{32'h418fe464, 32'h42beba78, 32'hc29590ad, 32'h42032591, 32'h4273fa31, 32'hc0c04fe5, 32'h4217b629, 32'h427d0d72};
test_weights[14912:14919] = '{32'h41c6d8e9, 32'h41af9894, 32'hc24123a4, 32'h429dd2b9, 32'hc2c35cb4, 32'h42823279, 32'hc2b52b46, 32'h4260ce37};
test_bias[1864:1864] = '{32'hc2385602};
test_output[1864:1864] = '{32'h4519edf9};
test_input[14920:14927] = '{32'hc214ebeb, 32'h42ab9aab, 32'h424a8c92, 32'hc2c0ca75, 32'hc29fcefc, 32'hc27b9782, 32'hc264630b, 32'hc2b60383};
test_weights[14920:14927] = '{32'h40f64d55, 32'h421bd087, 32'h42aa1966, 32'hc12f7441, 32'hc26b7c21, 32'h4285fc12, 32'h419e1ad8, 32'hc19f5536};
test_bias[1865:1865] = '{32'h42191326};
test_output[1865:1865] = '{32'h46168119};
test_input[14928:14935] = '{32'h4236af6c, 32'h42ad68c0, 32'hc28f7c8d, 32'h429ac11e, 32'hc0504088, 32'hc24ff66d, 32'h4264babc, 32'h421db10a};
test_weights[14928:14935] = '{32'hc279b2da, 32'hc2b9f50f, 32'hc2b30e04, 32'h416c525a, 32'h42a0f7b9, 32'hc1b331fe, 32'h4201f93c, 32'hc29573c8};
test_bias[1866:1866] = '{32'hc1f91da7};
test_output[1866:1866] = '{32'hc55eb2d0};
test_input[14936:14943] = '{32'h4128c74e, 32'h42c74f56, 32'hc2a969f3, 32'h426d9a81, 32'hc2bbeb6e, 32'h42549d06, 32'h427b5bab, 32'hc25363e2};
test_weights[14936:14943] = '{32'hc1fcf7c6, 32'h3e90417a, 32'h428d934d, 32'h4241f564, 32'h4282c823, 32'h4248fcb2, 32'h4283d7cc, 32'h40f74755};
test_bias[1867:1867] = '{32'h40a82fff};
test_output[1867:1867] = '{32'hc545357a};
test_input[14944:14951] = '{32'hc1ebe334, 32'h425a45e9, 32'hc244012d, 32'h429fa5bc, 32'h42b1d034, 32'h41a6ead4, 32'h429d3e2e, 32'hc2a93939};
test_weights[14944:14951] = '{32'h4298619f, 32'h426b79c4, 32'h4122900b, 32'h42936704, 32'h40c77505, 32'h42c7a1dd, 32'hc141ca3a, 32'hc24af084};
test_bias[1868:1868] = '{32'hc24dbfb7};
test_output[1868:1868] = '{32'h463fd3b8};
test_input[14952:14959] = '{32'h41673142, 32'h426d124b, 32'h428de619, 32'h427d2b9f, 32'hc29d6a3b, 32'hc2bc38c8, 32'hc284b6eb, 32'hc29a2bd0};
test_weights[14952:14959] = '{32'h42b1c89b, 32'hc2790bf0, 32'h41f8f5d6, 32'h42115688, 32'h42543730, 32'hc12db003, 32'hc2c6cb26, 32'h42a6c383};
test_bias[1869:1869] = '{32'h427d6023};
test_output[1869:1869] = '{32'hc44d289b};
test_input[14960:14967] = '{32'h3eb4c441, 32'h40cec229, 32'hc0839181, 32'h423782f5, 32'hc28c946c, 32'hc1c925e7, 32'h426c2857, 32'h4235f3ae};
test_weights[14960:14967] = '{32'h4295b576, 32'h42255334, 32'h427d1ffc, 32'h428c8c23, 32'h42be22d7, 32'hbfb9a668, 32'h41fc537c, 32'hc2b870ae};
test_bias[1870:1870] = '{32'hc2be62c3};
test_output[1870:1870] = '{32'hc5b5c3fc};
test_input[14968:14975] = '{32'h42b06493, 32'hc29823bd, 32'hc27f0249, 32'h42af793c, 32'hc1e44317, 32'h4225aa44, 32'h4204036e, 32'h41948bdd};
test_weights[14968:14975] = '{32'hc1db78bc, 32'h429bd204, 32'h427cad5a, 32'hc23c5f03, 32'hc2b86632, 32'hc222b41d, 32'hc17f4761, 32'h428e8ecb};
test_bias[1871:1871] = '{32'hc1279fa3};
test_output[1871:1871] = '{32'hc666d25e};
test_input[14976:14983] = '{32'h4185dc47, 32'h419ef3f5, 32'h42267a26, 32'hc27143d4, 32'hc2a5f1de, 32'h4299e834, 32'hc167d0c0, 32'hbf9ba5e7};
test_weights[14976:14983] = '{32'hc252f6de, 32'hc28e9c7f, 32'h429fc700, 32'hc1161b43, 32'h425feeb0, 32'h42390606, 32'h425786ef, 32'hc256c96b};
test_bias[1872:1872] = '{32'h4131490b};
test_output[1872:1872] = '{32'hc3464905};
test_input[14984:14991] = '{32'h427db14d, 32'hc280bb96, 32'h4164004e, 32'h409a2b9c, 32'h41cdb097, 32'hc269113d, 32'h4263e15e, 32'hc2504fcd};
test_weights[14984:14991] = '{32'h42a38d0b, 32'h422ed39c, 32'hc22577e2, 32'hc270e4ad, 32'hc214c18c, 32'hc186867b, 32'hc091d051, 32'h427455f3};
test_bias[1873:1873] = '{32'hc2b08059};
test_output[1873:1873] = '{32'hc4fb784e};
test_input[14992:14999] = '{32'h4237ff57, 32'hc2aede18, 32'h42c33bfa, 32'h41a473ce, 32'hc2c6bce7, 32'h42479431, 32'hc2c737c2, 32'h41e6cd6e};
test_weights[14992:14999] = '{32'hc27220ac, 32'hc21533e8, 32'h408c6829, 32'h42448e60, 32'h4208abfc, 32'h4205cdc5, 32'h42c3fa39, 32'h42797313};
test_bias[1874:1874] = '{32'hc202b64f};
test_output[1874:1874] = '{32'hc5f3e73c};
test_input[15000:15007] = '{32'hc128b8b9, 32'hc1de1118, 32'hc22f2409, 32'h42aa8b4d, 32'hc2947b47, 32'h42b126d8, 32'h41c59d7b, 32'hc068cd03};
test_weights[15000:15007] = '{32'hc21eec90, 32'hc28af61f, 32'hc298a0d0, 32'h422b5006, 32'h41de4d56, 32'h425b316b, 32'hc22b246c, 32'h42b5d5bb};
test_bias[1875:1875] = '{32'h42198c10};
test_output[1875:1875] = '{32'h46287add};
test_input[15008:15015] = '{32'hc1afa0ef, 32'hbfa23db7, 32'h42c2b42b, 32'h42156582, 32'h41ff00f7, 32'hc26cef56, 32'hc29050b4, 32'h420d1f36};
test_weights[15008:15015] = '{32'hc2a06d94, 32'h4290adba, 32'h40ff9d5f, 32'hc2ab914f, 32'h4253e02a, 32'h42ab1e41, 32'hc2b66c8d, 32'hc2514134};
test_bias[1876:1876] = '{32'hc23b69eb};
test_output[1876:1876] = '{32'h440a232c};
test_input[15016:15023] = '{32'h41b93233, 32'hc0512f76, 32'h427509f7, 32'h4202dcc8, 32'hc09bea19, 32'h41f84ca7, 32'hc20ddcab, 32'h4271563c};
test_weights[15016:15023] = '{32'hc2281ef9, 32'h40208a22, 32'h3b19dda9, 32'hc1ee5566, 32'hc2860c3e, 32'hc0f546a8, 32'hc165bcd0, 32'hc253ccb6};
test_bias[1877:1877] = '{32'h420757b4};
test_output[1877:1877] = '{32'hc58d3528};
test_input[15024:15031] = '{32'h4233f691, 32'h4257d017, 32'h42824cde, 32'hc2bc770a, 32'h424836a1, 32'h42c502bf, 32'h41f4ca5f, 32'h42802a49};
test_weights[15024:15031] = '{32'hc24cdb3b, 32'hc1c1614b, 32'h422eb630, 32'h4256a956, 32'hc22af5f4, 32'hc213c31e, 32'hc27c83f2, 32'h4284ee74};
test_bias[1878:1878] = '{32'hc09b9793};
test_output[1878:1878] = '{32'hc610ec73};
test_input[15032:15039] = '{32'h42b672f6, 32'h420bb9f2, 32'h41daa4ee, 32'hc25b80c1, 32'h413bfa66, 32'h4235e331, 32'h423f0c2a, 32'h42c65395};
test_weights[15032:15039] = '{32'hc216c9c4, 32'hc2236a09, 32'hc24bcb3d, 32'h426036db, 32'h40e1688d, 32'h42bc0692, 32'h42027dd7, 32'hc2bec659};
test_bias[1879:1879] = '{32'hc1c4b8f1};
test_output[1879:1879] = '{32'hc649985d};
test_input[15040:15047] = '{32'hc24335d5, 32'h428df28b, 32'h41ae6cc7, 32'h42427c91, 32'hc21dc778, 32'hc1a1e38e, 32'h408abfff, 32'hc2a7824b};
test_weights[15040:15047] = '{32'hc2174d7c, 32'hc2a53198, 32'hc14acabd, 32'hc206fc78, 32'hc2b15965, 32'hc2c3c8e4, 32'hc2c0f998, 32'h410cc0fc};
test_bias[1880:1880] = '{32'hc2ade696};
test_output[1880:1880] = '{32'hc4d418b7};
test_input[15048:15055] = '{32'hc2c76942, 32'h42a702d8, 32'hc2c7a183, 32'hc19f7623, 32'hc28e2ef8, 32'h427c9ab7, 32'h41c081eb, 32'h41f35a0f};
test_weights[15048:15055] = '{32'h42a0a389, 32'h41fa7965, 32'h420e7dba, 32'h42518bc3, 32'hc299437a, 32'h41ba54fa, 32'h42b57ff8, 32'hc2569a01};
test_bias[1881:1881] = '{32'hc24d7e30};
test_output[1881:1881] = '{32'hc520e8a4};
test_input[15056:15063] = '{32'h40b1f9f5, 32'h4278c189, 32'h41e61556, 32'h40fe950f, 32'hc26cc420, 32'h424fa782, 32'h4237b6ee, 32'h42a4c760};
test_weights[15056:15063] = '{32'h42135dba, 32'h41be7cf6, 32'h42741563, 32'h42a65241, 32'h414c2cce, 32'h42c755d9, 32'hc22135b8, 32'hbfdb84d7};
test_bias[1882:1882] = '{32'hc1bdee83};
test_output[1882:1882] = '{32'h45cb47b8};
test_input[15064:15071] = '{32'h42a8563c, 32'h421931c2, 32'h427c93a6, 32'h41a4ca3d, 32'hc063ecc5, 32'hc28de711, 32'hc2ae4f0c, 32'hc211e1dd};
test_weights[15064:15071] = '{32'h4195895f, 32'h41c99787, 32'hc2568c3a, 32'hbffc733e, 32'hc18873dc, 32'hc2177486, 32'hc2816268, 32'h42af0c90};
test_bias[1883:1883] = '{32'hc14c664d};
test_output[1883:1883] = '{32'h45861bcc};
test_input[15072:15079] = '{32'hc1c98289, 32'hc2b1be81, 32'hc26aec9d, 32'hc2c06ef0, 32'hc2b5d2f0, 32'hc2aa3120, 32'h4248c893, 32'h426548a6};
test_weights[15072:15079] = '{32'h41a33680, 32'hc21c352a, 32'hc2bc4f04, 32'h4299ddc8, 32'h42badd46, 32'hc2a98ce6, 32'h41ad9f64, 32'h4247115c};
test_bias[1884:1884] = '{32'h42791712};
test_output[1884:1884] = '{32'h456e089f};
test_input[15080:15087] = '{32'hc2b9df4b, 32'h41bff120, 32'hc1ff5e85, 32'h41c62422, 32'h428c01ad, 32'hc136aa47, 32'hc28650fe, 32'hc1b6ab30};
test_weights[15080:15087] = '{32'h42282429, 32'hc1e94877, 32'hc28bef0a, 32'hc2b8121f, 32'h42b577e0, 32'hc26950ff, 32'hc2628da2, 32'h42a0ebe9};
test_bias[1885:1885] = '{32'hc27b2394};
test_output[1885:1885] = '{32'h45856834};
test_input[15088:15095] = '{32'h422d6f01, 32'hc0cde6eb, 32'hc28ce15d, 32'h41af5ace, 32'h429dc5bb, 32'h42bd673f, 32'hc16cce7c, 32'h41dc7b1d};
test_weights[15088:15095] = '{32'hc2451a19, 32'hc2742597, 32'h4274ebe6, 32'h418e5451, 32'hc1a1a9e2, 32'hc2292408, 32'h42a8dd78, 32'hc295b500};
test_bias[1886:1886] = '{32'h428b4b87};
test_output[1886:1886] = '{32'hc662b1c4};
test_input[15096:15103] = '{32'hc28e5071, 32'h41e2796f, 32'h423c0ad2, 32'hc2b6eb8f, 32'hc188577e, 32'hc21d3835, 32'hc2049664, 32'hc249bc5d};
test_weights[15096:15103] = '{32'hc2b3073f, 32'h41a2ca3e, 32'h42ac5a63, 32'h42bdb8b9, 32'h42768000, 32'hc2b26590, 32'hc268581f, 32'h409a692c};
test_bias[1887:1887] = '{32'hc2596235};
test_output[1887:1887] = '{32'h45c82198};
test_input[15104:15111] = '{32'hc269ce30, 32'h422cfa95, 32'h4206f69f, 32'h42405a98, 32'h42952246, 32'hc1f7ff8f, 32'h4286b1b6, 32'h42a71aea};
test_weights[15104:15111] = '{32'h413e69fb, 32'h418750bd, 32'hc1d410b8, 32'hc2a18c7a, 32'hc27721c1, 32'hc23dea88, 32'hc218a8c1, 32'h42b8bc5f};
test_bias[1888:1888] = '{32'h428fedff};
test_output[1888:1888] = '{32'hc5262c2b};
test_input[15112:15119] = '{32'h4203fd50, 32'hc279bf05, 32'hc2b62811, 32'h42ba63be, 32'h42b401a0, 32'hc0e8eafc, 32'h4191b348, 32'hc2b0b3e9};
test_weights[15112:15119] = '{32'hc23806b0, 32'hc28b6915, 32'hc105e7fd, 32'hc1a8af1c, 32'h424d3aaa, 32'hc1ca8b84, 32'h413a97e2, 32'h42830611};
test_bias[1889:1889] = '{32'h42c62f36};
test_output[1889:1889] = '{32'h446f3186};
test_input[15120:15127] = '{32'hc2880c5d, 32'h42656ae9, 32'hc25209de, 32'h42906346, 32'hc2870c92, 32'hc28bc294, 32'hc21eab5f, 32'hc1caedf6};
test_weights[15120:15127] = '{32'h42b74403, 32'hc2588310, 32'hc22cff74, 32'hc2a85412, 32'hc1c64cb9, 32'h4293b4c9, 32'hc27910d2, 32'hc2bfe514};
test_bias[1890:1890] = '{32'h42c4d056};
test_output[1890:1890] = '{32'hc635af19};
test_input[15128:15135] = '{32'h428b6994, 32'h3e85dcfa, 32'h429852c6, 32'hc1bb1249, 32'hc2aa735b, 32'h42bed102, 32'h41e320ef, 32'hc10bc122};
test_weights[15128:15135] = '{32'hc038a099, 32'h41c75a20, 32'hc2a55a93, 32'hc1a01fa0, 32'hc267a906, 32'h42bc677a, 32'h41b51f2d, 32'h4195780b};
test_bias[1891:1891] = '{32'hc1d01664};
test_output[1891:1891] = '{32'h460286db};
test_input[15136:15143] = '{32'h4278c8a9, 32'h42c2e3dc, 32'hc195d63f, 32'h41856a26, 32'hc23b634e, 32'h421cf3c2, 32'hbfb53e32, 32'h4101119e};
test_weights[15136:15143] = '{32'h42c4568c, 32'hc1bc99e7, 32'h422168bc, 32'h42b849ce, 32'hc267dd11, 32'hc267b0e8, 32'h41e7796e, 32'hc1dfeec5};
test_bias[1892:1892] = '{32'h423e4ea0};
test_output[1892:1892] = '{32'h4596670c};
test_input[15144:15151] = '{32'hc2b08a96, 32'hc27467a7, 32'hc240ee51, 32'h425e862e, 32'hc140d093, 32'h414c2f3b, 32'h42ae6380, 32'h426f41dc};
test_weights[15144:15151] = '{32'hc1a8e079, 32'hc1bec623, 32'h42b1153c, 32'h41c90433, 32'h41802db8, 32'hc213c76c, 32'h42ac3e0f, 32'h40f0aa20};
test_bias[1893:1893] = '{32'h42c15326};
test_output[1893:1893] = '{32'h45f4f746};
test_input[15152:15159] = '{32'hbfc01930, 32'hc2bb5b00, 32'h41f5a8a5, 32'hc26c8b66, 32'hc241ebbb, 32'hc278f804, 32'h42bd3ead, 32'h41e11f94};
test_weights[15152:15159] = '{32'hc22028dc, 32'h4276b1bb, 32'h41fc32ec, 32'hc2acc661, 32'hc1172832, 32'hc145970d, 32'h4114b802, 32'hc1e4e733};
test_bias[1894:1894] = '{32'hc12c109e};
test_output[1894:1894] = '{32'h44ce31a6};
test_input[15160:15167] = '{32'h4212804f, 32'h3ee55858, 32'h425e80d0, 32'hc2554391, 32'h429dcb05, 32'h42930ec7, 32'hc1f87866, 32'hc2262ad9};
test_weights[15160:15167] = '{32'h4263b4ef, 32'h428f46ee, 32'h41064e73, 32'h41650248, 32'h4296b4d4, 32'h425ab0b2, 32'h42c1d0de, 32'h41e94362};
test_bias[1895:1895] = '{32'h427b7299};
test_output[1895:1895] = '{32'h45ee5dcb};
test_input[15168:15175] = '{32'hc2acf951, 32'h41a58d8b, 32'hc1e7a35d, 32'hc25aa41a, 32'hc21a5c2a, 32'h427804a7, 32'hc2b8b842, 32'hc27af267};
test_weights[15168:15175] = '{32'h40bef690, 32'h42aeac4b, 32'hc1f4fa91, 32'h41ac960f, 32'hc15c63b2, 32'hc2307757, 32'hc2719d22, 32'h41514237};
test_bias[1896:1896] = '{32'hc0d752f7};
test_output[1896:1896] = '{32'h455da6f3};
test_input[15176:15183] = '{32'h42210ac5, 32'h40b029eb, 32'h419b1162, 32'h42a78526, 32'h42bac7b1, 32'hc2b8ddbe, 32'h41c396a4, 32'h4271aa75};
test_weights[15176:15183] = '{32'hc0827d3e, 32'h41bd17b5, 32'hc210cfa6, 32'hc187e99b, 32'h411906dd, 32'hc2827f67, 32'h41bed44b, 32'h3f44133a};
test_bias[1897:1897] = '{32'hc2504019};
test_output[1897:1897] = '{32'h45a6f7a6};
test_input[15184:15191] = '{32'h423f7ad1, 32'hc2286193, 32'hc2403788, 32'hc142fa5b, 32'h4250fa4b, 32'h428e20cf, 32'hc1fe134c, 32'h429c78f0};
test_weights[15184:15191] = '{32'h42c720c9, 32'hc2a3f6f0, 32'hc2a08883, 32'hc23aaa7d, 32'h42329dc2, 32'hc20997fc, 32'hc25b2cca, 32'hc1fc2b5b};
test_bias[1898:1898] = '{32'hc142b094};
test_output[1898:1898] = '{32'h463845a7};
test_input[15192:15199] = '{32'hc059a619, 32'hc10be1cb, 32'h417287eb, 32'h4145b636, 32'hc23cd863, 32'h413739fd, 32'hc2252a78, 32'h42a0e77e};
test_weights[15192:15199] = '{32'h42455889, 32'hc2246df3, 32'h42880535, 32'hc2b65da3, 32'hc2aa7579, 32'hc1d1be08, 32'hc2ae2b25, 32'h42c14d76};
test_bias[1899:1899] = '{32'h42c70604};
test_output[1899:1899] = '{32'h466ee9ea};
test_input[15200:15207] = '{32'hc2212f78, 32'h42aacfa5, 32'hc28efd47, 32'h42b8d49a, 32'h424b5b2a, 32'hc2961cc0, 32'hc274bef8, 32'hc225a713};
test_weights[15200:15207] = '{32'hc282371e, 32'hc2a080df, 32'h4211a1f1, 32'hc12e9cec, 32'hc035ac74, 32'h424eddc7, 32'hc08077f8, 32'hc2655682};
test_bias[1900:1900] = '{32'h4292a805};
test_output[1900:1900] = '{32'hc60f59e6};
test_input[15208:15215] = '{32'hc23a9a1c, 32'hc1d1fe70, 32'h41724b62, 32'h425de251, 32'hc26e40ad, 32'hc1f19c73, 32'h42604b2c, 32'h41f1157a};
test_weights[15208:15215] = '{32'h4294be0a, 32'h416b343a, 32'h416c4ddc, 32'h42172d17, 32'h4241f81f, 32'hc1f6307c, 32'hc27eb39b, 32'h428b94ac};
test_bias[1901:1901] = '{32'h429975fa};
test_output[1901:1901] = '{32'hc598a5f0};
test_input[15216:15223] = '{32'hc22f15f8, 32'h42b55192, 32'hc2468c88, 32'hc25fd9be, 32'h429bb827, 32'hc1bd4d93, 32'hc0a22ffd, 32'hc2be4917};
test_weights[15216:15223] = '{32'hc2822e88, 32'h4217c9cc, 32'hc23af2b0, 32'hc08ef50f, 32'hc219c309, 32'hc1aca4d7, 32'h42c58f6f, 32'hc29a6f78};
test_bias[1902:1902] = '{32'h4217e6cf};
test_output[1902:1902] = '{32'h464f3405};
test_input[15224:15231] = '{32'hc28a9915, 32'h4222603c, 32'hc09ac364, 32'h42ba0f05, 32'h42656e6e, 32'hc235934d, 32'h4120455a, 32'hc2bc9466};
test_weights[15224:15231] = '{32'hc10beded, 32'hc1d3f258, 32'h41061d91, 32'h42b4b675, 32'hc0526843, 32'hc2c1fd32, 32'h42352f68, 32'h41b773b3};
test_bias[1903:1903] = '{32'hc2ac7d5a};
test_output[1903:1903] = '{32'h46212e07};
test_input[15232:15239] = '{32'hc2c11410, 32'h42a47cd3, 32'h42c61aab, 32'hc164e11f, 32'h423157fd, 32'hc2253a2d, 32'hc2b5b238, 32'hc233161d};
test_weights[15232:15239] = '{32'hc21cf5ce, 32'hc0b1317c, 32'h41899a28, 32'h421c644a, 32'hc0a1c0d7, 32'h413a8218, 32'h41e44709, 32'h42b64447};
test_bias[1904:1904] = '{32'hc2b3c8db};
test_output[1904:1904] = '{32'hc53aeca2};
test_input[15240:15247] = '{32'h42337d70, 32'hc2bcf20d, 32'h422591c5, 32'h420b5d1e, 32'h422a05b2, 32'hc1fd9bcf, 32'hc2391e1f, 32'hc247a9e8};
test_weights[15240:15247] = '{32'hc21ca83c, 32'hc25fe1c3, 32'hc2bbeb6e, 32'hc2486247, 32'hc09d7ed2, 32'hc29b8328, 32'h42bdb664, 32'h42a1b239};
test_bias[1905:1905] = '{32'h421fe690};
test_output[1905:1905] = '{32'hc600a860};
test_input[15248:15255] = '{32'h424ad55e, 32'hc221e1d8, 32'h41e2046f, 32'h4210a7f0, 32'hc2851a04, 32'h4281ebf8, 32'hc27f4be4, 32'hc1f2f0c0};
test_weights[15248:15255] = '{32'hc210d7c4, 32'hc181c1a3, 32'h42a48334, 32'h41f75d0b, 32'h42bac1eb, 32'h41919ed0, 32'hc27c650a, 32'h42439137};
test_bias[1906:1906] = '{32'h41fc63f6};
test_output[1906:1906] = '{32'hc34395e0};
test_input[15256:15263] = '{32'h409f64b8, 32'hc1e8011a, 32'h40b7037f, 32'h41d6a5b0, 32'hc2448348, 32'hc2b0c97d, 32'hc1ae718c, 32'hc25a9bdc};
test_weights[15256:15263] = '{32'h42a44c08, 32'h42c4d1bf, 32'hc27107db, 32'h3ecd9ba5, 32'hc28d2d95, 32'hc1ce20ab, 32'hc1bc970b, 32'h428156dc};
test_bias[1907:1907] = '{32'h425978cd};
test_output[1907:1907] = '{32'h3f6c4b64};
test_input[15264:15271] = '{32'h42699bfd, 32'hc29112ed, 32'hc29d59e2, 32'h425eb45e, 32'h4228aa2a, 32'hc24744d6, 32'h4246f1aa, 32'h4180d3df};
test_weights[15264:15271] = '{32'hc27f287a, 32'h41e55e1a, 32'hc29f3a3a, 32'h42c53e49, 32'h42b5eaa0, 32'hc0a1ace1, 32'h410d0767, 32'hc2baf910};
test_bias[1908:1908] = '{32'h3f5a074e};
test_output[1908:1908] = '{32'h460c28d4};
test_input[15272:15279] = '{32'hc217fa6e, 32'hc01d7e3d, 32'hc2bbaad6, 32'h428f86f1, 32'h42876a14, 32'h41fdc3a1, 32'h42910f04, 32'h4271e604};
test_weights[15272:15279] = '{32'h4226cf45, 32'h412b7517, 32'hc23e863a, 32'h42af4a1b, 32'hc20fb650, 32'hc2ba8b90, 32'hc2b7dcd9, 32'hc24e6959};
test_bias[1909:1909] = '{32'hc2ad5c3e};
test_output[1909:1909] = '{32'hc5bf3056};
test_input[15280:15287] = '{32'hc2b838f9, 32'hc239ff13, 32'hc2291fa4, 32'hc291516e, 32'hc247b8a5, 32'hc21360c9, 32'h41f34a7c, 32'hc2b8b990};
test_weights[15280:15287] = '{32'h42c18c6f, 32'h422c0a58, 32'h429e75b5, 32'hc157d49b, 32'h419a0d65, 32'h426df008, 32'h42887e57, 32'hc22b11e6};
test_bias[1910:1910] = '{32'hc286e218};
test_output[1910:1910] = '{32'hc623baef};
test_input[15288:15295] = '{32'h42bc5225, 32'h412a804a, 32'hc160c91d, 32'h4221a8b7, 32'h42aabe3f, 32'h426e60ee, 32'hc2840f21, 32'hc1ec6a5c};
test_weights[15288:15295] = '{32'h42c0e1ec, 32'hc2c79381, 32'hc2b2a2c7, 32'hc259cf52, 32'h41608dfd, 32'hc153ae17, 32'h41db5ff1, 32'h41dc8438};
test_bias[1911:1911] = '{32'h3fd673be};
test_output[1911:1911] = '{32'h4597cf21};
test_input[15296:15303] = '{32'hc1d73558, 32'h42b6190f, 32'hc243bd9e, 32'hc1bede42, 32'hc1b34c89, 32'hc1cc7230, 32'hc20bb506, 32'hc2a977c2};
test_weights[15296:15303] = '{32'hc0bcdac6, 32'h4294b230, 32'hc20bb3a9, 32'hc290727c, 32'h4282805a, 32'hc23aad2e, 32'h423b165d, 32'hc2a3a9e1};
test_bias[1912:1912] = '{32'h425f0619};
test_output[1912:1912] = '{32'h46715a8d};
test_input[15304:15311] = '{32'hc28ad277, 32'h4288d70d, 32'hc1900544, 32'hc2a40a46, 32'hc1c7f935, 32'h4032b739, 32'hc25b00b1, 32'h41fbdae0};
test_weights[15304:15311] = '{32'hc25a9f38, 32'hc2b72aa5, 32'h4212eadf, 32'h42b7c383, 32'hc1c4196a, 32'hc2791a1d, 32'hc1f7292b, 32'hc2c255f9};
test_bias[1913:1913] = '{32'h42b9e37a};
test_output[1913:1913] = '{32'hc633c62a};
test_input[15312:15319] = '{32'hc2495699, 32'h42b67936, 32'h428db074, 32'h42bf0394, 32'hc209244d, 32'hc2199c5d, 32'h428a54f4, 32'h42495d71};
test_weights[15312:15319] = '{32'h425eec5a, 32'hc217e121, 32'hc1c127d4, 32'h41a0f0bb, 32'h42a3006d, 32'h42bd44eb, 32'h428382d7, 32'hc2a70750};
test_bias[1914:1914] = '{32'hc2beaaac};
test_output[1914:1914] = '{32'hc63f3a5d};
test_input[15320:15327] = '{32'h41edee4f, 32'h423b6719, 32'hc293ee88, 32'hc2a24a65, 32'h4079d6dc, 32'hc24bdad4, 32'hc2442538, 32'hc2a3cb2d};
test_weights[15320:15327] = '{32'hc2c572f9, 32'h41384812, 32'h41db509d, 32'h417f1174, 32'h42bb5c30, 32'h428c2897, 32'hc1bb2b07, 32'h42b504c1};
test_bias[1915:1915] = '{32'h4209a2c1};
test_output[1915:1915] = '{32'hc66cc9ea};
test_input[15328:15335] = '{32'hc2419210, 32'hc2955a6f, 32'h42019b72, 32'hc219f320, 32'h42abc74e, 32'h428d9f6f, 32'h421d2e07, 32'hc233a533};
test_weights[15328:15335] = '{32'h4294994a, 32'h4226b944, 32'hc2bd9df0, 32'h4290a1be, 32'h41878412, 32'h426395b5, 32'hc2abea58, 32'h41820d66};
test_bias[1916:1916] = '{32'h421e0cb0};
test_output[1916:1916] = '{32'hc62e2f50};
test_input[15336:15343] = '{32'hc133978d, 32'hc1c031df, 32'h40d539ab, 32'hc2211f2f, 32'h42a38e0b, 32'hc0a43128, 32'hc261ac68, 32'hc215417c};
test_weights[15336:15343] = '{32'hbf884048, 32'h42bc9ba3, 32'hc2357fde, 32'hc2629934, 32'h425221f6, 32'hc2ac152d, 32'hc2647bff, 32'h428dfa84};
test_bias[1917:1917] = '{32'hc200bf45};
test_output[1917:1917] = '{32'h459c67e9};
test_input[15344:15351] = '{32'hc29e7d26, 32'hc21cc2fe, 32'h4286f913, 32'h421eca7b, 32'hc1ee3623, 32'hc2c08691, 32'h4158a3bc, 32'h4282042a};
test_weights[15344:15351] = '{32'hc246612e, 32'hc291978e, 32'hc2b2e135, 32'h42b39128, 32'h4179222a, 32'hc285cd01, 32'hc0dab126, 32'h42689a85};
test_bias[1918:1918] = '{32'hc081f7b5};
test_output[1918:1918] = '{32'h465a4d3e};
test_input[15352:15359] = '{32'hc2ba0794, 32'hc0f1cd57, 32'hc2492334, 32'hc292ec7f, 32'h41e72be7, 32'hc24dd759, 32'hc204a701, 32'hc1d54318};
test_weights[15352:15359] = '{32'hc17117fb, 32'hc1a2296f, 32'hc230a2ff, 32'hc0ad9f6c, 32'h41aa24b5, 32'h42807335, 32'h41d313e5, 32'h422e1b29};
test_bias[1919:1919] = '{32'hc291464a};
test_output[1919:1919] = '{32'hc41c250a};
test_input[15360:15367] = '{32'h42670334, 32'h428df5df, 32'h3f7c0c72, 32'hc156e102, 32'h428aadff, 32'h424f7717, 32'h4211e2fb, 32'h423eb9f0};
test_weights[15360:15367] = '{32'h41a72a92, 32'h41eb2de8, 32'h4264b909, 32'hc238a8f0, 32'h3f8738d8, 32'hc20c1cb2, 32'hc0e81b42, 32'hc2af70ef};
test_bias[1920:1920] = '{32'h42c07540};
test_output[1920:1920] = '{32'hc504cc43};
test_input[15368:15375] = '{32'h420527b1, 32'hc2bd5bb8, 32'hc23096bb, 32'hc21e15f2, 32'hc017bb32, 32'h42bd059c, 32'hc296a33d, 32'h4242bc8b};
test_weights[15368:15375] = '{32'hc2893e67, 32'h41cae099, 32'h4237ff7c, 32'hc230fae4, 32'hc18715ec, 32'h42573145, 32'hc06ed947, 32'hc18ef535};
test_bias[1921:1921] = '{32'h409e233d};
test_output[1921:1921] = '{32'hc3d5718e};
test_input[15376:15383] = '{32'h423e6446, 32'hc1540010, 32'hc0931ea4, 32'h4282d678, 32'h42c3f708, 32'hc297e567, 32'h41c1e872, 32'h40d5ea40};
test_weights[15376:15383] = '{32'h427d163c, 32'hc1bbc96c, 32'h42a1d804, 32'h428ba8ed, 32'hc1830200, 32'hc1ddf01e, 32'h4233f871, 32'hc26b542c};
test_bias[1922:1922] = '{32'hc22793f0};
test_output[1922:1922] = '{32'h46079247};
test_input[15384:15391] = '{32'hc2c457ac, 32'hc2015eeb, 32'hc282ec69, 32'h42954059, 32'hc2adf8e0, 32'h42837b51, 32'h42054c4d, 32'h422dc9cd};
test_weights[15384:15391] = '{32'hc285188e, 32'h4253d125, 32'h3fa96282, 32'hc28a0b60, 32'hc29f59be, 32'hc11d79e5, 32'hc297d8db, 32'hc2098010};
test_bias[1923:1923] = '{32'h40f05f91};
test_output[1923:1923] = '{32'h44e74ea9};
test_input[15392:15399] = '{32'hc0ce0d68, 32'h42ba2ac6, 32'hc2aa65f3, 32'h401fcda5, 32'h408e2bd6, 32'h41cf3853, 32'h426f28f0, 32'hc22135cd};
test_weights[15392:15399] = '{32'hc2992b86, 32'h41dbf305, 32'hc0188452, 32'hc1430311, 32'h4239420b, 32'h42840a22, 32'h410b1f35, 32'hc20bce31};
test_bias[1924:1924] = '{32'hc1babef8};
test_output[1924:1924] = '{32'h45dc2fb6};
test_input[15400:15407] = '{32'h40f47ab5, 32'h4031d685, 32'h428db4fa, 32'hc2460c8d, 32'hc296d3f4, 32'hc26f49d1, 32'h42b3a6b0, 32'hc20e00ce};
test_weights[15400:15407] = '{32'h401c28c0, 32'h429998a9, 32'hc28fb6d2, 32'h41f97600, 32'hc25ca666, 32'hc20d01fc, 32'hc2584a70, 32'h422507b3};
test_bias[1925:1925] = '{32'hc10d2fb6};
test_output[1925:1925] = '{32'hc5ca078d};
test_input[15408:15415] = '{32'h41b428b2, 32'h42ad3b09, 32'h42825396, 32'hc0a76a6d, 32'hc25ab558, 32'h425bfdc5, 32'h42b3fab4, 32'h4240fc62};
test_weights[15408:15415] = '{32'h426a52dd, 32'hc1daeccd, 32'h41b26d55, 32'h418b558d, 32'hc1182a1e, 32'hc29e08cc, 32'hc14ab951, 32'hc2963328};
test_bias[1926:1926] = '{32'h425e0be8};
test_output[1926:1926] = '{32'hc6007a47};
test_input[15416:15423] = '{32'h42232027, 32'hc199f563, 32'hc2bfd29d, 32'h40a44e5c, 32'hc0b25df5, 32'hc2bee7c5, 32'hc2706352, 32'h41e9d49c};
test_weights[15416:15423] = '{32'h40ca6aa5, 32'h4291dfec, 32'hc263432a, 32'h41a98364, 32'h425348ec, 32'hc1c6825b, 32'h41f1a60f, 32'h41864b09};
test_bias[1927:1927] = '{32'h424d317e};
test_output[1927:1927] = '{32'h45a2e8f1};
test_input[15424:15431] = '{32'h41af83a2, 32'hc2abee98, 32'hc29ed78a, 32'h41881132, 32'hc1c9512b, 32'h42bc4254, 32'h42c5d22b, 32'h425b16c7};
test_weights[15424:15431] = '{32'hc28f338a, 32'h42b9780e, 32'hc2454ff5, 32'h41853476, 32'hc1fdc48f, 32'h400173a1, 32'hc20b4f39, 32'hc24e48f4};
test_bias[1928:1928] = '{32'h418f36ca};
test_output[1928:1928] = '{32'hc625b3aa};
test_input[15432:15439] = '{32'hc1f8f259, 32'hc2733d1a, 32'h422cdec0, 32'h4237ba6e, 32'h412d1d77, 32'hc2ba6654, 32'h41de836e, 32'h423682a8};
test_weights[15432:15439] = '{32'hc227812a, 32'hc18d773a, 32'hc2bbca61, 32'h42ba7f91, 32'hc2495ff9, 32'h41d7e6ab, 32'hc23aad94, 32'hc2a8275b};
test_bias[1929:1929] = '{32'h4210bdc2};
test_output[1929:1929] = '{32'hc5ad9372};
test_input[15440:15447] = '{32'hc2ab868e, 32'h4176ecf2, 32'hc172fc0a, 32'hc2b6d1ca, 32'h41fbe5b0, 32'hc11864b8, 32'hc2abdc1e, 32'hc276e15b};
test_weights[15440:15447] = '{32'h42a5949d, 32'h428c9645, 32'h41501c17, 32'hc1dfb9b7, 32'h42bd2b59, 32'hc1bcd1a2, 32'h42a972a3, 32'hc26970f4};
test_bias[1930:1930] = '{32'h41eac7f0};
test_output[1930:1930] = '{32'hc5803538};
test_input[15448:15455] = '{32'h427a27e4, 32'hc2b844ca, 32'hc220df79, 32'h424d9b23, 32'h42b8157d, 32'hc0c56454, 32'hc2b6c384, 32'hc29b0329};
test_weights[15448:15455] = '{32'h42c3d1e1, 32'h42724111, 32'h427eddf6, 32'h41f5c061, 32'hc2103fc9, 32'hc1beb470, 32'hc2170f64, 32'h42c6bd48};
test_bias[1931:1931] = '{32'h40e42131};
test_output[1931:1931] = '{32'hc5f5815b};
test_input[15456:15463] = '{32'hc228caac, 32'h41d3e7a9, 32'h419f2674, 32'hc22d7d6d, 32'h4224d3af, 32'hc2bc4d16, 32'hc2354b8f, 32'h42897901};
test_weights[15456:15463] = '{32'h42786845, 32'hc209b99e, 32'h429d3074, 32'hc280417a, 32'hc2722e1a, 32'hc02e37df, 32'hc2769887, 32'h42026955};
test_bias[1932:1932] = '{32'h42b3a0fc};
test_output[1932:1932] = '{32'h45672c0f};
test_input[15464:15471] = '{32'h4273c4d6, 32'h4221a3bc, 32'hc24d0614, 32'hc2245d1c, 32'h42a021a8, 32'hc1382577, 32'hc22d3c89, 32'hc1fc1457};
test_weights[15464:15471] = '{32'hc103fe51, 32'h426c06d7, 32'hc1a19966, 32'hc2ae6de4, 32'hc211ca8f, 32'h429f5120, 32'h419ece0e, 32'hc29bd4e6};
test_bias[1933:1933] = '{32'h40fc7912};
test_output[1933:1933] = '{32'h458568a0};
test_input[15472:15479] = '{32'h419ff666, 32'h411ca691, 32'hc272fb25, 32'h425c249f, 32'h42a82576, 32'h42a22d5d, 32'h4254fcdd, 32'h428f9f22};
test_weights[15472:15479] = '{32'hc2acb4d6, 32'hc2c00001, 32'hc28f3eba, 32'h419363b0, 32'hc228c6d8, 32'hc2b4808f, 32'hc2a3397a, 32'hc1d90145};
test_bias[1934:1934] = '{32'h42695208};
test_output[1934:1934] = '{32'hc6610b2b};
test_input[15480:15487] = '{32'hc282407a, 32'h42288592, 32'hc2aaa345, 32'hc2c511d0, 32'h3fae5586, 32'hc0be88d0, 32'hc26464ae, 32'h41ba3cfd};
test_weights[15480:15487] = '{32'h426f9ccc, 32'hc1e0f7d8, 32'hc283a416, 32'hc25b34a9, 32'h3fb1019e, 32'h41c50d3e, 32'hc1a2ce6d, 32'hc28a187f};
test_bias[1935:1935] = '{32'h41ec9700};
test_output[1935:1935] = '{32'h45a7c7a2};
test_input[15488:15495] = '{32'hc22bdfd5, 32'h4242e250, 32'h42bfdb86, 32'hc28a9887, 32'h4294afd5, 32'hc1b270be, 32'hc2b9dd2d, 32'hc25ddc86};
test_weights[15488:15495] = '{32'h400ae0d5, 32'h412d5fe1, 32'hc2b375f8, 32'h424ff19e, 32'h4208f949, 32'h411d510c, 32'hc20b1fe7, 32'h4281e31b};
test_bias[1936:1936] = '{32'hc106c80f};
test_output[1936:1936] = '{32'hc6198d60};
test_input[15496:15503] = '{32'h42b46086, 32'h4283f755, 32'h42b2d0d8, 32'hc297d8f7, 32'h41e5f06b, 32'hc2c3f30d, 32'hc21a1e42, 32'hc0428b2b};
test_weights[15496:15503] = '{32'h42095ff8, 32'h42976278, 32'h41edc3c5, 32'h42771617, 32'h424b1838, 32'hbf13e883, 32'h42a2522b, 32'h41efde8a};
test_bias[1937:1937] = '{32'hc2628ae3};
test_output[1937:1937] = '{32'h45866209};
test_input[15504:15511] = '{32'h4237e747, 32'hc205de0e, 32'hc27ec441, 32'hc2ba13f7, 32'h41697105, 32'h4280f3cb, 32'h40b6800d, 32'hc2b2948c};
test_weights[15504:15511] = '{32'hc1a69829, 32'h41b27e0a, 32'h42c7d21f, 32'hc14847a7, 32'h4280f2b4, 32'hc269e1b3, 32'h4120ed7b, 32'hc2af2f89};
test_bias[1938:1938] = '{32'h42b4d5c0};
test_output[1938:1938] = '{32'hc4dc687b};
test_input[15512:15519] = '{32'hc28bbbbc, 32'hc1dbf2a0, 32'h42680b6a, 32'hc2222bf7, 32'hc1041c3d, 32'hc2af6dfa, 32'hc07b2b0b, 32'hc2b6ed1c};
test_weights[15512:15519] = '{32'hc225ff30, 32'h424fb726, 32'hc297cf87, 32'hc2a5a502, 32'hbec59e9a, 32'hc112207e, 32'hc2b7be28, 32'hc28bc46c};
test_bias[1939:1939] = '{32'hc2c3331d};
test_output[1939:1939] = '{32'h45f669b6};
test_input[15520:15527] = '{32'hc2b1cd6b, 32'hc2a7dbab, 32'hc2c2c3e6, 32'hc26e0620, 32'h41b12b43, 32'h41a08744, 32'h425deb10, 32'hc2c3be34};
test_weights[15520:15527] = '{32'h4264c364, 32'h413c1280, 32'h4262834b, 32'hbfe87eda, 32'hc2b039ec, 32'h42171133, 32'h42b2502b, 32'h42514909};
test_bias[1940:1940] = '{32'hc21de5a0};
test_output[1940:1940] = '{32'hc6495337};
test_input[15528:15535] = '{32'hc2870e72, 32'h422f2f91, 32'hc2c22a72, 32'h415d7618, 32'h428b24fc, 32'h42a0bb48, 32'h41199be0, 32'hc23e4e6d};
test_weights[15528:15535] = '{32'hc24af262, 32'hc2532d6f, 32'hc26b9d95, 32'h426fe28f, 32'h4280b7e0, 32'hc24663cb, 32'h42a4c7ef, 32'h40b2a933};
test_bias[1941:1941] = '{32'h4288a6f0};
test_output[1941:1941] = '{32'h4608afd5};
test_input[15536:15543] = '{32'h400f83f0, 32'hc28a0058, 32'h429848a3, 32'hc225955e, 32'hc24520dc, 32'h42a07937, 32'h42c6bd05, 32'hc2bfeb1e};
test_weights[15536:15543] = '{32'h41d48702, 32'hc2882b62, 32'hc1f5bede, 32'h42351315, 32'hc2a2b598, 32'h41dc88de, 32'h426be282, 32'h4225fac7};
test_bias[1942:1942] = '{32'hc2104e74};
test_output[1942:1942] = '{32'h46067f43};
test_input[15544:15551] = '{32'h41b6cc34, 32'hc1e2722e, 32'hc0872abf, 32'hc16a4c68, 32'h42beb8de, 32'hc2adeb50, 32'hc2883395, 32'hc20002ed};
test_weights[15544:15551] = '{32'h426c916d, 32'h41d0615c, 32'h42a0d522, 32'hc1d9757b, 32'h403e0c91, 32'h4271daa8, 32'h42be4121, 32'h41f017dc};
test_bias[1943:1943] = '{32'h41e50959};
test_output[1943:1943] = '{32'hc6370142};
test_input[15552:15559] = '{32'h42ac144a, 32'h41b7ef00, 32'h42be1a31, 32'hc256d168, 32'h41c5c6a1, 32'h41fd3187, 32'h411de0a3, 32'h42b1fdbc};
test_weights[15552:15559] = '{32'h42090689, 32'hc298d125, 32'hc28ea5b9, 32'hc118ebfd, 32'hc27f9c21, 32'h41558719, 32'hc2c4157b, 32'hc2550271};
test_bias[1944:1944] = '{32'hc2573c44};
test_output[1944:1944] = '{32'hc63b6558};
test_input[15560:15567] = '{32'h422f4dd9, 32'h41c3a17f, 32'h4211fe42, 32'h41d267cb, 32'hc1aad46c, 32'hc22757ff, 32'hc2c1d2ae, 32'hc18ab545};
test_weights[15560:15567] = '{32'h41d96457, 32'hc296d25a, 32'hc21b694a, 32'h41b4b60a, 32'h412542c5, 32'hc236177f, 32'hc22e6629, 32'hc115f60d};
test_bias[1945:1945] = '{32'h4241b1c2};
test_output[1945:1945] = '{32'h4591188b};
test_input[15568:15575] = '{32'hc1f37b2e, 32'h42aa8127, 32'hc2070deb, 32'h4225e943, 32'hc29da0c0, 32'h428e7c2a, 32'h4154716a, 32'hc188945b};
test_weights[15568:15575] = '{32'hc2127f11, 32'h42b3806f, 32'hc2405a7a, 32'hc2b29b4d, 32'hc204cac8, 32'h42a40184, 32'hc22b1988, 32'hc29f8763};
test_bias[1946:1946] = '{32'h4243f702};
test_output[1946:1946] = '{32'h4679cc1d};
test_input[15576:15583] = '{32'h42a693af, 32'hc28d79b6, 32'h42b8fdf6, 32'h4203d64a, 32'h41a2fe34, 32'hc097a15a, 32'hc25ffc9b, 32'hc1b25a16};
test_weights[15576:15583] = '{32'h428d6e03, 32'hc1101d3c, 32'hc0fb2ad4, 32'hc206281f, 32'hc2482bfb, 32'hc2be6355, 32'hc29caa73, 32'h429ce785};
test_bias[1947:1947] = '{32'hc1e554f1};
test_output[1947:1947] = '{32'h45d27d28};
test_input[15584:15591] = '{32'h41f3e40d, 32'h426734bb, 32'hc26e0077, 32'hc29f3556, 32'hc19adad7, 32'hc2b22c2c, 32'h42a93bdb, 32'hc0d90db5};
test_weights[15584:15591] = '{32'h426a8a20, 32'hc095eb5c, 32'hc2017827, 32'hc28f0a29, 32'h41540a57, 32'h426e031c, 32'hc0a0e4eb, 32'h42a6648c};
test_bias[1948:1948] = '{32'h4236ae14};
test_output[1948:1948] = '{32'h4524a63b};
test_input[15592:15599] = '{32'h4290dbff, 32'h4200b9a1, 32'h42bec4a1, 32'hc22c2735, 32'hc267bdbc, 32'h4281bfa4, 32'hc29db808, 32'hc2c60876};
test_weights[15592:15599] = '{32'h42a06790, 32'hc2904757, 32'hc225f6cc, 32'hc2ae28ba, 32'h42ba9f1f, 32'hc086985a, 32'h41041969, 32'h428368fc};
test_bias[1949:1949] = '{32'h418e20bc};
test_output[1949:1949] = '{32'hc6151190};
test_input[15600:15607] = '{32'h429a344c, 32'hc1821443, 32'h42368834, 32'hc29d5dd4, 32'hc2a355a1, 32'h410de44d, 32'hc2b226bb, 32'h428fb95b};
test_weights[15600:15607] = '{32'h41a4edb6, 32'hc2adc77b, 32'hc217ca8b, 32'h429b5811, 32'hc26f5364, 32'hc2b25b89, 32'h4252d2bd, 32'hc2c176f9};
test_bias[1950:1950] = '{32'hc190c1e9};
test_output[1950:1950] = '{32'hc641e6b0};
test_input[15608:15615] = '{32'hc22bed71, 32'hc12c61fa, 32'h422fd228, 32'h42bc3908, 32'h42b333cb, 32'hc2b0049b, 32'hc2212f6c, 32'h4296e251};
test_weights[15608:15615] = '{32'h42728954, 32'hc1e73a31, 32'h42447a3d, 32'hc1343329, 32'h4098072c, 32'hc1b2f2c3, 32'hc2246ff5, 32'hc2311022};
test_bias[1951:1951] = '{32'h42482cf4};
test_output[1951:1951] = '{32'hc3d91c9d};
test_input[15616:15623] = '{32'hc234b143, 32'h42ad6fc1, 32'hc278c0fc, 32'hc01d7d5a, 32'hc2917a83, 32'hc23090a1, 32'hbfbb923c, 32'h42ad8831};
test_weights[15616:15623] = '{32'h42b5775a, 32'hc2a2eeb9, 32'h4293dcec, 32'h40d66195, 32'h41588b7e, 32'hc18762d4, 32'hc2356ed3, 32'hc223731c};
test_bias[1952:1952] = '{32'hc215d268};
test_output[1952:1952] = '{32'hc69896c3};
test_input[15624:15631] = '{32'h42879c4c, 32'h42a7ff9f, 32'hc2851ad3, 32'hc170edd7, 32'hc1d3bf61, 32'h4106fd4b, 32'h4157d2b4, 32'hc1cf7ea6};
test_weights[15624:15631] = '{32'h422ee334, 32'h420c56cb, 32'h4194333a, 32'h4221d362, 32'h429bf55f, 32'h42984c58, 32'h419a53a3, 32'hc2ab0ace};
test_bias[1953:1953] = '{32'h42af6109};
test_output[1953:1953] = '{32'h45a2f0d9};
test_input[15632:15639] = '{32'hc262c461, 32'h42c4d64c, 32'h41ee6b32, 32'h41e50a50, 32'h4283f812, 32'hc14a9b48, 32'hc29ac185, 32'h42b8595d};
test_weights[15632:15639] = '{32'hc250a095, 32'hc1816176, 32'h4294a6b0, 32'h41b30d93, 32'h419eb3df, 32'h42836afd, 32'h420505a0, 32'hc065b193};
test_bias[1954:1954] = '{32'h424cf8b7};
test_output[1954:1954] = '{32'h44e6a4f3};
test_input[15640:15647] = '{32'h42c2077e, 32'h41a54a6b, 32'hc284b3bb, 32'h422daf13, 32'hc2275d10, 32'h416bfc93, 32'h42c5f0ba, 32'hc2bb03bc};
test_weights[15640:15647] = '{32'h424f17e5, 32'hc29d37fa, 32'hc18afdba, 32'hc1d804b5, 32'h42947f2f, 32'h41d472a6, 32'h41b318eb, 32'hc28973c8};
test_bias[1955:1955] = '{32'hc084b5cf};
test_output[1955:1955] = '{32'h46115781};
test_input[15648:15655] = '{32'h40e0ba68, 32'hc283bfb5, 32'hc2205fa6, 32'h42bdae61, 32'hc1ac1f99, 32'h4212b2e0, 32'h41976ede, 32'hc11cc615};
test_weights[15648:15655] = '{32'h41e95434, 32'h4277979b, 32'h42b82fdc, 32'hc1becc1d, 32'hc28a11f6, 32'hc24ba5f3, 32'h42b4d665, 32'h429e4f5a};
test_bias[1956:1956] = '{32'hc25d8f86};
test_output[1956:1956] = '{32'hc611c0e6};
test_input[15656:15663] = '{32'hc11ae685, 32'h413a63c5, 32'hc20b40e5, 32'hc1f63d1e, 32'h42b67bce, 32'hc247193c, 32'h42a66a29, 32'h4254cdc8};
test_weights[15656:15663] = '{32'h41d9fbcb, 32'h416cf36d, 32'h427593f3, 32'h4237cc9b, 32'hc01af7be, 32'hc2791861, 32'h417f5ce8, 32'hc1f2c069};
test_bias[1957:1957] = '{32'h4227af87};
test_output[1957:1957] = '{32'hc47c281e};
test_input[15664:15671] = '{32'h42c3b3fb, 32'h4290fa4a, 32'h42c08320, 32'hc0c45045, 32'h42aff079, 32'h414ba589, 32'h42c5472a, 32'hc0892c6e};
test_weights[15664:15671] = '{32'hc28d3dde, 32'h41e342f0, 32'h4262d314, 32'hc22bd447, 32'h41aace3d, 32'hc20975bc, 32'hc0ffc9e3, 32'hc122bb4a};
test_bias[1958:1958] = '{32'hc0143535};
test_output[1958:1958] = '{32'h44c38beb};
test_input[15672:15679] = '{32'h4148d6d2, 32'h42153071, 32'h41f67f5e, 32'h41962c11, 32'h424898bf, 32'hc2c2d9aa, 32'h42c40696, 32'hc1da2df8};
test_weights[15672:15679] = '{32'h42a2c1ea, 32'hc1eb410a, 32'h41b13106, 32'hc2510ceb, 32'hc2984cfd, 32'hc1dfb857, 32'hc265de83, 32'h42999b2a};
test_bias[1959:1959] = '{32'h42aaf1f5};
test_output[1959:1959] = '{32'hc60e57bc};
test_input[15680:15687] = '{32'hc29a3d53, 32'h4219e4cb, 32'hc246f373, 32'hc2a7eb1a, 32'h428fa14d, 32'h41a68adb, 32'hc29b7aae, 32'h42320141};
test_weights[15680:15687] = '{32'hc2c311f9, 32'hc2b2cb0c, 32'h4216f094, 32'hc293a669, 32'hc1b337fe, 32'hc1c5aaa9, 32'h429e1d0e, 32'h42ac81c3};
test_bias[1960:1960] = '{32'h425cb8f4};
test_output[1960:1960] = '{32'h457bc74d};
test_input[15688:15695] = '{32'hc2c62356, 32'h41c57b96, 32'hc1cda8b1, 32'h421e6f2c, 32'h4294a75a, 32'hc0f5dd94, 32'h41d8cf73, 32'hc2481345};
test_weights[15688:15695] = '{32'hc2b31049, 32'hc1266e3f, 32'h41bd096c, 32'hc27f7cd9, 32'h40271118, 32'h3f44d4e3, 32'hc2ace4f5, 32'h429e53f9};
test_bias[1961:1961] = '{32'hc29a8c6a};
test_output[1961:1961] = '{32'hc432fd1c};
test_input[15696:15703] = '{32'h425ce240, 32'h429fc238, 32'hc1cb0be0, 32'hc2688492, 32'hc23f8629, 32'hc1e7a466, 32'hc1c21657, 32'h4201ff43};
test_weights[15696:15703] = '{32'hc1badef0, 32'h41dae62b, 32'h42b26859, 32'hc232d86a, 32'hc1db225b, 32'hc298d262, 32'h40a43ded, 32'hc26489be};
test_bias[1962:1962] = '{32'h40ab037f};
test_output[1962:1962] = '{32'h452dacfb};
test_input[15704:15711] = '{32'hc0719d22, 32'h407bc35e, 32'hc2b220b8, 32'hc2288105, 32'hc19ea8bb, 32'h42852fc6, 32'h3fa48b1b, 32'hc2845efa};
test_weights[15704:15711] = '{32'hc20f2a62, 32'h4294e63c, 32'h421e771b, 32'h42a48391, 32'h42a6a010, 32'hc2c2d7bf, 32'h429addae, 32'hc291b9e0};
test_bias[1963:1963] = '{32'h4217d584};
test_output[1963:1963] = '{32'hc61845e6};
test_input[15712:15719] = '{32'hc264eff7, 32'hc2368895, 32'hc284a795, 32'hc12ca179, 32'h41a8f618, 32'h414b4a05, 32'hc1dde6c1, 32'hc20c24f4};
test_weights[15712:15719] = '{32'h4206400a, 32'hc251e29d, 32'h42b2af09, 32'h429a7e6f, 32'hc225e3e5, 32'h428fcbcc, 32'hc29263f8, 32'hc2a874a6};
test_bias[1964:1964] = '{32'h4241780a};
test_output[1964:1964] = '{32'hc4984fea};
test_input[15720:15727] = '{32'h3e01d906, 32'hc284bba5, 32'h4137b1e7, 32'hc2346354, 32'hc20d059d, 32'hc2b3e5cb, 32'h42a6012f, 32'h42b352a2};
test_weights[15720:15727] = '{32'hc292382a, 32'hc21a22b5, 32'h4081431e, 32'hc2a1111e, 32'h429c9fb5, 32'hc2b63dac, 32'h420553d7, 32'hc19de96b};
test_bias[1965:1965] = '{32'h42c520e2};
test_output[1965:1965] = '{32'h46475396};
test_input[15728:15735] = '{32'hc2c67391, 32'hc23c2f51, 32'hc2b1964f, 32'h41c84bb4, 32'h42a376aa, 32'hc176c55b, 32'h41376f06, 32'hc281e5b7};
test_weights[15728:15735] = '{32'h42bf8b5d, 32'h425dfa11, 32'h41d2e049, 32'h42a2b3f9, 32'h42ac2efd, 32'hc294251b, 32'hc2937cf2, 32'h40aa3480};
test_bias[1966:1966] = '{32'h420fa902};
test_output[1966:1966] = '{32'hc5a88de8};
test_input[15736:15743] = '{32'hc1c71fa0, 32'h420321bc, 32'hc2b04343, 32'h429ae5a4, 32'hc1f0cefe, 32'h41d9c806, 32'h41160b6f, 32'hc28f6a68};
test_weights[15736:15743] = '{32'h42c5e665, 32'h41996447, 32'hc29f048c, 32'hc2aa62c2, 32'hc2834307, 32'hc1f90018, 32'h42198cfd, 32'hc1d2568c};
test_bias[1967:1967] = '{32'h4254a380};
test_output[1967:1967] = '{32'h44fa3333};
test_input[15744:15751] = '{32'h41d08528, 32'hc2643aae, 32'hc263b6d3, 32'h4292a820, 32'hc2bf6a2c, 32'hc2bed115, 32'h41107381, 32'hc219d416};
test_weights[15744:15751] = '{32'h40ccdfed, 32'hc2b13b07, 32'h42a493e9, 32'hc20bb966, 32'h4236c2a4, 32'h42c428d0, 32'hc14ff4c3, 32'h41aba50c};
test_bias[1968:1968] = '{32'hc2a27363};
test_output[1968:1968] = '{32'hc6831260};
test_input[15752:15759] = '{32'hc22c9ef7, 32'h42c030d1, 32'h41dfecf5, 32'h4172fd09, 32'hc1b2e529, 32'h41c6ccf0, 32'hc2232c1c, 32'h4292a5a3};
test_weights[15752:15759] = '{32'hc2352ad4, 32'h42476a4e, 32'h42a2fda8, 32'h4207d86f, 32'hc1b4d98a, 32'hc295ef20, 32'hc2c2953c, 32'hc1da970f};
test_bias[1969:1969] = '{32'h429c2778};
test_output[1969:1969] = '{32'h461fd0b8};
test_input[15760:15767] = '{32'h4251acba, 32'h42c7267a, 32'hc2807966, 32'h426ec56d, 32'hc29f0a5f, 32'hc2b58279, 32'hc2915948, 32'hc149f20f};
test_weights[15760:15767] = '{32'h41927e57, 32'hc227ad41, 32'h4285d5c8, 32'hc13fab88, 32'hc1a5c19b, 32'hc1900cb7, 32'h42464df3, 32'h420189ee};
test_bias[1970:1970] = '{32'hc1ae779a};
test_output[1970:1970] = '{32'hc60c4e69};
test_input[15768:15775] = '{32'hc0ad2b1a, 32'hc2c420bf, 32'h406417a8, 32'hc2690c1a, 32'h41a93511, 32'h41dea9b2, 32'hc2192bfe, 32'hc2bb0f31};
test_weights[15768:15775] = '{32'hc26bc318, 32'hc2226d91, 32'hc2aff31c, 32'hc2931339, 32'h40176abe, 32'h413c09bb, 32'h415bf8b7, 32'hc2ad4a1b};
test_bias[1971:1971] = '{32'hc2449f76};
test_output[1971:1971] = '{32'h467cc542};
test_input[15776:15783] = '{32'hc1b999f6, 32'h42c536ee, 32'hc24f184d, 32'h41fab402, 32'h42b54f4d, 32'h42aa4d3c, 32'h41ca015c, 32'hc2b7da77};
test_weights[15776:15783] = '{32'hc2b3f748, 32'hc2b25228, 32'hc2885ac7, 32'h42bafe6f, 32'hc2244a78, 32'h422ca1fa, 32'hc2bda5f8, 32'hc23a37db};
test_bias[1972:1972] = '{32'h421891e3};
test_output[1972:1972] = '{32'h44cbcdad};
test_input[15784:15791] = '{32'hc2970527, 32'h4289d5e4, 32'h42b4be16, 32'hc201ccf5, 32'hc2a9554e, 32'h4266f472, 32'h412fea3e, 32'hc0c4b534};
test_weights[15784:15791] = '{32'h420d21a5, 32'h4219e8ec, 32'h422a689f, 32'h412eda67, 32'h3ffd7ff3, 32'h424dc938, 32'h42a36765, 32'hc24a407d};
test_bias[1973:1973] = '{32'hbff319be};
test_output[1973:1973] = '{32'h45ea277d};
test_input[15792:15799] = '{32'h428e4915, 32'h42bdd7ff, 32'hc2ba8999, 32'hc2a3370e, 32'h40f33bb4, 32'hc24584e4, 32'hc2bb0bae, 32'hc10673df};
test_weights[15792:15799] = '{32'h41bf6c84, 32'h42720677, 32'h42988a94, 32'h41037751, 32'h4290be48, 32'hc243de7f, 32'h42c5495c, 32'hc1b9bce9};
test_bias[1974:1974] = '{32'hc1e6c4f9};
test_output[1974:1974] = '{32'hc5c8eca9};
test_input[15800:15807] = '{32'h4296faa9, 32'hc17529dc, 32'hc22a6da9, 32'hc285b645, 32'hc1e68e8e, 32'h4127e793, 32'hc23bcd15, 32'h41663686};
test_weights[15800:15807] = '{32'h4234a147, 32'hbfe9fa8d, 32'h41ec1e68, 32'hc1145558, 32'hc0a7b6b7, 32'hc28a3b2a, 32'h426de730, 32'hc058d08d};
test_bias[1975:1975] = '{32'hc2426965};
test_output[1975:1975] = '{32'hc42633b1};
test_input[15808:15815] = '{32'hc2533108, 32'hc031f8e9, 32'h42708e03, 32'h42abefc4, 32'h41023d14, 32'h428e9d6a, 32'h428a6c88, 32'h429ee325};
test_weights[15808:15815] = '{32'hc2950046, 32'h41ef0ccd, 32'hc12af436, 32'hc1af377d, 32'h42466c93, 32'h41aaa7aa, 32'h42221916, 32'h427c4e24};
test_bias[1976:1976] = '{32'hc1ad7917};
test_output[1976:1976] = '{32'h462c8fcc};
test_input[15816:15823] = '{32'h42aca879, 32'hc2040f92, 32'hc2542e42, 32'hc2a44407, 32'hc2c54764, 32'h40c657af, 32'hc1b2ff92, 32'hc23137bd};
test_weights[15816:15823] = '{32'hc2b85f69, 32'hc22ce443, 32'hbf6dcc60, 32'hc1b5709c, 32'h4293a87c, 32'h40af02f8, 32'h42a06d11, 32'h42b60f9a};
test_bias[1977:1977] = '{32'hc1e68cd2};
test_output[1977:1977] = '{32'hc68a78f6};
test_input[15824:15831] = '{32'hc1bc3fad, 32'hc29c3b42, 32'h42b03c56, 32'h4293265b, 32'h428c6961, 32'hc2ad0c55, 32'hc297317e, 32'hc1e65bf3};
test_weights[15824:15831] = '{32'h4261f382, 32'hc26e9782, 32'hc22f8c30, 32'hc275aa07, 32'hc1c5c926, 32'hc20021f7, 32'hc2ab6c0f, 32'h410841d8};
test_bias[1978:1978] = '{32'h41e7e2fa};
test_output[1978:1978] = '{32'h450c37ce};
test_input[15832:15839] = '{32'h4226ecc3, 32'h42a38f21, 32'h41e628dc, 32'hc29bec14, 32'h420ebc13, 32'h4242e262, 32'hc0c14820, 32'h3f730a34};
test_weights[15832:15839] = '{32'h428b5c56, 32'h416b9075, 32'h428c5ba7, 32'h429a0b31, 32'h421d4a95, 32'hc24a4e18, 32'h42bc16cd, 32'h428d745f};
test_bias[1979:1979] = '{32'h4271f229};
test_output[1979:1979] = '{32'hc4abe491};
test_input[15840:15847] = '{32'h401d8bbd, 32'h42c01c81, 32'hc259a02e, 32'h424c7826, 32'hc2b118e5, 32'hc1db0fc7, 32'hc2c6c4d5, 32'h40e30b59};
test_weights[15840:15847] = '{32'h42ba1d9f, 32'h40b41b35, 32'hc163dbd7, 32'hc26bd4ac, 32'h4281dbe4, 32'hc2bc6665, 32'h4285a85f, 32'hc1ee45a8};
test_bias[1980:1980] = '{32'hc168673d};
test_output[1980:1980] = '{32'hc633cb33};
test_input[15848:15855] = '{32'h428fcfbf, 32'h417028ae, 32'h415b62a9, 32'hc14b666d, 32'h42008d64, 32'hc2512f06, 32'hc107c65a, 32'h415f2305};
test_weights[15848:15855] = '{32'hc26536df, 32'hc1ac1b4e, 32'hc13fff60, 32'h426ff3a2, 32'h419bb215, 32'hc211a495, 32'hc299aaf3, 32'h41e55a1e};
test_bias[1981:1981] = '{32'h3f33cda3};
test_output[1981:1981] = '{32'hc4df8bfd};
test_input[15856:15863] = '{32'hc285cf76, 32'h422d6931, 32'h42a006ef, 32'h42966433, 32'hc241f34c, 32'hc0e501bd, 32'hc2942093, 32'h42948841};
test_weights[15856:15863] = '{32'hc08294b9, 32'h41fd98b9, 32'hc202ea2b, 32'h4256b508, 32'h42b99570, 32'hc209cdcd, 32'h41a5e8df, 32'hc2900b87};
test_bias[1982:1982] = '{32'hc193eee3};
test_output[1982:1982] = '{32'hc5fcd9ad};
test_input[15864:15871] = '{32'hc10c0513, 32'h41b21171, 32'hc2570075, 32'hc2b41aa6, 32'hc284592a, 32'hc2a150aa, 32'h429748e7, 32'hc2bcb099};
test_weights[15864:15871] = '{32'hc1d1fcde, 32'hc20564ce, 32'h4274a58e, 32'h42190d3e, 32'h40805432, 32'hc1df0dce, 32'h41030ea5, 32'hc270e8d7};
test_bias[1983:1983] = '{32'h422bc25f};
test_output[1983:1983] = '{32'h44874f23};
test_input[15872:15879] = '{32'h421cefc4, 32'hc2924834, 32'hc24fee2b, 32'h428da3a2, 32'hc0095c18, 32'hc2744297, 32'hc14c4342, 32'h420e3a03};
test_weights[15872:15879] = '{32'hc2800312, 32'h42a219e1, 32'h41c8325d, 32'hc2a82f48, 32'hc1873c9a, 32'h41daf9a3, 32'hc28b5e19, 32'hc258e46c};
test_bias[1984:1984] = '{32'hc2935433};
test_output[1984:1984] = '{32'hc6901598};
test_input[15880:15887] = '{32'hc17c45a2, 32'h419a23f2, 32'hc28a5697, 32'h419c3a95, 32'h42b33505, 32'h416f16d4, 32'hc2b3e5a4, 32'hc1e10836};
test_weights[15880:15887] = '{32'hc1e88b20, 32'hc2c1a2b0, 32'h42aa0386, 32'h4101210e, 32'hc2c4d543, 32'hc15f35f6, 32'h4284b4c7, 32'hc2501860};
test_bias[1985:1985] = '{32'hc1b46153};
test_output[1985:1985] = '{32'hc6a197ad};
test_input[15888:15895] = '{32'h4282e17b, 32'h41d9d716, 32'hc229a551, 32'h41785bc9, 32'h41c3e6f6, 32'h4182ee20, 32'hc18b9aa6, 32'hc29ee4af};
test_weights[15888:15895] = '{32'hc29a5207, 32'hc0b20937, 32'h4242d444, 32'h42222143, 32'hc0c3f53f, 32'h429dab6b, 32'hc2a9c66a, 32'hc283566d};
test_bias[1986:1986] = '{32'hc089b85a};
test_output[1986:1986] = '{32'h44959fc2};
test_input[15896:15903] = '{32'hc24e5247, 32'hc260577b, 32'hc2878555, 32'hc2426cae, 32'h425f569e, 32'h4140cb3f, 32'hc1b92be0, 32'h41a637d8};
test_weights[15896:15903] = '{32'hc24f8ca8, 32'hc2398a8a, 32'h42c547fe, 32'h427d9f16, 32'hc1805027, 32'h42b67d36, 32'hc2a97590, 32'h429f1cd7};
test_bias[1987:1987] = '{32'h41b68a0c};
test_output[1987:1987] = '{32'hc421c141};
test_input[15904:15911] = '{32'hc140aa30, 32'hc2a9b36b, 32'h41d5144e, 32'hc281e09b, 32'h4289464c, 32'h4026b0a1, 32'h42b55522, 32'hc29a2344};
test_weights[15904:15911] = '{32'h4279d1c8, 32'hc1fd6133, 32'hc1978b59, 32'hc24f4c2d, 32'h4281d537, 32'h427b710c, 32'hc2651f98, 32'hc1dd4d50};
test_bias[1988:1988] = '{32'h42b2eebc};
test_output[1988:1988] = '{32'h45c95cd2};
test_input[15912:15919] = '{32'h42ad3e5d, 32'hc253bd5d, 32'h429c5b89, 32'hc2b945d5, 32'hc2a14bbb, 32'h41a4a8a0, 32'h4222c9df, 32'h4214eeae};
test_weights[15912:15919] = '{32'h42b963a9, 32'hc1b3433b, 32'hc23b4d0b, 32'h42a4dfee, 32'hc2c4c12f, 32'hc27a7230, 32'hc100e153, 32'h42bd7f13};
test_bias[1989:1989] = '{32'h41e4986e};
test_output[1989:1989] = '{32'h45f37ed5};
test_input[15920:15927] = '{32'hc2adace5, 32'hc201f9f5, 32'hc2b2f353, 32'h412809b0, 32'h4288179b, 32'hc290ad2a, 32'hc2b95ff8, 32'hc2275f3b};
test_weights[15920:15927] = '{32'hc237de95, 32'h42110758, 32'hc1f0ba62, 32'h4212ec89, 32'h425364f4, 32'hc1e6f706, 32'hc189e19e, 32'h42b5f198};
test_bias[1990:1990] = '{32'h4134d662};
test_output[1990:1990] = '{32'h46128a3b};
test_input[15928:15935] = '{32'hc2757c4c, 32'h41dd5b0c, 32'hc2669501, 32'h3fec2cff, 32'h426f69bc, 32'h41fccf82, 32'h42aa6c11, 32'hc1cf0389};
test_weights[15928:15935] = '{32'hc1910934, 32'h422a6d6e, 32'h426222b0, 32'hc1c9b0d4, 32'h428d8f88, 32'hc2911378, 32'h42561065, 32'hc23aef80};
test_bias[1991:1991] = '{32'h426a722b};
test_output[1991:1991] = '{32'h45d33295};
test_input[15936:15943] = '{32'h41b340f1, 32'hc2bc8d7b, 32'hc098c051, 32'hc272e3c2, 32'hbfcbdecf, 32'hc2b7876a, 32'hc2646f43, 32'h41aafe64};
test_weights[15936:15943] = '{32'h417f8feb, 32'hc2981e90, 32'h41955c45, 32'hc21d0ca7, 32'hc28377b8, 32'h4046581b, 32'hc29a3453, 32'h4279e2d5};
test_bias[1992:1992] = '{32'hc2a7c63a};
test_output[1992:1992] = '{32'h466f09a2};
test_input[15944:15951] = '{32'hc2559787, 32'h420b70f4, 32'h42395d81, 32'hc20b16b8, 32'hc26b8423, 32'h429da7d2, 32'hc292550e, 32'h428f5d38};
test_weights[15944:15951] = '{32'hc1e72250, 32'h42c3527d, 32'h41d31ffc, 32'hc257799e, 32'hc2690abd, 32'hc1908c3b, 32'hc217dedd, 32'h4299f638};
test_bias[1993:1993] = '{32'h42988804};
test_output[1993:1993] = '{32'h468feb81};
test_input[15952:15959] = '{32'h4218abaa, 32'h419e0660, 32'h42c0383f, 32'h42999c4c, 32'h419d251e, 32'hc2b7a018, 32'hc20a9535, 32'h416b26f1};
test_weights[15952:15959] = '{32'h42b38e55, 32'h424731c5, 32'h41eea873, 32'h42a982d5, 32'hc25699fd, 32'hc2058724, 32'h428daebd, 32'hc2b2648d};
test_bias[1994:1994] = '{32'h4247e9cb};
test_output[1994:1994] = '{32'h463ccb80};
test_input[15960:15967] = '{32'h4233363c, 32'hc2bc9ebd, 32'hc239923e, 32'h410dd2fe, 32'hc28008ba, 32'h41d54e47, 32'h41dd197b, 32'h4295a181};
test_weights[15960:15967] = '{32'hc18ad914, 32'hc1fd2bdf, 32'h41bf99c9, 32'h42a2eeb8, 32'h428b9608, 32'h418f0bfb, 32'h42abec78, 32'h42c47bfd};
test_bias[1995:1995] = '{32'hc2c2f2f2};
test_output[1995:1995] = '{32'h45e8f8f6};
test_input[15968:15975] = '{32'hc28df168, 32'h427bbe74, 32'hc2508aa7, 32'hc1e889d5, 32'h4209d397, 32'hc24d4751, 32'hbf8d819a, 32'h4154f324};
test_weights[15968:15975] = '{32'hc19fc38e, 32'h40fa2421, 32'h41923de5, 32'h4210b978, 32'hc27f1e87, 32'hc11525bb, 32'h42a9bccf, 32'h42b29fcc};
test_bias[1996:1996] = '{32'h423f0fd0};
test_output[1996:1996] = '{32'hc4280396};
test_input[15976:15983] = '{32'hc2a0e2ed, 32'hc24cf10d, 32'h3f90fe43, 32'h429275af, 32'hc2334f20, 32'hc13fd6d6, 32'h4182cc51, 32'h42886fa2};
test_weights[15976:15983] = '{32'h42388a1a, 32'h42a8bedd, 32'h4282fb77, 32'h4298de72, 32'h429c9c20, 32'h42be7ad0, 32'hc2607d06, 32'hc298ba09};
test_bias[1997:1997] = '{32'h42c715d0};
test_output[1997:1997] = '{32'hc64bc89f};
test_input[15984:15991] = '{32'hc0c25910, 32'hc2905cee, 32'hc2614529, 32'hc2ab62b7, 32'hbf04f36f, 32'hc232e508, 32'hc210db9e, 32'hc13d2e9a};
test_weights[15984:15991] = '{32'h41816980, 32'h4238dd6a, 32'h429ccf9b, 32'hc26f6a3d, 32'hc24c2f85, 32'hc28df856, 32'h4296db1e, 32'h42c6228c};
test_bias[1998:1998] = '{32'hc29a6ca7};
test_output[1998:1998] = '{32'hc55abb51};
test_input[15992:15999] = '{32'h42169622, 32'hc20b7de6, 32'hc02b9229, 32'h404c3529, 32'h42b04493, 32'h42199838, 32'hc24c4e78, 32'hc1ef93f3};
test_weights[15992:15999] = '{32'hc2b22006, 32'hc2391466, 32'h42c22398, 32'h427f3033, 32'hc1473482, 32'h4232b05f, 32'h42adc870, 32'hc2899976};
test_bias[1999:1999] = '{32'hc1744f06};
test_output[1999:1999] = '{32'hc55f2f8c};
test_input[16000:16007] = '{32'h4288c404, 32'hc20956db, 32'hc1cbf8b8, 32'hc2835a43, 32'h4266f3ab, 32'h428bf0d7, 32'hc08e7461, 32'hbfaf2a03};
test_weights[16000:16007] = '{32'h429905a7, 32'h41ee1187, 32'h413b1568, 32'h40c61bb2, 32'h4271d1e1, 32'h42a2bbaa, 32'hc234a186, 32'h40c65d0c};
test_bias[2000:2000] = '{32'h429f5a27};
test_output[2000:2000] = '{32'h464a865a};
test_input[16008:16015] = '{32'hc2be6dae, 32'hc2853a2f, 32'h4292ebb7, 32'hc0dc114f, 32'h41f16c8b, 32'hc197baeb, 32'hc18bb41e, 32'hc2a9a661};
test_weights[16008:16015] = '{32'hc2b93fcd, 32'hc2997b89, 32'h42abd9a9, 32'hc2994c37, 32'h40a8ad44, 32'h427a0546, 32'hc284dbd3, 32'hc1200803};
test_bias[2001:2001] = '{32'h4202b4a2};
test_output[2001:2001] = '{32'h46aa3247};
test_input[16016:16023] = '{32'hc1a330aa, 32'hc284756d, 32'hc1a6dbd4, 32'hc2488e70, 32'hc21fd38b, 32'h424d8390, 32'hc1257cf7, 32'hc2b89347};
test_weights[16016:16023] = '{32'hc192faf7, 32'hc23082a8, 32'h41032b65, 32'hc0ecb331, 32'h41e1c269, 32'h42af5989, 32'h40e84524, 32'h40af7cd3};
test_bias[2002:2002] = '{32'h424215e4};
test_output[2002:2002] = '{32'h45c62c97};
test_input[16024:16031] = '{32'h41e4d363, 32'h4277913c, 32'h41e597f4, 32'hc265d53d, 32'hc004b8de, 32'h41394b2c, 32'hc1b6ca84, 32'h42a27471};
test_weights[16024:16031] = '{32'h4233035d, 32'hc25bf59a, 32'h42692138, 32'hc2150144, 32'hc2ac15a0, 32'h41d3cfb9, 32'hc2b5c60a, 32'hc1d5bf1e};
test_bias[2003:2003] = '{32'h42b68bde};
test_output[2003:2003] = '{32'h4507c715};
test_input[16032:16039] = '{32'hc22ceca2, 32'hc10573ab, 32'h42266bd0, 32'h425b8fc3, 32'h42744b31, 32'hc24d41dd, 32'h418e6df8, 32'hc28a44ed};
test_weights[16032:16039] = '{32'h426cac2d, 32'h4290c5ee, 32'h426ef16d, 32'hc2bf7dbc, 32'hc2a806d2, 32'h42c43199, 32'h421e9193, 32'h41b821a7};
test_bias[2004:2004] = '{32'h42af3a23};
test_output[2004:2004] = '{32'hc683fce5};
test_input[16040:16047] = '{32'h4295695a, 32'h42c401de, 32'hc244127d, 32'h416f54ee, 32'h427a4a77, 32'h428a7b7f, 32'h427f9081, 32'h42488534};
test_weights[16040:16047] = '{32'h3f8a5bf6, 32'hc22a7a99, 32'hc1c9b02d, 32'h42aea390, 32'h41913fe2, 32'h411001c3, 32'h3fdf0137, 32'h42bc979f};
test_bias[2005:2005] = '{32'hc1917e8f};
test_output[2005:2005] = '{32'h459d0a48};
test_input[16048:16055] = '{32'hc2a948ce, 32'h41e7582f, 32'hc23764ee, 32'h419f269d, 32'hc14b18a3, 32'h408ff0d4, 32'hbe58e9cd, 32'h42c5476a};
test_weights[16048:16055] = '{32'hc225d1d7, 32'h42bb09cb, 32'hc27cae5b, 32'h424b44a2, 32'h4278d2f4, 32'h429ac05b, 32'hc2a1d400, 32'h41808fd6};
test_bias[2006:2006] = '{32'h4244160c};
test_output[2006:2006] = '{32'h463108c8};
test_input[16056:16063] = '{32'h4231331e, 32'h4140bdf5, 32'hc2bd035b, 32'hc297137a, 32'hc240f1b2, 32'h42113cd7, 32'h42ba343f, 32'hc115c7fb};
test_weights[16056:16063] = '{32'h4250bd8d, 32'h41b714a7, 32'h42afacc8, 32'hc29e2d89, 32'hc28c04c4, 32'hc1257b69, 32'h429ca08d, 32'h42a4fb01};
test_bias[2007:2007] = '{32'hc19f7d97};
test_output[2007:2007] = '{32'h461883b0};
test_input[16064:16071] = '{32'h4293c266, 32'h42541d40, 32'hc2231729, 32'hc1fcb855, 32'h42051f23, 32'h41d5b31a, 32'hc08fc7e7, 32'h42b1098e};
test_weights[16064:16071] = '{32'hc0ee2c30, 32'h4237fa80, 32'h429bc40e, 32'hc2b78fa0, 32'hc22aed3b, 32'h427f2450, 32'hbfa8a8f3, 32'h42a0a0ce};
test_bias[2008:2008] = '{32'hc28c90be};
test_output[2008:2008] = '{32'h460baeb6};
test_input[16072:16079] = '{32'h429d4499, 32'h427a2268, 32'h42860224, 32'hc265b33a, 32'hc163a9e5, 32'h426c386a, 32'hc26660f7, 32'hc1f821e6};
test_weights[16072:16079] = '{32'h41d5e568, 32'hc114ea1e, 32'hc27e8dda, 32'h42b66975, 32'h3e978e6c, 32'h42a96df3, 32'hc280d429, 32'h42027d37};
test_bias[2009:2009] = '{32'hc20b6436};
test_output[2009:2009] = '{32'hc39fa040};
test_input[16080:16087] = '{32'h4201d210, 32'hc258bcd3, 32'hc1b78555, 32'hc188286d, 32'h421509b0, 32'h423f92cc, 32'hc173a153, 32'h42a0a757};
test_weights[16080:16087] = '{32'h4217ab30, 32'h42182e98, 32'h42001240, 32'h428b021f, 32'h41cb911d, 32'hc26433e7, 32'hc1f1ccc6, 32'h425554f4};
test_bias[2010:2010] = '{32'h42971b78};
test_output[2010:2010] = '{32'h438fa6e5};
test_input[16088:16095] = '{32'hc18c908d, 32'h3e5ea484, 32'hc274406a, 32'h3fec7d1d, 32'h423a4290, 32'hc0e507ec, 32'h414e67d2, 32'hc1002c71};
test_weights[16088:16095] = '{32'h42994507, 32'h41bb5e04, 32'hc29953a9, 32'h4158dd0e, 32'h400f4606, 32'h41f500c1, 32'h40c27680, 32'hc25fcc0e};
test_bias[2011:2011] = '{32'hc2a2c0e7};
test_output[2011:2011] = '{32'h4566f2ce};
test_input[16096:16103] = '{32'h42834f6e, 32'h42962207, 32'hc1895158, 32'hc1dbfb7d, 32'h42b8a8a5, 32'hc28227c6, 32'hc249c1dc, 32'hc2996518};
test_weights[16096:16103] = '{32'h41017fc8, 32'h428f80ef, 32'h423087cb, 32'h415ba9a7, 32'hc1523cd8, 32'h41eb1a0f, 32'h3e836850, 32'hc2aad89b};
test_bias[2012:2012] = '{32'hc2236d21};
test_output[2012:2012] = '{32'h45fed612};
test_input[16104:16111] = '{32'h42972cf8, 32'h42a3a940, 32'h4218e045, 32'hc26a8722, 32'hc242f7a6, 32'hc20eb97b, 32'h4275c1a1, 32'hc2973262};
test_weights[16104:16111] = '{32'h4285bf4d, 32'h428b4950, 32'hc2b5df33, 32'h4248f9cf, 32'h424631df, 32'hbfebe90a, 32'hc13e8701, 32'h42667b95};
test_bias[2013:2013] = '{32'h42969fbf};
test_output[2013:2013] = '{32'hc53d546b};
test_input[16112:16119] = '{32'h4213d2c5, 32'h42991be9, 32'hc2b0c122, 32'hc2bfd932, 32'hc12c57a8, 32'hc29b8c5c, 32'hc26fd122, 32'h420e16b7};
test_weights[16112:16119] = '{32'hc2665d15, 32'hc2c40a7d, 32'hc2beebe9, 32'hc2683edc, 32'hc0f51eb7, 32'h4272395a, 32'h42619f3d, 32'h425aa036};
test_bias[2014:2014] = '{32'hc19a6210};
test_output[2014:2014] = '{32'hc4d61c99};
test_input[16120:16127] = '{32'hc1cbb7e6, 32'h427ea08a, 32'h41a7ad71, 32'h428a4906, 32'hc2c35f8e, 32'h41c1524b, 32'hc1b5a06c, 32'hc20c27ed};
test_weights[16120:16127] = '{32'hc247f08d, 32'h4096fd50, 32'hc215b57c, 32'h42830429, 32'h42859169, 32'h4216549e, 32'hc2b19f68, 32'hc2865dba};
test_bias[2015:2015] = '{32'hc1ddc088};
test_output[2015:2015] = '{32'h457cd103};
test_input[16128:16135] = '{32'hc2880f85, 32'h4264469f, 32'hc23d8425, 32'h42aed35b, 32'h42a590b3, 32'hc2103702, 32'hc1f874ad, 32'hc1fa4a6d};
test_weights[16128:16135] = '{32'hc2a91486, 32'hc2bf4164, 32'h42a8e86c, 32'h423aeac4, 32'h4283a06f, 32'h4215dc37, 32'h421e287a, 32'h41dca943};
test_bias[2016:2016] = '{32'h42892be0};
test_output[2016:2016] = '{32'h45194654};
test_input[16136:16143] = '{32'h42806de5, 32'hc21bc1db, 32'h4160424f, 32'h42023f0f, 32'hc2a4d0a0, 32'h429e6814, 32'hc0b53126, 32'h4278d4a2};
test_weights[16136:16143] = '{32'hc1aab882, 32'h41619f53, 32'h418907c8, 32'h429e04ab, 32'hc1dc6a10, 32'h40c558ef, 32'hbfeaa8bb, 32'hc289d9c3};
test_bias[2017:2017] = '{32'h4033b407};
test_output[2017:2017] = '{32'hc41b9127};
test_input[16144:16151] = '{32'h42c01a68, 32'hc21b63f5, 32'hc1bddb5d, 32'h40e2d728, 32'hc2a023f0, 32'h422f4a52, 32'hc1379e5f, 32'h41d17daa};
test_weights[16144:16151] = '{32'hc19bfddf, 32'hc29b656e, 32'h427f0c75, 32'hc2ad96b1, 32'h41e4dc4c, 32'hc28b1048, 32'hc2257038, 32'hc2babe52};
test_bias[2018:2018] = '{32'h42ae3b23};
test_output[2018:2018] = '{32'hc6002fe2};
test_input[16152:16159] = '{32'hc24a1099, 32'hc101d59a, 32'h4221cf26, 32'hc2809972, 32'hc23d0b49, 32'h429eaac9, 32'hc2717963, 32'h42a53775};
test_weights[16152:16159] = '{32'h41db2900, 32'hc0cbba02, 32'hc1518d30, 32'hc289b372, 32'hc1348f67, 32'h428c278d, 32'hc11bdcf7, 32'hc0ac14c8};
test_bias[2019:2019] = '{32'hc2bc1971};
test_output[2019:2019] = '{32'h46080e98};
test_input[16160:16167] = '{32'h428935ab, 32'h42302b13, 32'hc1b41a57, 32'hc13dadf4, 32'hc28a2b16, 32'h42bb0f2a, 32'h4229f14e, 32'h42b1e045};
test_weights[16160:16167] = '{32'hc22d84cb, 32'hc2bf8217, 32'hc2addf1f, 32'h429875cc, 32'hc2712eb4, 32'h42711b73, 32'hc0cd170b, 32'h422ae15c};
test_bias[2020:2020] = '{32'h428b106f};
test_output[2020:2020] = '{32'h45e2e02b};
test_input[16168:16175] = '{32'hc20aeee5, 32'h42aab892, 32'h42b46525, 32'h41442a50, 32'hc282d916, 32'h418bca25, 32'hc2bb050e, 32'h42b788fa};
test_weights[16168:16175] = '{32'hc2ae01c0, 32'h4288c0fb, 32'h40aba793, 32'hc2b80739, 32'h40dfac14, 32'hc2bbc430, 32'h40fd9a2a, 32'h42781581};
test_bias[2021:2021] = '{32'hc1dce1e8};
test_output[2021:2021] = '{32'h462c7d75};
test_input[16176:16183] = '{32'hc26b9272, 32'h42489842, 32'h41de20df, 32'hc2112582, 32'h42afc3df, 32'h4287617d, 32'h4272cb46, 32'h414a9258};
test_weights[16176:16183] = '{32'hc2495bd1, 32'h41c3d74f, 32'hc29c7cda, 32'h41c1b3da, 32'h3fad5bc8, 32'h42220da6, 32'hc287ed3a, 32'h42ad74be};
test_bias[2022:2022] = '{32'h42b666d4};
test_output[2022:2022] = '{32'h4485510d};
test_input[16184:16191] = '{32'hc1b822a4, 32'h40d468de, 32'h40fa46ca, 32'h4225cf9c, 32'hc2ba8712, 32'hc114e121, 32'hc2b0917d, 32'h422a74d2};
test_weights[16184:16191] = '{32'hc2c757cc, 32'h4290f101, 32'h42864bd5, 32'hc285acff, 32'h4076dcb8, 32'hc25a2828, 32'hc2aa1017, 32'hc2ae7aad};
test_bias[2023:2023] = '{32'h410a782b};
test_output[2023:2023] = '{32'h458bdb71};
test_input[16192:16199] = '{32'h41941118, 32'h41a2d68a, 32'hc0b07a62, 32'h421a4543, 32'hbf105671, 32'h42227605, 32'hc20cfeaa, 32'hc200a493};
test_weights[16192:16199] = '{32'h42aeaa05, 32'hc27ae49c, 32'h42a2b07f, 32'h4297d85c, 32'hc2850f22, 32'hbff18619, 32'h41398924, 32'hc2822788};
test_bias[2024:2024] = '{32'h419c1165};
test_output[2024:2024] = '{32'h458c1e24};
test_input[16200:16207] = '{32'h420baf09, 32'hc23e58f5, 32'h426b8cec, 32'h423a98a0, 32'h41ee99bc, 32'h414cc323, 32'hc284180a, 32'hc2c74aca};
test_weights[16200:16207] = '{32'h428924b0, 32'h42a34a34, 32'hc23b9fdc, 32'hc0ba12f3, 32'h42134926, 32'hc16eb699, 32'hc2c379e4, 32'h4214d2d6};
test_bias[2025:2025] = '{32'hc2a3a31d};
test_output[2025:2025] = '{32'hc46db07b};
test_input[16208:16215] = '{32'h40af58db, 32'h41d17dfc, 32'h42a72c49, 32'h41146d37, 32'h42684f8b, 32'h42177ab8, 32'hc162f28f, 32'h4260d04d};
test_weights[16208:16215] = '{32'hc0f1fbed, 32'hc1d570b7, 32'h41ba742e, 32'h3f930b10, 32'hc2c7505b, 32'h4295866c, 32'hc16276f9, 32'h428e0a70};
test_bias[2026:2026] = '{32'hc14ca5b8};
test_output[2026:2026] = '{32'h45189a78};
test_input[16216:16223] = '{32'h428760f3, 32'h411e04bd, 32'hc0a759b8, 32'h42c12f51, 32'h42a86d46, 32'h40028f09, 32'h427dca10, 32'h425aaa5b};
test_weights[16216:16223] = '{32'h422d1f82, 32'h42955b30, 32'h42565082, 32'h428ed78e, 32'hc1547375, 32'hc22332ed, 32'h429e3661, 32'h414ff7d5};
test_bias[2027:2027] = '{32'h42a2b939};
test_output[2027:2027] = '{32'h4668bd12};
test_input[16224:16231] = '{32'hc2a4557c, 32'hc28a88cb, 32'hc2aa3f93, 32'h4293bb15, 32'h42827047, 32'hc298697f, 32'hc2c09c53, 32'hc205ec0f};
test_weights[16224:16231] = '{32'h4108bb98, 32'hc2ba8533, 32'h4287bafe, 32'h420ccba9, 32'h4189ea4f, 32'hc252c299, 32'hc2bb1b9d, 32'hc2253a3c};
test_bias[2028:2028] = '{32'h41f13abd};
test_output[2028:2028] = '{32'h468dbe6a};
test_input[16232:16239] = '{32'h4199d2b9, 32'h42264542, 32'hc25d17d1, 32'hc29f9914, 32'h41b8b298, 32'hc2b7b10f, 32'h429402e5, 32'hc2ba1f88};
test_weights[16232:16239] = '{32'hc0cbd87d, 32'hc1f80fa0, 32'h42878f98, 32'h42a1be18, 32'hc283c509, 32'hc1308006, 32'hc288ee26, 32'h41dee308};
test_bias[2029:2029] = '{32'hc26cc194};
test_output[2029:2029] = '{32'hc69afbf8};
test_input[16240:16247] = '{32'hc22c84f0, 32'hc2b474f8, 32'h429697cf, 32'hc1412f66, 32'hc2ab8041, 32'hc2836ece, 32'h41d5a790, 32'hc0a5d0a5};
test_weights[16240:16247] = '{32'h420088ae, 32'h4157e1ad, 32'hc2bd1495, 32'h42369879, 32'hc28977f5, 32'h42a379fe, 32'hc1e73b9b, 32'h42a5675d};
test_bias[2030:2030] = '{32'hc29fc838};
test_output[2030:2030] = '{32'hc62c5bd0};
test_input[16248:16255] = '{32'h41b106b5, 32'hc1f55867, 32'h42b4d2c8, 32'h42a46128, 32'hc22a843d, 32'h41f66edd, 32'hc0138668, 32'h4168704d};
test_weights[16248:16255] = '{32'h4220d2af, 32'h4168f3a8, 32'h42b2cae0, 32'h416ba67a, 32'hc22d9682, 32'h429d4590, 32'h4291a84f, 32'hc20e6b46};
test_bias[2031:2031] = '{32'h428d247a};
test_output[2031:2031] = '{32'h4651477f};
test_input[16256:16263] = '{32'hc21c21e6, 32'hc24bb7d6, 32'hc2aa6c84, 32'h42b82029, 32'hc00fd598, 32'hc169295c, 32'h42692325, 32'h41150091};
test_weights[16256:16263] = '{32'hc201cc5c, 32'h42bea6c7, 32'hc1f4961f, 32'hc0cb7222, 32'hc2ab7d63, 32'h42264998, 32'h41acee69, 32'h41a25472};
test_bias[2032:2032] = '{32'h4258b213};
test_output[2032:2032] = '{32'hc3ef39e6};
test_input[16264:16271] = '{32'h41f28dd7, 32'h427843d8, 32'h42015eaa, 32'hc1c18e17, 32'hc22c0384, 32'hc29f0fee, 32'h428508b1, 32'hc26d9347};
test_weights[16264:16271] = '{32'hc2610dbe, 32'hc1e07b35, 32'hc2767a76, 32'hc2ad19d2, 32'h42be41b9, 32'hc0f19ec9, 32'hc25eba13, 32'h408725a8};
test_bias[2033:2033] = '{32'h41baac0d};
test_output[2033:2033] = '{32'hc6283fe2};
test_input[16272:16279] = '{32'hc2277a95, 32'h4274b6eb, 32'hc2bc6a61, 32'h42bd246b, 32'h42960e84, 32'h42bbcfc6, 32'hc0ae84cf, 32'h3e54250b};
test_weights[16272:16279] = '{32'h426cf14c, 32'h4243219b, 32'h41584209, 32'hc0e093ba, 32'hc042df43, 32'h4202d75b, 32'hc1bc0fe8, 32'h429a6f8d};
test_bias[2034:2034] = '{32'hc2a3c339};
test_output[2034:2034] = '{32'h44b81a1e};
test_input[16280:16287] = '{32'hc284522b, 32'hc284870b, 32'hc2688908, 32'hc2b6773b, 32'h42bd73e9, 32'hc287d341, 32'hc0bf05c0, 32'hc2a9a1db};
test_weights[16280:16287] = '{32'hc2bb7ea8, 32'h42ad8420, 32'h42322264, 32'h4204fbf8, 32'h41a0eda5, 32'hc14e81c8, 32'h42aa81f1, 32'h42b0e864};
test_bias[2035:2035] = '{32'hc1920687};
test_output[2035:2035] = '{32'hc622c01a};
test_input[16288:16295] = '{32'hc1e01c81, 32'h429b95fb, 32'hc2b155d8, 32'h41fdf29b, 32'h41f18a42, 32'h42b3058d, 32'h42442797, 32'h4100cc86};
test_weights[16288:16295] = '{32'h429fa070, 32'h429718e6, 32'h4223987b, 32'hc2ac51ff, 32'h427ce76e, 32'h425f13e1, 32'hc2abf670, 32'hc18eec3e};
test_bias[2036:2036] = '{32'hc29c0b39};
test_output[2036:2036] = '{32'hc380bf4c};
test_input[16296:16303] = '{32'h4201ca85, 32'h4100a999, 32'h4224c474, 32'hc18fbb6e, 32'h40bdfbb1, 32'h426e9d23, 32'h42109226, 32'h426a5249};
test_weights[16296:16303] = '{32'h42bca521, 32'h421e8962, 32'hc2179ee7, 32'h42775161, 32'h41200335, 32'hc2612490, 32'h41bf2b9f, 32'hc2990bd4};
test_bias[2037:2037] = '{32'h41e4d13e};
test_output[2037:2037] = '{32'hc5c12dab};
test_input[16304:16311] = '{32'hc1f92512, 32'h41644683, 32'h423b0698, 32'h42b3b976, 32'h428aaca8, 32'h42c0e798, 32'h40061dcb, 32'h42441930};
test_weights[16304:16311] = '{32'hc24bf185, 32'h422a2ec5, 32'hc1c1c0ae, 32'hc191f9dd, 32'hc219bb72, 32'hc23e8fe7, 32'h423c7236, 32'h401518f3};
test_bias[2038:2038] = '{32'h415f516c};
test_output[2038:2038] = '{32'hc5edd1e5};
test_input[16312:16319] = '{32'hc1b8d8f6, 32'h425a30f1, 32'hc27a71cf, 32'hc2b23720, 32'h42a71df7, 32'h42a4b173, 32'hc2aaf04d, 32'hc1005000};
test_weights[16312:16319] = '{32'hbf97f5df, 32'h425acc72, 32'hc29c6106, 32'h42722f47, 32'h41a60f6d, 32'h42a08f58, 32'hc21b8cdb, 32'hc2c2f5eb};
test_bias[2039:2039] = '{32'h42abaae9};
test_output[2039:2039] = '{32'h466b206d};
test_input[16320:16327] = '{32'h42ac2e29, 32'h4205d267, 32'hc15726d5, 32'hc27981ae, 32'h419536fb, 32'h42502245, 32'h409a9fc1, 32'hc2b1bd4a};
test_weights[16320:16327] = '{32'h4269b963, 32'hc25f6dc7, 32'hc2ad996d, 32'hc23b82f8, 32'h419cef75, 32'hc154b961, 32'h42199774, 32'hc287f749};
test_bias[2040:2040] = '{32'hc13b68a0};
test_output[2040:2040] = '{32'h464d59bc};
test_input[16328:16335] = '{32'h42b68965, 32'h4250fcf3, 32'h418a06a2, 32'hc2aca526, 32'hc261373b, 32'hc1bca315, 32'hc28de321, 32'h409d5dc4};
test_weights[16328:16335] = '{32'hc0c87daa, 32'hc253f583, 32'h41d0012a, 32'h4269209b, 32'hc2b192d3, 32'hbece5319, 32'h4206bb42, 32'h41855ce8};
test_bias[2041:2041] = '{32'h410bb559};
test_output[2041:2041] = '{32'hc5a2e93c};
test_input[16336:16343] = '{32'h42597e28, 32'h428369ba, 32'h424b15ce, 32'h426a0ef3, 32'hc250eca8, 32'hc1e92a69, 32'h41e60e01, 32'hc28aae90};
test_weights[16336:16343] = '{32'hc299d185, 32'h4211113b, 32'h42139193, 32'hc20b3b45, 32'h41cb9d0a, 32'h41e63733, 32'h4293b439, 32'hc245fd24};
test_bias[2042:2042] = '{32'hc20b5582};
test_output[2042:2042] = '{32'h44adcede};
test_input[16344:16351] = '{32'hc2902546, 32'hc205076f, 32'hc2c7e94d, 32'hc20b29b1, 32'hc27111e8, 32'hc29bccb9, 32'h42437ddd, 32'hc2b48f9c};
test_weights[16344:16351] = '{32'h41990ca4, 32'h42afaa0f, 32'h426ea023, 32'hc1d3de9d, 32'hc2c72a56, 32'h4231ab80, 32'h42297a1c, 32'h4220b310};
test_bias[2043:2043] = '{32'hc2a12d1a};
test_output[2043:2043] = '{32'hc603d39c};
test_input[16352:16359] = '{32'h42bec723, 32'hc2b16a65, 32'h419486b9, 32'h4222621f, 32'hc2b91c8f, 32'h4298f03d, 32'hc2a0b620, 32'hc103d513};
test_weights[16352:16359] = '{32'hc295e9ad, 32'h418ea336, 32'hc23dc848, 32'hc24df9cf, 32'hc2b72d18, 32'hc21a4bb9, 32'hc299e721, 32'hc138e44b};
test_bias[2044:2044] = '{32'hc25f02bf};
test_output[2044:2044] = '{32'h423d237f};
test_input[16360:16367] = '{32'h42504914, 32'h4130c7c0, 32'h42997c6b, 32'h42980ec3, 32'h42840302, 32'hc2946e3a, 32'hc23f2f6b, 32'hc1e4e3e0};
test_weights[16360:16367] = '{32'h42b790bf, 32'h42bffc5a, 32'hc1bfc43c, 32'hc18d4f04, 32'hc1e2af9e, 32'h4197ce4c, 32'h42c72717, 32'h41ea6338};
test_bias[2045:2045] = '{32'hc273f6c0};
test_output[2045:2045] = '{32'hc5c43f78};
test_input[16368:16375] = '{32'h42c2e9bb, 32'h42908851, 32'hc1d7e220, 32'h42973cdd, 32'h42985783, 32'h4291102c, 32'h4263f0c3, 32'hc10715f4};
test_weights[16368:16375] = '{32'h42942ee3, 32'h4125f996, 32'h42a40206, 32'hc28c8039, 32'h42c2fd89, 32'hc204b508, 32'hc28eb9fb, 32'h425aaaeb};
test_bias[2046:2046] = '{32'h4176df45};
test_output[2046:2046] = '{32'h446e1711};
test_input[16376:16383] = '{32'h42b5e29b, 32'h40f07f83, 32'hc216dd1f, 32'h422bd9a2, 32'hc0225c5e, 32'h4156d21c, 32'hc1e5c5f8, 32'h42209eb1};
test_weights[16376:16383] = '{32'h41fc031f, 32'h4295b381, 32'h41c20ba6, 32'h425a5202, 32'hc29b5f23, 32'hc014cb96, 32'h429beb63, 32'h411f8833};
test_bias[2047:2047] = '{32'hc0fd98fe};
test_output[2047:2047] = '{32'h45468a11};
test_input[16384:16391] = '{32'hc282ebe0, 32'hc26ff4c2, 32'hc29a9c76, 32'h42486d06, 32'hc1d2bd92, 32'hc18d1a94, 32'h42bc1291, 32'h4016e327};
test_weights[16384:16391] = '{32'h4232f0dd, 32'h421a4610, 32'hc2733940, 32'hc24f8e1a, 32'h42403f86, 32'hc2b81762, 32'h429e5c61, 32'h42ae3210};
test_bias[2048:2048] = '{32'h4284d791};
test_output[2048:2048] = '{32'h459a2ce3};
test_input[16392:16399] = '{32'hc2a5eb22, 32'h422376d4, 32'hc145b562, 32'h426fac8f, 32'h42b48e47, 32'h42579abf, 32'hc2844e04, 32'h427d4e73};
test_weights[16392:16399] = '{32'hc29afb16, 32'h3fb54bf0, 32'h4232d8f6, 32'h42927972, 32'h425b3e7e, 32'hc090fbf4, 32'h424ab7d6, 32'h41ed357f};
test_bias[2049:2049] = '{32'hc236df0e};
test_output[2049:2049] = '{32'h4653067e};
test_input[16400:16407] = '{32'hc1057232, 32'hc1b11ecb, 32'hc0834cea, 32'h42803a76, 32'hc2bc587f, 32'h4212f927, 32'hc298314c, 32'h4282adea};
test_weights[16400:16407] = '{32'h40a5ebaf, 32'hc0f3e5fc, 32'hc2940a56, 32'hc28db12f, 32'h42065507, 32'h409fcff7, 32'hc02b922f, 32'hc27c1efb};
test_bias[2050:2050] = '{32'h423392fc};
test_output[2050:2050] = '{32'hc62b4674};
test_input[16408:16415] = '{32'h403e0a7e, 32'h41e1222c, 32'h421759ab, 32'h410c0b9d, 32'hc2443519, 32'h4210ea8b, 32'h41dc8747, 32'h42161416};
test_weights[16408:16415] = '{32'hc2b9f076, 32'hc293d4c3, 32'h42843ab5, 32'h42892edc, 32'h40d363b6, 32'h42ae6e45, 32'h4224df8f, 32'h419d1833};
test_bias[2051:2051] = '{32'hc2bcc13c};
test_output[2051:2051] = '{32'h45a78107};
test_input[16416:16423] = '{32'h4255cabe, 32'hbfc66846, 32'h42c0f338, 32'hc2c3e92c, 32'h425851a6, 32'h41dffa4a, 32'h42b092f9, 32'hc20ae595};
test_weights[16416:16423] = '{32'h422d26fe, 32'hc2a1dc7b, 32'hc26723bd, 32'hc273927a, 32'h425e89bc, 32'h429060ea, 32'h419649c7, 32'h4279b80b};
test_bias[2052:2052] = '{32'h42bae8f4};
test_output[2052:2052] = '{32'h45e898d5};
test_input[16424:16431] = '{32'h424f21d7, 32'hc26975ef, 32'hc1a53dd3, 32'hc246b766, 32'h42733ebc, 32'hc19d0b93, 32'h41d3ee45, 32'h4220c83c};
test_weights[16424:16431] = '{32'h42c315ea, 32'hc2bdec6e, 32'h4263c0ee, 32'hc263dbb4, 32'h413838dd, 32'hc13629be, 32'h4227ff3f, 32'hc04b8f7d};
test_bias[2053:2053] = '{32'h42a0dd53};
test_output[2053:2053] = '{32'h465e7117};
test_input[16432:16439] = '{32'h4115cbcc, 32'h42489317, 32'h42a01570, 32'hc1ad3e61, 32'hc2700b1a, 32'h4293e966, 32'h4225131f, 32'h42b2c27d};
test_weights[16432:16439] = '{32'h417bb8ff, 32'hc1f2e91b, 32'h41e99d8b, 32'hc20f9615, 32'hc2c60da5, 32'hc122f9ac, 32'h421026f7, 32'hc19a37c9};
test_bias[2054:2054] = '{32'hc25d0291};
test_output[2054:2054] = '{32'h45cf6ea1};
test_input[16440:16447] = '{32'hc23d1748, 32'hc217ceb9, 32'hc23d3ecf, 32'hc1f4a93d, 32'h4289ba33, 32'hc234867f, 32'h40b99fcd, 32'hc2b7359d};
test_weights[16440:16447] = '{32'hc244a05e, 32'hc1c43b78, 32'hc2ba2c8e, 32'hc2312338, 32'h4171aead, 32'hc1e67f8e, 32'hc137c80c, 32'hc280add3};
test_bias[2055:2055] = '{32'hc2a7cc68};
test_output[2055:2055] = '{32'h468591cd};
test_input[16448:16455] = '{32'h419aa890, 32'h42250405, 32'h41e67d2e, 32'h422f3972, 32'hc12d9855, 32'hc1fad5d2, 32'h40bc3c61, 32'hc2901427};
test_weights[16448:16455] = '{32'h42b5f69c, 32'h42a16b84, 32'h4213cc19, 32'h42b2dd51, 32'hc218e283, 32'hc0d1dbd5, 32'hc21a8759, 32'h42099a6b};
test_bias[2056:2056] = '{32'h424c7ede};
test_output[2056:2056] = '{32'h45fb2591};
test_input[16456:16463] = '{32'h420b1ce2, 32'h3fdd96b8, 32'h420cfe66, 32'h3e221289, 32'h420ef670, 32'h4209ea6c, 32'hc24eecee, 32'h426d55a7};
test_weights[16456:16463] = '{32'hc2b2a747, 32'hc24c65dc, 32'h4271db78, 32'h41a6f4d0, 32'h42907abd, 32'hc288f770, 32'h4011d896, 32'hc24816fd};
test_bias[2057:2057] = '{32'hc1931d5b};
test_output[2057:2057] = '{32'hc5768226};
test_input[16464:16471] = '{32'h4145babb, 32'h41e85b5f, 32'hc2b5cac0, 32'h41c4ea0d, 32'hc24fbeb7, 32'hc21c261c, 32'hc2b64481, 32'hc2814412};
test_weights[16464:16471] = '{32'hc2b7e3f5, 32'h4019c064, 32'h4136fada, 32'hc2334f17, 32'h41574618, 32'h4296134e, 32'hc0cb49c8, 32'h419d0a99};
test_bias[2058:2058] = '{32'hc2bfac30};
test_output[2058:2058] = '{32'hc5ee389e};
test_input[16472:16479] = '{32'h42061432, 32'hc1e54049, 32'hc29d7c7a, 32'h41bf4f4f, 32'hc272703a, 32'h42263256, 32'h41c90aec, 32'hc23f5854};
test_weights[16472:16479] = '{32'h429aaf7f, 32'hc135664c, 32'hc299861e, 32'h402c6139, 32'hc26d5fda, 32'h40be270d, 32'hc1d92d99, 32'hc02737b6};
test_bias[2059:2059] = '{32'hc1b00adc};
test_output[2059:2059] = '{32'h46400aee};
test_input[16480:16487] = '{32'hc28f9b43, 32'hc1613035, 32'h41ca6c17, 32'h41f997b9, 32'h4290c967, 32'hc2afff9b, 32'hc2a1f03d, 32'h4289778d};
test_weights[16480:16487] = '{32'h42a24e57, 32'hc1c121e1, 32'hc2a2f973, 32'h428c06ba, 32'h418cef11, 32'h42bae6e4, 32'h42c5b82e, 32'h41ec3809};
test_bias[2060:2060] = '{32'h42a7e96a};
test_output[2060:2060] = '{32'hc68e385c};
test_input[16488:16495] = '{32'hc1c88122, 32'hc291bada, 32'h4237ea8c, 32'hc2a2e4b6, 32'hc11a006d, 32'hc1b0fae9, 32'h424d7373, 32'hc28325e5};
test_weights[16488:16495] = '{32'hc1b6534f, 32'hc108023b, 32'h428bd813, 32'hc2a6bdd1, 32'hc15e2171, 32'hc2707dc0, 32'h41e47c19, 32'h429231ed};
test_bias[2061:2061] = '{32'hc2aae59d};
test_output[2061:2061] = '{32'h46107edb};
test_input[16496:16503] = '{32'h42bf9ede, 32'hc2938d14, 32'h4209a2f6, 32'h4231b5cb, 32'h4298d2b1, 32'hc27fb7f1, 32'hc26a078b, 32'hc2253bd9};
test_weights[16496:16503] = '{32'hc29db38c, 32'h42117a0b, 32'h42b35f07, 32'hc2a7a9c0, 32'hc22f260b, 32'hc2bc821f, 32'hc114fbca, 32'h426438ea};
test_bias[2062:2062] = '{32'h4200e943};
test_output[2062:2062] = '{32'hc61be16d};
test_input[16504:16511] = '{32'hc2afc47f, 32'h42472fa5, 32'h41a35428, 32'h42c3e9e6, 32'hc2a38c11, 32'h42800909, 32'hc0263432, 32'h4294289f};
test_weights[16504:16511] = '{32'hc1e492d7, 32'hc2507e3d, 32'hc2aaa12e, 32'h418bcf15, 32'hc2bd9970, 32'hc201c4a2, 32'h4262ba83, 32'h4293398e};
test_bias[2063:2063] = '{32'h42c4cb4b};
test_output[2063:2063] = '{32'h462b5492};
test_input[16512:16519] = '{32'h413a2c87, 32'hc1e391b4, 32'hc2be18d1, 32'h42bbdde6, 32'h42c1b15d, 32'h42b836db, 32'h42a8c991, 32'hc263936e};
test_weights[16512:16519] = '{32'h41eeb52f, 32'h429bb394, 32'h42808c98, 32'h4297a63c, 32'h422bdef2, 32'h42510a1e, 32'hc069cce4, 32'hc1caaf3b};
test_bias[2064:2064] = '{32'h3fb38310};
test_output[2064:2064] = '{32'h46109ceb};
test_input[16520:16527] = '{32'hc29cda20, 32'h428613c4, 32'hc2c2be47, 32'h429f7548, 32'hc2c07542, 32'h3f546bcd, 32'hc23ab05f, 32'h410f9258};
test_weights[16520:16527] = '{32'h3e9bd389, 32'hc2584e2c, 32'h42645291, 32'hc2528435, 32'hc1b40b21, 32'h41a858a5, 32'hc26b8bdd, 32'h427514e2};
test_bias[2065:2065] = '{32'h41c3c8c6};
test_output[2065:2065] = '{32'hc5f6cb3a};
test_input[16528:16535] = '{32'hc2b57c64, 32'hc1a413fc, 32'hc292fe21, 32'hc25a2b20, 32'hc287453e, 32'h42384479, 32'hc1891d2e, 32'h41ea4dbf};
test_weights[16528:16535] = '{32'hc29e58dd, 32'h422909bc, 32'h420b223d, 32'hc11e4d88, 32'hc0e991f2, 32'h4231fc3c, 32'h42ac293f, 32'h42a01ebb};
test_bias[2066:2066] = '{32'hc2c3754d};
test_output[2066:2066] = '{32'h45ee00a4};
test_input[16536:16543] = '{32'h41fd9e07, 32'h424eeffe, 32'hc2afb7cc, 32'hc280c3c7, 32'h42b3a8e9, 32'hc260a30b, 32'hbfe925ba, 32'h4135ebda};
test_weights[16536:16543] = '{32'hc2a73ebb, 32'hc2922338, 32'h41565555, 32'hc18fb7b1, 32'h423cda76, 32'h411dfdc0, 32'h42036613, 32'h413eb90f};
test_bias[2067:2067] = '{32'h4227f44a};
test_output[2067:2067] = '{32'hc5257339};
test_input[16544:16551] = '{32'h42212cc5, 32'h42c00fa2, 32'h42b99ba8, 32'hc1961049, 32'hc1c7a129, 32'h4218a799, 32'hc1fb157f, 32'h42b26664};
test_weights[16544:16551] = '{32'hc2a9bd85, 32'hc201e77d, 32'h4277b4a5, 32'h429a38f5, 32'h4269ba8c, 32'hc286c4fb, 32'h4297c5be, 32'h426ea36c};
test_bias[2068:2068] = '{32'hc1adc71d};
test_output[2068:2068] = '{32'hc55156b0};
test_input[16552:16559] = '{32'hc27621db, 32'hc1b169e1, 32'h41e53666, 32'hc26bf740, 32'hc2877e39, 32'h42aaa13f, 32'h429cbb0f, 32'h41cd22d4};
test_weights[16552:16559] = '{32'h42421a16, 32'h40a71bbe, 32'h42832a85, 32'hc19e71eb, 32'hc0904db6, 32'h4196ef00, 32'hc2c4634e, 32'hc20b6115};
test_bias[2069:2069] = '{32'h42abeaff};
test_output[2069:2069] = '{32'hc5cf8dde};
test_input[16560:16567] = '{32'h419383a4, 32'hc261704a, 32'h421f8f14, 32'hc1d38411, 32'h42a10313, 32'h4297ddd9, 32'hc1ef1a82, 32'h42799011};
test_weights[16560:16567] = '{32'h42c032b4, 32'hc2b07f6e, 32'h42b89d3b, 32'hc24d5fcd, 32'hc2c421e6, 32'hc2becb75, 32'h42926820, 32'h41b094b7};
test_bias[2070:2070] = '{32'hc2ab6614};
test_output[2070:2070] = '{32'hc584cf9d};
test_input[16568:16575] = '{32'hc28d0834, 32'h42634059, 32'hc21665c2, 32'h4285bf06, 32'hc2b00c54, 32'h42c5bc04, 32'h40dbfe86, 32'hc27b12dd};
test_weights[16568:16575] = '{32'hbfe54aee, 32'h40565990, 32'h426cba56, 32'hc18f15e9, 32'h42a95d26, 32'h421321b8, 32'h42757631, 32'h411b8e64};
test_bias[2071:2071] = '{32'h42489361};
test_output[2071:2071] = '{32'hc5dca2ac};
test_input[16576:16583] = '{32'hc2a15d65, 32'hc1fd8114, 32'hc20da56a, 32'hc2af42ec, 32'h424bb301, 32'h426c2409, 32'hc2bb7c33, 32'hc159fc8e};
test_weights[16576:16583] = '{32'hc250eb4d, 32'h42816ad2, 32'h42b796c3, 32'h428855b1, 32'h4250963d, 32'h42c4cac9, 32'h422eaedb, 32'h40844953};
test_bias[2072:2072] = '{32'hc06b7c00};
test_output[2072:2072] = '{32'hc52be051};
test_input[16584:16591] = '{32'hc0e93ebf, 32'h422cb327, 32'h404b1aba, 32'hc23bc3ef, 32'hc2886c69, 32'hc2367a78, 32'h4298ed01, 32'h421d27e2};
test_weights[16584:16591] = '{32'h41949aa0, 32'h42b07822, 32'h42894cbd, 32'hc1823399, 32'h42c21013, 32'h41e9ef3d, 32'hc2bdba66, 32'h3e1a6ff0};
test_bias[2073:2073] = '{32'hc09178ed};
test_output[2073:2073] = '{32'hc624d3a4};
test_input[16592:16599] = '{32'h42abc245, 32'hc26cb1ec, 32'hc20634c1, 32'hc2a42e8e, 32'h427cc65d, 32'h428c894e, 32'hc214ec9e, 32'h424da9c7};
test_weights[16592:16599] = '{32'hc2956777, 32'h42ab8904, 32'hc1ce3c99, 32'h429ddbde, 32'h42b23cb2, 32'h425f4b50, 32'hc2acc624, 32'h41f83766};
test_bias[2074:2074] = '{32'h41da2efd};
test_output[2074:2074] = '{32'hc5297d2e};
test_input[16600:16607] = '{32'h422e5c14, 32'h42092e84, 32'hc2903bb3, 32'hc0c4c6e4, 32'hc216ba91, 32'h42637413, 32'hc2250e30, 32'hc15ef083};
test_weights[16600:16607] = '{32'hc2b4ebc9, 32'hc292f92f, 32'h40ec832f, 32'h42a9daf6, 32'h41b3cef0, 32'hc245898f, 32'h4226e175, 32'h42b32d63};
test_bias[2075:2075] = '{32'h4230afb5};
test_output[2075:2075] = '{32'hc65c4dd1};
test_input[16608:16615] = '{32'hc1f9156e, 32'h42ad8e6f, 32'hc20961a7, 32'hc2a5dfdb, 32'hc26f368e, 32'h4234dd9d, 32'hc19a2136, 32'h41e1804e};
test_weights[16608:16615] = '{32'h40fb0a4d, 32'hc278981c, 32'h42c69583, 32'hc2376b84, 32'hc267e8c3, 32'hc22dd0cf, 32'hc2abd4c2, 32'hc2163fb8};
test_bias[2076:2076] = '{32'h4242bce2};
test_output[2076:2076] = '{32'hc5418f7a};
test_input[16616:16623] = '{32'hc21c8fe7, 32'hc2806964, 32'h420cd1fd, 32'hc2be96d3, 32'hc2b09e17, 32'h40e3f200, 32'hc2a1e892, 32'h4226afa4};
test_weights[16616:16623] = '{32'hc209be37, 32'h42a37d30, 32'h42c6ab09, 32'h42811747, 32'h41428595, 32'h40a28b13, 32'h42a9f318, 32'hc29c6fef};
test_bias[2077:2077] = '{32'h428ece25};
test_output[2077:2077] = '{32'hc689f604};
test_input[16624:16631] = '{32'hc28dcd1b, 32'h41f2d044, 32'h42304678, 32'h427c3c21, 32'h419531dc, 32'h422185c0, 32'hc21ba35f, 32'hc22650e1};
test_weights[16624:16631] = '{32'hc2950084, 32'h42a0c7be, 32'hc210fd5f, 32'hc2c121fe, 32'hc2c12270, 32'h425376d5, 32'hc2911310, 32'hbe6e9725};
test_bias[2078:2078] = '{32'hc29b805c};
test_output[2078:2078] = '{32'h45433951};
test_input[16632:16639] = '{32'h424f341f, 32'h42a8ab07, 32'hc2b33fd2, 32'h423314af, 32'hc28ac61d, 32'hc0ad37cf, 32'hc0eb3828, 32'hc2af0988};
test_weights[16632:16639] = '{32'h42a25287, 32'h42c1998e, 32'hc2a64688, 32'hc1b09e10, 32'hc2b71ba1, 32'h42c67056, 32'h4280a2af, 32'hc267d805};
test_bias[2079:2079] = '{32'h422efe0f};
test_output[2079:2079] = '{32'h46e4d37f};
test_input[16640:16647] = '{32'hc2b0f5c4, 32'hc1f87d69, 32'hc2aacdc7, 32'hc21a7805, 32'h42178f59, 32'hc2366195, 32'hc2c68fbd, 32'hc28b32a3};
test_weights[16640:16647] = '{32'hc268675f, 32'h414a6d28, 32'h4144f023, 32'hc22c1a07, 32'h4281dea0, 32'h42705550, 32'h413496f7, 32'h41f916a6};
test_bias[2080:2080] = '{32'hc28ab5ea};
test_output[2080:2080] = '{32'h44d7415e};
test_input[16648:16655] = '{32'h42ad1929, 32'h426fb5c7, 32'h42856845, 32'h4231699d, 32'hc29a98a1, 32'hc2466481, 32'h41aff520, 32'h420c562a};
test_weights[16648:16655] = '{32'h42a43f14, 32'hc18056e9, 32'hc20d9605, 32'hc24c3e28, 32'h4211c5f5, 32'hc24fa948, 32'h42bac9a7, 32'h426aa60d};
test_bias[2081:2081] = '{32'h421a6e81};
test_output[2081:2081] = '{32'h45a9aa96};
test_input[16656:16663] = '{32'hc140c9d9, 32'hc2be8287, 32'hc297509c, 32'hc2382a67, 32'hc1be1d35, 32'h40cd4889, 32'hc1e701eb, 32'h4247490c};
test_weights[16656:16663] = '{32'hc28af44b, 32'hc222fd9c, 32'hc27a1c9c, 32'h3f9da531, 32'h421ccfe7, 32'h42851cbc, 32'hc2350615, 32'hc1f4f70e};
test_bias[2082:2082] = '{32'h4225ebea};
test_output[2082:2082] = '{32'h46081a81};
test_input[16664:16671] = '{32'h428de640, 32'h416eba27, 32'h42839ae7, 32'h4219a262, 32'h4283f524, 32'h427cd9ee, 32'h40da023e, 32'h42608b26};
test_weights[16664:16671] = '{32'hc1ec7d7a, 32'hc10834bf, 32'h41b52df2, 32'h42174b69, 32'hc2b3c41a, 32'hc2a7c507, 32'h429de407, 32'h41258473};
test_bias[2083:2083] = '{32'h41771fd7};
test_output[2083:2083] = '{32'hc612915a};
test_input[16672:16679] = '{32'h42330391, 32'hc21149b1, 32'hc10d11ae, 32'h42c417b4, 32'hc1472573, 32'hc21dd354, 32'hc1b0e04a, 32'hc21d431a};
test_weights[16672:16679] = '{32'hc23551e5, 32'hc2767ee6, 32'h42aa2a5e, 32'hc29502e0, 32'h41cda0e6, 32'h4291efe6, 32'hc26eeaad, 32'hc1e29f0f};
test_bias[2084:2084] = '{32'h4287640f};
test_output[2084:2084] = '{32'hc6057a21};
test_input[16680:16687] = '{32'h4284c31c, 32'h42c54a1b, 32'h42c2c353, 32'h426c5199, 32'h42c588ef, 32'h4296545b, 32'h4235abbb, 32'hc2987a70};
test_weights[16680:16687] = '{32'hc22f1f7f, 32'hc2284bae, 32'h41fb879c, 32'h4288f9c6, 32'h42aa0c63, 32'hc2488ec2, 32'hc2a01645, 32'h413690b9};
test_bias[2085:2085] = '{32'hc26ff4d1};
test_output[2085:2085] = '{32'h42e61ea7};
test_input[16688:16695] = '{32'hc20a7241, 32'h41704395, 32'hc09d4cc5, 32'h42c5f906, 32'hc2a42474, 32'hc294711e, 32'hc2c66ccf, 32'hc1341745};
test_weights[16688:16695] = '{32'hc2aa7b83, 32'hc2c7d8e7, 32'h4206a699, 32'hc25bb91d, 32'hc2262bf4, 32'h42b5f075, 32'hc1cb56a7, 32'h428913ba};
test_bias[2086:2086] = '{32'h424b42db};
test_output[2086:2086] = '{32'hc5b1f2a9};
test_input[16696:16703] = '{32'h4251415e, 32'hc2162051, 32'hc2be9eae, 32'hc27e7d5a, 32'h4118c4f8, 32'h415980d9, 32'h42953408, 32'h42a5612b};
test_weights[16696:16703] = '{32'h42349dbb, 32'h42c1a064, 32'hc18b068b, 32'hc2945d1d, 32'h427f957f, 32'h42447ce2, 32'h42926744, 32'h4208d0c7};
test_bias[2087:2087] = '{32'h3f368030};
test_output[2087:2087] = '{32'h466541a1};
test_input[16704:16711] = '{32'h42a145cb, 32'hc186797e, 32'h42683216, 32'hc2092bca, 32'h4210f618, 32'h42ba2473, 32'h42bcfdfb, 32'hc2a00181};
test_weights[16704:16711] = '{32'hc2673a85, 32'h42a479a9, 32'hc28c71e5, 32'h42769c2e, 32'h4203f2fd, 32'h4184dc23, 32'hc240869b, 32'hc2bda4b8};
test_bias[2088:2088] = '{32'hc2b245cf};
test_output[2088:2088] = '{32'hc5cc83ea};
test_input[16712:16719] = '{32'h427e1ea1, 32'h40cb78e4, 32'hc25f4b3d, 32'h3ffce28a, 32'h42a98ab2, 32'h42bb9913, 32'hc2c0ac2a, 32'h422742cf};
test_weights[16712:16719] = '{32'hc236b9c8, 32'h42bd5909, 32'h412d361b, 32'h4244abda, 32'hc18750cc, 32'hc2c1e0c2, 32'hc244adbb, 32'hc1130d71};
test_bias[2089:2089] = '{32'h4253278a};
test_output[2089:2089] = '{32'hc60b82b5};
test_input[16720:16727] = '{32'hc1941ffd, 32'hc1cee5ae, 32'h429d1d94, 32'h42bdfaa1, 32'hc2887d77, 32'hc1147da6, 32'h42a706df, 32'h4206c92a};
test_weights[16720:16727] = '{32'h4275949c, 32'hc18e9f4c, 32'h421310ae, 32'hbfbbcba4, 32'h41403d5d, 32'hc1c4aed7, 32'hc155aa53, 32'hc2c59607};
test_bias[2090:2090] = '{32'hc28a872b};
test_output[2090:2090] = '{32'hc53d8116};
test_input[16728:16735] = '{32'h42a8b746, 32'h429be10f, 32'hc27b43e5, 32'h42c5bc0a, 32'hc2b67392, 32'h419d495c, 32'hc1e72123, 32'hc2714de1};
test_weights[16728:16735] = '{32'hc18b2de4, 32'hc0b6667b, 32'h429faa93, 32'h42818771, 32'h4238a5a3, 32'h42b30897, 32'h4285af2a, 32'hc29d82f0};
test_bias[2091:2091] = '{32'h40dbc04e};
test_output[2091:2091] = '{32'hc3140558};
test_input[16736:16743] = '{32'h42654159, 32'hc2b03754, 32'h41dba271, 32'h41ef9007, 32'hc21abf27, 32'h41272c33, 32'h4244b8b2, 32'hc2afddb2};
test_weights[16736:16743] = '{32'hbfd9894a, 32'h422301dd, 32'h41806bb2, 32'hc20e24c3, 32'h42a4bf63, 32'h429660d3, 32'h426d27b0, 32'hc245e9ef};
test_bias[2092:2092] = '{32'h421bc5c3};
test_output[2092:2092] = '{32'h441440e5};
test_input[16744:16751] = '{32'hc27b124a, 32'hc2a8ed2c, 32'h41aa2766, 32'h4282ec4c, 32'h42abe540, 32'hc2114821, 32'hc23fb24f, 32'h422dcb60};
test_weights[16744:16751] = '{32'h42b96be4, 32'h4216c034, 32'h42c3f814, 32'h4297bb35, 32'h41396dbd, 32'hc2689381, 32'hc2a5f3d6, 32'h408d5865};
test_bias[2093:2093] = '{32'hc2b126e3};
test_output[2093:2093] = '{32'h45a39d35};
test_input[16752:16759] = '{32'hc1dac45c, 32'hc1bf8c8c, 32'hc2a8a27d, 32'h428bb0b0, 32'h420e997a, 32'hc21e02c8, 32'h423033db, 32'hc261e857};
test_weights[16752:16759] = '{32'h4242608a, 32'hc271c162, 32'hc1c00e3b, 32'hc23f4513, 32'hc282ef15, 32'h41f392eb, 32'h4140f8ae, 32'h42ac2905};
test_bias[2094:2094] = '{32'h4283ffab};
test_output[2094:2094] = '{32'hc60c98db};
test_input[16760:16767] = '{32'h42ac1c9a, 32'hc276b9a1, 32'h4206e038, 32'h4209dc8d, 32'h425d9fd7, 32'h42c4a57a, 32'h42a64e8c, 32'hc2af3813};
test_weights[16760:16767] = '{32'h41a87657, 32'hc2c2562a, 32'hc2c3c664, 32'h42bfdb0b, 32'h40c192eb, 32'h42c716c0, 32'h425bc69b, 32'h42b049fe};
test_bias[2095:2095] = '{32'hc2968813};
test_output[2095:2095] = '{32'h4665c423};
test_input[16768:16775] = '{32'h42726a97, 32'h4188f228, 32'h41fde15f, 32'hc1f346b4, 32'h424b58e4, 32'h4296ee44, 32'hc084fd81, 32'h4177ccfd};
test_weights[16768:16775] = '{32'h41a7500a, 32'hc20f5f52, 32'hc211ae47, 32'h42ad7383, 32'h421b61da, 32'h420972ce, 32'h424cc104, 32'h4278855f};
test_bias[2096:2096] = '{32'h425e1194};
test_output[2096:2096] = '{32'h450b9c96};
test_input[16776:16783] = '{32'hc2a00ab9, 32'hc26f6ef8, 32'h4133c239, 32'h4122a357, 32'hbf97f415, 32'h428f271a, 32'h40d820d5, 32'hc2a1744a};
test_weights[16776:16783] = '{32'hc2ab08ef, 32'h41ae69b2, 32'hc2c31bf7, 32'h420b4ebb, 32'hc2c470fd, 32'hc1064ccb, 32'h422fe851, 32'hc20b6f45};
test_bias[2097:2097] = '{32'hc262050c};
test_output[2097:2097] = '{32'h45e63445};
test_input[16784:16791] = '{32'h428ba247, 32'hc2c70a99, 32'h422108db, 32'h41a5fbe3, 32'hc24e701f, 32'h42a7b88c, 32'h4260486e, 32'hc16a6786};
test_weights[16784:16791] = '{32'h41be9d96, 32'h4128b173, 32'hc280d68c, 32'hc1d1aaea, 32'hc281c3d1, 32'h428d5c03, 32'h42331a3e, 32'h423b74e4};
test_bias[2098:2098] = '{32'h4204d8d5};
test_output[2098:2098] = '{32'h4606884c};
test_input[16792:16799] = '{32'hc220eabf, 32'hc2c7b93e, 32'h42b5e33d, 32'hc2396b06, 32'hc051c201, 32'h413bccbd, 32'hc2a28051, 32'hc2c5acfb};
test_weights[16792:16799] = '{32'hc2644c26, 32'hc12877ce, 32'h4239d2af, 32'hc216a402, 32'hc1570278, 32'hc22a9564, 32'hc18553dd, 32'h4136e7c9};
test_bias[2099:2099] = '{32'h42260d8e};
test_output[2099:2099] = '{32'h460e9d6c};
test_input[16800:16807] = '{32'hc2b8af99, 32'h417d4cd9, 32'h4282f69d, 32'hc26ff7b8, 32'h3fc414cf, 32'hc1398cb0, 32'h42b599b8, 32'hc14a55da};
test_weights[16800:16807] = '{32'hc2248482, 32'hc232b61f, 32'hc01a5b5a, 32'h424a75d2, 32'h429bc005, 32'h42b7ccb1, 32'hc075371a, 32'h42583393};
test_bias[2100:2100] = '{32'hc1e12d66};
test_output[2100:2100] = '{32'hc503dbd1};
test_input[16808:16815] = '{32'hc0ee1a56, 32'h424cf1c2, 32'h422b8e15, 32'hc174afb2, 32'hc23eb0cd, 32'h4226b00f, 32'hc287fa94, 32'hc29c73ce};
test_weights[16808:16815] = '{32'h41fcdcda, 32'hc1b89bc7, 32'hc2865f5b, 32'hc21058b4, 32'hc2905386, 32'hc2162264, 32'hc214d451, 32'h425bc8d7};
test_bias[2101:2101] = '{32'hc122fe5a};
test_output[2101:2101] = '{32'hc5641c61};
test_input[16816:16823] = '{32'hc2807044, 32'hc2407452, 32'hc1e518fc, 32'hc29ef493, 32'h40ccf7e3, 32'hc292a412, 32'h4281843b, 32'hc18f86a9};
test_weights[16816:16823] = '{32'h407a2fe8, 32'hc21ad48b, 32'hc2b5a38e, 32'hc2ad6578, 32'hc2805fa0, 32'h42ba8261, 32'hc2a67563, 32'hc20e8e2f};
test_bias[2102:2102] = '{32'hc2957a8c};
test_output[2102:2102] = '{32'hc472c281};
test_input[16824:16831] = '{32'hc1e82231, 32'h41d8cf65, 32'hc22f4b99, 32'hc2a030c4, 32'h426995f1, 32'hc0a708d5, 32'hc28c33ca, 32'hc28e27a0};
test_weights[16824:16831] = '{32'h426686d2, 32'h42c1fe66, 32'h42a0e062, 32'hc2bb5e1f, 32'h3e7f43ae, 32'hc2a55234, 32'h4204d7d0, 32'h424f2396};
test_bias[2103:2103] = '{32'hc28ec460};
test_output[2103:2103] = '{32'hc42ecdb6};
test_input[16832:16839] = '{32'h41945315, 32'hc18abe3d, 32'hc28e8f51, 32'h418738a1, 32'h4281c079, 32'hc230ccc6, 32'hc21365f7, 32'hc2bd2e28};
test_weights[16832:16839] = '{32'hc2c67e64, 32'hc25bc83b, 32'h4200eee9, 32'hc283b3ee, 32'hc289ffbd, 32'hc293f07b, 32'h4294414f, 32'h418ed964};
test_bias[2104:2104] = '{32'h42c47fd4};
test_output[2104:2104] = '{32'hc6198c73};
test_input[16840:16847] = '{32'hc28287e4, 32'h42527ad7, 32'h423cda16, 32'h4210e131, 32'hc28e59b3, 32'h429a928d, 32'h42b2f369, 32'hc1b62922};
test_weights[16840:16847] = '{32'hc0d8e4e9, 32'h40648b88, 32'hc199ea3b, 32'h424c9fe8, 32'hc23810ba, 32'h42a17868, 32'h40b18604, 32'hc2a4da49};
test_bias[2105:2105] = '{32'hc2c3f850};
test_output[2105:2105] = '{32'h4650d3ea};
test_input[16848:16855] = '{32'h42c38f0b, 32'h421708c8, 32'hc23e8bec, 32'h42b7f295, 32'h40a0a0b0, 32'h42bd64ae, 32'h42ab3b48, 32'h428dfded};
test_weights[16848:16855] = '{32'hc144bc1d, 32'hc25a7419, 32'hc22357d9, 32'hc0cb0b29, 32'h4290692a, 32'hc2365f2a, 32'h42a461da, 32'hc2476eb8};
test_bias[2106:2106] = '{32'hc266ade3};
test_output[2106:2106] = '{32'hc51724eb};
test_input[16856:16863] = '{32'h42a1837b, 32'hc2bf2600, 32'h41caae2e, 32'hc0e2ab62, 32'hc1bbae42, 32'hc259683f, 32'hc107a356, 32'h4229dc82};
test_weights[16856:16863] = '{32'hc2905946, 32'h4039720e, 32'h42239f8d, 32'h4262738a, 32'hc2a04767, 32'h41dfec07, 32'hc28f8039, 32'hc27e4c32};
test_bias[2107:2107] = '{32'hc287ac3c};
test_output[2107:2107] = '{32'hc5e33596};
test_input[16864:16871] = '{32'h42ad0155, 32'h41cbceec, 32'h42654432, 32'h42c0f3bb, 32'hc26d9464, 32'hc246429e, 32'hc120d623, 32'h41b717d0};
test_weights[16864:16871] = '{32'h424f3a3e, 32'h42b95c58, 32'h40964a5c, 32'h42719cc0, 32'hc2ad8114, 32'h427eda0d, 32'hc23142ae, 32'h428fa667};
test_bias[2108:2108] = '{32'h41fbe080};
test_output[2108:2108] = '{32'h46853d5d};
test_input[16872:16879] = '{32'hc1f09f94, 32'h422cc754, 32'hc294d0dc, 32'h42c016e8, 32'hc25b9503, 32'h40fd86de, 32'h42c5100b, 32'hc246999f};
test_weights[16872:16879] = '{32'hc0e1f9ff, 32'h428a767b, 32'h4012547f, 32'hc1d72cc3, 32'h421448b7, 32'hc28fcca1, 32'h420de8b4, 32'hc23023a4};
test_bias[2109:2109] = '{32'hc1850fa4};
test_output[2109:2109] = '{32'h455b60bc};
test_input[16880:16887] = '{32'h41aa33a3, 32'hbf994aac, 32'hc1a1b2e9, 32'hc2849db0, 32'hc2b0238d, 32'hc1f783fb, 32'h42950881, 32'hc28a5b98};
test_weights[16880:16887] = '{32'h411cec70, 32'h424371c6, 32'h41a6bdfd, 32'hc10cec45, 32'h4185ee1f, 32'h3e1ab082, 32'hc177a2d9, 32'hbf5e03ff};
test_bias[2110:2110] = '{32'hc0e905b7};
test_output[2110:2110] = '{32'hc50dac89};
test_input[16888:16895] = '{32'h42a03c79, 32'h429a7f30, 32'hc2b21d70, 32'h42a6812a, 32'h42bc40ad, 32'h4218f336, 32'hc20b19b1, 32'h420501a4};
test_weights[16888:16895] = '{32'hc28088d0, 32'hc206a4e2, 32'h414c84b8, 32'hc2ad73f3, 32'hc23b213e, 32'h425227a1, 32'h427f5cc8, 32'h41e82994};
test_bias[2111:2111] = '{32'hc2036498};
test_output[2111:2111] = '{32'hc69a9c72};
test_input[16896:16903] = '{32'h42c3cf8a, 32'h429fe384, 32'h41b06582, 32'h4047d67a, 32'h42bb018d, 32'h418da57e, 32'hc1b4c45b, 32'h42426415};
test_weights[16896:16903] = '{32'h42ba53b8, 32'hc1c77933, 32'h42b0c637, 32'h418bc0e7, 32'hc26de3bb, 32'h40d2a183, 32'hc29224b6, 32'hc1524557};
test_bias[2112:2112] = '{32'h429a6cc0};
test_output[2112:2112] = '{32'h4595454b};
test_input[16904:16911] = '{32'h42bc03a5, 32'hc283b8d1, 32'hc29cf373, 32'h4262d029, 32'hc2b8d43c, 32'h42bdfb4a, 32'h4110ce2f, 32'h41674418};
test_weights[16904:16911] = '{32'h4001a70d, 32'h42178f3f, 32'h42b8752f, 32'hc215e100, 32'h421d35fb, 32'hc2af557d, 32'hc1fc3d50, 32'h429238a1};
test_bias[2113:2113] = '{32'h420818be};
test_output[2113:2113] = '{32'hc6b24b55};
test_input[16912:16919] = '{32'hbf7b8a1d, 32'h4286e78c, 32'hc1ccb7a6, 32'hc17cdb75, 32'hc238d4af, 32'hc2030f01, 32'hc2a53e5b, 32'hc0b7c526};
test_weights[16912:16919] = '{32'hc18943eb, 32'h424bd39e, 32'h428fc634, 32'h42c30a3b, 32'hc201d522, 32'hc19b93f2, 32'hc1ba686f, 32'hc1d20e0f};
test_bias[2114:2114] = '{32'h428f80b6};
test_output[2114:2114] = '{32'h45882fcc};
test_input[16920:16927] = '{32'hc18aa31b, 32'hc2c43fbf, 32'hc23f8f7c, 32'hc2780b43, 32'h4288e919, 32'hc271db04, 32'hc2b17d02, 32'h4259f837};
test_weights[16920:16927] = '{32'h425590b1, 32'h42715bad, 32'hc1c3087b, 32'h4190b6d9, 32'hc262f99d, 32'hc2ba85e1, 32'h42a7acf1, 32'hc2994d45};
test_bias[2115:2115] = '{32'h41f2664e};
test_output[2115:2115] = '{32'hc681f0d5};
test_input[16928:16935] = '{32'h421bbb55, 32'h429fa7a2, 32'h42be590a, 32'hc1724d39, 32'h42438365, 32'h42b895d3, 32'hc10e1420, 32'h42ad005d};
test_weights[16928:16935] = '{32'h42b05ece, 32'hc2adb341, 32'h412a8c03, 32'h41284955, 32'h42a850b0, 32'hc1c5443a, 32'hc1ec9f5f, 32'h4234055c};
test_bias[2116:2116] = '{32'hc27bd51a};
test_output[2116:2116] = '{32'h454d5dc1};
test_input[16936:16943] = '{32'hc1db8c7b, 32'hc265243a, 32'h421682f6, 32'hc22a3cdb, 32'h429e0f4a, 32'hc283ae6c, 32'h40d82cf8, 32'h412f31f7};
test_weights[16936:16943] = '{32'hc131fbd3, 32'hc288ab94, 32'hc2a9cc8e, 32'h41ddc218, 32'h41721e22, 32'h42056ebc, 32'h42b86216, 32'hc2ad881e};
test_bias[2117:2117] = '{32'hc244f890};
test_output[2117:2117] = '{32'hc4bf6b89};
test_input[16944:16951] = '{32'h429bc21b, 32'hc112e720, 32'h4249430d, 32'h427b9578, 32'h425ee5e0, 32'hc29f682b, 32'hc0db36cd, 32'h417a556b};
test_weights[16944:16951] = '{32'h422a5177, 32'hc1e9dd7e, 32'h42893a00, 32'h40f20bbc, 32'h427a6ad7, 32'h427d1e10, 32'h42bde1a7, 32'h41434e32};
test_bias[2118:2118] = '{32'hc1e2644f};
test_output[2118:2118] = '{32'h45aaee90};
test_input[16952:16959] = '{32'h409837b3, 32'hc2a193f4, 32'h4274ba7b, 32'h4269aa76, 32'hc2a6edbc, 32'hc08c10dc, 32'hc21191b0, 32'hc2098542};
test_weights[16952:16959] = '{32'hc2792382, 32'h42a6cdda, 32'h42b01f31, 32'h4296d046, 32'h424da704, 32'h3f8e2e79, 32'h42547f89, 32'h4249a908};
test_bias[2119:2119] = '{32'h4204a262};
test_output[2119:2119] = '{32'hc5a197a3};
test_input[16960:16967] = '{32'hc188535b, 32'hc1dbfc6c, 32'hc2b70777, 32'hc2724493, 32'hc05b992e, 32'h41f76784, 32'h42c2bc4d, 32'hc20ed163};
test_weights[16960:16967] = '{32'hc26d83e1, 32'h4151ccb6, 32'hc24a9658, 32'h428152b3, 32'h42c2223d, 32'hc294f836, 32'hc29a915f, 32'h4294bbfb};
test_bias[2120:2120] = '{32'h4289e81d};
test_output[2120:2120] = '{32'hc631c7be};
test_input[16968:16975] = '{32'h429d5b18, 32'hc113739f, 32'h41d4fd9c, 32'h423f2c9e, 32'h4227707b, 32'hc2b012fe, 32'h424b6fb6, 32'h41e18929};
test_weights[16968:16975] = '{32'h4205a757, 32'hc2abd1c2, 32'hc101b6a5, 32'hc2203970, 32'hc18a0592, 32'h417bd1a7, 32'hc1c36fb4, 32'hc2a2479b};
test_bias[2121:2121] = '{32'h4258c8eb};
test_output[2121:2121] = '{32'hc5862989};
test_input[16976:16983] = '{32'hc051aae4, 32'hc2b051f8, 32'h42b812c7, 32'hc26abb55, 32'hc292d4e8, 32'hc2b6c2f7, 32'hc2357f6b, 32'hc2b027de};
test_weights[16976:16983] = '{32'h407cdd73, 32'hbff445ef, 32'h42977790, 32'hc0d5361b, 32'hc2ae8b47, 32'h42846c05, 32'hc29e193c, 32'h42bca7b8};
test_bias[2122:2122] = '{32'h41b27c15};
test_output[2122:2122] = '{32'h454663ff};
test_input[16984:16991] = '{32'hc217f841, 32'hc1e33f49, 32'h428b4915, 32'h4201d5f0, 32'hc2bd1a1a, 32'hc079f1f8, 32'hc0ff891d, 32'h40c94783};
test_weights[16984:16991] = '{32'hc228dc16, 32'h42a3e4da, 32'h427683e6, 32'h41265d29, 32'h420289f6, 32'hc25206fa, 32'hc0afa313, 32'hc25130c2};
test_bias[2123:2123] = '{32'h42a714c6};
test_output[2123:2123] = '{32'h444dd9c4};
test_input[16992:16999] = '{32'hc16b86de, 32'hc2315e38, 32'hc09f790a, 32'h41dff432, 32'hc29abf4a, 32'hc22ed18c, 32'hc2133dff, 32'hc22e0962};
test_weights[16992:16999] = '{32'hc1d2d3a9, 32'h424f6585, 32'h4270728b, 32'h41d7dd8d, 32'hc23cf62a, 32'hc1d03a30, 32'hc1ec4a0e, 32'hc1965dd4};
test_bias[2124:2124] = '{32'h420c8b91};
test_output[2124:2124] = '{32'h45a4ec43};
test_input[17000:17007] = '{32'h4074c94d, 32'hc211124f, 32'h422a0ea8, 32'h40bf60de, 32'hc1cbd7c3, 32'hbff5495b, 32'hc15874fa, 32'hc2474288};
test_weights[17000:17007] = '{32'hc29b5727, 32'hbfd43bda, 32'h4222e628, 32'hc22fa734, 32'hc2aeb374, 32'hc2c61bf9, 32'h40a1da38, 32'h41d33ea2};
test_bias[2125:2125] = '{32'hc2156141};
test_output[2125:2125] = '{32'h450b2328};
test_input[17008:17015] = '{32'hc270571e, 32'h42b43331, 32'h41d5ae34, 32'hc2779171, 32'h4233c7c4, 32'hc2aeeb92, 32'h418e25a4, 32'hc27ffd0d};
test_weights[17008:17015] = '{32'h418af747, 32'hc220e572, 32'h40fffdd5, 32'hc2b07c70, 32'h424c6e8d, 32'hc2acbddd, 32'h42a4ca5a, 32'h41394ade};
test_bias[2126:2126] = '{32'h42833687};
test_output[2126:2126] = '{32'h4635fb6c};
test_input[17016:17023] = '{32'hc11b704e, 32'hc2763b5a, 32'hc2c300be, 32'hc231bdf8, 32'h4252d338, 32'h42287f43, 32'h42039e3e, 32'h40f8a9a1};
test_weights[17016:17023] = '{32'h3eb5a118, 32'h41afe6ae, 32'hc2c31a0c, 32'h41d108f9, 32'h42b60ba3, 32'hc2992770, 32'hc2a7c02d, 32'hc14f4c14};
test_bias[2127:2127] = '{32'h410536c2};
test_output[2127:2127] = '{32'h45b2866e};
test_input[17024:17031] = '{32'hc2660c0b, 32'h41fb732a, 32'hc2b3c0ca, 32'hc2925e1a, 32'h413e44c9, 32'h4288c2d0, 32'hbd9ac42f, 32'hc2a8f5eb};
test_weights[17024:17031] = '{32'hc26615a0, 32'hc08cc02e, 32'hc247a85b, 32'h426cb987, 32'h423a5823, 32'hc158dcc0, 32'h4241fdf6, 32'hc1be77ac};
test_bias[2128:2128] = '{32'hc22b2dc8};
test_output[2128:2128] = '{32'h4599a7d1};
test_input[17032:17039] = '{32'h429ec076, 32'hbf5fa82d, 32'h41fe9092, 32'hc25f0f23, 32'h421844e3, 32'hc2a3441e, 32'h4185a621, 32'hc2794b2a};
test_weights[17032:17039] = '{32'h42665954, 32'h4144757b, 32'hc23cba3f, 32'h427eae53, 32'h41fb615b, 32'h42befe18, 32'h42afaa62, 32'h41287551};
test_bias[2129:2129] = '{32'h428622ab};
test_output[2129:2129] = '{32'hc5c226ce};
test_input[17040:17047] = '{32'hc2832669, 32'h42521401, 32'hc29ef0bd, 32'h42b7ff63, 32'h414277d0, 32'hc28249dd, 32'h42621996, 32'h41bf9f2b};
test_weights[17040:17047] = '{32'h425c6282, 32'hc26e636e, 32'hc294bd79, 32'hc2c20ba9, 32'hc2a843fd, 32'h42905b23, 32'h41837f81, 32'hc1cff4f5};
test_bias[2130:2130] = '{32'hc2226edb};
test_output[2130:2130] = '{32'hc66dc5a3};
test_input[17048:17055] = '{32'hc2a31412, 32'h41272557, 32'h427b6c25, 32'h4292f15e, 32'h4115735f, 32'hc2a7c79b, 32'h420b7efa, 32'h41e1cdc7};
test_weights[17048:17055] = '{32'h40d64b99, 32'h4249ccc9, 32'hc1872781, 32'h425468d3, 32'hc231b5d8, 32'h4225f913, 32'h42329eb8, 32'h420e7f35};
test_bias[2131:2131] = '{32'hc09a5f4d};
test_output[2131:2131] = '{32'h44b95766};
test_input[17056:17063] = '{32'h428f7a4b, 32'h42c44846, 32'hc0d7c2e6, 32'hc25d12ce, 32'hc19912a4, 32'hc2a55bfd, 32'h42867a17, 32'h41dc0427};
test_weights[17056:17063] = '{32'h3f4df693, 32'h40dd2a4a, 32'h428163a7, 32'hc23df587, 32'hc24f1286, 32'h41d2418f, 32'hc1caba54, 32'h420938ba};
test_bias[2132:2132] = '{32'h41840871};
test_output[2132:2132] = '{32'h44798796};
test_input[17064:17071] = '{32'h428b4cbd, 32'h424349b3, 32'h4282dd14, 32'h42b2a377, 32'hc24c587e, 32'hc101d1e6, 32'h421a8ae4, 32'hc2c762a8};
test_weights[17064:17071] = '{32'hc2a3a227, 32'h4211c984, 32'hc2b961d0, 32'h427e1d56, 32'h4294cfdd, 32'hc214bd2f, 32'hc2023380, 32'hc2a604db};
test_bias[2133:2133] = '{32'hc28f61db};
test_output[2133:2133] = '{32'hc457c09f};
test_input[17072:17079] = '{32'hc285734f, 32'h42abcfff, 32'hc2b2f6eb, 32'h403d9cee, 32'hc13968fb, 32'hc1be419a, 32'hc24b5d77, 32'h42b6172d};
test_weights[17072:17079] = '{32'hc2a84954, 32'h41183392, 32'h41c7c88f, 32'hc19cf0e2, 32'hc1c06747, 32'h4258ece5, 32'hc29a4653, 32'h4242f65d};
test_bias[2134:2134] = '{32'hc2a6ee92};
test_output[2134:2134] = '{32'h46322f18};
test_input[17080:17087] = '{32'hc08a49ed, 32'hc25d7c4a, 32'h42945f84, 32'h4276420d, 32'h427dfcb4, 32'hc2b685cf, 32'hc14cbbab, 32'h41a80b0f};
test_weights[17080:17087] = '{32'h40e42d09, 32'hc20618af, 32'hc1389c77, 32'hc2badd8c, 32'hc281937f, 32'h42c7ba89, 32'h42260fc0, 32'hc261b338};
test_bias[2135:2135] = '{32'hc1f8d4ad};
test_output[2135:2135] = '{32'hc69a5b9a};
test_input[17088:17095] = '{32'hc29dead5, 32'h422b4201, 32'h429df5c9, 32'hc2899578, 32'h41e3fbe7, 32'h42a8c71d, 32'h3fc4d7e7, 32'hc243643e};
test_weights[17088:17095] = '{32'h42522ed6, 32'h40075a24, 32'h42a29cd6, 32'h41708ca1, 32'hc1851e5e, 32'hc2238368, 32'hc25dbdec, 32'h41ca1b79};
test_bias[2136:2136] = '{32'h42371189};
test_output[2136:2136] = '{32'hc571c7c0};
test_input[17096:17103] = '{32'hc23a41ce, 32'hc2a492cd, 32'hc29410b4, 32'h4297c623, 32'h42b18c65, 32'hc2984388, 32'hc180e864, 32'h428bd61e};
test_weights[17096:17103] = '{32'hc0bd5d92, 32'hc0dbb82e, 32'h4288564d, 32'h40ffbfa0, 32'h42391e32, 32'h41e912a5, 32'hc29f6c93, 32'hc2a9f5d6};
test_bias[2137:2137] = '{32'hc0eb84cd};
test_output[2137:2137] = '{32'hc5c72eb0};
test_input[17104:17111] = '{32'hc2491986, 32'h4144a7d8, 32'hc233f206, 32'h3fd37d5e, 32'hc2ac9c53, 32'h4049d694, 32'h42302e57, 32'hc019be52};
test_weights[17104:17111] = '{32'h423e3a26, 32'h428059f0, 32'hc2c760b3, 32'h4245e398, 32'hc1104d55, 32'h42a54b47, 32'hc25d8028, 32'h411cd8ce};
test_bias[2138:2138] = '{32'hc1a3653d};
test_output[2138:2138] = '{32'h44be0918};
test_input[17112:17119] = '{32'h42bf5408, 32'hc19e8262, 32'hc27d1461, 32'hc28be742, 32'hc2961280, 32'hc1a20aea, 32'hc18208c2, 32'h42567be4};
test_weights[17112:17119] = '{32'h427955f8, 32'h418829a8, 32'hc2a6e5f2, 32'h427a1093, 32'hc23af65b, 32'hbf2fee8c, 32'hc2609b5d, 32'h422636d9};
test_bias[2139:2139] = '{32'h42c4ee0c};
test_output[2139:2139] = '{32'h464fb43c};
test_input[17120:17127] = '{32'hc1f24eb9, 32'hc1f066cb, 32'hc27ef28a, 32'h4198a89f, 32'h42c7e5e8, 32'hc26ce0c7, 32'h41d6a9d7, 32'hc257ecf7};
test_weights[17120:17127] = '{32'h420c99d0, 32'hc29855c7, 32'h427c67f5, 32'hc28a1102, 32'hc28eaa8e, 32'h42657554, 32'h4248a5e7, 32'h41ba1f93};
test_bias[2140:2140] = '{32'hc22f554f};
test_output[2140:2140] = '{32'hc6640e16};
test_input[17128:17135] = '{32'h42b49b3a, 32'h42209cd7, 32'h40f25321, 32'h4226a36b, 32'hc13836b1, 32'h422422e1, 32'h40ab0930, 32'h411cf059};
test_weights[17128:17135] = '{32'h4232e249, 32'hc2c0cdd1, 32'h42664110, 32'hc11cf60f, 32'hc1d8cf19, 32'hc25a1936, 32'hc1759d9a, 32'hc24a36b1};
test_bias[2141:2141] = '{32'h42bec893};
test_output[2141:2141] = '{32'hc50a508c};
test_input[17136:17143] = '{32'h412ccd53, 32'h422d9ac0, 32'hc28053b6, 32'hc0fd1448, 32'h4287dbf1, 32'hc0746559, 32'h40c1675c, 32'h41e8646f};
test_weights[17136:17143] = '{32'h42aa738c, 32'h425f0cb6, 32'h40cb8e51, 32'hc20fde96, 32'hc280ac33, 32'h42429510, 32'hc2108d92, 32'hc209b86b};
test_bias[2142:2142] = '{32'h41f3c527};
test_output[2142:2142] = '{32'hc51df4d6};
test_input[17144:17151] = '{32'hc27bbd73, 32'h41980faa, 32'h42a9c322, 32'h42207b2b, 32'h427285bf, 32'h411f3589, 32'hc2c0f3e5, 32'hc2aed76c};
test_weights[17144:17151] = '{32'h414758a5, 32'hc225ca15, 32'h4270e4c5, 32'h4214308b, 32'h42a1f758, 32'hc22be171, 32'hc2661bf2, 32'hc0ffed1c};
test_bias[2143:2143] = '{32'hc267a4d9};
test_output[2143:2143] = '{32'h46755004};
test_input[17152:17159] = '{32'h4204e28d, 32'hc1d9f637, 32'hc2bd94a3, 32'hc1c019c6, 32'h41fd2d5e, 32'h42b53eaf, 32'hc25ba7d6, 32'hc1af0e2a};
test_weights[17152:17159] = '{32'hc2ab139d, 32'hc27617c0, 32'h424c3ddb, 32'hc1d25616, 32'h42ac5d61, 32'hc294977d, 32'h42519ee9, 32'hc09748ff};
test_bias[2144:2144] = '{32'hc1da9300};
test_output[2144:2144] = '{32'hc63e5508};
test_input[17160:17167] = '{32'h420580d6, 32'h4120b92d, 32'hc29cf73b, 32'hc2b05f2d, 32'hc26a341e, 32'hc2088aa2, 32'h42350ec4, 32'h4283787b};
test_weights[17160:17167] = '{32'hc234e564, 32'h4286803e, 32'hc1d128eb, 32'h429cacce, 32'h4214b8a7, 32'h4259aac9, 32'h42813ee8, 32'hc2598ada};
test_bias[2145:2145] = '{32'hc2825dc4};
test_output[2145:2145] = '{32'hc6231f18};
test_input[17168:17175] = '{32'h41df0b01, 32'h42376b3f, 32'h429cf2a4, 32'h42b8d93c, 32'hc00836bb, 32'hc1bcd51b, 32'h41b417e6, 32'h42515529};
test_weights[17168:17175] = '{32'h4113013a, 32'hc122e468, 32'h42c544f3, 32'hc2902fef, 32'hc2986b21, 32'hc19a0b99, 32'h41d50e09, 32'hc232485e};
test_bias[2146:2146] = '{32'h42a5931f};
test_output[2146:2146] = '{32'hc32720e2};
test_input[17176:17183] = '{32'hc2bbf381, 32'h419d1fc9, 32'h42c15a39, 32'h4281b106, 32'h429f5868, 32'hc2ad038e, 32'hc247f016, 32'hc2936ce0};
test_weights[17176:17183] = '{32'hc2c29938, 32'hc2849818, 32'h4266a6fe, 32'h429c06f2, 32'h41d9fa17, 32'hc296a49f, 32'h41d3b6f8, 32'h41a79594};
test_bias[2147:2147] = '{32'h410e5333};
test_output[2147:2147] = '{32'h46bddf91};
test_input[17184:17191] = '{32'hc28aab2a, 32'hc1b83253, 32'h424cf70d, 32'hc2456d42, 32'h429b6832, 32'hc1ebfcb8, 32'h426b794e, 32'h410733db};
test_weights[17184:17191] = '{32'h4299c5f6, 32'hc230c9b0, 32'h4185a8a2, 32'h4299329c, 32'h42bcb1c5, 32'hc2807b1d, 32'h42247077, 32'hc2a9a51b};
test_bias[2148:2148] = '{32'hc28f64d5};
test_output[2148:2148] = '{32'h45623e28};
test_input[17192:17199] = '{32'h426bcbbf, 32'h42a6ab0e, 32'hc13c2af3, 32'h42840460, 32'hc2a39288, 32'h42731c36, 32'h41da3760, 32'h4281ef0c};
test_weights[17192:17199] = '{32'hc213a47b, 32'hc25764ac, 32'h423ce3c7, 32'hc2105e9d, 32'hc2181a53, 32'hc2a89297, 32'h42af3423, 32'h425ee194};
test_bias[2149:2149] = '{32'hc22970b2};
test_output[2149:2149] = '{32'hc5b074ea};
test_input[17200:17207] = '{32'h414fa19d, 32'h4286313e, 32'hc24d6c0a, 32'hc26cb573, 32'h41b90d22, 32'h42772da6, 32'h415be3e8, 32'h429d4dc1};
test_weights[17200:17207] = '{32'hc0f476c4, 32'hc1d8b30d, 32'h4295a4a8, 32'h41fac7ef, 32'hc1e9a58b, 32'hc2ba89d7, 32'h420379ea, 32'hc2a992ae};
test_bias[2150:2150] = '{32'h42a52b4c};
test_output[2150:2150] = '{32'hc69db727};
test_input[17208:17215] = '{32'hc222906d, 32'hc262ac83, 32'h4138ce9a, 32'hc2a5be2d, 32'hc2bf0aa2, 32'h41633829, 32'hc2c54f17, 32'h41fd33e3};
test_weights[17208:17215] = '{32'h42868c41, 32'h42974989, 32'hc2c62edf, 32'hc06025fb, 32'hc10b9d72, 32'hc25ca34a, 32'hc18d1afd, 32'hc2b4ea8e};
test_bias[2151:2151] = '{32'hc2b04911};
test_output[2151:2151] = '{32'hc60d2fa3};
test_input[17216:17223] = '{32'h3df0ea36, 32'h4222d2f5, 32'hc2852fd5, 32'hc2530d3b, 32'hc02b3c25, 32'h416071f9, 32'h3f901de0, 32'h416f9492};
test_weights[17216:17223] = '{32'h424786ae, 32'hc1b33cfc, 32'hc0b1770c, 32'h409a779a, 32'hc2c044bb, 32'hc21e88e9, 32'h4257d101, 32'h42848d33};
test_bias[2152:2152] = '{32'hc2a66b3f};
test_output[2152:2152] = '{32'hc2f0b1c0};
test_input[17224:17231] = '{32'hc23a6e22, 32'h41136037, 32'hc27be9fb, 32'hc28b14fd, 32'h4287e2b5, 32'hc2188bf3, 32'h41905c94, 32'h42b799d9};
test_weights[17224:17231] = '{32'h422d619a, 32'h42808a19, 32'hc1a3ad1c, 32'h3e1ed26d, 32'h41ff6624, 32'hc23f5e04, 32'hc1157789, 32'h42a987f3};
test_bias[2153:2153] = '{32'h42a2bf0e};
test_output[2153:2153] = '{32'h4634459c};
test_input[17232:17239] = '{32'h42c281bc, 32'h429d96f9, 32'h417bdb95, 32'h41bda5fb, 32'hc28bdc5b, 32'hc255e9bd, 32'h4298d920, 32'hc222cdac};
test_weights[17232:17239] = '{32'h42056525, 32'h427057ed, 32'hc29c1bfd, 32'h42a31ddd, 32'hc2aa41e9, 32'hc27e854b, 32'hc2b9ca49, 32'h423696d3};
test_bias[2154:2154] = '{32'h41afde32};
test_output[2154:2154] = '{32'h460e3c5e};
test_input[17240:17247] = '{32'hbeffef3f, 32'h42893ffe, 32'hc25fc381, 32'hc288c7a2, 32'hc1b98003, 32'h42133605, 32'hc0374c98, 32'hc16609a4};
test_weights[17240:17247] = '{32'hc23b2e2f, 32'hc0a0d3e1, 32'hc1986cab, 32'hc28fbbb0, 32'hc16d1243, 32'hc26cf083, 32'hc2c5a7d8, 32'h4244d655};
test_bias[2155:2155] = '{32'hc295ccd5};
test_output[2155:2155] = '{32'h454fb7ef};
test_input[17248:17255] = '{32'h4284bd25, 32'hc242b9ac, 32'h42308838, 32'hc290db4f, 32'hc1dd949e, 32'hc08f074e, 32'hc08d9bd0, 32'h42bf2807};
test_weights[17248:17255] = '{32'h423e693f, 32'hc2934d92, 32'h422ef0df, 32'h42c4affc, 32'hc10e1243, 32'h4216ba8b, 32'h42a2e4f8, 32'hc1a9d546};
test_bias[2156:2156] = '{32'hc2874f5e};
test_output[2156:2156] = '{32'hc44edf8b};
test_input[17256:17263] = '{32'h4295b86f, 32'h42c4adac, 32'h42bce8b3, 32'h42579ccc, 32'hc2842c4b, 32'h421c9629, 32'h4273f6db, 32'h40311f39};
test_weights[17256:17263] = '{32'hc213fecc, 32'hc1834012, 32'hc01a3fdb, 32'hc224749d, 32'h424e2616, 32'hc16f10d5, 32'h41624f0c, 32'hc2681496};
test_bias[2157:2157] = '{32'h42803a6b};
test_output[2157:2157] = '{32'hc61d0e2f};
test_input[17264:17271] = '{32'hc29edea5, 32'hc1ad0b04, 32'hc2c39073, 32'hc1242ec7, 32'h41cd5884, 32'hc13a37fc, 32'hc2761e33, 32'hc284adab};
test_weights[17264:17271] = '{32'hc27b449d, 32'hc26c96a0, 32'h410df3f5, 32'h42c23ca5, 32'hc24f37b0, 32'hc224062d, 32'h421d832e, 32'hc2ad6c7b};
test_bias[2158:2158] = '{32'hc2a8f945};
test_output[2158:2158] = '{32'h45d46d3f};
test_input[17272:17279] = '{32'hc235900d, 32'h41da2dc1, 32'hc223dad3, 32'h41222879, 32'h41f55022, 32'h40a27b7a, 32'h42c1e5db, 32'h427cedc3};
test_weights[17272:17279] = '{32'hc1e41d8a, 32'h42579aa6, 32'hc2a931ce, 32'h42569e03, 32'hc2a1c3a6, 32'hc21e7ab9, 32'h420fb436, 32'hc1609135};
test_bias[2159:2159] = '{32'hc223bb0d};
test_output[2159:2159] = '{32'h45cfb59e};
test_input[17280:17287] = '{32'hc28cd0d3, 32'hc247ef90, 32'h41c87cce, 32'h41d27d75, 32'hc2a83763, 32'h421ba554, 32'h410c2481, 32'h42bf93a7};
test_weights[17280:17287] = '{32'h42c06aa0, 32'hc21c9b07, 32'hc2afc8dc, 32'hc22397cb, 32'h4145f8ea, 32'hc247b791, 32'hc2b16dfd, 32'h42a7aa12};
test_bias[2160:2160] = '{32'h41c3786a};
test_output[2160:2160] = '{32'hc56d999b};
test_input[17288:17295] = '{32'hc1af4892, 32'hc2936526, 32'hc239c5a6, 32'h4282d2dd, 32'h42911c24, 32'hbf8ed73f, 32'hc1859f4c, 32'hc207cd46};
test_weights[17288:17295] = '{32'h429160f8, 32'hc28b3337, 32'hc28b6e7f, 32'hc286d5fd, 32'h41a54fd9, 32'h42bd1943, 32'h418a8703, 32'h41bf29f2};
test_bias[2161:2161] = '{32'h424915e1};
test_output[2161:2161] = '{32'h452941fc};
test_input[17296:17303] = '{32'hc246eb83, 32'hc0fb53d5, 32'h42add618, 32'hc287cae3, 32'h420f8d87, 32'hc2329749, 32'h3fa84a0d, 32'hc14c81a5};
test_weights[17296:17303] = '{32'hc0aac41d, 32'hc01ee744, 32'h42848e6e, 32'hc2a03e11, 32'h41a529b7, 32'hc10873ce, 32'h42448424, 32'h42c2fd04};
test_bias[2162:2162] = '{32'h42a46153};
test_output[2162:2162] = '{32'h4633cfb9};
test_input[17304:17311] = '{32'h40161ba9, 32'h41accdc8, 32'h41aa9f11, 32'h4148617e, 32'hc135a69e, 32'hc286af85, 32'hc08f7c74, 32'hc1c3f94a};
test_weights[17304:17311] = '{32'h420c38d4, 32'hc28d1e3a, 32'hc1fb2c64, 32'hc295cf8e, 32'hc22b973e, 32'hc23d6e9f, 32'h427dc5c3, 32'h425a7a30};
test_bias[2163:2163] = '{32'h42aaa1b2};
test_output[2163:2163] = '{32'hc463a0ca};
test_input[17312:17319] = '{32'h422bcf7f, 32'hc19cebd8, 32'hc2603d52, 32'h429daf73, 32'hc22a8d80, 32'hc0921802, 32'hc214f80e, 32'hc299e49d};
test_weights[17312:17319] = '{32'hc2941deb, 32'h422a9aef, 32'hc1c6c714, 32'hc2bced55, 32'hc2970b56, 32'h424f4a42, 32'hc18828f8, 32'hc2ad70f3};
test_bias[2164:2164] = '{32'h422f3ff2};
test_output[2164:2164] = '{32'h4382cead};
test_input[17320:17327] = '{32'hc18fcc13, 32'h4294acb4, 32'h4210105f, 32'hc1a7d2a3, 32'hc199d8f3, 32'h423fe877, 32'h424a382c, 32'h4249547d};
test_weights[17320:17327] = '{32'h41fc532f, 32'hc2663050, 32'h42186838, 32'hc2721d4a, 32'h415f8d03, 32'hc1739706, 32'h4233c9d7, 32'h42b22eb1};
test_bias[2165:2165] = '{32'hc2adbad3};
test_output[2165:2165] = '{32'h4558bb2f};
test_input[17328:17335] = '{32'h4200c862, 32'hc235780b, 32'hc2c2f22b, 32'hc06f5ad6, 32'hc2682b0c, 32'h41f9e0f6, 32'hc20315c7, 32'h41a9610c};
test_weights[17328:17335] = '{32'h42843baa, 32'h42978b46, 32'hc229d80c, 32'h41bc09de, 32'h4233626e, 32'h429b572e, 32'h4224f190, 32'hc0da8e13};
test_bias[2166:2166] = '{32'h42616a47};
test_output[2166:2166] = '{32'h448cae5c};
test_input[17336:17343] = '{32'hc09545d8, 32'hc2157f47, 32'h42ad06d1, 32'h42840549, 32'hc0ea6bfd, 32'hc21a811a, 32'hc29f0c61, 32'hc201d5af};
test_weights[17336:17343] = '{32'h4267f304, 32'h42bd62ae, 32'hc272c0d3, 32'hc20d8b68, 32'h3f3e05b0, 32'h4281a182, 32'h42ae4ca7, 32'hc225f14c};
test_bias[2167:2167] = '{32'hc28c9768};
test_output[2167:2167] = '{32'hc698ce04};
test_input[17344:17351] = '{32'h425f2bc3, 32'h42a98f12, 32'h42941dc5, 32'h4293cc1d, 32'hc23895ce, 32'hc057bf54, 32'h42c4cf0d, 32'hc18fe817};
test_weights[17344:17351] = '{32'h4105fc21, 32'hc21d074b, 32'hc25dea41, 32'h41a5975b, 32'hc293ead5, 32'hc2c0f932, 32'hc2c379b5, 32'hc1d92e59};
test_bias[2168:2168] = '{32'hc0ba08a2};
test_output[2168:2168] = '{32'hc6295487};
test_input[17352:17359] = '{32'hc2aa11fd, 32'h42b6d5eb, 32'h42c4fd2d, 32'hc2a0cd48, 32'hc28738b0, 32'h3f8add71, 32'hc2af3f0a, 32'h42b5b2d0};
test_weights[17352:17359] = '{32'h429863e0, 32'hc2bb49e4, 32'hc1706cf1, 32'h42631a24, 32'h4283bef0, 32'h42c3767c, 32'hc1741d82, 32'hc1220cbd};
test_bias[2169:2169] = '{32'hc21a5c3b};
test_output[2169:2169] = '{32'hc6c3bcc5};
test_input[17360:17367] = '{32'h41b81107, 32'h41df83e2, 32'h40c6f2ae, 32'h420dc31f, 32'h4195d927, 32'hc22fcf72, 32'h40e3feae, 32'hc1868f17};
test_weights[17360:17367] = '{32'hc287d8e9, 32'hc29383f7, 32'hc26d0219, 32'h4264e5c0, 32'hc22b1403, 32'h42901bf5, 32'h42203db6, 32'h41754c57};
test_bias[2170:2170] = '{32'h41b45e35};
test_output[2170:2170] = '{32'hc5b7cefb};
test_input[17368:17375] = '{32'hc2833956, 32'hc298f4b5, 32'hc200d773, 32'h40a85dc5, 32'h4237b465, 32'h421cb8a0, 32'hc2323fad, 32'hc2088436};
test_weights[17368:17375] = '{32'hc2a4eb53, 32'h4231299c, 32'hc08ecdec, 32'h42bd61da, 32'h426eedef, 32'hc1481749, 32'hc1880a49, 32'h42413d45};
test_bias[2171:2171] = '{32'h427864e3};
test_output[2171:2171] = '{32'h457f9728};
test_input[17376:17383] = '{32'h42c2e8a9, 32'hc2c476b4, 32'hc1fe3aa5, 32'hc29c8293, 32'h42a9640d, 32'h411ac924, 32'hc1cbd22c, 32'h41ec9ed9};
test_weights[17376:17383] = '{32'h41db5f8c, 32'h4284c511, 32'hc258d20e, 32'hc28af441, 32'h4082634a, 32'h42c61147, 32'h4219441e, 32'hc292387a};
test_bias[2172:2172] = '{32'hc27ccf74};
test_output[2172:2172] = '{32'h44b08231};
test_input[17384:17391] = '{32'h423b1300, 32'hc222a1ae, 32'hc19af746, 32'h423835ac, 32'hc28f1e2c, 32'h414d14b1, 32'hc28d19b7, 32'hc241bcf6};
test_weights[17384:17391] = '{32'hc23c9aee, 32'hc2a7167d, 32'hc29a559b, 32'h42885b07, 32'hc244baca, 32'hc2a89e83, 32'hc233a66f, 32'hc1538fc6};
test_bias[2173:2173] = '{32'h421880a9};
test_output[2173:2173] = '{32'h463d4002};
test_input[17392:17399] = '{32'hc1c193ee, 32'hc2b35893, 32'hc29d3a35, 32'h42bfd825, 32'hc2994d4e, 32'h426ec6b3, 32'hc28fae06, 32'hc1df3e6b};
test_weights[17392:17399] = '{32'hc27408dc, 32'hc18a33c6, 32'h42b53b06, 32'h42862b46, 32'h42185c41, 32'hc2078770, 32'hc2ac7b93, 32'h4296140c};
test_bias[2174:2174] = '{32'h428fe816};
test_output[2174:2174] = '{32'h44c3fedc};
test_input[17400:17407] = '{32'h428c1e2d, 32'hc27300a5, 32'h42a1fbd9, 32'hc2162bee, 32'h424a61ee, 32'h42c7360a, 32'h42760b41, 32'h42677332};
test_weights[17400:17407] = '{32'h4290e277, 32'hc1e52cb9, 32'h41eb2828, 32'hbfbe3b1c, 32'h428f01df, 32'hc227a5e1, 32'hc239c7e6, 32'h4210ba0a};
test_bias[2175:2175] = '{32'h4298d1d6};
test_output[2175:2175] = '{32'h45fa4204};
test_input[17408:17415] = '{32'h42a14b41, 32'h41e713a9, 32'h41b48eea, 32'h426d1f24, 32'hc28a85b5, 32'hc29565dd, 32'hc2943a37, 32'hc1da0899};
test_weights[17408:17415] = '{32'hc2b79f66, 32'hc0d8e6a0, 32'hc2672c9e, 32'h41c5ff63, 32'hc20c40c2, 32'h41ed2187, 32'hc2a3c764, 32'hc13c1a1e};
test_bias[2176:2176] = '{32'hc079421f};
test_output[2176:2176] = '{32'hc4515475};
test_input[17416:17423] = '{32'hc1851fbb, 32'hc0539bbd, 32'hc0cb7188, 32'hc24fc0b5, 32'h42c34691, 32'h4275ddbb, 32'hc25a7eb2, 32'h42b95dd5};
test_weights[17416:17423] = '{32'hc1f65fa9, 32'h426e24dc, 32'hc2ad4a3b, 32'h4223cade, 32'h42a495a6, 32'hc2178313, 32'h42b00de5, 32'hc2976434};
test_bias[2177:2177] = '{32'hc12caa9f};
test_output[2177:2177] = '{32'hc5e6e48f};
test_input[17424:17431] = '{32'h429f1918, 32'hc242dad8, 32'hc11f0b61, 32'hc190b941, 32'h4219d182, 32'h418d07f0, 32'hc1b5e2f3, 32'h4274c6bd};
test_weights[17424:17431] = '{32'h42612eec, 32'h419b8d20, 32'h4257d38d, 32'hc238608b, 32'hc185d7bb, 32'hc2b9e578, 32'h401c3f72, 32'h40a85175};
test_bias[2178:2178] = '{32'hc28f2d46};
test_output[2178:2178] = '{32'h44d9aef4};
test_input[17432:17439] = '{32'h425f2617, 32'h429063e0, 32'h42288599, 32'hbfcfbb9b, 32'h42032381, 32'h4296af60, 32'hbe32d8eb, 32'hc1d141bd};
test_weights[17432:17439] = '{32'h425dc388, 32'h42b718c1, 32'hc1ebfe36, 32'h41fe88fb, 32'h422620e4, 32'h42244d85, 32'hc2c1985f, 32'hc2b20e63};
test_bias[2179:2179] = '{32'hc0a54822};
test_output[2179:2179] = '{32'h466d926f};
test_input[17440:17447] = '{32'h42a1037d, 32'hc2b049d8, 32'hc29e6673, 32'hc29f0cde, 32'h422419a5, 32'h40d632a9, 32'hc24c4c9d, 32'hc12cf58d};
test_weights[17440:17447] = '{32'h41a5ff30, 32'h42b3ee3c, 32'hc1267486, 32'h4269f940, 32'h42b933f4, 32'h428583b4, 32'h42035f1d, 32'h41a813d3};
test_bias[2180:2180] = '{32'hc09d54f5};
test_output[2180:2180] = '{32'hc5f23695};
test_input[17448:17455] = '{32'h42c33c74, 32'h41f3ff1f, 32'h42aacbf1, 32'h428a3b06, 32'hc28f6251, 32'hc2026fef, 32'hc27cfb11, 32'hc2758da1};
test_weights[17448:17455] = '{32'h4199fc99, 32'h4245b2d1, 32'h426418bf, 32'h422a0163, 32'h4149a3ae, 32'h41a593a6, 32'h42926b55, 32'h41afb123};
test_bias[2181:2181] = '{32'h426e4342};
test_output[2181:2181] = '{32'h456707e4};
test_input[17456:17463] = '{32'hc2329ec2, 32'h41d5e009, 32'h422da73d, 32'hc2a8589a, 32'h4270a964, 32'hc22cbc79, 32'hc20555b8, 32'hc2a951be};
test_weights[17456:17463] = '{32'hc189e10e, 32'hc2644f8a, 32'h4208e649, 32'hc223f10c, 32'h420b3200, 32'h4293f2de, 32'hc13470c3, 32'h40c2234c};
test_bias[2182:2182] = '{32'h418fca30};
test_output[2182:2182] = '{32'h4538ed33};
test_input[17464:17471] = '{32'h41944765, 32'h42925b3c, 32'hc28df3a5, 32'hc2ae4ba5, 32'h4143fa5d, 32'hc2a4a63e, 32'hc005f918, 32'h42259c90};
test_weights[17464:17471] = '{32'h42818705, 32'hc2863625, 32'hc05056f5, 32'hc281ac54, 32'hbf961f8e, 32'hc2bb05b8, 32'h41f2ad58, 32'h42b5e8a6};
test_bias[2183:2183] = '{32'h41c49f7e};
test_output[2183:2183] = '{32'h46543788};
test_input[17472:17479] = '{32'hc2958e16, 32'h410773be, 32'hc1f0b0bc, 32'h429b6310, 32'h428ddab0, 32'hc191e2e1, 32'hc271c002, 32'h426b6573};
test_weights[17472:17479] = '{32'hc2a4b5c4, 32'hc242ffc3, 32'h4297f312, 32'h4282c358, 32'h415e0808, 32'hc21c2b20, 32'h42816d1d, 32'h3eb17509};
test_bias[2184:2184] = '{32'h429b300d};
test_output[2184:2184] = '{32'h45c8b503};
test_input[17480:17487] = '{32'hc28fba20, 32'h3f36592e, 32'hc28f6397, 32'h3edd3ea1, 32'hc1ca5a28, 32'hc05fa4eb, 32'h42c61307, 32'h415a70cd};
test_weights[17480:17487] = '{32'hc238b579, 32'hc181ffe8, 32'h41c2335e, 32'h41d9dabf, 32'h42803001, 32'hc275978e, 32'h42bd54a3, 32'h4276871e};
test_bias[2185:2185] = '{32'hc2bdfdb0};
test_output[2185:2185] = '{32'h4620d5c6};
test_input[17488:17495] = '{32'h42bbad83, 32'h426f9bc3, 32'hc2aa8ccc, 32'h41e56c57, 32'h41fca0d8, 32'hc19b3183, 32'hc1efda7a, 32'h41c33890};
test_weights[17488:17495] = '{32'h42c0b0c1, 32'hc27ecb3a, 32'h42567ee6, 32'hc1d895b0, 32'h42b8b698, 32'hc279a092, 32'hc284868d, 32'h42176a94};
test_bias[2186:2186] = '{32'hc10abbe5};
test_output[2186:2186] = '{32'h45d7c78a};
test_input[17496:17503] = '{32'h40936de3, 32'h3f8483f3, 32'h41b99ce0, 32'h42a18820, 32'h42a3a872, 32'h423eab9d, 32'h422ec1d8, 32'h41d626f6};
test_weights[17496:17503] = '{32'h42687a5b, 32'hc2a11079, 32'hc2c15340, 32'h419e9aba, 32'h41491a81, 32'h4057d9f6, 32'h413319f9, 32'hc2b21627};
test_bias[2187:2187] = '{32'hc09ee44f};
test_output[2187:2187] = '{32'hc491eb23};
test_input[17504:17511] = '{32'hc19d0f43, 32'h409bbd8e, 32'h418f0e06, 32'h42acfb6d, 32'hc2bcfdf9, 32'hc2bfa153, 32'hc2684906, 32'h42a102d5};
test_weights[17504:17511] = '{32'hc2b08053, 32'hc089a359, 32'h428ba086, 32'h418f4e72, 32'hc2bbc207, 32'h4170396b, 32'hc0f48309, 32'hc269aa6d};
test_bias[2188:2188] = '{32'h41a7e683};
test_output[2188:2188] = '{32'h45f0bee9};
test_input[17512:17519] = '{32'h4239d58b, 32'h420dea5c, 32'hc2b27a38, 32'h41859485, 32'h428bf0ec, 32'hc2739444, 32'h4295d76e, 32'h42c715c6};
test_weights[17512:17519] = '{32'h42b922ed, 32'h422e2ec1, 32'hc2b471d9, 32'h4212b026, 32'h413488ff, 32'hc187201e, 32'hc23f7a16, 32'h423a55de};
test_bias[2189:2189] = '{32'hc2bc32f6};
test_output[2189:2189] = '{32'h468707aa};
test_input[17520:17527] = '{32'h42285b22, 32'hc2b64950, 32'h424a6046, 32'hc29cacda, 32'hc25e6642, 32'h41c73b40, 32'h42962987, 32'h40c0530b};
test_weights[17520:17527] = '{32'hc241bc9d, 32'h417a7895, 32'h416e7ca6, 32'hc2c44933, 32'h428650ad, 32'h3f6d422e, 32'h428319c7, 32'hc24b1aca};
test_bias[2190:2190] = '{32'hc016cba3};
test_output[2190:2190] = '{32'h45b7c217};
test_input[17528:17535] = '{32'hc296835a, 32'hc2588446, 32'hc1866412, 32'h4289ac3f, 32'h42a8b992, 32'hc28f3ca2, 32'hc2c0c98a, 32'h428d46aa};
test_weights[17528:17535] = '{32'h4230d942, 32'h4190fd50, 32'hc1e024d5, 32'h4197319e, 32'h3fe72bf5, 32'hc206193a, 32'hc1877254, 32'h4230d50f};
test_bias[2191:2191] = '{32'hc2b99d36};
test_output[2191:2191] = '{32'h4592356f};
test_input[17536:17543] = '{32'hc27bf9d4, 32'h41964867, 32'hc273dd29, 32'h421ca888, 32'h40b318d1, 32'h4259b6ea, 32'h42b47727, 32'hc27779fd};
test_weights[17536:17543] = '{32'hc1dad4aa, 32'hc2bd712f, 32'hc1e4ae47, 32'h42928644, 32'h415bd1a4, 32'h4299c171, 32'hc0574105, 32'h41c2278b};
test_bias[2192:2192] = '{32'h4222baab};
test_output[2192:2192] = '{32'h45dc657c};
test_input[17544:17551] = '{32'hc224716b, 32'h4234e534, 32'h3b6176a0, 32'hc212617c, 32'h42a2a3ca, 32'h428d01fc, 32'hc224429a, 32'h42a58d9a};
test_weights[17544:17551] = '{32'h42233824, 32'hc15d2d0b, 32'hc1f75e28, 32'hc29fc627, 32'h428e025e, 32'hc1513de0, 32'h4088c5e2, 32'h42b08b4b};
test_bias[2193:2193] = '{32'h41eae113};
test_output[2193:2193] = '{32'h464565e4};
test_input[17552:17559] = '{32'h421b961e, 32'h4212cbf9, 32'hc22bc7e1, 32'h4289a41e, 32'hc21e4f10, 32'h423a4d5d, 32'hc18d780d, 32'h42b5a0b5};
test_weights[17552:17559] = '{32'h427ab2b9, 32'hc26b33c8, 32'h40fb2441, 32'hc22054a7, 32'h42815670, 32'h429e41d0, 32'hbfa7a3d5, 32'hc23ef88c};
test_bias[2194:2194] = '{32'hc2777057};
test_output[2194:2194] = '{32'hc5bd8024};
test_input[17560:17567] = '{32'hc1a10603, 32'hc20eb578, 32'hc0a4e559, 32'hc2bd493c, 32'h41f93b6a, 32'hc25f3e34, 32'h4269dbea, 32'hc294e213};
test_weights[17560:17567] = '{32'hc2222792, 32'hc10f4a97, 32'h420c43d6, 32'hc2051cda, 32'hc294272c, 32'h4294face, 32'h42c177b8, 32'h41e68a64};
test_bias[2195:2195] = '{32'hc27f5476};
test_output[2195:2195] = '{32'h4487b58c};
test_input[17568:17575] = '{32'hc234b3b6, 32'h429228db, 32'h42c3fbb8, 32'h421f9d55, 32'hc24f8315, 32'hc2bf666c, 32'h42ba4d93, 32'h41ce1e63};
test_weights[17568:17575] = '{32'hc2485612, 32'hc162f987, 32'h422db911, 32'h409d0305, 32'hc29d14bf, 32'hc12b88d9, 32'hc2c0cf33, 32'hc23205df};
test_bias[2196:2196] = '{32'h427d6da8};
test_output[2196:2196] = '{32'h44329d3f};
test_input[17576:17583] = '{32'h422072a9, 32'hc222c86a, 32'h425233c7, 32'hc238d1f7, 32'h427d891d, 32'h3f68c568, 32'hc2aeeaaa, 32'hc23b16c9};
test_weights[17576:17583] = '{32'hc2a9b0b1, 32'h423394c2, 32'hc2be1982, 32'hc2c0dfd7, 32'h410d0e47, 32'hc255d0e4, 32'hc226c913, 32'hc1df48a0};
test_bias[2197:2197] = '{32'hc2739b06};
test_output[2197:2197] = '{32'hc3b7fc4a};
test_input[17584:17591] = '{32'hc1fe609f, 32'h4173f830, 32'hbf55cb8f, 32'h41c58048, 32'hc2bf5532, 32'hc2a9506a, 32'hc273b681, 32'hc292ebd5};
test_weights[17584:17591] = '{32'hc2271e5a, 32'h418b46d6, 32'h426f6361, 32'h429a6d9c, 32'hc2bb6544, 32'hc268cfd6, 32'h42156087, 32'h42027b8a};
test_bias[2198:2198] = '{32'h42c4082d};
test_output[2198:2198] = '{32'h46477e4c};
test_input[17592:17599] = '{32'h41b26458, 32'h3e902764, 32'h41d03ca8, 32'hc2b89b3c, 32'hc23a76c4, 32'h429d73bf, 32'hc22b7c97, 32'h42b767e8};
test_weights[17592:17599] = '{32'hc23c8b40, 32'h42973c31, 32'hc20c98ee, 32'hc1edde2e, 32'hc08a5439, 32'h4246be96, 32'h4291a4c5, 32'hc1296a02};
test_bias[2199:2199] = '{32'hc13a795e};
test_output[2199:2199] = '{32'h444a0fce};
test_input[17600:17607] = '{32'h4214f6db, 32'hc162e465, 32'h41cf5dfb, 32'hc264769f, 32'h418f7784, 32'hc252c16d, 32'h41306057, 32'hc2a3c26a};
test_weights[17600:17607] = '{32'h429ea2d6, 32'h428b9cd8, 32'h42ab7d66, 32'hc1e762f5, 32'h4210ed3e, 32'h4218519d, 32'h42b12c4a, 32'hc2c7a57d};
test_bias[2200:2200] = '{32'hc244f83f};
test_output[2200:2200] = '{32'h46543adb};
test_input[17608:17615] = '{32'h41dcc91a, 32'hc2c5b230, 32'h41c0065d, 32'h423036fd, 32'h4296fd73, 32'h4249cd47, 32'h40852df4, 32'hc2710b52};
test_weights[17608:17615] = '{32'hc1fe4225, 32'h41478897, 32'h41558be4, 32'h415058d8, 32'hc18db5ad, 32'hc0b3df71, 32'hc2815956, 32'hc24be171};
test_bias[2201:2201] = '{32'h42aab7d0};
test_output[2201:2201] = '{32'h424bf601};
test_input[17616:17623] = '{32'hc2020379, 32'h4240ffb1, 32'hc249f9cf, 32'hc10f3f23, 32'hc12badd1, 32'hc12733af, 32'h42902275, 32'hc2bbd4aa};
test_weights[17616:17623] = '{32'hc1c7e38e, 32'hc16fbee1, 32'h4226b1dc, 32'h420ca639, 32'h426a071b, 32'hc1e4b927, 32'hc256a1eb, 32'hc29561ff};
test_bias[2202:2202] = '{32'hc17d3767};
test_output[2202:2202] = '{32'h43ec7675};
test_input[17624:17631] = '{32'hc28e26a8, 32'hc22e5498, 32'h416ef683, 32'h421d3533, 32'hc183cca5, 32'h40ed03da, 32'hc291e52e, 32'h41801c62};
test_weights[17624:17631] = '{32'hc250f7c2, 32'hc2b4f7e3, 32'hc2a68f73, 32'h420a7bc4, 32'h3f3c8e86, 32'h421bff77, 32'hc241bd48, 32'h423e0292};
test_bias[2203:2203] = '{32'hc1653eba};
test_output[2203:2203] = '{32'h4640a74a};
test_input[17632:17639] = '{32'h428154bd, 32'h413c3582, 32'h42ab9ea6, 32'hc28ce9c1, 32'h4292ca54, 32'hc272761a, 32'h41a74de1, 32'hc214578d};
test_weights[17632:17639] = '{32'hc22e7c88, 32'h42ad948c, 32'h428b5907, 32'hc23fd9bd, 32'h3fd8c2cf, 32'hc0c0b306, 32'hc129ddfb, 32'hc294aba8};
test_bias[2204:2204] = '{32'hc2c495b2};
test_output[2204:2204] = '{32'h4623cf5c};
test_input[17640:17647] = '{32'h424485db, 32'hc2a64342, 32'h42988513, 32'hc109596c, 32'hc25d5bad, 32'hc2556c7a, 32'h42a8c83d, 32'hc2975ae8};
test_weights[17640:17647] = '{32'hc27260a8, 32'h429d0c8d, 32'h418547ed, 32'h42586b81, 32'hc2c1aab3, 32'h3f562f6d, 32'hc21a0c26, 32'hc2c16b18};
test_bias[2205:2205] = '{32'hc0864164};
test_output[2205:2205] = '{32'h4429eba0};
test_input[17648:17655] = '{32'h412f445d, 32'hc2bffcb5, 32'hc23d268a, 32'h428ac6c9, 32'h42b5f54d, 32'h428f3135, 32'hc156ed35, 32'hc13af690};
test_weights[17648:17655] = '{32'h40194775, 32'h4201de3b, 32'hc2434459, 32'hc2a43193, 32'h42ba5db9, 32'hc2082d5b, 32'hc2b2542f, 32'h41894cf2};
test_bias[2206:2206] = '{32'hc21b5833};
test_output[2206:2206] = '{32'h440206ef};
test_input[17656:17663] = '{32'h42beedd9, 32'h42805d65, 32'h42a10323, 32'h3f8e6d79, 32'h427c0d7c, 32'hc2ba0952, 32'hc1a26fc2, 32'h41d16626};
test_weights[17656:17663] = '{32'h403c8e0a, 32'hc23e7c00, 32'hc1c800b7, 32'h41efab79, 32'h42ae9163, 32'hc29c0364, 32'hc1d4541f, 32'h41872b6b};
test_bias[2207:2207] = '{32'h423cf008};
test_output[2207:2207] = '{32'h460d17c5};
test_input[17664:17671] = '{32'h429e0a29, 32'hc120bea4, 32'hc2916df0, 32'hc237fc88, 32'h41a6b79d, 32'h40dff7de, 32'h41cb13de, 32'h41e5dea4};
test_weights[17664:17671] = '{32'h42808889, 32'h429f680a, 32'h42482fd7, 32'h4232cee3, 32'hc20c1eb7, 32'h4244879f, 32'h41b9d6e2, 32'hc2436e37};
test_bias[2208:2208] = '{32'hc1c97d82};
test_output[2208:2208] = '{32'hc52532c3};
test_input[17672:17679] = '{32'hc287be2c, 32'h4130ac51, 32'hc2c5dfbe, 32'h42882ff2, 32'h410e9998, 32'h42703158, 32'hc16dfd78, 32'hc1043e8d};
test_weights[17672:17679] = '{32'h42b4261f, 32'hc141298e, 32'hc1b61366, 32'h42a89117, 32'hc2bc7ef4, 32'hc2c7f18a, 32'h4215153a, 32'h4212f560};
test_bias[2209:2209] = '{32'h41bfb5fe};
test_output[2209:2209] = '{32'hc5b9687a};
test_input[17680:17687] = '{32'hc0e535dd, 32'h3f988c98, 32'hc08d96a6, 32'h42ad3e3f, 32'hc2904b99, 32'hc2c52399, 32'hc2819971, 32'hc28a813f};
test_weights[17680:17687] = '{32'h419db61c, 32'h425f2740, 32'h42a938b1, 32'hc195bf62, 32'h41919c5d, 32'h41113383, 32'h42b85680, 32'hc25cb5e0};
test_bias[2210:2210] = '{32'h4265cb89};
test_output[2210:2210] = '{32'hc5c720e1};
test_input[17688:17695] = '{32'h40a7d5dd, 32'h4240400c, 32'hc2af8e7e, 32'h41ae1339, 32'hc15f7abe, 32'hc268ccaa, 32'h4290edba, 32'hc2c5a6b4};
test_weights[17688:17695] = '{32'hc29cf411, 32'h42b87cf4, 32'h41267ef0, 32'hc13cde15, 32'hc2b412c2, 32'hc2076f1e, 32'hc2375577, 32'h426cebb8};
test_bias[2211:2211] = '{32'hc24e81c8};
test_output[2211:2211] = '{32'hc544a9e9};
test_input[17696:17703] = '{32'h42b977f4, 32'hc18676bf, 32'h4282e264, 32'hc2694119, 32'hc1cf5dd9, 32'h409e800c, 32'h41a06b06, 32'h42951881};
test_weights[17696:17703] = '{32'hc226a81c, 32'hc2935c25, 32'h42a34411, 32'hc152441b, 32'hc2a1448a, 32'h415aff8a, 32'h426c896d, 32'h4202e8e4};
test_bias[2212:2212] = '{32'h41c0652a};
test_output[2212:2212] = '{32'h46112b0c};
test_input[17704:17711] = '{32'h42800aa6, 32'hc2c111a1, 32'hc29f7562, 32'h412aec27, 32'hc295f19f, 32'hc236ec3f, 32'hc186c4e2, 32'h41c74a37};
test_weights[17704:17711] = '{32'h425d2ee3, 32'hc2c48013, 32'h410ab582, 32'hc233a62a, 32'hc196dae8, 32'hc18cc6cc, 32'hc2b460fb, 32'h4186e247};
test_bias[2213:2213] = '{32'h418f8bb0};
test_output[2213:2213] = '{32'h467a758d};
test_input[17712:17719] = '{32'h42a570a4, 32'h419b2aff, 32'hc2200a8d, 32'hc2163069, 32'hc1db35d4, 32'hc2831c5c, 32'h427975e7, 32'h42630ec6};
test_weights[17712:17719] = '{32'h427244da, 32'hc2b1dc0a, 32'h428f6c2c, 32'h4204b9f6, 32'h4278ee28, 32'h426c88c7, 32'h42a45d99, 32'hc09150ac};
test_bias[2214:2214] = '{32'hc235acb8};
test_output[2214:2214] = '{32'hc4c6ae86};
test_input[17720:17727] = '{32'hc21af4e0, 32'h423bc938, 32'hc2a8d3c7, 32'h42c3ad29, 32'h42103f45, 32'hc22d5644, 32'hc29eb559, 32'hc1fc6311};
test_weights[17720:17727] = '{32'h427d94fe, 32'h4214cac7, 32'h422a9f01, 32'h419b97e6, 32'hc22cb2e2, 32'h42c57e7d, 32'h42711ef8, 32'hc26c60cd};
test_bias[2215:2215] = '{32'h422b9d34};
test_output[2215:2215] = '{32'hc62dbee1};
test_input[17728:17735] = '{32'h42ad6c1c, 32'h42ade758, 32'hc24d477c, 32'hc1c2035e, 32'hc14e9845, 32'h42388c54, 32'hc11059b7, 32'h4285fae5};
test_weights[17728:17735] = '{32'h4125d708, 32'h426c362d, 32'hc2765eee, 32'hc29dc3a1, 32'h41fe71ac, 32'hc180ab78, 32'h428b4d46, 32'hc29c7784};
test_bias[2216:2216] = '{32'hc193d4d2};
test_output[2216:2216] = '{32'h457e3027};
test_input[17736:17743] = '{32'h429dcf79, 32'hc25f2ed9, 32'h429faa47, 32'hc23d1ccb, 32'h42b7cefa, 32'hc085e712, 32'h41cadcb4, 32'h3f758f3b};
test_weights[17736:17743] = '{32'h42705766, 32'h42115d32, 32'hc28bf0ac, 32'hc2b4071b, 32'h41aaf459, 32'h41a44814, 32'h42c0cb32, 32'h40f511ae};
test_bias[2217:2217] = '{32'h42388f1d};
test_output[2217:2217] = '{32'h45b3f88b};
test_input[17744:17751] = '{32'hc2332691, 32'h4191de23, 32'hc287a539, 32'hc15452e6, 32'hc1ac0c64, 32'h411156af, 32'h42c51fd7, 32'h42ad0ef7};
test_weights[17744:17751] = '{32'h42c38e89, 32'h420694e1, 32'h4294a36e, 32'hc2abfc7b, 32'hc2bf574f, 32'h42985d51, 32'h41f86742, 32'hc20196c6};
test_bias[2218:2218] = '{32'h41ee2b8c};
test_output[2218:2218] = '{32'hc590a66e};
test_input[17752:17759] = '{32'h417431b1, 32'hc28bf53b, 32'hc0d466d6, 32'h41797844, 32'h4176f069, 32'h425efeaf, 32'h428cc3a5, 32'hc1644ce6};
test_weights[17752:17759] = '{32'h41b51c39, 32'hc1ac4a45, 32'hc2a98c84, 32'h40d88ce6, 32'h4201dd20, 32'h42b0b8ea, 32'h42842236, 32'hc09e57d1};
test_bias[2219:2219] = '{32'hbf1e33ad};
test_output[2219:2219] = '{32'h4645ef3d};
test_input[17760:17767] = '{32'h41c0fb1c, 32'hc052f064, 32'h425172fc, 32'h422a1f03, 32'hc20bbc32, 32'h40d65c0d, 32'hc200448b, 32'h42351381};
test_weights[17760:17767] = '{32'h42b24044, 32'hc28f1010, 32'h42aba002, 32'h4075777c, 32'hc253e5fe, 32'h4285e22b, 32'h41eed05f, 32'h42c02c64};
test_bias[2220:2220] = '{32'h421c92fd};
test_output[2220:2220] = '{32'h46479357};
test_input[17768:17775] = '{32'hc224f694, 32'hc2b35df9, 32'h42220f89, 32'hc251a677, 32'h4288e765, 32'hc2aa371b, 32'h42966fb6, 32'hc2a4f2e7};
test_weights[17768:17775] = '{32'hc2b5af36, 32'h42887b7d, 32'h4190c409, 32'h3f903009, 32'h429f2645, 32'hc24ca1a0, 32'h42575821, 32'hc0d717a2};
test_bias[2221:2221] = '{32'h425cf884};
test_output[2221:2221] = '{32'h464761b7};
test_input[17776:17783] = '{32'hc1be22d7, 32'hc27f83db, 32'h411677ee, 32'h42bd4ba1, 32'hc129451d, 32'h42917dd1, 32'hc2ae6498, 32'h42a5fbd6};
test_weights[17776:17783] = '{32'h429e7301, 32'hc19a9d70, 32'hbfb9928f, 32'hc2176760, 32'hc24acdf4, 32'hc2b5dd9e, 32'hc2b1b83a, 32'h3f2989ae};
test_bias[2222:2222] = '{32'hc1fd9243};
test_output[2222:2222] = '{32'hc51f78ef};
test_input[17784:17791] = '{32'hc2b2390e, 32'h428d80d4, 32'hc21d3dd5, 32'h429bc436, 32'hc1fe1166, 32'hc2b01a7a, 32'h421e4246, 32'hc19d4b0b};
test_weights[17784:17791] = '{32'hc29814e3, 32'h422ab52e, 32'h426d4c5d, 32'hc13d6f84, 32'hc2208b97, 32'hc2be0da9, 32'h414550e7, 32'h421a2a9e};
test_bias[2223:2223] = '{32'hc286a8d0};
test_output[2223:2223] = '{32'h46779871};
test_input[17792:17799] = '{32'h4298efc4, 32'h417fa6f2, 32'h4202c356, 32'hc11abc31, 32'h41e123ea, 32'h42c70a67, 32'hc1262fde, 32'h4277b3b6};
test_weights[17792:17799] = '{32'hc245c602, 32'hc23e9f6f, 32'h4292860d, 32'h41fed5e9, 32'h42877eec, 32'h4210dbec, 32'h428a4339, 32'hc28c83ce};
test_bias[2224:2224] = '{32'h42797386};
test_output[2224:2224] = '{32'hc4f3e2db};
test_input[17800:17807] = '{32'hc2b50afd, 32'h42bcfab8, 32'h424fd5c8, 32'hc2ba8929, 32'hc2a2294d, 32'hc06cdbc5, 32'h41df652c, 32'hc0838bcc};
test_weights[17800:17807] = '{32'h423cb63d, 32'hc24e5c85, 32'hc2b9c21f, 32'hc2b92c27, 32'hc13b1021, 32'h4223a5cf, 32'h428d7b4f, 32'hc2c3bea7};
test_bias[2225:2225] = '{32'h42ad7e8f};
test_output[2225:2225] = '{32'hc501aec0};
test_input[17808:17815] = '{32'h42aeb406, 32'h420f9d1a, 32'hc22448a8, 32'h428d404e, 32'h4060f8cc, 32'h423127f5, 32'hc2c09916, 32'h42b4745a};
test_weights[17808:17815] = '{32'hc2b3bfe7, 32'hc23d5343, 32'hbff03eb2, 32'h42c14403, 32'hc2c7a0ad, 32'hc081cac4, 32'h42c625e4, 32'hc1f63331};
test_bias[2226:2226] = '{32'hc2ab6def};
test_output[2226:2226] = '{32'hc67377a6};
test_input[17816:17823] = '{32'h42ac4636, 32'h3ef30681, 32'h429801f9, 32'hc2bdd84e, 32'h408bb3d8, 32'h42a5813f, 32'h41f09cbe, 32'h4254fbd4};
test_weights[17816:17823] = '{32'hc2719211, 32'h429756ba, 32'h42b2f030, 32'hc1876d58, 32'hc28244ca, 32'hc2580e55, 32'h42219ca2, 32'hc172608c};
test_bias[2227:2227] = '{32'h42be67e1};
test_output[2227:2227] = '{32'hc47c6728};
test_input[17824:17831] = '{32'hc289ad00, 32'hc0c8f9bb, 32'hc2bc87a2, 32'h42a493d6, 32'h4270b7b3, 32'h42b13faf, 32'hc28943ad, 32'hc21f0e3d};
test_weights[17824:17831] = '{32'h42aace27, 32'h4155842a, 32'h42456980, 32'h427f2566, 32'hc1888a37, 32'h41c02c73, 32'hc1ead4bd, 32'hc1a86d0c};
test_bias[2228:2228] = '{32'h41efa07e};
test_output[2228:2228] = '{32'hc4acd216};
test_input[17832:17839] = '{32'hc20c956e, 32'hc29fb550, 32'hc2b211fa, 32'hbf86b35d, 32'h41b33ff9, 32'h41c2f8e0, 32'h4190dab3, 32'hc20d544a};
test_weights[17832:17839] = '{32'hc2a7eb44, 32'hc2a08607, 32'hc2c2c1a0, 32'h41d36213, 32'h4274baa1, 32'hc2c3290f, 32'h40a4b678, 32'h3f94d5aa};
test_bias[2229:2229] = '{32'h3ea5676b};
test_output[2229:2229] = '{32'h46852eee};
test_input[17840:17847] = '{32'hc2ae3ce5, 32'hc2ad70ea, 32'h428798ba, 32'hc1b1f246, 32'h4290d488, 32'hc1e071d4, 32'hc2b622ab, 32'h42b08274};
test_weights[17840:17847] = '{32'hc0f6a08a, 32'hc1ba9b7b, 32'hc1d82528, 32'h41429507, 32'h41633660, 32'hc1ab62a7, 32'h41fbb450, 32'hc21720f7};
test_bias[2230:2230] = '{32'hc2a191b1};
test_output[2230:2230] = '{32'hc57db24e};
test_input[17848:17855] = '{32'hc2899a8e, 32'h426dec6c, 32'hbf3c6e77, 32'h428a4503, 32'hc2c77dde, 32'h41b96b22, 32'hc2b286bb, 32'hc0f8d42d};
test_weights[17848:17855] = '{32'h429e77bb, 32'h424bba21, 32'hc1eb54a9, 32'hc28250fb, 32'hc272b384, 32'h4200caf5, 32'hc21dbe52, 32'h42a60d0f};
test_bias[2231:2231] = '{32'hc297c9e0};
test_output[2231:2231] = '{32'h4528409f};
test_input[17856:17863] = '{32'hc1b85bca, 32'h42b1eab4, 32'hc29800b9, 32'hc282eafb, 32'h42bd19d5, 32'h42a6e2a5, 32'hc27b0404, 32'hc2b2cc63};
test_weights[17856:17863] = '{32'hbf24265a, 32'hc2b8aa01, 32'hc2a080b2, 32'h420ac2da, 32'hc20b4b10, 32'hc296225f, 32'h42abebad, 32'hc13ebdcb};
test_bias[2232:2232] = '{32'h428f7034};
test_output[2232:2232] = '{32'hc68e0f79};
test_input[17864:17871] = '{32'h42038d67, 32'hc093209c, 32'hc2172fd5, 32'h429b83f0, 32'hc27c6ff4, 32'h427a9018, 32'hc2b33dbe, 32'hc294ed33};
test_weights[17864:17871] = '{32'h42709c48, 32'h4287a783, 32'h416c2e34, 32'h4192a93e, 32'hc0b479d0, 32'h42afd5f5, 32'hc1e3cd43, 32'hc2a4dfd3};
test_bias[2233:2233] = '{32'h41ef126e};
test_output[2233:2233] = '{32'h4685bb2d};
test_input[17872:17879] = '{32'h42ab3fab, 32'hc25c009f, 32'h4102b3e0, 32'hc2c31444, 32'hc23d730b, 32'h42380efa, 32'hbfffd8fc, 32'hc23ad15f};
test_weights[17872:17879] = '{32'h42b723e9, 32'h42c70615, 32'hc21f729c, 32'h4280637b, 32'hc2b005ee, 32'hc1861de9, 32'hc0a3106a, 32'h42bcb881};
test_bias[2234:2234] = '{32'h417bb19e};
test_output[2234:2234] = '{32'hc5a29e79};
test_input[17880:17887] = '{32'h429a80d7, 32'hc28b8dc9, 32'hc1d75b7d, 32'hc235e7a7, 32'h422be882, 32'h4211ec6a, 32'h4296e350, 32'hc28dd17e};
test_weights[17880:17887] = '{32'hc281c56a, 32'hc280fb6a, 32'h4295b7ce, 32'hc25678a9, 32'hbea622e1, 32'h4238dba1, 32'hc2b0d915, 32'h425e56ae};
test_bias[2235:2235] = '{32'h420723e8};
test_output[2235:2235] = '{32'hc60c906d};
test_input[17888:17895] = '{32'h40cfbb84, 32'hc29ec982, 32'hc208fc07, 32'hc2a0623d, 32'hc287832c, 32'hc21a7928, 32'h42b98c5a, 32'hc23e8d2a};
test_weights[17888:17895] = '{32'h42944fe3, 32'hc2c2b6f1, 32'h3f826391, 32'hc2a126c9, 32'h4248fe08, 32'h423320a1, 32'h42b2891d, 32'h424ad73d};
test_bias[2236:2236] = '{32'h428d5939};
test_output[2236:2236] = '{32'h467140fc};
test_input[17896:17903] = '{32'h413a6bec, 32'h42bea488, 32'hc24d88f9, 32'hc27831bb, 32'h42983ca4, 32'hc2b52271, 32'hc1dcc4f8, 32'h4190b69f};
test_weights[17896:17903] = '{32'hc2a17c6a, 32'h42c41ed4, 32'h42a5935b, 32'hc107cdf6, 32'hc1fa4027, 32'h413da85a, 32'hc2874071, 32'hc091637b};
test_bias[2237:2237] = '{32'hc179e1f9};
test_output[2237:2237] = '{32'h453b0f36};
test_input[17904:17911] = '{32'hc29b2ee3, 32'hc1ee4b7d, 32'hc294285c, 32'hc147aa90, 32'h4246d79d, 32'h42901e02, 32'hc2ab1516, 32'hc1a5b5a4};
test_weights[17904:17911] = '{32'hc210ffba, 32'hc2aa910a, 32'hc2ab58f2, 32'h4234fb2b, 32'hc258d3e3, 32'hc25bda68, 32'hc2843db0, 32'hc1bacd3f};
test_bias[2238:2238] = '{32'hc1946d08};
test_output[2238:2238] = '{32'h4625a38d};
test_input[17912:17919] = '{32'h425d302c, 32'h424dfd51, 32'h42832556, 32'hc147dc05, 32'h41fa8fb3, 32'hc29c17c1, 32'h4248fb2b, 32'hc2b427aa};
test_weights[17912:17919] = '{32'h4196b1aa, 32'h42b7e0ab, 32'h42298a7f, 32'h42513228, 32'hc2c297ff, 32'h427cee49, 32'hc0d878ac, 32'h42a245fb};
test_bias[2239:2239] = '{32'hc23c1885};
test_output[2239:2239] = '{32'hc5f2fd64};
test_input[17920:17927] = '{32'h41bf6b47, 32'hc1b7af34, 32'h428c64b0, 32'h41c4c787, 32'hc28feb92, 32'hc2c64403, 32'h4223deb0, 32'hc242d4e0};
test_weights[17920:17927] = '{32'h4235eb6b, 32'hc1ea6a14, 32'hc2a08fb4, 32'h41a8e202, 32'h423fdd71, 32'hc23ff1a2, 32'hc29c7afd, 32'hc116842c};
test_bias[2240:2240] = '{32'h42c5eb33};
test_output[2240:2240] = '{32'hc592cfd7};
test_input[17928:17935] = '{32'h42685fec, 32'hc27c4873, 32'h427d8e43, 32'hc2211708, 32'hc24e69be, 32'hc14bde1b, 32'hc243fc67, 32'h4284e715};
test_weights[17928:17935] = '{32'h42678d39, 32'hc267ce0d, 32'hc2b02807, 32'hc2a62d9e, 32'h4257f630, 32'hc1f2187d, 32'h4295a3a7, 32'hc1da4fad};
test_bias[2241:2241] = '{32'h40dd5891};
test_output[2241:2241] = '{32'hc5413e2d};
test_input[17936:17943] = '{32'hc289c8bf, 32'h40e1eeaf, 32'hc277551f, 32'h41de23cd, 32'hc255bcf1, 32'hc1d05241, 32'hc180fd30, 32'hc2380290};
test_weights[17936:17943] = '{32'h3e3f8c63, 32'hc29a0a87, 32'h4157b9c3, 32'h3f830fee, 32'h42a6f18d, 32'h428282af, 32'h42c20cf5, 32'hc29c4038};
test_bias[2242:2242] = '{32'h4227255d};
test_output[2242:2242] = '{32'hc5aa50ee};
test_input[17944:17951] = '{32'h425c0f4e, 32'hc13116fe, 32'h423290fb, 32'hc28c9b6d, 32'hc24fa712, 32'h42346903, 32'h42693265, 32'hc24674ec};
test_weights[17944:17951] = '{32'h428bcd23, 32'h42a8762d, 32'hc2825bb0, 32'h42a7aae5, 32'h41d76b81, 32'hc20fa4d1, 32'h41e9292a, 32'hc295efec};
test_bias[2243:2243] = '{32'hc23117e0};
test_output[2243:2243] = '{32'hc55cd676};
test_input[17952:17959] = '{32'h414bfa6e, 32'hc2a14ff6, 32'hc1de7a7e, 32'hc279beff, 32'h419ee360, 32'hc2b23b1c, 32'h409ae62e, 32'hc13468bd};
test_weights[17952:17959] = '{32'hc298d7b1, 32'h415e0183, 32'hc216108c, 32'h41d88cde, 32'hc1bea346, 32'h416a5c1e, 32'hc2702814, 32'hc2906d5d};
test_bias[2244:2244] = '{32'h428189fb};
test_output[2244:2244] = '{32'hc575a5f1};
test_input[17960:17967] = '{32'h42908cd7, 32'hc0ccca26, 32'hc2bdcabc, 32'h3f9bcf28, 32'hc27b1eb9, 32'hc212f05a, 32'hc2210af0, 32'hc270d301};
test_weights[17960:17967] = '{32'h3f33c730, 32'h405be0c5, 32'hc130d029, 32'h4285cb38, 32'hc18e165f, 32'hc27a8cd2, 32'hc1f504ca, 32'hc1e0671f};
test_bias[2245:2245] = '{32'h42bfce8c};
test_output[2245:2245] = '{32'h45ed454d};
test_input[17968:17975] = '{32'hc280c452, 32'hc2a7d8e0, 32'h4289a66d, 32'hc2671358, 32'hc2a69583, 32'hc29f70ea, 32'h428cbd1f, 32'h417a7af1};
test_weights[17968:17975] = '{32'hc26a8b1f, 32'h420d074a, 32'hc2953199, 32'h4190444c, 32'h41c9844b, 32'h42c2bb04, 32'hc0e1d0c9, 32'hc21c4d41};
test_bias[2246:2246] = '{32'hc20db8a1};
test_output[2246:2246] = '{32'hc67faddb};
test_input[17976:17983] = '{32'hc2b22b86, 32'h420641ce, 32'hc2b76928, 32'h41053305, 32'hc2b9d1f3, 32'h42b11e6e, 32'hc2963571, 32'hc230c8cf};
test_weights[17976:17983] = '{32'hc138ec90, 32'h429ad3b3, 32'hc203144d, 32'h42c71593, 32'hc1c95a7f, 32'hc1b7da91, 32'hc2be7177, 32'h41d497f4};
test_bias[2247:2247] = '{32'hc13a07a2};
test_output[2247:2247] = '{32'h465689ed};
test_input[17984:17991] = '{32'hc1ec4297, 32'hc226edf2, 32'h42c13da3, 32'hc1ce3cc2, 32'h4263cb78, 32'h42987690, 32'h42949575, 32'h4275365e};
test_weights[17984:17991] = '{32'h425a8ee5, 32'h425c0823, 32'h4276f176, 32'h427104fa, 32'hc09c8273, 32'hc28039ec, 32'h429c622c, 32'h428d01fe};
test_bias[2248:2248] = '{32'h428f8b68};
test_output[2248:2248] = '{32'h45ad19fc};
test_input[17992:17999] = '{32'h42b3ed19, 32'hc188c55b, 32'h42ac7f1f, 32'hc292ecc6, 32'h42a059f4, 32'h429bd36b, 32'hc2b55e96, 32'hc2483681};
test_weights[17992:17999] = '{32'hc27857f6, 32'h41513b33, 32'h425f5a05, 32'hc2162144, 32'hc16e2613, 32'hc2626587, 32'hc28b1a77, 32'h4126081a};
test_bias[2249:2249] = '{32'h41e83b19};
test_output[2249:2249] = '{32'h44f73c55};
test_input[18000:18007] = '{32'h4223216a, 32'hc20b99ed, 32'hc23c363c, 32'hc2c43110, 32'hc2ae2ecc, 32'h41eb69f5, 32'hc1eda8b4, 32'hc287cf53};
test_weights[18000:18007] = '{32'hc2aeebbf, 32'hc1f0625e, 32'hc23c8766, 32'hc2ba6f51, 32'h42618132, 32'h4288f02f, 32'h3ff4e822, 32'h40882242};
test_bias[2250:2250] = '{32'h41831dc6};
test_output[2250:2250] = '{32'h45af9b0d};
test_input[18008:18015] = '{32'hc08d6718, 32'h41039feb, 32'hc20eaae3, 32'h42980b64, 32'hc2a3517a, 32'hc20965d4, 32'hc2b56753, 32'h426b1b42};
test_weights[18008:18015] = '{32'h40b11bf7, 32'h41a1e912, 32'hc2a04e9a, 32'h40f93f5a, 32'hc26819da, 32'hc29aa80d, 32'h425f7608, 32'hc1fb530d};
test_bias[2251:2251] = '{32'hc267c1ca};
test_output[2251:2251] = '{32'h457aff43};
test_input[18016:18023] = '{32'hc2c42cf0, 32'h42886306, 32'hc2b91e42, 32'hc1831b43, 32'hc24018fd, 32'h4257eb24, 32'hc23723d0, 32'hc2b6f11d};
test_weights[18016:18023] = '{32'hc2b64374, 32'h4205ab69, 32'h413d435c, 32'h426cd6c3, 32'h41b05caa, 32'h41f6b830, 32'h420b3258, 32'hc286f258};
test_bias[2252:2252] = '{32'h41ea3c5a};
test_output[2252:2252] = '{32'h46607998};
test_input[18024:18031] = '{32'h422ba9de, 32'hc1d370e9, 32'h424d6afe, 32'h42a8cf82, 32'hc2b89a62, 32'h4203290f, 32'hc20b4aa1, 32'h429a2561};
test_weights[18024:18031] = '{32'hc2be0555, 32'hc25cc86c, 32'h429b96e8, 32'hc2c7ed7f, 32'h4221d360, 32'hc2810604, 32'hc1c578b6, 32'h426f92bb};
test_bias[2253:2253] = '{32'hc2adb57c};
test_output[2253:2253] = '{32'hc5eb0d4f};
test_input[18032:18039] = '{32'h4296a3f9, 32'hc20ea899, 32'h420c651f, 32'hc26b5729, 32'h4277e8e0, 32'h428c44fe, 32'hc18f568b, 32'hc2881c72};
test_weights[18032:18039] = '{32'hc0deaadd, 32'h41e76739, 32'hc218576e, 32'hc2bcd4b7, 32'h41be8dfb, 32'hc0881f8c, 32'h428e07cb, 32'hc06f0405};
test_bias[2254:2254] = '{32'h422bd944};
test_output[2254:2254] = '{32'h453311e8};
test_input[18040:18047] = '{32'hc2bfd8f3, 32'h4272d312, 32'hc2af7400, 32'h428252a3, 32'h428fe80f, 32'h4240d23c, 32'h41c07f6a, 32'hc11144bf};
test_weights[18040:18047] = '{32'hc23a2ede, 32'hc1271791, 32'hc1d421de, 32'h426092f6, 32'h42bfd7f8, 32'hc281be3e, 32'h42a47cc9, 32'h421dc527};
test_bias[2255:2255] = '{32'hc21f2c2e};
test_output[2255:2255] = '{32'h466d0d0e};
test_input[18048:18055] = '{32'hc2a55ea1, 32'h40edd9da, 32'hc2653656, 32'h42bd22f5, 32'hc2c37757, 32'hc2c0ff88, 32'hc1b23dc7, 32'hc1a4749d};
test_weights[18048:18055] = '{32'h42b888bc, 32'h42010d4d, 32'h418cc589, 32'h4227b885, 32'h427eaa10, 32'hc2b9229a, 32'hc27dc128, 32'h411ebff1};
test_bias[2256:2256] = '{32'hc113d592};
test_output[2256:2256] = '{32'hc4026dfc};
test_input[18056:18063] = '{32'hc2be7792, 32'h426d1a12, 32'h4225238f, 32'h4272b704, 32'hbf87e4b2, 32'h4244841f, 32'hc1188381, 32'h41421a12};
test_weights[18056:18063] = '{32'hc2c3105f, 32'hc247ed66, 32'h42ad60b8, 32'hc1d06fa4, 32'h419e9da1, 32'hc29cedf8, 32'h425751a7, 32'h423908bd};
test_bias[2257:2257] = '{32'h428e22a2};
test_output[2257:2257] = '{32'h458eb63c};
test_input[18064:18071] = '{32'hc1febdab, 32'hbf567366, 32'hc1387d2e, 32'hc0e3de73, 32'hc1a35625, 32'hc2175079, 32'hc29600cd, 32'hc29bcfc7};
test_weights[18064:18071] = '{32'hc1a59bfa, 32'hc0f18f5c, 32'hc286bb58, 32'hc2b34d66, 32'hc2ad48fc, 32'hc2a5eff6, 32'h428588ca, 32'h42997fcc};
test_bias[2258:2258] = '{32'h42a7fa4b};
test_output[2258:2258] = '{32'hc574aa70};
test_input[18072:18079] = '{32'h41d22cd9, 32'h429e472c, 32'h428c4843, 32'hc1eb32f0, 32'h429848a2, 32'h42bb0ff7, 32'hc2a2f90e, 32'hc21e0878};
test_weights[18072:18079] = '{32'hc25f13e2, 32'h421c487e, 32'hbffa992a, 32'hc288f471, 32'hc2c4d65a, 32'hc190caf9, 32'h4290e107, 32'hc158e9a7};
test_bias[2259:2259] = '{32'h42c18ca6};
test_output[2259:2259] = '{32'hc62b2930};
test_input[18080:18087] = '{32'hc0c55f3e, 32'h425b3b35, 32'hc28b465a, 32'hc2c72ba8, 32'hc11d5f2e, 32'hc2aac5bb, 32'h41b69c48, 32'hc0e94a3d};
test_weights[18080:18087] = '{32'h40d94acb, 32'h42be2856, 32'hc291363b, 32'hc247ecf9, 32'h42434399, 32'h4183dec6, 32'hc1918acb, 32'hc19caed4};
test_bias[2260:2260] = '{32'hc03ac28c};
test_output[2260:2260] = '{32'h464bbe92};
test_input[18088:18095] = '{32'hc244599b, 32'hc2bdee60, 32'h42bda8b1, 32'h42c54cf0, 32'h4285ca0a, 32'hc10dcef6, 32'h42c502d6, 32'h42ae741a};
test_weights[18088:18095] = '{32'hc1f52b52, 32'hc2b0041d, 32'hc0b40bd6, 32'hc2a418ec, 32'h4136fd55, 32'hc14b38b7, 32'h40b72c63, 32'hc2821fce};
test_bias[2261:2261] = '{32'hc1f4c81e};
test_output[2261:2261] = '{32'hc53d5dbb};
test_input[18096:18103] = '{32'h4293fa27, 32'hc219760b, 32'hc16c2c56, 32'hc2703a4e, 32'hc2203529, 32'h4102b0e0, 32'h417fcf1b, 32'h426941cb};
test_weights[18096:18103] = '{32'hc15711c8, 32'hc2591947, 32'h41828472, 32'h42327781, 32'h42b80bfc, 32'hc2774ca2, 32'hc1e812e8, 32'hc2680ec9};
test_bias[2262:2262] = '{32'h426bc3a4};
test_output[2262:2262] = '{32'hc6194d1e};
test_input[18104:18111] = '{32'hc21733de, 32'h42c7d172, 32'h428a9954, 32'h42ae496c, 32'h42065d7a, 32'h42b1a564, 32'h42ac890b, 32'h42a6fb06};
test_weights[18104:18111] = '{32'h422e881e, 32'hc11a32ac, 32'hc29180db, 32'h41ffb57f, 32'h42a5bed1, 32'hc032f1fa, 32'hc0f5eb9d, 32'h422ab122};
test_bias[2263:2263] = '{32'hc26da718};
test_output[2263:2263] = '{32'h43fdb337};
test_input[18112:18119] = '{32'hc1eabd97, 32'h41a9b7c8, 32'h41fbe1ae, 32'hc28d017b, 32'h42679e9c, 32'h428dbc38, 32'h42bf44fa, 32'h424347b1};
test_weights[18112:18119] = '{32'h429679e6, 32'hc2c58255, 32'hc29273e0, 32'hc2231d7a, 32'h41da360f, 32'hc1593e63, 32'h4215230b, 32'h4239bb4b};
test_bias[2264:2264] = '{32'h410da538};
test_output[2264:2264] = '{32'h452a555d};
test_input[18120:18127] = '{32'hc284364b, 32'hc2b7c2f1, 32'hc243eea7, 32'hc154de48, 32'hbf3dcc79, 32'h42aecfee, 32'hc28dfc0a, 32'h41757a03};
test_weights[18120:18127] = '{32'h424d7370, 32'h3f9afc7b, 32'hc25345b0, 32'h42382325, 32'hc239c136, 32'hc29febe8, 32'h42a5e47a, 32'hc2417b0f};
test_bias[2265:2265] = '{32'h428b81bd};
test_output[2265:2265] = '{32'hc66b1db7};
test_input[18128:18135] = '{32'h42c42822, 32'hc207be38, 32'h411010e2, 32'hc1e2ff24, 32'h41b63688, 32'hc261b244, 32'hc23380fc, 32'h429c27d1};
test_weights[18128:18135] = '{32'hc2890fde, 32'hc2a00f41, 32'h4162b4f4, 32'hc2187359, 32'hc2862f47, 32'hc0bcc15b, 32'hc200444c, 32'h417d576a};
test_bias[2266:2266] = '{32'hc24f689c};
test_output[2266:2266] = '{32'hc4ab0cb3};
test_input[18136:18143] = '{32'h429f9284, 32'hc20663f9, 32'hc248f170, 32'h42bf3986, 32'h42b763a5, 32'h427f71b5, 32'h40c26244, 32'h412cb5dd};
test_weights[18136:18143] = '{32'hc2a8ab60, 32'h3da0abbf, 32'hc2b00222, 32'hc28d5d12, 32'h42c24de2, 32'h422d7c1a, 32'hc29ba870, 32'hc29bdfa2};
test_bias[2267:2267] = '{32'hc1e72a10};
test_output[2267:2267] = '{32'h449e5454};
test_input[18144:18151] = '{32'hc204c456, 32'hc20fce08, 32'hc2800491, 32'h42ba4423, 32'h42aa9fae, 32'h40bf593d, 32'hc28e216f, 32'hc2a21390};
test_weights[18144:18151] = '{32'hc2baf82e, 32'hc242a8a3, 32'hc1d61e12, 32'h42bb0ceb, 32'hc26cae07, 32'h424f6fa8, 32'h41e982c9, 32'hc1d68b9a};
test_bias[2268:2268] = '{32'hc0dd21de};
test_output[2268:2268] = '{32'h462618dd};
test_input[18152:18159] = '{32'h42b5193d, 32'h42a86ef0, 32'h42a76380, 32'h420d6be7, 32'h4289f9fe, 32'h41b8ac55, 32'h42963fa8, 32'hc1d6d279};
test_weights[18152:18159] = '{32'h41c5da9c, 32'h4259519e, 32'hc2b2c5a4, 32'hc1de2328, 32'h42652550, 32'h42b159e3, 32'h41e10766, 32'h42595137};
test_bias[2269:2269] = '{32'h40977ea9};
test_output[2269:2269] = '{32'h459c914f};
test_input[18160:18167] = '{32'hc26d5e43, 32'h4272e838, 32'hc210b67e, 32'h42a7d8b6, 32'hc1032239, 32'hc2aadb44, 32'hc2479392, 32'h42c13645};
test_weights[18160:18167] = '{32'hc2a47508, 32'hc16691f9, 32'h41bda58c, 32'hc2a4a306, 32'h42bdd9d1, 32'h4298443a, 32'hc1f73ade, 32'h4105a2b2};
test_bias[2270:2270] = '{32'hc25fc0eb};
test_output[2270:2270] = '{32'hc608ba8e};
test_input[18168:18175] = '{32'h42c2eaf4, 32'h42bb100e, 32'h42947942, 32'h4239fc30, 32'hc0f66774, 32'h41ea81be, 32'hc2c76b60, 32'hc2be9bcb};
test_weights[18168:18175] = '{32'hc2b168df, 32'hc2bda95d, 32'hc2887b00, 32'h41a1dddc, 32'h42178c79, 32'hc2c6b07c, 32'hc24c5fc0, 32'h42beeff1};
test_bias[2271:2271] = '{32'hc19f351e};
test_output[2271:2271] = '{32'hc6e18769};
test_input[18176:18183] = '{32'hc2b6602c, 32'h42b2cea4, 32'h4091feaf, 32'hc28d8ac0, 32'hc239344f, 32'hc0daa1f3, 32'h428f3ac3, 32'hc22643ff};
test_weights[18176:18183] = '{32'h424eea5d, 32'h42907a89, 32'hc199a1e0, 32'h42bdaf1c, 32'hc2a1a5f7, 32'h42c323ea, 32'h424fdcf9, 32'hbfb7fd9c};
test_bias[2272:2272] = '{32'h419f22c4};
test_output[2272:2272] = '{32'h44e35063};
test_input[18184:18191] = '{32'h42a8ce09, 32'hc2ac2eb2, 32'h416bf4e4, 32'h41c49596, 32'h4138dccb, 32'hc1644c9e, 32'h42bd04b1, 32'hc20d6c57};
test_weights[18184:18191] = '{32'hc2c40bb1, 32'h42714568, 32'hc234b9a5, 32'h41b47add, 32'hc2207ef2, 32'hc27cf915, 32'hc190fe98, 32'h42a05402};
test_bias[2273:2273] = '{32'h41fbbcfe};
test_output[2273:2273] = '{32'hc689ee0f};
test_input[18192:18199] = '{32'hbfbe7ec4, 32'hc1c309bd, 32'h412f37a1, 32'h429dea5f, 32'hc2a9f1f8, 32'hc222963f, 32'hc0a5f28c, 32'hc2be4974};
test_weights[18192:18199] = '{32'h41c5915a, 32'h42c7f09e, 32'h4286f0af, 32'hc2b60d93, 32'h41eda319, 32'hc1852848, 32'h42bb305d, 32'hc271e1d3};
test_bias[2274:2274] = '{32'hc29fb75f};
test_output[2274:2274] = '{32'hc5ae6e08};
test_input[18200:18207] = '{32'hc1963b8c, 32'hc2555870, 32'h4294f489, 32'hc284c434, 32'hc1a95af1, 32'hc27a408d, 32'hc202976b, 32'h427ad3a6};
test_weights[18200:18207] = '{32'h42ba1f98, 32'h418b8425, 32'hc1d5af0c, 32'h427bb7a4, 32'hc19c8680, 32'hc219b8a7, 32'hc283523b, 32'hc1c31070};
test_bias[2275:2275] = '{32'h42619d0d};
test_output[2275:2275] = '{32'hc5a75789};
test_input[18208:18215] = '{32'h3f8f75b6, 32'hc2b3b7c4, 32'hc241ed81, 32'h427f67e6, 32'h40964d08, 32'hc2673d2e, 32'h421f14ee, 32'hc24989bd};
test_weights[18208:18215] = '{32'hc28ff67c, 32'h42bdd6fa, 32'hc20c9ff0, 32'hc215b7ff, 32'h42784d92, 32'h41bf3005, 32'hc2374457, 32'h421e16d1};
test_bias[2276:2276] = '{32'h421a0dc3};
test_output[2276:2276] = '{32'hc65d4215};
test_input[18216:18223] = '{32'hc248835e, 32'hc2b0fe84, 32'hc087a535, 32'h426596ef, 32'h42823b4d, 32'h4283bde7, 32'hc2b10eb1, 32'hc2a7d2e8};
test_weights[18216:18223] = '{32'hc0eb15a1, 32'h423acf6a, 32'hc2c4f351, 32'h42c49792, 32'h42822963, 32'h429211f1, 32'hc043296e, 32'h42a09848};
test_bias[2277:2277] = '{32'hc2ad4c44};
test_output[2277:2277] = '{32'h4595a54b};
test_input[18224:18231] = '{32'hc223e54b, 32'h417f404c, 32'h419cd67d, 32'hc2883f3a, 32'h4140b9b0, 32'h4297cebd, 32'h42769f7a, 32'hc2b6f92f};
test_weights[18224:18231] = '{32'hc2988a63, 32'hc203206e, 32'hc1df363f, 32'h427f2b3a, 32'h412b7017, 32'h41e7c5de, 32'hc2747cd6, 32'h3f9ec91a};
test_bias[2278:2278] = '{32'h428363e1};
test_output[2278:2278] = '{32'hc56c2d24};
test_input[18232:18239] = '{32'hc2707bb0, 32'hc2abca01, 32'hc1d90f81, 32'hc2b49b0e, 32'hc1febe02, 32'hc2b4c417, 32'h4108f78a, 32'h416aee9a};
test_weights[18232:18239] = '{32'hc26c2831, 32'h42bf7aad, 32'h40cac393, 32'h42b2faeb, 32'h426aea24, 32'hc25d3145, 32'h42ac38b5, 32'h428c6814};
test_bias[2279:2279] = '{32'hc187e489};
test_output[2279:2279] = '{32'hc5fb820c};
test_input[18240:18247] = '{32'hc1983642, 32'h424e5192, 32'hc259608d, 32'h40977aec, 32'hc1b65487, 32'hc23c2dae, 32'hc2c5187a, 32'h42748fb8};
test_weights[18240:18247] = '{32'h418174a9, 32'hc20ff2ea, 32'h4272477a, 32'h415d9a70, 32'h427a6ffe, 32'h425bfed3, 32'hc1e5619a, 32'hc294ae54};
test_bias[2280:2280] = '{32'hc27547a0};
test_output[2280:2280] = '{32'hc62ec596};
test_input[18248:18255] = '{32'hc2822cbd, 32'h429d2634, 32'hc1b8fc75, 32'hc21aafa6, 32'h4227594b, 32'h429cea06, 32'h4298d58d, 32'h4129543f};
test_weights[18248:18255] = '{32'hc0d86c0c, 32'hc2477b4d, 32'h414d23e2, 32'hc242d2cb, 32'hc1938015, 32'h41fb03ed, 32'hc29a9294, 32'h429ca4c6};
test_bias[2281:2281] = '{32'hc110fdff};
test_output[2281:2281] = '{32'hc5a538c0};
test_input[18256:18263] = '{32'h42b17d39, 32'h41c68118, 32'hc25b3429, 32'h41d063b4, 32'h42a660f6, 32'h4227325d, 32'h425c347d, 32'hc2aae272};
test_weights[18256:18263] = '{32'h42bb148a, 32'hc2afeac4, 32'h42a502eb, 32'hc2903fc7, 32'h40beb5c7, 32'hc2c70e03, 32'hc286030c, 32'h42ae5a3b};
test_bias[2282:2282] = '{32'h423cf895};
test_output[2282:2282] = '{32'hc66aefa8};
test_input[18264:18271] = '{32'h42c52e84, 32'hc2174fc5, 32'h41b25633, 32'hc285b285, 32'hc26c5a34, 32'hc2ad8a3f, 32'hc26f1602, 32'h42bde699};
test_weights[18264:18271] = '{32'h428f52b0, 32'hc1f2b090, 32'h42b58084, 32'h40dcffe3, 32'hc2c47ffe, 32'hc24ee72f, 32'hc1e3f690, 32'h4217e7c9};
test_bias[2283:2283] = '{32'hc260f1e7};
test_output[2283:2283] = '{32'h46c5d126};
test_input[18272:18279] = '{32'hc199ac3b, 32'hc2b278d3, 32'hc29791e3, 32'h420a722f, 32'hc10ded83, 32'h41933f61, 32'hc1157f91, 32'hc22c032d};
test_weights[18272:18279] = '{32'h422f2d64, 32'h3f303fdb, 32'hc2674460, 32'h42bc3f6f, 32'h3fd4346c, 32'hc1cd6212, 32'h41dbd8e1, 32'h4288b755};
test_bias[2284:2284] = '{32'h413f6bcb};
test_output[2284:2284] = '{32'h453f9114};
test_input[18280:18287] = '{32'h421a99e3, 32'hc1bc5bfd, 32'h42864961, 32'hc189a0fd, 32'h424cd1e2, 32'hc1eb601b, 32'h41bc20ea, 32'hc2bc49ad};
test_weights[18280:18287] = '{32'hc16e1ce5, 32'h425eac1a, 32'h426aedd3, 32'hc28c1052, 32'hc20c7b8d, 32'h42a5bbbd, 32'hc264b84e, 32'h416bc152};
test_bias[2285:2285] = '{32'h42ac81af};
test_output[2285:2285] = '{32'hc5623a48};
test_input[18288:18295] = '{32'h42921a11, 32'h427157bd, 32'hc1c8e6a3, 32'h42101723, 32'h40461f08, 32'h42c2138e, 32'h404aa4bc, 32'hc2abf291};
test_weights[18288:18295] = '{32'hc29d35af, 32'hc1d34171, 32'h429b90d0, 32'hc156dd30, 32'hc16c9250, 32'hc22e6d38, 32'h42075aa8, 32'h42a622e9};
test_bias[2286:2286] = '{32'h41b6ebe0};
test_output[2286:2286] = '{32'hc6a48af3};
test_input[18296:18303] = '{32'hc1f3b364, 32'h421cbd78, 32'hc2428c4c, 32'hc28f0ec8, 32'h4200a9e2, 32'h42b0db1e, 32'h410e18eb, 32'hc1c9bcbf};
test_weights[18296:18303] = '{32'hc29f907b, 32'h42881008, 32'hc20d1286, 32'hc25157a1, 32'h41918181, 32'h42ade5d1, 32'h42968ad3, 32'hc1902018};
test_bias[2287:2287] = '{32'h42b04b60};
test_output[2287:2287] = '{32'h469c8f6d};
test_input[18304:18311] = '{32'hc1b8dae5, 32'h426d5738, 32'h41308b61, 32'h42599ee0, 32'h41e6e4de, 32'hc226ba90, 32'hc185e946, 32'hc0f63115};
test_weights[18304:18311] = '{32'h41501162, 32'hc299752e, 32'h41bd2e3e, 32'hc24ce5fa, 32'h41935f8c, 32'hc2535afe, 32'hc1b2b7ae, 32'hc2a6a4b1};
test_bias[2288:2288] = '{32'hc28af42b};
test_output[2288:2288] = '{32'hc56738ab};
test_input[18312:18319] = '{32'hc2401b76, 32'hc20c4f55, 32'hc223803c, 32'hc27e47bb, 32'h41ef3aba, 32'hc1d8824d, 32'hc2834869, 32'h419364dd};
test_weights[18312:18319] = '{32'h42773985, 32'h41a0189b, 32'hc0cb9f9b, 32'hc25a415b, 32'hc1e81a9f, 32'h40dedb6b, 32'h427f4512, 32'hc1535707};
test_bias[2289:2289] = '{32'hc1ca2828};
test_output[2289:2289] = '{32'hc5aa7aff};
test_input[18320:18327] = '{32'h41512cea, 32'h40fe8330, 32'h4226888f, 32'h42b45e6e, 32'hc28a9d2e, 32'h4205e20a, 32'hc244a75c, 32'hc298a38c};
test_weights[18320:18327] = '{32'h4165909d, 32'h4246c855, 32'h42610c0d, 32'hc23709b7, 32'hc2b65392, 32'h3f1ce8aa, 32'h41e2b20d, 32'hc19fa693};
test_bias[2290:2290] = '{32'hc106e8c8};
test_output[2290:2290] = '{32'h45a45533};
test_input[18328:18335] = '{32'h42b3995b, 32'h422a2da4, 32'hc240c024, 32'h42819f06, 32'h42bb50c0, 32'hbf2e7804, 32'h41dcba60, 32'hc019d45d};
test_weights[18328:18335] = '{32'hc2470aca, 32'h40e63114, 32'h42779285, 32'h41dcadc3, 32'hc0eba106, 32'h4245bb74, 32'hc0ad0519, 32'hc2bac9fa};
test_bias[2291:2291] = '{32'hc23a8d9a};
test_output[2291:2291] = '{32'hc5bd1e4c};
test_input[18336:18343] = '{32'h42071bc6, 32'h4106e20c, 32'h429aa0d5, 32'h424d694e, 32'h42b40e5e, 32'hc18a0733, 32'h42961ef0, 32'h42a80ff7};
test_weights[18336:18343] = '{32'h410d707f, 32'h41f61b5f, 32'hc2a4798d, 32'h3f8363df, 32'hc18e34b0, 32'hc1403646, 32'hc22dc109, 32'h42bb751b};
test_bias[2292:2292] = '{32'h42b15c6c};
test_output[2292:2292] = '{32'hc518435f};
test_input[18344:18351] = '{32'h420e4192, 32'hc2793609, 32'hc2a0a5cc, 32'h424d49dd, 32'h42967893, 32'h421140c4, 32'hc19570b3, 32'hc212c36e};
test_weights[18344:18351] = '{32'h428423d5, 32'hc1d8789f, 32'h429041fd, 32'h42779ffa, 32'h42c16216, 32'h42b7dc4f, 32'h41345a28, 32'h427c37fb};
test_bias[2293:2293] = '{32'h4230dbc6};
test_output[2293:2293] = '{32'h46154068};
test_input[18352:18359] = '{32'hc1f40e50, 32'h41fb6903, 32'hc0fbd3ac, 32'hc292605d, 32'h41f706aa, 32'hc2c664bd, 32'h41ff3173, 32'h42bf6d67};
test_weights[18352:18359] = '{32'h42a8ecdb, 32'h42b9fc49, 32'h4264062a, 32'h3ea6b226, 32'hc2c478b3, 32'hc1da13e7, 32'hc2279847, 32'h4211dbd4};
test_bias[2294:2294] = '{32'h4280c10e};
test_output[2294:2294] = '{32'h44dc406b};
test_input[18360:18367] = '{32'hc2af0d37, 32'hc203a7a5, 32'hc20d3901, 32'hc2c6b83f, 32'hc1b62746, 32'h41746574, 32'hc2aece60, 32'hc2ab8a30};
test_weights[18360:18367] = '{32'h42b61339, 32'hc29a2de2, 32'hc2b730dd, 32'hc27e27ef, 32'hc21ab14f, 32'hbf99ece8, 32'h41c07f2a, 32'h428b6f39};
test_bias[2295:2295] = '{32'hc2c13a62};
test_output[2295:2295] = '{32'hc5480eec};
test_input[18368:18375] = '{32'hc25d80a0, 32'h41f0fd14, 32'hc1b0864f, 32'hc196dda1, 32'h42ab7e2d, 32'h42009add, 32'h4067c9db, 32'hc2539d36};
test_weights[18368:18375] = '{32'hc25c4aa7, 32'hc2458b46, 32'hc1b6c35f, 32'h426eb372, 32'h4107f5a2, 32'hc28d03cb, 32'hc24b8acd, 32'h4118a03a};
test_bias[2296:2296] = '{32'hc1431065};
test_output[2296:2296] = '{32'hc4a25562};
test_input[18376:18383] = '{32'h4267fd91, 32'hc2b9373c, 32'h42649b2a, 32'hc2b51e12, 32'h42ab67ce, 32'h424426be, 32'h4249c4ca, 32'h40fd2249};
test_weights[18376:18383] = '{32'h42c67b01, 32'h42c21243, 32'hc28f6d96, 32'hc07a2a80, 32'h41940610, 32'hc253a686, 32'hc2a0f9c4, 32'h4215ec98};
test_bias[2297:2297] = '{32'hc128214a};
test_output[2297:2297] = '{32'hc637b87b};
test_input[18384:18391] = '{32'h42954707, 32'hc1cf478c, 32'h424b5d1d, 32'h4221df5a, 32'hc28126a8, 32'h42064003, 32'hc210f685, 32'hc2ba35df};
test_weights[18384:18391] = '{32'h4119999d, 32'h423bf16d, 32'hc076376b, 32'h428764ae, 32'h42be553e, 32'h42ad8a2e, 32'h40dbd0f5, 32'h42c6f9d3};
test_bias[2298:2298] = '{32'h42b472f7};
test_output[2298:2298] = '{32'hc625ceb8};
test_input[18392:18399] = '{32'h4135a3e1, 32'hc2479a09, 32'h424f4c4a, 32'hc21aeef1, 32'hc2b9bd6b, 32'hc1983216, 32'hc0684a13, 32'h4174aacd};
test_weights[18392:18399] = '{32'h415cad28, 32'h42afea87, 32'h40a570c0, 32'h42ac2e6c, 32'h425907a8, 32'hc2c20a38, 32'hc24820c7, 32'hc262a51d};
test_bias[2299:2299] = '{32'h428e1405};
test_output[2299:2299] = '{32'hc62d88aa};
test_input[18400:18407] = '{32'hc293f39a, 32'hc2c4f17b, 32'h41f4d3d0, 32'h41b9597c, 32'h42bab665, 32'hc21c4412, 32'hc2808d2d, 32'hc2a47482};
test_weights[18400:18407] = '{32'h425b4dc2, 32'hc11eaf06, 32'hc2b64aed, 32'hc2c12a88, 32'h42946b7e, 32'h41e57718, 32'hc234d176, 32'hc2ae7359};
test_bias[2300:2300] = '{32'h4225f146};
test_output[2300:2300] = '{32'h45f4640b};
test_input[18408:18415] = '{32'h427d3a48, 32'h42c0989e, 32'h4293f42a, 32'h429a17d9, 32'hc2b7fba2, 32'hc2b37d06, 32'hc2a2bb08, 32'hc29ccf16};
test_weights[18408:18415] = '{32'hc28ed2db, 32'h4210f613, 32'hc1fd4f6c, 32'hc21b85e5, 32'hc2b1c3c0, 32'hc1a58892, 32'hc2a118de, 32'hc2aa39bf};
test_bias[2301:2301] = '{32'hc1ad1bf1};
test_output[2301:2301] = '{32'h4683cb9e};
test_input[18416:18423] = '{32'h4286cbea, 32'hc227840c, 32'h414a4c6c, 32'hc1ab8062, 32'h42554e25, 32'h42c055e7, 32'h427ad40f, 32'hc2c32300};
test_weights[18416:18423] = '{32'hc00bff47, 32'hc22cf2aa, 32'h429467c5, 32'hc0dae30d, 32'hc16f7110, 32'h42868a42, 32'h403bba46, 32'hc2812428};
test_bias[2302:2302] = '{32'hc2af079e};
test_output[2302:2302] = '{32'h46677f10};
test_input[18424:18431] = '{32'h429d315c, 32'hc0bd61bd, 32'hc28c64e1, 32'hc20fb5df, 32'h42942a3f, 32'h41057f0d, 32'h413616f2, 32'h415cbc51};
test_weights[18424:18431] = '{32'hc21ba1fc, 32'hc2bc352a, 32'h4203c5d7, 32'hc1b65480, 32'hc2c451fa, 32'hc1bdc3a9, 32'hc25ae498, 32'h4291b424};
test_bias[2303:2303] = '{32'hc293a963};
test_output[2303:2303] = '{32'hc62e50d9};
test_input[18432:18439] = '{32'h428fed43, 32'h4246f845, 32'h4236b0cb, 32'hc28b6d6b, 32'h429c9aec, 32'hc28a72b9, 32'h41d55751, 32'hc266ce58};
test_weights[18432:18439] = '{32'hc107093e, 32'hc07e77a2, 32'h41813709, 32'hc203bc33, 32'hc2155a48, 32'hc155310c, 32'hc29b39cb, 32'hc2c4248d};
test_bias[2304:2304] = '{32'h4102fb0b};
test_output[2304:2304] = '{32'h456f0810};
test_input[18440:18447] = '{32'hc2aa23e8, 32'hc210277c, 32'hc26ce264, 32'hc2adfddc, 32'hc21a59eb, 32'hc260929f, 32'hc2adebda, 32'hc2839d4b};
test_weights[18440:18447] = '{32'h42051a2b, 32'hc097cabe, 32'hc2266843, 32'h42168a18, 32'h41b08252, 32'h427c6f42, 32'hc29dbcdb, 32'hc17130c3};
test_bias[2305:2305] = '{32'hc233c087};
test_output[2305:2305] = '{32'hc26c86aa};
test_input[18448:18455] = '{32'hc2b6e690, 32'h4110abe6, 32'h420a50d0, 32'hc2737f33, 32'hc22eeb5a, 32'hc2294b35, 32'hc2b39ba9, 32'h40e8297e};
test_weights[18448:18455] = '{32'hc1017afb, 32'h41825aa3, 32'hc25c7521, 32'h429507de, 32'hc28b62cf, 32'hc23e203e, 32'hc104a94a, 32'hc2bd1dfe};
test_bias[2306:2306] = '{32'hbfe4ef4d};
test_output[2306:2306] = '{32'hc3db29fd};
test_input[18456:18463] = '{32'hc2c478fb, 32'h42bef1c3, 32'hc27df507, 32'h429ed653, 32'h4125b16f, 32'h427c6418, 32'h4228b6bd, 32'h4261d1a9};
test_weights[18456:18463] = '{32'h4281b36b, 32'h428e9ffe, 32'hc21c17ca, 32'hc2903bed, 32'h421829e4, 32'hc201b690, 32'h41556802, 32'h422fd133};
test_bias[2307:2307] = '{32'h3f83706b};
test_output[2307:2307] = '{32'hc4b16b9c};
test_input[18464:18471] = '{32'h41d99340, 32'h42bf34e9, 32'h4186a2b9, 32'h428bd1aa, 32'h42913c4a, 32'hc2bf6432, 32'hc22c9fbb, 32'h4200378b};
test_weights[18464:18471] = '{32'hc28f01d8, 32'h420c967e, 32'h415673f1, 32'hc1c8d6a7, 32'h42211ee8, 32'hc1d2194f, 32'h426c80e7, 32'h411a15b5};
test_bias[2308:2308] = '{32'h42976abe};
test_output[2308:2308] = '{32'h45455030};
test_input[18472:18479] = '{32'hc2b62372, 32'hc2bafb5f, 32'h417edd9a, 32'h42a92e15, 32'hc14f1452, 32'h41ee9cea, 32'h4281eb04, 32'h4166a3f1};
test_weights[18472:18479] = '{32'h41977c84, 32'h4261af04, 32'hc2a1d453, 32'hc227ba42, 32'hc0ec9006, 32'hc2a4baab, 32'hc1265b94, 32'h42158168};
test_bias[2309:2309] = '{32'hc28e3da3};
test_output[2309:2309] = '{32'hc6610fce};
test_input[18480:18487] = '{32'hc219a769, 32'hc1b24dfb, 32'h3ea197b8, 32'h4277dacc, 32'h4110bc05, 32'h41841c17, 32'hc2952573, 32'hc29c903b};
test_weights[18480:18487] = '{32'h4131e47b, 32'hc22e9149, 32'hc23bf083, 32'hc26be734, 32'h42c1e514, 32'hc29e7f88, 32'h4237db96, 32'hc0ef78c4};
test_bias[2310:2310] = '{32'hc1fd3f02};
test_output[2310:2310] = '{32'hc5c8e6cf};
test_input[18488:18495] = '{32'h40ddfcae, 32'hc26edef2, 32'hc2694390, 32'h41da619f, 32'hc283e130, 32'hc2977011, 32'hc1a001c1, 32'h4285c06b};
test_weights[18488:18495] = '{32'hc29abb02, 32'h428f6eea, 32'h41f263a6, 32'h4243bd92, 32'hc2c5a2c0, 32'hc1da1bfe, 32'h42701825, 32'hc27ba7a1};
test_bias[2311:2311] = '{32'h42670246};
test_output[2311:2311] = '{32'hc4fc8965};
test_input[18496:18503] = '{32'hc0f66133, 32'hc26b7a2a, 32'h42abe261, 32'h3f908b6d, 32'hc297f61f, 32'hc26f403e, 32'h42c1b2c0, 32'h428e2b6b};
test_weights[18496:18503] = '{32'hc223b982, 32'h4192494b, 32'h41a5177a, 32'hc22c7128, 32'h4210e7a1, 32'h424f5726, 32'h42b0cd80, 32'hc1c9f5df};
test_bias[2312:2312] = '{32'h422285ef};
test_output[2312:2312] = '{32'h44efca6f};
test_input[18504:18511] = '{32'hc28fc396, 32'hc22b1f1f, 32'h420ed21e, 32'hc2b59a7d, 32'hc1ab3dae, 32'h426ece8b, 32'h4259542f, 32'h41bed175};
test_weights[18504:18511] = '{32'hc2b8da49, 32'hc225ba98, 32'h41a016a9, 32'hc21bceb4, 32'hc181f4fe, 32'h41e810f3, 32'h42c2526a, 32'h42b390ea};
test_bias[2313:2313] = '{32'h416afe99};
test_output[2313:2313] = '{32'h46ad4cd7};
test_input[18512:18519] = '{32'h42612244, 32'h4151bd82, 32'hc25230a4, 32'hc2bd5050, 32'h40dae254, 32'hbddc3fb1, 32'h42b2665f, 32'h428be005};
test_weights[18512:18519] = '{32'hc20f272a, 32'hc276b0bd, 32'h42b84997, 32'h420e4490, 32'h42a7161a, 32'h42349f69, 32'hc1b1c309, 32'h4244999f};
test_bias[2314:2314] = '{32'hc24e5896};
test_output[2314:2314] = '{32'hc60d93b4};
test_input[18520:18527] = '{32'hc23407f2, 32'hc246bb2e, 32'h4286cee2, 32'h42ac1f89, 32'hc2beca46, 32'hc0e37f4c, 32'hc1758ba4, 32'hc1a61948};
test_weights[18520:18527] = '{32'hc1b24e19, 32'hc213e882, 32'hc282b8ee, 32'hc1b0c9bd, 32'hc1e6d165, 32'h429352b0, 32'hbf7ea078, 32'hc200a816};
test_bias[2315:2315] = '{32'h427d9508};
test_output[2315:2315] = '{32'hc3f604a1};
test_input[18528:18535] = '{32'hc2ab30db, 32'h424f7d4c, 32'h42ae05cc, 32'h42891138, 32'hc2acc88c, 32'hc1ebe2e6, 32'hc2c5bb70, 32'h40af242f};
test_weights[18528:18535] = '{32'hc20ff00b, 32'h42a15ac1, 32'h42ab8152, 32'hc297a6d8, 32'h4286a9f6, 32'h4103bfef, 32'h42a334bd, 32'h40eb2475};
test_bias[2316:2316] = '{32'h426b93ee};
test_output[2316:2316] = '{32'hc58c9442};
test_input[18536:18543] = '{32'h42559d82, 32'hc2981047, 32'hc0177cb2, 32'h42167d54, 32'h414e3862, 32'hc2be4eb7, 32'h419ce753, 32'h41cbe36c};
test_weights[18536:18543] = '{32'h420bb3f9, 32'hc2821351, 32'hc1fdca6e, 32'h4291f2f1, 32'h40a57fd2, 32'hc2bc5ad3, 32'hc29bc8a9, 32'hc28f1fd9};
test_bias[2317:2317] = '{32'hc2972648};
test_output[2317:2317] = '{32'h466dfe38};
test_input[18544:18551] = '{32'hc2baf7ab, 32'hc251390b, 32'hc2410c64, 32'hc06d66cd, 32'h41aab2e2, 32'h42be63c0, 32'hc275929f, 32'hc28a10d3};
test_weights[18544:18551] = '{32'h42b78eee, 32'hc2ae1691, 32'h410cca26, 32'hc2999941, 32'h429f844d, 32'hc2a87d5e, 32'hc1a5bfa0, 32'h42831dbb};
test_bias[2318:2318] = '{32'h4276f03c};
test_output[2318:2318] = '{32'hc655b22a};
test_input[18552:18559] = '{32'hc281efe9, 32'h42a332ae, 32'h423a0411, 32'h429a42a6, 32'h42aff969, 32'hc076b006, 32'h42c7c6b5, 32'h42a1c00e};
test_weights[18552:18559] = '{32'h415fde94, 32'hc1fb52dd, 32'h425c1cc8, 32'hc2028948, 32'h423e5f58, 32'h40917eeb, 32'hc2245e4e, 32'h425a8741};
test_bias[2319:2319] = '{32'h41d6333c};
test_output[2319:2319] = '{32'h44870196};
test_input[18560:18567] = '{32'h4202dbb6, 32'h421165bf, 32'hc2b8c421, 32'h40b99bfc, 32'h421400bb, 32'hc2afa682, 32'h4134b7eb, 32'h416518b6};
test_weights[18560:18567] = '{32'h41cf089a, 32'hc2b5bda5, 32'h42970cdf, 32'hc2823ffd, 32'h42af8562, 32'hc2a7003b, 32'hc1f086f0, 32'hc087bbc6};
test_bias[2320:2320] = '{32'h42a82f5d};
test_output[2320:2320] = '{32'h43e27c50};
test_input[18568:18575] = '{32'hc2181e33, 32'h420ba3cb, 32'h422be632, 32'hc201dc73, 32'h42892ee5, 32'h41235bd9, 32'h429864c6, 32'hc2397c07};
test_weights[18568:18575] = '{32'hc20e5b4d, 32'hc2b035e1, 32'hc10a7c4e, 32'h425a580b, 32'hc28385dc, 32'h42962552, 32'h4233f717, 32'h41ecc4d4};
test_bias[2321:2321] = '{32'hc1967964};
test_output[2321:2321] = '{32'hc5ae2d18};
test_input[18576:18583] = '{32'h4247df9f, 32'h4248f81d, 32'h4250b884, 32'hc229d26a, 32'h4170b13e, 32'hc22f68f6, 32'h407980fc, 32'hc26115cb};
test_weights[18576:18583] = '{32'h4209a074, 32'h40a7be0c, 32'h42bfb657, 32'hc240cefc, 32'hc28ec389, 32'hc2ab4ad0, 32'h423de86c, 32'hc20467b3};
test_bias[2322:2322] = '{32'h42a9d855};
test_output[2322:2322] = '{32'h465855f7};
test_input[18584:18591] = '{32'hc25f97ef, 32'h42715c1d, 32'h427de29f, 32'hc217dd1c, 32'h4251ae3c, 32'h42875b55, 32'h428d109e, 32'h41c2caed};
test_weights[18584:18591] = '{32'h4150e88a, 32'hc1f751b2, 32'h42006d3a, 32'h42517832, 32'hc295415a, 32'hc21aa8e5, 32'h40d483d0, 32'hc2a5600b};
test_bias[2323:2323] = '{32'h420b63da};
test_output[2323:2323] = '{32'hc62561d6};
test_input[18592:18599] = '{32'hc29f0932, 32'hc1c54c3b, 32'h42a01730, 32'h420cd826, 32'hc131804f, 32'hc2c04aa2, 32'hc2b14445, 32'h422c33bd};
test_weights[18592:18599] = '{32'hc1e5b194, 32'hc22a6842, 32'h3fac40c4, 32'hc0ad71a3, 32'h42923884, 32'hc22251e5, 32'hc1d4ce5b, 32'hc2aacf68};
test_bias[2324:2324] = '{32'h42be6559};
test_output[2324:2324] = '{32'h459fea8e};
test_input[18600:18607] = '{32'hc0636be8, 32'hc1e26e57, 32'h4198c0e8, 32'h3f4cc8ce, 32'h42c5030b, 32'h41b12357, 32'h42be9227, 32'hbfc73680};
test_weights[18600:18607] = '{32'h426f6a74, 32'hc249c940, 32'hc25bd8ef, 32'h42b68d58, 32'h42b574a0, 32'hc2c7625d, 32'h42a5e03f, 32'hc296b671};
test_bias[2325:2325] = '{32'hc0faf51e};
test_output[2325:2325] = '{32'h466a12fb};
test_input[18608:18615] = '{32'h42c06d0e, 32'hc1e9a983, 32'h4277b45c, 32'hc203293e, 32'h42c126cc, 32'h4155a0c2, 32'hc0d20533, 32'hc2c6664c};
test_weights[18608:18615] = '{32'h4295c513, 32'hc2532085, 32'h420cc877, 32'h426d8085, 32'h3f65f227, 32'hc1ac8d3d, 32'hc18d3878, 32'hc2b3cbe3};
test_bias[2326:2326] = '{32'h4245d0f5};
test_output[2326:2326] = '{32'h468b8a32};
test_input[18616:18623] = '{32'h3e9520d3, 32'hc191a850, 32'hc280faa8, 32'hc1f14cae, 32'h41d30579, 32'hc1176522, 32'h42871ff4, 32'hbfbe905c};
test_weights[18616:18623] = '{32'hc1e6f053, 32'hc1915335, 32'h42b8312f, 32'h429afd88, 32'hc2a1514d, 32'hc2922fe2, 32'hc283efce, 32'hc233dc08};
test_bias[2327:2327] = '{32'hc2c2809c};
test_output[2327:2327] = '{32'hc658d664};
test_input[18624:18631] = '{32'hc11bf2f8, 32'hc2b0d8a1, 32'h403408c5, 32'hc1e51b1f, 32'h42295aab, 32'h42b721a4, 32'hc25b061e, 32'h41b3e56c};
test_weights[18624:18631] = '{32'hc2c2d2db, 32'h4227d714, 32'h4200e230, 32'hc2491af6, 32'hc20722b5, 32'hc1e0e325, 32'hc2362596, 32'hc0f1ac4a};
test_bias[2328:2328] = '{32'h41085173};
test_output[2328:2328] = '{32'hc5356934};
test_input[18632:18639] = '{32'h429e9f9d, 32'hc188b240, 32'h42b62513, 32'h4282622f, 32'hc2abf53f, 32'h4299f771, 32'h4134b674, 32'h42c20850};
test_weights[18632:18639] = '{32'h422d8dbf, 32'h42995217, 32'h42816a6a, 32'h4212d9d3, 32'h42c11ff0, 32'h4289feea, 32'hc2b4317a, 32'hc2bd8b82};
test_bias[2329:2329] = '{32'hc209e236};
test_output[2329:2329] = '{32'hc530369e};
test_input[18640:18647] = '{32'h427be2c1, 32'hc1ba947c, 32'hc13b9d4c, 32'h426bc043, 32'hc19ab070, 32'h41071345, 32'hc26d557c, 32'h42b0d75c};
test_weights[18640:18647] = '{32'hc0f8f140, 32'h4210ebec, 32'hc291d8f4, 32'hc2689510, 32'h42ad199c, 32'hc28e89ed, 32'hc2a83c70, 32'h42228346};
test_bias[2330:2330] = '{32'h423f4075};
test_output[2330:2330] = '{32'h451913ed};
test_input[18648:18655] = '{32'h41f7bc41, 32'hc2a4f7f3, 32'h4273f5db, 32'h4291e137, 32'h42715e95, 32'hc2220791, 32'h41ca6d9c, 32'h42608b37};
test_weights[18648:18655] = '{32'hc1e7f68d, 32'h424da24c, 32'hc2bf4df9, 32'h41c22f09, 32'hc2bcc8db, 32'h41c0f00c, 32'h4229192e, 32'hc1f67749};
test_bias[2331:2331] = '{32'h4122ee0c};
test_output[2331:2331] = '{32'hc6811808};
test_input[18656:18663] = '{32'h413b62df, 32'hc1c2d4bd, 32'hc07f54a0, 32'h41e0a716, 32'hc1b6b8de, 32'h4215e444, 32'hc153b1dd, 32'h429c6551};
test_weights[18656:18663] = '{32'h424b6c07, 32'h41fee029, 32'hc2c5b851, 32'hc12c10e0, 32'h42864e3d, 32'hc2bb0ffe, 32'h41ac3092, 32'hc2663aed};
test_bias[2332:2332] = '{32'h424682e4};
test_output[2332:2332] = '{32'hc61a1a5e};
test_input[18664:18671] = '{32'h424d6a71, 32'hc2b5186e, 32'h426ab64a, 32'h422a85f8, 32'h42bbb5b2, 32'h42045118, 32'h415e90ee, 32'h4116ea0d};
test_weights[18664:18671] = '{32'h42928926, 32'h421ea0df, 32'hc2b2ada1, 32'h422946d6, 32'hc295f401, 32'hc19df56e, 32'h42614eca, 32'h425f70a5};
test_bias[2333:2333] = '{32'h42a1e283};
test_output[2333:2333] = '{32'hc6157476};
test_input[18672:18679] = '{32'h4293473b, 32'hc2087041, 32'h429c13ab, 32'hc24a1b36, 32'hc2330ea5, 32'hc19a7eec, 32'h42ae66ec, 32'h42299d98};
test_weights[18672:18679] = '{32'hc1cdc35f, 32'h42b5baaa, 32'hc23299d8, 32'h41c0bdff, 32'hc27eddad, 32'hc1d72094, 32'h423f47aa, 32'hc22703dd};
test_bias[2334:2334] = '{32'h4293b249};
test_output[2334:2334] = '{32'hc570a538};
test_input[18680:18687] = '{32'hc21dcb63, 32'hc2ba23ea, 32'h41b6150a, 32'h41d2b8e7, 32'hc24372b7, 32'hc20a917c, 32'hbff9f689, 32'hc24b6fef};
test_weights[18680:18687] = '{32'h4250a9fd, 32'h42046b83, 32'hc17b3338, 32'h42a930d3, 32'hc2143283, 32'h421c2e18, 32'hc2bd8474, 32'hc19e1602};
test_bias[2335:2335] = '{32'hc1dd8211};
test_output[2335:2335] = '{32'hc4cdfe72};
test_input[18688:18695] = '{32'h419413b4, 32'hc2321922, 32'hc29e1b74, 32'hc28c0497, 32'hc2477686, 32'h42ba0d42, 32'hc1c0aedf, 32'h410f21f7};
test_weights[18688:18695] = '{32'h4296d90b, 32'h4156603d, 32'hc2b6254c, 32'h42b4d161, 32'h42768f6b, 32'hc1e42f7e, 32'hc2b82ae2, 32'hc2abca2f};
test_bias[2336:2336] = '{32'hc1ccb20d};
test_output[2336:2336] = '{32'hc524986e};
test_input[18696:18703] = '{32'hc2ae75fc, 32'hc0d7e545, 32'hc15dd57c, 32'h4207efc6, 32'hc1ad2894, 32'hc165c5bd, 32'h423a4d9f, 32'h4269aa9c};
test_weights[18696:18703] = '{32'hc298413b, 32'hc299f7e1, 32'h42a4e095, 32'h42465edc, 32'hc1ed05a9, 32'h42a8c042, 32'h415592da, 32'hc21f8c93};
test_bias[2337:2337] = '{32'hc28f738e};
test_output[2337:2337] = '{32'h45a73f2b};
test_input[18704:18711] = '{32'h424db154, 32'hc1287b5d, 32'hc276c64d, 32'hc20d852f, 32'hc169254e, 32'h401e06f8, 32'hc1f4c5cb, 32'h4141320c};
test_weights[18704:18711] = '{32'h4167836e, 32'hc20dab73, 32'h4218a6a5, 32'hc29fcfe6, 32'hc2c33dd9, 32'h40eec4ba, 32'h409e784f, 32'hc265b0bb};
test_bias[2338:2338] = '{32'hc2ad987e};
test_output[2338:2338] = '{32'h45032f0c};
test_input[18712:18719] = '{32'h4239a40b, 32'hc23c883e, 32'hc296ea69, 32'hc1997676, 32'hc1b2744f, 32'h40e95028, 32'h41348b23, 32'hc1a33d5c};
test_weights[18712:18719] = '{32'h41e33263, 32'hc29dc737, 32'hc09938a0, 32'hc284b4d2, 32'h41c85215, 32'h41c98c8f, 32'h429ce220, 32'hc102dd14};
test_bias[2339:2339] = '{32'h4299a6a3};
test_output[2339:2339] = '{32'h45e8037c};
test_input[18720:18727] = '{32'h41c3af15, 32'h40564c38, 32'hc268ae73, 32'hc1cefd0c, 32'hc1a342d0, 32'hc262e83e, 32'h42957f1f, 32'hc2ac4ce7};
test_weights[18720:18727] = '{32'hc1b8af9e, 32'hc1e344ee, 32'hc152df34, 32'h41c2f64c, 32'hc21be440, 32'hc160f065, 32'hc289201a, 32'hc2b07e95};
test_bias[2340:2340] = '{32'h4240a809};
test_output[2340:2340] = '{32'h4560ae24};
test_input[18728:18735] = '{32'h42b33131, 32'h428e2b5e, 32'hc2ad5db0, 32'hc22c05ad, 32'h41f9bf5c, 32'hc2c568d6, 32'hc1a25443, 32'hc29ba6a6};
test_weights[18728:18735] = '{32'h421ed643, 32'h42a5ce39, 32'h4269355b, 32'hc0ccaab2, 32'hc20feef2, 32'hc2209644, 32'hc15c403e, 32'h41e56d4f};
test_bias[2341:2341] = '{32'h42a26eaf};
test_output[2341:2341] = '{32'h45b04106};
test_input[18736:18743] = '{32'hc24dc3a5, 32'h4250ecbb, 32'hc28cfbd2, 32'hc2a3f7ea, 32'h428baa7e, 32'h42a6e76d, 32'h42a1be83, 32'h422ce391};
test_weights[18736:18743] = '{32'h41212652, 32'h3e733a1a, 32'h41e95db7, 32'hc2ba284d, 32'hc18981f5, 32'hc0acde1e, 32'hbf5e0252, 32'h42609fa7};
test_bias[2342:2342] = '{32'h41c87621};
test_output[2342:2342] = '{32'h45b53f9f};
test_input[18744:18751] = '{32'h421b8fc1, 32'hc22f53dd, 32'h42507e9d, 32'h4201682e, 32'hc2bdd2ab, 32'h413b0245, 32'h42b1a08f, 32'h422294d7};
test_weights[18744:18751] = '{32'hc2c31a32, 32'h4139aa09, 32'hc299035b, 32'h42a2f9d6, 32'h429059df, 32'hc2200e5e, 32'hc2b5628a, 32'hc294008f};
test_bias[2343:2343] = '{32'hc116c884};
test_output[2343:2343] = '{32'hc6bbd7bd};
test_input[18752:18759] = '{32'hc1ed9f37, 32'hc0833873, 32'h41c49d1e, 32'h42c6b6fb, 32'h42b5e5f8, 32'hbe3aa4c1, 32'hc1604a76, 32'h4287ff51};
test_weights[18752:18759] = '{32'hc2a9b569, 32'hc2b24223, 32'hbcb24e55, 32'h413993c8, 32'hc1c77999, 32'h42944662, 32'h42b530d4, 32'h41d61cbe};
test_bias[2344:2344] = '{32'h41f74f70};
test_output[2344:2344] = '{32'h4512156d};
test_input[18760:18767] = '{32'hbff04e9c, 32'h42149b5b, 32'h42a51243, 32'hc2a656ca, 32'h40816ba3, 32'hc17c60b0, 32'h42aa28d2, 32'h42962fd6};
test_weights[18760:18767] = '{32'hc1808c73, 32'hc2adab57, 32'hc297bdc9, 32'hc292d3fb, 32'hc13fc18d, 32'h4267b3f8, 32'hc2bc1099, 32'hc256ec0a};
test_bias[2345:2345] = '{32'hc2961080};
test_output[2345:2345] = '{32'hc68050c2};
test_input[18768:18775] = '{32'hc2a80cda, 32'h424cffb7, 32'hc29d8a01, 32'hc1e3c3c9, 32'h42178200, 32'h425f53c9, 32'h42071eaf, 32'h42844941};
test_weights[18768:18775] = '{32'hc2be51df, 32'hc24ea44e, 32'hc1c19455, 32'hc1c9e970, 32'hc282fee9, 32'hc2b206cf, 32'h42b9b671, 32'hbf319edf};
test_bias[2346:2346] = '{32'hc27e8646};
test_output[2346:2346] = '{32'h455dd5a3};
test_input[18776:18783] = '{32'hc2a70e1f, 32'hc17f2c62, 32'hc2b0c0cb, 32'hc1b0481e, 32'h429a62c3, 32'hc20e02e4, 32'hc101abc4, 32'hc0d57efd};
test_weights[18776:18783] = '{32'h4232fe2c, 32'hc1920515, 32'h41f5e7cb, 32'h424d2760, 32'hc26ce389, 32'hc277d14e, 32'h4268908a, 32'h429d3987};
test_bias[2347:2347] = '{32'h4249265a};
test_output[2347:2347] = '{32'hc625cab1};
test_input[18784:18791] = '{32'h41e32124, 32'hc2baef5a, 32'h42595c7b, 32'hc21ea1cc, 32'h422e53c4, 32'h41db1f84, 32'hc1e73742, 32'hc224403b};
test_weights[18784:18791] = '{32'hc28b22bf, 32'h425c6128, 32'h424832e3, 32'h421cf61f, 32'h427cc4a6, 32'h42031ae5, 32'h3f9703f0, 32'h4296411e};
test_bias[2348:2348] = '{32'h4112c2a1};
test_output[2348:2348] = '{32'hc5a959fa};
test_input[18792:18799] = '{32'hc23ef084, 32'hc1cf9209, 32'h42a6add7, 32'hc2a993fb, 32'hc245b851, 32'h41627436, 32'hc24ec4f8, 32'h420d65c3};
test_weights[18792:18799] = '{32'hc231911b, 32'hc0b9ee22, 32'hc160ca02, 32'h4268438e, 32'h4193ec30, 32'hc24b7ef8, 32'h420fbb09, 32'hc2bb1bcc};
test_bias[2349:2349] = '{32'hc29bd1e8};
test_output[2349:2349] = '{32'hc627338c};
test_input[18800:18807] = '{32'h4209f79b, 32'h420028a8, 32'h42b2c928, 32'hbf0dcf24, 32'hc2979b03, 32'hc1a8a908, 32'hc2144f32, 32'hc230894f};
test_weights[18800:18807] = '{32'h41c1a459, 32'h426bf186, 32'hbf8bd6a5, 32'hc29cb358, 32'h40d42e13, 32'h42512ac9, 32'h429f2b6a, 32'h41bf4b5c};
test_bias[2350:2350] = '{32'hc2a3c635};
test_output[2350:2350] = '{32'hc53ce8e0};
test_input[18808:18815] = '{32'h418b90de, 32'hc259b336, 32'hc2606e25, 32'h42c0e58a, 32'hc27706f2, 32'h423b606e, 32'hc2a0a2b7, 32'hc1f541e1};
test_weights[18808:18815] = '{32'hc29096d7, 32'hc2ae34f9, 32'h428015ea, 32'h4292352a, 32'hbf4e89e4, 32'h41ff5a8c, 32'h42343a81, 32'h42119a0d};
test_bias[2351:2351] = '{32'hc2a626f8};
test_output[2351:2351] = '{32'h4564ffbe};
test_input[18816:18823] = '{32'h42074a7b, 32'h42010155, 32'hbdd4a89d, 32'hc195d061, 32'hc230e7e4, 32'hc0cfb168, 32'h42a8f8aa, 32'h42b86261};
test_weights[18816:18823] = '{32'hc2aa7d7d, 32'hc2a2e55d, 32'h41b0c14d, 32'h424ae696, 32'hc1ad22aa, 32'hc2b55ffe, 32'hc21b677a, 32'hc1d50df5};
test_bias[2352:2352] = '{32'h42907004};
test_output[2352:2352] = '{32'hc6255781};
test_input[18824:18831] = '{32'hc1e9cfe9, 32'hc22822ef, 32'h4296f12e, 32'hc2b2a666, 32'hc244a1d6, 32'hc1fcaa11, 32'hc2a95e80, 32'h41ce8796};
test_weights[18824:18831] = '{32'hc27c8cfe, 32'h42c2ee0c, 32'h4068deec, 32'hc268430a, 32'h42ac21d8, 32'h41fa64e5, 32'h4250c54f, 32'hc2ac88a7};
test_bias[2353:2353] = '{32'hc2a2caf2};
test_output[2353:2353] = '{32'hc608880d};
test_input[18832:18839] = '{32'hc0d41205, 32'hc22523a9, 32'hc26ab9ff, 32'h42858242, 32'h4188a9e0, 32'h423745c3, 32'hc2a48ff4, 32'hc2c7ee6a};
test_weights[18832:18839] = '{32'h401f22e2, 32'h42b3149c, 32'hc286aef0, 32'h42c79b51, 32'hc20f21c0, 32'h41e25faa, 32'h411d1f47, 32'h423e768d};
test_bias[2354:2354] = '{32'hc277a25b};
test_output[2354:2354] = '{32'h44f48868};
test_input[18840:18847] = '{32'hc299fefe, 32'hc13ad240, 32'h414b0e4a, 32'hc008b6fe, 32'h4220c530, 32'hc1bc5c35, 32'hc26275dc, 32'h42770eab};
test_weights[18840:18847] = '{32'h405fba1d, 32'h428fe8ab, 32'h4284b974, 32'h428b88c3, 32'h4244ea9e, 32'hc1b041e3, 32'hc18c3b2f, 32'hc2269c2b};
test_bias[2355:2355] = '{32'hc25ac8c5};
test_output[2355:2355] = '{32'h43df2606};
test_input[18848:18855] = '{32'hc29cd435, 32'hc1cc4c87, 32'h41f59cf9, 32'hc28d4699, 32'h4120c5ba, 32'h421b5d37, 32'hc25cb372, 32'h40a9df45};
test_weights[18848:18855] = '{32'hc109cf02, 32'h42693a0f, 32'h41436b84, 32'hc2b59403, 32'h41293785, 32'h42c1489a, 32'h42c088fb, 32'h42bf9ef3};
test_bias[2356:2356] = '{32'h40bf7956};
test_output[2356:2356] = '{32'h459d6bba};
test_input[18856:18863] = '{32'hc191df40, 32'hc2820917, 32'hc2215403, 32'hbf47c0da, 32'hc26a7821, 32'h4299df50, 32'h42877a60, 32'hc2508eff};
test_weights[18856:18863] = '{32'h4112dce3, 32'h4189a096, 32'hc1d097d0, 32'h420e9d5c, 32'hc2840b82, 32'h42bd74c5, 32'hc20e77da, 32'h42964ca4};
test_bias[2357:2357] = '{32'hc1a612c8};
test_output[2357:2357] = '{32'h458e023d};
test_input[18864:18871] = '{32'hc13a1365, 32'hc299ab48, 32'hc2968f6c, 32'h4215c463, 32'hc2afe274, 32'hc28655b0, 32'h41ce0bff, 32'hc2a409ae};
test_weights[18864:18871] = '{32'hc250b17a, 32'h42c646d1, 32'hc2b69749, 32'h41dedbb5, 32'hbfaaf8a2, 32'hc1baf9b2, 32'hc2b69bcf, 32'hc298ecaa};
test_bias[2358:2358] = '{32'hc20931ea};
test_output[2358:2358] = '{32'h45ca7002};
test_input[18872:18879] = '{32'h414eba6b, 32'h41fc79f3, 32'h429bc2a9, 32'h422626c9, 32'hc2b3a1e1, 32'hc154868b, 32'hc2a68b26, 32'hc2a7cec0};
test_weights[18872:18879] = '{32'h42869ecc, 32'hc222cf5d, 32'h428542f3, 32'hc26a4b52, 32'h4136cd81, 32'hc22ec7fa, 32'hc279c508, 32'hc2700d48};
test_bias[2359:2359] = '{32'hc18bf3f2};
test_output[2359:2359] = '{32'h463d4448};
test_input[18880:18887] = '{32'h406eb036, 32'h42a4f0e8, 32'hc2a4f5ae, 32'h4191dd04, 32'hc29b7402, 32'h41d4ed75, 32'h4281bab8, 32'hc2ac0f16};
test_weights[18880:18887] = '{32'h42b954de, 32'h422f4c96, 32'hc188a98e, 32'h42a7bb04, 32'h40464e2c, 32'h4193d39d, 32'hc2ba9704, 32'h42174560};
test_bias[2360:2360] = '{32'hc0cbb5b1};
test_output[2360:2360] = '{32'hc50726da};
test_input[18888:18895] = '{32'hc0dd25a0, 32'h42237245, 32'hc2aa670c, 32'h4259ef31, 32'h4298a887, 32'hc28de56a, 32'h41ee2c1d, 32'hc2a87e7a};
test_weights[18888:18895] = '{32'hc218081f, 32'h4280ba36, 32'hc2a924a0, 32'h427888c0, 32'hc10030bc, 32'hc2be2f89, 32'hc243584c, 32'hc280e27e};
test_bias[2361:2361] = '{32'hc28c4938};
test_output[2361:2361] = '{32'h46b7c74b};
test_input[18896:18903] = '{32'hc28cf47f, 32'h42750383, 32'hc20f930c, 32'hc104f435, 32'hc1cc9eb7, 32'h4161fca4, 32'hc1f2a64f, 32'hc1903b2a};
test_weights[18896:18903] = '{32'hc2c55dc4, 32'hc1089eee, 32'hc14b3783, 32'hc2af742e, 32'h41b41aad, 32'hc2c7efcc, 32'h41031289, 32'hc22f6aa0};
test_bias[2362:2362] = '{32'hc2b04811};
test_output[2362:2362] = '{32'h45be180c};
test_input[18904:18911] = '{32'h404096f9, 32'h42afca9a, 32'h4202e1fe, 32'h420242c6, 32'h413519f6, 32'h41fe02cd, 32'h425a9a88, 32'h42aaa400};
test_weights[18904:18911] = '{32'hc28c7b42, 32'h4290ca6c, 32'hc2a7018a, 32'hc2c665e8, 32'h41e1a9fb, 32'hc27e1b16, 32'h410c8788, 32'h424f0c8f};
test_bias[2363:2363] = '{32'hc10b156b};
test_output[2363:2363] = '{32'h45533125};
test_input[18912:18919] = '{32'hc2698c37, 32'hc2b43c26, 32'h4159e394, 32'hc2bef277, 32'hc22911f4, 32'hc23de9d7, 32'hc28c0ea2, 32'hc2b6c338};
test_weights[18912:18919] = '{32'h42761508, 32'hc1e99cf7, 32'hc27fb84b, 32'hc1e03642, 32'h41c18937, 32'hc2806efe, 32'hc29a6af1, 32'h42349fe5};
test_bias[2364:2364] = '{32'hc1c8f0e0};
test_output[2364:2364] = '{32'h4580f365};
test_input[18920:18927] = '{32'h42984876, 32'h41e828b9, 32'hc20d46ac, 32'hbfefc137, 32'hc297a938, 32'hc14c7c9f, 32'hc23863a1, 32'hc040f7c1};
test_weights[18920:18927] = '{32'h4030752e, 32'hc131d6d0, 32'hc0a30486, 32'hc2c4d41b, 32'h418fe1a7, 32'h422b65f6, 32'h425ff38a, 32'hc2c3c1cc};
test_bias[2365:2365] = '{32'h40d70ba4};
test_output[2365:2365] = '{32'hc5762de9};
test_input[18928:18935] = '{32'h418912b8, 32'h411e7838, 32'hc1fd13b1, 32'h40efc281, 32'hc26eb05d, 32'hc2aecf26, 32'h426569eb, 32'h42160c54};
test_weights[18928:18935] = '{32'h423419ad, 32'hc1941b2e, 32'h4216fcc7, 32'h41eb0223, 32'hc1cc2bc5, 32'h42845d42, 32'h429911af, 32'h42b0c647};
test_bias[2366:2366] = '{32'hc23208a2};
test_output[2366:2366] = '{32'h453c4fcd};
test_input[18936:18943] = '{32'hc224c0c4, 32'h420c7065, 32'hc25b05b1, 32'h41fa2e0c, 32'hc26049d8, 32'hc21d773a, 32'h42819d9a, 32'hc1b99093};
test_weights[18936:18943] = '{32'h41973f6a, 32'h40ed5515, 32'h41c9c318, 32'h423196f6, 32'hc25c0241, 32'hc2243ed2, 32'hc24d1b80, 32'h42066abf};
test_bias[2367:2367] = '{32'hc1b18ccf};
test_output[2367:2367] = '{32'h4281c4ac};
test_input[18944:18951] = '{32'h41556e45, 32'hc0b1d9c8, 32'h4292efe6, 32'hc1ef478f, 32'hc2131f57, 32'hc2bd3aa4, 32'h42a6020f, 32'hc2c569d9};
test_weights[18944:18951] = '{32'h42a8b8ca, 32'hc291ed21, 32'h41730681, 32'h42461f1f, 32'hc179eecc, 32'h41e6849f, 32'hc2ac90b2, 32'h4143e206};
test_bias[2368:2368] = '{32'hc23784d8};
test_output[2368:2368] = '{32'hc612ea3c};
test_input[18952:18959] = '{32'h42955d28, 32'h429922cb, 32'hc2248863, 32'hc1b7fa4a, 32'hc0b4b980, 32'h4293e186, 32'h4150eaf0, 32'h4283938c};
test_weights[18952:18959] = '{32'hc2878f1c, 32'hc1bbfcd3, 32'hc194d8e1, 32'hc202417e, 32'hc1f6d5d7, 32'h42c3b23c, 32'h428b6bda, 32'h3f397616};
test_bias[2369:2369] = '{32'hc29566b4};
test_output[2369:2369] = '{32'h45381744};
test_input[18960:18967] = '{32'h423b825d, 32'h42a23923, 32'hc24d7916, 32'hc29d2696, 32'hc1e7fe8f, 32'h42835b44, 32'hc0f67d96, 32'hc2ab17b3};
test_weights[18960:18967] = '{32'h428b667b, 32'h41540e53, 32'hc2715287, 32'h41b160bd, 32'h4250ced1, 32'h422043f2, 32'hc155fa31, 32'hbff345aa};
test_bias[2370:2370] = '{32'hc250feb5};
test_output[2370:2370] = '{32'h45dbb22f};
test_input[18968:18975] = '{32'h42a2a2f7, 32'hc1870f2d, 32'hc2a4b430, 32'hc2704ef4, 32'hc07992a7, 32'hc279e0a4, 32'h42622ace, 32'hc1b2690c};
test_weights[18968:18975] = '{32'hc2446518, 32'hc0c11722, 32'hc27f6bd6, 32'hc1a853c9, 32'hc21e72d5, 32'hc247251c, 32'hc1fbae99, 32'hc2b62df8};
test_bias[2371:2371] = '{32'hc2bdb964};
test_output[2371:2371] = '{32'h45bd3208};
test_input[18976:18983] = '{32'h42900166, 32'h42721133, 32'hc183abbb, 32'h4202bd39, 32'hc2160248, 32'h41c4b626, 32'h4283870c, 32'hc1582949};
test_weights[18976:18983] = '{32'h4126aa5f, 32'h40ea7a3e, 32'h42bbea79, 32'h419e45d0, 32'hc23efe50, 32'hc2a70e60, 32'hc2a642c7, 32'hc2b56c49};
test_bias[2372:2372] = '{32'h41cd2055};
test_output[2372:2372] = '{32'hc582cad3};
test_input[18984:18991] = '{32'hc288d4a4, 32'h42937416, 32'hc2110f18, 32'hc1ab1cab, 32'h42a30f75, 32'hc27b801b, 32'h405c48d7, 32'h425f05e5};
test_weights[18984:18991] = '{32'h4171492c, 32'hc227c9e5, 32'hc24379a1, 32'h42730579, 32'hc2190a72, 32'h4255e471, 32'h42398542, 32'hc161cf65};
test_bias[2373:2373] = '{32'hc2397c50};
test_output[2373:2373] = '{32'hc628dafd};
test_input[18992:18999] = '{32'hc28e414f, 32'h414c35f3, 32'h4242cc46, 32'hc255b0cc, 32'h429aa44d, 32'hc2301ebb, 32'h4204ac79, 32'h4076f17e};
test_weights[18992:18999] = '{32'hc0f0cb32, 32'h4124cf47, 32'h41f9972d, 32'h42b18c7e, 32'h41c329a4, 32'h42a4a862, 32'hc28d62f5, 32'h42429b7d};
test_bias[2374:2374] = '{32'hc21a9905};
test_output[2374:2374] = '{32'hc5cad724};
test_input[19000:19007] = '{32'h422ab3de, 32'hc0c6ebd8, 32'hc272e018, 32'h42a4a7e3, 32'h421f74b8, 32'h3eee9243, 32'hc1f33e0e, 32'h42be4921};
test_weights[19000:19007] = '{32'h41e1093d, 32'h429c4347, 32'h42213c7e, 32'h42b54ee7, 32'h42570db3, 32'hc2bbf037, 32'h403b2629, 32'hc2b93046};
test_bias[2375:2375] = '{32'h42bca4e6};
test_output[2375:2375] = '{32'hc4738f08};
test_input[19008:19015] = '{32'hc21e9a1b, 32'hc1eafa92, 32'h416a574e, 32'h42b992e3, 32'hc235786a, 32'hc29495cc, 32'h415e3178, 32'hc2212c13};
test_weights[19008:19015] = '{32'h42b0fb93, 32'h40976bdb, 32'h409e7264, 32'h42b2e0bc, 32'hbfd1fe33, 32'h40b4d2e7, 32'hc202e1ce, 32'hc1b21495};
test_bias[2376:2376] = '{32'h420bbf69};
test_output[2376:2376] = '{32'h4597bd42};
test_input[19016:19023] = '{32'hc2a7e9d4, 32'hc2bd744b, 32'hc28c9344, 32'h4278bf05, 32'h42c582ba, 32'h428e4475, 32'h4253bbe0, 32'h42aa70af};
test_weights[19016:19023] = '{32'hc25ee699, 32'h4297618d, 32'h4286a118, 32'hc2af69a5, 32'hc0f53b4c, 32'hc29e26ea, 32'hc2758830, 32'hc2bea449};
test_bias[2377:2377] = '{32'hc1104d2d};
test_output[2377:2377] = '{32'hc6edd080};
test_input[19024:19031] = '{32'hc25f9ffd, 32'h42a66025, 32'h4291dc19, 32'hc27978bc, 32'hc298d957, 32'hc2570e2e, 32'hc28e9c24, 32'h42218551};
test_weights[19024:19031] = '{32'hc14e34c0, 32'h420d0f04, 32'hc248ca96, 32'hc09c98dc, 32'hc2858aec, 32'hc28c0723, 32'hc24d7f79, 32'h425f100e};
test_bias[2378:2378] = '{32'h4283d26e};
test_output[2378:2378] = '{32'h466caa44};
test_input[19032:19039] = '{32'h42bf9de4, 32'h42b7b399, 32'hc1d4eb70, 32'h41145572, 32'h4289202b, 32'hc2a8767e, 32'h42909a5a, 32'h428b71c4};
test_weights[19032:19039] = '{32'h41a1291e, 32'hc2a56104, 32'h42949c2f, 32'h4220a09a, 32'h42bf0b36, 32'h42b0f9de, 32'hc1d2f350, 32'hc2c1c610};
test_bias[2379:2379] = '{32'hc103ccb1};
test_output[2379:2379] = '{32'hc68398fa};
test_input[19040:19047] = '{32'hc2a59bb4, 32'h4230b2d4, 32'h422bcda1, 32'h42055f47, 32'hc2c4d4ea, 32'h41bac3d5, 32'hc261effc, 32'h42853efb};
test_weights[19040:19047] = '{32'h42676ad8, 32'hc21dd8be, 32'h427a36d3, 32'hc2c49650, 32'hc2ba2ceb, 32'h4239d3b1, 32'h41d4fb7d, 32'h426df215};
test_bias[2380:2380] = '{32'h428ca1cd};
test_output[2380:2380] = '{32'h45b098e8};
test_input[19048:19055] = '{32'h4221ffe5, 32'hc13f9636, 32'hc1c4ba94, 32'h42312819, 32'hc28a9bca, 32'hc234a7eb, 32'h426d5714, 32'hc243d872};
test_weights[19048:19055] = '{32'h42044876, 32'hc2821008, 32'hc1026a52, 32'hc106dc39, 32'hc1e3d5cf, 32'h4294b0c8, 32'hc164861b, 32'hc10211a1};
test_bias[2381:2381] = '{32'h419fec06};
test_output[2381:2381] = '{32'h4303c1e0};
test_input[19056:19063] = '{32'h42a48eee, 32'hc2626048, 32'hc0f7d6ec, 32'hc2aa81b3, 32'h42997604, 32'h42827774, 32'hc2c099c8, 32'h42c3799a};
test_weights[19056:19063] = '{32'hc2a467f7, 32'hc2b4e9c5, 32'h42af2588, 32'hc2b3d249, 32'h409dfda6, 32'hc2864910, 32'hc28c2894, 32'hc1b323a5};
test_bias[2382:2382] = '{32'h4286b90f};
test_output[2382:2382] = '{32'h45ba87c5};
test_input[19064:19071] = '{32'hc2c53f1d, 32'h42a4ed66, 32'h429275e8, 32'hc09829bc, 32'hc1e31fe3, 32'hc0631026, 32'h42c693e6, 32'h427dbbde};
test_weights[19064:19071] = '{32'hc15eee49, 32'h42bf324f, 32'hc2910750, 32'h41c2ac67, 32'h3fc43a76, 32'hc2a0c0f5, 32'h428ea6ab, 32'hc29fcb26};
test_bias[2383:2383] = '{32'hc149ab11};
test_output[2383:2383] = '{32'h45bdd26f};
test_input[19072:19079] = '{32'h42a9a662, 32'h4226e680, 32'hc2b85e43, 32'hc2808cb8, 32'hc2b28292, 32'h418e6db4, 32'h42789c54, 32'h41c2f861};
test_weights[19072:19079] = '{32'hc1cfa0d5, 32'hc1a17160, 32'h42add59b, 32'hc2b68601, 32'h4237147d, 32'h42b02bf8, 32'hc25a19d1, 32'h41679c18};
test_bias[2384:2384] = '{32'hc22301b4};
test_output[2384:2384] = '{32'hc6287f95};
test_input[19080:19087] = '{32'hc1acca52, 32'h42475c7c, 32'hc25d7183, 32'h42565142, 32'hc274f4a7, 32'h42332d75, 32'hc220ee64, 32'hc291bda6};
test_weights[19080:19087] = '{32'h429eb8d2, 32'h4287bc2b, 32'h40c50e06, 32'h41adfff2, 32'h419592fe, 32'hc1544ec3, 32'hc2bf8377, 32'h4274f5e5};
test_bias[2385:2385] = '{32'hc2a5b5f7};
test_output[2385:2385] = '{32'h4272893c};
test_input[19088:19095] = '{32'h42b37706, 32'h426f8846, 32'hc2a7ab26, 32'h42ab709e, 32'hc2280ac4, 32'h3fcf4df8, 32'hc25b0467, 32'hc1ad8edc};
test_weights[19088:19095] = '{32'hc2985e22, 32'hc1c47282, 32'hc17b90ec, 32'hc13e2619, 32'h41822ca8, 32'hc1faa17c, 32'h40888db2, 32'h4240f8ef};
test_bias[2386:2386] = '{32'hc2a6c28a};
test_output[2386:2386] = '{32'hc61de4f1};
test_input[19096:19103] = '{32'hc1d5e17c, 32'h416857aa, 32'h41a52247, 32'h42529d60, 32'hc220b1ce, 32'hc1ddfed6, 32'hc0f48c30, 32'hc286b0e2};
test_weights[19096:19103] = '{32'h4249644f, 32'h424b44fb, 32'hc229c8ff, 32'h4259aa65, 32'hc2017da5, 32'hc2a39f68, 32'h4296ddbd, 32'h42b4e357};
test_bias[2387:2387] = '{32'hc1936065};
test_output[2387:2387] = '{32'hc4d8c657};
test_input[19104:19111] = '{32'hc214a604, 32'h42267873, 32'hc1e5b797, 32'hc290b530, 32'hc2b7b24e, 32'hc1435146, 32'h422429f2, 32'hc26c8677};
test_weights[19104:19111] = '{32'h4286bfd3, 32'h425fe4b1, 32'hc27ebdaa, 32'h42a071d3, 32'hc2a7945f, 32'hc2825e58, 32'hc28c4dfe, 32'h42702d19};
test_bias[2388:2388] = '{32'h42ac9009};
test_output[2388:2388] = '{32'hc4fa34f1};
test_input[19112:19119] = '{32'hc22f7b81, 32'h411ef68a, 32'hc0e26377, 32'hc1cf04b7, 32'h4288f6bf, 32'h422a57fe, 32'hc186dc3c, 32'hc1df50d5};
test_weights[19112:19119] = '{32'h42a3bc73, 32'hbfcd8f3c, 32'hc20966c3, 32'hc2b19149, 32'h42383229, 32'hc2100d0e, 32'h424df7ca, 32'hc266bb15};
test_bias[2389:2389] = '{32'h42201e03};
test_output[2389:2389] = '{32'h44a6e06d};
test_input[19120:19127] = '{32'hc2017506, 32'hc2b845e3, 32'hc28b5e14, 32'h401df595, 32'h425e6ee9, 32'h4253a8e8, 32'h4209a7be, 32'h429b82d9};
test_weights[19120:19127] = '{32'hc23a496e, 32'hc2c6f3d0, 32'h4183bf7b, 32'h4185f4ad, 32'h41433ded, 32'h41f6add8, 32'h4137446d, 32'hc26c880c};
test_bias[2390:2390] = '{32'h402846bc};
test_output[2390:2390] = '{32'h45efdbe2};
test_input[19128:19135] = '{32'hc2c4df39, 32'h41b4db85, 32'hc2bb1a26, 32'hc2004802, 32'hc1a55198, 32'hc281b758, 32'hc2ad06cd, 32'h42117209};
test_weights[19128:19135] = '{32'hc2c15a79, 32'hc1ecadd3, 32'hc2bf8589, 32'h42a7a99e, 32'hc170cbca, 32'hc2b5e200, 32'hc29fd364, 32'h42b540d3};
test_bias[2391:2391] = '{32'hc2a51eaa};
test_output[2391:2391] = '{32'h46f5ba73};
test_input[19136:19143] = '{32'h41d37547, 32'hc29d6767, 32'h42b5230f, 32'hc20c244e, 32'hc2ae6216, 32'h42a99215, 32'h42786f06, 32'hc1aea7f5};
test_weights[19136:19143] = '{32'h428cf51a, 32'hc28eeb4e, 32'hc2b91510, 32'h42b864a8, 32'h413c3fab, 32'h418d0754, 32'hc0873e91, 32'hc131dee7};
test_bias[2392:2392] = '{32'h42323881};
test_output[2392:2392] = '{32'hc562efbf};
test_input[19144:19151] = '{32'hc1cae68c, 32'h41bad7fd, 32'h42b7f402, 32'hc28cfaee, 32'h41800ca5, 32'h4122ce3d, 32'hc2919d6f, 32'hc2accffe};
test_weights[19144:19151] = '{32'h42c7677d, 32'hc24c5d50, 32'h4198c106, 32'h422cd917, 32'h42167a7a, 32'h3f4c9fe4, 32'h41a57528, 32'hbf24dfc8};
test_bias[2393:2393] = '{32'hc2998681};
test_output[2393:2393] = '{32'hc5b94343};
test_input[19152:19159] = '{32'h42a43943, 32'h42a4ae47, 32'h42222008, 32'h4167056a, 32'hc2a85d2f, 32'hc281fa56, 32'h428df92e, 32'hc1a9c184};
test_weights[19152:19159] = '{32'hc262e198, 32'h42190f51, 32'h41cc89ce, 32'hc1694d79, 32'h3fcc6b28, 32'h427d5412, 32'h4219e380, 32'h41af08ec};
test_bias[2394:2394] = '{32'hc29e66cb};
test_output[2394:2394] = '{32'hc52b7b48};
test_input[19160:19167] = '{32'h427e7587, 32'h424a4e84, 32'hc299f674, 32'hc29fbc3c, 32'h4295d90b, 32'h41865ab3, 32'hc1b4870b, 32'hc2ac7daf};
test_weights[19160:19167] = '{32'hc181a4b0, 32'hc2aefd3d, 32'h419e9c57, 32'hc29943ba, 32'h42863cb0, 32'hc06ab2fa, 32'hc26fe55e, 32'hc2a193ae};
test_bias[2395:2395] = '{32'h41fdcab9};
test_output[2395:2395] = '{32'h4642a812};
test_input[19168:19175] = '{32'hc2a66e57, 32'hc1ae6f0c, 32'h42265986, 32'hc2acf9de, 32'h427c57ad, 32'h429f64c4, 32'hc283b652, 32'hc17aeeea};
test_weights[19168:19175] = '{32'h428561eb, 32'h429080b4, 32'hc1787f40, 32'h41444400, 32'hc2aa60cf, 32'hc198944b, 32'h427379a6, 32'h42a75cfb};
test_bias[2396:2396] = '{32'h4237c30b};
test_output[2396:2396] = '{32'hc6a41269};
test_input[19176:19183] = '{32'h42b8aed2, 32'h427c36d2, 32'hc2b14826, 32'h41d177b8, 32'hc22a96b4, 32'hc1085aa5, 32'hc202c75e, 32'hc190c0f2};
test_weights[19176:19183] = '{32'h40c49225, 32'h425711e4, 32'hc1d659dd, 32'hc26f7695, 32'hc1e08fc9, 32'h42230ea6, 32'hc2a29692, 32'hc21f3552};
test_bias[2397:2397] = '{32'h41aef1af};
test_output[2397:2397] = '{32'h460cdaa9};
test_input[19184:19191] = '{32'h42ae1f07, 32'h421ab12b, 32'h42c42385, 32'hc253e7a2, 32'hc2c6fecb, 32'hc28b0c0f, 32'h3dce4056, 32'h41e1b9f4};
test_weights[19184:19191] = '{32'h419b954c, 32'hc2c699f5, 32'h4270e6ee, 32'h410e333d, 32'h41c2b887, 32'hc24a4a7f, 32'hc231ee41, 32'h41e7a7f6};
test_bias[2398:2398] = '{32'h422c5235};
test_output[2398:2398] = '{32'h45a3b19c};
test_input[19192:19199] = '{32'hc2ba01c6, 32'hc24846a5, 32'hc230fe9c, 32'h428d4ec9, 32'hc1cfda9a, 32'h42c28ab3, 32'h42846240, 32'hc28e7836};
test_weights[19192:19199] = '{32'h42915b18, 32'h4296a11f, 32'hc080c28b, 32'hc1d03580, 32'h41a6fe2f, 32'hc2158b20, 32'hc21e2552, 32'hc280a9ad};
test_bias[2399:2399] = '{32'h42b33db8};
test_output[2399:2399] = '{32'hc65faaad};
test_input[19200:19207] = '{32'h4278b6bf, 32'hc118c094, 32'h42716f9c, 32'hc1354f32, 32'h42422edd, 32'h42620cbf, 32'hc035a831, 32'h4287c683};
test_weights[19200:19207] = '{32'hc1c15b69, 32'hc22758a3, 32'h428cd963, 32'hc2a572d8, 32'hc2b81614, 32'hc03ebb5f, 32'hc2c2386a, 32'h429e0686};
test_bias[2400:2400] = '{32'h4295505e};
test_output[2400:2400] = '{32'h45a1529b};
test_input[19208:19215] = '{32'hc274adf7, 32'hc2a026c9, 32'hc01e09e2, 32'h42bf8ca3, 32'hc2adb577, 32'hc2373451, 32'h41788d2b, 32'h42123922};
test_weights[19208:19215] = '{32'hc1a88782, 32'hc28e6d73, 32'h3fdeafb1, 32'h425ac8aa, 32'hc288a87e, 32'hc2c050d9, 32'hc15aca18, 32'h4159c215};
test_bias[2401:2401] = '{32'hc2c29481};
test_output[2401:2401] = '{32'h46b1bfdc};
test_input[19216:19223] = '{32'hbfbd32cc, 32'hc2b83c4e, 32'h429263ee, 32'h429e370f, 32'h428dd2a6, 32'hc238fae1, 32'h42c708ec, 32'hc297e244};
test_weights[19216:19223] = '{32'hc2ba211e, 32'h427b226e, 32'hc2afa583, 32'h40f00765, 32'h42547cc1, 32'h4213d086, 32'hc1e3f353, 32'hc26f9f22};
test_bias[2402:2402] = '{32'h426463b8};
test_output[2402:2402] = '{32'hc5ef1fbc};
test_input[19224:19231] = '{32'hc225a508, 32'h3fd47854, 32'hc21e7531, 32'h42540ae5, 32'hc22fdfb6, 32'h4289aa89, 32'hc286bf27, 32'hc1cfdad4};
test_weights[19224:19231] = '{32'h4204eaca, 32'h4199386b, 32'hc216ea5a, 32'hc1c9669c, 32'h4233e472, 32'h41fd732c, 32'hc2a8063a, 32'hc2b50c88};
test_bias[2403:2403] = '{32'h428e6f22};
test_output[2403:2403] = '{32'h45ddf3fa};
test_input[19232:19239] = '{32'h410dc624, 32'h40523751, 32'h42650eaf, 32'hc2a8a08d, 32'hc25f099f, 32'h4228633d, 32'h40b1e7a0, 32'h429454fc};
test_weights[19232:19239] = '{32'hc1f1858a, 32'hc204555e, 32'hc29ec0c1, 32'h4209c3b6, 32'hc179a67a, 32'hc2b2837f, 32'h41ec1135, 32'hc2b36ac1};
test_bias[2404:2404] = '{32'hc18e705a};
test_output[2404:2404] = '{32'hc68687ec};
test_input[19240:19247] = '{32'hc139e688, 32'h41bc3217, 32'h42693d26, 32'h42b5cb87, 32'hc19b4f79, 32'h42b4c211, 32'h42052300, 32'hc11783c9};
test_weights[19240:19247] = '{32'h42204f45, 32'h423a8ea4, 32'hc287339b, 32'hc03ad554, 32'h424c90d1, 32'hc18fc426, 32'h41a1152a, 32'hc28307ff};
test_bias[2405:2405] = '{32'h42afc371};
test_output[2405:2405] = '{32'hc5967163};
test_input[19248:19255] = '{32'hc299923e, 32'h41709a77, 32'hc11f47c8, 32'hc26944da, 32'hc146c4ff, 32'hc2234460, 32'hc0f82b0e, 32'h4281c22e};
test_weights[19248:19255] = '{32'h42902e3d, 32'hc2c59e26, 32'hc21056aa, 32'h42a2d6ff, 32'h42699934, 32'h425f6f03, 32'h421a72ec, 32'h41aa3b72};
test_bias[2406:2406] = '{32'hc2a6bc1d};
test_output[2406:2406] = '{32'hc651a820};
test_input[19256:19263] = '{32'h409552dd, 32'hc2c272b7, 32'hc22f3d79, 32'h422e55e2, 32'h4250594d, 32'hc1e84efc, 32'hc22d75dc, 32'h405599eb};
test_weights[19256:19263] = '{32'h42a6e33e, 32'hc24a19c1, 32'hc18cd73a, 32'h4290c19d, 32'h42c256f2, 32'hc2a211ff, 32'h42b1b59f, 32'hc28db7f1};
test_bias[2407:2407] = '{32'h4297c956};
test_output[2407:2407] = '{32'h4645505f};
test_input[19264:19271] = '{32'h424c5ea2, 32'hc28fc009, 32'h428197af, 32'hc1b44d47, 32'h420260d6, 32'h403f9346, 32'h42529e93, 32'h41eba962};
test_weights[19264:19271] = '{32'h427457c2, 32'h42bed7ce, 32'hc2169fc9, 32'hc1816396, 32'hc04771be, 32'hbfaf567c, 32'hc27161bd, 32'hc2b7ac29};
test_bias[2408:2408] = '{32'h4217f2d8};
test_output[2408:2408] = '{32'hc637cd46};
test_input[19272:19279] = '{32'hc2053fce, 32'h425a37c1, 32'h42669bb8, 32'h42adb2db, 32'hc1d8d562, 32'h4281e430, 32'hc25d62c6, 32'h41951a0b};
test_weights[19272:19279] = '{32'h4014bac4, 32'h421f2890, 32'h429ff607, 32'hc127993b, 32'hc2ababc5, 32'hc2b92266, 32'hc1bb4f89, 32'h4000bec9};
test_bias[2409:2409] = '{32'h42a38791};
test_output[2409:2409] = '{32'h455c461e};
test_input[19280:19287] = '{32'hc190d406, 32'hc1626b5c, 32'hc2491350, 32'h425a41d2, 32'h4041d4a6, 32'hc1f06fc2, 32'hc2a66a68, 32'hc2c3c955};
test_weights[19280:19287] = '{32'h4184e0b2, 32'hc2bee473, 32'hc2a292e9, 32'hc2c01f6b, 32'hc2bd0f90, 32'h41fa13d5, 32'hc28b906e, 32'hc14487a2};
test_bias[2410:2410] = '{32'hc2a4f320};
test_output[2410:2410] = '{32'h45aeda00};
test_input[19288:19295] = '{32'h4293732a, 32'h427a00dd, 32'hc29afba5, 32'hc286273a, 32'h41aec1df, 32'h41f5f458, 32'hc277e6f9, 32'h428ec964};
test_weights[19288:19295] = '{32'hc2b0a5e6, 32'hc2246077, 32'hc1c557b3, 32'hc2972325, 32'hc289f996, 32'hc2a03a52, 32'h39f0d6f0, 32'hc29ec21b};
test_bias[2411:2411] = '{32'hc2b8dc56};
test_output[2411:2411] = '{32'hc638d54a};
test_input[19296:19303] = '{32'hc2a21591, 32'h42b15fe8, 32'hc291d05d, 32'hc1c152b3, 32'hc2866c7f, 32'hc28f5ea3, 32'h423d5408, 32'hc2c2f3df};
test_weights[19296:19303] = '{32'hc198688b, 32'hc231e2e5, 32'h42c713fd, 32'hc2637ee5, 32'h42a5a410, 32'hc1a10f31, 32'h429f09ac, 32'h4244bf24};
test_bias[2412:2412] = '{32'hc20943bb};
test_output[2412:2412] = '{32'hc6527ce5};
test_input[19304:19311] = '{32'h42393fa2, 32'h421cc57a, 32'hc29ad377, 32'h424f6a54, 32'hc200a8fa, 32'h3fe2ca24, 32'h42abbd8d, 32'hc14feb2c};
test_weights[19304:19311] = '{32'h42b6940a, 32'hc2bc010a, 32'hc2b7e1af, 32'hc185d33f, 32'h40a2f015, 32'hc232fc38, 32'h42297d10, 32'h42a4dd2f};
test_bias[2413:2413] = '{32'hc25c45a0};
test_output[2413:2413] = '{32'h460d9b0e};
test_input[19312:19319] = '{32'h423fcd16, 32'hc29b1e4b, 32'hc2075aa5, 32'hc1c8e5b8, 32'hc21670cf, 32'h3fdd3a58, 32'hc1e6b0c3, 32'h418a0924};
test_weights[19312:19319] = '{32'hc22b517a, 32'h4210e5ad, 32'h4279df76, 32'h4292a0fc, 32'hc2111a16, 32'hc2a73700, 32'hc28f954e, 32'h42830409};
test_bias[2414:2414] = '{32'hc2a5641d};
test_output[2414:2414] = '{32'hc58c03f5};
test_input[19320:19327] = '{32'h41df469d, 32'h4181427a, 32'h41d85ff4, 32'h429e9665, 32'h413a2a78, 32'hc2b5d7b7, 32'hc2c620ce, 32'h42667db1};
test_weights[19320:19327] = '{32'hc2376292, 32'h3f1e2a08, 32'h42a5d5df, 32'h42431198, 32'h42ab1414, 32'hc2988367, 32'hc2aa1f4f, 32'hc29657f3};
test_bias[2415:2415] = '{32'h425fdb6f};
test_output[2415:2415] = '{32'h46842f10};
test_input[19328:19335] = '{32'hc1999533, 32'hc0603ab5, 32'h420ab3ab, 32'hc22a8dc3, 32'h42b14f1e, 32'h421e0df9, 32'hc10d475d, 32'hc21e3fd5};
test_weights[19328:19335] = '{32'hc1c69c3d, 32'h42961d5f, 32'h42920923, 32'hc1842635, 32'h429be8d1, 32'hc1ca01f6, 32'h428b6a24, 32'hc224b3cd};
test_bias[2416:2416] = '{32'h423e0d4b};
test_output[2416:2416] = '{32'h4622e0be};
test_input[19336:19343] = '{32'h41b46065, 32'hc2447444, 32'hc28efb1d, 32'h41c3988f, 32'h428e4565, 32'h429b3c99, 32'hc25e5575, 32'hc154919f};
test_weights[19336:19343] = '{32'hc24c5313, 32'hc1ff0d9f, 32'h42b91917, 32'h41fc5878, 32'h4280b639, 32'h4150316c, 32'h42a5212b, 32'hc2618a88};
test_bias[2417:2417] = '{32'h4229c4d7};
test_output[2417:2417] = '{32'hc5638c7f};
test_input[19344:19351] = '{32'hc29da2da, 32'hc2a9bc82, 32'hc0af0d4c, 32'h4261dddb, 32'hc2b8a1fa, 32'h42972b44, 32'h42bd3356, 32'hc235eefc};
test_weights[19344:19351] = '{32'h4182cfa9, 32'hc28a9e67, 32'h425ce21a, 32'hc289c2ad, 32'hc24cf1f8, 32'h42029918, 32'hc20afc03, 32'h42beae1e};
test_bias[2418:2418] = '{32'hc150961c};
test_output[2418:2418] = '{32'hc2133e19};
test_input[19352:19359] = '{32'hc2877ccb, 32'hbf07e59a, 32'h424e0b15, 32'hc268d3b2, 32'hc23157fa, 32'hc2b3d5e4, 32'h4213f398, 32'h429ac4fc};
test_weights[19352:19359] = '{32'h42b6ca50, 32'hbf38bbbf, 32'hc29f4e46, 32'hc2c65597, 32'h4279f6f2, 32'h4288c853, 32'h42722be1, 32'hbf6bc76d};
test_bias[2419:2419] = '{32'h420fc7c5};
test_output[2419:2419] = '{32'hc62f9815};
test_input[19360:19367] = '{32'hc2a317ab, 32'h42bfe267, 32'hc0ed728c, 32'h428010e1, 32'h41bfb4f3, 32'hc280b6b2, 32'hc2c79dbd, 32'hc258f9ed};
test_weights[19360:19367] = '{32'hc2b39005, 32'h414d0e6d, 32'hc2b9ea51, 32'h4094c278, 32'h42687f14, 32'hc1bd01a7, 32'hc261c179, 32'hc1e51493};
test_bias[2420:2420] = '{32'h42825bc5};
test_output[2420:2420] = '{32'h4699ee6e};
test_input[19368:19375] = '{32'h41656bb2, 32'hc2c5b0ea, 32'hc2392e3e, 32'hc29b4b4c, 32'h41c683d4, 32'h4195620c, 32'hc24c30dd, 32'hc2243e09};
test_weights[19368:19375] = '{32'h427ada7c, 32'hc29732e7, 32'hc2936a55, 32'h410f9042, 32'h420543b4, 32'h41cff050, 32'h4223b5c8, 32'hc205e2de};
test_bias[2421:2421] = '{32'hc2bb0230};
test_output[2421:2421] = '{32'h46351cb1};
test_input[19376:19383] = '{32'hc18186ed, 32'h427c8889, 32'hc283cbf6, 32'h42aadb99, 32'h42b19f92, 32'h4240986a, 32'h426703a4, 32'h40d43b81};
test_weights[19376:19383] = '{32'h42756e62, 32'hc1e27906, 32'hc1165047, 32'hc1ba0350, 32'hc2903528, 32'h42978441, 32'h41d575dd, 32'hc2b47edd};
test_bias[2422:2422] = '{32'hc200696a};
test_output[2422:2422] = '{32'hc5bb4ca2};
test_input[19384:19391] = '{32'hc12cec7f, 32'h41cbb62d, 32'h428207c2, 32'hc26b3b00, 32'hc2a5ee29, 32'hc2adffe6, 32'h42aeeca2, 32'h423a76b2};
test_weights[19384:19391] = '{32'hc2b46cc3, 32'hc00afbd6, 32'hc23a94a7, 32'h426383f7, 32'h42a9918a, 32'hc2238ce2, 32'h428ee1e6, 32'hc280a20d};
test_bias[2423:2423] = '{32'hc2a54b02};
test_output[2423:2423] = '{32'hc5b4399f};
test_input[19392:19399] = '{32'h429fc35c, 32'h41fc8534, 32'h3e8bd6b1, 32'h428950ca, 32'hc19f2c51, 32'h42920f91, 32'hc28614f4, 32'hc1851246};
test_weights[19392:19399] = '{32'hc2910508, 32'h424c008f, 32'h3f9da51d, 32'h41f2af5c, 32'h42a82fd2, 32'hc1b01992, 32'hc01b2442, 32'hc20a4e3b};
test_bias[2424:2424] = '{32'h4259eb07};
test_output[2424:2424] = '{32'hc58f5efd};
test_input[19400:19407] = '{32'hc291d27d, 32'hc1a8ba98, 32'hc20f9ef1, 32'h4194a194, 32'h41a93c38, 32'h4084f7a0, 32'h4299d112, 32'h426d80ca};
test_weights[19400:19407] = '{32'hc2b503c5, 32'hc26df859, 32'hc2ba1fc5, 32'h41ebde0f, 32'hc2a95579, 32'h422ad9f0, 32'h42099d10, 32'hc2c102cd};
test_bias[2425:2425] = '{32'h40b3332e};
test_output[2425:2425] = '{32'h45dc5619};
test_input[19408:19415] = '{32'hc299bb6e, 32'h42bc4dd8, 32'h42913d06, 32'h42a2874f, 32'hc252b9de, 32'hc2368d4c, 32'h41812b73, 32'hc028fe72};
test_weights[19408:19415] = '{32'h4257219e, 32'hc2adc802, 32'hc24ea873, 32'hc28b3365, 32'hc292c14d, 32'hc281798f, 32'hc2625c71, 32'h4112a0ca};
test_bias[2426:2426] = '{32'h42be6365};
test_output[2426:2426] = '{32'hc67605d9};
test_input[19416:19423] = '{32'hc2bdb4f2, 32'hc0a529df, 32'hc22ce956, 32'h410366bb, 32'h40bd1ee8, 32'hc0fb8a17, 32'hc23d7c42, 32'h426885a1};
test_weights[19416:19423] = '{32'h41c9daeb, 32'hc206111d, 32'h420d4ad7, 32'h42718127, 32'hc2bfbf5e, 32'h42a99a33, 32'h4280756d, 32'hc1ed79db};
test_bias[2427:2427] = '{32'h429971c5};
test_output[2427:2427] = '{32'hc60f6080};
test_input[19424:19431] = '{32'h42a5f81e, 32'h423d538c, 32'hc2956d3e, 32'h40472323, 32'hc196d96d, 32'hbdaafe98, 32'h41033efe, 32'h42abf9c5};
test_weights[19424:19431] = '{32'h41c2bb39, 32'h428641ed, 32'h40eaa54d, 32'hc18dffb7, 32'h4219079a, 32'h42c755da, 32'hc1db6af9, 32'hc050af95};
test_bias[2428:2428] = '{32'hc2b44a93};
test_output[2428:2428] = '{32'h454c4f9e};
test_input[19432:19439] = '{32'h427317be, 32'hc254bc15, 32'hc28784aa, 32'hc25d383a, 32'h429cf298, 32'hc1a5dd22, 32'hc2822680, 32'h428f3f18};
test_weights[19432:19439] = '{32'hc2465847, 32'hc1b85590, 32'h41abcb67, 32'h41dab5a4, 32'hc23a82c2, 32'hc2a6df61, 32'hc203213a, 32'hc2c044a0};
test_bias[2429:2429] = '{32'hc223d174};
test_output[2429:2429] = '{32'hc633555d};
test_input[19440:19447] = '{32'h423d23c7, 32'hc2025097, 32'hc25c099d, 32'h42c133a1, 32'h42b6f33d, 32'hc2c0fb78, 32'hc25839dd, 32'hc1a7c2d2};
test_weights[19440:19447] = '{32'h42a83cf9, 32'hc11a6dbe, 32'hc19ae051, 32'h4241fe6e, 32'hc26d31f9, 32'h42a4ad61, 32'hc2bdc508, 32'h3fde8a35};
test_bias[2430:2430] = '{32'h424ae161};
test_output[2430:2430] = '{32'h44e30196};
test_input[19448:19455] = '{32'h42c2c467, 32'h4278d4d2, 32'hc2586196, 32'h42982bb3, 32'hc245a546, 32'h428b9b24, 32'h42121113, 32'hc094d7ee};
test_weights[19448:19455] = '{32'hc2833737, 32'h427a43a5, 32'hc1282031, 32'h41d5e2c9, 32'hc0552aea, 32'hc13e3411, 32'hc2476ac6, 32'h42953299};
test_bias[2431:2431] = '{32'h41851ffc};
test_output[2431:2431] = '{32'hc52967bf};
test_input[19456:19463] = '{32'hc24f3970, 32'hc2987bf7, 32'hc2bb3495, 32'h42059243, 32'hc29b4516, 32'h4163137d, 32'hc2195640, 32'hc104d2dd};
test_weights[19456:19463] = '{32'hc2c0d448, 32'hc225e0ab, 32'hc28050c5, 32'hc22d5306, 32'hc278e5ea, 32'hc291b9c6, 32'hc2c2d28e, 32'h421bf90f};
test_bias[2432:2432] = '{32'hc26f5ed0};
test_output[2432:2432] = '{32'h469b2ca4};
test_input[19464:19471] = '{32'hc25f7017, 32'h41bc6060, 32'hc273bfc6, 32'hc26e4400, 32'h428f058f, 32'h429b1368, 32'h4249f37f, 32'h42802be2};
test_weights[19464:19471] = '{32'h4238582e, 32'hc221d95d, 32'h4205fa4c, 32'h4192c98c, 32'hc247539c, 32'hc29d4b2d, 32'h42b6c87e, 32'hc156558b};
test_bias[2433:2433] = '{32'hc245dd24};
test_output[2433:2433] = '{32'hc645221b};
test_input[19472:19479] = '{32'h428be8c5, 32'h4260485f, 32'h408d43c0, 32'h425188d6, 32'hc28c8bfc, 32'hc1b40c09, 32'h41e0ff5a, 32'h42161b6a};
test_weights[19472:19479] = '{32'hc2b5fd33, 32'h418061ca, 32'h428fcd6d, 32'hc1a7fd7e, 32'hc1cfe7f9, 32'h421d5393, 32'h42436173, 32'hc2026d6d};
test_bias[2434:2434] = '{32'h42bbbcc2};
test_output[2434:2434] = '{32'hc59e396d};
test_input[19480:19487] = '{32'h4268672c, 32'hc200b8f9, 32'h40d73e0d, 32'h41367e28, 32'h42abab50, 32'h42228aa0, 32'h423d7910, 32'hc10edc39};
test_weights[19480:19487] = '{32'hc2c3ef9c, 32'h40b80da7, 32'hc282933e, 32'h4216b974, 32'h42188615, 32'h4282eb92, 32'hc2592e9b, 32'h3f88550c};
test_bias[2435:2435] = '{32'h41b6b90c};
test_output[2435:2435] = '{32'hc51d0123};
test_input[19488:19495] = '{32'h42a51601, 32'h4037f340, 32'hc21ceed1, 32'h42a7f9b4, 32'h40b76b4d, 32'hc252fca0, 32'h41660d30, 32'h42be7714};
test_weights[19488:19495] = '{32'h4296603d, 32'hc256392a, 32'hc2a27b9d, 32'hc2389f21, 32'hc2b3d42a, 32'h4281044a, 32'h429bbe25, 32'h427ac057};
test_bias[2436:2436] = '{32'hc21466b7};
test_output[2436:2436] = '{32'h4604c6b8};
test_input[19496:19503] = '{32'hc2118806, 32'hc213b405, 32'h421b3684, 32'h42151f73, 32'h427b8605, 32'hc2527b70, 32'h40a1c562, 32'hc28e186b};
test_weights[19496:19503] = '{32'h4294dcb1, 32'h423cc4b6, 32'hc1d287bc, 32'h42b0ee01, 32'h42479509, 32'h42823b04, 32'hc26ce307, 32'hc24d9666};
test_bias[2437:2437] = '{32'h41a91ec9};
test_output[2437:2437] = '{32'h4463adca};
test_input[19504:19511] = '{32'h42993948, 32'hc2679d58, 32'hc2bac1ce, 32'hc2af06e0, 32'h42982121, 32'h42c5885a, 32'hc1d504c8, 32'h42321aae};
test_weights[19504:19511] = '{32'hc2861b9e, 32'h426263ba, 32'h428acac7, 32'hc1b90865, 32'hc258ba92, 32'hc20f0d0d, 32'hc288922d, 32'h426e4e9b};
test_bias[2438:2438] = '{32'h4278ed34};
test_output[2438:2438] = '{32'hc679da76};
test_input[19512:19519] = '{32'hc26ee7b0, 32'h40d44b90, 32'h41156a60, 32'hc2c12afe, 32'h41ebcd7f, 32'h42a315fc, 32'hc287d3fb, 32'hc27a0fed};
test_weights[19512:19519] = '{32'hc278023b, 32'h427c8859, 32'h42a9a3be, 32'h424e74f9, 32'h4226058a, 32'hc2152139, 32'hc0730e14, 32'hc26f7282};
test_bias[2439:2439] = '{32'hc1cbf2d2};
test_output[2439:2439] = '{32'h45026f6e};
test_input[19520:19527] = '{32'h4224c9dc, 32'h41ab43ed, 32'h42774019, 32'hc2191d91, 32'h42188536, 32'hc15de6f5, 32'h421441e7, 32'h42aebf57};
test_weights[19520:19527] = '{32'hc127f522, 32'h41eafd9d, 32'hc2b3a649, 32'h42c70fb9, 32'h42263c40, 32'hc22f6a1e, 32'h42c08ad7, 32'h42879e4e};
test_bias[2440:2440] = '{32'hc07d7fee};
test_output[2440:2440] = '{32'h451d4015};
test_input[19528:19535] = '{32'h421983a6, 32'h4249ad07, 32'hc15ed388, 32'h419d0c89, 32'h40521994, 32'hc299cb0c, 32'hc27ddb4e, 32'hc297a2c8};
test_weights[19528:19535] = '{32'h42c0898e, 32'h42473fd4, 32'hc2157411, 32'h42a5cffb, 32'hc2470bf2, 32'hc239bfea, 32'hc1dadb5b, 32'h411cf65f};
test_bias[2441:2441] = '{32'h428b674d};
test_output[2441:2441] = '{32'h46485ea3};
test_input[19536:19543] = '{32'hc1f893c8, 32'hc20a1e1e, 32'hc278ed91, 32'hc295f740, 32'hc2a1498d, 32'h42612eb0, 32'h425ddee6, 32'hc259bae9};
test_weights[19536:19543] = '{32'h41ddb74a, 32'hc25bdc42, 32'h428f1a0c, 32'h41dea166, 32'hc1cff6df, 32'hc170f271, 32'hc28e0316, 32'hc1951f25};
test_bias[2442:2442] = '{32'hc272d0d8};
test_output[2442:2442] = '{32'hc5e23567};
test_input[19544:19551] = '{32'hc2879f21, 32'hc0853b1e, 32'h42617aeb, 32'h42946e59, 32'h428e0b4b, 32'hc20c4751, 32'h4271ec28, 32'hc213178f};
test_weights[19544:19551] = '{32'hc0b1d8df, 32'h419b0b4c, 32'h4012e494, 32'h42c197b4, 32'hc1f22ba1, 32'h4205da2e, 32'hc281e72e, 32'h428032db};
test_bias[2443:2443] = '{32'hc1c4f67c};
test_output[2443:2443] = '{32'hc4fd0571};
test_input[19552:19559] = '{32'h42415b9f, 32'h42a2b503, 32'h42a311da, 32'h42975d80, 32'hc158103d, 32'h3e0b4a0e, 32'h41aa027f, 32'hc2277fd3};
test_weights[19552:19559] = '{32'h420a3872, 32'hc2c6b79d, 32'hc17e955b, 32'hc275a511, 32'hc1a5a946, 32'hbeb19931, 32'h410afdcd, 32'hc25c7353};
test_bias[2444:2444] = '{32'h421d8c28};
test_output[2444:2444] = '{32'hc61529ee};
test_input[19560:19567] = '{32'hc0d7ee87, 32'h42b1d649, 32'hc2aa8067, 32'hc2736357, 32'hc2bbdfb4, 32'hc2aaec42, 32'h41d81e5f, 32'hc1238761};
test_weights[19560:19567] = '{32'h41dcb571, 32'hc28f510e, 32'hc24fef72, 32'h42b99a36, 32'h41b729b4, 32'h4294af7c, 32'hc184f941, 32'hc25e7d94};
test_bias[2445:2445] = '{32'h41f93777};
test_output[2445:2445] = '{32'hc67bf9e4};
test_input[19568:19575] = '{32'hc2037c08, 32'hc2bd7d3c, 32'hc2c3eae7, 32'hc2a49ed9, 32'hc283d10c, 32'h42723714, 32'hc092e01f, 32'h41d5b786};
test_weights[19568:19575] = '{32'hc23159e9, 32'hc1cb725f, 32'hc2873eb9, 32'hc21fd12f, 32'h41f0ce7e, 32'h424e3261, 32'hc2c01ca4, 32'h429cb25f};
test_bias[2446:2446] = '{32'h429a5718};
test_output[2446:2446] = '{32'h4688f0e1};
test_input[19576:19583] = '{32'hc10bd0c2, 32'h420278fb, 32'hc21689a4, 32'h427ef146, 32'h41a3d719, 32'hc282c235, 32'hc1edffb7, 32'hc18f88ec};
test_weights[19576:19583] = '{32'h42b6c3da, 32'hc106c7c9, 32'h429f117f, 32'h42b4440a, 32'h4255f875, 32'hc27e5056, 32'hc2af3b73, 32'hc2b6ac14};
test_bias[2447:2447] = '{32'hc2b25ab2};
test_output[2447:2447] = '{32'h462d3a12};
test_input[19584:19591] = '{32'hc2a1c7ae, 32'hc29a1ac9, 32'hc1d14925, 32'h41fdeef3, 32'hc1f0417d, 32'hc2a9360c, 32'hc2b0de1b, 32'hc256a079};
test_weights[19584:19591] = '{32'h41e5ccde, 32'hc2260f75, 32'h413c67a5, 32'h42c60923, 32'h428ee6d8, 32'h425629b0, 32'hc27c132f, 32'hc2967bb9};
test_bias[2448:2448] = '{32'h42b1bc5b};
test_output[2448:2448] = '{32'h45d26d07};
test_input[19592:19599] = '{32'hc2904eda, 32'hc2b57c43, 32'hc1c8719e, 32'hc2324394, 32'h4246a271, 32'hc0c715a3, 32'h420b0306, 32'hc1c2bef0};
test_weights[19592:19599] = '{32'hc2024bd3, 32'h41b7fc34, 32'hc268183a, 32'hc2514c4f, 32'h41a08138, 32'hc17e9418, 32'h424bb9e8, 32'h428b2b32};
test_bias[2449:2449] = '{32'h40517e89};
test_output[2449:2449] = '{32'h45a33e91};
test_input[19600:19607] = '{32'hc1b95275, 32'hc16f2fee, 32'h410a5349, 32'hc21940a7, 32'hc1994cab, 32'h426957cf, 32'hc1ccdb83, 32'hc23e5a15};
test_weights[19600:19607] = '{32'hc296bfe8, 32'hc275cbea, 32'h42b96ada, 32'h419a872c, 32'hc23abf2c, 32'h413f7909, 32'h41d53aaa, 32'hc158d31c};
test_bias[2450:2450] = '{32'hc11f5d54};
test_output[2450:2450] = '{32'h45857a36};
test_input[19608:19615] = '{32'h41fe385c, 32'hc298c7a5, 32'hc2009e06, 32'h428f170e, 32'hc2b34e76, 32'h42165ade, 32'hc2566b64, 32'hc297748d};
test_weights[19608:19615] = '{32'hc28bb3d3, 32'hc2b5132b, 32'hc2c1a6ed, 32'h3f6a5390, 32'hc2beab29, 32'h424cf914, 32'h42a85893, 32'hc1434eec};
test_bias[2451:2451] = '{32'h429d0de5};
test_output[2451:2451] = '{32'h4667dd61};
test_input[19616:19623] = '{32'h41be5726, 32'h424b12fa, 32'hc11669f9, 32'hbf8b806b, 32'hc259aebd, 32'hc11f0f05, 32'hc2bbeb78, 32'hc287f178};
test_weights[19616:19623] = '{32'hc2af4298, 32'hc28741e1, 32'hc2bb68eb, 32'hc2a1a779, 32'hc24c8406, 32'h42a056a0, 32'h41122b18, 32'hc2ae6ea5};
test_bias[2452:2452] = '{32'hc2bd5968};
test_output[2452:2452] = '{32'h4516b502};
test_input[19624:19631] = '{32'h411c0f58, 32'h410927eb, 32'hc29b7439, 32'h412cc4d6, 32'h4286363e, 32'hc1e24fb2, 32'h4245eef9, 32'hc14b1ecd};
test_weights[19624:19631] = '{32'hc15df86d, 32'h4044e4b9, 32'hc2ab2e1d, 32'hc0d9f989, 32'hc19c315b, 32'hc2c52678, 32'hc2b9b812, 32'h4237c71b};
test_bias[2453:2453] = '{32'hc2c14ca7};
test_output[2453:2453] = '{32'h45271a56};
test_input[19632:19639] = '{32'hc1486f16, 32'hc20c859b, 32'hc1696a89, 32'h42574919, 32'h418c6ac0, 32'h42b325a7, 32'h424d6a5d, 32'hc2837c80};
test_weights[19632:19639] = '{32'hc2a3a831, 32'h4294ff22, 32'hc24d2678, 32'h4268a7b9, 32'h41b92af0, 32'hc1f12662, 32'hc1549827, 32'h4124ab7a};
test_bias[2454:2454] = '{32'h422ce145};
test_output[2454:2454] = '{32'hc4a55f98};
test_input[19640:19647] = '{32'hc16b5e30, 32'hc0ccf1d9, 32'h42c53d6e, 32'h40d2289b, 32'hc2b3052e, 32'h42acc002, 32'hc2788229, 32'hc23049ae};
test_weights[19640:19647] = '{32'hc29d8cc1, 32'h4296c5f6, 32'hc2bc34fc, 32'hc0372015, 32'hbe093501, 32'hc23aa37f, 32'hc283841e, 32'hc1e61a2b};
test_bias[2455:2455] = '{32'h41ba9a15};
test_output[2455:2455] = '{32'hc5e3098e};
test_input[19648:19655] = '{32'hc0e6c6a0, 32'hc2acaaa6, 32'hc25591b4, 32'hc24f9cd5, 32'h428c432d, 32'h416b250b, 32'hc23d4e27, 32'h427de07c};
test_weights[19648:19655] = '{32'h4269fe4c, 32'h42571190, 32'h42873d18, 32'h42c6b6b2, 32'h4289dcc0, 32'h421d68b8, 32'hc296bbbb, 32'hc284f920};
test_bias[2456:2456] = '{32'h41cb76f0};
test_output[2456:2456] = '{32'hc60d5850};
test_input[19656:19663] = '{32'h429e6361, 32'hc2b0f945, 32'hc0c2c57b, 32'h422b38b6, 32'h428483ca, 32'hc2171eec, 32'h42302424, 32'hc27bb840};
test_weights[19656:19663] = '{32'h428744f4, 32'h42bf115c, 32'h41f005e6, 32'hc23ed424, 32'hc22d205b, 32'h42adb986, 32'hc1b07651, 32'hc1b17c7b};
test_bias[2457:2457] = '{32'h42bed9a1};
test_output[2457:2457] = '{32'hc62b1c77};
test_input[19664:19671] = '{32'hc27ea85f, 32'hc1e02071, 32'h411e53ce, 32'hc2a43da6, 32'h3feab359, 32'hc2885f5b, 32'hc2c66df9, 32'h4123e7f7};
test_weights[19664:19671] = '{32'h42b989e1, 32'h4244297d, 32'h4288b886, 32'hc233e512, 32'h424b07cf, 32'h4281a142, 32'hc20f3ebb, 32'hc24108ae};
test_bias[2458:2458] = '{32'h42900345};
test_output[2458:2458] = '{32'hc5805091};
test_input[19672:19679] = '{32'h42c1d95f, 32'hc1f09bce, 32'h429e31be, 32'hc2ab166a, 32'h4245844c, 32'h4286406e, 32'h427fafeb, 32'hc2bccf0d};
test_weights[19672:19679] = '{32'h4286402a, 32'hc1b1263b, 32'h42016f90, 32'hc036e573, 32'hc2b68e23, 32'h42a07d52, 32'h4169241e, 32'h4291ae29};
test_bias[2459:2459] = '{32'hc2058825};
test_output[2459:2459] = '{32'h4598678c};
test_input[19680:19687] = '{32'hc217e883, 32'h410b9c4f, 32'hc0e150b9, 32'h41de5224, 32'h413616ee, 32'hc217972b, 32'hc1e071c7, 32'hc1b7d034};
test_weights[19680:19687] = '{32'h4074858a, 32'h4285ab94, 32'hc204bdbf, 32'h427d5d41, 32'h4232e725, 32'hc21cec9a, 32'hc297b1b8, 32'h42814d2e};
test_bias[2460:2460] = '{32'h423283ab};
test_output[2460:2460] = '{32'h459fd6fa};
test_input[19688:19695] = '{32'hc1afa500, 32'hc2863242, 32'h42aaeabb, 32'hc1a565ff, 32'hc18fc115, 32'h4275d8fb, 32'h4163c79a, 32'hc21362ef};
test_weights[19688:19695] = '{32'h4223d628, 32'h42c4f0ee, 32'hc21847f0, 32'h427f3c12, 32'hbfcd514f, 32'hc12b4122, 32'h41dbc7e4, 32'hc2b06b54};
test_bias[2461:2461] = '{32'hc230e13b};
test_output[2461:2461] = '{32'hc60e5c30};
test_input[19696:19703] = '{32'h4286259a, 32'hc2acc884, 32'hc19f4470, 32'h425a2d0f, 32'h427b58f7, 32'hc204d8ff, 32'h41e8d139, 32'hc2b30a68};
test_weights[19696:19703] = '{32'hc2a949cd, 32'hc2b7ede8, 32'h41e1fb88, 32'h40ceaa67, 32'h428988e5, 32'hc09b7729, 32'h421ef8b6, 32'hc1f92bb4};
test_bias[2462:2462] = '{32'h4290be90};
test_output[2462:2462] = '{32'h4624f4ba};
test_input[19704:19711] = '{32'h429cd539, 32'h42173de8, 32'h4263e44d, 32'h4245491a, 32'hc2925a17, 32'hc0c31f20, 32'hc29564c9, 32'h41a382a6};
test_weights[19704:19711] = '{32'h4115245f, 32'hc22d7106, 32'hc28a3d5a, 32'hc1147937, 32'hbf9e3d67, 32'h41ee34ab, 32'h4219c9aa, 32'hc2c35cac};
test_bias[2463:2463] = '{32'hc2a3ac1d};
test_output[2463:2463] = '{32'hc621a5ca};
test_input[19712:19719] = '{32'h4280644f, 32'h41467dec, 32'h42b94273, 32'hc292e6be, 32'hc1fe5c95, 32'hc1837be8, 32'h42872373, 32'hc16feba6};
test_weights[19712:19719] = '{32'hc24f056a, 32'hc121cae6, 32'hc1780f7b, 32'h42accbbb, 32'hc2c184af, 32'hc296580f, 32'h42190dd2, 32'h40e7f145};
test_bias[2464:2464] = '{32'h4219437c};
test_output[2464:2464] = '{32'hc58997ee};
test_input[19720:19727] = '{32'hc2c113ee, 32'h41aa21fa, 32'hc2c5da3e, 32'hc1365f53, 32'h421f6cdb, 32'hc1bf9185, 32'h423eabc4, 32'h4296d55f};
test_weights[19720:19727] = '{32'h4182fa18, 32'h42bb033d, 32'h4281b0eb, 32'hc2ba30a1, 32'hc2ae5e97, 32'hc29c9e33, 32'hc200977d, 32'hc1d61a21};
test_bias[2465:2465] = '{32'hc124da26};
test_output[2465:2465] = '{32'hc61dea2d};
test_input[19728:19735] = '{32'hc29c562b, 32'hc286c23e, 32'hc260d73a, 32'h41d79b2d, 32'hc1a5d2a3, 32'h424726be, 32'hc12bb5cf, 32'h3f8ca67c};
test_weights[19728:19735] = '{32'hc22e2c19, 32'h41cf6271, 32'hc236b95c, 32'hc2ad2533, 32'h41dd4746, 32'hc2477d8b, 32'h4215500b, 32'hc258df3d};
test_bias[2466:2466] = '{32'h42972aeb};
test_output[2466:2466] = '{32'hc4c1ad9f};
test_input[19736:19743] = '{32'h4072871a, 32'hc1e98544, 32'h4275fda6, 32'hc2bef00b, 32'h4134ab83, 32'hc2490dde, 32'h425a2d3d, 32'hc24b74c7};
test_weights[19736:19743] = '{32'hc23c1ae3, 32'hc290e505, 32'hc222e33b, 32'h42240e78, 32'hc2b6edf3, 32'h42c0124c, 32'hc22858d3, 32'h42aa3937};
test_bias[2467:2467] = '{32'hc2084417};
test_output[2467:2467] = '{32'hc684d40c};
test_input[19744:19751] = '{32'h41c2171d, 32'h401635f8, 32'hc1f7e7b5, 32'hc23c41ec, 32'hc2b6b5ea, 32'h41bcdf17, 32'hc2260d17, 32'hc29165a6};
test_weights[19744:19751] = '{32'h42b290df, 32'hc21a9aba, 32'hc29824a0, 32'hc291a553, 32'hc180169f, 32'h423ddb0c, 32'hc2664d83, 32'h42a67630};
test_bias[2468:2468] = '{32'hc20aec8e};
test_output[2468:2468] = '{32'h45d2dfe3};
test_input[19752:19759] = '{32'hc29ae8d8, 32'hc23f6b30, 32'h410f94c7, 32'h41fd0d8a, 32'hc1f0d742, 32'hc00bd539, 32'h41f9025b, 32'hc230c73d};
test_weights[19752:19759] = '{32'h428551d9, 32'hc2a9f68b, 32'hc0292c0a, 32'h42b68863, 32'hc18e49a6, 32'hc1d61653, 32'h426863fb, 32'h41b31135};
test_bias[2469:2469] = '{32'h4188b5bf};
test_output[2469:2469] = '{32'h4547cf56};
test_input[19760:19767] = '{32'h42436ec6, 32'h42535963, 32'h42445039, 32'hc2833acd, 32'h41ff6118, 32'h42b38bf1, 32'h42637c3e, 32'h41fc06e3};
test_weights[19760:19767] = '{32'hc277b056, 32'hc22a3908, 32'h427292d3, 32'hc23672bf, 32'hc289a36b, 32'hc116d91c, 32'hc1ebd778, 32'hc28570df};
test_bias[2470:2470] = '{32'hc21840ec};
test_output[2470:2470] = '{32'hc5c0a52d};
test_input[19768:19775] = '{32'h42bc4878, 32'h418e020d, 32'hc25d541d, 32'h41ad1c0b, 32'h41944ee1, 32'hc1c66674, 32'hc12199df, 32'hc2a065b2};
test_weights[19768:19775] = '{32'h4160027c, 32'h42b892ae, 32'hc239e59d, 32'h428ba486, 32'hc0ac428f, 32'h421ad81e, 32'h42c353e8, 32'hc286fa01};
test_bias[2471:2471] = '{32'h419ecc35};
test_output[2471:2471] = '{32'h4622e29d};
test_input[19776:19783] = '{32'h42073946, 32'hc2bb3008, 32'h42b47708, 32'h41f661a9, 32'hc18c1983, 32'h42671b9e, 32'hc21afdb9, 32'hc24900db};
test_weights[19776:19783] = '{32'h42672cc2, 32'hc218613d, 32'h418b4da9, 32'h42c29527, 32'h42725a49, 32'h42a9eac2, 32'h42508a94, 32'h42837eef};
test_bias[2472:2472] = '{32'hc1880695};
test_output[2472:2472] = '{32'h46064570};
test_input[19784:19791] = '{32'hc2bdf537, 32'hc246096d, 32'hc29b5a91, 32'hc281e153, 32'h4299f51f, 32'hc25e6521, 32'hc259d7bf, 32'h420f70bb};
test_weights[19784:19791] = '{32'hc1f0da0d, 32'h428e047a, 32'h421ec030, 32'h4189c3c9, 32'h42b573d2, 32'hc0973617, 32'hc18bce5d, 32'hc1bc1ec0};
test_bias[2473:2473] = '{32'h4289673a};
test_output[2473:2473] = '{32'h45206adc};
test_input[19792:19799] = '{32'h42a080ea, 32'h42a0e73e, 32'h4236d28e, 32'h419c0926, 32'hc2a853b1, 32'h41c8811b, 32'h41082651, 32'hc2b2ec74};
test_weights[19792:19799] = '{32'hc23e299b, 32'h426e6cb6, 32'h41f038c0, 32'hc293a694, 32'hc09c8f99, 32'hbfd0d379, 32'h42adfe97, 32'h41e847d9};
test_bias[2474:2474] = '{32'hc1d983a7};
test_output[2474:2474] = '{32'hc41635f2};
test_input[19800:19807] = '{32'hc212d414, 32'h41ff97c5, 32'hc23d1630, 32'hbf691095, 32'hc2befa25, 32'hc2b8ab5f, 32'hc207eace, 32'hc297a0f7};
test_weights[19800:19807] = '{32'hc2182f97, 32'h41a36415, 32'hc2a1625c, 32'h42a62d32, 32'hc2805aca, 32'h429ec4a2, 32'h4226e64e, 32'h42658362};
test_bias[2475:2475] = '{32'h419ddb9e};
test_output[2475:2475] = '{32'hc4913e55};
test_input[19808:19815] = '{32'h41076c33, 32'hc2a87955, 32'h41c6e013, 32'hc2a513b5, 32'hc2a252e9, 32'h417e53b5, 32'h423efc87, 32'hc10fa6cb};
test_weights[19808:19815] = '{32'h42c22147, 32'hc0e97dd3, 32'h42af1abd, 32'h427b7cd3, 32'h42a33aad, 32'hc291f7a9, 32'hc2c1383e, 32'h41e2725b};
test_bias[2476:2476] = '{32'hc1c2d3fe};
test_output[2476:2476] = '{32'hc65eb033};
test_input[19816:19823] = '{32'hc147624c, 32'h4284b35c, 32'h4220b091, 32'hc25cc0e0, 32'h42829445, 32'h42895450, 32'hbfa8f2bc, 32'hc2ace3ea};
test_weights[19816:19823] = '{32'hc11d26cc, 32'h414a7f40, 32'hc2b02173, 32'hc1ae879e, 32'h42122ef3, 32'hc1e8d172, 32'h4195ca10, 32'hc268a73c};
test_bias[2477:2477] = '{32'h42c672fb};
test_output[2477:2477] = '{32'h4580b45f};
test_input[19824:19831] = '{32'hc2521a1e, 32'hc29fa7ca, 32'h41873008, 32'hc297069b, 32'h4230961e, 32'h3ef278e9, 32'h42038b0d, 32'hc247d688};
test_weights[19824:19831] = '{32'h413f1dc2, 32'hc21b2c4f, 32'h428614e0, 32'hc0faf1ec, 32'h422e96bb, 32'h414fa38c, 32'h4299c022, 32'h429eecd4};
test_bias[2478:2478] = '{32'h428b2eb1};
test_output[2478:2478] = '{32'h459499eb};
test_input[19832:19839] = '{32'hc2b41905, 32'h42650dcc, 32'hc13dec27, 32'h421a5c50, 32'hc1ce8c55, 32'hc20bf9f4, 32'h4269d2e1, 32'h41630230};
test_weights[19832:19839] = '{32'h42c5d36d, 32'h421f7613, 32'h41e9e8dc, 32'h4250e72a, 32'h4216c72b, 32'h425e4f3e, 32'hc1f09116, 32'hc218ca2d};
test_bias[2479:2479] = '{32'h410de897};
test_output[2479:2479] = '{32'hc61ed355};
test_input[19840:19847] = '{32'hbfc00c8d, 32'hc1f5afd2, 32'hc2810a9b, 32'h429a6cfc, 32'hbfcca954, 32'hc18e7e52, 32'h428f2f7a, 32'h418db6a6};
test_weights[19840:19847] = '{32'h42060938, 32'hc21d8424, 32'hc26fa3c1, 32'h3e4facb9, 32'h42b9d619, 32'h42c26fbf, 32'h42a9c2cf, 32'h40c03cc3};
test_bias[2480:2480] = '{32'hc18f67ed};
test_output[2480:2480] = '{32'h4611b538};
test_input[19848:19855] = '{32'h42bc5ee6, 32'h427cab3d, 32'hc1a61c48, 32'hbeafb356, 32'hc12120d0, 32'h4152de4f, 32'hc2aa1213, 32'h415dde1c};
test_weights[19848:19855] = '{32'hc219fc72, 32'hc2213933, 32'h4289e66a, 32'hc1df4925, 32'hc2acb1cf, 32'h41b49c16, 32'hc1936209, 32'h41c5aeb3};
test_bias[2481:2481] = '{32'hc29b73a8};
test_output[2481:2481] = '{32'hc58f9a4b};
test_input[19856:19863] = '{32'hc2788185, 32'h42b83e8d, 32'h42bec68e, 32'h42b88d9d, 32'h42169129, 32'h42b1aaa0, 32'h419c3344, 32'h41719be2};
test_weights[19856:19863] = '{32'h4284362d, 32'hc07fdbd6, 32'h41f477b6, 32'hc21a612c, 32'h42c0d593, 32'hc2998928, 32'hc18df74f, 32'hc13e127f};
test_bias[2482:2482] = '{32'hc18a8cb3};
test_output[2482:2482] = '{32'hc60a5c87};
test_input[19864:19871] = '{32'hc28b8fd0, 32'h41c10c4e, 32'h41b1086b, 32'hc28dbedc, 32'hc2ab7583, 32'h429aad0d, 32'hc1c0bea8, 32'hc291138b};
test_weights[19864:19871] = '{32'hc2a52a59, 32'hc1289362, 32'h42c2c757, 32'hc1101870, 32'h41a306aa, 32'hc287f9f8, 32'hc18a0403, 32'h42495fac};
test_bias[2483:2483] = '{32'hc27bef2d};
test_output[2483:2483] = '{32'hc4fa4bf3};
test_input[19872:19879] = '{32'hc271e6d7, 32'hc225785f, 32'h42a24523, 32'hc29666f6, 32'h4285eb02, 32'h42aa18c8, 32'h4292c14b, 32'h421200b9};
test_weights[19872:19879] = '{32'hc2190d7d, 32'hc18d0339, 32'hc2086694, 32'hc2aa1399, 32'h422eeaf8, 32'hc2a914d5, 32'hc1a15253, 32'h40847751};
test_bias[2484:2484] = '{32'hc285e2e0};
test_output[2484:2484] = '{32'h447d7a96};
test_input[19880:19887] = '{32'h42b02d3c, 32'hc229e5f1, 32'hc1a358e2, 32'hc1fb9f68, 32'hc29ca81c, 32'h41e67ea6, 32'hc14ca4e8, 32'h41b7760a};
test_weights[19880:19887] = '{32'h412a4f5a, 32'hc28613c9, 32'hc1c6a1e5, 32'hc2c1d747, 32'h41ffd19a, 32'h4251bf96, 32'h4235759e, 32'hc101fa90};
test_bias[2485:2485] = '{32'hc2b210c4};
test_output[2485:2485] = '{32'h45ab97f1};
test_input[19888:19895] = '{32'h4225bc2e, 32'h426656b9, 32'hc0686a5d, 32'hc294d64b, 32'hc25d4f2b, 32'h42c14049, 32'hc2a8842f, 32'hc1cebf6e};
test_weights[19888:19895] = '{32'h4214b580, 32'h3d850986, 32'h42c17cd2, 32'hc18a17c4, 32'h422809ab, 32'h42455d52, 32'h42a9a77a, 32'h42bebcfa};
test_bias[2486:2486] = '{32'h4189aa6a};
test_output[2486:2486] = '{32'hc59210ca};
test_input[19896:19903] = '{32'hc1b12b69, 32'hc2653a9c, 32'h4209c882, 32'h42c34f1a, 32'h411f731c, 32'h429ef92c, 32'hc2124805, 32'h429cfdb9};
test_weights[19896:19903] = '{32'h4211af45, 32'hc27ef3bf, 32'hc24aeeb5, 32'h41c002c3, 32'h41f9d091, 32'hc225c198, 32'hc2bfea59, 32'h42ad4565};
test_bias[2487:2487] = '{32'hc2adec10};
test_output[2487:2487] = '{32'h4626e9ca};
test_input[19904:19911] = '{32'hc283fe3a, 32'h41eb7b6b, 32'hc13e9800, 32'hc28e84b3, 32'hc200c00a, 32'h42828d49, 32'hc170bc52, 32'hc2a0abac};
test_weights[19904:19911] = '{32'h423d039d, 32'hc2ac8d9e, 32'h4218f770, 32'h429f2479, 32'hc243400e, 32'h42a219f6, 32'h42248bdd, 32'h4205794f};
test_bias[2488:2488] = '{32'h408c7876};
test_output[2488:2488] = '{32'hc600650c};
test_input[19912:19919] = '{32'hc280f9c0, 32'h418c8aba, 32'hc206299f, 32'h42b1e4e8, 32'hc23322ca, 32'hc23d1d10, 32'hc1bc60cd, 32'hc28d6dda};
test_weights[19912:19919] = '{32'hc25360e3, 32'hc27c9a33, 32'h42772a02, 32'h42b5cd77, 32'h423bb434, 32'h42976304, 32'hc1d66e0c, 32'hc2b641b9};
test_bias[2489:2489] = '{32'h42b79740};
test_output[2489:2489] = '{32'h461918b2};
test_input[19920:19927] = '{32'hc2920011, 32'hc1e73e19, 32'hc239c390, 32'hc287bdb4, 32'hc1f10981, 32'hc2419d01, 32'h421e13b0, 32'hc254ec11};
test_weights[19920:19927] = '{32'hc2a6bf32, 32'h427680c9, 32'hc29d5fc7, 32'h428a2739, 32'h429b2e32, 32'hc141a9ad, 32'h42949617, 32'h42ad21c8};
test_bias[2490:2490] = '{32'h40814969};
test_output[2490:2490] = '{32'hc314cd9b};
test_input[19928:19935] = '{32'h428d729a, 32'hc251065a, 32'hc124f68a, 32'h42814ace, 32'hc24ef069, 32'h42bc7ab5, 32'hc28f3629, 32'hc1ae022f};
test_weights[19928:19935] = '{32'h428b1b7f, 32'h40e9026b, 32'h42ab99f3, 32'h424bf6f0, 32'hc274f420, 32'hc2a54d9c, 32'hc058e6be, 32'hc1a7ef41};
test_bias[2491:2491] = '{32'h42a9d2e8};
test_output[2491:2491] = '{32'h45429a36};
test_input[19936:19943] = '{32'hc28729c2, 32'hc2a6424f, 32'hc28bebe3, 32'h429a9fb5, 32'h42195498, 32'hc2c685c0, 32'h4287ec05, 32'hc11841d3};
test_weights[19936:19943] = '{32'hc106774e, 32'hbf48efeb, 32'h428e50b3, 32'h42ab79ea, 32'h4258220b, 32'hc2c6b61f, 32'hc224b069, 32'h42b5ec92};
test_bias[2492:2492] = '{32'hc28476fb};
test_output[2492:2492] = '{32'h4623dc13};
test_input[19944:19951] = '{32'h4116459f, 32'hc176d0fc, 32'h42a7c5d6, 32'h42381398, 32'h42900dfe, 32'hc201bb1c, 32'hc0f91863, 32'hc209e5fd};
test_weights[19944:19951] = '{32'hc2aabdcb, 32'h42a5291f, 32'hc0b76f27, 32'h420fd16c, 32'h429c3229, 32'h42462c6f, 32'hc29534b8, 32'h42013eb6};
test_bias[2493:2493] = '{32'h4253b2e4};
test_output[2493:2493] = '{32'h4524c23d};
test_input[19952:19959] = '{32'h41a3768e, 32'hc198bb8f, 32'hc21ad1fa, 32'h42b8690b, 32'h42c783ce, 32'hc1cfb011, 32'hc2409eda, 32'h411125d7};
test_weights[19952:19959] = '{32'h416eb7ef, 32'h424c76dc, 32'hc2857a6a, 32'h4250fde9, 32'hc2ae67f4, 32'hc20a51dc, 32'hc21fe57e, 32'hc1020b12};
test_bias[2494:2494] = '{32'h42b98cbe};
test_output[2494:2494] = '{32'h445a0e2b};
test_input[19960:19967] = '{32'h41f9f567, 32'hc277631c, 32'hc16f4113, 32'hc1c25ef0, 32'hc2c7dbb6, 32'hc24f44b7, 32'hc298b88f, 32'hc2b1cca1};
test_weights[19960:19967] = '{32'hbfbfd8e8, 32'hc24916f7, 32'hc2affa48, 32'h4185ab97, 32'hc2b8d35d, 32'hc2a9a231, 32'hc2108c20, 32'h42aec0d5};
test_bias[2495:2495] = '{32'h4286b558};
test_output[2495:2495] = '{32'h4645d361};
test_input[19968:19975] = '{32'h4253d021, 32'hc1b0c26f, 32'h42a6980c, 32'h4210da38, 32'h3fea5f01, 32'h428a9259, 32'hc2c5d94e, 32'hc2a8831d};
test_weights[19968:19975] = '{32'hc28bc9ef, 32'h42b3eddb, 32'h41fc077d, 32'hc24844a5, 32'hc1909b57, 32'h42c2676f, 32'hc100e6f1, 32'h4291cf9b};
test_bias[2496:2496] = '{32'hc2c063ec};
test_output[2496:2496] = '{32'hc562225c};
test_input[19976:19983] = '{32'hc2aed541, 32'hc29db9e9, 32'hc29c4461, 32'hc2b1d7f9, 32'h42af8e78, 32'hc2b635b8, 32'hc0dfa544, 32'hc246d799};
test_weights[19976:19983] = '{32'h427efcf3, 32'hc1cf0a06, 32'hc2939f4f, 32'hc0f4374a, 32'hc2c2d4b3, 32'hbf75eab5, 32'h42b746c6, 32'h42981fd8};
test_bias[2497:2497] = '{32'h4203afee};
test_output[2497:2497] = '{32'hc61b4787};
test_input[19984:19991] = '{32'hc1046aae, 32'h41bc93ab, 32'hc2662df7, 32'hc282be5f, 32'h42445bb0, 32'h428f82be, 32'h427506bb, 32'hc29237f0};
test_weights[19984:19991] = '{32'h421b2dbe, 32'h428533d0, 32'h426c2d93, 32'h42b6d494, 32'hc146a210, 32'hc1bdf47a, 32'hc2248df2, 32'hc203f8d6};
test_bias[2498:2498] = '{32'h428ce5d9};
test_output[2498:2498] = '{32'hc623ae02};
test_input[19992:19999] = '{32'hc2a955fb, 32'hc18878d2, 32'h3ff91821, 32'hc20b59dc, 32'hc2bef963, 32'h423f7bbb, 32'hc03c2a34, 32'h423eb93f};
test_weights[19992:19999] = '{32'hc1971b13, 32'hc25a495b, 32'h4187c15f, 32'h4293055c, 32'hc280507a, 32'h417c65c8, 32'hc285c0bf, 32'h429964fe};
test_bias[2499:2499] = '{32'h42a476a9};
test_output[2499:2499] = '{32'h46290dbb};
test_input[20000:20007] = '{32'h42b28f0c, 32'hc1ac62c1, 32'hc27f4722, 32'h4048fba7, 32'hc2a1a3f6, 32'hc2290cdb, 32'h4296ef49, 32'hc27e7fbd};
test_weights[20000:20007] = '{32'hc11e9493, 32'h41bb4af2, 32'h425a9047, 32'hc1892ed4, 32'hc2900801, 32'hc124de45, 32'h42bc7e4c, 32'hc1dfface};
test_bias[2500:2500] = '{32'h412e3ff3};
test_output[2500:2500] = '{32'h461fd8e2};
test_input[20008:20015] = '{32'hc2199ad5, 32'hc1227bc2, 32'hc2423488, 32'h4250f410, 32'h41b82688, 32'h421884c1, 32'h428550a4, 32'hc29f4282};
test_weights[20008:20015] = '{32'hc2b1dc0b, 32'h42391468, 32'hc2aa029e, 32'hc2a78034, 32'h4299c4b7, 32'hc2a1189c, 32'h4180120f, 32'h3f8a32f5};
test_bias[2501:2501] = '{32'hc2b3bdc7};
test_output[2501:2501] = '{32'h450ef086};
test_input[20016:20023] = '{32'hc2b4c065, 32'h410fd64d, 32'h427cacb6, 32'hc229d446, 32'h41d61d40, 32'h42921ff2, 32'h42c4d2c0, 32'hc27b7cfd};
test_weights[20016:20023] = '{32'hc0c6f834, 32'h42277f9b, 32'hc23ded91, 32'hc23b23f2, 32'h42b0ce16, 32'hc2b1d22a, 32'h42b2ddfb, 32'hc1ac4c78};
test_bias[2502:2502] = '{32'h4275b853};
test_output[2502:2502] = '{32'h45bbe1cb};
test_input[20024:20031] = '{32'h42a97c64, 32'hc22f47c4, 32'h423e6fdc, 32'hc2afc4e2, 32'hc288c264, 32'h42ad1685, 32'hc2941c8c, 32'hc2859742};
test_weights[20024:20031] = '{32'hc00314d4, 32'h4102799c, 32'hc1e2930f, 32'h41ab7d20, 32'hc23d9037, 32'h429a60a3, 32'h41362959, 32'h418c53b3};
test_bias[2503:2503] = '{32'h421dddab};
test_output[2503:2503] = '{32'h4582b250};
test_input[20032:20039] = '{32'h421ce9c4, 32'hc27aeeed, 32'h42a53026, 32'h4210f5c7, 32'hc25b0d19, 32'hc2527191, 32'h4276407d, 32'hc22a9302};
test_weights[20032:20039] = '{32'h42ba2e16, 32'h421a0ebe, 32'hc235703d, 32'hc261f7d1, 32'h42832a9f, 32'hc24a5cd8, 32'hc2163f0d, 32'h422ae1ea};
test_bias[2504:2504] = '{32'h42327411};
test_output[2504:2504] = '{32'hc615a61d};
test_input[20040:20047] = '{32'hc2786638, 32'h41a7f689, 32'hc043dd39, 32'h42be19d8, 32'h42b7a144, 32'h42aec477, 32'hc241ebdc, 32'hc25a0031};
test_weights[20040:20047] = '{32'hc2bbfeb1, 32'hc2a30098, 32'h40947d6f, 32'hc24059a6, 32'hc082021f, 32'h42282c74, 32'hc2b8a66d, 32'h42a72703};
test_bias[2505:2505] = '{32'hc22cea1c};
test_output[2505:2505] = '{32'h4529fd23};
test_input[20048:20055] = '{32'hc2846616, 32'hc0d6ba81, 32'h42282b58, 32'hc16705ad, 32'hc100877a, 32'hc132b71c, 32'hc23fb45b, 32'hbf8884b1};
test_weights[20048:20055] = '{32'hc2bb2dca, 32'hc26bb7bc, 32'hc1d3e8ce, 32'h417c09af, 32'hc28d5ac0, 32'h420d4c30, 32'h42159795, 32'hc1e28492};
test_bias[2506:2506] = '{32'hc08a4b95};
test_output[2506:2506] = '{32'h45648a14};
test_input[20056:20063] = '{32'hc1bc7e46, 32'hc1ce7ce3, 32'h410316d0, 32'hc28f8bdb, 32'h427b91b3, 32'h42ae4faf, 32'hc25cdb0b, 32'h42a09aa3};
test_weights[20056:20063] = '{32'hc29ea7f8, 32'h410bb001, 32'h42b0f9e8, 32'h4115977c, 32'hc24c2a9f, 32'h41fd6b06, 32'hc15d1946, 32'hc218ebd4};
test_bias[2507:2507] = '{32'hc1a791e7};
test_output[2507:2507] = '{32'hc486f007};
test_input[20064:20071] = '{32'hc23a0144, 32'hc285ac08, 32'hc1b7a1b4, 32'h428b88aa, 32'hc2297a19, 32'h411c0676, 32'h421cca79, 32'h4199a9ab};
test_weights[20064:20071] = '{32'h428f3d16, 32'hc2971b34, 32'hc2776981, 32'h4192f496, 32'hc2c191fb, 32'h425580b8, 32'h409df5b4, 32'h4112cc90};
test_bias[2508:2508] = '{32'h4229a491};
test_output[2508:2508] = '{32'h4613b7e4};
test_input[20072:20079] = '{32'hc24a8539, 32'hc298a3fc, 32'hc21c45de, 32'hc2bab60d, 32'h4172eac8, 32'hc25aee60, 32'h3ffa06ed, 32'h3f35217f};
test_weights[20072:20079] = '{32'h4207ec1c, 32'h42973200, 32'h42567fb6, 32'hc21551ce, 32'h429a228a, 32'hc295fb93, 32'h426e0afd, 32'hc2ae387f};
test_bias[2509:2509] = '{32'h424e954a};
test_output[2509:2509] = '{32'hc433d5c4};
test_input[20080:20087] = '{32'hc21abdcd, 32'h424a45a4, 32'h41575959, 32'hc299d0e8, 32'hc2ada9d2, 32'hc297f08f, 32'h424eb02d, 32'hc0bf8c4a};
test_weights[20080:20087] = '{32'hc2644df5, 32'hc25d9da7, 32'h4281a98f, 32'h4205da4b, 32'h425e34e7, 32'h426fd751, 32'hc234ddb8, 32'hc16a937b};
test_bias[2510:2510] = '{32'hc2c549ec};
test_output[2510:2510] = '{32'hc65b132d};
test_input[20088:20095] = '{32'hc29c5d65, 32'h41ae20b3, 32'h41cac971, 32'hc2972c3e, 32'hc151f357, 32'hc10dc4de, 32'hc28f99ba, 32'hc27f270f};
test_weights[20088:20095] = '{32'h3fd5f729, 32'h425a4fa1, 32'h4229f59a, 32'h4229a5a1, 32'hc21d80ae, 32'hc1d0d678, 32'h4125cbf8, 32'h41817edf};
test_bias[2511:2511] = '{32'hc21c0800};
test_output[2511:2511] = '{32'hc505b075};
test_input[20096:20103] = '{32'h40f36f6f, 32'h41f11ede, 32'h420176b6, 32'h42c62a46, 32'h42973c74, 32'hc12a104c, 32'h4288dd08, 32'hc1e9a7f0};
test_weights[20096:20103] = '{32'hc29805f4, 32'hc28665f8, 32'h4292a71d, 32'h41ccaf0f, 32'hc2892497, 32'h42a92a83, 32'hc23b85f5, 32'hc29c8e0e};
test_bias[2512:2512] = '{32'hc29fae77};
test_output[2512:2512] = '{32'hc5956a41};
test_input[20104:20111] = '{32'h42aed6a5, 32'hc1127037, 32'h424d26f8, 32'hc07cc232, 32'hc2b2aa88, 32'h42aa9270, 32'hc2a518e4, 32'h42195316};
test_weights[20104:20111] = '{32'hc0f135c6, 32'h423221c4, 32'h429d1c6d, 32'hc2be8e58, 32'hc25d552a, 32'hc269f497, 32'hc288bc13, 32'h41d72b02};
test_bias[2513:2513] = '{32'h42272a48};
test_output[2513:2513] = '{32'h461c678d};
test_input[20112:20119] = '{32'hc1e6da7e, 32'hc246a137, 32'h422393c5, 32'hc23d3d8e, 32'hc20add4c, 32'h4111c339, 32'hc2c3f306, 32'hc28b2ca2};
test_weights[20112:20119] = '{32'hc22852e5, 32'hc1779147, 32'hc102292b, 32'h425dae38, 32'hc2b4fc9b, 32'hc286786e, 32'h41d5c949, 32'hc24aaf1a};
test_bias[2514:2514] = '{32'hc0d2cf28};
test_output[2514:2514] = '{32'h4519a5e3};
test_input[20120:20127] = '{32'hc2b14a04, 32'hc23531c0, 32'h42a9f8dc, 32'h41e09c59, 32'h427868e0, 32'hc27170c7, 32'h429ad6c4, 32'hc1e65647};
test_weights[20120:20127] = '{32'hc2ba9608, 32'h415fd992, 32'h41a174ad, 32'h427b0355, 32'h41b36b43, 32'h3e9e7ef8, 32'hc2bcc881, 32'h40edcb46};
test_bias[2515:2515] = '{32'h42be74dc};
test_output[2515:2515] = '{32'h459e26ed};
test_input[20128:20135] = '{32'h4298b816, 32'hc27d4c75, 32'hc25fc55e, 32'h4281f2de, 32'h429bf622, 32'hc1d81387, 32'hc212ec53, 32'h42b3eb75};
test_weights[20128:20135] = '{32'hc21fda1a, 32'h421bd622, 32'h4224a081, 32'hc1dc8af6, 32'h405e01cc, 32'hc18bf816, 32'h42834acc, 32'hc2ae6c9d};
test_bias[2516:2516] = '{32'h42c233d9};
test_output[2516:2516] = '{32'hc694a9d2};
test_input[20136:20143] = '{32'h4212c703, 32'hc225d281, 32'h4215ae9d, 32'h42975e44, 32'hc20f5bf4, 32'h41677220, 32'h42634ae4, 32'h427e80df};
test_weights[20136:20143] = '{32'h4264a8f4, 32'h429f89ec, 32'hc29e47e5, 32'h422e4056, 32'hc24b69d2, 32'h4226288e, 32'h4072b2c5, 32'h42350527};
test_bias[2517:2517] = '{32'hc2a5519c};
test_output[2517:2517] = '{32'h458e8fa9};
test_input[20144:20151] = '{32'h421436a5, 32'hc2442da6, 32'hc2b9be23, 32'hc18ec4a0, 32'h4258eb45, 32'h4290b13a, 32'h42bf8ea7, 32'hc1a2f9c9};
test_weights[20144:20151] = '{32'hc201d281, 32'hc2a287b7, 32'h429468b8, 32'hc29474ef, 32'hc268c120, 32'hc264f149, 32'h4273ecb4, 32'hc1588283};
test_bias[2518:2518] = '{32'hc21b98a1};
test_output[2518:2518] = '{32'hc57a2a3f};
test_input[20152:20159] = '{32'hc2adae1c, 32'hc210427d, 32'h42b72db4, 32'h42054085, 32'h421504ef, 32'hc2a2917a, 32'h429ac4e0, 32'hc2b2f400};
test_weights[20152:20159] = '{32'h42920bb3, 32'h42aadfe7, 32'h410910a3, 32'hc1bc1f8a, 32'hc2a0cf6e, 32'hc23d12dc, 32'h4110071c, 32'h4294e58f};
test_bias[2519:2519] = '{32'h42bbbbdf};
test_output[2519:2519] = '{32'hc661b65c};
test_input[20160:20167] = '{32'hc29853a9, 32'h42beded3, 32'h42901c53, 32'h42a0e161, 32'h426dc4ce, 32'h4296c441, 32'hc1e49ebe, 32'hc1c89516};
test_weights[20160:20167] = '{32'h415f41dc, 32'hc28cebf0, 32'h42b6301e, 32'h42ab747c, 32'hc2621963, 32'hc2496445, 32'hc2c029ae, 32'h42c547a7};
test_bias[2520:2520] = '{32'hc2336c7a};
test_output[2520:2520] = '{32'hc49ce23b};
test_input[20168:20175] = '{32'hc2bf935a, 32'hbf317788, 32'h405ecca6, 32'hc0bc7b0a, 32'h4299f490, 32'h40b42edc, 32'hc293699b, 32'hc2c6f07a};
test_weights[20168:20175] = '{32'h42709b7a, 32'hc2900904, 32'h40ef872e, 32'h3fd35a39, 32'hc24200bc, 32'hc2bdac59, 32'h42577870, 32'hc26c098f};
test_bias[2521:2521] = '{32'hc108c1c0};
test_output[2521:2521] = '{32'hc5fc4281};
test_input[20176:20183] = '{32'hc1e4198a, 32'h424e2219, 32'h41a0731b, 32'h429a7f07, 32'h420564f0, 32'h41e50420, 32'h426f82d2, 32'h4284ee1f};
test_weights[20176:20183] = '{32'h421e70bd, 32'h41cb27f8, 32'h4259c312, 32'hc2ba8233, 32'h3d0cfd63, 32'h429285de, 32'h42a4dbd0, 32'hc2bbb7e7};
test_bias[2522:2522] = '{32'hc220144a};
test_output[2522:2522] = '{32'hc5a1c6da};
test_input[20184:20191] = '{32'hc19385ce, 32'h4248d73a, 32'h410894a8, 32'hc1c47286, 32'hc2aa1a96, 32'hc2b89b51, 32'h4186f654, 32'hc125485d};
test_weights[20184:20191] = '{32'hc1b07bf3, 32'hc257b3ad, 32'hc2b37474, 32'h4294bb23, 32'h4294afda, 32'hc2a0eccd, 32'h42679727, 32'hc2b9679f};
test_bias[2523:2523] = '{32'h42619e4a};
test_output[2523:2523] = '{32'hc4e0c567};
test_input[20192:20199] = '{32'h411bcce1, 32'hc2936633, 32'hc271cdcc, 32'hc1dfccf3, 32'hc2ad1d69, 32'hc286f0c0, 32'hc1e74973, 32'hc23a4187};
test_weights[20192:20199] = '{32'h429a976d, 32'h42457409, 32'h418662eb, 32'hc1fac91a, 32'hbfa682b1, 32'h4233ce6a, 32'h41a68536, 32'hc2bd103e};
test_bias[2524:2524] = '{32'h41d31052};
test_output[2524:2524] = '{32'hc5045cf6};
test_input[20200:20207] = '{32'h41e24691, 32'hc11a45ad, 32'h41a29c00, 32'h4135612a, 32'h42a52bf1, 32'hc2a20e42, 32'h41235902, 32'h41e9cb5c};
test_weights[20200:20207] = '{32'h41f0377c, 32'hc16ede78, 32'hc22baa40, 32'h42a88f4e, 32'h4299b2a9, 32'hc218c0b0, 32'h42316ce4, 32'h428408f3};
test_bias[2525:2525] = '{32'h4230c34a};
test_output[2525:2525] = '{32'h464a3e84};
test_input[20208:20215] = '{32'h4231906f, 32'h4279c075, 32'h42870eb5, 32'hc1401544, 32'hc28649ed, 32'h428794bb, 32'h42acd728, 32'hc2833dab};
test_weights[20208:20215] = '{32'hc0bc25c9, 32'hc11bf676, 32'hc2b746f0, 32'h42955ad6, 32'h4273ce4f, 32'h423ac177, 32'hc2747fd2, 32'h42687a36};
test_bias[2526:2526] = '{32'h414bcd59};
test_output[2526:2526] = '{32'hc68c5aba};
test_input[20216:20223] = '{32'h4174abe1, 32'hc27c5cb9, 32'hc2847e56, 32'hc21526c6, 32'hbfca00ea, 32'hc166ce0b, 32'h4128f12d, 32'h42a2e1b3};
test_weights[20216:20223] = '{32'h4234348a, 32'h428326ef, 32'h425ce8e7, 32'hc25bcb3c, 32'h41787c7c, 32'hc288e96a, 32'hc1a73d35, 32'hc0d16d6f};
test_bias[2527:2527] = '{32'hc2c79b84};
test_output[2527:2527] = '{32'hc59aa4a4};
test_input[20224:20231] = '{32'hc2a2ddeb, 32'hc21123fe, 32'hc15e1a5b, 32'h41558534, 32'hc1b363c9, 32'h425e363f, 32'hc2a0d206, 32'hc24cd5c5};
test_weights[20224:20231] = '{32'hc07aae36, 32'hc284dfb3, 32'hc201b830, 32'h4068735f, 32'hc1d8063c, 32'hc256a1b4, 32'h425aa39b, 32'hc2aff2b5};
test_bias[2528:2528] = '{32'h429ac125};
test_output[2528:2528] = '{32'h448204c3};
test_input[20232:20239] = '{32'h4241ec67, 32'hc2c4592f, 32'hc28a8739, 32'hc2994a59, 32'h419d5d8d, 32'h42b17003, 32'hc2329494, 32'hc1c55e56};
test_weights[20232:20239] = '{32'h4136dbf1, 32'hc2b9efa7, 32'h401c6b35, 32'hc2c22875, 32'hc2b7add3, 32'h42afc780, 32'h420fc4a8, 32'hc2c6468d};
test_bias[2529:2529] = '{32'h4280f866};
test_output[2529:2529] = '{32'h46ba5230};
test_input[20240:20247] = '{32'h429f2865, 32'h418eee86, 32'hc2a3f776, 32'hc28e072a, 32'hc2851ab0, 32'hc2853c39, 32'hc2a5765d, 32'hc24ff4b4};
test_weights[20240:20247] = '{32'h4217a2aa, 32'h425602ce, 32'h42b3c192, 32'h422306be, 32'hc2423fb5, 32'h42c48e4e, 32'hc20c88f4, 32'h41e15b8b};
test_bias[2530:2530] = '{32'h422942e3};
test_output[2530:2530] = '{32'hc5fdc674};
test_input[20248:20255] = '{32'h42c53a4d, 32'hc1e3f9db, 32'hc148b2e5, 32'hc25fae5c, 32'h4263eef1, 32'h42846b98, 32'h41cb0965, 32'hc28d3a6b};
test_weights[20248:20255] = '{32'h42acff9f, 32'hc2b16bda, 32'hc201581c, 32'hc276275f, 32'hc183be0e, 32'hc2311008, 32'h42364981, 32'hc0e19abb};
test_bias[2531:2531] = '{32'h4243bfb2};
test_output[2531:2531] = '{32'h46470c12};
test_input[20256:20263] = '{32'h42ac489c, 32'hc19a91ef, 32'hc2b5dd76, 32'h411d4eba, 32'h42a82be3, 32'hc2646eaa, 32'hc2ac1707, 32'h41e2471d};
test_weights[20256:20263] = '{32'h4291c53d, 32'hc28b3cce, 32'hc1b0ccf2, 32'h415a1ac0, 32'h4274b3b9, 32'hc23ac7fe, 32'hc22652b0, 32'hc2039c0a};
test_bias[2532:2532] = '{32'h42a78060};
test_output[2532:2532] = '{32'h469ea9a4};
test_input[20264:20271] = '{32'hc283e181, 32'h41c849b4, 32'hc180f870, 32'h42765e86, 32'h424647e2, 32'h42c7fa3f, 32'h42628e72, 32'h422f583b};
test_weights[20264:20271] = '{32'h41d2defe, 32'hc2b8827e, 32'h40762015, 32'h42c06b6f, 32'h3f88567e, 32'h42b04e74, 32'h425aa671, 32'h42ba709b};
test_bias[2533:2533] = '{32'h4125d2e9};
test_output[2533:2533] = '{32'h468ba7d5};
test_input[20272:20279] = '{32'h410fd0c6, 32'hc2a8ef41, 32'hc2b6c114, 32'h42ae336b, 32'h42b35eab, 32'h42358ed9, 32'h42b29b8c, 32'hc2c22835};
test_weights[20272:20279] = '{32'h41f4e07f, 32'h4200908b, 32'h424c4b32, 32'h42a433fa, 32'h42288a56, 32'h403adf17, 32'h41621edb, 32'hc22949af};
test_bias[2534:2534] = '{32'h3fb028f7};
test_output[2534:2534] = '{32'h4611bf4b};
test_input[20280:20287] = '{32'hc2b53e0a, 32'h42881456, 32'h4280f03f, 32'hc19f9faa, 32'h42631e58, 32'hc1357d65, 32'hc25b436e, 32'hc2b9a3c4};
test_weights[20280:20287] = '{32'h42b56ecf, 32'h41485b19, 32'hc2bbe86b, 32'h427077d4, 32'h429b49cd, 32'hc29fe0e5, 32'h426d8df1, 32'hc285d5b6};
test_bias[2535:2535] = '{32'h42b8e983};
test_output[2535:2535] = '{32'hc5c3ae94};
test_input[20288:20295] = '{32'hc28ada0b, 32'h429e9613, 32'hc22fa718, 32'hc2ae5fd9, 32'h42b1bac2, 32'h41f37234, 32'hc23bd5ab, 32'h40d9a1af};
test_weights[20288:20295] = '{32'h418b6071, 32'h4287d248, 32'h42893678, 32'hc16a2ca2, 32'hc285e2ae, 32'h41291205, 32'h42b4905f, 32'h42822584};
test_bias[2536:2536] = '{32'h424e9a66};
test_output[2536:2536] = '{32'hc5d8af9f};
test_input[20296:20303] = '{32'h41052235, 32'hc237295f, 32'h4252550e, 32'h41ac4bf7, 32'hc29aec94, 32'h41d9090a, 32'h421b0f25, 32'h42851fe4};
test_weights[20296:20303] = '{32'hc0ed07b2, 32'h4299689f, 32'hc24afe68, 32'h42c4b213, 32'hc046e4b5, 32'hc28ac59e, 32'hc2927cec, 32'hc2820633};
test_bias[2537:2537] = '{32'h41ce2b18};
test_output[2537:2537] = '{32'hc649ab87};
test_input[20304:20311] = '{32'h4199ff46, 32'h42549805, 32'h4298a4ca, 32'hc2904a4b, 32'h41b40843, 32'hc2a3dd40, 32'h4277e476, 32'h4173e7a6};
test_weights[20304:20311] = '{32'h41db3c0a, 32'h41fbb61a, 32'h411a6a2e, 32'hc025fd52, 32'hc224f7d7, 32'h428fb0bc, 32'hc11a98ae, 32'h418e4acd};
test_bias[2538:2538] = '{32'h42793672};
test_output[2538:2538] = '{32'hc57746d8};
test_input[20312:20319] = '{32'hbfc87659, 32'h4212027e, 32'h427c43b0, 32'hc290a545, 32'hc1c3d500, 32'hc27e1698, 32'h42b6066b, 32'hc1456165};
test_weights[20312:20319] = '{32'h42bc8a44, 32'h4206e245, 32'hc1609cfd, 32'h42953b82, 32'h426efc5b, 32'h4234bfbb, 32'hc2186c75, 32'h41819255};
test_bias[2539:2539] = '{32'hc28b587a};
test_output[2539:2539] = '{32'hc64f5432};
test_input[20320:20327] = '{32'h41ec5a93, 32'hc16d9310, 32'h42338d67, 32'hc2c21f44, 32'h42c09dc4, 32'h427dae77, 32'hc232eea7, 32'hc2b1df9d};
test_weights[20320:20327] = '{32'hc1c62e61, 32'h4245f23f, 32'h4227e062, 32'h429d18b1, 32'hc2b8d929, 32'h4254ded9, 32'hc2106dd4, 32'h407854ab};
test_bias[2540:2540] = '{32'h42b61d79};
test_output[2540:2540] = '{32'hc631aed3};
test_input[20328:20335] = '{32'hc177f583, 32'h42850c35, 32'hc2bcd6c4, 32'hc0a287da, 32'h419bbe05, 32'hc0a81ed6, 32'h41ccb20d, 32'h42af83da};
test_weights[20328:20335] = '{32'h424d38ff, 32'hc212c749, 32'h42a3b939, 32'hc2ad276b, 32'h4253deee, 32'hc1ad76e4, 32'h42aa5446, 32'hbf7868cf};
test_bias[2541:2541] = '{32'h42be9d85};
test_output[2541:2541] = '{32'hc5e0bb99};
test_input[20336:20343] = '{32'hc27e7afd, 32'hc2b03716, 32'hc2716285, 32'hc2b3cbcd, 32'hc0dad756, 32'hc29638a8, 32'hc10be565, 32'hc1b68829};
test_weights[20336:20343] = '{32'hc1c5b011, 32'hc2b3eb69, 32'h4217f20b, 32'hc1e55ea5, 32'hc2ae3288, 32'hc2592100, 32'h3e49954c, 32'hc223b699};
test_bias[2542:2542] = '{32'h41651c77};
test_output[2542:2542] = '{32'h4670aaad};
test_input[20344:20351] = '{32'h421b6426, 32'h423e64ef, 32'hc25be48c, 32'hc113f279, 32'h423734a4, 32'hc2a46ac0, 32'h4255b125, 32'h412cec91};
test_weights[20344:20351] = '{32'h4143ac87, 32'hc220060a, 32'h42868edc, 32'hc28ddc81, 32'hc02e5e41, 32'h421f79ec, 32'h42c423f6, 32'hc28f9432};
test_bias[2543:2543] = '{32'h409155f1};
test_output[2543:2543] = '{32'hc554e4b7};
test_input[20352:20359] = '{32'hc0a12646, 32'hc2c38073, 32'hc15aa78e, 32'h4295efa9, 32'hc2c482a5, 32'h421ac55c, 32'hc271edfd, 32'h42a4ce38};
test_weights[20352:20359] = '{32'h42b444d2, 32'hc2c7769b, 32'hc29d54a6, 32'hc022029a, 32'h42683f71, 32'hc2ae36e5, 32'hc2ba916c, 32'hc271a0d3};
test_bias[2544:2544] = '{32'h42009585};
test_output[2544:2544] = '{32'h44e12c31};
test_input[20360:20367] = '{32'h41633def, 32'h42b8b307, 32'h429e8204, 32'hc253d78f, 32'hc2a56c96, 32'h40aade50, 32'h42c4e5b3, 32'h4280569c};
test_weights[20360:20367] = '{32'h41715d26, 32'h42a9e16f, 32'h411be1ff, 32'h429aa6cf, 32'hc26a8dc1, 32'h42b475be, 32'hc2bf9b96, 32'h42c1ecf5};
test_bias[2545:2545] = '{32'hc2482b59};
test_output[2545:2545] = '{32'h45d4bc16};
test_input[20368:20375] = '{32'hc28590b6, 32'hc17ce295, 32'h42ab7665, 32'hc2b79d1c, 32'h40696b71, 32'hc2b9f200, 32'hc295d701, 32'hc18d0e9a};
test_weights[20368:20375] = '{32'hc14d5db6, 32'h42c40e8d, 32'h417131c7, 32'h42a43297, 32'hc28612d1, 32'h4207c894, 32'hc284ca00, 32'hc299d0ef};
test_bias[2546:2546] = '{32'hc246b854};
test_output[2546:2546] = '{32'hc57d8f0f};
test_input[20376:20383] = '{32'hc1d5cf59, 32'hc1c649e7, 32'hc206be97, 32'hc29144ce, 32'h422cfeb4, 32'hc2c315d4, 32'hc285b2ac, 32'h41758ed9};
test_weights[20376:20383] = '{32'hc10ffdfc, 32'h42a5a3cd, 32'h429a5096, 32'h41ff3aba, 32'h4294f59a, 32'hc264db4e, 32'h42273680, 32'hc22038b1};
test_bias[2547:2547] = '{32'hc1fe7060};
test_output[2547:2547] = '{32'hc4aaf8ce};
test_input[20384:20391] = '{32'hc29cf1c1, 32'h42ac8e16, 32'h429d97be, 32'hc1d03586, 32'hc29ba245, 32'h42b2a723, 32'h4249c41a, 32'hc28f6c21};
test_weights[20384:20391] = '{32'hc1001328, 32'h429088c2, 32'hc2baaf01, 32'hc1ab5a01, 32'h429d6517, 32'h42611158, 32'h4185ccad, 32'hc10b78c6};
test_bias[2548:2548] = '{32'hc17750e4};
test_output[2548:2548] = '{32'h43d284e5};
test_input[20392:20399] = '{32'hc176164a, 32'h41cc22cc, 32'h428ef9be, 32'hc29f3be1, 32'hc1e44467, 32'h421ccd59, 32'h4064867a, 32'h4216f0a6};
test_weights[20392:20399] = '{32'hc049fa4c, 32'hc16f5595, 32'hc270c1b8, 32'h42c0e089, 32'h42c35a9f, 32'hc10123b5, 32'hc27c42c2, 32'h41a60d0d};
test_bias[2549:2549] = '{32'h423ee72d};
test_output[2549:2549] = '{32'hc6676f0a};
test_input[20400:20407] = '{32'h42381ca2, 32'h4289057e, 32'h42510fdc, 32'hc2560734, 32'h41007d02, 32'h42ba6d4f, 32'hc2777652, 32'h42ab8691};
test_weights[20400:20407] = '{32'hc2a864df, 32'hc103e05e, 32'h42b9864d, 32'h428c164c, 32'hc2afe789, 32'hc22182b3, 32'hc1e54543, 32'h42834164};
test_bias[2550:2550] = '{32'hc1b029a7};
test_output[2550:2550] = '{32'hc3d72756};
test_input[20408:20415] = '{32'hc193506e, 32'h4193f41e, 32'h41484548, 32'h42ad0abf, 32'hc22dfd37, 32'hc1fbe0c6, 32'hc15b9d1c, 32'hc1c148d3};
test_weights[20408:20415] = '{32'hc275ad01, 32'hc0227995, 32'h41410b2c, 32'h419a667b, 32'h4231f342, 32'hc2b4965a, 32'h41eff2bc, 32'h4251359c};
test_bias[2551:2551] = '{32'hc22dbc43};
test_output[2551:2551] = '{32'h4502dec5};
test_input[20416:20423] = '{32'h427c5d19, 32'h4257b726, 32'h410158ad, 32'h426c2c9f, 32'hc2af33b1, 32'h407b1e15, 32'h429ae636, 32'h4295bda8};
test_weights[20416:20423] = '{32'h42968663, 32'h4291e5de, 32'hc24e29bc, 32'h42a53fca, 32'h42b5a4e8, 32'hc2b1d0fb, 32'h42b8acb7, 32'hc2b29171};
test_bias[2552:2552] = '{32'hc279502e};
test_output[2552:2552] = '{32'h45a3dd93};
test_input[20424:20431] = '{32'hc2afb411, 32'h41e70475, 32'hc2398134, 32'hc2b98894, 32'h423590c4, 32'h42810da9, 32'hc241caa2, 32'h42b4772d};
test_weights[20424:20431] = '{32'h41e8e067, 32'hc2b5e50f, 32'hc181e7f9, 32'hc2a28543, 32'h425e9bcb, 32'h42bd0bee, 32'h4252756a, 32'h42588784};
test_bias[2553:2553] = '{32'hc245d8d7};
test_output[2553:2553] = '{32'h465b0c4b};
test_input[20432:20439] = '{32'hc2689f14, 32'h420269a0, 32'hc28045c3, 32'hc2a6168a, 32'h41b870ff, 32'hc1bf8f39, 32'h410c6a13, 32'h42a6d2ea};
test_weights[20432:20439] = '{32'h423a4e69, 32'hc24d6481, 32'h42c6e787, 32'hc1f59789, 32'hc2879c2c, 32'h40abc89b, 32'h42c042cd, 32'hc254f577};
test_bias[2554:2554] = '{32'h428400ea};
test_output[2554:2554] = '{32'hc651eb9f};
test_input[20440:20447] = '{32'hc2ba52b0, 32'hbf09c612, 32'h40ae22d7, 32'hc282c5f5, 32'h428ca187, 32'hc2c2647d, 32'h423ac035, 32'hc2c23035};
test_weights[20440:20447] = '{32'hc29b8b63, 32'h424b4d2c, 32'h4236ecf9, 32'h4236b1c2, 32'hc2438e89, 32'h42a218b3, 32'h41f0c5dd, 32'h42629395};
test_bias[2555:2555] = '{32'h42bda77f};
test_output[2555:2555] = '{32'hc6294aa0};
test_input[20448:20455] = '{32'hc142dc56, 32'h422dfdad, 32'hc2435250, 32'h418d441f, 32'hc2175b78, 32'h41a1891e, 32'h42c67a3d, 32'hc0c96028};
test_weights[20448:20455] = '{32'hc1fa233d, 32'h429d4bef, 32'hc22315ef, 32'hc054bc1a, 32'hc2bdee90, 32'hc1e82397, 32'h42c7ed51, 32'h42bfd482};
test_bias[2556:2556] = '{32'h4115e4f3};
test_output[2556:2556] = '{32'h468d2722};
test_input[20456:20463] = '{32'h42afc47c, 32'h3f9510d5, 32'hc290af7f, 32'hc23f37f9, 32'h41bb6f64, 32'h42b16029, 32'hbfb3c92d, 32'h4276f0dc};
test_weights[20456:20463] = '{32'hc1b79b58, 32'h4234a958, 32'hc21c26ff, 32'h42992a93, 32'hc2c7c583, 32'h42c50dc0, 32'h42c2aa7a, 32'hc29e441c};
test_bias[2557:2557] = '{32'hc2acdc7f};
test_output[2557:2557] = '{32'hc4bcfc50};
test_input[20464:20471] = '{32'h42bd39f5, 32'hc23341f2, 32'hc16f2788, 32'hc24b0994, 32'hc16c7135, 32'hc2c0d09f, 32'hc2a49184, 32'h4180cfac};
test_weights[20464:20471] = '{32'h4216448b, 32'h42953fb9, 32'h4254e2b3, 32'hc258a95d, 32'hc2acf027, 32'h42bfebdd, 32'h42b02442, 32'hc1f79906};
test_bias[2558:2558] = '{32'h41b493c7};
test_output[2558:2558] = '{32'hc6537095};
test_input[20472:20479] = '{32'hc1ca3259, 32'h41adc5ae, 32'h42334526, 32'hc2c470c4, 32'hc2a93ebc, 32'hc1ed192b, 32'h429345a8, 32'hc2c2bb94};
test_weights[20472:20479] = '{32'hc283989c, 32'hc199dc36, 32'h42a379c2, 32'hc1ff12e1, 32'h419abc1d, 32'h42932a6b, 32'h42852472, 32'h4294d010};
test_bias[2559:2559] = '{32'hc2a471fd};
test_output[2559:2559] = '{32'h44e0b9cc};
test_input[20480:20487] = '{32'hc28cca7f, 32'h427ef36c, 32'h426e71e4, 32'hc2c30ee5, 32'h420ad517, 32'h423b18c8, 32'hc28cd4dc, 32'h41a70cf3};
test_weights[20480:20487] = '{32'hc2958cb2, 32'h42846d3e, 32'h42342942, 32'hc27f8da6, 32'h42916f6a, 32'hc0df2d3e, 32'hc1df4223, 32'hc1e9ff48};
test_bias[2560:2560] = '{32'h42318513};
test_output[2560:2560] = '{32'h46abd8be};
test_input[20488:20495] = '{32'hc294c56f, 32'h41fda142, 32'hc2553f5a, 32'h42b21aad, 32'h41ef61af, 32'hc0a94d77, 32'h41bd8007, 32'h42bbe2f2};
test_weights[20488:20495] = '{32'hc106c7fe, 32'hc18de9d5, 32'h42b010c3, 32'h4287c0b1, 32'hc29c45f0, 32'h3fdd513e, 32'hc24c17c8, 32'h42784c3f};
test_bias[2561:2561] = '{32'h42768eca};
test_output[2561:2561] = '{32'h456a8da5};
test_input[20496:20503] = '{32'hc10e59b9, 32'hc22eaa62, 32'hc2c56fea, 32'h4282c77a, 32'hc2b7b990, 32'hc1879faa, 32'h42b65853, 32'hc27f3aae};
test_weights[20496:20503] = '{32'hc2abd422, 32'h425c72ac, 32'hc2c67389, 32'hc11612be, 32'h410b27e2, 32'h41c61b99, 32'hc28a8716, 32'h42ada99d};
test_bias[2562:2562] = '{32'hc0d802ca};
test_output[2562:2562] = '{32'hc5ad282e};
test_input[20504:20511] = '{32'hc2762299, 32'hc1a4053b, 32'hc2564797, 32'h3fb0dfe1, 32'h424fd717, 32'h40c5e05a, 32'h423a1bea, 32'h42bbaf6f};
test_weights[20504:20511] = '{32'hc0a4ee11, 32'hc1bae6e4, 32'hc26e0288, 32'h42a8611e, 32'hc111e3e1, 32'hc21a09cd, 32'h4261f989, 32'hc2415109};
test_bias[2563:2563] = '{32'hc2ad9e49};
test_output[2563:2563] = '{32'h44ae4efc};
test_input[20512:20519] = '{32'h42475966, 32'hc2b1bcce, 32'h4130ed4f, 32'h4073c121, 32'hc1b0873c, 32'h41d93c95, 32'hc16044d5, 32'h41938846};
test_weights[20512:20519] = '{32'hc2591d33, 32'hc2c4541f, 32'hc13e961c, 32'hc290bb3e, 32'hbfa03c57, 32'h42811b64, 32'hc2a3d59e, 32'hc230e0a3};
test_bias[2564:2564] = '{32'hc25a70c5};
test_output[2564:2564] = '{32'h45efafec};
test_input[20520:20527] = '{32'hc191834b, 32'h42a4eac3, 32'hc2a6229d, 32'hc22b71b2, 32'h41576ad9, 32'hc152844a, 32'hc226e225, 32'hc1fe0e63};
test_weights[20520:20527] = '{32'h4238b746, 32'h42426679, 32'h42c06946, 32'h40013f7d, 32'hc2aa6ae5, 32'hc2baa8b9, 32'h424e8ea4, 32'h42241a7d};
test_bias[2565:2565] = '{32'h42822727};
test_output[2565:2565] = '{32'hc600783f};
test_input[20528:20535] = '{32'hc22a4bad, 32'h429cd0c1, 32'h42a22322, 32'h41bb0b2a, 32'hc29d1979, 32'hc2871ce7, 32'hc269a6d8, 32'h41aaff35};
test_weights[20528:20535] = '{32'h4290046a, 32'h42a79513, 32'hc29c528d, 32'h42c465c5, 32'hc1c6778d, 32'hc094e87f, 32'h412d8fa7, 32'h42c3c5f0};
test_bias[2566:2566] = '{32'h42c164c3};
test_output[2566:2566] = '{32'h454d2192};
test_input[20536:20543] = '{32'hc2c065c6, 32'hc2a094ba, 32'hc25fca39, 32'h427d790c, 32'h4284b7e6, 32'hc29b2cf5, 32'hc254eda9, 32'hc1bba193};
test_weights[20536:20543] = '{32'h4194ff1c, 32'h408d0e27, 32'h3ffa22ec, 32'h42bf5bd7, 32'hc2c084af, 32'hc234abc4, 32'hc1c74245, 32'hc2918de2};
test_bias[2567:2567] = '{32'hc2938308};
test_output[2567:2567] = '{32'h4572bee1};
test_input[20544:20551] = '{32'h42943e62, 32'h42bbe418, 32'h4218e0ba, 32'h423b2192, 32'h429e70fd, 32'hc2a3ce35, 32'h429e45a3, 32'h41e647e0};
test_weights[20544:20551] = '{32'h41b2859e, 32'h424ba775, 32'hc16a60a6, 32'h42acfc9b, 32'hc1e53814, 32'h4109df29, 32'hc2a52a37, 32'h42a98d01};
test_bias[2568:2568] = '{32'hc29e03f4};
test_output[2568:2568] = '{32'h452d6150};
test_input[20552:20559] = '{32'hc223744b, 32'hc192cedd, 32'h42beea9a, 32'hc1d51fad, 32'hc2a9e8ba, 32'hc1c15a72, 32'h42c6bc39, 32'hc258753b};
test_weights[20552:20559] = '{32'hc14ca6ed, 32'hc1d2b0fc, 32'h42a292b9, 32'hc1a29317, 32'h42856770, 32'hc29958b2, 32'h42c45ff9, 32'h4293b195};
test_bias[2569:2569] = '{32'h42347baa};
test_output[2569:2569] = '{32'h46308ba1};
test_input[20560:20567] = '{32'hbf36525c, 32'hc200c9ee, 32'hc2858cdf, 32'hc0b5892c, 32'h4199f14e, 32'h4261d4a2, 32'hc295d6d9, 32'h4222474b};
test_weights[20560:20567] = '{32'hc12cfb1c, 32'hc29c6b59, 32'h42084247, 32'h42c7b882, 32'hc08d52e9, 32'h3ff51efc, 32'h42c05e7f, 32'h416fb26e};
test_bias[2570:2570] = '{32'hc2c76207};
test_output[2570:2570] = '{32'hc5da71f8};
test_input[20568:20575] = '{32'h429ff488, 32'h41fbf95e, 32'h41a1001c, 32'hc1da84b8, 32'h4279d26b, 32'hc1c90b69, 32'h42b59ada, 32'h4288f721};
test_weights[20568:20575] = '{32'h42c7555f, 32'hc0e4b32e, 32'h42c72bc9, 32'hc1c8660f, 32'hc28962a0, 32'h4288787a, 32'hc14d182b, 32'h424695ba};
test_bias[2571:2571] = '{32'hc25a1d01};
test_output[2571:2571] = '{32'h45ce967b};
test_input[20576:20583] = '{32'h42b6acf8, 32'hc2abc6aa, 32'hc2ac1aa8, 32'h417977ff, 32'h4125ad3b, 32'hc2864808, 32'h428aaaab, 32'hc1f5bbd3};
test_weights[20576:20583] = '{32'h428dc43a, 32'hc2a6e30c, 32'hc047aa22, 32'h41e97054, 32'h4236a2ae, 32'hc29356b7, 32'hc1635ab5, 32'h41cd47db};
test_bias[2572:2572] = '{32'hc29a0b25};
test_output[2572:2572] = '{32'h468c1a40};
test_input[20584:20591] = '{32'hc23c6e14, 32'h41b0dfc0, 32'h40cbeec6, 32'h41e24cb8, 32'h428002c4, 32'h411c4557, 32'h42950833, 32'hc2c09d9d};
test_weights[20584:20591] = '{32'hc2a3a0bb, 32'h426b5c58, 32'h42b95363, 32'h41956a7c, 32'h42553ee7, 32'h41a24bca, 32'hc1f704fb, 32'hc14e9dc9};
test_bias[2573:2573] = '{32'hc24d85cc};
test_output[2573:2573] = '{32'h46091e6e};
test_input[20592:20599] = '{32'h4205a773, 32'hc131f166, 32'h4144de98, 32'hc0d6de05, 32'h41e5bd81, 32'hc1318406, 32'hc2968eb8, 32'hc1acff9c};
test_weights[20592:20599] = '{32'h42005c10, 32'h42a9e21b, 32'h41b16ba9, 32'h4188ebbd, 32'h416937aa, 32'h42c38bee, 32'hc233886d, 32'hc0f48f6f};
test_bias[2574:2574] = '{32'h41c6ed00};
test_output[2574:2574] = '{32'h454743b2};
test_input[20600:20607] = '{32'h41b8f0ad, 32'h419e8782, 32'hc1da3a8c, 32'hc10e30ac, 32'h42645dd9, 32'h427c022f, 32'hc2983f49, 32'hc2325311};
test_weights[20600:20607] = '{32'h422b519d, 32'hc15d79f3, 32'hc2acbce0, 32'h429eafde, 32'h427ecfce, 32'hc10c89f1, 32'h408fbf48, 32'h41e25621};
test_bias[2575:2575] = '{32'hc0ff4c6c};
test_output[2575:2575] = '{32'h456ff02f};
test_input[20608:20615] = '{32'h42120af4, 32'hc260458e, 32'h42c35243, 32'h422a5fc7, 32'h41e5245c, 32'h425a41d6, 32'hc2bf742c, 32'h4296ed6f};
test_weights[20608:20615] = '{32'h422e12ae, 32'hc2ae936b, 32'h428211e7, 32'h427d1636, 32'h41ff3582, 32'h410cb581, 32'hc29f8bf5, 32'h408aa25b};
test_bias[2576:2576] = '{32'hc1bfb130};
test_output[2576:2576] = '{32'h46c23c8e};
test_input[20616:20623] = '{32'h417e44ae, 32'h4259f220, 32'h40c17e51, 32'h42c56b04, 32'hc0a22c27, 32'hc2b21b3c, 32'h41d8e979, 32'h42b7a1c4};
test_weights[20616:20623] = '{32'h425a2f60, 32'hc2797518, 32'hc201d79d, 32'hc1492558, 32'h424834f5, 32'hc2284b14, 32'hc19ffff9, 32'h42999ed6};
test_bias[2577:2577] = '{32'h4250044f};
test_output[2577:2577] = '{32'h45be36cc};
test_input[20624:20631] = '{32'hc2b5b9eb, 32'hc2019a94, 32'h426afa49, 32'h424ddead, 32'h428da3d2, 32'h429b7b01, 32'h40ac3035, 32'hc2a81279};
test_weights[20624:20631] = '{32'h427cab5c, 32'hc0977606, 32'hc29427b2, 32'h42000586, 32'hc24ae795, 32'h4208a653, 32'h4260ba49, 32'h411638bb};
test_bias[2578:2578] = '{32'h3f5b37d9};
test_output[2578:2578] = '{32'hc617c461};
test_input[20632:20639] = '{32'h42446a50, 32'h41682f7c, 32'hc22cb01a, 32'hc1c2a606, 32'hc1682b9c, 32'hc1ab80ff, 32'h41e7de93, 32'hc218e045};
test_weights[20632:20639] = '{32'hc233257f, 32'hc29158dc, 32'h41de11ca, 32'hc2bfbf80, 32'hc299bfb6, 32'h420bf366, 32'hc2a067b2, 32'hc28a0ce8};
test_bias[2579:2579] = '{32'hc280984d};
test_output[2579:2579] = '{32'hc4bc1acb};
test_input[20640:20647] = '{32'hc28aa1d6, 32'hc2b3d61b, 32'h429f8478, 32'hc014551a, 32'h42b37cf1, 32'hc251c9ba, 32'hc2576d19, 32'hc29ec107};
test_weights[20640:20647] = '{32'h41595848, 32'h425d2108, 32'hc1228642, 32'hc1de8f5c, 32'h428df620, 32'h4131e449, 32'hc236f373, 32'hc1581a91};
test_bias[2580:2580] = '{32'hc2a542de};
test_output[2580:2580] = '{32'h452158fb};
test_input[20648:20655] = '{32'h4212e09a, 32'hc2adacaf, 32'h42682088, 32'hc2014db0, 32'h4269a52b, 32'hc1b4e955, 32'hc232b4c8, 32'hc20987b9};
test_weights[20648:20655] = '{32'hc2044973, 32'h42b38230, 32'hc0fa74ab, 32'hc15e002f, 32'h41920bb4, 32'h42702aaf, 32'h42a27108, 32'hc210dc4d};
test_bias[2581:2581] = '{32'h427af39e};
test_output[2581:2581] = '{32'hc635a90a};
test_input[20656:20663] = '{32'hc29ee3ed, 32'h428a7601, 32'hc2bb4af3, 32'hc2149cd3, 32'hc22fead3, 32'h42af8a8b, 32'h42afb261, 32'hc28e4f1b};
test_weights[20656:20663] = '{32'h42aed191, 32'h427eddf9, 32'hc2a762fb, 32'h413322eb, 32'h41b0d486, 32'hc18c517b, 32'hc2b62a3b, 32'h40c422a0};
test_bias[2582:2582] = '{32'hc2944189};
test_output[2582:2582] = '{32'hc5bfb643};
test_input[20664:20671] = '{32'hc080a3c8, 32'h424e2f7c, 32'hc163ba09, 32'hc2a4ff5f, 32'hc1ab7a92, 32'hc152213c, 32'h42c3c79f, 32'h42bf1404};
test_weights[20664:20671] = '{32'hc2b708c3, 32'h424cca18, 32'hc290321e, 32'hc28881cd, 32'h419cddac, 32'h427a30e5, 32'h42bb7d88, 32'h419f5861};
test_bias[2583:2583] = '{32'h413ac870};
test_output[2583:2583] = '{32'h4698730d};
test_input[20672:20679] = '{32'hc046e13d, 32'hc2baf280, 32'hc2a3a9c1, 32'hc28f7059, 32'hc221ff57, 32'h4268ea83, 32'hc25c2262, 32'h42a1e364};
test_weights[20672:20679] = '{32'h4278a57f, 32'h4283d0d4, 32'hc2691abb, 32'hc211e60d, 32'h424ad264, 32'h42a1d560, 32'h4220a4ad, 32'hc2bda6de};
test_bias[2584:2584] = '{32'hc2abbd8f};
test_output[2584:2584] = '{32'hc5c45463};
test_input[20680:20687] = '{32'h4189fae5, 32'hc271228b, 32'hc2babe06, 32'hc1b10a25, 32'hc28ec6fb, 32'h42c13632, 32'hc24e90f5, 32'hc25e254d};
test_weights[20680:20687] = '{32'hc1058ebe, 32'hc12ff894, 32'hc27df77c, 32'hc28e25c1, 32'h406719a9, 32'hc2c3b9e3, 32'hc27222c7, 32'hc2a4e521};
test_bias[2585:2585] = '{32'h42a973c7};
test_output[2585:2585] = '{32'h45be8f36};
test_input[20688:20695] = '{32'hc2250f52, 32'h428be51a, 32'hc246c3b8, 32'h427ceda7, 32'h424e545f, 32'hc1e51599, 32'h4299922b, 32'hc2b714ca};
test_weights[20688:20695] = '{32'hbfca6f52, 32'hc27ab213, 32'hc2b20f16, 32'h41b461a3, 32'hc2b0f0a9, 32'h420f1e06, 32'hc2bbca8e, 32'h42958561};
test_bias[2586:2586] = '{32'hc29a2e7a};
test_output[2586:2586] = '{32'hc68e16ff};
test_input[20696:20703] = '{32'h42164ecc, 32'hc2aef4f3, 32'h4299baa1, 32'hc2bd788e, 32'h41b93387, 32'hc29db403, 32'hc29a4bb3, 32'h428acfb0};
test_weights[20696:20703] = '{32'h42c05a92, 32'h428c67d1, 32'hc2b60152, 32'h4186059e, 32'h422657c4, 32'hc2bc1b6e, 32'h4232b07f, 32'hc2be0444};
test_bias[2587:2587] = '{32'h4298e045};
test_output[2587:2587] = '{32'hc64658d1};
test_input[20704:20711] = '{32'hc28c176f, 32'hc1960249, 32'h42b3c2c2, 32'hc253338d, 32'h41c86fc5, 32'hc22f62a0, 32'h42851b18, 32'hc1f61bf8};
test_weights[20704:20711] = '{32'h428557bf, 32'h424fc47f, 32'hc2146ffe, 32'h42194ba6, 32'h41e9357d, 32'h41c3ca32, 32'hc1cfba16, 32'hc2a489bd};
test_bias[2588:2588] = '{32'h4233b556};
test_output[2588:2588] = '{32'hc62407b7};
test_input[20712:20719] = '{32'h428a5a45, 32'h42ae97de, 32'hc2c544be, 32'hbfd164bc, 32'h42632cf9, 32'h42430c5b, 32'h41a4309a, 32'hc274e70a};
test_weights[20712:20719] = '{32'h4223bf7e, 32'h42204b4e, 32'hc2455a60, 32'hc2bc8f1f, 32'h42299252, 32'h42c42727, 32'h42add67f, 32'hc2c5261e};
test_bias[2589:2589] = '{32'h423b95d1};
test_output[2589:2589] = '{32'h46ce4df5};
test_input[20720:20727] = '{32'h4299424b, 32'h42436c52, 32'h40e927cc, 32'h4226ca60, 32'hc1cabdb1, 32'h420a11a9, 32'hc07dfbf8, 32'hc21fce54};
test_weights[20720:20727] = '{32'hc29224dc, 32'hc187f76f, 32'hc2ad854f, 32'h426a472b, 32'h42abd5a8, 32'h421ed0b8, 32'hc10ec588, 32'h425b4878};
test_bias[2590:2590] = '{32'hc2c5d6fe};
test_output[2590:2590] = '{32'hc5f002a6};
test_input[20728:20735] = '{32'h4226b8aa, 32'h41dd4089, 32'hc29337b1, 32'h42baac71, 32'h426b6a0b, 32'h415dca28, 32'h42875910, 32'hc217affa};
test_weights[20728:20735] = '{32'h423cce87, 32'h41658581, 32'h409e8568, 32'hc29c15fe, 32'hc29fad20, 32'hc2a09984, 32'hc2bfb932, 32'h42b22d48};
test_bias[2591:2591] = '{32'h42aaa607};
test_output[2591:2591] = '{32'hc6a31a2a};
test_input[20736:20743] = '{32'h40b104ec, 32'h41cdb763, 32'h41a7e3ae, 32'hc2470760, 32'h427f1820, 32'h426529e3, 32'hc2bd6524, 32'hc1cb3b52};
test_weights[20736:20743] = '{32'h42c51611, 32'hc2888422, 32'hc1a641d1, 32'hc289f2a2, 32'h41d1c31a, 32'hc1f5a179, 32'hc2b9cd9d, 32'hc1aa5656};
test_bias[2592:2592] = '{32'h4251237c};
test_output[2592:2592] = '{32'h462d463f};
test_input[20744:20751] = '{32'hc2c1cc0e, 32'h421b4ecf, 32'hc2a4d959, 32'h42c7db4b, 32'hc1ea62e6, 32'hc25413aa, 32'hc21a0e84, 32'hc258484d};
test_weights[20744:20751] = '{32'h418a9227, 32'h41442026, 32'hc208cf36, 32'h4260f7fb, 32'hc1f0f690, 32'h413e5498, 32'h427f25ea, 32'h421de196};
test_bias[2593:2593] = '{32'h4168e956};
test_output[2593:2593] = '{32'h4536043b};
test_input[20752:20759] = '{32'h41097856, 32'hc254af7f, 32'h40baee83, 32'h429a8b41, 32'h41c7f9e5, 32'h42a3cdbd, 32'h4250ee77, 32'h42b3ea5e};
test_weights[20752:20759] = '{32'h41c4dda2, 32'h417548b3, 32'hc280d06e, 32'h40f0e5e7, 32'hc22ff4b1, 32'h41b13bb5, 32'hc15569e8, 32'h42a2eb26};
test_bias[2594:2594] = '{32'h41260fc9};
test_output[2594:2594] = '{32'h45d971b3};
test_input[20760:20767] = '{32'hc1bab52f, 32'hc2abb0dc, 32'h41f3626b, 32'hc1f6d239, 32'hc2c114f6, 32'h4289398d, 32'hc1a5afa0, 32'h4233c3fd};
test_weights[20760:20767] = '{32'hc2a2dd00, 32'hc2291d1e, 32'h4208cfe0, 32'h42b04e55, 32'hbfe8f4c9, 32'h42903483, 32'hc130d215, 32'h428fb9c3};
test_bias[2595:2595] = '{32'hc2b4c48e};
test_output[2595:2595] = '{32'h4640d69a};
test_input[20768:20775] = '{32'h428a4014, 32'h424962d4, 32'h42baed83, 32'hc2940835, 32'hc257ae71, 32'h420b2461, 32'hc217beb8, 32'h420d359b};
test_weights[20768:20775] = '{32'hc1aa7165, 32'h426e4670, 32'h41f82a39, 32'h413db3b2, 32'hc29f285b, 32'h4288e727, 32'hc28d2123, 32'hc18895f8};
test_bias[2596:2596] = '{32'h427b36c4};
test_output[2596:2596] = '{32'h464114ac};
test_input[20776:20783] = '{32'h4200c4fd, 32'hc1ec4efd, 32'hc035063e, 32'hc28c72e0, 32'h40aea1d9, 32'hc2c70d0f, 32'h427d80f2, 32'hc291b5a3};
test_weights[20776:20783] = '{32'hc11276f8, 32'h420a0690, 32'h42889032, 32'hc28e1c75, 32'h42a8afbf, 32'hc1d09a8d, 32'h41ebefcd, 32'hc227b54e};
test_bias[2597:2597] = '{32'h42541713};
test_output[2597:2597] = '{32'h4633eb90};
test_input[20784:20791] = '{32'hc03613e1, 32'h4169f1ec, 32'hc241a518, 32'hc2c00e03, 32'hc277921e, 32'h42941b3e, 32'h42a8f511, 32'hc2988469};
test_weights[20784:20791] = '{32'hc259d0b9, 32'hbffcea0f, 32'h409f3da3, 32'hc2628fec, 32'h4279413d, 32'h4202f927, 32'hc2220861, 32'hc262cd14};
test_bias[2598:2598] = '{32'h411e7364};
test_output[2598:2598] = '{32'h45961ede};
test_input[20792:20799] = '{32'h42984987, 32'h42c28160, 32'h41ae422b, 32'h4225d0cb, 32'hc2755007, 32'h428713b0, 32'hc0528c19, 32'h419ed35f};
test_weights[20792:20799] = '{32'h42bb7e45, 32'hc2225919, 32'hc2b47310, 32'h41a084f8, 32'h42a8cbfe, 32'hc298a9cb, 32'h4108cb63, 32'hc10bce92};
test_bias[2599:2599] = '{32'hc1c68bfa};
test_output[2599:2599] = '{32'hc604d10e};
test_input[20800:20807] = '{32'hc2817503, 32'h42b0fb7e, 32'hc24b854c, 32'h3fbd8780, 32'h42806f53, 32'hc2610e59, 32'h429b27d1, 32'hc2c370ad};
test_weights[20800:20807] = '{32'h427672c5, 32'h4283cb90, 32'h42940e64, 32'h42918902, 32'hc236fe76, 32'hc2785a54, 32'hc2af46fe, 32'hc1e89afd};
test_bias[2600:2600] = '{32'hc28ba5d2};
test_output[2600:2600] = '{32'hc5a53b2c};
test_input[20808:20815] = '{32'h40f681a9, 32'h42bbb963, 32'h426cfcb2, 32'hc2a38cda, 32'hc1ac3bea, 32'hc1f73139, 32'hc24648bd, 32'hc2c236a7};
test_weights[20808:20815] = '{32'hc23a2f7b, 32'hc1da722c, 32'hc2b96354, 32'hc2aa9960, 32'hc2576af1, 32'h4253e914, 32'hc2a26b9e, 32'h42476500};
test_bias[2601:2601] = '{32'h42c0a736};
test_output[2601:2601] = '{32'hc524a207};
test_input[20816:20823] = '{32'h4101aa91, 32'h42b5634d, 32'h408833f3, 32'hc2493829, 32'h4118aa00, 32'hc284036b, 32'hc1a7704c, 32'hc00afed1};
test_weights[20816:20823] = '{32'hc297eee4, 32'h428db577, 32'hc1c65cf3, 32'hc29ba24b, 32'h421ec590, 32'hc28a4c01, 32'hc1ce66e5, 32'h427030cb};
test_bias[2602:2602] = '{32'h428e8891};
test_output[2602:2602] = '{32'h466b0d2f};
test_input[20824:20831] = '{32'h4234659b, 32'h42a43396, 32'h42c294a7, 32'hc1eaa101, 32'h4250cd9d, 32'h42216eb2, 32'h41d0027d, 32'hc20fa1cb};
test_weights[20824:20831] = '{32'h42ba95e7, 32'hc246d08d, 32'hc0fb93df, 32'h40db9867, 32'h408b7f34, 32'h422fcf2d, 32'hc28ab68a, 32'hc2760a1f};
test_bias[2603:2603] = '{32'hc25d70c6};
test_output[2603:2603] = '{32'h44bcfe9a};
test_input[20832:20839] = '{32'h42b5fd65, 32'hc2a2ecbc, 32'hc2a13fd9, 32'hc2200575, 32'h41844325, 32'hc2c71559, 32'h42c2ce91, 32'hc1e13cc7};
test_weights[20832:20839] = '{32'hc14a80e8, 32'h42593412, 32'h42165878, 32'hc208049c, 32'hc2ac9d0e, 32'h41da73a1, 32'h412a1a64, 32'h4280648b};
test_bias[2604:2604] = '{32'hc28b59f3};
test_output[2604:2604] = '{32'hc63f1f13};
test_input[20840:20847] = '{32'h424d0ba0, 32'hc2a4f128, 32'hc00a6836, 32'hc1b99d12, 32'h423ece12, 32'hc2423d63, 32'h420819e5, 32'hc0cd1a86};
test_weights[20840:20847] = '{32'hc2bad07c, 32'hc1f15b57, 32'hc27ec8c2, 32'hc20b0a5c, 32'hc1cb8f3f, 32'hc211ce88, 32'hc2be4c19, 32'hc26ffc40};
test_bias[2605:2605] = '{32'h42519382};
test_output[2605:2605] = '{32'hc5610005};
test_input[20848:20855] = '{32'hc2a39b19, 32'h41ad871b, 32'h41a150c3, 32'h4258e9a5, 32'hc2a4fbd5, 32'hc08c7104, 32'hc215b937, 32'h4290f9ab};
test_weights[20848:20855] = '{32'hc2005deb, 32'h4235bc40, 32'hc220d468, 32'h42c178b7, 32'h41ca9a80, 32'h42b09ee6, 32'hc1904517, 32'hc1fc0677};
test_bias[2606:2606] = '{32'hc032ce6f};
test_output[2606:2606] = '{32'h45775a93};
test_input[20856:20863] = '{32'h42a3658c, 32'hc26a26ad, 32'hc0a4981c, 32'h407aeac5, 32'hc1f7a600, 32'h40aa6b7a, 32'hc2964ef6, 32'hc2c112a6};
test_weights[20856:20863] = '{32'hc29a5888, 32'h422176b2, 32'h40e5b744, 32'hc121360d, 32'h42690b87, 32'h42432418, 32'h4299fc75, 32'hc2c4e9a0};
test_bias[2607:2607] = '{32'hc224a9c4};
test_output[2607:2607] = '{32'hc5ce9711};
test_input[20864:20871] = '{32'hc288ba0c, 32'h421b4e13, 32'h41d7939f, 32'hc1b38d74, 32'h40fff521, 32'hc16ffe2c, 32'hc1fa2850, 32'h427f6d5f};
test_weights[20864:20871] = '{32'hc2b096df, 32'hc2b8cb34, 32'hc222097d, 32'hc29eafea, 32'hc230a058, 32'h42c7b220, 32'hc2b34edd, 32'h4235ca59};
test_bias[2608:2608] = '{32'hc2bdd72a};
test_output[2608:2608] = '{32'h45d78d80};
test_input[20872:20879] = '{32'h41d112ef, 32'h41ceb33c, 32'hc15d388f, 32'h42c427bd, 32'h425d0f0d, 32'h4298a2b0, 32'h424a5345, 32'h4294f4e6};
test_weights[20872:20879] = '{32'hc196d636, 32'h42163e97, 32'h42ab06b1, 32'hbf8529e9, 32'h4249bb41, 32'hc1bf6a51, 32'h4245ed92, 32'hc1ad43c5};
test_bias[2609:2609] = '{32'h426a6d67};
test_output[2609:2609] = '{32'h4489dc9a};
test_input[20880:20887] = '{32'h421dcf7c, 32'hc2a23cf5, 32'h42ac55df, 32'hc1c7b70d, 32'h42702b41, 32'h426eec79, 32'hc2a1bb29, 32'h4252fd63};
test_weights[20880:20887] = '{32'hc2b5fe58, 32'h41c28252, 32'hc1bd8c05, 32'h420c8e8d, 32'hc29f0d15, 32'h42b5f702, 32'h42028114, 32'hc29c1218};
test_bias[2610:2610] = '{32'h42824180};
test_output[2610:2610] = '{32'hc662bbeb};
test_input[20888:20895] = '{32'hc26a978a, 32'hc29686a6, 32'h420e3516, 32'h4297a38a, 32'hc2983848, 32'hc2442b7c, 32'hc17f2631, 32'h42107f22};
test_weights[20888:20895] = '{32'hc2a36830, 32'hc2b0fde7, 32'hc207c01c, 32'h400ea492, 32'h4081d352, 32'hc28d77db, 32'hc2b0f419, 32'hc2a8b403};
test_bias[2611:2611] = '{32'hc2848adc};
test_output[2611:2611] = '{32'h46398179};
test_input[20896:20903] = '{32'h42bccc0a, 32'h429c070a, 32'h42495734, 32'h41e1d3e3, 32'hc2af6752, 32'hc2b61641, 32'h410fde52, 32'hc1bea75d};
test_weights[20896:20903] = '{32'h423a63d7, 32'h42c3cb6a, 32'hc2a82803, 32'h42baba0e, 32'hc236b866, 32'hc1ad4832, 32'hc24bee2c, 32'h4141a9a3};
test_bias[2612:2612] = '{32'h42ae3f4f};
test_output[2612:2612] = '{32'h467637ea};
test_input[20904:20911] = '{32'h41a38dd8, 32'hbfe26573, 32'h42a846b4, 32'hc2c02577, 32'hc2476987, 32'hc250ead8, 32'h42a1ebec, 32'h40bcd592};
test_weights[20904:20911] = '{32'hc2678a48, 32'hc235f30d, 32'h41cf35ad, 32'h4288afeb, 32'hc28b293e, 32'hc2bd0120, 32'h420c0062, 32'hc20f2c6f};
test_bias[2613:2613] = '{32'hc2b977c7};
test_output[2613:2613] = '{32'h45aa2500};
test_input[20912:20919] = '{32'h4212c961, 32'h40b97bf6, 32'h42428317, 32'h4289193a, 32'h427bed1a, 32'h4266f2b2, 32'h427b9d65, 32'hc28982af};
test_weights[20912:20919] = '{32'hc24a9f11, 32'h41b42a22, 32'h426c6e95, 32'hc23dade9, 32'h4242c1f0, 32'hc1420fc4, 32'h428794f8, 32'hc2987de5};
test_bias[2614:2614] = '{32'h41c77691};
test_output[2614:2614] = '{32'h4619049e};
test_input[20920:20927] = '{32'h4291fe85, 32'hc13b15ea, 32'h418766ac, 32'h429c15ce, 32'h408a8b2f, 32'hc187f936, 32'h429a0685, 32'h42c211c0};
test_weights[20920:20927] = '{32'h42233b0b, 32'h42580da3, 32'hc110f796, 32'hc2a3680c, 32'h42804520, 32'h4291460d, 32'hc2a10559, 32'hc2af8ca4};
test_bias[2615:2615] = '{32'h42631001};
test_output[2615:2615] = '{32'hc69ab025};
test_input[20928:20935] = '{32'h422b40f4, 32'h42719f05, 32'hc2c063fd, 32'h4282c61a, 32'hc1f13c6a, 32'hc27b2e8c, 32'h428a00cc, 32'hc0820b60};
test_weights[20928:20935] = '{32'h421a94c0, 32'hc2b8b7f2, 32'hc20fa2ed, 32'hc203494d, 32'h426477f8, 32'h42be7318, 32'hc226b3f3, 32'h424fa56e};
test_bias[2616:2616] = '{32'hc240f972};
test_output[2616:2616] = '{32'hc65234c0};
test_input[20936:20943] = '{32'h4115fe85, 32'h42b5c6e7, 32'hc28fc89c, 32'hc05a82da, 32'h400ed896, 32'hc2a35b8b, 32'hc2bd197c, 32'hc2552c30};
test_weights[20936:20943] = '{32'h42be1079, 32'h4235ff2b, 32'hc2b2f5de, 32'h41dc7d66, 32'hc07ee947, 32'h42936d85, 32'h42015192, 32'h42255900};
test_bias[2617:2617] = '{32'h42802371};
test_output[2617:2617] = '{32'h430b9e75};
test_input[20944:20951] = '{32'hc2399b20, 32'h411bcd69, 32'hc24daa0a, 32'hc101ef11, 32'hc215506e, 32'hc27e701f, 32'hc18dff96, 32'h4293d0ab};
test_weights[20944:20951] = '{32'h4287dd9f, 32'h42bc38a4, 32'h42354371, 32'h4196497e, 32'hbf58c07c, 32'h429f649b, 32'hc29e9d7e, 32'h42bc4bf5};
test_bias[2618:2618] = '{32'hbf0f0657};
test_output[2618:2618] = '{32'hc4add74d};
test_input[20952:20959] = '{32'h419a0bd5, 32'h429bb93e, 32'hc2691ecc, 32'hc2122833, 32'hc2c67005, 32'h4154781d, 32'hc14e9ead, 32'hc08d57c8};
test_weights[20952:20959] = '{32'hc268ec1b, 32'hc222aa03, 32'h42c0947f, 32'hc2b5e389, 32'hc2bed644, 32'h426cb3e6, 32'hc240f1b6, 32'hc200bf63};
test_bias[2619:2619] = '{32'hc2b03702};
test_output[2619:2619] = '{32'h45880dde};
test_input[20960:20967] = '{32'hc24ca3b2, 32'h419a1de9, 32'h4223d5e8, 32'h42b63695, 32'hc1c60358, 32'h4269cf10, 32'h41fcf2a8, 32'hc2a29268};
test_weights[20960:20967] = '{32'hc1cd0299, 32'h42969f17, 32'hc27b2ba4, 32'h429b4ed1, 32'h418bbb69, 32'hc270d950, 32'hc26e5f29, 32'h42a39faa};
test_bias[2620:2620] = '{32'hc06966b9};
test_output[2620:2620] = '{32'hc5a3494c};
test_input[20968:20975] = '{32'hc2b54566, 32'hc0adf033, 32'hc29213eb, 32'hc27d3f02, 32'h42ad6808, 32'hc1a2a5b5, 32'h42575a9f, 32'hc28e4a6a};
test_weights[20968:20975] = '{32'h4186966a, 32'h4270772e, 32'h428952b6, 32'hc2c584ce, 32'hc155084a, 32'h4273da18, 32'hc2912b3b, 32'hc2b336f2};
test_bias[2621:2621] = '{32'h4296defe};
test_output[2621:2621] = '{32'hc3e88392};
test_input[20976:20983] = '{32'hc19fb922, 32'hc1170dcd, 32'h42a65d83, 32'hc2c1c4b4, 32'hc289a483, 32'h42c2cbfb, 32'h424b76a7, 32'h42c4b7fd};
test_weights[20976:20983] = '{32'h415fdb73, 32'hc15d7556, 32'h42b0a6f1, 32'h3d2960c8, 32'h409ba6e2, 32'h41c0a8e5, 32'h42acbe98, 32'h42116e64};
test_bias[2622:2622] = '{32'h42b4e6a3};
test_output[2622:2622] = '{32'h4686e2af};
test_input[20984:20991] = '{32'hc2b9fd81, 32'h42bdc2bf, 32'h41a630ac, 32'hc2ada729, 32'hc299bd7f, 32'h42473dd9, 32'h428d45ae, 32'hc202666b};
test_weights[20984:20991] = '{32'h41c9338b, 32'hc2a77b97, 32'h40e2efd6, 32'hc165a890, 32'h4241b91e, 32'h423da29d, 32'h42918cfa, 32'h42b44da7};
test_bias[2623:2623] = '{32'hc2a3613b};
test_output[2623:2623] = '{32'hc5fe213a};
test_input[20992:20999] = '{32'h419e6ec3, 32'hc2a52ae3, 32'h418cd188, 32'h421c958f, 32'hc011de6f, 32'hc2991563, 32'h41d43799, 32'h428de388};
test_weights[20992:20999] = '{32'hc282e2ea, 32'h41d4a86a, 32'h4253f968, 32'hc1813101, 32'h42c61447, 32'hc2b0ad27, 32'hc2c03d78, 32'h42b603b0};
test_bias[2624:2624] = '{32'hc2b8d26d};
test_output[2624:2624] = '{32'h45dfbb57};
test_input[21000:21007] = '{32'hc2a733af, 32'hc2b0f0c9, 32'h4119271a, 32'h424de62d, 32'hc2a0a269, 32'hc26b16ce, 32'hc22f7c62, 32'hc21e771e};
test_weights[21000:21007] = '{32'h429ca44d, 32'h4277790d, 32'hc1107244, 32'hc1c6213f, 32'hc2b8c71b, 32'hc2742da1, 32'hc298f0a4, 32'h42a926b0};
test_bias[2625:2625] = '{32'h418539cf};
test_output[2625:2625] = '{32'hc5131605};
test_input[21008:21015] = '{32'h429859aa, 32'hc2649590, 32'h42bd88ed, 32'h42b46918, 32'hc2a0d603, 32'hc220cfa4, 32'hc22da109, 32'hc2468d89};
test_weights[21008:21015] = '{32'hc1d92ffe, 32'hc28b3726, 32'h424bebe3, 32'h425a7f1d, 32'h424c990a, 32'hc215fe01, 32'hc22c2d60, 32'hc25ec315};
test_bias[2626:2626] = '{32'h4114a163};
test_output[2626:2626] = '{32'h465622e6};
test_input[21016:21023] = '{32'hc2b6a803, 32'h41191de6, 32'h42af26c7, 32'h427f99f2, 32'hc29ce624, 32'h4285ee0a, 32'hc2c44fa1, 32'hc25c910f};
test_weights[21016:21023] = '{32'h409eee07, 32'hc294e22b, 32'hc23e5cc4, 32'hc2236d20, 32'hc28bdec3, 32'h428450cf, 32'hc2499a7b, 32'h42a3abb9};
test_bias[2627:2627] = '{32'hc22766ce};
test_output[2627:2627] = '{32'h4513cd99};
test_input[21024:21031] = '{32'hc2b06b4a, 32'h425c1879, 32'h4234098e, 32'h41985708, 32'h421a2519, 32'h429c617f, 32'h42bb156e, 32'hc2c18cf0};
test_weights[21024:21031] = '{32'hc244143f, 32'hc2994e84, 32'h42572e8f, 32'hc17c5606, 32'h41fffa07, 32'hc2949af3, 32'h420d28a3, 32'hc1ac494e};
test_bias[2628:2628] = '{32'h42531ae0};
test_output[2628:2628] = '{32'h454107d0};
test_input[21032:21039] = '{32'h42c467ef, 32'hc2245872, 32'hc27b7c95, 32'h429e24a0, 32'hc2b2fc0d, 32'hc282e3e3, 32'h42a64b63, 32'hc2834947};
test_weights[21032:21039] = '{32'hc1971ff2, 32'hc1430c33, 32'hc2368d44, 32'hc12a2ee7, 32'hc27fd771, 32'hc24ee7aa, 32'h424d78b9, 32'h4196e9f4};
test_bias[2629:2629] = '{32'h42061b6b};
test_output[2629:2629] = '{32'h4648c634};
test_input[21040:21047] = '{32'h42a87453, 32'hc1c39c26, 32'h41d21962, 32'hc1a8120c, 32'hc29a9edf, 32'h41ad0a58, 32'hc27027a8, 32'hc24a40fd};
test_weights[21040:21047] = '{32'hc28a282a, 32'hc0e0b4ec, 32'h418e019b, 32'hc1294746, 32'hc25a7bee, 32'hc1241fd9, 32'h420cdf30, 32'hc0373b33};
test_bias[2630:2630] = '{32'h429e6521};
test_output[2630:2630] = '{32'hc531fb9d};
test_input[21048:21055] = '{32'hc28e1ddb, 32'h429f0fca, 32'h42b89e62, 32'hc2bb1114, 32'hc25e1479, 32'hc1207d3d, 32'h42c1f70a, 32'h3f8bc871};
test_weights[21048:21055] = '{32'h42c49566, 32'h423f020e, 32'hc2b81a61, 32'hc2a82aec, 32'hc12adaa1, 32'hc1f9179d, 32'h42b6b79e, 32'hc18f395a};
test_bias[2631:2631] = '{32'h4235500f};
test_output[2631:2631] = '{32'h45ba9f0f};
test_input[21056:21063] = '{32'h4267d9a7, 32'h421a6fb4, 32'h4211f2f2, 32'h4176f0d3, 32'hc1869b03, 32'hc1e204ea, 32'h41814439, 32'hc1851f83};
test_weights[21056:21063] = '{32'hc26b97db, 32'hc2a6a221, 32'h42a7419e, 32'h423c4ca2, 32'h41d89c89, 32'h42984179, 32'h420b0fae, 32'h4293da51};
test_bias[2632:2632] = '{32'hc254452d};
test_output[2632:2632] = '{32'hc5c12506};
test_input[21064:21071] = '{32'hc1a02789, 32'hc2722f75, 32'h428e9986, 32'h429d202a, 32'hc25d0ab2, 32'hc21ade19, 32'h418fb166, 32'hc1fbb9de};
test_weights[21064:21071] = '{32'h40451e00, 32'h4256ed55, 32'h41d054d8, 32'h42250cfc, 32'h41829b20, 32'h4263fdec, 32'hc26df4b8, 32'h41c0aa1f};
test_bias[2633:2633] = '{32'h428e15bd};
test_output[2633:2633] = '{32'hc5408adb};
test_input[21072:21079] = '{32'h42812f04, 32'h42abaceb, 32'h42a26830, 32'hc291acdf, 32'hc2a25df5, 32'hc2253412, 32'hc09f28fa, 32'hc1eacbef};
test_weights[21072:21079] = '{32'h42c032cb, 32'h419cd08d, 32'hc04ebc53, 32'hc050308e, 32'h425ff764, 32'h418b2044, 32'hc28dc55c, 32'h4273d1f5};
test_bias[2634:2634] = '{32'hc29c83f2};
test_output[2634:2634] = '{32'h4487bc72};
test_input[21080:21087] = '{32'h42b892e3, 32'h4219ae6e, 32'hc20aa978, 32'h41268df5, 32'h4150fe19, 32'hc1bd5921, 32'h416e7cfc, 32'hc2435a40};
test_weights[21080:21087] = '{32'h429b56dc, 32'hc11db21d, 32'hc294d0f9, 32'h42aa4d2c, 32'hc22fb62e, 32'hc296c315, 32'hc2b4a9ef, 32'h4083f671};
test_bias[2635:2635] = '{32'hc1eb5715};
test_output[2635:2635] = '{32'h461a8074};
test_input[21088:21095] = '{32'h4283d06b, 32'hc27b1aac, 32'h42251315, 32'hc238dd6f, 32'h4094a79e, 32'h42771386, 32'hc1a38ee4, 32'h426e1a2c};
test_weights[21088:21095] = '{32'h41076daa, 32'h42923d79, 32'hc28260da, 32'hc253c2b1, 32'h427a7cf3, 32'hc220ddc3, 32'h41cafb82, 32'h419474b2};
test_bias[2636:2636] = '{32'h42ad14ab};
test_output[2636:2636] = '{32'hc5b525cd};
test_input[21096:21103] = '{32'hc2973571, 32'h42830e70, 32'hc21bc20b, 32'hc2b02328, 32'hc261c753, 32'hc281b635, 32'h420a34fe, 32'hc180d1bd};
test_weights[21096:21103] = '{32'hc2a19d75, 32'hbeb44809, 32'h41fa2769, 32'hc2bed940, 32'hc14b6e79, 32'h4065dcfd, 32'hc246a39c, 32'h42b65b87};
test_bias[2637:2637] = '{32'h4222bd58};
test_output[2637:2637] = '{32'h4625d7fa};
test_input[21104:21111] = '{32'h41c0c68c, 32'h41992090, 32'hc2b11880, 32'hc23a5ce7, 32'hc1a8218a, 32'h42bf94bc, 32'hc2713fd0, 32'hc191fa70};
test_weights[21104:21111] = '{32'h416cfd68, 32'h3fdf0d7c, 32'h42c55930, 32'h412bba93, 32'hc1cb54b9, 32'h4236fa8a, 32'hc1ba1d3f, 32'hc1c3e99b};
test_bias[2638:2638] = '{32'h41cdb4db};
test_output[2638:2638] = '{32'hc50076a0};
test_input[21112:21119] = '{32'hc29cf5c1, 32'h41b9f8f9, 32'hc2c547b5, 32'h424b2b52, 32'h42920b08, 32'hc0db1f9a, 32'h42454970, 32'hc153a069};
test_weights[21112:21119] = '{32'hc2682dde, 32'hc2811912, 32'hc19e8c91, 32'h41e50701, 32'h3f5c9501, 32'hc224338f, 32'h4295805b, 32'hc2c65b74};
test_bias[2639:2639] = '{32'h40df003f};
test_output[2639:2639] = '{32'h463895c9};
test_input[21120:21127] = '{32'h408bb1f7, 32'hc1aa9355, 32'hc0717a8b, 32'h429c2e31, 32'h40b75c80, 32'hc23fd33b, 32'h3f8e78ba, 32'h420292ce};
test_weights[21120:21127] = '{32'h42ab6571, 32'hc2a10e9a, 32'h41ba4bb6, 32'h42812cdf, 32'hc25a342d, 32'h41904fb3, 32'hc2484c4d, 32'h429a7b4d};
test_bias[2640:2640] = '{32'hc1bc60f9};
test_output[2640:2640] = '{32'h4601dd94};
test_input[21128:21135] = '{32'h42823a35, 32'hc2bb88b7, 32'hc298afbc, 32'hc2b22b1f, 32'h42aacc64, 32'hc1b622c5, 32'hc287f64b, 32'hc2b687c0};
test_weights[21128:21135] = '{32'hc263975b, 32'h4216da8e, 32'h42ae8e2f, 32'h424ca044, 32'h40ee005b, 32'h425019c1, 32'h427c93b7, 32'hc2119aa9};
test_bias[2641:2641] = '{32'hc1aca9dd};
test_output[2641:2641] = '{32'hc69c457e};
test_input[21136:21143] = '{32'hc1a07822, 32'h4206dd9a, 32'hc1286dfb, 32'hc2c00b1e, 32'hc1ec8adf, 32'h4048e2cd, 32'hc2038c38, 32'h42c0ac4c};
test_weights[21136:21143] = '{32'hc200f915, 32'hc28ac8e5, 32'hc26cf056, 32'h429abc76, 32'h42214ac8, 32'hc24adbec, 32'h41b7c8cc, 32'h426802a6};
test_bias[2642:2642] = '{32'hc25a8646};
test_output[2642:2642] = '{32'hc59e818c};
test_input[21144:21151] = '{32'h40191eef, 32'hc212f990, 32'hc20747df, 32'h4261cffb, 32'hc265b01c, 32'h42247c06, 32'hc1980b06, 32'hc24282a2};
test_weights[21144:21151] = '{32'hc074efc6, 32'hc051915a, 32'hc23bce0f, 32'hc283a724, 32'h420bde11, 32'hc2996348, 32'hc29a08fe, 32'hc15afb51};
test_bias[2643:2643] = '{32'hc2592848};
test_output[2643:2643] = '{32'hc59f7d48};
test_input[21152:21159] = '{32'hc24b19f7, 32'hc210c2f5, 32'hc03a5eaa, 32'h42bce7bd, 32'hc0b8ca24, 32'h40b9bd15, 32'h41be851f, 32'hc23bf542};
test_weights[21152:21159] = '{32'hc13a2122, 32'hc2116d7a, 32'h401af7de, 32'h42af857e, 32'hc1f25f71, 32'hc2c26d2e, 32'h3f5caefa, 32'h425956f2};
test_bias[2644:2644] = '{32'hc288cd1a};
test_output[2644:2644] = '{32'h45e0f238};
test_input[21160:21167] = '{32'h41ac085e, 32'h42b5efc1, 32'h422dc413, 32'hc2bcb5ac, 32'h40744a1d, 32'h420c5f8b, 32'hc2b262db, 32'hc0ad741f};
test_weights[21160:21167] = '{32'h420903ab, 32'h42c55c5b, 32'h4298362e, 32'hc252ef45, 32'hc1d04443, 32'hc2ae08b4, 32'hbff19c68, 32'hc25dde46};
test_bias[2645:2645] = '{32'h4258ee58};
test_output[2645:2645] = '{32'h46701575};
test_input[21168:21175] = '{32'hc1bc50f4, 32'hc2c604d6, 32'h42658a1d, 32'h412c307c, 32'h42260433, 32'h42725702, 32'hc02aa8d4, 32'hbfc3b253};
test_weights[21168:21175] = '{32'hc2b52071, 32'hc09bb569, 32'h424eff4f, 32'h41fb9edb, 32'hc24b69ae, 32'hc1bf5cb6, 32'h42b64eb8, 32'h4129bbc4};
test_bias[2646:2646] = '{32'h42c7b4d6};
test_output[2646:2646] = '{32'h4509a728};
test_input[21176:21183] = '{32'h42b53d57, 32'hc14d27df, 32'h427cc243, 32'h423a1812, 32'h42bb0717, 32'h41927251, 32'hc2b66eb8, 32'hc2ad0e64};
test_weights[21176:21183] = '{32'hc1e08aad, 32'h42c23d49, 32'hc1bb6550, 32'hc2ae9913, 32'h42b3041a, 32'hc2a4c18e, 32'hc27f93ec, 32'hc29b2520};
test_bias[2647:2647] = '{32'h41cfea90};
test_output[2647:2647] = '{32'h461dc8e5};
test_input[21184:21191] = '{32'hc297495d, 32'hbff57168, 32'hc299ceae, 32'h42c1453b, 32'h42ade0bd, 32'hc2366286, 32'h42bd603b, 32'hc221b7bb};
test_weights[21184:21191] = '{32'hc27522bb, 32'h427277ae, 32'h42ad8c17, 32'hc1a6da32, 32'h429b487e, 32'h428c2082, 32'h4230b780, 32'h42878d00};
test_bias[2648:2648] = '{32'hc2c46e41};
test_output[2648:2648] = '{32'h4436c966};
test_input[21192:21199] = '{32'hc1d0a425, 32'h429d65ab, 32'hc21a7660, 32'h3f6b9c72, 32'h429cddd7, 32'h41526a7f, 32'hc2436c3d, 32'h4276b4f9};
test_weights[21192:21199] = '{32'h40970b3e, 32'hc186e647, 32'hc2955eb7, 32'hc282569e, 32'hc2853b29, 32'h4087f6a4, 32'hc27c882e, 32'hc1d480e4};
test_bias[2649:2649] = '{32'h40c1ebbf};
test_output[2649:2649] = '{32'hc5126f8d};
test_input[21200:21207] = '{32'hc29d00e9, 32'h4149dea8, 32'hc1ac648b, 32'h422a847b, 32'h4280df16, 32'h4196ed02, 32'hc252d063, 32'hc2a62a20};
test_weights[21200:21207] = '{32'h42c1e781, 32'h41a5b373, 32'hc279f98c, 32'hc1f9dc33, 32'h3f2fb28a, 32'hc19cc5b0, 32'hc1d2f9db, 32'hc0b1b261};
test_bias[2650:2650] = '{32'h40d5ae3e};
test_output[2650:2650] = '{32'hc5b54f02};
test_input[21208:21215] = '{32'h4284f69c, 32'h406b5dc7, 32'hc2809bb5, 32'hc2aebd0d, 32'hc286f5a6, 32'h42a01703, 32'hc172065c, 32'h4249b15a};
test_weights[21208:21215] = '{32'h428d42d5, 32'h429d0343, 32'h42af4bc0, 32'hc21ac848, 32'hc1b92dd5, 32'hc0475345, 32'h4199b0cd, 32'h4283d124};
test_bias[2651:2651] = '{32'h42aba68b};
test_output[2651:2651] = '{32'h45dfc209};
test_input[21216:21223] = '{32'hc24bd35a, 32'hc2b3780b, 32'hc24fe1ac, 32'hc1950f37, 32'hc1ff0177, 32'hc2a941ab, 32'hc2b69adf, 32'hc27e7fd0};
test_weights[21216:21223] = '{32'hc1d909a6, 32'hc24f8cb2, 32'hc2058d34, 32'h428316b4, 32'h4166978b, 32'hc185c95e, 32'hc27d0d19, 32'hc26e0521};
test_bias[2652:2652] = '{32'h416e98f2};
test_output[2652:2652] = '{32'h46857a90};
test_input[21224:21231] = '{32'hc1dc5265, 32'h421a01e6, 32'h42a5a6dc, 32'hc0287330, 32'h41ab1366, 32'h41fc6315, 32'hc2ac4a9f, 32'h4231b173};
test_weights[21224:21231] = '{32'hc1a77dbf, 32'h428bb3ad, 32'h42775990, 32'hc1eafd33, 32'h41f43320, 32'h4260a652, 32'hc1ecb095, 32'h41a68477};
test_bias[2653:2653] = '{32'h42ad15aa};
test_output[2653:2653] = '{32'h4661c63c};
test_input[21232:21239] = '{32'hc1c5465e, 32'h428630f5, 32'h403bbbed, 32'h41fffcc6, 32'hc1e86cc0, 32'hc0c0206a, 32'h42363bd6, 32'hc202f260};
test_weights[21232:21239] = '{32'h40da3d50, 32'hc207b333, 32'h4280d5ac, 32'h42422978, 32'hc2a760c7, 32'hc1aeb4f0, 32'hc2539d23, 32'hc10a545a};
test_bias[2654:2654] = '{32'hc28baf34};
test_output[2654:2654] = '{32'hc3a85816};
test_input[21240:21247] = '{32'hc22abb34, 32'hc2bd28fe, 32'h41d85120, 32'hc188d5c6, 32'h4281a3c8, 32'hc2a4ac29, 32'hc1c55c89, 32'hc1bd08ca};
test_weights[21240:21247] = '{32'h4288869c, 32'h406a0886, 32'h429f667a, 32'h428eba1a, 32'h4225d4aa, 32'hc2b76ca3, 32'h3f9e9d90, 32'hc25d95d8};
test_bias[2655:2655] = '{32'h42af3d59};
test_output[2655:2655] = '{32'h4610fdde};
test_input[21248:21255] = '{32'h4248be3d, 32'h4294bb96, 32'h40b1b3a5, 32'h419039d6, 32'h429482c1, 32'hbfd8897c, 32'hc29bee9e, 32'h4225d7c2};
test_weights[21248:21255] = '{32'hc2b01675, 32'h4250eabe, 32'hc1bc4ade, 32'h4240baac, 32'h4255cffa, 32'h42bdd811, 32'h417c85e7, 32'h42b8c9c3};
test_bias[2656:2656] = '{32'h42c6ed27};
test_output[2656:2656] = '{32'h45d1be19};
test_input[21256:21263] = '{32'h4221927b, 32'hc26cd30d, 32'hc17745ce, 32'h4202b005, 32'hc1b97f16, 32'h427354bb, 32'hc1ad9766, 32'h42207a84};
test_weights[21256:21263] = '{32'h428858e2, 32'hc1c7d0ca, 32'hc2addb73, 32'hc054e7ec, 32'h429ebbbc, 32'hc2660667, 32'hc239001e, 32'h42bcdd5a};
test_bias[2657:2657] = '{32'h4148b611};
test_output[2657:2657] = '{32'h459a2b9d};
test_input[21264:21271] = '{32'h419ac4b5, 32'h42a23584, 32'h429c9841, 32'h4176dd0a, 32'h420bb7e3, 32'h41f66eea, 32'hc208eb57, 32'h4250db14};
test_weights[21264:21271] = '{32'h4294c72a, 32'hc29dfb33, 32'hc15a51ec, 32'hc2a1ea4e, 32'h3fc20edc, 32'hc2a6998b, 32'hc2084ba1, 32'h41a19868};
test_bias[2658:2658] = '{32'h42826a4b};
test_output[2658:2658] = '{32'hc5eabce0};
test_input[21272:21279] = '{32'h41a9cae2, 32'h41632a43, 32'h426c7d8a, 32'hc2b7597d, 32'hc2bd3541, 32'hc2306ba1, 32'hc106ed9e, 32'hc2413704};
test_weights[21272:21279] = '{32'hc1b280ca, 32'hc19b5900, 32'hc1d127bf, 32'h4235b5ac, 32'hc2a5e284, 32'h423829f8, 32'hc155416e, 32'h4289bcd5};
test_bias[2659:2659] = '{32'hc27f1833};
test_output[2659:2659] = '{32'hc57517ef};
test_input[21280:21287] = '{32'h426c0f03, 32'h42801e57, 32'hc2c2f873, 32'hc21795df, 32'hc2aa70e6, 32'h42a87dbb, 32'hc0a940d5, 32'h4227786c};
test_weights[21280:21287] = '{32'h429cb73c, 32'h42b1c170, 32'hc2a92892, 32'h42025dd6, 32'h42210922, 32'h41ada517, 32'hc21e8998, 32'hc19ec039};
test_bias[2660:2660] = '{32'h41a0cc7a};
test_output[2660:2660] = '{32'h466c51df};
test_input[21288:21295] = '{32'h42322085, 32'hc246299c, 32'h426c83d1, 32'hc29df309, 32'h41564f60, 32'hc24bda01, 32'h423847f1, 32'h41f9a447};
test_weights[21288:21295] = '{32'hc28bff7d, 32'hc209855d, 32'h4033c08a, 32'h424797aa, 32'hc2a4962d, 32'h40c9352f, 32'h426fae2c, 32'h429af2d4};
test_bias[2661:2661] = '{32'hc2490aa0};
test_output[2661:2661] = '{32'hc4b96d25};
test_input[21296:21303] = '{32'h40d3610d, 32'h41abc52e, 32'h418dc9b5, 32'hc2be4c1b, 32'h427db943, 32'h428ce67e, 32'hbcde239b, 32'h417275ca};
test_weights[21296:21303] = '{32'hc2312981, 32'hc2804189, 32'h41772744, 32'hc206af10, 32'hc2576ca2, 32'hc132b1a0, 32'hc19704a4, 32'hc2c521aa};
test_bias[2662:2662] = '{32'h423aed61};
test_output[2662:2662] = '{32'hc57014e3};
test_input[21304:21311] = '{32'h40998214, 32'h3fa2f27d, 32'h4219d6db, 32'h42aa6472, 32'hbf8ef577, 32'h424887d7, 32'h41e191f0, 32'h4254ac5c};
test_weights[21304:21311] = '{32'hc22acbdb, 32'h41cb2089, 32'h4241cb8b, 32'hc22f8bf4, 32'hc143c466, 32'hc14f8fb8, 32'h4221dc84, 32'hc17feac7};
test_bias[2663:2663] = '{32'h4276ae75};
test_output[2663:2663] = '{32'hc511c9de};
test_input[21312:21319] = '{32'hc1af2f45, 32'hc2bc8e3a, 32'h42911dfa, 32'h42171201, 32'h42073439, 32'hc2a3298d, 32'hc1be528e, 32'hc266a864};
test_weights[21312:21319] = '{32'hc2861d52, 32'hc2bfe079, 32'hc2990b5b, 32'hc18f7df9, 32'hc29afcda, 32'h422af1c6, 32'h41b72afb, 32'hc1d653ce};
test_bias[2664:2664] = '{32'h41d0d77e};
test_output[2664:2664] = '{32'hc44700e3};
test_input[21320:21327] = '{32'hc27f5ba8, 32'h423ae0ca, 32'hc2a5a902, 32'hc09dc8f8, 32'h411623b0, 32'h408b151f, 32'hc25dfac7, 32'hc2a13ab9};
test_weights[21320:21327] = '{32'h42be0c5d, 32'hc1c2750c, 32'h412f284f, 32'hc13dc4ae, 32'hc2322fdd, 32'h4255c2ba, 32'hc2a0c4d3, 32'hc11c2073};
test_bias[2665:2665] = '{32'hc237c1ec};
test_output[2665:2665] = '{32'hc53da541};
test_input[21328:21335] = '{32'hc1d9d87c, 32'hc2892ccd, 32'h429b0ab1, 32'hc21e500e, 32'h42830c71, 32'h424f9a1b, 32'h4236097d, 32'hc29747da};
test_weights[21328:21335] = '{32'hc2642b8a, 32'h41910993, 32'h41b79878, 32'h41a24d88, 32'hc1ee75bb, 32'hc2a025e6, 32'hc27c7697, 32'h41735ea0};
test_bias[2666:2666] = '{32'hc04d6040};
test_output[2666:2666] = '{32'hc60a449a};
test_input[21336:21343] = '{32'h42bda245, 32'h40e970cc, 32'hc040e24c, 32'h4264b96e, 32'hc1b32190, 32'hc2a4d46f, 32'h42794bc4, 32'h42560a22};
test_weights[21336:21343] = '{32'hc2937e19, 32'h41637e40, 32'h42a2ac90, 32'h428c0fec, 32'h42968c8b, 32'h42b16c81, 32'hc1d4bb5b, 32'hc264c997};
test_bias[2667:2667] = '{32'h42c346b9};
test_output[2667:2667] = '{32'hc682d493};
test_input[21344:21351] = '{32'hc220572b, 32'h40da0b99, 32'hc244a21d, 32'h42b41572, 32'h42bb9b0b, 32'h41feda2d, 32'h4278d4a5, 32'hc2c2f6ef};
test_weights[21344:21351] = '{32'hc28ec0b6, 32'h42867d3f, 32'h4280ffa5, 32'h41d10fcb, 32'h42a99003, 32'h41abfae4, 32'h41474ff7, 32'hc1c67590};
test_bias[2668:2668] = '{32'h42088be1};
test_output[2668:2668] = '{32'h46607a5e};
test_input[21352:21359] = '{32'h405b8058, 32'h429793e9, 32'h42656c81, 32'hc15903df, 32'h42142374, 32'h41c37447, 32'hc2a8dfed, 32'h42a488e5};
test_weights[21352:21359] = '{32'h4296cb98, 32'hc213447f, 32'hc1e2a6ec, 32'hc29df00c, 32'h41730a04, 32'h41d5e534, 32'hbfe6297f, 32'hc1e81ec7};
test_bias[2669:2669] = '{32'hc1f5d2e3};
test_output[2669:2669] = '{32'hc5813db6};
test_input[21360:21367] = '{32'hc2bb3ff9, 32'h42b0d665, 32'h429ef656, 32'h41aced6e, 32'h41c50676, 32'hc28efc49, 32'h429f7a34, 32'h42c351e3};
test_weights[21360:21367] = '{32'hbfd0682d, 32'h4289ce49, 32'hc2b58e7c, 32'hc207d3dc, 32'h41ba5dc5, 32'h4216f665, 32'h3feaeccf, 32'hc2ba5595};
test_bias[2670:2670] = '{32'hc1ba43c5};
test_output[2670:2670] = '{32'hc6481206};
test_input[21368:21375] = '{32'h428eab77, 32'hc2a449b1, 32'hc2b97637, 32'h422a7301, 32'hc2277569, 32'hc29514d9, 32'h42af5663, 32'hc1f2d721};
test_weights[21368:21375] = '{32'h42b4201a, 32'hc19eaf3b, 32'h4186a510, 32'h41a5f798, 32'hc216436d, 32'h426d20ff, 32'hc2bb26f6, 32'h42c00d1d};
test_bias[2671:2671] = '{32'h420cd363};
test_output[2671:2671] = '{32'hc5ccc280};
test_input[21376:21383] = '{32'h41d945cc, 32'hc28466d1, 32'hc0155fbd, 32'hc287b969, 32'h41e649d3, 32'hc2ad6e00, 32'hc2bd4549, 32'hc2550100};
test_weights[21376:21383] = '{32'h42c644c0, 32'hc2226946, 32'hc157a3cd, 32'hc0384816, 32'h40ea07ed, 32'h42b7c508, 32'hc1aa553a, 32'h42b09534};
test_bias[2672:2672] = '{32'hc299122e};
test_output[2672:2672] = '{32'hc5998a15};
test_input[21384:21391] = '{32'hc19e4290, 32'hc287435f, 32'hc167380d, 32'hc1bd971a, 32'hc1d4d7fb, 32'hc2bc2060, 32'hc287ef4d, 32'h420ad7e9};
test_weights[21384:21391] = '{32'h41565d98, 32'hc2985e54, 32'h41a04fff, 32'h411dba17, 32'hc221c6b8, 32'h42631313, 32'h4261ae25, 32'h42820f2f};
test_bias[2673:2673] = '{32'hc1c309a6};
test_output[2673:2673] = '{32'hc4bbaf01};
test_input[21392:21399] = '{32'hc22c14a2, 32'h4298a8b0, 32'hc125b95f, 32'hc233f449, 32'h41251ec9, 32'h41776cf5, 32'hc2a84a1f, 32'h420b2314};
test_weights[21392:21399] = '{32'hc20e9812, 32'h41829cb9, 32'hc146e21f, 32'h42c4e3f0, 32'h429b7e66, 32'h429e871c, 32'h424b2fea, 32'h424fd2f4};
test_bias[2674:2674] = '{32'h40bf8b69};
test_output[2674:2674] = '{32'hc4f42a03};
test_input[21400:21407] = '{32'hc28168c2, 32'h42c0a6f9, 32'h42c4f501, 32'h423856bc, 32'hc2c00fd9, 32'h429ff419, 32'hc2bd9af4, 32'h42a7390b};
test_weights[21400:21407] = '{32'hc002d359, 32'h4226f358, 32'hc1b20e76, 32'hc1657490, 32'hc2a3406a, 32'h4299368d, 32'hc2866e48, 32'hc29359f8};
test_bias[2675:2675] = '{32'hc1c2991f};
test_output[2675:2675] = '{32'h46717426};
test_input[21408:21415] = '{32'hc1b7a703, 32'hbf930f73, 32'h426208d9, 32'hc18a9b31, 32'hc084785a, 32'h4239b1e6, 32'h41a4c064, 32'h42886947};
test_weights[21408:21415] = '{32'h4291245c, 32'hc2b9a9d9, 32'hc2baf3e6, 32'hc283de20, 32'hc1bf58a9, 32'hc263df85, 32'h4126398f, 32'h4210cd7a};
test_bias[2676:2676] = '{32'hc1d9b576};
test_output[2676:2676] = '{32'hc5aea840};
test_input[21416:21423] = '{32'hbf918ffc, 32'h415c9cfa, 32'h4231f297, 32'hc12039e9, 32'h4276a8d1, 32'hc1a3e599, 32'hc284a8c4, 32'h410563fa};
test_weights[21416:21423] = '{32'h4297ef76, 32'h41f56f0e, 32'h40ac86ae, 32'h41f8257e, 32'hbfa5f741, 32'h42b97cd7, 32'hc2848ac6, 32'h42014320};
test_bias[2677:2677] = '{32'hc1d64c8e};
test_output[2677:2677] = '{32'h4536c335};
test_input[21424:21431] = '{32'hc1bc0cd9, 32'hc2898493, 32'hc27b9149, 32'hc28221ec, 32'hc1211bc6, 32'hc23b0d5c, 32'h425346b1, 32'hc2c55258};
test_weights[21424:21431] = '{32'hc1e0e433, 32'h423eee13, 32'h429b1daf, 32'h420ade7b, 32'h42b7fb59, 32'hc14da9d8, 32'hc2820b9e, 32'hc2943604};
test_bias[2678:2678] = '{32'hc298a310};
test_output[2678:2678] = '{32'hc5c45486};
test_input[21432:21439] = '{32'h42546be6, 32'h424656d1, 32'hc24ebb3a, 32'hc03389f4, 32'h4165651a, 32'h42be024e, 32'hc2901459, 32'hc24d53fe};
test_weights[21432:21439] = '{32'h41e72e12, 32'h426dba3a, 32'h429333a1, 32'hc270d803, 32'hc24b7579, 32'hc1912b49, 32'hc29c6f09, 32'hc1553c4c};
test_bias[2679:2679] = '{32'hc10f3c62};
test_output[2679:2679] = '{32'h4592f999};
test_input[21440:21447] = '{32'hc25aa901, 32'h423fc319, 32'h4216d7e2, 32'hc2a7c793, 32'h425e9d08, 32'h4203dfe9, 32'hc08b5f59, 32'h423d0209};
test_weights[21440:21447] = '{32'hc07971e5, 32'hc26a2977, 32'h42157e09, 32'hc2aecfa3, 32'h4217ec79, 32'h422fad5f, 32'hc2baf8c3, 32'hc248ea44};
test_bias[2680:2680] = '{32'h42c18d07};
test_output[2680:2680] = '{32'h45f5054b};
test_input[21448:21455] = '{32'hc16d061a, 32'hc23ebf3f, 32'h419072d5, 32'hc0c2b003, 32'hc2c5d03e, 32'h426fa2ea, 32'h4277e6c5, 32'hc2aba917};
test_weights[21448:21455] = '{32'hc1ebeb24, 32'h429b7923, 32'h41d52ddd, 32'h425c2e23, 32'hc132fd75, 32'hc2c11509, 32'hc24b2936, 32'h424a3d04};
test_bias[2681:2681] = '{32'h418ee6a0};
test_output[2681:2681] = '{32'hc66e9a2e};
test_input[21456:21463] = '{32'hc11b4c0b, 32'hc1eab68a, 32'hc212520d, 32'h41a07326, 32'hc2c0c530, 32'h42c1ff7d, 32'h42c2d75f, 32'h4252b56e};
test_weights[21456:21463] = '{32'hc21e5a37, 32'hc28f1c72, 32'h41d67690, 32'hc0a95ab1, 32'hc264e032, 32'h41cad4e7, 32'h426d00e3, 32'h4221d31e};
test_bias[2682:2682] = '{32'hc28a6780};
test_output[2682:2682] = '{32'h46866ac2};
test_input[21464:21471] = '{32'hc286a9f2, 32'h427af22a, 32'hc298daab, 32'h3f5cba2f, 32'hc29e6d63, 32'hc162a461, 32'h41d890e2, 32'hc27828c4};
test_weights[21464:21471] = '{32'h41d7c8c4, 32'h41e4b698, 32'hc2568ade, 32'hc2b10965, 32'h41a00c1f, 32'hc197e420, 32'h42b96b90, 32'hc08b2686};
test_bias[2683:2683] = '{32'h42b5cb08};
test_output[2683:2683] = '{32'h45ad977d};
test_input[21472:21479] = '{32'hc285e20e, 32'hc2c53146, 32'h41f940ba, 32'hc0d313eb, 32'h421e7046, 32'h42689575, 32'hc2b4e0ea, 32'h41b00303};
test_weights[21472:21479] = '{32'hc2b106c7, 32'h4083dabd, 32'h427b5da5, 32'hc2a89583, 32'hbf193a83, 32'h425c833e, 32'h429b2d55, 32'h41a57850};
test_bias[2684:2684] = '{32'h428d25ba};
test_output[2684:2684] = '{32'h459399f9};
test_input[21480:21487] = '{32'h42b8384d, 32'h42302f56, 32'hc21f8369, 32'hc0e63d34, 32'h42b812c6, 32'h4218916c, 32'hc1b0da08, 32'hc27fda4d};
test_weights[21480:21487] = '{32'h426c22ba, 32'hc2b66026, 32'hc164ff7c, 32'hc298f2f0, 32'hc18d8e91, 32'h427c6258, 32'hc2bf39d3, 32'h418a9da4};
test_bias[2685:2685] = '{32'hc27331f3};
test_output[2685:2685] = '{32'h45854604};
test_input[21488:21495] = '{32'h42c72535, 32'h420311bc, 32'h41824d8d, 32'h426a5fab, 32'hc2bc604e, 32'hc19d9d98, 32'hc1d2b6dc, 32'hc1635f94};
test_weights[21488:21495] = '{32'hc1f5b206, 32'hc2923e28, 32'h42ad079f, 32'hc2a07a78, 32'h41a99967, 32'h42b4de8e, 32'h42a3bc0e, 32'hc2857740};
test_bias[2686:2686] = '{32'hc1fa1fde};
test_output[2686:2686] = '{32'hc65710c0};
test_input[21496:21503] = '{32'hc08e9db1, 32'h42809344, 32'hc1cb4c9c, 32'hc258287f, 32'h40e731df, 32'h41f55e1a, 32'h42a9c919, 32'h40d0b75e};
test_weights[21496:21503] = '{32'h3f87148e, 32'hc2aa6675, 32'h40f09206, 32'h42c12029, 32'hc1998f1e, 32'hc1788273, 32'hc2156535, 32'hc265d4a7};
test_bias[2687:2687] = '{32'hc265496d};
test_output[2687:2687] = '{32'hc66c143b};
test_input[21504:21511] = '{32'h42b8621e, 32'h421f13f3, 32'hc1a50175, 32'h42b76217, 32'h41388129, 32'hc26c4dbb, 32'hc0b5504c, 32'hc10f9f5e};
test_weights[21504:21511] = '{32'hc058585a, 32'hc1d6193e, 32'h421464dc, 32'hc295baab, 32'h40846edd, 32'hc23aa0a0, 32'h42587758, 32'h42438b3e};
test_bias[2688:2688] = '{32'h41931343};
test_output[2688:2688] = '{32'hc5d8852b};
test_input[21512:21519] = '{32'hc29aabfe, 32'h42a4a830, 32'hc04a2f38, 32'hc0cb28d5, 32'hc12bed97, 32'hc285b6ee, 32'hc22a4188, 32'hc1edc7d9};
test_weights[21512:21519] = '{32'hc2b538fb, 32'hc27744f3, 32'hc22173b3, 32'hc23d8c84, 32'h40fe4faa, 32'h4251c01e, 32'h3fcc94fe, 32'h426747d7};
test_bias[2689:2689] = '{32'h42919950};
test_output[2689:2689] = '{32'hc538e7ce};
test_input[21520:21527] = '{32'h419d01fb, 32'hc2409aa6, 32'h4285deae, 32'hc2a7cfbd, 32'h426ac06d, 32'h42694356, 32'h42bc9de3, 32'hc23215ad};
test_weights[21520:21527] = '{32'hc254f2cd, 32'h425a7b86, 32'hc2370a17, 32'hc21426e0, 32'hc29fdc4b, 32'hc2657681, 32'hc21ad451, 32'hbf1bbbad};
test_bias[2690:2690] = '{32'h3fc5a9ea};
test_output[2690:2690] = '{32'hc66ee0ac};
test_input[21528:21535] = '{32'hc1d268db, 32'hc203397f, 32'hc11013fe, 32'h426b3603, 32'hc2156cc3, 32'hc2934c3a, 32'hc1d7d674, 32'hc23f63ef};
test_weights[21528:21535] = '{32'h41bfc31c, 32'hc0f415e1, 32'h426c87e6, 32'h42a7edd0, 32'h417cd0b5, 32'h41b3a056, 32'h408a507c, 32'hc2a000ef};
test_bias[2691:2691] = '{32'h41bf3904};
test_output[2691:2691] = '{32'h45ac5f3f};
test_input[21536:21543] = '{32'hc21bd4db, 32'hc24d2212, 32'h420ab521, 32'h4282c9fa, 32'hc2848d1d, 32'h4210ffc7, 32'h42a506b5, 32'h42595b32};
test_weights[21536:21543] = '{32'h42250085, 32'hc22d8aa0, 32'hc2c52ea0, 32'hc2c5fabc, 32'hc22874c5, 32'hc27fc4c9, 32'h4244243f, 32'h41eda825};
test_bias[2692:2692] = '{32'h423943f3};
test_output[2692:2692] = '{32'hc54166c4};
test_input[21544:21551] = '{32'hc2964647, 32'h426e7b3b, 32'h429dbe93, 32'h423da3b5, 32'h427b8afe, 32'h42552199, 32'h42b3ce41, 32'h42485069};
test_weights[21544:21551] = '{32'h4282e419, 32'h4288c7f8, 32'hc0a8d0a5, 32'hc21f43eb, 32'hc290b6b1, 32'h42034841, 32'hc2a699bf, 32'h40bed8bb};
test_bias[2693:2693] = '{32'hc290aadf};
test_output[2693:2693] = '{32'hc64e5ef7};
test_input[21552:21559] = '{32'hc2b57b30, 32'h425ff13d, 32'hc294cda1, 32'hc1b486bb, 32'h40a5e895, 32'hc21e89f9, 32'hc218e720, 32'h423f4024};
test_weights[21552:21559] = '{32'hc150b9c5, 32'h42a6b271, 32'hc23e0c0f, 32'hc2b24fb3, 32'h42aed965, 32'h41622a3b, 32'hc2c5e310, 32'hc2b7bd22};
test_bias[2694:2694] = '{32'h427077f3};
test_output[2694:2694] = '{32'h4627ceb7};
test_input[21560:21567] = '{32'h428683b1, 32'hc1f262d0, 32'hc1634165, 32'h420cf775, 32'hc2402986, 32'h41784e1a, 32'hc238ce55, 32'h4278bbfc};
test_weights[21560:21567] = '{32'h427a0181, 32'hc26fe77a, 32'hc283192d, 32'h41d213d5, 32'hc29d9ec9, 32'h429e0864, 32'hc2844bc9, 32'h421f1929};
test_bias[2695:2695] = '{32'h42aa2e2a};
test_output[2695:2695] = '{32'h46909066};
test_input[21568:21575] = '{32'hc2c13954, 32'h423e0f65, 32'h426e4502, 32'hc2c4c4e0, 32'h4175fb7b, 32'hc263de6c, 32'h419772b0, 32'hc2a115a6};
test_weights[21568:21575] = '{32'hc2c1abc8, 32'hc185fd5d, 32'h42297616, 32'h422ba3e8, 32'hc1aabe9d, 32'hbd9f5cca, 32'hc2baca24, 32'h42c2576f};
test_bias[2696:2696] = '{32'hc2b56e63};
test_output[2696:2696] = '{32'hc544b437};
test_input[21576:21583] = '{32'h42b6c78a, 32'hbf8632d6, 32'h421ea921, 32'h4060bc3e, 32'h40bb3fac, 32'h42346af0, 32'h42b8ba76, 32'hc29dddc6};
test_weights[21576:21583] = '{32'h429107e2, 32'hc1b61c6c, 32'h42804d0c, 32'hbfb30270, 32'h4237d078, 32'h429e5469, 32'h41399462, 32'h42506284};
test_bias[2697:2697] = '{32'hc116277c};
test_output[2697:2697] = '{32'h461bf030};
test_input[21584:21591] = '{32'h3fed803b, 32'h42c01114, 32'h4204c222, 32'h41200105, 32'h422a6719, 32'h427bdc57, 32'h428b2c9a, 32'hc24d736e};
test_weights[21584:21591] = '{32'hc29ffd4a, 32'hc2be6ef9, 32'hc098f841, 32'h41106853, 32'hc19c6a2a, 32'hc1241961, 32'h427b3d67, 32'hc21d59cc};
test_bias[2698:2698] = '{32'h42259746};
test_output[2698:2698] = '{32'hc589b6e7};
test_input[21592:21599] = '{32'h41ffbe0f, 32'hc27139ff, 32'hc1190f3d, 32'h42b0371f, 32'hc230e157, 32'hc218d431, 32'h41c35738, 32'h425711b6};
test_weights[21592:21599] = '{32'hc2281d5a, 32'h426d07d8, 32'h420bd67c, 32'hc2837e32, 32'h42931d5c, 32'h41effbe8, 32'h42af2170, 32'h4119965b};
test_bias[2699:2699] = '{32'h41aa26c9};
test_output[2699:2699] = '{32'hc6477ede};
test_input[21600:21607] = '{32'h429c49e8, 32'hbf22c282, 32'hc2626ee0, 32'hc280bcac, 32'hc1407024, 32'hc191b430, 32'h4234014e, 32'hc1f74db3};
test_weights[21600:21607] = '{32'h42bbb9fb, 32'hc1f845ff, 32'hc281b09f, 32'hc153d13b, 32'h425771cc, 32'h428d2c18, 32'h422cd6d0, 32'h42bdc710};
test_bias[2700:2700] = '{32'hc147cc92};
test_output[2700:2700] = '{32'h460bbb62};
test_input[21608:21615] = '{32'hc1750068, 32'hc1f78068, 32'h412a5130, 32'hc20554d8, 32'hc1a53287, 32'h4215be61, 32'h428d9988, 32'hc1a5d842};
test_weights[21608:21615] = '{32'h42403a54, 32'h42219260, 32'hc19fc88b, 32'hc12288ba, 32'h42a4b0e7, 32'hc1a72fec, 32'hc280bf59, 32'h4288574a};
test_bias[2701:2701] = '{32'h4172e4a1};
test_output[2701:2701] = '{32'hc620e7f1};
test_input[21616:21623] = '{32'hc13c40d6, 32'hc190162d, 32'h42686f01, 32'hc2c6aeb4, 32'h4290483c, 32'h429b60bf, 32'hc2c55ace, 32'h41987284};
test_weights[21616:21623] = '{32'h422bfeb3, 32'h42c25134, 32'h400212d9, 32'h4295ad34, 32'h42771ece, 32'h41a366a4, 32'h41df18a0, 32'hc249e0c6};
test_bias[2702:2702] = '{32'h429ea1dc};
test_output[2702:2702] = '{32'hc5dfd672};
test_input[21624:21631] = '{32'h42b7485c, 32'hc29fc0ce, 32'hc1aeeef6, 32'hc198d562, 32'hc2c10f97, 32'hc2c25c6e, 32'hc18b10ec, 32'h4204f2dc};
test_weights[21624:21631] = '{32'hc2305ce8, 32'hc26cddef, 32'h42a07c06, 32'h425dff42, 32'hc2bd73dc, 32'hc1f22c62, 32'hc1a3dc2d, 32'hc26af506};
test_bias[2703:2703] = '{32'hc20d5953};
test_output[2703:2703] = '{32'h46022318};
test_input[21632:21639] = '{32'hc2875882, 32'hc15ac475, 32'hc202af62, 32'h427d9947, 32'h41b34881, 32'hc1654e1e, 32'hc29a7a18, 32'h42af218c};
test_weights[21632:21639] = '{32'hc2b7e8f2, 32'hc23f6695, 32'h42335854, 32'h42997010, 32'h4203e34c, 32'hc2c466e9, 32'h42c12269, 32'hc09987e3};
test_bias[2704:2704] = '{32'hc23df0e3};
test_output[2704:2704] = '{32'h458c8173};
test_input[21640:21647] = '{32'hc0b6b3e3, 32'h422d4cc5, 32'hc2a0eb48, 32'h42be5755, 32'h42b747ea, 32'h421b74b7, 32'h428a13e7, 32'h42ad2cd9};
test_weights[21640:21647] = '{32'h42b018fd, 32'hc2a335ea, 32'hc26f7203, 32'hc2a606a0, 32'h4262a389, 32'hc2a3ddbb, 32'h42775af1, 32'hc0f70f2b};
test_bias[2705:2705] = '{32'h428ef3e7};
test_output[2705:2705] = '{32'hc4b43d03};
test_input[21648:21655] = '{32'hc2192f14, 32'hc2a57ebe, 32'hc2ad2bbc, 32'hc276fd00, 32'hc28e1d2f, 32'hc2adb814, 32'hc205f1d1, 32'h424bd5c6};
test_weights[21648:21655] = '{32'hc1aca15c, 32'hc179a5a0, 32'hc1cc8394, 32'hc20be89b, 32'hc29e347d, 32'h41d65274, 32'h4107536a, 32'hc22ac390};
test_bias[2706:2706] = '{32'hc20f8476};
test_output[2706:2706] = '{32'h45e3cf72};
test_input[21656:21663] = '{32'h4265e677, 32'h42380f56, 32'h429fd718, 32'h423ab2e1, 32'hc281f7d8, 32'h42400172, 32'h42006373, 32'h4294850d};
test_weights[21656:21663] = '{32'hc2544478, 32'h4215b008, 32'h42a28a94, 32'h4242fb05, 32'h4276ae56, 32'h42b9cc2f, 32'h42a8e771, 32'h42870fe1};
test_bias[2707:2707] = '{32'h40e19949};
test_output[2707:2707] = '{32'h46742a15};
test_input[21664:21671] = '{32'h4196a918, 32'hc28b7623, 32'h42626299, 32'hc19274be, 32'hc1f15f09, 32'h4157de70, 32'hc1e7f2cb, 32'h41c9ee76};
test_weights[21664:21671] = '{32'h4247f3b3, 32'h42b98839, 32'hc2189a05, 32'h42c3e556, 32'h40cdfdc2, 32'h42aaf611, 32'h4287e835, 32'h420e8260};
test_bias[2708:2708] = '{32'h417a4cdc};
test_output[2708:2708] = '{32'hc6159f10};
test_input[21672:21679] = '{32'h421304b0, 32'h420d27ac, 32'hc25023bd, 32'hc27e7c5e, 32'h42874201, 32'hc2726859, 32'hc2a3e2c3, 32'h410ee2cf};
test_weights[21672:21679] = '{32'h42b753ad, 32'hc1c810a9, 32'hc2916cb5, 32'hc2b012d1, 32'hc24099cb, 32'hbf9a444a, 32'h421f5a07, 32'hc2be13d2};
test_bias[2709:2709] = '{32'h4001e3a6};
test_output[2709:2709] = '{32'h458f05a7};
test_input[21680:21687] = '{32'hc23163ea, 32'h4045fefa, 32'hc14f80b2, 32'h4290771d, 32'h4212e53a, 32'hc28f9c01, 32'h4218bb55, 32'h41892187};
test_weights[21680:21687] = '{32'h41442b68, 32'hc1a11602, 32'h424e076f, 32'h4123df82, 32'hc104c3dc, 32'h42aa2036, 32'h41f343b1, 32'h423809d5};
test_bias[2710:2710] = '{32'h42a71217};
test_output[2710:2710] = '{32'hc5998c9b};
test_input[21688:21695] = '{32'h42b4ec09, 32'h423c5be3, 32'h4143a881, 32'hc287f156, 32'hc1e87a38, 32'h421cbb7e, 32'h42862641, 32'hc2c1e4ed};
test_weights[21688:21695] = '{32'hc2c4789e, 32'hc22aa537, 32'h419598dd, 32'hc2420522, 32'h428b43fb, 32'hc0f311a3, 32'h4213b53c, 32'h4230a277};
test_bias[2711:2711] = '{32'hc29bddf6};
test_output[2711:2711] = '{32'hc634d425};
test_input[21696:21703] = '{32'h428f911c, 32'hc2b5507e, 32'hc0ff4e4b, 32'hc2309787, 32'hc29a62c8, 32'h4284ac32, 32'h42906b46, 32'h42a744dc};
test_weights[21696:21703] = '{32'hc2b980c4, 32'h42968ee3, 32'hc2b8b67e, 32'h42008a94, 32'hc27f968e, 32'hc20e972d, 32'h42718cee, 32'h423b9b43};
test_bias[2712:2712] = '{32'hc1452c69};
test_output[2712:2712] = '{32'hc54fdf9a};
test_input[21704:21711] = '{32'h40acc1c0, 32'hc22897f5, 32'hc23bc082, 32'h40f512f7, 32'hc10a39cd, 32'h422276b2, 32'h42b11b20, 32'h42c34c70};
test_weights[21704:21711] = '{32'hc1e2c978, 32'hc261e8ed, 32'h42c78052, 32'hc24cbf26, 32'h424e0298, 32'h42853ef9, 32'h42a97bbb, 32'hc29e2b26};
test_bias[2713:2713] = '{32'h4258c9cf};
test_output[2713:2713] = '{32'hc43b79a7};
test_input[21712:21719] = '{32'h426a92f8, 32'hc29a0762, 32'hc2941408, 32'h429a374f, 32'h41a94bc2, 32'hc18f6eb9, 32'hc1fb5a6b, 32'h42816414};
test_weights[21712:21719] = '{32'h42216338, 32'hc011ab02, 32'hc2a35138, 32'hc299ff3b, 32'hc28b254e, 32'h42358f57, 32'h42bd2c24, 32'h42899cd8};
test_bias[2714:2714] = '{32'h427e7d76};
test_output[2714:2714] = '{32'h44ee688c};
test_input[21720:21727] = '{32'h426c6c66, 32'hc2ba4c3b, 32'h421beb87, 32'h424e8844, 32'h42239caa, 32'h40e83957, 32'hc27af7dc, 32'h427be6d5};
test_weights[21720:21727] = '{32'hc1b04fce, 32'h42b41d3d, 32'hc28a0ea9, 32'h4258623b, 32'h4291aa37, 32'h4299e8e2, 32'h416a564f, 32'h41d02eba};
test_bias[2715:2715] = '{32'h42575be5};
test_output[2715:2715] = '{32'hc5a4edae};
test_input[21728:21735] = '{32'hc27d338b, 32'h42bc85ab, 32'hc29e4aed, 32'hc2b82c5f, 32'h4235b8ec, 32'h429e5416, 32'h427009c8, 32'hc2ba2537};
test_weights[21728:21735] = '{32'hc2958463, 32'hc21e21d1, 32'hc28ba52c, 32'hc0c62704, 32'h42265cd2, 32'h42c0c0ea, 32'h4278f5ba, 32'hc2a76f9e};
test_bias[2716:2716] = '{32'hc28dbfef};
test_output[2716:2716] = '{32'h46db5a9c};
test_input[21736:21743] = '{32'hc1db37c0, 32'hc2c13ba9, 32'h424f285a, 32'hc2c3c7d8, 32'hc2816301, 32'h429f6174, 32'hc2714f66, 32'hc10d1d37};
test_weights[21736:21743] = '{32'hc255766b, 32'hc294b225, 32'hc27597b4, 32'h420cfc8a, 32'h41c53e6b, 32'hc2aea84d, 32'h42033f58, 32'h42542498};
test_bias[2717:2717] = '{32'h4293bd17};
test_output[2717:2717] = '{32'hc60b4095};
test_input[21744:21751] = '{32'h42903382, 32'h42a62f1e, 32'hc20cdf0e, 32'h417eadb0, 32'h42965ea0, 32'h42316ceb, 32'h423c15a6, 32'hc292f11e};
test_weights[21744:21751] = '{32'h4295edff, 32'hc2c44975, 32'h42b4230e, 32'hc2907dfd, 32'h41bb6d0a, 32'hc22bee60, 32'hc2c22981, 32'h4280fa86};
test_bias[2718:2718] = '{32'h42153f94};
test_output[2718:2718] = '{32'hc680c555};
test_input[21752:21759] = '{32'hc1dbcd5d, 32'h3f8600d1, 32'h420c8d34, 32'hc2930b3f, 32'h42b64736, 32'hc2191558, 32'h42b40082, 32'h41b9e529};
test_weights[21752:21759] = '{32'hc2a09968, 32'hc1fa8c12, 32'hc244e263, 32'h42605ce3, 32'hc1fdbb87, 32'h4033c759, 32'h42187754, 32'h41fed401};
test_bias[2719:2719] = '{32'h41f94410};
test_output[2719:2719] = '{32'hc51ac384};
test_input[21760:21767] = '{32'h42a9b2f6, 32'h40f42a23, 32'hc24bb959, 32'h41c782f1, 32'hc24f54da, 32'hc2ab5413, 32'hc21eaac2, 32'h41f5901c};
test_weights[21760:21767] = '{32'h424fb531, 32'h421368e0, 32'hc2022947, 32'h426d8242, 32'h429ed524, 32'hc0b6963a, 32'h4260e692, 32'h429de6df};
test_bias[2720:2720] = '{32'h4294afcf};
test_output[2720:2720] = '{32'h458b898e};
test_input[21768:21775] = '{32'h4225214c, 32'hc2878c7d, 32'hc221dd3e, 32'h4253715a, 32'hc28973cd, 32'hc207419a, 32'hc2ab8e3f, 32'hc1a364be};
test_weights[21768:21775] = '{32'hc24afc7f, 32'hc291d8a1, 32'h4298183d, 32'hc220799d, 32'hc1176e0a, 32'hc250556e, 32'h42bc5381, 32'h42c3d3e4};
test_bias[2721:2721] = '{32'hc24819a8};
test_output[2721:2721] = '{32'hc61d4809};
test_input[21776:21783] = '{32'hc2be6fc0, 32'hc2c70965, 32'hc17c94a4, 32'hc2519977, 32'hc2318735, 32'hc20bbe55, 32'h414eeca5, 32'hc275d6ea};
test_weights[21776:21783] = '{32'h4209abbc, 32'hc256df5b, 32'h428ead9a, 32'hc2c420f1, 32'hc0a3c178, 32'hc21bceed, 32'h42a44312, 32'hc13b403c};
test_bias[2722:2722] = '{32'h42a445ee};
test_output[2722:2722] = '{32'h4614f2a6};
test_input[21784:21791] = '{32'h42659b9f, 32'hc2c26f28, 32'h42b51dfd, 32'hc09ce767, 32'h421fdd4f, 32'h40f844f5, 32'hc206df17, 32'hc2621a25};
test_weights[21784:21791] = '{32'h42966f2d, 32'h42947001, 32'h42428f0e, 32'hc2bd614c, 32'h42c71db0, 32'hc2baa742, 32'hc2ba6fcd, 32'h42b342cc};
test_bias[2723:2723] = '{32'hc1e55fcd};
test_output[2723:2723] = '{32'h454ca3b5};
test_input[21792:21799] = '{32'h4244e0a5, 32'hc2bb5d02, 32'h42a4eb92, 32'hc22c599b, 32'hc2347e28, 32'h419da552, 32'hc20169c0, 32'h41cc32fe};
test_weights[21792:21799] = '{32'hc2971748, 32'h42c1d4c9, 32'h42a08ef2, 32'hc1c2889e, 32'hc1c00830, 32'hc28e3e6c, 32'h427a61ed, 32'h42744797};
test_bias[2724:2724] = '{32'hc2c76aa6};
test_output[2724:2724] = '{32'hc5bbf31d};
test_input[21800:21807] = '{32'h42c4af38, 32'hc27d2c58, 32'hc18895ce, 32'h4089356c, 32'hc215756c, 32'h4265d1f5, 32'h41fd3530, 32'hc2856fcd};
test_weights[21800:21807] = '{32'h42983021, 32'h4290b7c6, 32'h421d86ae, 32'h417140fc, 32'hc2bd3fd4, 32'hc295659c, 32'h429ed2da, 32'hc08af30f};
test_bias[2725:2725] = '{32'h4292404d};
test_output[2725:2725] = '{32'h4589fe79};
test_input[21808:21815] = '{32'hc2693aaf, 32'hc1db9bfe, 32'h41d0502a, 32'hc26be1a7, 32'h412f0386, 32'hc085ddc6, 32'hc222990d, 32'h41d9f26e};
test_weights[21808:21815] = '{32'h42815a39, 32'hc2c4c56a, 32'h411e94c3, 32'h41db6f75, 32'hc25be1c2, 32'h41930d0b, 32'h42ba04b7, 32'h4276a2c6};
test_bias[2726:2726] = '{32'h4292f41f};
test_output[2726:2726] = '{32'hc5a07b5c};
test_input[21816:21823] = '{32'hc1c95d76, 32'hc2b1c259, 32'hc269a70b, 32'hc26bd315, 32'hc22f6be1, 32'hc28fd07f, 32'h428bc377, 32'hc1a171ee};
test_weights[21816:21823] = '{32'h4282cb21, 32'h423e3987, 32'hc20edcf1, 32'h42c6a2e4, 32'hc20e722b, 32'h422ca005, 32'hc252a156, 32'hc132eeaa};
test_bias[2727:2727] = '{32'hc2c23d04};
test_output[2727:2727] = '{32'hc6663ae6};
test_input[21824:21831] = '{32'hc18d6a15, 32'hc177c94e, 32'h42bc31ea, 32'h42bc2dc3, 32'h4224a594, 32'hc2c5e8e6, 32'h422b535e, 32'h42b53a2b};
test_weights[21824:21831] = '{32'hc25ad1e6, 32'h4255fbea, 32'hbee126fa, 32'hc22ceaf7, 32'hc1a07d22, 32'h42767a66, 32'hc19b2f84, 32'h4262c0af};
test_bias[2728:2728] = '{32'h423c4f2d};
test_output[2728:2728] = '{32'hc5cc6515};
test_input[21832:21839] = '{32'h42a0ca34, 32'h426d640f, 32'h41f69015, 32'h41cad66c, 32'hc12e6ad6, 32'h42671fc4, 32'h41d1972b, 32'hc221dbc8};
test_weights[21832:21839] = '{32'hc2a7a947, 32'hc0507d77, 32'h42c2de69, 32'h400e56a6, 32'h421dcb27, 32'hc1befd9a, 32'hc2b04bf3, 32'h42acdbe7};
test_bias[2729:2729] = '{32'hc2a65108};
test_output[2729:2729] = '{32'hc634d39a};
test_input[21840:21847] = '{32'h41f392ce, 32'hc2bd7688, 32'hc21ec692, 32'h41c674df, 32'h426b5ab8, 32'hc2292547, 32'hc219f155, 32'hc0dd79b5};
test_weights[21840:21847] = '{32'hc2c3a9a2, 32'hc232fe90, 32'h41a14f5e, 32'h42499c45, 32'hc24d88d5, 32'h424ae582, 32'hc27a35dc, 32'hc229d238};
test_bias[2730:2730] = '{32'h4279fbd0};
test_output[2730:2730] = '{32'hc42d8926};
test_input[21848:21855] = '{32'hc1884fdc, 32'hc26d1444, 32'hc1d288f8, 32'hc2635a37, 32'h426cb38b, 32'hc2c32287, 32'hc145fede, 32'h421cb2cf};
test_weights[21848:21855] = '{32'h422e3e13, 32'hc1750f46, 32'h4179bb4e, 32'hc29472ec, 32'hc2053a87, 32'hc20145f7, 32'hc0526705, 32'hc1999613};
test_bias[2731:2731] = '{32'hc2c21e7b};
test_output[2731:2731] = '{32'h4587daf4};
test_input[21856:21863] = '{32'hc2b71324, 32'hc20b724f, 32'hc0cadc3a, 32'hc28e59ef, 32'hc20dd2c5, 32'hc1dd476d, 32'hc1e83a7b, 32'h41afaa54};
test_weights[21856:21863] = '{32'hc2b45f7c, 32'hc2081862, 32'hc28baf5a, 32'hc2410e07, 32'hc1d40422, 32'h4203a35b, 32'hc219f333, 32'hc240246d};
test_bias[2732:2732] = '{32'hc2c1e31b};
test_output[2732:2732] = '{32'h465009ab};
test_input[21864:21871] = '{32'hc2bac56a, 32'hc26dc5b9, 32'h42796942, 32'hc250ccc2, 32'hc2c17a3d, 32'h41822d55, 32'hc06c7900, 32'h4131bf2f};
test_weights[21864:21871] = '{32'h421c3ce1, 32'hc07522fa, 32'hc2b013e1, 32'hc282e1fd, 32'h41d91a48, 32'h42a5df4f, 32'h423deed9, 32'hc20a116e};
test_bias[2733:2733] = '{32'hc0112874};
test_output[2733:2733] = '{32'hc5e511e4};
test_input[21872:21879] = '{32'h42138520, 32'hc18a8e12, 32'hc2759e23, 32'hc1cdd688, 32'hc0a2fe6d, 32'h415c5f62, 32'hc2ab0f9c, 32'hc25972f4};
test_weights[21872:21879] = '{32'h4298366f, 32'hc12247f0, 32'h41deae63, 32'hc034a78b, 32'h41bbeeeb, 32'hc2bca4ca, 32'h409af6fd, 32'h41b9554d};
test_bias[2734:2734] = '{32'h41d0528c};
test_output[2734:2734] = '{32'hc4d70dd9};
test_input[21880:21887] = '{32'h4290f04f, 32'hc11c6269, 32'hc14bab6b, 32'hc2244b8d, 32'hc1d4edc7, 32'hc275fddd, 32'h42a468cc, 32'h40ef5fb3};
test_weights[21880:21887] = '{32'hc2bee717, 32'hc22516b1, 32'h42a3a898, 32'h4299af79, 32'h4216c3d5, 32'h42aa0d7b, 32'h422312b0, 32'hc2bca4e7};
test_bias[2735:2735] = '{32'hc2b428f3};
test_output[2735:2735] = '{32'hc660d0ce};
test_input[21888:21895] = '{32'h41232444, 32'h41cb5f0e, 32'hc22e08aa, 32'hc2ae39f7, 32'h40fe0d8f, 32'hc1fe7b6a, 32'hc26328ce, 32'hc291c449};
test_weights[21888:21895] = '{32'hc2a48950, 32'hc2495abc, 32'h40b8b1c8, 32'hc22ae182, 32'h4278c586, 32'hbeeaff10, 32'hc28653f1, 32'h428f5275};
test_bias[2736:2736] = '{32'hc297333c};
test_output[2736:2736] = '{32'h43bbfa3f};
test_input[21896:21903] = '{32'h428ca5a6, 32'hc2aa983b, 32'h42c39b77, 32'h429004be, 32'hc2c3ae1b, 32'hc2a008e8, 32'h42adddb6, 32'h424cd2e6};
test_weights[21896:21903] = '{32'hc162d134, 32'hc106cef1, 32'hc2a7b246, 32'h428e9e67, 32'hc2b7c95d, 32'h42999399, 32'h4241c56f, 32'hc2832681};
test_bias[2737:2737] = '{32'h422e362a};
test_output[2737:2737] = '{32'h43c7bd26};
test_input[21904:21911] = '{32'h42a96d45, 32'h4223843b, 32'h426ca796, 32'hc2234c99, 32'hc2574dde, 32'hc293a08a, 32'h42c541fa, 32'hc24daf4f};
test_weights[21904:21911] = '{32'hc289cf64, 32'hc2832856, 32'h41c64578, 32'h42ab71ab, 32'h40dfb7f5, 32'h42a91d94, 32'h428a0a5d, 32'hc19fcc21};
test_bias[2738:2738] = '{32'hc194f9ef};
test_output[2738:2738] = '{32'hc61224c7};
test_input[21912:21919] = '{32'h42913f11, 32'hc0c9fc94, 32'h4280b08c, 32'h41134b37, 32'h41475d01, 32'h429b81e1, 32'hc284ccaf, 32'hc27f20df};
test_weights[21912:21919] = '{32'h4198fddf, 32'hc28dafcb, 32'hc1975ca8, 32'hc2b813d7, 32'hc20ef1f2, 32'hc2914f1b, 32'h42b4fde4, 32'hc29bf974};
test_bias[2739:2739] = '{32'hc26b9674};
test_output[2739:2739] = '{32'hc5e7c608};
test_input[21920:21927] = '{32'hc23728c9, 32'h42821b6b, 32'h42181948, 32'hc2c2be1e, 32'h42a8e996, 32'hbf42718d, 32'h426310d7, 32'h4245a0b5};
test_weights[21920:21927] = '{32'hc0d0bdd4, 32'hc2a38a38, 32'h42897ec4, 32'h41018fad, 32'hc2b88e14, 32'hc259ba7c, 32'h42552f64, 32'h41fc31fd};
test_bias[2740:2740] = '{32'h417b66a7};
test_output[2740:2740] = '{32'hc5c663e0};
test_input[21928:21935] = '{32'hc17f88f9, 32'h4270649a, 32'h4138e01a, 32'hc1b2c776, 32'hc1f9de76, 32'h42984097, 32'h429a38e4, 32'hc0c4105d};
test_weights[21928:21935] = '{32'h42602c4f, 32'hc266096c, 32'hc1a7c213, 32'hc10d9b21, 32'h42c2aba9, 32'h41d91ae2, 32'h3febb9ef, 32'h4213967e};
test_bias[2741:2741] = '{32'h425bf78a};
test_output[2741:2741] = '{32'hc5a8b87f};
test_input[21936:21943] = '{32'hc08bae28, 32'h42413e76, 32'hc1c89198, 32'h42abffad, 32'h428bc63a, 32'hc1d769d9, 32'h41a3e762, 32'h4283e628};
test_weights[21936:21943] = '{32'hc2a2688e, 32'hc228ed11, 32'h41d64bf3, 32'hc215ffec, 32'hc18be846, 32'hc2684f6c, 32'h418ce5e9, 32'h418e2dcd};
test_bias[2742:2742] = '{32'hc22d0f91};
test_output[2742:2742] = '{32'hc56a7111};
test_input[21944:21951] = '{32'hc2be5200, 32'hc2a45ae7, 32'h429b4ede, 32'hc2a9801d, 32'h42b14137, 32'h423e8e6e, 32'hc1313e1e, 32'h41b8d66e};
test_weights[21944:21951] = '{32'hc12569c7, 32'hc132b0ad, 32'h41e76b20, 32'h4108c01c, 32'h40f3efa9, 32'hc2bf6ab4, 32'hc264a2b9, 32'h4128331a};
test_bias[2743:2743] = '{32'h42ab74a3};
test_output[2743:2743] = '{32'h43fabe0f};
test_input[21952:21959] = '{32'h41fbd3d2, 32'h42bd7335, 32'hc285e4f9, 32'h417a18e3, 32'h4229a5ba, 32'h41a73e7d, 32'h42b641e2, 32'h4214e531};
test_weights[21952:21959] = '{32'h412931e8, 32'h42bf6a5f, 32'hc2b18f8b, 32'h41b0ea71, 32'hc1d73e52, 32'hc230234f, 32'hc28009ba, 32'hc28be384};
test_bias[2744:2744] = '{32'h41d743a3};
test_output[2744:2744] = '{32'h45a2fde3};
test_input[21960:21967] = '{32'h42b0bbcb, 32'hc239e632, 32'h429cc1b4, 32'h4288f608, 32'hc1e7a12d, 32'h42c419af, 32'hc190ae8b, 32'hc217287f};
test_weights[21960:21967] = '{32'h42b8c413, 32'hc281fea1, 32'hc252266c, 32'hc2a64390, 32'h408eed45, 32'hc2ad5192, 32'h4081318a, 32'hc2893dfc};
test_bias[2745:2745] = '{32'hc2548a39};
test_output[2745:2745] = '{32'hc5958d63};
test_input[21968:21975] = '{32'hc1942028, 32'hc024a08c, 32'hc29b3f26, 32'h41ef48ee, 32'hc1f45262, 32'hc286302c, 32'hc2c4cd6b, 32'h428a1e3b};
test_weights[21968:21975] = '{32'h41b03f6b, 32'h42a8a347, 32'h424de7d4, 32'h41c86d8f, 32'hc28745c8, 32'h42c67d0b, 32'h411af2b7, 32'hc29a3fb5};
test_bias[2746:2746] = '{32'h422ea70d};
test_output[2746:2746] = '{32'hc665aed5};
test_input[21976:21983] = '{32'h42962bae, 32'h4233dd07, 32'hc0bb53c7, 32'hc2433d3d, 32'hc204df74, 32'h424e0db9, 32'hc2014eeb, 32'hc2c7e112};
test_weights[21976:21983] = '{32'h42bcae7e, 32'h41817d5e, 32'h42c6473f, 32'h42b34474, 32'hc288b4bb, 32'hc1d532ef, 32'hc2c76ec1, 32'h42306327};
test_bias[2747:2747] = '{32'h42b37c65};
test_output[2747:2747] = '{32'h4526412a};
test_input[21984:21991] = '{32'hc2a95dd0, 32'hc2828c43, 32'hc2a0f47f, 32'hc233c834, 32'hc1cc5986, 32'hc21118e5, 32'hc13d51d6, 32'hc1d3eb07};
test_weights[21984:21991] = '{32'hc18643a6, 32'h422bf80e, 32'h41da6ce3, 32'hc24479f5, 32'hc248d577, 32'hc2a21567, 32'h4234999a, 32'hc2b1ae5d};
test_bias[2748:2748] = '{32'hc2a90b21};
test_output[2748:2748] = '{32'h458f31b2};
test_input[21992:21999] = '{32'h418eafa1, 32'h420aebac, 32'hc2841e25, 32'hc2b62eed, 32'hc1a19c25, 32'h427c2f4a, 32'hc225b8d6, 32'hc2952c45};
test_weights[21992:21999] = '{32'hc2c23965, 32'h4276156d, 32'h42b585bc, 32'hc1016312, 32'hc1b37395, 32'h41e594f3, 32'h42a352a4, 32'h425a4b3a};
test_bias[2749:2749] = '{32'h408bf285};
test_output[2749:2749] = '{32'hc61ce539};
test_input[22000:22007] = '{32'h40f4bd04, 32'h4279c3d1, 32'hc25fb8d0, 32'h4297d86e, 32'h42c4ea88, 32'hc10fe108, 32'h42520c33, 32'h429bff09};
test_weights[22000:22007] = '{32'h428fa0e1, 32'h4058907b, 32'h41c339cd, 32'hc2186176, 32'h42c5e10f, 32'h42bf3f72, 32'h4232443a, 32'h41e0c0bc};
test_bias[2750:2750] = '{32'hbf857d9c};
test_output[2750:2750] = '{32'h461aed8c};
test_input[22008:22015] = '{32'hc20e4478, 32'h429097ab, 32'h42ac847d, 32'hc2661172, 32'h4291149a, 32'h42ace352, 32'h41d09f61, 32'hc20271d7};
test_weights[22008:22015] = '{32'h4293aa3d, 32'hc1f3e01b, 32'h427a8736, 32'h42818089, 32'hc2bdc05c, 32'hc28ef757, 32'hc1cb2d12, 32'hc199b17e};
test_bias[2751:2751] = '{32'h42084ea0};
test_output[2751:2751] = '{32'hc67d5bae};
test_input[22016:22023] = '{32'h417094c8, 32'hc10010d4, 32'hc2ae4537, 32'h42b50dd6, 32'h429e81fd, 32'hc28e3dc6, 32'h40809fc4, 32'h40ae0351};
test_weights[22016:22023] = '{32'hc18260a3, 32'h42a3062d, 32'h42567c6d, 32'h420be8ce, 32'hc25ff178, 32'h4278021e, 32'hbf4cf48b, 32'hc191b2ac};
test_bias[2752:2752] = '{32'hc0216c24};
test_output[2752:2752] = '{32'hc6316b9d};
test_input[22024:22031] = '{32'h4258327e, 32'hc26bbf3f, 32'h420358c8, 32'h42848b59, 32'h420954b6, 32'hc0e3744f, 32'hc293e8c9, 32'h421e9152};
test_weights[22024:22031] = '{32'h428221c7, 32'h4293b1b4, 32'h424f5086, 32'h42c7ad97, 32'h414aeb99, 32'h42b55175, 32'h428d3162, 32'h4251d8c0};
test_bias[2753:2753] = '{32'h4240cc8b};
test_output[2753:2753] = '{32'h4582a6ea};
test_input[22032:22039] = '{32'hc16d2356, 32'h425706f1, 32'h42957458, 32'hc27480e9, 32'h42b9219b, 32'h4283e240, 32'h42b11d81, 32'hc28a2e7a};
test_weights[22032:22039] = '{32'hc2a81ff5, 32'hc0dc7fef, 32'h42b53f97, 32'hc176295b, 32'h4285ab7a, 32'h424caf73, 32'hc08b9f37, 32'hc1e726f1};
test_bias[2754:2754] = '{32'hc2497dea};
test_output[2754:2754] = '{32'h4699f900};
test_input[22040:22047] = '{32'hc20686b8, 32'hc2b2e253, 32'hc221fac7, 32'h421c2fff, 32'h40273e1e, 32'hc0956f86, 32'h4261dcbc, 32'h4159aa05};
test_weights[22040:22047] = '{32'hc29eb946, 32'hc2c66eb9, 32'h42577c7d, 32'hc2bdefc1, 32'h422557a4, 32'hc25664e7, 32'hbf5406cd, 32'hc2ae8036};
test_bias[2755:2755] = '{32'hc2357d37};
test_output[2755:2755] = '{32'h4593e534};
test_input[22048:22055] = '{32'h4238f188, 32'hc1642db1, 32'hc265f825, 32'h3f8fb30f, 32'hc29a3c3c, 32'h4142aa62, 32'hc1be0aac, 32'hc21100d0};
test_weights[22048:22055] = '{32'h422d01b0, 32'hc23cd8a7, 32'h42701530, 32'hc2b9ed7a, 32'h42350220, 32'hc29757e4, 32'h425cbbdb, 32'hc1aad038};
test_bias[2756:2756] = '{32'h41d88cad};
test_output[2756:2756] = '{32'hc5b551e6};
test_input[22056:22063] = '{32'h42b73eb1, 32'hc2a3fcd6, 32'h42068a96, 32'hc1d70e77, 32'hc19c37b7, 32'h4272717f, 32'h42a49038, 32'h4280a89e};
test_weights[22056:22063] = '{32'hc1e40676, 32'h4247c190, 32'hc200598e, 32'h4252a37d, 32'hc153c0dc, 32'hc2c00e91, 32'hc18d223f, 32'h428d940c};
test_bias[2757:2757] = '{32'h4296d3f0};
test_output[2757:2757] = '{32'hc6350586};
test_input[22064:22071] = '{32'hc2b50a73, 32'h423fc386, 32'hc14c522d, 32'hc1b4190f, 32'hbe0fccc4, 32'h42355a09, 32'hc2320cff, 32'hc2a42467};
test_weights[22064:22071] = '{32'hc1f28614, 32'h429c286b, 32'h41efc9ef, 32'h41f4659b, 32'h42835541, 32'h41aa1f34, 32'hc28140a0, 32'hc053b252};
test_bias[2758:2758] = '{32'h42360b14};
test_output[2758:2758] = '{32'h461575a5};
test_input[22072:22079] = '{32'hc0cb96f6, 32'h42076fac, 32'h40cdba67, 32'h42954ea9, 32'h40adb6d1, 32'hc2761511, 32'hc0ad0ff9, 32'hc19ff729};
test_weights[22072:22079] = '{32'hc1f16b19, 32'h42c1cd6e, 32'hc189d9cf, 32'h4200143b, 32'h429f6eaf, 32'h4288c10b, 32'h4287edc3, 32'hc1a64289};
test_bias[2759:2759] = '{32'hc2afd255};
test_output[2759:2759] = '{32'h44f25a54};
test_input[22080:22087] = '{32'hc2b88609, 32'h4213dff6, 32'hc25d1b31, 32'hc14f7bd7, 32'hc2421657, 32'hc29b2709, 32'hbf0366eb, 32'h426450b2};
test_weights[22080:22087] = '{32'h41c7921d, 32'hc0a2213d, 32'h4232f25c, 32'h3e425cd0, 32'hc1e63dc5, 32'h42a55bbe, 32'h4210f948, 32'hc09e7da9};
test_bias[2760:2760] = '{32'hc24fb079};
test_output[2760:2760] = '{32'hc6217bce};
test_input[22088:22095] = '{32'h41ab1fc7, 32'hc02524bd, 32'hc1961a82, 32'hc2b8789e, 32'hc26b3a43, 32'hc162ec0e, 32'h42753564, 32'h4269a54e};
test_weights[22088:22095] = '{32'hc288c4b4, 32'hc1ef7b8b, 32'h4253407c, 32'h4206aed0, 32'hc277f7e0, 32'h3f437dfd, 32'h42793bdf, 32'h41deeca9};
test_bias[2761:2761] = '{32'h4282c818};
test_output[2761:2761] = '{32'h45651565};
test_input[22096:22103] = '{32'h42330612, 32'h420a72de, 32'hc2bc93fa, 32'hc119d49a, 32'hc225aae9, 32'hc27e52bd, 32'hc28781be, 32'h42022619};
test_weights[22096:22103] = '{32'hc1d677ce, 32'hc27273c8, 32'h4186abd5, 32'hc1c7d4af, 32'h427011f6, 32'h42163aa2, 32'h4299314b, 32'h4183425e};
test_bias[2762:2762] = '{32'h42755843};
test_output[2762:2762] = '{32'hc65c8411};
test_input[22104:22111] = '{32'hc2996646, 32'h42934920, 32'hc1a68d34, 32'h41eae38b, 32'hc15d7ce6, 32'hc26b6c50, 32'hc2567780, 32'h4180b8fb};
test_weights[22104:22111] = '{32'h42c2d3f9, 32'h420eceb5, 32'hc294af73, 32'h42906c80, 32'hc20938b9, 32'hc1a70059, 32'h41bce313, 32'h4235b646};
test_bias[2763:2763] = '{32'h42b01a4e};
test_output[2763:2763] = '{32'h42a42ede};
test_input[22112:22119] = '{32'hc2a90d36, 32'h429e7bab, 32'hc2205b95, 32'hc2b8785e, 32'h42af2669, 32'h42690f6c, 32'hc2801beb, 32'hc13c7da7};
test_weights[22112:22119] = '{32'h42503cf1, 32'h41b55be9, 32'h4295bc1c, 32'hc1f6efbb, 32'hc191f0da, 32'hc2bc225c, 32'hc298c746, 32'hc27be0c2};
test_bias[2764:2764] = '{32'hc0e2cfea};
test_output[2764:2764] = '{32'hc58387a4};
test_input[22120:22127] = '{32'h42a0e9ff, 32'h42a98f37, 32'h42aae93c, 32'h42359695, 32'h42aa8e7e, 32'h41de2f1b, 32'h4265e85d, 32'hc21cd565};
test_weights[22120:22127] = '{32'hc283e9a1, 32'h41e4c4b7, 32'h42af0314, 32'h41984c73, 32'h422605a8, 32'h42105dce, 32'h4271a121, 32'hc2bea3bf};
test_bias[2765:2765] = '{32'hc21dd101};
test_output[2765:2765] = '{32'h46862744};
test_input[22128:22135] = '{32'h42344d0b, 32'hc29ead9c, 32'hc2832069, 32'hc29df4fa, 32'h42631d6b, 32'h41dbf2ab, 32'hc29e0171, 32'hc2c3e910};
test_weights[22128:22135] = '{32'h41eef482, 32'hbc92c58a, 32'hc1812cdd, 32'hc2c711e7, 32'hc1ebd34c, 32'hc1d538f4, 32'hc206b765, 32'h40c0d846};
test_bias[2766:2766] = '{32'hc26b410b};
test_output[2766:2766] = '{32'h461a429f};
test_input[22136:22143] = '{32'h426164dc, 32'h428ee297, 32'hc2851a3a, 32'h42a58c62, 32'h41b51240, 32'hc1f253e8, 32'h409a968e, 32'hc2b9d2d3};
test_weights[22136:22143] = '{32'hc2be955d, 32'hc22df595, 32'h42c39845, 32'h40e268e8, 32'h41ba9133, 32'h42912ab9, 32'hc23be4f9, 32'hbff269e0};
test_bias[2767:2767] = '{32'hc29aaa85};
test_output[2767:2767] = '{32'hc67d1a1d};
test_input[22144:22151] = '{32'h3fcdbc2e, 32'h427eeea3, 32'h4201eb09, 32'h41aacac6, 32'hc124cf0e, 32'h42ae690b, 32'hc1c20d4c, 32'hc191e8f2};
test_weights[22144:22151] = '{32'h42995d8c, 32'h42c4face, 32'h42a7a4b5, 32'hc1c756f5, 32'h417543c7, 32'hc29cf4b0, 32'hc2ae0494, 32'hc2509cbf};
test_bias[2768:2768] = '{32'hc242f508};
test_output[2768:2768] = '{32'h458fd213};
test_input[22152:22159] = '{32'h420c0404, 32'h421cce78, 32'h42c52143, 32'h41fb8021, 32'h42b5afb5, 32'hc2ab0ef9, 32'h429cc633, 32'h416b3086};
test_weights[22152:22159] = '{32'hc1f95348, 32'h42544540, 32'hc19a0a65, 32'h42b5834f, 32'hc20d5763, 32'hc23285c2, 32'hc12b685b, 32'hc1adcd1b};
test_bias[2769:2769] = '{32'hc2bf23b0};
test_output[2769:2769] = '{32'h44a228e1};
test_input[22160:22167] = '{32'hc239bf4a, 32'hc2ad1492, 32'hc2ba6cc6, 32'h426aee24, 32'h420af966, 32'h42897a42, 32'hc1fef2a9, 32'hc27a5942};
test_weights[22160:22167] = '{32'h42b64673, 32'hc2b8a0bc, 32'hc24a2ed7, 32'hc28c1646, 32'h424ce99f, 32'hc2254709, 32'h4243c862, 32'h4276c621};
test_bias[2770:2770] = '{32'hc1618bac};
test_output[2770:2770] = '{32'hc505d277};
test_input[22168:22175] = '{32'hc2446735, 32'h41c61d53, 32'hc2a9e149, 32'hc24f8ff7, 32'hc2816c52, 32'hc2061ade, 32'h40fadcdb, 32'h411d7d55};
test_weights[22168:22175] = '{32'h4288853f, 32'h42910887, 32'hc1ede8ac, 32'hc171ecd1, 32'hc1275528, 32'hc28f8282, 32'h423ee61a, 32'h41bc9a2c};
test_bias[2771:2771] = '{32'hc186663a};
test_output[2771:2771] = '{32'h45a99506};
test_input[22176:22183] = '{32'hc203a1cb, 32'hc23a2321, 32'hc2a55780, 32'h419d0cdc, 32'hc293c12c, 32'hc2c3dd09, 32'h4298f1b6, 32'hc2c1d1e8};
test_weights[22176:22183] = '{32'h42a95cc1, 32'hc264ead1, 32'hc114f1e5, 32'h425af15f, 32'hc26299c7, 32'hc2c73323, 32'h41c8619f, 32'h422640d0};
test_bias[2772:2772] = '{32'hc2181cb7};
test_output[2772:2772] = '{32'h465314e9};
test_input[22184:22191] = '{32'h4205b7d6, 32'hc2c23423, 32'hc1e913c6, 32'h42a08dfe, 32'h4295043c, 32'h42b7b04f, 32'hc2253b75, 32'h42142770};
test_weights[22184:22191] = '{32'h42a4e529, 32'hc229de7d, 32'hc2ad359c, 32'h428c2e82, 32'hc24d391a, 32'hc1d347af, 32'h4249d441, 32'hc23cb113};
test_bias[2773:2773] = '{32'hc2c22903};
test_output[2773:2773] = '{32'h4597a6b1};
test_input[22192:22199] = '{32'hc1a3ccac, 32'h4201baa4, 32'h42c07184, 32'h42c2d9bb, 32'hc27aaa99, 32'hc2430da8, 32'hc2c26267, 32'hc25a5a69};
test_weights[22192:22199] = '{32'h42859b2e, 32'hc1cfaae2, 32'hc269ebd3, 32'h4209a53a, 32'hc254195c, 32'h41f111e2, 32'h41e686ab, 32'hc199e7f7};
test_bias[2774:2774] = '{32'h426b8256};
test_output[2774:2774] = '{32'hc58712ea};
test_input[22200:22207] = '{32'h3f28413f, 32'hc2b8adea, 32'h425a22a3, 32'hc1d7003a, 32'h42b523c5, 32'h41ad4f4c, 32'h428c141a, 32'hc0dcd610};
test_weights[22200:22207] = '{32'h42c509ab, 32'h419ff7d0, 32'h41a4237d, 32'h427483ef, 32'hc28d97ab, 32'h41a088d7, 32'h4299e0cf, 32'h429d448e};
test_bias[2775:2775] = '{32'hc0c3d311};
test_output[2775:2775] = '{32'hc5572f04};
test_input[22208:22215] = '{32'h418c9d75, 32'h41df5d0f, 32'hc202de46, 32'hc271fc98, 32'h424e9f25, 32'hc2b6ebc3, 32'hc2bdf17e, 32'hc2406faf};
test_weights[22208:22215] = '{32'hc2ba0263, 32'hc2a476cb, 32'hc2809638, 32'h41bdb1df, 32'hc2198a30, 32'hc29b7b9c, 32'hc26b6073, 32'h4294a6f4};
test_bias[2776:2776] = '{32'h42b0c616};
test_output[2776:2776] = '{32'h4577ef41};
test_input[22216:22223] = '{32'hc1639c6d, 32'h402fb21d, 32'hc25068e6, 32'hc1b52978, 32'h42ab24f7, 32'h42748acc, 32'h41047083, 32'hc2832fce};
test_weights[22216:22223] = '{32'hc2a5407d, 32'hc18f908e, 32'h42343a13, 32'hc25fad6b, 32'h41d6c237, 32'hc2063dd5, 32'hc2a99f7c, 32'h420abf37};
test_bias[2777:2777] = '{32'hc23881e7};
test_output[2777:2777] = '{32'hc52ad0b0};
test_input[22224:22231] = '{32'hc0336028, 32'hc22dd6e2, 32'hc00680f2, 32'h42a5df8e, 32'h41e9f85e, 32'hc195e4bf, 32'h42c33e0e, 32'hbe0935c6};
test_weights[22224:22231] = '{32'h42705dec, 32'h42abb183, 32'h421e24bc, 32'h42022b86, 32'hc292ba6a, 32'hc099c873, 32'hc2abf847, 32'hc20c54bc};
test_bias[2778:2778] = '{32'hc22bee2a};
test_output[2778:2778] = '{32'hc637ecfb};
test_input[22232:22239] = '{32'h429e7d8e, 32'h4286c53c, 32'h42bc05e7, 32'hc180452a, 32'h423af3a7, 32'hc283b879, 32'h42a3bc13, 32'h429b7129};
test_weights[22232:22239] = '{32'hc2536491, 32'hc1dab38b, 32'hc1cc564e, 32'hc13f648c, 32'h4232abbb, 32'h4250426e, 32'hc1c6c145, 32'hc1a36796};
test_bias[2779:2779] = '{32'hc1b71837};
test_output[2779:2779] = '{32'hc64ea4f5};
test_input[22240:22247] = '{32'hc2531335, 32'h425157c6, 32'h42236d88, 32'h42129afc, 32'h4278a316, 32'hc2196f7f, 32'h42be4d21, 32'hc27f84a6};
test_weights[22240:22247] = '{32'hc207fe52, 32'hc2975ff6, 32'hc2a020e8, 32'h42816dc4, 32'hc2580217, 32'h41a469e1, 32'h4083d1db, 32'h4283a030};
test_bias[2780:2780] = '{32'h429c5bde};
test_output[2780:2780] = '{32'hc62b05c3};
test_input[22248:22255] = '{32'hc20b4b0b, 32'h42b7bb16, 32'h422e1d26, 32'h4141a896, 32'h42abd657, 32'hc2c3c5de, 32'hc126d9aa, 32'hc23d3c43};
test_weights[22248:22255] = '{32'h41886015, 32'h424db222, 32'h4212dd16, 32'h41affe33, 32'hc247b371, 32'h42124b38, 32'hc1f873db, 32'hc24085d3};
test_bias[2781:2781] = '{32'h4229478e};
test_output[2781:2781] = '{32'h444022ec};
test_input[22256:22263] = '{32'h425a6e3c, 32'h429ba8e9, 32'h42b2c9ca, 32'h426e6342, 32'h428de01f, 32'hc1f37b38, 32'hc249c657, 32'h428e820f};
test_weights[22256:22263] = '{32'h4153be12, 32'h41d3619d, 32'h426a1c2b, 32'hc2b849e9, 32'hc297c63c, 32'hc2846868, 32'hc2532d15, 32'h42a193cf};
test_bias[2782:2782] = '{32'h42a3a486};
test_output[2782:2782] = '{32'h45ef2625};
test_input[22264:22271] = '{32'hc1222a41, 32'h412e56ef, 32'hc2924e79, 32'hc1023afd, 32'hc27c303d, 32'h42b6667e, 32'h420bdb35, 32'hc2983898};
test_weights[22264:22271] = '{32'h42b4b55e, 32'h41f1041d, 32'h429f50c4, 32'h418382cf, 32'h4235ef99, 32'h42bbd3e3, 32'h42308368, 32'hc290e590};
test_bias[2783:2783] = '{32'hc2826a93};
test_output[2783:2783] = '{32'h45bfe4a8};
test_input[22272:22279] = '{32'h422917c7, 32'hc199eec8, 32'h41a14572, 32'hc18d2758, 32'hc282d11d, 32'h42429676, 32'h41da5caf, 32'h422ad822};
test_weights[22272:22279] = '{32'h41d49602, 32'hc20b989c, 32'h4245ec07, 32'h4285e6d5, 32'h42599d7f, 32'hc2aa3f82, 32'h41d39c42, 32'h420772c2};
test_bias[2784:2784] = '{32'hc2789454};
test_output[2784:2784] = '{32'hc578e540};
test_input[22280:22287] = '{32'h42bcc6c0, 32'hc2a44532, 32'hc2c2bda2, 32'h421347f3, 32'h422c1088, 32'h41a65d80, 32'hc2b9239c, 32'h41d6eff6};
test_weights[22280:22287] = '{32'h428c3cab, 32'h42c5444d, 32'h42006dcc, 32'h425d3ff5, 32'h4203bb34, 32'hc28b7351, 32'h42b059ba, 32'h42bf5afb};
test_bias[2785:2785] = '{32'hc103978e};
test_output[2785:2785] = '{32'hc600379e};
test_input[22288:22295] = '{32'h40ef49a2, 32'h428bd556, 32'hc22a19db, 32'hc211a0cf, 32'hc2945e18, 32'hc24f02df, 32'hc2b066b4, 32'h42346b67};
test_weights[22288:22295] = '{32'h42851d48, 32'hc219eeaa, 32'hc28fb3a1, 32'h42543dc0, 32'h42b55b8c, 32'h42659c2f, 32'hc251262d, 32'h4182d176};
test_bias[2786:2786] = '{32'hc1f2a7dc};
test_output[2786:2786] = '{32'hc5aa3eb3};
test_input[22296:22303] = '{32'h4279ee28, 32'h410cba19, 32'hc0d7184d, 32'hc2c135a7, 32'h421d5655, 32'h42830d44, 32'hc2b7eb4c, 32'h42a7f347};
test_weights[22296:22303] = '{32'h4003fd47, 32'hc25993d6, 32'hc1ac6867, 32'h419eb96f, 32'h4296c793, 32'hc2aa6f7e, 32'hc0c85b65, 32'h4280d832};
test_bias[2787:2787] = '{32'h41e7a839};
test_output[2787:2787] = '{32'h449f5477};
test_input[22304:22311] = '{32'h40f32d5b, 32'h3f88c013, 32'h42055587, 32'h42b737e4, 32'hc2c02cc4, 32'h4277325e, 32'hc2a778bb, 32'h41f55bb4};
test_weights[22304:22311] = '{32'hc19e3ef4, 32'h421e2a08, 32'h4243095b, 32'hc226dfd1, 32'hc2452e15, 32'h41ab04dc, 32'h40e5678d, 32'h4282cab5};
test_bias[2788:2788] = '{32'hc04f7988};
test_output[2788:2788] = '{32'h45a11a82};
test_input[22312:22319] = '{32'hc08d8c6a, 32'hc1d3d217, 32'h42a5597b, 32'h41c3483a, 32'h4235a25a, 32'h4286fffb, 32'hc0b68850, 32'hc2b24b23};
test_weights[22312:22319] = '{32'hc236aae0, 32'hc24c6173, 32'hc23aeecb, 32'hc16d6093, 32'hc0b83a46, 32'h4275cf5c, 32'h426ee099, 32'hc28024ce};
test_bias[2789:2789] = '{32'h428dd585};
test_output[2789:2789] = '{32'h45d00e13};
test_input[22320:22327] = '{32'h4283ccb4, 32'hbf56dd04, 32'h42a39f64, 32'h422d134d, 32'h419653a0, 32'hc10d4fde, 32'hc26f8ad0, 32'h42a5e91a};
test_weights[22320:22327] = '{32'h428ae633, 32'h4270f706, 32'h428b3fca, 32'h4198d171, 32'h4131bc85, 32'h415ba19b, 32'hc11259b0, 32'hc1255c95};
test_bias[2790:2790] = '{32'h40fdfd15};
test_output[2790:2790] = '{32'h46294a7d};
test_input[22328:22335] = '{32'h41dbd33a, 32'h3ffb3383, 32'h421b3f40, 32'h42301f10, 32'h428e2667, 32'hc2c17c44, 32'h42972be1, 32'h41393dfa};
test_weights[22328:22335] = '{32'hc28126bd, 32'hc2a7ca98, 32'h4230f5ae, 32'h4253ff3f, 32'hc21dfc4e, 32'hc21731d9, 32'h4022fba3, 32'hc2846994};
test_bias[2791:2791] = '{32'hc24d97f7};
test_output[2791:2791] = '{32'h4511fa86};
test_input[22336:22343] = '{32'hc2189d32, 32'h4262bfad, 32'h41f96a06, 32'hc2ae1b7b, 32'h411379ea, 32'h40fc05cd, 32'hc217cf0e, 32'h41d09427};
test_weights[22336:22343] = '{32'hc1e2f5f9, 32'h4292a520, 32'hc1fa7d5a, 32'h4064bcbe, 32'h41ef63df, 32'hc11d7eae, 32'h416e3422, 32'h42acea29};
test_bias[2792:2792] = '{32'hc2a1e812};
test_output[2792:2792] = '{32'h45b3f01b};
test_input[22344:22351] = '{32'hc2193dcf, 32'hc184b9b0, 32'h425efaaf, 32'h4246daaf, 32'hc2b31163, 32'hc2887d5c, 32'hc24d0c3c, 32'h429e9011};
test_weights[22344:22351] = '{32'h42b2f84f, 32'hc21ff283, 32'hc26811df, 32'h424f95aa, 32'hc2bb8e51, 32'hc2a733de, 32'hc13ee84c, 32'h4104f914};
test_bias[2793:2793] = '{32'hc1fe23fe};
test_output[2793:2793] = '{32'h463a45a9};
test_input[22352:22359] = '{32'hc246be81, 32'h429c3234, 32'h42ae9de0, 32'hc2a11270, 32'h41a4721b, 32'h42443237, 32'hc1b7223e, 32'h4296c66c};
test_weights[22352:22359] = '{32'h42af16f2, 32'hc26a3fa6, 32'hc1fa50be, 32'h424c4961, 32'hc2c7d8f9, 32'hbfd9859f, 32'h42821cf1, 32'h4151ba24};
test_bias[2794:2794] = '{32'hc2379c04};
test_output[2794:2794] = '{32'hc690293e};
test_input[22360:22367] = '{32'h41dea7a2, 32'hc01bd68a, 32'h429e3da7, 32'h3fdd7906, 32'h427cf3b5, 32'hc27c4284, 32'h421882e8, 32'hc242acd8};
test_weights[22360:22367] = '{32'hc1f0642a, 32'hc2b38730, 32'hc2c022e8, 32'hc1ccf76f, 32'h42013bf3, 32'hc2aa9c70, 32'h412c1349, 32'h419d54c7};
test_bias[2795:2795] = '{32'hc2c0e594};
test_output[2795:2795] = '{32'hc4b974a4};
test_input[22368:22375] = '{32'h426fa753, 32'hbfea4ecd, 32'h42610bd0, 32'hc1e08f06, 32'hc1801aa8, 32'hc2498814, 32'h414dfd24, 32'hc2bcfc34};
test_weights[22368:22375] = '{32'hc2c386ff, 32'h418c1923, 32'hc217036f, 32'hc29ccb31, 32'hc1a3feb0, 32'hc2b8263b, 32'h417d1315, 32'h409eb1c7};
test_bias[2796:2796] = '{32'hc2c6d608};
test_output[2796:2796] = '{32'hc4974103};
test_input[22376:22383] = '{32'h42b309a7, 32'h426f5db1, 32'hc2b1f75c, 32'hc1f05e7c, 32'hc0f84185, 32'h421346d9, 32'hc28c7bbc, 32'h4206512b};
test_weights[22376:22383] = '{32'hc234d28b, 32'h428df428, 32'hc2afcc7e, 32'h42afc531, 32'hc2800603, 32'h425ca747, 32'hc20e91c6, 32'hbfe5db71};
test_bias[2797:2797] = '{32'h40f1ef51};
test_output[2797:2797] = '{32'h4621e04c};
test_input[22384:22391] = '{32'hc2ad536b, 32'h4255accb, 32'hc21a2465, 32'h41a10848, 32'hbf96826f, 32'hc2af1286, 32'h4261e143, 32'hc1a852e5};
test_weights[22384:22391] = '{32'h42c5b80b, 32'h427af6dd, 32'h41f8c181, 32'hc2a07dc1, 32'h42622539, 32'h42b8cf58, 32'hc05109d0, 32'hc2846b41};
test_bias[2798:2798] = '{32'h42981b79};
test_output[2798:2798] = '{32'hc668cfea};
test_input[22392:22399] = '{32'h424fc25a, 32'h41a71d96, 32'hc10bdb4d, 32'hc2a4c82b, 32'hc2c7cdfa, 32'hc1dd6d74, 32'hc1c16655, 32'h411b76f2};
test_weights[22392:22399] = '{32'h42aa53d0, 32'h421de886, 32'h425255d9, 32'h42087db2, 32'hc2162415, 32'hc1cc872e, 32'hc23effc7, 32'h42a36046};
test_bias[2799:2799] = '{32'hc1510ba1};
test_output[2799:2799] = '{32'h4602c5f5};
test_input[22400:22407] = '{32'h4187169e, 32'h4117ae0c, 32'hc2bd5a60, 32'h415a631a, 32'hc0fa21d9, 32'hc0f52235, 32'h428830bb, 32'hc23be25a};
test_weights[22400:22407] = '{32'h423edbe9, 32'hbfe109e0, 32'h41ece4fa, 32'hc1586d26, 32'h42bd5fe4, 32'h423538c4, 32'h40b647a8, 32'h42332ac1};
test_bias[2800:2800] = '{32'h415510c6};
test_output[2800:2800] = '{32'hc59be83e};
test_input[22408:22415] = '{32'h421d6c92, 32'hc28f4844, 32'hc1b02da7, 32'h42b78332, 32'h42be2182, 32'hc29ebc96, 32'h42816fe5, 32'h4254dd20};
test_weights[22408:22415] = '{32'h42a9fc8a, 32'hc275d320, 32'hc2985712, 32'h42ae82c3, 32'h4234c54d, 32'hc25bc151, 32'hc1a2986c, 32'hc298cdcd};
test_bias[2801:2801] = '{32'hc2595589};
test_output[2801:2801] = '{32'h46a15939};
test_input[22416:22423] = '{32'hc28ebb29, 32'hc23858d5, 32'hc1327730, 32'hc21ab65c, 32'hc29640f6, 32'h42bf8447, 32'hc17e29c4, 32'h42442925};
test_weights[22416:22423] = '{32'h41a6def2, 32'h42c79866, 32'h42948e9b, 32'hc251b751, 32'hc128a3c0, 32'h42963ab3, 32'hc0e32044, 32'hc108f42a};
test_bias[2802:2802] = '{32'h426de42d};
test_output[2802:2802] = '{32'h45320899};
test_input[22424:22431] = '{32'h410216bb, 32'h40b4d959, 32'h42105dc0, 32'hc1d38fbc, 32'h41035b0e, 32'h42a42284, 32'h421b498b, 32'h428dce59};
test_weights[22424:22431] = '{32'hc19c3e4c, 32'h40bee9be, 32'hc17ab3a9, 32'hc29a997e, 32'hc1e7daf8, 32'hc25a81e0, 32'h42bc9fbb, 32'hc26a4491};
test_bias[2803:2803] = '{32'hc28bbf17};
test_output[2803:2803] = '{32'hc57587c1};
test_input[22432:22439] = '{32'h42426fdc, 32'hc25cdaba, 32'h415bb272, 32'h3fbc81ff, 32'hc13a394a, 32'h4211e53c, 32'hc2bac4c3, 32'h42aded8d};
test_weights[22432:22439] = '{32'h42998b56, 32'h428c7e07, 32'h424a692c, 32'hc10bf102, 32'h42b87c82, 32'hc28c7e63, 32'hc2133fa5, 32'h41eb331f};
test_bias[2804:2804] = '{32'h41981e7d};
test_output[2804:2804] = '{32'h45360e10};
test_input[22440:22447] = '{32'hc1fe9527, 32'hc25159c8, 32'hc1b948d9, 32'h3f598879, 32'hc2096102, 32'hc2c5af4c, 32'h416738ad, 32'hc0e4de94};
test_weights[22440:22447] = '{32'h418b2baa, 32'hc2a02dd1, 32'h412c3548, 32'hc206ec5f, 32'hc18807ae, 32'h41aec1be, 32'h420766d8, 32'hc28cb38b};
test_bias[2805:2805] = '{32'h41820233};
test_output[2805:2805] = '{32'h452e991e};
test_input[22448:22455] = '{32'h41d3c037, 32'hc2626f8d, 32'h42390298, 32'hc199b3e7, 32'hc2aec067, 32'hc28325df, 32'hc29086fb, 32'hc29ec4bd};
test_weights[22448:22455] = '{32'hc216f4aa, 32'h4186ba4e, 32'hc1d788ab, 32'h417064dc, 32'h427cbaeb, 32'h41c0378f, 32'h42a9b9fb, 32'h41a2ac77};
test_bias[2806:2806] = '{32'hc2b0ef8e};
test_output[2806:2806] = '{32'hc68fe4de};
test_input[22456:22463] = '{32'h42b6daff, 32'h42ac0c7c, 32'hc29ea12d, 32'hc28f0dd4, 32'hc26fa932, 32'hc2363b09, 32'h42a09dba, 32'hc260eaae};
test_weights[22456:22463] = '{32'h42588b43, 32'hc2b7e743, 32'hc2c34ce0, 32'h42196d62, 32'h41b7021c, 32'h424c29a3, 32'hc1aa9a7c, 32'hc21496c5};
test_bias[2807:2807] = '{32'h429e8d06};
test_output[2807:2807] = '{32'hc495ef9b};
test_input[22464:22471] = '{32'hc233bb0f, 32'hc2b9dee6, 32'hc27800c7, 32'hc2b48be1, 32'h426482dc, 32'hc29bad87, 32'hc2162918, 32'hc2a87d1c};
test_weights[22464:22471] = '{32'h4204961f, 32'h424cfab5, 32'hc2c34cfc, 32'h42af2bdf, 32'h429f720d, 32'h425dce09, 32'hc297db31, 32'hc2c44f37};
test_bias[2808:2808] = '{32'h4248dab5};
test_output[2808:2808] = '{32'h454e79a0};
test_input[22472:22479] = '{32'hc2c5db84, 32'h4141b951, 32'h4219d815, 32'h4249f4ca, 32'hc1a3f569, 32'h428b0a4a, 32'hc18e2527, 32'hc24a4a0c};
test_weights[22472:22479] = '{32'hc29b870b, 32'h424745bd, 32'h4287db62, 32'hc1c8224c, 32'h40832a16, 32'h42b67f9f, 32'h4248e576, 32'h42535b5c};
test_bias[2809:2809] = '{32'hc1b20aef};
test_output[2809:2809] = '{32'h46407a5a};
test_input[22480:22487] = '{32'hc247000a, 32'hc201dd91, 32'hc2c69bce, 32'h4256c158, 32'h427fc3e8, 32'h41e02c13, 32'hc1967c11, 32'h42779fee};
test_weights[22480:22487] = '{32'h4286a7a4, 32'h4264a06b, 32'h42768664, 32'h411be9d3, 32'h42c762c2, 32'h41735539, 32'h42891494, 32'h41df4cdc};
test_bias[2810:2810] = '{32'h40048664};
test_output[2810:2810] = '{32'hc55e8e1c};
test_input[22488:22495] = '{32'hc2b88fda, 32'hc1988205, 32'hc2bce8e0, 32'h415c775f, 32'h42b17aba, 32'h4297600b, 32'hc29ddc85, 32'hc109a58d};
test_weights[22488:22495] = '{32'hc2414330, 32'h41d1b6f3, 32'hc239e8e0, 32'hc1675f74, 32'hc29f5e25, 32'h429e53e6, 32'hc248b51a, 32'h42596de1};
test_bias[2811:2811] = '{32'h4214a985};
test_output[2811:2811] = '{32'h4625a10b};
test_input[22496:22503] = '{32'h42737978, 32'h422aed8f, 32'h42ba1a08, 32'h42102363, 32'h4281deea, 32'hc2b8167c, 32'hc14d3b95, 32'h3f9b48bb};
test_weights[22496:22503] = '{32'hc0c8c972, 32'h420bd943, 32'hc127aaf8, 32'hc251f4b5, 32'h4290c576, 32'h408c52b0, 32'hc22420d1, 32'h426fca1f};
test_bias[2812:2812] = '{32'h424cc974};
test_output[2812:2812] = '{32'h45478921};
test_input[22504:22511] = '{32'hc286c3ed, 32'h42a0ce41, 32'h4293124e, 32'hc29d7b18, 32'h42a8ef70, 32'h4269ad92, 32'hc2a896e9, 32'hbef4b67d};
test_weights[22504:22511] = '{32'h42bc10dd, 32'h4113868d, 32'hc1c23af5, 32'h4252f5b1, 32'h429240ba, 32'h423f7e53, 32'h418233e6, 32'h40ba2f29};
test_bias[2813:2813] = '{32'hc260bdd2};
test_output[2813:2813] = '{32'hc57964f0};
test_input[22512:22519] = '{32'h42b4d22a, 32'h4286f255, 32'hc01eb80a, 32'h429ba5ed, 32'hc2b43fc0, 32'h41cabf30, 32'h42b55b79, 32'h429792a1};
test_weights[22512:22519] = '{32'hc2051477, 32'h3ff019f7, 32'hc180ab3d, 32'hc24cb4f9, 32'hc287b0aa, 32'h42217346, 32'hc2be99b2, 32'hc284aac5};
test_bias[2814:2814] = '{32'hc1e912ac};
test_output[2814:2814] = '{32'hc6512376};
test_input[22520:22527] = '{32'h42ab48a4, 32'hc1df30c4, 32'hc2552e1a, 32'hc2a25b1b, 32'hc29227e4, 32'h4246e1fc, 32'hc2c353f3, 32'h40fe6aa0};
test_weights[22520:22527] = '{32'hc2bb8480, 32'hc1915eab, 32'h42a6c9b9, 32'hc2acb1c7, 32'hbe3b70d0, 32'h4129e3fe, 32'h41adaedc, 32'h4283bd5b};
test_bias[2815:2815] = '{32'h42c45e2c};
test_output[2815:2815] = '{32'hc5b8d6b3};
test_input[22528:22535] = '{32'hc145cc80, 32'hc286b8ae, 32'h42bb3b25, 32'hc28cbcc9, 32'hc277fb32, 32'h4211ec8d, 32'h41df9155, 32'hc2c70d13};
test_weights[22528:22535] = '{32'hc274909e, 32'h42bcc879, 32'h426ea28a, 32'h42b6acb8, 32'hc26fa14e, 32'h40ad6cae, 32'hc013c54f, 32'h411ea14b};
test_bias[2816:2816] = '{32'h42ac0ecb};
test_output[2816:2816] = '{32'hc55aa455};
test_input[22536:22543] = '{32'h410ddda7, 32'h3feda886, 32'h41b1bc4f, 32'hc2305fbd, 32'hc281896d, 32'hc1828873, 32'h40c679ad, 32'h41f55c41};
test_weights[22536:22543] = '{32'hc1cad28d, 32'h428bfb83, 32'h420aef21, 32'hc1468c7a, 32'hbfa1f95c, 32'h4117acfa, 32'h42a362ee, 32'h42b3574e};
test_bias[2817:2817] = '{32'hc29b79fd};
test_output[2817:2817] = '{32'h4587537a};
test_input[22544:22551] = '{32'h42c1360d, 32'hc2acea87, 32'hc2b1e9d0, 32'h42144a40, 32'hc231665b, 32'h42bd075e, 32'hc2be3996, 32'h42abca48};
test_weights[22544:22551] = '{32'hc220ed35, 32'hc187e8e4, 32'h4282d966, 32'hc21223c5, 32'h4287c7a5, 32'h41ce9230, 32'hc29fcc46, 32'hc2105c62};
test_bias[2818:2818] = '{32'hc2762d3b};
test_output[2818:2818] = '{32'hc5b2e5e7};
test_input[22552:22559] = '{32'h4273473b, 32'h42be9617, 32'hc24d307e, 32'h423a0dd6, 32'h42b31630, 32'h42b811d4, 32'hc2952a1e, 32'h422723a2};
test_weights[22552:22559] = '{32'hc261153b, 32'hbee94855, 32'hc152ab97, 32'h42b4d224, 32'h42b48fa2, 32'hc1a7f496, 32'hc0216b9e, 32'hc278ed59};
test_bias[2819:2819] = '{32'h41cfe819};
test_output[2819:2819] = '{32'h45a1e419};
test_input[22560:22567] = '{32'hc2a10014, 32'h404dbf87, 32'h4264766f, 32'h425f3f3b, 32'h42a84e12, 32'h4216bf78, 32'hc09e92de, 32'hc1acf833};
test_weights[22560:22567] = '{32'h4274270b, 32'h3f2275b6, 32'h42b0ef9b, 32'h4259687b, 32'hc2922a56, 32'h42a8a641, 32'h422e7822, 32'hc23215e0};
test_bias[2820:2820] = '{32'hc293e029};
test_output[2820:2820] = '{32'h445aceb3};
test_input[22568:22575] = '{32'h40d029bb, 32'hc2a42936, 32'h42b4b408, 32'hbe8397ad, 32'h42a78e4c, 32'h42b68b36, 32'hc21d012c, 32'h42667e2e};
test_weights[22568:22575] = '{32'hc2b820dc, 32'h427695e9, 32'hc2a70ea2, 32'h4213b190, 32'h4289df79, 32'h417c5545, 32'h4282ab18, 32'h4299cae3};
test_bias[2821:2821] = '{32'hc2320118};
test_output[2821:2821] = '{32'hc5829371};
test_input[22576:22583] = '{32'hc29bc6db, 32'hc285c528, 32'hc2a0781b, 32'h4281b0ce, 32'hc2ac72d1, 32'h4218e111, 32'h427a1cac, 32'h4293477d};
test_weights[22576:22583] = '{32'hc2019774, 32'hc1a44175, 32'hc25a4bcd, 32'h42a9e7d9, 32'hc2bf1b7b, 32'hc23f70a7, 32'h4258f773, 32'hc1837f91};
test_bias[2822:2822] = '{32'h42c69c1d};
test_output[2822:2822] = '{32'h46af951c};
test_input[22584:22591] = '{32'h40bbc92c, 32'h421d908b, 32'hc1882ea5, 32'hc209b877, 32'hc1c5f239, 32'h423af458, 32'h414b5496, 32'hc262a03c};
test_weights[22584:22591] = '{32'h4255e8ec, 32'h412149fa, 32'hc298b4e6, 32'h4288a4f5, 32'hc295593f, 32'h428e7758, 32'h42777698, 32'hc26d61b7};
test_bias[2823:2823] = '{32'h426706a3};
test_output[2823:2823] = '{32'h460d465f};
test_input[22592:22599] = '{32'hc1756298, 32'hc26f22a9, 32'hc100cc19, 32'h417920af, 32'hc2628efb, 32'hc1deffb4, 32'hc2837b09, 32'hc1f9c9e4};
test_weights[22592:22599] = '{32'hc28ad27d, 32'hc23aa4a8, 32'hc157e2db, 32'h42b1a1ef, 32'h424ebae2, 32'hc1cb7286, 32'h422e0721, 32'h42a97068};
test_bias[2824:2824] = '{32'h41f57523};
test_output[2824:2824] = '{32'hc512b80c};
test_input[22600:22607] = '{32'h42c56b3b, 32'hc29bb5b4, 32'h40939ae9, 32'h42a406cc, 32'h420d4fe8, 32'h4298d245, 32'hc252daa7, 32'hc23a7755};
test_weights[22600:22607] = '{32'h42a6e3a4, 32'hc290ad04, 32'h40b87c5a, 32'hc21c64d2, 32'hc25decd5, 32'h427e939e, 32'hc19df6b9, 32'h41dfc09e};
test_bias[2825:2825] = '{32'hc23d8d31};
test_output[2825:2825] = '{32'h464f854d};
test_input[22608:22615] = '{32'h42469d33, 32'hc22c40e2, 32'h42a7fc74, 32'hc25bdabd, 32'hc28adbb3, 32'hc2519eac, 32'h42aa72d1, 32'h429b2b23};
test_weights[22608:22615] = '{32'hc1459c4a, 32'hc291c55f, 32'hc1a8a180, 32'h42140cbf, 32'h4289cf6e, 32'h41e509fa, 32'hc2bf396e, 32'h429f7b0c};
test_bias[2826:2826] = '{32'h414954d3};
test_output[2826:2826] = '{32'hc614a42b};
test_input[22616:22623] = '{32'hc12465f9, 32'hc2080bd4, 32'hc0aee473, 32'h41895e6b, 32'hc246309d, 32'h4285417a, 32'hc1e0a6e7, 32'h4059430f};
test_weights[22616:22623] = '{32'hc2566542, 32'hc28ad5b0, 32'hc2b0edbb, 32'hc27923e3, 32'h423ec744, 32'h4256ac4c, 32'hc2c750c6, 32'h426cafba};
test_bias[2827:2827] = '{32'h41dc11ad};
test_output[2827:2827] = '{32'h45cd2a39};
test_input[22624:22631] = '{32'hc2961b54, 32'h4197bc6f, 32'h429adfdc, 32'hc28aa8bb, 32'h401a8b61, 32'hc20a9e3f, 32'hc228169c, 32'h42861dd8};
test_weights[22624:22631] = '{32'hc2782973, 32'hc162362b, 32'h405b94e2, 32'hc1f5293f, 32'hc1d688da, 32'h421b2102, 32'h42bdf083, 32'h42c07e8b};
test_bias[2828:2828] = '{32'hc2b87838};
test_output[2828:2828] = '{32'h45f1e6dc};
test_input[22632:22639] = '{32'h421118f6, 32'hc23d5d32, 32'hc1d98bbf, 32'hc25f6169, 32'hc281cb1c, 32'hc1783174, 32'h40c16da5, 32'h42af01e2};
test_weights[22632:22639] = '{32'hc17e7667, 32'h4205a447, 32'h41cf2c0e, 32'hc1d32522, 32'h41c1e85d, 32'hc2a3f3ff, 32'h428b9423, 32'hc29e0293};
test_bias[2829:2829] = '{32'h42b4a247};
test_output[2829:2829] = '{32'hc5fcda6a};
test_input[22640:22647] = '{32'hc227089b, 32'hc1abdb7c, 32'hc09e985a, 32'h42a046a0, 32'hc23e512b, 32'h42b80685, 32'h42112170, 32'hc1f4dcb2};
test_weights[22640:22647] = '{32'h42918391, 32'h42ab0caf, 32'hc02a541d, 32'h42158271, 32'hc2bd03c5, 32'h4286f59a, 32'h4200add9, 32'hc13cd60f};
test_bias[2830:2830] = '{32'h42c71a88};
test_output[2830:2830] = '{32'h46238a93};
test_input[22648:22655] = '{32'hc2ab708f, 32'h3f31957b, 32'h4290e2fa, 32'h41529dc8, 32'h416e11c8, 32'h42b2f129, 32'hc116a290, 32'hc201a449};
test_weights[22648:22655] = '{32'h419bac83, 32'hc22eac18, 32'h429c9ec4, 32'h42a5b335, 32'hc2b2afb2, 32'hc1b8c164, 32'hc20cceb5, 32'h4280a5f2};
test_bias[2831:2831] = '{32'hc29e4cf4};
test_output[2831:2831] = '{32'hc322d9fd};
test_input[22656:22663] = '{32'hc1f19cfb, 32'h42221faf, 32'h4293d4b3, 32'hc2392216, 32'h42071662, 32'h42b39e48, 32'hc20d8ec8, 32'hc2b44a9e};
test_weights[22656:22663] = '{32'h4205313e, 32'h4224cf99, 32'hc2602d0b, 32'h424734b6, 32'h3f934829, 32'h42a67734, 32'hc1039b4c, 32'hc295fa65};
test_bias[2832:2832] = '{32'hc15e5933};
test_output[2832:2832] = '{32'h4608ff9d};
test_input[22664:22671] = '{32'hc29f26fc, 32'hc29bf04b, 32'h42c533c6, 32'hc2b347fd, 32'hc2b7c6bf, 32'hc0a6e8a4, 32'hc2b8eba7, 32'hc184c563};
test_weights[22664:22671] = '{32'hc1e444a3, 32'hc26187d9, 32'h40abe520, 32'h3fa51b0a, 32'h428ae6d5, 32'hc28c3e75, 32'h42172569, 32'hc2134f03};
test_bias[2833:2833] = '{32'h428fdc46};
test_output[2833:2833] = '{32'hc4da3b3e};
test_input[22672:22679] = '{32'h4282b4f4, 32'h42ba00be, 32'h410b68c4, 32'hc2830354, 32'hc2701772, 32'hc17251f8, 32'hc214d4aa, 32'h41c8e121};
test_weights[22672:22679] = '{32'hc08702f3, 32'h42433ca0, 32'h4292fc9e, 32'h42c7e175, 32'h42b2a8d2, 32'h4186d427, 32'h420ad91f, 32'hc18f5b4d};
test_bias[2834:2834] = '{32'h4098a663};
test_output[2834:2834] = '{32'hc60c9276};
test_input[22680:22687] = '{32'hc1e6e0ee, 32'hc2bf1499, 32'hc28fcf44, 32'hc1238dbf, 32'hc2793e7c, 32'hc228cd95, 32'h4289c525, 32'h415e74b4};
test_weights[22680:22687] = '{32'hc27f2113, 32'hc0aafadc, 32'hc0dc3bbc, 32'h40ed0891, 32'hc10a635f, 32'h429861de, 32'hc29a1a50, 32'h42bbf647};
test_bias[2835:2835] = '{32'hc2a3eb59};
test_output[2835:2835] = '{32'hc5794fbc};
test_input[22688:22695] = '{32'h4046fba4, 32'hc2a6485b, 32'hc1aeceb2, 32'h42295bb0, 32'h42a53971, 32'hc27c45af, 32'h422ac0e5, 32'h41a22943};
test_weights[22688:22695] = '{32'h42b9c143, 32'hc1b6f0c6, 32'hc00a168e, 32'hc1e6c53a, 32'hc2641e4a, 32'hc22587b4, 32'hc141fc00, 32'hc1a666f8};
test_bias[2836:2836] = '{32'hc05d7e3d};
test_output[2836:2836] = '{32'hc4fd8808};
test_input[22696:22703] = '{32'hc23fdc73, 32'hc2a23296, 32'hc29c8a0e, 32'hc276e0cf, 32'hc20fcfd7, 32'h42c36b85, 32'h41adcd53, 32'h42530a19};
test_weights[22696:22703] = '{32'hc26fed9b, 32'hc2bb46d5, 32'hc2aefaf8, 32'hc2303354, 32'h4293b5df, 32'h424cba9c, 32'hc28741d3, 32'hc1e5994e};
test_bias[2837:2837] = '{32'h4235128b};
test_output[2837:2837] = '{32'h4697ea39};
test_input[22704:22711] = '{32'h4266d0ae, 32'hc240840a, 32'h424fbb25, 32'hc0fbd04b, 32'hc21d91d7, 32'hc2804b1b, 32'hc1214724, 32'h41c1ef1e};
test_weights[22704:22711] = '{32'hc223f9fb, 32'hc0c50530, 32'h4258a594, 32'h429ff5df, 32'hc2642869, 32'h42b15878, 32'hc212428b, 32'hc26aa3eb};
test_bias[2838:2838] = '{32'h42068202};
test_output[2838:2838] = '{32'hc587d631};
test_input[22712:22719] = '{32'h4107245c, 32'h41214b96, 32'h4270a0c4, 32'hc049c6ac, 32'h428e2bc2, 32'hc2026b18, 32'hc21d1f54, 32'h42a8253b};
test_weights[22712:22719] = '{32'hc28d599e, 32'h422abf64, 32'hc29f0d42, 32'h428fd8c3, 32'hc1048747, 32'hc241d186, 32'hc2a636f6, 32'hc197e607};
test_bias[2839:2839] = '{32'hc22a87de};
test_output[2839:2839] = '{32'hc5200d22};
test_input[22720:22727] = '{32'h42b06bee, 32'h4260c243, 32'h41b0aa1b, 32'h420c5150, 32'h40ef7e90, 32'hc29eb382, 32'hc15a9718, 32'h4208ec96};
test_weights[22720:22727] = '{32'h4076deb4, 32'hc22d7c0d, 32'hc237eef0, 32'h4295e5ef, 32'hc1f4b14e, 32'h42bce051, 32'h42649e50, 32'hc281452b};
test_bias[2840:2840] = '{32'h421d1c53};
test_output[2840:2840] = '{32'hc62e5f0c};
test_input[22728:22735] = '{32'hc234530a, 32'h42a52fef, 32'h420704b8, 32'h42badc86, 32'h4276bf52, 32'h424948c0, 32'hc2845275, 32'h4180fbd2};
test_weights[22728:22735] = '{32'hc299b3f5, 32'hc234fdbc, 32'hc24cf567, 32'h42186300, 32'hc21bcea4, 32'h4121d232, 32'hc2547e56, 32'hc2a70e48};
test_bias[2841:2841] = '{32'hc24f2765};
test_output[2841:2841] = '{32'h44de7068};
test_input[22736:22743] = '{32'h41bedd2c, 32'h41f65e8f, 32'hc2157cb6, 32'h429cf190, 32'h42b3ed36, 32'h42c75b27, 32'hc2c0bf39, 32'h4205f570};
test_weights[22736:22743] = '{32'h42b07a76, 32'h41c3fc0f, 32'h422c9e00, 32'h42b0730d, 32'h425e61a8, 32'hc265b9d4, 32'h3f624877, 32'hc1964ceb};
test_bias[2842:2842] = '{32'hc1c420c1};
test_output[2842:2842] = '{32'h45d1a067};
test_input[22744:22751] = '{32'hc286e5f3, 32'h424c35fe, 32'h411d0407, 32'h427ae4fd, 32'h41ad0ce7, 32'hc27c4006, 32'h41a5e678, 32'hc244624f};
test_weights[22744:22751] = '{32'h42408394, 32'hc234e4d8, 32'hc1f9c77a, 32'hc29654bf, 32'hc279bce4, 32'h422fb1ab, 32'h421de06b, 32'hc10e3629};
test_bias[2843:2843] = '{32'h40effcd3};
test_output[2843:2843] = '{32'hc651e8a1};
test_input[22752:22759] = '{32'hc2650072, 32'hc2b74fdf, 32'h4171d190, 32'hc2abb8ed, 32'hc2860fba, 32'h414143b3, 32'h428228f2, 32'h4284ada6};
test_weights[22752:22759] = '{32'h420bf7d7, 32'hc25a315e, 32'h428b1b62, 32'hc27549fb, 32'h41bad359, 32'hc15c4267, 32'hc2b52a77, 32'hc297cde3};
test_bias[2844:2844] = '{32'h42036674};
test_output[2844:2844] = '{32'hc54f4760};
test_input[22760:22767] = '{32'h426579c1, 32'hc21037a4, 32'h4235d6d6, 32'hc1c0863a, 32'h42af8607, 32'h42428c66, 32'hc25fa615, 32'h429c58fd};
test_weights[22760:22767] = '{32'h42c5c4be, 32'h40fc16d3, 32'hc19f4c7a, 32'h42423754, 32'h420d8886, 32'h415a7257, 32'hc231498b, 32'h4226eb44};
test_bias[2845:2845] = '{32'hbfd431be};
test_output[2845:2845] = '{32'h46485c99};
test_input[22768:22775] = '{32'hc2bbe600, 32'hc183406f, 32'hc2905c74, 32'hc1ba559f, 32'hc0a6a236, 32'hc2986884, 32'hc2149a3d, 32'hc1559a9b};
test_weights[22768:22775] = '{32'hc2a439e3, 32'hc1fc8353, 32'h42529153, 32'h42a42ef1, 32'hc295e1bc, 32'h42b0bd4e, 32'h41c81764, 32'hc22f0d14};
test_bias[2846:2846] = '{32'h420f1c79};
test_output[2846:2846] = '{32'hc5812455};
test_input[22776:22783] = '{32'hc1eeed6b, 32'hc19c5414, 32'hc19ca027, 32'hc29c6232, 32'h41fbac5c, 32'hc275f2a5, 32'h429d212b, 32'h4257c09b};
test_weights[22776:22783] = '{32'hc2631fd0, 32'hc229263a, 32'hc2b102b6, 32'hc205672c, 32'hc2b06b2c, 32'hbcaa4c3b, 32'hc2b64007, 32'h4125a150};
test_bias[2847:2847] = '{32'h42028880};
test_output[2847:2847] = '{32'hc51af405};
test_input[22784:22791] = '{32'h42b90f15, 32'hc00bc7de, 32'h42801764, 32'h41e07864, 32'h3f321567, 32'hbf032942, 32'h410cd546, 32'hc1b99129};
test_weights[22784:22791] = '{32'h42827bf7, 32'hc29e3e01, 32'h42b76a5f, 32'h42ab017d, 32'hc27da11e, 32'h421c3f60, 32'hc2b94e5b, 32'hc2a5d72c};
test_bias[2848:2848] = '{32'hc2ad4e48};
test_output[2848:2848] = '{32'h46713d40};
test_input[22792:22799] = '{32'hc2bb8474, 32'hc1dbc3a3, 32'hc07d4dbc, 32'h42129b15, 32'hc23f39b2, 32'h4283b8d0, 32'hc2a54dc2, 32'h422f6da2};
test_weights[22792:22799] = '{32'hc25485f5, 32'h41db7f76, 32'h42c36bc3, 32'h429e71ab, 32'h424b7dba, 32'h4270d25c, 32'hc2a8782d, 32'h42a876eb};
test_bias[2849:2849] = '{32'h401cd2bc};
test_output[2849:2849] = '{32'h4693f123};
test_input[22800:22807] = '{32'h421685d8, 32'h41f3702e, 32'h42156a59, 32'hc1604223, 32'hc1f9e13d, 32'hc1b82dc6, 32'h42448b0f, 32'hc290f6e4};
test_weights[22800:22807] = '{32'h42c41780, 32'hc2bf3bc9, 32'hc190a2e1, 32'hc2bd280c, 32'h4293de0c, 32'h428390e0, 32'hc1b21927, 32'hc2922ed7};
test_bias[2850:2850] = '{32'h42a66d5b};
test_output[2850:2850] = '{32'h44ecb31e};
test_input[22808:22815] = '{32'hc180f5a2, 32'h424725a2, 32'h41dd5c72, 32'h42b6cb9a, 32'hc2929adc, 32'h4209820f, 32'hc29a71b2, 32'hc2b2da32};
test_weights[22808:22815] = '{32'h426b53e3, 32'hc2a027da, 32'h42a6bae0, 32'h41bcf5fc, 32'hc24ee321, 32'h41da3eeb, 32'h42215101, 32'h4197f0e5};
test_bias[2851:2851] = '{32'hc28f7fdc};
test_output[2851:2851] = '{32'hc41c3d42};
test_input[22816:22823] = '{32'hc2965f48, 32'h42bf0a32, 32'h428e2896, 32'hc28b6905, 32'h41fec958, 32'hc2816f99, 32'h42c27dc8, 32'hc0f50b98};
test_weights[22816:22823] = '{32'hc229e812, 32'hc2924373, 32'h425b1695, 32'hc27a4c95, 32'h42008612, 32'hc280a0fb, 32'h4205385a, 32'hc2c1d756};
test_bias[2852:2852] = '{32'h4272ffd0};
test_output[2852:2852] = '{32'h4655e97e};
test_input[22824:22831] = '{32'h4208343c, 32'hc2a5d06d, 32'hc245ed8c, 32'h425e5e99, 32'h428747da, 32'h422c0d40, 32'hc2a23f8e, 32'hc287c6b7};
test_weights[22824:22831] = '{32'h42ac9010, 32'hbfe932eb, 32'hc2232b2c, 32'h41a03168, 32'hc2aaf83d, 32'hc1d26056, 32'hbea06e22, 32'h42322145};
test_bias[2853:2853] = '{32'h420474b9};
test_output[2853:2853] = '{32'hc564959c};
test_input[22832:22839] = '{32'hc2aac277, 32'hc127e41d, 32'h42304567, 32'h410d3ffb, 32'hc2ab9676, 32'hc13f34d0, 32'hc297ec2c, 32'h42ad8db2};
test_weights[22832:22839] = '{32'hbfeaa2eb, 32'hc295855e, 32'h424531aa, 32'hc2aa29b9, 32'h42966e6a, 32'h4233f348, 32'h42595735, 32'h413433df};
test_bias[2854:2854] = '{32'hc1a0b421};
test_output[2854:2854] = '{32'hc5f3b36d};
test_input[22840:22847] = '{32'h422d75fe, 32'h4219977d, 32'h428a7423, 32'h42825001, 32'h4032f00f, 32'h428310ea, 32'h40d89cd3, 32'hc215a9a5};
test_weights[22840:22847] = '{32'h422f349b, 32'hc2add432, 32'hc2849479, 32'h421940ba, 32'hc2ae38d6, 32'h42961be3, 32'h41770d22, 32'h425b6df4};
test_bias[2855:2855] = '{32'h4286ff5a};
test_output[2855:2855] = '{32'hc43805e1};
test_input[22848:22855] = '{32'h42b697c5, 32'h4026979e, 32'h421a152c, 32'hc2a4bebd, 32'hc208a404, 32'hc2bf53c2, 32'h42152678, 32'h425574bd};
test_weights[22848:22855] = '{32'h4244becc, 32'h42880c1e, 32'hc2368496, 32'hc2579328, 32'hc27320ce, 32'h416dc4b0, 32'h4288f283, 32'hc29863c5};
test_bias[2856:2856] = '{32'hc29f6c68};
test_output[2856:2856] = '{32'h45c85b86};
test_input[22856:22863] = '{32'h40b07a76, 32'hbd0cb3c9, 32'hc18ccea7, 32'h42a3d1d5, 32'hc2645c01, 32'hc26ea03a, 32'hc2476f85, 32'h41827f0d};
test_weights[22856:22863] = '{32'hc2697f49, 32'hc29ba0d5, 32'hc2650a39, 32'hc293fb07, 32'h41eab376, 32'h42bfadf9, 32'h42215b56, 32'h41e2e19b};
test_bias[2857:2857] = '{32'hc108bdfc};
test_output[2857:2857] = '{32'hc65fc60a};
test_input[22864:22871] = '{32'h41e3ab41, 32'hc2921fd2, 32'h41622297, 32'hc06d4bdc, 32'h4247f3c7, 32'hc246c2d9, 32'hc1d38eae, 32'hc205a436};
test_weights[22864:22871] = '{32'hc1790dfb, 32'h425b3232, 32'hc205b4af, 32'h42748cb6, 32'hc2287cfe, 32'h425f3d84, 32'hc22b497b, 32'hc1ee55f5};
test_bias[2858:2858] = '{32'hc1f74e23};
test_output[2858:2858] = '{32'hc5f7be5e};
test_input[22872:22879] = '{32'hc2c4c502, 32'h42887396, 32'h42b6fc57, 32'hc1a14b40, 32'hc2c47e1a, 32'hc214afc2, 32'hc29d5598, 32'h42696dd1};
test_weights[22872:22879] = '{32'h42117680, 32'h423abb8f, 32'h429df4cf, 32'hc265afbe, 32'h4222aed8, 32'hc1518b62, 32'hc2a72a87, 32'hc23da8d1};
test_bias[2859:2859] = '{32'h42b687af};
test_output[2859:2859] = '{32'h4602f593};
test_input[22880:22887] = '{32'h4272ddbe, 32'h4154fdb7, 32'hc22bb656, 32'h428affe8, 32'h425c9cf2, 32'hc299d935, 32'hc28e19c4, 32'hc290c24c};
test_weights[22880:22887] = '{32'hc29132a1, 32'h3e50e430, 32'h42bf4764, 32'hc18636f3, 32'hc23b6259, 32'h42695862, 32'hc186e219, 32'h429a7d2c};
test_bias[2860:2860] = '{32'hc2b70b19};
test_output[2860:2860] = '{32'hc6a5e10f};
test_input[22888:22895] = '{32'h421c34df, 32'h417883cd, 32'hc1907f1a, 32'h42088de8, 32'h424a197d, 32'hc2b6b57b, 32'hc29bc81d, 32'hc207d7e6};
test_weights[22888:22895] = '{32'h408d5ef9, 32'hc26e0540, 32'h401bb9c6, 32'hc1f8d87a, 32'hc217271d, 32'h42721502, 32'h40fa5fbe, 32'hc2a1800c};
test_bias[2861:2861] = '{32'hc2757b08};
test_output[2861:2861] = '{32'hc5e1c0ca};
test_input[22896:22903] = '{32'h4239fd10, 32'hc16f2e45, 32'hc2837d71, 32'hc13c97ac, 32'hc1ea315e, 32'hc15443f7, 32'hc2a5ecd3, 32'hc294009c};
test_weights[22896:22903] = '{32'hc2c7305b, 32'hc250b9db, 32'hc2c56e38, 32'h428d793a, 32'h423cb6c9, 32'hc2ab08f8, 32'hc2aca87b, 32'h42325d9a};
test_bias[2862:2862] = '{32'h42bb1594};
test_output[2862:2862] = '{32'h45ac5568};
test_input[22904:22911] = '{32'h41cd1ed6, 32'h429893e1, 32'h41d2e18b, 32'h427905ec, 32'hc2c487e0, 32'h42a35b01, 32'hc2ac6d5d, 32'h411a2f0e};
test_weights[22904:22911] = '{32'h4289b117, 32'hc19748da, 32'hc245b0e5, 32'hc1b94bd6, 32'h417b09c1, 32'hc2be3980, 32'hc19cbc00, 32'h414c73ec};
test_bias[2863:2863] = '{32'hc1747842};
test_output[2863:2863] = '{32'hc61b3e6d};
test_input[22912:22919] = '{32'h42afe90f, 32'hc1b31aac, 32'h411892e9, 32'hc1fee487, 32'h42102746, 32'h421d775d, 32'hc2817840, 32'h427f8d38};
test_weights[22912:22919] = '{32'h42400643, 32'hc299a908, 32'hc2103bf6, 32'h42731a72, 32'hc2a54ecd, 32'hc281f2dd, 32'h41534bca, 32'hc2ab85c1};
test_bias[2864:2864] = '{32'hc1432a9b};
test_output[2864:2864] = '{32'hc6007217};
test_input[22920:22927] = '{32'hc2bc9a35, 32'hc1eee03e, 32'h42a61821, 32'h419dcd75, 32'h40006cdb, 32'hc24c6189, 32'h423953e9, 32'hc18d88b3};
test_weights[22920:22927] = '{32'hc255df4d, 32'h42570dc4, 32'h41e30cbd, 32'h425318b2, 32'hc286c57d, 32'h4270c73d, 32'h418a8281, 32'h418272da};
test_bias[2865:2865] = '{32'hc29e438d};
test_output[2865:2865] = '{32'h457da67e};
test_input[22928:22935] = '{32'hc19a3f57, 32'hc22698db, 32'hc299f3a5, 32'hc1dd2fff, 32'h42828065, 32'hc232a5bc, 32'h42c0191c, 32'hc23893a5};
test_weights[22928:22935] = '{32'h425103be, 32'h422f5837, 32'hc28c60ea, 32'hbfd6958c, 32'hc28fe24c, 32'h419134b9, 32'h4285f312, 32'hc2a02349};
test_bias[2866:2866] = '{32'hc2becb91};
test_output[2866:2866] = '{32'h45df3a02};
test_input[22936:22943] = '{32'h4292d6aa, 32'hc2b251d5, 32'hc1b8d8a9, 32'hc22e0622, 32'hc1f1bfba, 32'h42223c90, 32'hc1ef7cde, 32'hc2a4dbb1};
test_weights[22936:22943] = '{32'h4282e220, 32'h426ee57a, 32'h40ab436b, 32'hc2304327, 32'h42a74876, 32'h42b6ac2b, 32'hc2c42afb, 32'h42588305};
test_bias[2867:2867] = '{32'h42c48782};
test_output[2867:2867] = '{32'h447fbaad};
test_input[22944:22951] = '{32'h42befff7, 32'hc2a752ec, 32'h42af4221, 32'h422f9804, 32'hc012db67, 32'h42954c2d, 32'hc07b4e7d, 32'hc1de7a64};
test_weights[22944:22951] = '{32'h424f336f, 32'h41e10975, 32'hc2915d1d, 32'h41b47119, 32'h42869e8a, 32'hc1bdd8dd, 32'hc24f2275, 32'h429c1782};
test_bias[2868:2868] = '{32'hc1b507dd};
test_output[2868:2868] = '{32'hc5d16849};
test_input[22952:22959] = '{32'h423d63c2, 32'h426188bc, 32'h418b7295, 32'hc293ab35, 32'hc26f583c, 32'hc1038213, 32'h40dc3fef, 32'h42351067};
test_weights[22952:22959] = '{32'hc2c49000, 32'hc2168a45, 32'h42220e4b, 32'hc29c765c, 32'hc2aeede2, 32'h429f529f, 32'h42995362, 32'hbff56209};
test_bias[2869:2869] = '{32'h42a3d87f};
test_output[2869:2869] = '{32'h459644a2};
test_input[22960:22967] = '{32'h4265d405, 32'hc1a95a55, 32'h4281c0c5, 32'h42919a47, 32'h41c4a9cb, 32'h4239212c, 32'hc28893bb, 32'h42bcbfb8};
test_weights[22960:22967] = '{32'hc2479f6e, 32'h42493778, 32'h4238fdc4, 32'hc2c6cf3e, 32'hc25fd2da, 32'h42544a02, 32'h41c77008, 32'hc259a7c2};
test_bias[2870:2870] = '{32'h4142a3af};
test_output[2870:2870] = '{32'hc6596601};
test_input[22968:22975] = '{32'hc1d3dc2d, 32'h42c42960, 32'h42097702, 32'hc20e97e7, 32'h425960b8, 32'hc228f429, 32'h42054027, 32'hc1fba2ac};
test_weights[22968:22975] = '{32'hc2c724b7, 32'hc2a884d3, 32'h42815e5f, 32'h41e122fd, 32'hc2115db2, 32'h41c1a1d1, 32'h42bda78e, 32'h4217d169};
test_bias[2871:2871] = '{32'hc251abc8};
test_output[2871:2871] = '{32'hc5aba18d};
test_input[22976:22983] = '{32'hc20543b7, 32'h426efc54, 32'h424246de, 32'h4119d548, 32'hc0f4eed6, 32'h4296e49e, 32'h422a8003, 32'hc2b29a90};
test_weights[22976:22983] = '{32'hc21a8d1d, 32'hc2714b08, 32'hc2a47a57, 32'hc061efee, 32'hc2680df8, 32'h42909e27, 32'hc14e4bf7, 32'hc1e6012c};
test_bias[2872:2872] = '{32'h42ac5fb1};
test_output[2872:2872] = '{32'h44cf509c};
test_input[22984:22991] = '{32'h422b62df, 32'h422fc563, 32'hc1e18e21, 32'hc1a6b300, 32'hc2a70ca2, 32'hc2b1a6a9, 32'hc2aae82f, 32'hc2c53b4c};
test_weights[22984:22991] = '{32'h42a68603, 32'h42417fee, 32'hc295873f, 32'hc2a80472, 32'hc19338a3, 32'h41241262, 32'hc2908116, 32'hc23aed14};
test_bias[2873:2873] = '{32'h42274ad7};
test_output[2873:2873] = '{32'h46a414b9};
test_input[22992:22999] = '{32'hc22144a4, 32'hc164915f, 32'hc21c6c37, 32'hc28c1ef8, 32'h40ba45b8, 32'h428a6796, 32'h40e51ced, 32'hc260a6f8};
test_weights[22992:22999] = '{32'hc0b2e4d3, 32'hc278beba, 32'h42a5a5c2, 32'hc2772990, 32'h427fd76f, 32'hc1c91cca, 32'hc17971f4, 32'hc192bc31};
test_bias[2874:2874] = '{32'hc1517730};
test_output[2874:2874] = '{32'h44d9c029};
test_input[23000:23007] = '{32'hc1e9d13f, 32'h423509aa, 32'hc25a0a00, 32'hc2b448f1, 32'h429fed7a, 32'h41e04d50, 32'hc28ee51a, 32'h42ac1b99};
test_weights[23000:23007] = '{32'h421ab816, 32'hc27c96b0, 32'hc2b0d4f6, 32'hc1e02768, 32'hc1deff28, 32'hc283b4bf, 32'hbfde6ac8, 32'h41838041};
test_bias[2875:2875] = '{32'h4285aece};
test_output[2875:2875] = '{32'h445dbbc9};
test_input[23008:23015] = '{32'hc262a5d6, 32'hc2a9b9c6, 32'hc1ffa197, 32'hc20ee752, 32'hc0f91a7a, 32'h4266ecac, 32'hc256132e, 32'hc21924b2};
test_weights[23008:23015] = '{32'hc155bd61, 32'h41d4e362, 32'hc28236d3, 32'hc292105d, 32'h41a869c0, 32'h424eae9e, 32'hc1ff0ad3, 32'hc20325be};
test_bias[2876:2876] = '{32'h42a9ed93};
test_output[2876:2876] = '{32'h460d7702};
test_input[23016:23023] = '{32'hc2b3c3cd, 32'hc238fb5d, 32'hc17c361d, 32'hc18fe764, 32'hc2a7a630, 32'hc211ee4d, 32'hc23def29, 32'h419bf852};
test_weights[23016:23023] = '{32'hc1ee5f5e, 32'h427a19a8, 32'hc1cc2e45, 32'h4239c5ec, 32'hc2b45992, 32'h423372f6, 32'h4220ddfd, 32'h4203be99};
test_bias[2877:2877] = '{32'h42515cdc};
test_output[2877:2877] = '{32'h457dc998};
test_input[23024:23031] = '{32'hc226097d, 32'h41451f04, 32'h425b2849, 32'hc2943464, 32'h4292cf39, 32'hc2935955, 32'hc20cf543, 32'hc2b6ebcf};
test_weights[23024:23031] = '{32'h42480cb5, 32'h41924fe9, 32'h4295295d, 32'hc2543493, 32'h42bdf826, 32'h4287cf8b, 32'hc20a2be5, 32'hc23c93b2};
test_bias[2878:2878] = '{32'h426fcdd0};
test_output[2878:2878] = '{32'h46567533};
test_input[23032:23039] = '{32'hc1048eff, 32'hc2beae85, 32'hc250c5a5, 32'h4212ca89, 32'hc1ebfb99, 32'h420b1630, 32'h42564811, 32'h4280ae56};
test_weights[23032:23039] = '{32'hc286999c, 32'hbff92c42, 32'hc1a0791b, 32'hc25ecc06, 32'hc1a2f18d, 32'hc2c187b9, 32'h4288c57d, 32'hc20b6286};
test_bias[2879:2879] = '{32'h421f39c9};
test_output[2879:2879] = '{32'hc4c291f8};
test_input[23040:23047] = '{32'hc232c349, 32'h42960a81, 32'hc2c2dcd0, 32'h4267600e, 32'h42c6e016, 32'h3ffb3484, 32'hc27436fa, 32'h40c4f469};
test_weights[23040:23047] = '{32'hc1c516b5, 32'h404e941a, 32'h424e6024, 32'h3f922cab, 32'h420ad9f6, 32'h428300d3, 32'h3f218445, 32'h426c8101};
test_bias[2880:2880] = '{32'h4163bb43};
test_output[2880:2880] = '{32'h43972547};
test_input[23048:23055] = '{32'hc222c85c, 32'hc17feace, 32'hc2655c72, 32'h425c18b2, 32'hc29936a8, 32'hc2c7f31b, 32'h422294f0, 32'hc1ce17d0};
test_weights[23048:23055] = '{32'hc1fab1ea, 32'h42287c04, 32'hc2a07c34, 32'hc0fb0058, 32'hc22500f3, 32'hc2998f4c, 32'h40bb33d2, 32'h427f53f6};
test_bias[2881:2881] = '{32'h42419c9c};
test_output[2881:2881] = '{32'h465ea409};
test_input[23056:23063] = '{32'h4162877c, 32'hc2a2b709, 32'h4253e3a0, 32'h423ee703, 32'h42acec1a, 32'hc2454bf7, 32'hc15a5664, 32'hc098069e};
test_weights[23056:23063] = '{32'h41f5594d, 32'h42bf2dd1, 32'h4285890a, 32'h42bc5e99, 32'h421459bc, 32'h42878859, 32'hc28fbd77, 32'hc287b5d7};
test_bias[2882:2882] = '{32'h41b2f7a1};
test_output[2882:2882] = '{32'h44ead80b};
test_input[23064:23071] = '{32'hc1d4b072, 32'hc21b683e, 32'h41151e4e, 32'h4280f2be, 32'hc2be6e30, 32'hc180942b, 32'h412fe872, 32'h41f85750};
test_weights[23064:23071] = '{32'hc2699da0, 32'hc201df9c, 32'hc2839da7, 32'h42b3910e, 32'h42bf1aef, 32'h42b1cd7d, 32'hc01a6a97, 32'h42b82c98};
test_bias[2883:2883] = '{32'hc269c016};
test_output[2883:2883] = '{32'h436c5063};
test_input[23072:23079] = '{32'h42c3662b, 32'h4270bcb2, 32'h42bea96b, 32'hc2bd75c6, 32'hc2bd95cf, 32'hc2a724b2, 32'h421b9d2b, 32'hc2c53220};
test_weights[23072:23079] = '{32'hc28fec34, 32'hc07e22b4, 32'h42b14562, 32'h42821c31, 32'hc1533afa, 32'hc1c2c652, 32'h42650e45, 32'hc29fa472};
test_bias[2884:2884] = '{32'h42b56164};
test_output[2884:2884] = '{32'h4604b111};
test_input[23080:23087] = '{32'h42a2dd03, 32'h42458229, 32'h420e740d, 32'h41f4272f, 32'h429e36ed, 32'h42a62011, 32'h41c40e55, 32'h41baf3c1};
test_weights[23080:23087] = '{32'h4184b016, 32'hc2b3a483, 32'hc19056f0, 32'h4159144b, 32'hc1d16e20, 32'h42c4ec6c, 32'h42b645a2, 32'hc2b51a37};
test_bias[2885:2885] = '{32'hc29a7914};
test_output[2885:2885] = '{32'h45312b94};
test_input[23088:23095] = '{32'hc2133123, 32'hc269db06, 32'hc1a494ad, 32'hc23f188c, 32'h42c451d5, 32'hc1e4bc1a, 32'h42b1830c, 32'h418bf5ae};
test_weights[23088:23095] = '{32'hc253a633, 32'hc2b2fa61, 32'hc29027db, 32'hc1250cb6, 32'hc267e4a7, 32'hc1624066, 32'hc22a88da, 32'h41c6aa37};
test_bias[2886:2886] = '{32'h4279cde7};
test_output[2886:2886] = '{32'h44114a8a};
test_input[23096:23103] = '{32'h418c0414, 32'h420b8daf, 32'hc2344d47, 32'hc293401c, 32'hc24dc0b8, 32'hbf06e25a, 32'hc18ba126, 32'hc2963b40};
test_weights[23096:23103] = '{32'h424ca1e0, 32'hc2125bd9, 32'hc2b0cbb1, 32'hc1795ea2, 32'h428bf4f4, 32'hc28ffbc0, 32'hc1683183, 32'h4114bcc6};
test_bias[2887:2887] = '{32'h4261ae4a};
test_output[2887:2887] = '{32'h44482b3c};
test_input[23104:23111] = '{32'hc2ba9013, 32'hc077be9f, 32'hc290dbab, 32'h41c75829, 32'h42a9e510, 32'hc1d94a7f, 32'h42a41e2f, 32'hc1fffb7a};
test_weights[23104:23111] = '{32'h41bfbb0b, 32'hc1e6c19e, 32'h40dc9b9a, 32'h427a1d76, 32'h42956d9a, 32'h41c47bfa, 32'hc12a8f33, 32'hc2c4dfc7};
test_bias[2888:2888] = '{32'hc202869d};
test_output[2888:2888] = '{32'h45d646fc};
test_input[23112:23119] = '{32'hc29d1ae3, 32'hc226c3c6, 32'hc1502c88, 32'hc2becc72, 32'h41eea6fd, 32'hc1ebe385, 32'h41383788, 32'hc2a1478b};
test_weights[23112:23119] = '{32'hc07d1d07, 32'hc26dd386, 32'h41bb43dc, 32'h4187f498, 32'hc194ac11, 32'hc20d5200, 32'hc1e707cf, 32'hc2844422};
test_bias[2889:2889] = '{32'hc27cc002};
test_output[2889:2889] = '{32'h45c4824f};
test_input[23120:23127] = '{32'hc2a4fc65, 32'h42814939, 32'hc1ec7807, 32'h424da1ad, 32'h4280c050, 32'h41a5a8e5, 32'hc223d927, 32'h400bce0b};
test_weights[23120:23127] = '{32'hc2073fc3, 32'hc28a7f9a, 32'hc2260509, 32'h42c5d366, 32'hbea9a21e, 32'hc2177324, 32'hc27d2d4d, 32'h426d57c4};
test_bias[2890:2890] = '{32'h42aceb2a};
test_output[2890:2890] = '{32'h45cf1f33};
test_input[23128:23135] = '{32'hc0bc0636, 32'hc23c5d45, 32'hc2b13d61, 32'hc12a3f68, 32'h425c78a5, 32'h428a5bc6, 32'hc2b02bf3, 32'h42c72029};
test_weights[23128:23135] = '{32'h42c50bba, 32'h426c8a72, 32'hc29e2b3a, 32'h4230ec61, 32'h411aba3f, 32'hc24bcdc4, 32'hc296a66c, 32'hc2315334};
test_bias[2891:2891] = '{32'h41fa966c};
test_output[2891:2891] = '{32'h4518317f};
test_input[23136:23143] = '{32'hc28a937c, 32'hc1e3abfd, 32'hc2b46e01, 32'hc2152f5a, 32'hc2265e58, 32'hc0f3c456, 32'hc283893d, 32'hc23a4441};
test_weights[23136:23143] = '{32'h42c21712, 32'h413b3c6f, 32'hc21b9324, 32'hc26a33dd, 32'h427a40ff, 32'hc1663d12, 32'hc275a4ba, 32'hc2c7a237};
test_bias[2892:2892] = '{32'h42011421};
test_output[2892:2892] = '{32'h4597f142};
test_input[23144:23151] = '{32'h41aa80fc, 32'h40935b5e, 32'hc1822956, 32'h4295971d, 32'h429d3ea3, 32'h42af13f9, 32'hc23a7ddf, 32'h3f1cf9f3};
test_weights[23144:23151] = '{32'h423b67da, 32'h429a04a6, 32'hc2948323, 32'h42785e1b, 32'hc009c871, 32'h4128ddd3, 32'h42a9e504, 32'h429c2b06};
test_bias[2893:2893] = '{32'h42af1cbb};
test_output[2893:2893] = '{32'h458138a2};
test_input[23152:23159] = '{32'h42884500, 32'h418ab06e, 32'h4297d052, 32'h4278a88c, 32'hc2a434ef, 32'h418664f3, 32'hc28b3382, 32'h42847586};
test_weights[23152:23159] = '{32'h42b364b8, 32'h42c1689e, 32'hc106b8ba, 32'hc26cd724, 32'h42922e48, 32'h42bee730, 32'hc28dccba, 32'h42191990};
test_bias[2894:2894] = '{32'h414965db};
test_output[2894:2894] = '{32'h45ccc62e};
test_input[23160:23167] = '{32'h42af8574, 32'hc285a24b, 32'hc1f2e1f4, 32'hc28174ab, 32'h42c2572f, 32'hc22ea02f, 32'hc1acddde, 32'h419f9874};
test_weights[23160:23167] = '{32'hc28ceff1, 32'h429ce85c, 32'hc2501c91, 32'h427b6f69, 32'hc244ebc9, 32'h4242e7c9, 32'h42c06a2d, 32'h423f36b5};
test_bias[2895:2895] = '{32'hc2737dab};
test_output[2895:2895] = '{32'hc6abf92f};
test_input[23168:23175] = '{32'h42ab86d8, 32'h41fd0268, 32'h422c6794, 32'hc25ce814, 32'h41cc1627, 32'h42ba2d0b, 32'hc28e40aa, 32'h42c20be1};
test_weights[23168:23175] = '{32'hc1d5ec96, 32'h4288c642, 32'hc2a0978b, 32'h419f7eaf, 32'hc2907ac0, 32'h41bd13db, 32'h4034fd53, 32'hc288842b};
test_bias[2896:2896] = '{32'h41467214};
test_output[2896:2896] = '{32'hc62e2a4f};
test_input[23176:23183] = '{32'h41ba1cf5, 32'h420c9dd7, 32'hc2c35b18, 32'hc2c6d910, 32'h41eccf9c, 32'h41ab03a2, 32'hc2129111, 32'h428904b0};
test_weights[23176:23183] = '{32'h42af66c9, 32'hc1be9c85, 32'hc29ab2b4, 32'h42a0a899, 32'hc2a46929, 32'hc253381d, 32'hc1ceaa2f, 32'h4295818c};
test_bias[2897:2897] = '{32'hc1ebefa1};
test_output[2897:2897] = '{32'h454af799};
test_input[23184:23191] = '{32'h40c2638a, 32'h427fa3de, 32'hc28335e5, 32'hc0f93128, 32'hc2495d3a, 32'h4283fd31, 32'h4253c9bd, 32'hc1c7e86d};
test_weights[23184:23191] = '{32'hc229343b, 32'hc1b340c1, 32'hc2b5d4eb, 32'h423c4ca1, 32'h3dafb8bb, 32'h42ba39af, 32'hc2445d8c, 32'h41b34537};
test_bias[2898:2898] = '{32'hc2a12522};
test_output[2898:2898] = '{32'h45d4cead};
test_input[23192:23199] = '{32'hc253ee65, 32'h42003914, 32'hc0cb2dce, 32'h41e8c310, 32'h429e43ee, 32'h422a98fe, 32'h429e5188, 32'h42069203};
test_weights[23192:23199] = '{32'hc2a1f8e3, 32'h41cb713e, 32'h4290e4d5, 32'hc1c64f9f, 32'h4292c986, 32'h41d428bb, 32'h4231e081, 32'h415fa96b};
test_bias[2899:2899] = '{32'hc267f443};
test_output[2899:2899] = '{32'h466730aa};
test_input[23200:23207] = '{32'h41d585a9, 32'hc11d2e91, 32'h42b62e8f, 32'hc143112d, 32'h4280799c, 32'hc1551e98, 32'h41741bdd, 32'h4216fef1};
test_weights[23200:23207] = '{32'h4288493a, 32'h42809280, 32'hc1be9093, 32'h4148d33a, 32'h41874aa0, 32'hc22dfdb1, 32'hc222577e, 32'h4033b940};
test_bias[2900:2900] = '{32'hc1bdf120};
test_output[2900:2900] = '{32'hc0db417e};
test_input[23208:23215] = '{32'h4083db54, 32'hc1d0d146, 32'h426aafb3, 32'h41a14aef, 32'hc203631c, 32'h42765914, 32'h424463dc, 32'h42113ab3};
test_weights[23208:23215] = '{32'h42c401d0, 32'hc29fb0f9, 32'h415c35f0, 32'hc2c40c20, 32'h411b3868, 32'h423a09ab, 32'hc2803e47, 32'hc1ca71d1};
test_bias[2901:2901] = '{32'h42b65437};
test_output[2901:2901] = '{32'hc2dde13a};
test_input[23216:23223] = '{32'hc135a8f3, 32'hc1958ed8, 32'hc2b3f269, 32'h42aa5337, 32'hc2190ea6, 32'h42a0459b, 32'h42601790, 32'h41b2f54d};
test_weights[23216:23223] = '{32'h421f1a2e, 32'h42421e75, 32'hc291da92, 32'hc1ef4872, 32'h4237e950, 32'h42ad4876, 32'hbf161e46, 32'hc1b5f661};
test_bias[2902:2902] = '{32'h42b19d83};
test_output[2902:2902] = '{32'h45e6d29f};
test_input[23224:23231] = '{32'hc298b8d3, 32'hc2364e76, 32'hc262f3f4, 32'hc2beff59, 32'h41b5523f, 32'h414fce71, 32'h42c0746f, 32'hc28009df};
test_weights[23224:23231] = '{32'hbec7c34b, 32'hc16c93a0, 32'hc25cd119, 32'hc25453e0, 32'h42850a7e, 32'h4286b31f, 32'h4152843c, 32'h41d75ae4};
test_bias[2903:2903] = '{32'h41832bbc};
test_output[2903:2903] = '{32'h46297ac6};
test_input[23232:23239] = '{32'h41c48fc2, 32'h42825981, 32'h4278d936, 32'hc28aa7d8, 32'h427405c2, 32'h413d6522, 32'h4260cf4f, 32'hc01e8ce3};
test_weights[23232:23239] = '{32'hc25df9ef, 32'h42473296, 32'h408f7056, 32'hbfbd5212, 32'hc2811552, 32'hc2169fee, 32'h42a51ec7, 32'h3eb4b8e4};
test_bias[2904:2904] = '{32'h42813958};
test_output[2904:2904] = '{32'h452183e0};
test_input[23240:23247] = '{32'h407e9a02, 32'hc1b169de, 32'hc23952a2, 32'hc22fe02e, 32'h4279af13, 32'hc1a6cedb, 32'hc2c23e39, 32'h42a4a73d};
test_weights[23240:23247] = '{32'h41b2b456, 32'hc291eecd, 32'hbea547df, 32'h41ece11a, 32'h42a1ebc6, 32'hc018a7b8, 32'hc2bd27a0, 32'hc2c77d73};
test_bias[2905:2905] = '{32'h4284ce7a};
test_output[2905:2905] = '{32'h45cd1d43};
test_input[23248:23255] = '{32'h41cf0de1, 32'hc096866e, 32'h42aa4c39, 32'hc2bd6ce2, 32'h42bece9f, 32'hc1d0fe4e, 32'hc268e292, 32'hc22e6c4f};
test_weights[23248:23255] = '{32'hc252ace0, 32'hc2b41142, 32'hc06d55f6, 32'h427f44df, 32'h41b37f65, 32'h425b9327, 32'hc2853972, 32'hc218b6e0};
test_bias[2906:2906] = '{32'hc1b60403};
test_output[2906:2906] = '{32'hc4861c2c};
test_input[23256:23263] = '{32'hc20d067b, 32'hc227ed52, 32'hc2c06fc1, 32'hc2275c2b, 32'h42926e82, 32'h41f1ddfd, 32'hc2a8eff4, 32'h420854d4};
test_weights[23256:23263] = '{32'hc294ce50, 32'hc00ce791, 32'h427391db, 32'hc2a030c4, 32'h426c7969, 32'h424e7e13, 32'hc224e858, 32'hc2649115};
test_bias[2907:2907] = '{32'hc14553a7};
test_output[2907:2907] = '{32'h45ee1bd4};
test_input[23264:23271] = '{32'hc23d0c6c, 32'h42826701, 32'hc287523c, 32'h42800d68, 32'hc234296f, 32'h40f90725, 32'h428d04ef, 32'h411c08bc};
test_weights[23264:23271] = '{32'hc2aa779b, 32'hc292df2b, 32'hc18f2080, 32'h41cf2d69, 32'hc207ff56, 32'h4276bce6, 32'hc2a068d9, 32'h42368a38};
test_bias[2908:2908] = '{32'hc2493f17};
test_output[2908:2908] = '{32'hc48e88f9};
test_input[23272:23279] = '{32'hc231afcd, 32'h42bfa90c, 32'h42903e7d, 32'h420c87a0, 32'h42b99c81, 32'h418cb1dc, 32'h42848032, 32'h421b3ff1};
test_weights[23272:23279] = '{32'hc28727e9, 32'hc2ad79c2, 32'hc205a611, 32'h4250202b, 32'hc284e7ce, 32'hc2c11882, 32'hc21ccac3, 32'hc2b6d4d1};
test_bias[2909:2909] = '{32'h428cbbee};
test_output[2909:2909] = '{32'hc69aef5d};
test_input[23280:23287] = '{32'h42a50eba, 32'hc21b3264, 32'hc2853540, 32'h42038399, 32'hc12992a4, 32'h424e78d6, 32'h4280cb48, 32'h4202c040};
test_weights[23280:23287] = '{32'h41eb36ab, 32'hc1dfe80b, 32'h42b1b3cb, 32'hc2c08aa5, 32'h41b66fb5, 32'h423d747e, 32'hc2aac95a, 32'h4154ca22};
test_bias[2910:2910] = '{32'h42b99b8d};
test_output[2910:2910] = '{32'hc6024c56};
test_input[23288:23295] = '{32'hc2bc1f71, 32'hc2041ba8, 32'hc10f0b86, 32'h42bd0b04, 32'hc1e4ec02, 32'h427287f0, 32'h41adff86, 32'h41430f17};
test_weights[23288:23295] = '{32'h40dcd371, 32'hc1ea4da1, 32'hc284e9e5, 32'h41f60b49, 32'h42a928ca, 32'hbfd28741, 32'h42a4a24e, 32'hc28e2c91};
test_bias[2911:2911] = '{32'h424cc89a};
test_output[2911:2911] = '{32'h450e2566};
test_input[23296:23303] = '{32'hc2b1928f, 32'hc292d46d, 32'h426445de, 32'hc226acb7, 32'hc2908bac, 32'hc2815a56, 32'hc141c822, 32'hc2be6a2b};
test_weights[23296:23303] = '{32'hc2bc3772, 32'h41fd22ab, 32'hc256ee3b, 32'h4233a49d, 32'h42b2e452, 32'h429c470a, 32'h40ca6cd6, 32'hc298a803};
test_bias[2912:2912] = '{32'hc26c3bb3};
test_output[2912:2912] = '{32'hc54dc2de};
test_input[23304:23311] = '{32'hc26daac0, 32'h42c2a438, 32'hc181c9fa, 32'hc2582f42, 32'hc1d6ce87, 32'h42c6d540, 32'h40bc42c2, 32'hc2a29dd8};
test_weights[23304:23311] = '{32'h425024cc, 32'hc228e798, 32'hc28a761a, 32'h41d3475d, 32'h42c20f0e, 32'hc21796db, 32'hc26b86f0, 32'hc26b764a};
test_bias[2913:2913] = '{32'hc290197e};
test_output[2913:2913] = '{32'hc6149a73};
test_input[23312:23319] = '{32'h42ba75c8, 32'hc199e470, 32'h4266d5d6, 32'h42c61e1b, 32'h42283e51, 32'h4269e9d2, 32'h429a26e0, 32'hc243bb74};
test_weights[23312:23319] = '{32'h42b26eee, 32'hc28c3676, 32'hc2ad7401, 32'hc115dabb, 32'hc2b15acb, 32'h42a84dc7, 32'h42996fd4, 32'h4285f777};
test_bias[2914:2914] = '{32'h4258cc7c};
test_output[2914:2914] = '{32'h45edf3d0};
test_input[23320:23327] = '{32'hc0b0030d, 32'hc1ef8ff6, 32'h429cbda2, 32'hc2b24014, 32'h412067c9, 32'h4254ec26, 32'h400bfe34, 32'hc1bd0464};
test_weights[23320:23327] = '{32'h4289af85, 32'hc23111a2, 32'h4257e8b4, 32'h42a371bc, 32'hc28082c2, 32'h42818da0, 32'h41b22c1a, 32'hc2281004};
test_bias[2915:2915] = '{32'h427c8fca};
test_output[2915:2915] = '{32'h44e1445f};
test_input[23328:23335] = '{32'h4281e827, 32'h420e6a05, 32'hc285ad5f, 32'hc28f4021, 32'h4208754d, 32'hc236e0f1, 32'h40ea2fec, 32'h41f976a5};
test_weights[23328:23335] = '{32'hc2920e68, 32'h423ce27b, 32'h42bc78e0, 32'hc2b5326f, 32'hc004b203, 32'hc293c01a, 32'hc2918934, 32'h413a9e46};
test_bias[2916:2916] = '{32'hc2bba4e0};
test_output[2916:2916] = '{32'h432c813b};
test_input[23336:23343] = '{32'hc260a7fc, 32'hc287912d, 32'h426b0ad5, 32'h41dcd707, 32'hc2aedcb4, 32'h420cc58d, 32'hc0e868b8, 32'h42ad36a6};
test_weights[23336:23343] = '{32'h41cc5ec1, 32'hc2548cb6, 32'hc24f9adf, 32'hc28a9298, 32'hc1dd59b7, 32'hc1dbfb55, 32'h40e5c917, 32'h419e7d55};
test_bias[2917:2917] = '{32'h4124d507};
test_output[2917:2917] = '{32'h43a4fe37};
test_input[23344:23351] = '{32'hc290ba8c, 32'h42be1069, 32'h425dda07, 32'hc28d302d, 32'h42207fe4, 32'hc2bec6f2, 32'h41b2f127, 32'hc242b062};
test_weights[23344:23351] = '{32'hc242fd8e, 32'hc2bd5575, 32'h4262c823, 32'hc18e3d6f, 32'hc0a6cbca, 32'hc255173b, 32'hc293e6fd, 32'hc24f3273};
test_bias[2918:2918] = '{32'hc21f6cb7};
test_output[2918:2918] = '{32'h4590b434};
test_input[23352:23359] = '{32'h42437c08, 32'h42abf807, 32'hc284cb64, 32'hc2517826, 32'hc290cddb, 32'hc29cdfed, 32'h42717ca3, 32'hc2ae9512};
test_weights[23352:23359] = '{32'h42048591, 32'h4293ebc7, 32'h418d8397, 32'hc084f893, 32'h3f5d39d5, 32'hc2b3dd71, 32'h428d6515, 32'hc1a2dc6e};
test_bias[2919:2919] = '{32'hc19c32e0};
test_output[2919:2919] = '{32'h469c8d9a};
test_input[23360:23367] = '{32'h428aca2b, 32'hc280b2d2, 32'hc202fd0e, 32'h428f4b01, 32'h4211ad1b, 32'h4135cad1, 32'hc2726590, 32'hc2879a9b};
test_weights[23360:23367] = '{32'hc2c34a41, 32'h3e840424, 32'h41ee27a9, 32'hc26fbba4, 32'hc2bcaa06, 32'hc1078927, 32'hc2a06aa8, 32'h4230b481};
test_bias[2920:2920] = '{32'h41b75193};
test_output[2920:2920] = '{32'hc6562414};
test_input[23368:23375] = '{32'h42a67f44, 32'hc2c0dc81, 32'hc0e34230, 32'hc296e303, 32'h42914223, 32'h41eba579, 32'hc1dab0e0, 32'hc1d00d69};
test_weights[23368:23375] = '{32'h42c09487, 32'hc2ab5310, 32'h408df388, 32'hc283f029, 32'h41e9c203, 32'h425462e6, 32'h42b5f13c, 32'hc2b0bc2e};
test_bias[2921:2921] = '{32'hc28d1b9a};
test_output[2921:2921] = '{32'h46c091be};
test_input[23376:23383] = '{32'hc205f1a8, 32'hc2b40296, 32'hc1cbf77b, 32'h42818405, 32'h4216d0e6, 32'h421f7bf0, 32'hc29ff77d, 32'h419cc6a2};
test_weights[23376:23383] = '{32'hc1ca0f98, 32'h4187580a, 32'hc1abc312, 32'hc21b976b, 32'h4171f826, 32'hc2463301, 32'hc29a97bb, 32'h424a89e1};
test_bias[2922:2922] = '{32'h428a255f};
test_output[2922:2922] = '{32'h45475e99};
test_input[23384:23391] = '{32'h427c825f, 32'hc18cc31c, 32'hc2c26788, 32'hc0911593, 32'h418f7982, 32'hc1f14bc3, 32'hc268bd52, 32'h41d848a3};
test_weights[23384:23391] = '{32'hc26fb6ee, 32'h428d93a7, 32'h4102f6c6, 32'h423baad6, 32'h41a5dc12, 32'hc25a141d, 32'h42455a26, 32'hc281b844};
test_bias[2923:2923] = '{32'hc16f5db1};
test_output[2923:2923] = '{32'hc6074fe8};
test_input[23392:23399] = '{32'hc263cff3, 32'h4101a4ca, 32'h41512470, 32'hc24d5ee5, 32'h42378b8b, 32'hc1ebe8b5, 32'hc2a5e5dd, 32'hc195651f};
test_weights[23392:23399] = '{32'hc297b35f, 32'hc132fc2c, 32'h41f0b815, 32'h4219971e, 32'h41a12881, 32'h428da9aa, 32'h41aeb427, 32'h40a98bf2};
test_bias[2924:2924] = '{32'h42b40e6e};
test_output[2924:2924] = '{32'hc3a6c69a};
test_input[23400:23407] = '{32'hc07bff93, 32'h41b6f9b8, 32'h42bd282d, 32'h428a7079, 32'h42512bd0, 32'h429c7806, 32'h4214be9c, 32'hc2ae2ef5};
test_weights[23400:23407] = '{32'h42438bc6, 32'hc2277ec3, 32'hc29030f0, 32'h42a58980, 32'h40db1e58, 32'h4194fad8, 32'hc2c49e2a, 32'hc2a695ea};
test_bias[2925:2925] = '{32'hc22de020};
test_output[2925:2925] = '{32'h4543a347};
test_input[23408:23415] = '{32'h4284d764, 32'h42b722f8, 32'h42304e82, 32'hc2207e0f, 32'hc28e3ead, 32'h422b8e41, 32'h42ba05e0, 32'h423dc861};
test_weights[23408:23415] = '{32'hc25b8dab, 32'hc2994b9f, 32'hc28db37f, 32'h421bc9b4, 32'h3edc08cb, 32'hc2292841, 32'h415a8960, 32'hc279ce5a};
test_bias[2926:2926] = '{32'h429a2886};
test_output[2926:2926] = '{32'hc692f345};
test_input[23416:23423] = '{32'h42aa69ed, 32'h4265f3ba, 32'h41ea7a13, 32'hc21ae6a6, 32'hc267eb7d, 32'hc21b4cf8, 32'hc20a17d6, 32'h42603d22};
test_weights[23416:23423] = '{32'hc223ff8a, 32'hc1bbb9ea, 32'hc2b5e9e3, 32'hc28712f7, 32'hc2288d14, 32'hc2ac7bcd, 32'h428156fa, 32'h4299f1b2};
test_bias[2927:2927] = '{32'h4247c8f4};
test_output[2927:2927] = '{32'h453d6e50};
test_input[23424:23431] = '{32'hc212dcec, 32'h42289bd2, 32'hc25910d3, 32'h426d419d, 32'hc289f953, 32'h413db354, 32'h421a7231, 32'h42a00006};
test_weights[23424:23431] = '{32'hc14386b8, 32'hc185419e, 32'hc1862d34, 32'h42830820, 32'h42bd6962, 32'hc2c606cc, 32'hc1a18dd4, 32'h42a5de13};
test_bias[2928:2928] = '{32'hc2a7ad4a};
test_output[2928:2928] = '{32'h4522e760};
test_input[23432:23439] = '{32'hc2bcbbf3, 32'h4092926f, 32'h42b41287, 32'h42b95564, 32'hc1065cb9, 32'hc21737f3, 32'h42bb9ea9, 32'hc2ab548b};
test_weights[23432:23439] = '{32'hc222b948, 32'hc28d779e, 32'h41b144c1, 32'h418ee790, 32'h428e28c9, 32'hbe17ff6a, 32'h420d6250, 32'hc1797aaa};
test_bias[2929:2929] = '{32'hc0a14b57};
test_output[2929:2929] = '{32'h462f522e};
test_input[23440:23447] = '{32'h42ae1afb, 32'hc215e8a1, 32'h42494bde, 32'h3fff164c, 32'hc297cdd9, 32'hc24fedc0, 32'h42a6cd73, 32'h429b8cd9};
test_weights[23440:23447] = '{32'h405860f3, 32'hc11a1986, 32'h41f17a76, 32'hc2bbed6c, 32'h42a95a80, 32'hc287eb69, 32'h423cb271, 32'hc27c1021};
test_bias[2930:2930] = '{32'hc24cb01a};
test_output[2930:2930] = '{32'hc4f0a7c2};
test_input[23448:23455] = '{32'hc2a8260b, 32'hc2942db0, 32'hc0acefac, 32'hc1929e77, 32'hc10e9ae9, 32'hc1bbfd33, 32'h42921ac8, 32'hc135356c};
test_weights[23448:23455] = '{32'h4093a577, 32'hc2b686ed, 32'h422a35a1, 32'hc2428deb, 32'h42b415eb, 32'hc20f85ae, 32'hc2377c72, 32'h426f678a};
test_bias[2931:2931] = '{32'h4290d90a};
test_output[2931:2931] = '{32'h4542f596};
test_input[23456:23463] = '{32'h40e27b10, 32'h4218e2ef, 32'hc20761e0, 32'hc2678551, 32'h4266960d, 32'hc0c6412b, 32'hc1a1ea9b, 32'h42679ec0};
test_weights[23456:23463] = '{32'hc2720565, 32'hc2be1acb, 32'hc2346c2a, 32'h409c26af, 32'hc1016253, 32'hc2ab1d8d, 32'hc2038642, 32'h42a1bd52};
test_bias[2932:2932] = '{32'h41f3ae9e};
test_output[2932:2932] = '{32'h452418ab};
test_input[23464:23471] = '{32'hc28fae10, 32'hc04fc6e0, 32'h42b78e92, 32'hc0bee255, 32'h3e957a77, 32'hc22dff0a, 32'h429854ab, 32'hc18bae8e};
test_weights[23464:23471] = '{32'h42674cf4, 32'h41ceb27a, 32'hc2963664, 32'hc27b0c09, 32'hc0be54d2, 32'h42308294, 32'h4244ccee, 32'hc1d876a1};
test_bias[2933:2933] = '{32'h42b1a41c};
test_output[2933:2933] = '{32'hc602c5b6};
test_input[23472:23479] = '{32'h41ae2dd9, 32'h429bbfb5, 32'hc1312be5, 32'hc2b9e782, 32'hc2bbe6f3, 32'h42bb4285, 32'hc29fc167, 32'hc149c9aa};
test_weights[23472:23479] = '{32'hc2647cea, 32'h41d14740, 32'hc1c9b7eb, 32'hc25b0dc4, 32'h420e35c9, 32'hc29254bb, 32'hc2c0ae4c, 32'h40189738};
test_bias[2934:2934] = '{32'hc24951b0};
test_output[2934:2934] = '{32'h45603775};
test_input[23480:23487] = '{32'h42add92b, 32'hc2769141, 32'hc21cef2f, 32'hc27399f7, 32'hc2b0139e, 32'h42c3746f, 32'hc203fa75, 32'hc1a7b70f};
test_weights[23480:23487] = '{32'hc1633fdb, 32'hc2562825, 32'h420780f6, 32'hc24a9c0a, 32'hc287d860, 32'h4131400e, 32'h41156d7a, 32'hc1fc60eb};
test_bias[2935:2935] = '{32'hc1717b87};
test_output[2935:2935] = '{32'h462f579b};
test_input[23488:23495] = '{32'h4260f7ee, 32'h42383b84, 32'hc2c45549, 32'h41930c03, 32'h40f9b2d5, 32'h42828752, 32'hc2876782, 32'h417e825d};
test_weights[23488:23495] = '{32'hc2983eaa, 32'h42b7dcd6, 32'h41a3d11c, 32'h42b742e8, 32'hc28a9278, 32'h41dfcb15, 32'h4103fd6a, 32'hc0fef1fe};
test_bias[2936:2936] = '{32'h42704e77};
test_output[2936:2936] = '{32'h438f7303};
test_input[23496:23503] = '{32'h426b4e31, 32'hc2c561f1, 32'hc24c5828, 32'hc28268f3, 32'hc047d3ac, 32'hc0bca804, 32'hc197f1a1, 32'h42a71f85};
test_weights[23496:23503] = '{32'hc2bd7660, 32'hc2770c52, 32'hc20990e5, 32'h42171a5a, 32'hc1f6bafe, 32'hc2ab6d32, 32'hc29a67db, 32'hc231516f};
test_bias[2937:2937] = '{32'h42ab3672};
test_output[2937:2937] = '{32'hc4d8c864};
test_input[23504:23511] = '{32'hc29b95cc, 32'h426cac63, 32'hc23d7084, 32'h428518b0, 32'hc28e8c44, 32'hc2922186, 32'hc2a98703, 32'h4299c019};
test_weights[23504:23511] = '{32'hc28064e6, 32'h42b5b151, 32'hc2c0ffcf, 32'h41103561, 32'h428e6556, 32'hc20b059d, 32'hc29bf74e, 32'h41ebda7a};
test_bias[2938:2938] = '{32'h4242bcbc};
test_output[2938:2938] = '{32'h46ab52c5};
test_input[23512:23519] = '{32'hc1079731, 32'h428ac059, 32'hbfa63ced, 32'hc2839e36, 32'h42655df0, 32'h4260a597, 32'h42921aa9, 32'h42be9c0a};
test_weights[23512:23519] = '{32'h425d4526, 32'hc2615d94, 32'hc2a985f2, 32'h4209d7b2, 32'hc1e226f2, 32'hbfdd6b13, 32'hc1cd06ba, 32'hc141d3ea};
test_bias[2939:2939] = '{32'hbfc929db};
test_output[2939:2939] = '{32'hc63046d0};
test_input[23520:23527] = '{32'hc21d282e, 32'h42674bd8, 32'hc2656911, 32'h3f33b0f5, 32'h428e3c4e, 32'h4269b13d, 32'hc2a75f46, 32'h40359ee4};
test_weights[23520:23527] = '{32'h420e05ac, 32'h404f4018, 32'h4270fbad, 32'h421a45a0, 32'hbfc06a3e, 32'h429d16f4, 32'h4222b007, 32'hc2ba3fbb};
test_bias[2940:2940] = '{32'h425fdb14};
test_output[2940:2940] = '{32'hc56b5f85};
test_input[23528:23535] = '{32'h42117441, 32'h42b33d19, 32'hc2aa0578, 32'h42362687, 32'hc2083972, 32'hc119fabf, 32'hc294711f, 32'h42369693};
test_weights[23528:23535] = '{32'h42afa80e, 32'hc21ee083, 32'hc2a79886, 32'hc1df424f, 32'h426e5817, 32'hc29d11b4, 32'hc1c06158, 32'h419af4b6};
test_bias[2941:2941] = '{32'h42b57f37};
test_output[2941:2941] = '{32'h45d9ea39};
test_input[23536:23543] = '{32'hc20b876a, 32'h421dc0ac, 32'hc2734bc1, 32'h42b7241d, 32'hc246b0ad, 32'h4143aecf, 32'h428de688, 32'h42880420};
test_weights[23536:23543] = '{32'hc21894a7, 32'h4228bbc4, 32'hc27ad1d6, 32'hc292ed34, 32'hc23e4f6f, 32'h424bfa31, 32'hc2c58af8, 32'hc1d30e32};
test_bias[2942:2942] = '{32'h426bc6bb};
test_output[2942:2942] = '{32'hc5b1581f};
test_input[23544:23551] = '{32'h4267190f, 32'hc2440da5, 32'h42c07df3, 32'hc2a0f154, 32'h4282f4e2, 32'hc2515dcc, 32'hc29e5a30, 32'h429c1676};
test_weights[23544:23551] = '{32'h425cf8d0, 32'h41d1b11a, 32'hc0e4b2ee, 32'hc2a9408e, 32'h420738f4, 32'hc2c11a8c, 32'h3fd2eec9, 32'h422e5e34};
test_bias[2943:2943] = '{32'h42c3f48e};
test_output[2943:2943] = '{32'h4691d3b0};
test_input[23552:23559] = '{32'h41afd7b8, 32'hc2a12f35, 32'h427da223, 32'hc2c6334f, 32'hc2b7af2a, 32'hc27e0a8b, 32'hc299c996, 32'h424531e4};
test_weights[23552:23559] = '{32'h42567a2f, 32'h428251f3, 32'hc283e57d, 32'hc292c7ce, 32'hc298dc30, 32'h42bc8f8b, 32'h42889c39, 32'h42887008};
test_bias[2944:2944] = '{32'h42a9c68a};
test_output[2944:2944] = '{32'hc4db40ba};
test_input[23560:23567] = '{32'hc2ab1b21, 32'h42c08413, 32'h4236867e, 32'h41009190, 32'hc215bf1f, 32'hc243108e, 32'h42c7d55f, 32'h42bc4697};
test_weights[23560:23567] = '{32'h4282862e, 32'h42bf9d84, 32'hbffdcbce, 32'hc2194723, 32'h423af8c0, 32'h42a6276b, 32'h425b8082, 32'hc1fc27be};
test_bias[2945:2945] = '{32'hc1a0ccb9};
test_output[2945:2945] = '{32'hc28216be};
test_input[23568:23575] = '{32'h42a1d368, 32'hc2b155c2, 32'hc2bf956d, 32'h42a65928, 32'h429bb6c2, 32'hc28da4a4, 32'h421a44c3, 32'h41abb4e0};
test_weights[23568:23575] = '{32'h42129469, 32'h410789d4, 32'hc2acb1df, 32'hc25f412b, 32'hc1ae9323, 32'hc2b3e5f8, 32'hc004f600, 32'h428ba55f};
test_bias[2946:2946] = '{32'h42bcca34};
test_output[2946:2946] = '{32'h463bed48};
test_input[23576:23583] = '{32'h41b8c375, 32'hc245773e, 32'hc03a78f1, 32'h428bf951, 32'hc2ab5dc4, 32'h4091e82d, 32'h40366f83, 32'h4229dc55};
test_weights[23576:23583] = '{32'h42a95852, 32'h42c422e4, 32'hc2a53959, 32'hc2bbe4ed, 32'hc2a1b00e, 32'hc0ee3df5, 32'h4247c5b5, 32'h42a449e0};
test_bias[2947:2947] = '{32'h416c14d6};
test_output[2947:2947] = '{32'h44a4c9aa};
test_input[23584:23591] = '{32'hc18962d3, 32'h425097e0, 32'h42c356a8, 32'hc24deb48, 32'h41241db6, 32'hc0830530, 32'h3ece0b73, 32'hc23bc762};
test_weights[23584:23591] = '{32'hbfbc3ff7, 32'hc292c44c, 32'h40fb5431, 32'hc2439258, 32'h4215479e, 32'hc17bcc6b, 32'hc2198d78, 32'h428f34b2};
test_bias[2948:2948] = '{32'h420d74c6};
test_output[2948:2948] = '{32'hc5553b2e};
test_input[23592:23599] = '{32'hc29aed5f, 32'h421d4d5a, 32'hc1935929, 32'h42c10e50, 32'h428545c2, 32'hc28c5af0, 32'hc2bbe2ea, 32'h4195b7e3};
test_weights[23592:23599] = '{32'h429bfb02, 32'hc233ae6c, 32'hc1a765d4, 32'h42a66d79, 32'hc292f8db, 32'hc211362e, 32'hc25d1685, 32'h42a91686};
test_bias[2949:2949] = '{32'h41fc6951};
test_output[2949:2949] = '{32'h459e57a9};
test_input[23600:23607] = '{32'hc22a0043, 32'hc2ba102b, 32'hc24a5bf3, 32'h4260eae2, 32'hc29c9760, 32'h416f4fe7, 32'h40e6ac55, 32'h42b18f43};
test_weights[23600:23607] = '{32'h42ac2669, 32'hc1def16a, 32'hc2bb603f, 32'h4279cdc7, 32'hc0a934e8, 32'hc2b4b479, 32'hc2bacb16, 32'hc19e3601};
test_bias[2950:2950] = '{32'hc04bce9c};
test_output[2950:2950] = '{32'h456e809d};
test_input[23608:23615] = '{32'h4296cc00, 32'h4233daa9, 32'hc14f71ec, 32'hc073d896, 32'hc0902175, 32'h424e32fb, 32'hc28688ad, 32'h423fce3a};
test_weights[23608:23615] = '{32'hc1b3db4b, 32'h428642b5, 32'h42ad25e4, 32'h40298713, 32'hc28964ff, 32'hc231dd87, 32'h4141538b, 32'h422f5212};
test_bias[2951:2951] = '{32'hc236e849};
test_output[2951:2951] = '{32'hc409367e};
test_input[23616:23623] = '{32'h4221efb7, 32'h4266cec3, 32'h42825380, 32'h4000b750, 32'h42bf7c58, 32'h41ac123c, 32'h421d5cb5, 32'hc2b7c8af};
test_weights[23616:23623] = '{32'hc1307384, 32'h4255fb1b, 32'hc19033c6, 32'h4218c9ea, 32'hc27da2b6, 32'h41b4b1b1, 32'hc085494d, 32'hc145a2f5};
test_bias[2952:2952] = '{32'hc2869c52};
test_output[2952:2952] = '{32'hc5442acc};
test_input[23624:23631] = '{32'h419838f6, 32'h4278eefa, 32'hc227b992, 32'h4082c214, 32'hc28cfb9a, 32'h42b92f80, 32'hbe90168c, 32'h42880745};
test_weights[23624:23631] = '{32'h42a6f8a5, 32'hc1d57686, 32'hc2a2eed5, 32'h4299909b, 32'h417e454d, 32'hc232e529, 32'h4238d6d2, 32'hc2bf99eb};
test_bias[2953:2953] = '{32'h42a54651};
test_output[2953:2953] = '{32'hc5fb8e58};
test_input[23632:23639] = '{32'h42472919, 32'h4081f531, 32'hc1bd1b28, 32'h42a60e61, 32'hc28eb036, 32'hc1bafbab, 32'hc2947392, 32'h41acad74};
test_weights[23632:23639] = '{32'hbf8d410d, 32'h41ab403d, 32'hc28fe770, 32'h41169719, 32'h42a71b8e, 32'hc08c7bed, 32'h42270f08, 32'hc25bb7a3};
test_bias[2954:2954] = '{32'hc2a80928};
test_output[2954:2954] = '{32'hc5f10ef6};
test_input[23640:23647] = '{32'h42655e7e, 32'h4125af4a, 32'hc09d8f42, 32'hc195edad, 32'hc28eaca6, 32'hc1a2e193, 32'hc25f24f4, 32'hc2ba3055};
test_weights[23640:23647] = '{32'hc245507b, 32'hc2b707de, 32'h422a79b4, 32'hc25c5e48, 32'h429c03cb, 32'hc14d912e, 32'hc2a91a84, 32'hc2b2c719};
test_bias[2955:2955] = '{32'h405bfd2d};
test_output[2955:2955] = '{32'h459587ba};
test_input[23648:23655] = '{32'h41c5d757, 32'h42a510da, 32'h42af866d, 32'h420b1aa0, 32'hc2b930a4, 32'hc23ad2c9, 32'h404e74f7, 32'hc2a92210};
test_weights[23648:23655] = '{32'h42b63dd5, 32'h422333cc, 32'h4279a919, 32'h428be565, 32'hc1c48035, 32'h420a97ab, 32'h41c2024a, 32'h3e7e05fe};
test_bias[2956:2956] = '{32'h417dfa17};
test_output[2956:2956] = '{32'h465ed11c};
test_input[23656:23663] = '{32'hc13ab3b1, 32'hc0b5bfb1, 32'h426f4a3f, 32'h41576d17, 32'h41cb02fa, 32'hc090c32f, 32'h42197577, 32'h426816bf};
test_weights[23656:23663] = '{32'h40cfe275, 32'h42a6af93, 32'hc22a0faa, 32'h42361da3, 32'h423067ed, 32'hc25d5db1, 32'h40bc99f0, 32'hc241bff2};
test_bias[2957:2957] = '{32'hc1592b69};
test_output[2957:2957] = '{32'hc567bf0d};
test_input[23664:23671] = '{32'h42536af3, 32'hc2a86119, 32'h42924317, 32'h4258f5e9, 32'hc2a6d4a0, 32'hc292751f, 32'hc1eb64a6, 32'h4288349d};
test_weights[23664:23671] = '{32'h42a12f2c, 32'h42552ed5, 32'h424ba8d7, 32'h421024a7, 32'h4296b215, 32'h426bee65, 32'h42bd6c17, 32'hc05cadee};
test_bias[2958:2958] = '{32'hc236da5a};
test_output[2958:2958] = '{32'hc60073ed};
test_input[23672:23679] = '{32'h42979d77, 32'hc2c25475, 32'hc1b2863b, 32'h42b59432, 32'hc2108ad3, 32'h41d22bed, 32'h42177f7b, 32'h42177a17};
test_weights[23672:23679] = '{32'h4219460a, 32'hc13c5fa9, 32'hc26fa7b7, 32'hc1ffd3d2, 32'h429958f3, 32'h422eb674, 32'hc1a933c3, 32'hc27a2483};
test_bias[2959:2959] = '{32'h42616486};
test_output[2959:2959] = '{32'hc50cd8f0};
test_input[23680:23687] = '{32'h3f8f554e, 32'hc2b3b7c3, 32'h42c77994, 32'hc28b6ffb, 32'h41db1b15, 32'hc292f315, 32'h4298baf5, 32'hc1750738};
test_weights[23680:23687] = '{32'hc27b93e6, 32'h414a69e4, 32'h41bc3a79, 32'hc1a7e7b0, 32'hc1f66f8a, 32'hc2431df2, 32'h429c78f9, 32'h429c2370};
test_bias[2960:2960] = '{32'h4282e5c9};
test_output[2960:2960] = '{32'h461f2df4};
test_input[23688:23695] = '{32'h42a731a6, 32'h411bf22e, 32'hc1af0cac, 32'hc2561323, 32'hc024a408, 32'hc1cd6675, 32'h42163ba6, 32'h411e71d8};
test_weights[23688:23695] = '{32'hc2816a06, 32'h41e1251b, 32'hc26d4fb2, 32'hc22826f5, 32'h42be573e, 32'hc26fd8f7, 32'hc2bf20a7, 32'h413db05e};
test_bias[2961:2961] = '{32'hc2c0e1fb};
test_output[2961:2961] = '{32'hc571494c};
test_input[23696:23703] = '{32'h40a4f6b1, 32'h424d6d1c, 32'hc1f373f7, 32'hc27df605, 32'h42a222fb, 32'hc295c14e, 32'h42abab86, 32'h42c7dc60};
test_weights[23696:23703] = '{32'hc2655c37, 32'hc299d079, 32'hc1e361f2, 32'hc0c2e411, 32'hc253f9bc, 32'hc23ee256, 32'hc2257a8b, 32'h41c7418f};
test_bias[2962:2962] = '{32'hc1299d3b};
test_output[2962:2962] = '{32'hc595a922};
test_input[23704:23711] = '{32'h425f148a, 32'h418dae3a, 32'hc268e816, 32'h428b547b, 32'h42954363, 32'h4142dd5d, 32'h4174404e, 32'h42b4a7fa};
test_weights[23704:23711] = '{32'hc17d24cf, 32'hc188fd09, 32'hc1537f23, 32'h42388788, 32'hc29bf3b0, 32'h4293e0cb, 32'hc1656156, 32'hc2c6b56c};
test_bias[2963:2963] = '{32'hc2137e9c};
test_output[2963:2963] = '{32'hc6315d49};
test_input[23712:23719] = '{32'hc1722bdc, 32'h423c7a18, 32'hc2c1ea91, 32'hc003121c, 32'hc27feb10, 32'h41be6daf, 32'h41178e3b, 32'hc2aa01d4};
test_weights[23712:23719] = '{32'h4158c56a, 32'hc28e03b3, 32'h4143eab5, 32'hc296b19b, 32'hc269e571, 32'h41f9562e, 32'h4268d3d4, 32'h4229d27a};
test_bias[2964:2964] = '{32'hc28acfbc};
test_output[2964:2964] = '{32'hc549bb0a};
test_input[23720:23727] = '{32'hc2b7c9d1, 32'h41cef631, 32'hc268b011, 32'h42bc1ca1, 32'h4221fb70, 32'hc2832aa2, 32'hc2999cbf, 32'hc28762a7};
test_weights[23720:23727] = '{32'hc26f7754, 32'hc1d70e3c, 32'hc2aede61, 32'hbf74184f, 32'hc2b85f26, 32'h42057023, 32'hc2b82875, 32'h4210130b};
test_bias[2965:2965] = '{32'h42c73c57};
test_output[2965:2965] = '{32'h46069ccf};
test_input[23728:23735] = '{32'h40f3f360, 32'h41abca46, 32'h42bae758, 32'h429c201a, 32'hc1c1e826, 32'h424ed473, 32'h429e0c2a, 32'hc204584a};
test_weights[23728:23735] = '{32'h40ce532a, 32'hc2a93d29, 32'h42bd8284, 32'h41bf92ae, 32'h40aad7e2, 32'h42c37c1b, 32'hc2a7c486, 32'h42afd227};
test_bias[2966:2966] = '{32'hc27c1595};
test_output[2966:2966] = '{32'h4585c47a};
test_input[23736:23743] = '{32'hc2706a00, 32'hc18da199, 32'h421573c8, 32'hc23dd6c1, 32'hc27aaf00, 32'h4289172b, 32'hc2c368aa, 32'h4297a561};
test_weights[23736:23743] = '{32'hc2acf44b, 32'hc2427bce, 32'hc26cded2, 32'h41578f33, 32'h41ade3dc, 32'h41e0495f, 32'h4204893a, 32'hc0f37ac9};
test_bias[2967:2967] = '{32'hc2846b40};
test_output[2967:2967] = '{32'hc2e5215f};
test_input[23744:23751] = '{32'h42b39bfa, 32'hbf43521c, 32'h42898aed, 32'hc103c472, 32'h427fb81d, 32'h4098e0fc, 32'h421268eb, 32'hbf893e1c};
test_weights[23744:23751] = '{32'hc113e195, 32'hc27313b5, 32'h42b6c94b, 32'h42c0ac68, 32'hc29c0c05, 32'h42aefd1b, 32'hc22be673, 32'h42b49072};
test_bias[2968:2968] = '{32'hc1f14cb8};
test_output[2968:2968] = '{32'hc4c3393e};
test_input[23752:23759] = '{32'h4294b5d5, 32'hc241221e, 32'hc2692f28, 32'h41ab09b0, 32'hc1a64980, 32'h428c62e4, 32'hc14b596d, 32'h4141c629};
test_weights[23752:23759] = '{32'hc0466bed, 32'hc2963897, 32'h429387a6, 32'h4276ae0e, 32'hc28f42be, 32'hc284f55f, 32'h42611412, 32'hc2527ea9};
test_bias[2969:2969] = '{32'hc21d5b67};
test_output[2969:2969] = '{32'hc581d79d};
test_input[23760:23767] = '{32'h41e78492, 32'h4240c2f2, 32'hc260413b, 32'h42bd72dc, 32'hc2c03b7b, 32'h424782dd, 32'hc1abb57b, 32'h422d07c8};
test_weights[23760:23767] = '{32'h411e0cb3, 32'hc24610e8, 32'h42c62806, 32'hc268a208, 32'h420d576c, 32'hc18ff0a5, 32'h429f11be, 32'hc11644ff};
test_bias[2970:2970] = '{32'hc2212aea};
test_output[2970:2970] = '{32'hc69936db};
test_input[23768:23775] = '{32'hc2c0391f, 32'h4106657a, 32'hc22f9a18, 32'hc1c47608, 32'hc2c3b1c5, 32'h42955f47, 32'h424a4438, 32'h41a319a4};
test_weights[23768:23775] = '{32'h42a46537, 32'hc213df30, 32'hc1d01f03, 32'h422a9cad, 32'hc28e0224, 32'hc13e0d6d, 32'hc1a45de6, 32'h4184afb4};
test_bias[2971:2971] = '{32'h41b47d6a};
test_output[2971:2971] = '{32'hc52addc6};
test_input[23776:23783] = '{32'h42609682, 32'h4226888e, 32'h4109a66f, 32'h42149aa7, 32'hc13bb3ab, 32'hc2bb2fb6, 32'hc274ab3a, 32'hc1a62232};
test_weights[23776:23783] = '{32'h42a1f455, 32'h42b464e1, 32'hc26774f7, 32'h42a25091, 32'hc199c6eb, 32'hc18fb582, 32'hc275e8c5, 32'h424d14e1};
test_bias[2972:2972] = '{32'hc26aa4b5};
test_output[2972:2972] = '{32'h46700b8f};
test_input[23784:23791] = '{32'h42486547, 32'hc2b96e9d, 32'hc2a29d32, 32'h42a216ef, 32'hc1829950, 32'hc25168ae, 32'hc218a791, 32'hc2b250da};
test_weights[23784:23791] = '{32'hc22636be, 32'hc1903e5f, 32'hc246c65e, 32'hc25a50de, 32'hc28d9e95, 32'hc123a87f, 32'hc2826dee, 32'h4003d8fe};
test_bias[2973:2973] = '{32'h428b19f6};
test_output[2973:2973] = '{32'h454c9314};
test_input[23792:23799] = '{32'h41b4ca78, 32'h4208c0ac, 32'hc2c79dc4, 32'hc26703f9, 32'hc20131cc, 32'hc15a88f2, 32'h42c7d1b8, 32'h42414bc6};
test_weights[23792:23799] = '{32'h42170699, 32'hc2321cf5, 32'hc1c74099, 32'h428531bd, 32'h420818a4, 32'h40884c59, 32'hc18ad82c, 32'hc23938ab};
test_bias[2974:2974] = '{32'hc16d3a7a};
test_output[2974:2974] = '{32'hc5e02846};
test_input[23800:23807] = '{32'h42c50def, 32'h4242b92a, 32'h41bdb897, 32'hc28330a2, 32'h3fe90c88, 32'h42326b7a, 32'hc289f698, 32'hc29d2d34};
test_weights[23800:23807] = '{32'hc24d0f12, 32'hc2a88eca, 32'hc27683d5, 32'hc29dc4e2, 32'hc2c1b9a3, 32'h416a8b35, 32'h41075e69, 32'h42a07565};
test_bias[2975:2975] = '{32'h416c60ff};
test_output[2975:2975] = '{32'hc638f50e};
test_input[23808:23815] = '{32'h4291dd89, 32'h4123e1ab, 32'hc29ce1f1, 32'h42bfcaed, 32'hc2245da4, 32'hc20556c9, 32'h428c055c, 32'hc27961d9};
test_weights[23808:23815] = '{32'h4238e654, 32'hc17f2d44, 32'hc25752ca, 32'hc2a9de92, 32'hc2340338, 32'h42b0a3ed, 32'hc042a789, 32'hc242c27b};
test_bias[2976:2976] = '{32'hc29be5bf};
test_output[2976:2976] = '{32'h4469daa8};
test_input[23816:23823] = '{32'h427b255b, 32'hc282b0c4, 32'hc268b8ef, 32'hc2a478ef, 32'hc2c675be, 32'h42c75008, 32'hc2c6ee11, 32'hc204e597};
test_weights[23816:23823] = '{32'h4243d7c6, 32'hc24a3721, 32'hc212c5ce, 32'hc26d2e2b, 32'hc2a745e8, 32'hc24755f5, 32'hc2c47a10, 32'hc1a053a6};
test_bias[2977:2977] = '{32'h42c0852e};
test_output[2977:2977] = '{32'h46d4edd8};
test_input[23824:23831] = '{32'hc2005b13, 32'hc221ae7c, 32'hc2c489ff, 32'h41c3b2d1, 32'hc0724053, 32'hc27d2b03, 32'hbeee2b5e, 32'h42abf77d};
test_weights[23824:23831] = '{32'hc23d189f, 32'hc2b98013, 32'h42b28d12, 32'h408c849c, 32'hc28271c1, 32'hc2bf0f6a, 32'hc24730d9, 32'hc2a09d1d};
test_bias[2978:2978] = '{32'hc265c399};
test_output[2978:2978] = '{32'hc57cdd60};
test_input[23832:23839] = '{32'h423f6808, 32'h4206e9ac, 32'hc297f555, 32'h4154907a, 32'h428ea1a4, 32'h42892786, 32'hc29717e4, 32'h426602ce};
test_weights[23832:23839] = '{32'h413bdd84, 32'h42977273, 32'h4284ea30, 32'h429a2f16, 32'hc1bab1c3, 32'h41e6dc29, 32'h428c1a08, 32'h4285a271};
test_bias[2979:2979] = '{32'h41a4cf8d};
test_output[2979:2979] = '{32'hc4fcfec9};
test_input[23840:23847] = '{32'hc1ff9d0d, 32'h42862fc4, 32'h4220379b, 32'hc24d4b6c, 32'hbf869eb3, 32'h421d6e78, 32'hc0fbbaff, 32'h425f126b};
test_weights[23840:23847] = '{32'hc28c2e5a, 32'h4286ab70, 32'h428f20b8, 32'hc26e6c26, 32'h40d4b573, 32'h42a532af, 32'h42a7c067, 32'hc276024f};
test_bias[2980:2980] = '{32'h428d2173};
test_output[2980:2980] = '{32'h463a0eae};
test_input[23848:23855] = '{32'hc23a7d1f, 32'hc2be4f49, 32'hc2b70873, 32'hc2b460cb, 32'h41f99edf, 32'hc11598ef, 32'h420be5fe, 32'hc1da00f1};
test_weights[23848:23855] = '{32'h42093670, 32'hc2688673, 32'h410121a8, 32'hc21e95c8, 32'hc2b059c9, 32'h42853a54, 32'h42b68378, 32'hc0b6e252};
test_bias[2981:2981] = '{32'hc0479978};
test_output[2981:2981] = '{32'h45d29b3e};
test_input[23856:23863] = '{32'hc190b3b4, 32'h424871b6, 32'h4281584e, 32'hc2855a60, 32'h412ad606, 32'hc285b2dd, 32'hc2b4b30a, 32'hc0b5b73c};
test_weights[23856:23863] = '{32'h4209154a, 32'hc1cd9782, 32'h42b73315, 32'h3f5c93dc, 32'hc285ad85, 32'h421db802, 32'h421b8d3b, 32'h41a46f15};
test_bias[2982:2982] = '{32'hc1ecf24f};
test_output[2982:2982] = '{32'hc53ea816};
test_input[23864:23871] = '{32'hc206d780, 32'h4290fe88, 32'h42ab3810, 32'hc2780e72, 32'hc23ba81c, 32'h4250c58a, 32'hc2392b04, 32'hc18dda43};
test_weights[23864:23871] = '{32'h420ca847, 32'h41dec3db, 32'hc2b258cf, 32'hc15e72e6, 32'h41de0746, 32'hc2bd0242, 32'h41a37115, 32'h429c5e7f};
test_bias[2983:2983] = '{32'h42150dc1};
test_output[2983:2983] = '{32'hc6620fa3};
test_input[23872:23879] = '{32'h42a859ac, 32'h4213b7b3, 32'h422d607a, 32'hc2b564bf, 32'h41cc7aa5, 32'h42a73665, 32'hc2a11c4a, 32'h4282ad68};
test_weights[23872:23879] = '{32'hc23ade82, 32'hc24a696d, 32'h42328194, 32'h42b23cfa, 32'hc2a1d900, 32'h429a387d, 32'hc24e96c8, 32'hc2b13904};
test_bias[2984:2984] = '{32'h416071fc};
test_output[2984:2984] = '{32'hc60f89c9};
test_input[23880:23887] = '{32'hc2b49338, 32'h42987589, 32'h41d6ac41, 32'h428e51a8, 32'h421c9d76, 32'h4296e85f, 32'hc2886352, 32'h414fa35c};
test_weights[23880:23887] = '{32'hc10b1943, 32'hc2b5cec3, 32'h42a132b2, 32'h429d4bda, 32'hc14a175f, 32'hc2004e86, 32'hc2ae757f, 32'hc204f96a};
test_bias[2985:2985] = '{32'hc2ae459b};
test_output[2985:2985] = '{32'h45810ee6};
test_input[23888:23895] = '{32'hc26a4f15, 32'h41aabcf2, 32'hc0f08c62, 32'hc26265eb, 32'h42c618a3, 32'hc2c35be7, 32'h42ada818, 32'hc28b9181};
test_weights[23888:23895] = '{32'hc2969085, 32'h42b1f513, 32'hc11e4ec5, 32'hc2a4d25d, 32'h4282c3bd, 32'h3fbc5834, 32'hc291568f, 32'hc2b9de57};
test_bias[2986:2986] = '{32'h3fc14062};
test_output[2986:2986] = '{32'h46892a04};
test_input[23896:23903] = '{32'h42bcbefe, 32'hc2aa788f, 32'h42897df2, 32'hc227d1fe, 32'hc2b15b2a, 32'h41f69169, 32'hc28932e8, 32'hc2a99ce4};
test_weights[23896:23903] = '{32'hc16d03f3, 32'h42a7f14f, 32'hc2030d00, 32'h42c248b1, 32'hc24f0d9f, 32'hc2af9376, 32'h42b5a698, 32'h421d5314};
test_bias[2987:2987] = '{32'hc2abf085};
test_output[2987:2987] = '{32'hc6b0f57d};
test_input[23904:23911] = '{32'hc2097759, 32'hc1d3e1a1, 32'hc1d171fe, 32'hc0baebbb, 32'hc2659087, 32'h42893b46, 32'hc1739c30, 32'hc299149e};
test_weights[23904:23911] = '{32'h4299b9b7, 32'hc2afa402, 32'hc2a98832, 32'hc1951e20, 32'hc206e694, 32'h3eb0ca04, 32'h42ba9f63, 32'hc1d8a567};
test_bias[2988:2988] = '{32'h41736be8};
test_output[2988:2988] = '{32'h4590f823};
test_input[23912:23919] = '{32'h429d201b, 32'hc2777afc, 32'hc2a04279, 32'h41a3ff05, 32'h4231b69e, 32'hc28cd520, 32'hc2b5d307, 32'hc2a29e2c};
test_weights[23912:23919] = '{32'hc1bedfc8, 32'h41589801, 32'h4282f43c, 32'h42693605, 32'hc2b266b1, 32'h42b753c3, 32'h42277e3d, 32'hc0fd6702};
test_bias[2989:2989] = '{32'hc2206951};
test_output[2989:2989] = '{32'hc69f4047};
test_input[23920:23927] = '{32'h42609159, 32'h42c050d7, 32'hc20119bc, 32'h42a880c5, 32'hc1c7185c, 32'h42a6d3a0, 32'hc1d86713, 32'h4288976e};
test_weights[23920:23927] = '{32'hc277acb8, 32'hc1163475, 32'hc2819597, 32'h40ff42f1, 32'h427f7d93, 32'hc20c9645, 32'hc25ae983, 32'h41f1c808};
test_bias[2990:2990] = '{32'h429a9cdf};
test_output[2990:2990] = '{32'hc51d3341};
test_input[23928:23935] = '{32'hc236b7a4, 32'h414c864a, 32'hc2a9a823, 32'hc2567cc6, 32'hc1520c45, 32'h412e8378, 32'h4274924a, 32'hbffe12c8};
test_weights[23928:23935] = '{32'hc255b228, 32'h42162072, 32'h4150f674, 32'hc200ceee, 32'h4277706d, 32'hc236550e, 32'hc1e370bf, 32'h40838b43};
test_bias[2991:2991] = '{32'h42b1dcde};
test_output[2991:2991] = '{32'h440f0c98};
test_input[23936:23943] = '{32'h4295658c, 32'hc29b70ed, 32'h42c0fad5, 32'h41d94ef4, 32'h42bcb668, 32'h4211f4e9, 32'hc19ce325, 32'h41949514};
test_weights[23936:23943] = '{32'h4171052d, 32'h429dae29, 32'h424bbc09, 32'h42bc39bd, 32'h41edcd94, 32'hbdb1f95c, 32'hc2c5f7fb, 32'hc2888ec4};
test_bias[2992:2992] = '{32'hc2b5608f};
test_output[2992:2992] = '{32'h45b6e5b9};
test_input[23944:23951] = '{32'h41f94ab3, 32'hc274c084, 32'hc2583014, 32'hc248d44e, 32'hc2babfbb, 32'h424d9a62, 32'h41dde72a, 32'hc06002b1};
test_weights[23944:23951] = '{32'h426fd781, 32'hc18f82b7, 32'h425735bf, 32'hc127cd71, 32'h42b8ed7f, 32'hc192671e, 32'hc0616d1d, 32'hc293cc1b};
test_bias[2993:2993] = '{32'hc1f8dcfc};
test_output[2993:2993] = '{32'hc60a6f19};
test_input[23952:23959] = '{32'h42894ef8, 32'hc1070339, 32'hc1e9d91e, 32'h4113293c, 32'h41e2e3f9, 32'hc2b47322, 32'h42050763, 32'hc2a5eb63};
test_weights[23952:23959] = '{32'h4281ee5c, 32'h42ac7a2a, 32'h4282f1c4, 32'h428eef93, 32'hc28f07ac, 32'h419e509c, 32'h42816ccd, 32'h426d9831};
test_bias[2994:2994] = '{32'hc2705077};
test_output[2994:2994] = '{32'hc5826b34};
test_input[23960:23967] = '{32'h42c6ab26, 32'hc2289334, 32'h42623d43, 32'hc2bda196, 32'h3e8e5d3a, 32'hbf1aa0e5, 32'hc23b9aa6, 32'h42b06e3f};
test_weights[23960:23967] = '{32'h424103b9, 32'hc2c14b43, 32'hc18b9a21, 32'h42c30e2c, 32'h42740166, 32'h409b9af9, 32'h4275e523, 32'hc17bb33e};
test_bias[2995:2995] = '{32'hc2acc6fc};
test_output[2995:2995] = '{32'hc5b278da};
test_input[23968:23975] = '{32'hc2581b13, 32'h42aa676d, 32'h42946456, 32'h4079ec89, 32'h4232cbae, 32'h41c9d3ce, 32'hc22b2db8, 32'hc28ee563};
test_weights[23968:23975] = '{32'h42bdf0a1, 32'hc2b37e0d, 32'hc1f7493c, 32'h42811b8b, 32'h420a538f, 32'hc2a5bff0, 32'hc2b7ac79, 32'hc1e4b38c};
test_bias[2996:2996] = '{32'h40de08f0};
test_output[2996:2996] = '{32'hc612a108};
test_input[23976:23983] = '{32'h42b36770, 32'h42bcc351, 32'hc299453f, 32'hc25269cf, 32'h42b590dc, 32'h42b986aa, 32'hc1e5d049, 32'hc20ac918};
test_weights[23976:23983] = '{32'h42822275, 32'h42817f75, 32'hc219dbef, 32'hc25c5802, 32'h42a6e41c, 32'h42394cbf, 32'hc0ff38e9, 32'h42bcb895};
test_bias[2997:2997] = '{32'hc27f35c1};
test_output[2997:2997] = '{32'h46cf7a7e};
test_input[23984:23991] = '{32'h42861267, 32'h4289c18c, 32'h42901013, 32'h42b4471c, 32'h429b1257, 32'h418c5d60, 32'h429be221, 32'hc2c053b2};
test_weights[23984:23991] = '{32'hc2310e53, 32'h42b67fc3, 32'hc15a943e, 32'h42b0b769, 32'h425c757e, 32'h42606b6f, 32'h42b67759, 32'h42af458d};
test_bias[2998:2998] = '{32'hc26eb8e9};
test_output[2998:2998] = '{32'h465d8f71};
test_input[23992:23999] = '{32'h427f5bc0, 32'h4240a4ca, 32'hc2bbd92d, 32'h424bcfde, 32'h42196ffe, 32'h425129b8, 32'h4286204d, 32'hc2a3d6c5};
test_weights[23992:23999] = '{32'h402b3d9e, 32'hc23dcc08, 32'h42b87283, 32'h42ac23ef, 32'h42a1a14c, 32'h41e0e64c, 32'h42956fa9, 32'h42033f89};
test_bias[2999:2999] = '{32'h42121e77};
test_output[2999:2999] = '{32'h4406a3bd};
test_input[24000:24007] = '{32'hc16447be, 32'h40e9cb31, 32'h4272375c, 32'h40a0e68d, 32'hc27cc403, 32'h42baabef, 32'hc0cb3ba8, 32'hc2c6c2b8};
test_weights[24000:24007] = '{32'h42c43a4d, 32'h4006fe49, 32'hc2b5e4fd, 32'h428512ff, 32'hc258a1a2, 32'hc205a373, 32'hc2653f6d, 32'h4295e046};
test_bias[3000:3000] = '{32'h40a48e17};
test_output[3000:3000] = '{32'hc6504d55};
test_input[24008:24015] = '{32'h40845333, 32'h42b16631, 32'hc27b1a8f, 32'h426d3f00, 32'h42919802, 32'h4267603a, 32'hc2a79504, 32'hc28a82a6};
test_weights[24008:24015] = '{32'h419306e9, 32'hc01e14ca, 32'h42b4c407, 32'h42af56dc, 32'hc29bdf5f, 32'hc286d655, 32'h42af1c1c, 32'h421fa2c5};
test_bias[3001:3001] = '{32'h4278ba07};
test_output[3001:3001] = '{32'hc69e08ea};
test_input[24016:24023] = '{32'hc28b4d72, 32'h40440d7f, 32'hc26ca7eb, 32'h42b5c84c, 32'h40fedb48, 32'h420718c8, 32'hc1ee661b, 32'h4287d9e1};
test_weights[24016:24023] = '{32'hc0c3f93b, 32'hc26f2a50, 32'h42874775, 32'hc1bef96f, 32'h42944116, 32'hc2885020, 32'h41ad400d, 32'hc288d0ea};
test_bias[3002:3002] = '{32'h4286cede};
test_output[3002:3002] = '{32'hc6490153};
test_input[24024:24031] = '{32'h425c0a9c, 32'hc276ae73, 32'h42066f98, 32'h42c6836c, 32'h42c36d77, 32'hc2290d84, 32'hc2b71bf5, 32'h42ba76f2};
test_weights[24024:24031] = '{32'h41abe0ac, 32'hc2723ca5, 32'hc2887a36, 32'h42859fcf, 32'h42140a0d, 32'h42ac2a17, 32'h42461b1b, 32'h422694dc};
test_bias[3003:3003] = '{32'hc20568d1};
test_output[3003:3003] = '{32'h46058fbc};
test_input[24032:24039] = '{32'hc2ad086e, 32'hc2ae4901, 32'h41c92742, 32'hc203f508, 32'h4285f048, 32'hc1fcaede, 32'h409a5b9a, 32'h41a47744};
test_weights[24032:24039] = '{32'hc1f44cbb, 32'hc21704a4, 32'h42b9732c, 32'hc0cc59c5, 32'hc18d697c, 32'h41c3ef67, 32'h42bfa9ff, 32'hc2280570};
test_bias[3004:3004] = '{32'hc19b8495};
test_output[3004:3004] = '{32'h45be80a5};
test_input[24040:24047] = '{32'h428994dd, 32'hc243f2d8, 32'h42388baa, 32'h4251b41c, 32'h42b2470c, 32'h42615338, 32'hc0f03430, 32'h428fe5c4};
test_weights[24040:24047] = '{32'hc28e7820, 32'h423ada94, 32'h426f7aac, 32'hc2c5c7f0, 32'hc2b5493f, 32'h4257ebf1, 32'h42c56e05, 32'hc24dc477};
test_bias[3005:3005] = '{32'hc1c935c4};
test_output[3005:3005] = '{32'hc6955a77};
test_input[24048:24055] = '{32'hc283f2f3, 32'h42a9b660, 32'hc023fdac, 32'h42797c5c, 32'h42c1a7d6, 32'hc2011193, 32'h426af59e, 32'h4255299d};
test_weights[24048:24055] = '{32'hc282e194, 32'hc25d7817, 32'hc28c2674, 32'h425a999e, 32'hc212284a, 32'hc1839ef7, 32'hc25857ac, 32'h424f5660};
test_bias[3006:3006] = '{32'h414d3e1a};
test_output[3006:3006] = '{32'hc349b3cc};
test_input[24056:24063] = '{32'h42a26243, 32'h429921ce, 32'h428005f2, 32'h428a93c3, 32'h42bc1bb5, 32'h4254200c, 32'hc25bc254, 32'h4239ca15};
test_weights[24056:24063] = '{32'hc24a265f, 32'h426f502e, 32'hc2aa7698, 32'hc1ab4542, 32'hc2353bc2, 32'hc0bc11e6, 32'h420d6e6b, 32'h42b6ea5f};
test_bias[3007:3007] = '{32'h42bf2248};
test_output[3007:3007] = '{32'hc606e6fd};
test_input[24064:24071] = '{32'hc22412df, 32'hc2a2848c, 32'hc2551fd3, 32'hc2c775fb, 32'h40e8c35e, 32'h4284d05a, 32'h4291434d, 32'hc02fb433};
test_weights[24064:24071] = '{32'h4209e185, 32'hc17a144a, 32'h42a0e5cd, 32'hc1677d60, 32'h41a729ef, 32'hc2138bb5, 32'h42735257, 32'h4186f587};
test_bias[3008:3008] = '{32'h42491989};
test_output[3008:3008] = '{32'hc457ac7e};
test_input[24072:24079] = '{32'h417005e3, 32'hc25913cb, 32'hc1413ce1, 32'hc27dfaff, 32'hc2c134bd, 32'h41467e4e, 32'h41f08fe4, 32'h429733dc};
test_weights[24072:24079] = '{32'hc22710f2, 32'hc19899d9, 32'hc28e0175, 32'hc2c3a0f1, 32'h41f59fec, 32'hc29dd414, 32'hc29e9b57, 32'h42135f07};
test_bias[3009:3009] = '{32'hc2b3e927};
test_output[3009:3009] = '{32'h457029f4};
test_input[24080:24087] = '{32'hc115c8ec, 32'h42b8af02, 32'h42867334, 32'hc257f03f, 32'hc184a36c, 32'h42541dca, 32'hc105f686, 32'h42b8d8fa};
test_weights[24080:24087] = '{32'h420e8e00, 32'hc283c932, 32'hc28dd2d9, 32'h4249da4b, 32'h42b763af, 32'hc168a9b4, 32'h421b60cf, 32'h423d0b4c};
test_bias[3010:3010] = '{32'hc1c000b3};
test_output[3010:3010] = '{32'hc63e58b7};
test_input[24088:24095] = '{32'h42887599, 32'hc2b28df3, 32'hbdec343b, 32'h42910589, 32'hc26af757, 32'h425a849d, 32'h420b9834, 32'hc1871157};
test_weights[24088:24095] = '{32'h424f4371, 32'hc285cb59, 32'hc29d7bcb, 32'h41433122, 32'hc1a03205, 32'hc2acca3f, 32'h427a908b, 32'h421ac222};
test_bias[3011:3011] = '{32'hc2ababe0};
test_output[3011:3011] = '{32'h4601c42a};
test_input[24096:24103] = '{32'h42b61210, 32'hc20dc952, 32'h42ae5e08, 32'h427ba5e9, 32'hc29cfade, 32'hc265de9a, 32'hc29eee94, 32'hc241e349};
test_weights[24096:24103] = '{32'h40ea051e, 32'h425443ac, 32'hc245682b, 32'hc265adc5, 32'hc27fcdb4, 32'h42811bfc, 32'hc1f99cb2, 32'hc2aa0f8a};
test_bias[3012:3012] = '{32'h426e26e3};
test_output[3012:3012] = '{32'hc4910068};
test_input[24104:24111] = '{32'h41797c29, 32'hc24b29b4, 32'hc2835161, 32'h41969a86, 32'h41195811, 32'hc2455cb3, 32'hbe576762, 32'hc2369adc};
test_weights[24104:24111] = '{32'hc2ab6a2d, 32'h4282b753, 32'hc2a15c66, 32'h42c07568, 32'hc1b35b29, 32'hc26c0da4, 32'hc2930f6b, 32'hc0f6e4c5};
test_bias[3013:3013] = '{32'h4261edaf};
test_output[3013:3013] = '{32'h45ae3000};
test_input[24112:24119] = '{32'hc2996af5, 32'hc246d872, 32'hc22e3bcb, 32'hc219d89a, 32'h418ecf4c, 32'h41aea40b, 32'hc1874d59, 32'hc2c14c08};
test_weights[24112:24119] = '{32'hc1fc5a69, 32'hc2458bb3, 32'hbdf6b8fb, 32'hc2a2ca02, 32'h4284c093, 32'hc289b3c1, 32'hc22a5596, 32'h4255193d};
test_bias[3014:3014] = '{32'hc198161a};
test_output[3014:3014] = '{32'h454acbd4};
test_input[24120:24127] = '{32'h418732c2, 32'hc2c64f16, 32'h41d87412, 32'hc21105ef, 32'hc29db231, 32'h424cc950, 32'hc282ea01, 32'h427a2e9e};
test_weights[24120:24127] = '{32'h42057cac, 32'h4143d8cd, 32'hc20d2ff4, 32'h4215041e, 32'hc296f2ae, 32'h41f46fa6, 32'hc2ab896d, 32'h42c25800};
test_bias[3015:3015] = '{32'hc0a4472a};
test_output[3015:3015] = '{32'h467dda22};
test_input[24128:24135] = '{32'hc2c4b027, 32'hc2a66bd0, 32'h428c507f, 32'hc2aa83bf, 32'hc25a296c, 32'hc294acdd, 32'hc2b27ec9, 32'h4295d2fd};
test_weights[24128:24135] = '{32'hc295752c, 32'hc1780a5b, 32'h4274cf05, 32'h422f05c3, 32'h42761db9, 32'hc2a65efc, 32'h41b678f7, 32'hc14cd8ae};
test_bias[3016:3016] = '{32'hc1031da8};
test_output[3016:3016] = '{32'h460d0dcc};
test_input[24136:24143] = '{32'h42c2ba38, 32'h418e677f, 32'h423b1451, 32'hc2c58b80, 32'h412bd6ca, 32'h42b5687a, 32'hc2b89238, 32'hc238fa4f};
test_weights[24136:24143] = '{32'hc2800821, 32'h4266a56e, 32'h42c45a1c, 32'h41db2efd, 32'hc2203600, 32'hc14fde98, 32'hc2092df7, 32'h40b055b9};
test_bias[3017:3017] = '{32'h421df649};
test_output[3017:3017] = '{32'hc4f77c9e};
test_input[24144:24151] = '{32'hc2af66ca, 32'hc28e85a4, 32'h429a0772, 32'h4277eeae, 32'h428673bf, 32'hc25a5657, 32'h41e19887, 32'h4257426b};
test_weights[24144:24151] = '{32'hbff08345, 32'hc20bc9c9, 32'hc2aef5ae, 32'hc219c006, 32'h422ad55a, 32'h426e892e, 32'h42018e14, 32'h4236f203};
test_bias[3018:3018] = '{32'hc262c93c};
test_output[3018:3018] = '{32'hc55ca905};
test_input[24152:24159] = '{32'h42872c45, 32'hc2b8849d, 32'h428316f1, 32'hc2806335, 32'hc1e90fcd, 32'hc2ac1a37, 32'hc1c7db11, 32'h413eed1c};
test_weights[24152:24159] = '{32'h4202e665, 32'hc2203d31, 32'h42b1cd7e, 32'hc1514bda, 32'h42c3ef80, 32'hc00af107, 32'h4225d48c, 32'h42497cf4};
test_bias[3019:3019] = '{32'hc29d0e5b};
test_output[3019:3019] = '{32'h4612c7f9};
test_input[24160:24167] = '{32'h422fe7ab, 32'hc2841999, 32'hc0854935, 32'h4253d2b0, 32'hc2971665, 32'hc16d1cc0, 32'hc29547e8, 32'h41a6075b};
test_weights[24160:24167] = '{32'h42916cd1, 32'h423f8754, 32'hc2a92116, 32'h40716edc, 32'h41d4afb4, 32'h41e3025a, 32'hc2b18109, 32'hc2422d9f};
test_bias[3020:3020] = '{32'hc2843865};
test_output[3020:3020] = '{32'h4567cffe};
test_input[24168:24175] = '{32'hc229147b, 32'h4120ca4e, 32'hc168d223, 32'h4109676f, 32'h41d162c3, 32'hc2972757, 32'hc28db43b, 32'h422440a8};
test_weights[24168:24175] = '{32'h42b1f697, 32'hc23e569a, 32'hc29c8e28, 32'hc1ff3e38, 32'hc2a80205, 32'h42874d25, 32'hc1aeaf1c, 32'hc2311a1c};
test_bias[3021:3021] = '{32'hc1ce72bf};
test_output[3021:3021] = '{32'hc62b9ac1};
test_input[24176:24183] = '{32'hc21da294, 32'h410973c2, 32'h4046539f, 32'h42bbb0d8, 32'hc1b690ae, 32'h414e5361, 32'hc2707655, 32'h3e8e19f0};
test_weights[24176:24183] = '{32'h4292da0e, 32'h429c4874, 32'h42409b28, 32'h416c603b, 32'h423238ca, 32'h42b017a0, 32'h4247dc33, 32'hc219e812};
test_bias[3022:3022] = '{32'hc2b82d38};
test_output[3022:3022] = '{32'hc565a87e};
test_input[24184:24191] = '{32'hc25c4fe0, 32'hc0b51b7a, 32'hc245e024, 32'hc1a7653c, 32'h429ab459, 32'h4124f9e0, 32'h42b892f2, 32'hc296893c};
test_weights[24184:24191] = '{32'h424c4574, 32'h40d7bd69, 32'h4288712d, 32'h4224b36b, 32'h4167a448, 32'hc244df3c, 32'hc26afec2, 32'hc2354e86};
test_bias[3023:3023] = '{32'h4215d422};
test_output[3023:3023] = '{32'hc603fe0a};
test_input[24192:24199] = '{32'h42c308b3, 32'hc128e4be, 32'hc28d3174, 32'hc259a34e, 32'h415f91a0, 32'h428b1ff4, 32'h402f190a, 32'hc15827fb};
test_weights[24192:24199] = '{32'hc294e31d, 32'h41fbc0f1, 32'hc19599f4, 32'hc231fb50, 32'hc22e0e1d, 32'hc28f9f57, 32'hc231b577, 32'h422512da};
test_bias[3024:3024] = '{32'hc224d826};
test_output[3024:3024] = '{32'hc61ef8e6};
test_input[24200:24207] = '{32'hc2ac2640, 32'hc187cb3b, 32'hc24aa81b, 32'hc14cf841, 32'h42914ba8, 32'h427eefb2, 32'h4284e208, 32'hc18f1eb7};
test_weights[24200:24207] = '{32'hc2a5a3fe, 32'hc186667f, 32'hc296c62c, 32'h40874097, 32'hc2ab6b81, 32'h413a6e88, 32'h42abdd76, 32'hc23bfb37};
test_bias[3025:3025] = '{32'h42a6663f};
test_output[3025:3025] = '{32'h4640a264};
test_input[24208:24215] = '{32'hc20fab5b, 32'hc1c50281, 32'h41951855, 32'hc128f480, 32'hc2ac3cc4, 32'hc19805b7, 32'h42b8bdc5, 32'h4296e24a};
test_weights[24208:24215] = '{32'hc21aaf41, 32'h41a0f2f3, 32'hc21a3130, 32'hc2a2b9d6, 32'h3fe7b136, 32'hc2a05550, 32'hc219bfea, 32'h4267af3c};
test_bias[3026:3026] = '{32'hc0d2628d};
test_output[3026:3026] = '{32'h4548e661};
test_input[24216:24223] = '{32'hc16b699b, 32'hc2802047, 32'hc255799e, 32'h4231e492, 32'h42b70f70, 32'h428c3e26, 32'hc2b4598b, 32'h42a474bd};
test_weights[24216:24223] = '{32'h422f0329, 32'hc08ca008, 32'h421f2648, 32'h42a659c2, 32'h42aa4519, 32'hc1fb49d9, 32'hc145f51b, 32'hc1f821d7};
test_bias[3027:3027] = '{32'h42094f83};
test_output[3027:3027] = '{32'h45a8d6cb};
test_input[24224:24231] = '{32'hc1f090d7, 32'h429e3d20, 32'h42afa0b2, 32'hc2a1e82e, 32'h428c48c2, 32'hc2a61e63, 32'h4215ed1b, 32'hc16a42b1};
test_weights[24224:24231] = '{32'hc1539153, 32'hc088baa1, 32'h4279a833, 32'h429af079, 32'h42b1d062, 32'h41962abb, 32'h424aa432, 32'hc0f8ca2a};
test_bias[3028:3028] = '{32'h42b2280d};
test_output[3028:3028] = '{32'h45bcfdd5};
test_input[24232:24239] = '{32'hc1cd7b31, 32'h419726ed, 32'hc29bd44f, 32'h41e4429e, 32'h424e30fc, 32'h4262022b, 32'h420597fc, 32'h3f6cb9c3};
test_weights[24232:24239] = '{32'h42367d2f, 32'h42aa6d06, 32'h4185f001, 32'hc29f344c, 32'h42c7b56f, 32'hc05485a9, 32'h3f1c9adc, 32'hc2aea62c};
test_bias[3029:3029] = '{32'hc205965f};
test_output[3029:3029] = '{32'h44d80d8c};
test_input[24240:24247] = '{32'h42c4a5e8, 32'h40637e76, 32'hc24a00df, 32'h42214cbd, 32'h41f62427, 32'hc2ad1cea, 32'h42b55736, 32'h415d93b9};
test_weights[24240:24247] = '{32'hc1efd7ac, 32'hc284a0f8, 32'h422ba086, 32'hc2909f1d, 32'hc22fd7e9, 32'h42ad03f4, 32'h41809a43, 32'h426fbcf7};
test_bias[3030:3030] = '{32'h42312564};
test_output[3030:3030] = '{32'hc666db27};
test_input[24248:24255] = '{32'hc1fcbf13, 32'hc19f1d61, 32'hc21fe66a, 32'hc18102e1, 32'hc2b97258, 32'hc215d639, 32'h424486c9, 32'h404b035b};
test_weights[24248:24255] = '{32'h418fa3c8, 32'hc2c0bafb, 32'hc169a9e9, 32'hc2be550d, 32'h4260891f, 32'hc10f4b2d, 32'hc276552e, 32'h42a783f2};
test_bias[3031:3031] = '{32'hc2962cc7};
test_output[3031:3031] = '{32'hc584654a};
test_input[24256:24263] = '{32'h41e035c9, 32'hc234e050, 32'h4238f530, 32'h42bf5174, 32'hc296fc85, 32'hc1ca1d9a, 32'hc18da076, 32'h426ebffd};
test_weights[24256:24263] = '{32'hc22d7008, 32'hc1e16b04, 32'hc1306a4b, 32'h42372733, 32'hc2950c99, 32'hc23bae56, 32'h42b468ac, 32'h42824591};
test_bias[3032:3032] = '{32'h4208e33f};
test_output[3032:3032] = '{32'h464c272a};
test_input[24264:24271] = '{32'h4200ab0c, 32'hc2308bf2, 32'hc0d7c20b, 32'h4281de75, 32'h4290be43, 32'h42b61c39, 32'hc20f3ddb, 32'hc290e3c1};
test_weights[24264:24271] = '{32'h42b8ad2f, 32'h42b6ac76, 32'hc249c3c3, 32'h41d598c6, 32'hc0d0a6a2, 32'h41d41abc, 32'h4125df84, 32'hc2550c43};
test_bias[3033:3033] = '{32'h4262aa18};
test_output[3033:3033] = '{32'h45cb17fe};
test_input[24272:24279] = '{32'h42ad7d52, 32'hc139c76c, 32'h41b928a6, 32'h411cb079, 32'hc025ea9a, 32'h42822845, 32'hc256f3a3, 32'hc2b4428c};
test_weights[24272:24279] = '{32'h42b9b75e, 32'h42403291, 32'h42b5f659, 32'h402e188f, 32'h422adc8d, 32'hc23af77d, 32'hc2bd271a, 32'hc2c560dc};
test_bias[3034:3034] = '{32'h419e9ccf};
test_output[3034:3034] = '{32'h469ff3a7};
test_input[24280:24287] = '{32'hc14529f9, 32'h4246730c, 32'h42aedff6, 32'h41a14402, 32'h41c27a57, 32'h421db9a2, 32'h426889f7, 32'hc1fcc27c};
test_weights[24280:24287] = '{32'h3fe12936, 32'h42997d35, 32'hc244fff7, 32'hc1ccc0a9, 32'hc195e18b, 32'hc2c5b568, 32'hc0b5639f, 32'hc2ba4fc7};
test_bias[3035:3035] = '{32'hc2bcee53};
test_output[3035:3035] = '{32'hc53368f8};
test_input[24288:24295] = '{32'h42bb9c16, 32'hc2c29bef, 32'hc286871b, 32'h41d2fa5f, 32'hc2a67b62, 32'hc281c230, 32'hc2a9124d, 32'h42c24a23};
test_weights[24288:24295] = '{32'h41bdc72f, 32'hc292a735, 32'h42c423e1, 32'h42947ab9, 32'hc1e139fa, 32'hc293dce7, 32'h42af28cd, 32'h424a81dc};
test_bias[3036:3036] = '{32'h4132f097};
test_output[3036:3036] = '{32'h4612ad96};
test_input[24296:24303] = '{32'h4221147b, 32'hc0613e9d, 32'h4209222c, 32'h42b1f0d5, 32'hc29aa7a9, 32'h429559c5, 32'hc2b33984, 32'hc2220908};
test_weights[24296:24303] = '{32'h4294aee9, 32'hc29de712, 32'hc2b734fd, 32'hc1a34c44, 32'h428ef9fd, 32'hc2b627c3, 32'hc21cdd6d, 32'h42b8abe2};
test_bias[3037:3037] = '{32'hc2b5abad};
test_output[3037:3037] = '{32'hc65fecd3};
test_input[24304:24311] = '{32'hc27b5cbe, 32'hbe98da52, 32'h4267c1d9, 32'hc1a2e2cc, 32'hc2bd36e2, 32'hc2625cfb, 32'hc221fdd1, 32'h42985b4f};
test_weights[24304:24311] = '{32'h411a9e8c, 32'hc17e17f9, 32'hc2a6bb55, 32'h42415377, 32'hc2175561, 32'hc29ec474, 32'h41d3c966, 32'h41b1d803};
test_bias[3038:3038] = '{32'hc224350a};
test_output[3038:3038] = '{32'h450bb40d};
test_input[24312:24319] = '{32'hc29c4829, 32'h4287c76d, 32'h41a943fb, 32'h42a51fce, 32'hc1e3163a, 32'hc2c03f5f, 32'h41c8d98d, 32'hc1f8a085};
test_weights[24312:24319] = '{32'h4200f756, 32'hc2229c98, 32'hc28e5746, 32'hc29a5acf, 32'h42bf60e6, 32'hc13e3b3c, 32'hc1ff63cd, 32'h427e638d};
test_bias[3039:3039] = '{32'hc19b1047};
test_output[3039:3039] = '{32'hc688ef91};
test_input[24320:24327] = '{32'hc288d17d, 32'h419cb9d5, 32'h4292eeac, 32'hc1475776, 32'hc275fe29, 32'hc23360e8, 32'hc2a7186d, 32'h40b777ea};
test_weights[24320:24327] = '{32'hc1c69d88, 32'hc2c6f0c9, 32'hc286c539, 32'hc2a0af61, 32'hc28bff88, 32'h428adb93, 32'hc1a1c309, 32'hc10f7591};
test_bias[3040:3040] = '{32'h4279e5b9};
test_output[3040:3040] = '{32'hc4a3845c};
test_input[24328:24335] = '{32'h4067bd2e, 32'hc1e8f533, 32'h42c11427, 32'hc2588f5f, 32'h42b35682, 32'hc23d7d3a, 32'h426dd6ae, 32'h42a88107};
test_weights[24328:24335] = '{32'h40a57711, 32'h41c69ff7, 32'h419da93e, 32'h41edc115, 32'hc2383ffb, 32'hc2651ba5, 32'hc1ec4b14, 32'hc22abc90};
test_bias[3041:3041] = '{32'h404cd6b7};
test_output[3041:3041] = '{32'hc5e04800};
test_input[24336:24343] = '{32'hc205a187, 32'h429cb85d, 32'h40750cd3, 32'h41662877, 32'hc20bd73e, 32'h42431e2c, 32'h404a0572, 32'h42197f08};
test_weights[24336:24343] = '{32'hc21f66df, 32'hc19e1e11, 32'hc21c8148, 32'h4103ec4c, 32'hc25f6eb7, 32'h4237fc34, 32'hc2908cdc, 32'h42959c3c};
test_bias[3042:3042] = '{32'hc2964a96};
test_output[3042:3042] = '{32'h45cb98f8};
test_input[24344:24351] = '{32'hc299bf3d, 32'h42ad0ae5, 32'h425e8761, 32'h42aea21a, 32'hc2a09355, 32'hc1a23bd5, 32'hc19cc1a1, 32'h41f15820};
test_weights[24344:24351] = '{32'hc29b9446, 32'h412977c0, 32'hc2249170, 32'hc1a31b9f, 32'h42514c0a, 32'h4228f71c, 32'hc2116cd8, 32'h4253310b};
test_bias[3043:3043] = '{32'hc2b1961a};
test_output[3043:3043] = '{32'hc15ec717};
test_input[24352:24359] = '{32'hc2930a9d, 32'hc2a072ea, 32'hc2545337, 32'hc297b8e2, 32'h41e05f40, 32'hc271b11a, 32'h42286df6, 32'hc2a45786};
test_weights[24352:24359] = '{32'h423bfac1, 32'hc24eebbd, 32'hc28cb084, 32'h4267217a, 32'hc1fb9f05, 32'hbf5c1e88, 32'hc2b9b674, 32'hc2bba6a9};
test_bias[3044:3044] = '{32'hc2ac1e06};
test_output[3044:3044] = '{32'h4537102e};
test_input[24360:24367] = '{32'hc24c6960, 32'hc18c2596, 32'h4073560a, 32'hc2bc80c6, 32'h402694b7, 32'h42af1253, 32'h4222c153, 32'hc2a548d0};
test_weights[24360:24367] = '{32'hc28d3e62, 32'h41ce7cad, 32'hc2b6e010, 32'h4252e5ef, 32'hc229d96f, 32'hc2af9d66, 32'hbf72f244, 32'h40de213e};
test_bias[3045:3045] = '{32'hc1c4dace};
test_output[3045:3045] = '{32'hc62587a2};
test_input[24368:24375] = '{32'h4257f353, 32'hc22fb670, 32'hc2be46d1, 32'h426218ea, 32'hc28093b2, 32'hc22c2030, 32'hc0a36edf, 32'h418c35a1};
test_weights[24368:24375] = '{32'hc2862c09, 32'hc2b19af9, 32'hc2884c26, 32'h42c1fff3, 32'hc2c09978, 32'hc272f09d, 32'hc2715e56, 32'h41ba26be};
test_bias[3046:3046] = '{32'h425ea2f1};
test_output[3046:3046] = '{32'h46aa7b56};
test_input[24376:24383] = '{32'h400f8d69, 32'hc1827596, 32'hc084e5c0, 32'hc260c8eb, 32'hc279a0be, 32'h41ed4a82, 32'hc1f8ae60, 32'h422cda4a};
test_weights[24376:24383] = '{32'hc26f03e6, 32'hc21c013e, 32'h420a332b, 32'h416a8c88, 32'h42890163, 32'hc1e8404d, 32'hc2c67781, 32'h426f5df0};
test_bias[3047:3047] = '{32'h42122fbb};
test_output[3047:3047] = '{32'h42d370a2};
test_input[24384:24391] = '{32'hc2963c01, 32'hc2c32527, 32'h42b0057e, 32'h41c26be6, 32'hc2850616, 32'hc1d90a59, 32'hc23510c5, 32'hc1a07425};
test_weights[24384:24391] = '{32'hc268136c, 32'h428ee3c5, 32'hc20e892f, 32'h41124134, 32'h428a7ea0, 32'hc2750878, 32'hc224fee5, 32'hc1beb528};
test_bias[3048:3048] = '{32'h42c66cc6};
test_output[3048:3048] = '{32'hc5bc5153};
test_input[24392:24399] = '{32'h4246cd05, 32'hc25e2367, 32'h4291f1e2, 32'h42746752, 32'h426e08ee, 32'h42bfc050, 32'h42781fa9, 32'hc22f7f9a};
test_weights[24392:24399] = '{32'hc28d4976, 32'hc2b611f8, 32'hc2c6eaf2, 32'hc1df7d4a, 32'h41e2582a, 32'hc0a1dfd1, 32'hc1aa077a, 32'h42c1e5dd};
test_bias[3049:3049] = '{32'hc2424032};
test_output[3049:3049] = '{32'hc63907be};
test_input[24400:24407] = '{32'hc2ac9c10, 32'hc25aeb44, 32'h41cd736f, 32'hc2c65421, 32'hc25447c8, 32'h421ce9ef, 32'hc2b59683, 32'h42944ca7};
test_weights[24400:24407] = '{32'hc1cb2fd4, 32'h418d192f, 32'hc2b910db, 32'hc29bc2cc, 32'h424b0a54, 32'hc2902abb, 32'h42c7aef7, 32'h42746f34};
test_bias[3050:3050] = '{32'h4276dd75};
test_output[3050:3050] = '{32'hc555c626};
test_input[24408:24415] = '{32'hc25ff976, 32'h42a7ac66, 32'hc2851e72, 32'hc2c4f177, 32'h4257b5c2, 32'hc25e5638, 32'hc290535f, 32'h41a8c2f8};
test_weights[24408:24415] = '{32'h42b4a2ae, 32'h42a999a3, 32'h422c994f, 32'hc216b6fc, 32'h402d25df, 32'hc2c73a3f, 32'h4144b9c1, 32'h424bdbb9};
test_bias[3051:3051] = '{32'hc12b7ff3};
test_output[3051:3051] = '{32'h4608b97e};
test_input[24416:24423] = '{32'hc24f0671, 32'h4231b877, 32'h4298d3d2, 32'h40372409, 32'hc2c72f76, 32'hc14ab99f, 32'hc1eb55af, 32'hc20a51a6};
test_weights[24416:24423] = '{32'h42400d05, 32'h4271abd3, 32'hc2882276, 32'hc2177da5, 32'h42a56674, 32'h42a88338, 32'hc201b985, 32'h42553151};
test_bias[3052:3052] = '{32'hc286ebca};
test_output[3052:3052] = '{32'hc6702a61};
test_input[24424:24431] = '{32'hc2b90984, 32'h4284138f, 32'h42c4e899, 32'h41e4a3b0, 32'h423c95d5, 32'hc2331cb0, 32'h42c1c10c, 32'h423fff22};
test_weights[24424:24431] = '{32'hc2924b17, 32'h41b8bba3, 32'h42b366a9, 32'h4297c747, 32'h4268a452, 32'h40a34482, 32'hc15d3594, 32'hc27f16f3};
test_bias[3053:3053] = '{32'h428998db};
test_output[3053:3053] = '{32'h4688854b};
test_input[24432:24439] = '{32'h4166bfea, 32'hc2943667, 32'h425b6599, 32'h4071a2b5, 32'hc2c4e418, 32'h41b89cc1, 32'h410959c1, 32'h42881010};
test_weights[24432:24439] = '{32'h429266ad, 32'h4234d1ab, 32'h41d4fe27, 32'hc29d8f6d, 32'hc29c9e75, 32'hc2800f08, 32'h4187eb4a, 32'h422068d8};
test_bias[3054:3054] = '{32'hc288e2ec};
test_output[3054:3054] = '{32'h45f70ef7};
test_input[24440:24447] = '{32'h41e27320, 32'h41ea9ef7, 32'h419041d3, 32'hc11a391a, 32'h4283bbd5, 32'hc285019c, 32'hc2c53d91, 32'h42027403};
test_weights[24440:24447] = '{32'h421a8ede, 32'hc2b8156c, 32'h426766d1, 32'hc2c1e9a2, 32'hc1bcf815, 32'hc14da475, 32'hc2afb1db, 32'h422db6a7};
test_bias[3055:3055] = '{32'hc29bd3e2};
test_output[3055:3055] = '{32'h461723c6};
test_input[24448:24455] = '{32'hc18824cb, 32'hbf72cae3, 32'hbfca7b8f, 32'hc2010c2c, 32'hc2bdc33e, 32'h40f7d65d, 32'h41c04b7a, 32'hc1ebe1d1};
test_weights[24448:24455] = '{32'hc1e2c2f1, 32'h429ba044, 32'h42487644, 32'hc2c4e2e1, 32'hc1bd292a, 32'hc22b2429, 32'h420d7f20, 32'h4282d8fd};
test_bias[3056:3056] = '{32'h428fc77e};
test_output[3056:3056] = '{32'h4589d40e};
test_input[24456:24463] = '{32'h410800b6, 32'hc24be31b, 32'hc248ff46, 32'h429a1b89, 32'hc2552ca5, 32'h42112a7a, 32'hc229e80f, 32'h42b2e278};
test_weights[24456:24463] = '{32'h42a701fc, 32'h4299aad3, 32'h41c062b3, 32'hc1f4a1bd, 32'h42254e2d, 32'h42bbd77f, 32'hc2422b39, 32'h412fdfc5};
test_bias[3057:3057] = '{32'h41247f95};
test_output[3057:3057] = '{32'hc51cdbae};
test_input[24464:24471] = '{32'h42283970, 32'hc2a68f98, 32'h412ffae8, 32'h42990add, 32'h4170e2b4, 32'h4155a486, 32'h4285a234, 32'h41cdce73};
test_weights[24464:24471] = '{32'h41185b4e, 32'h41027436, 32'hc1635ece, 32'h429a94d2, 32'h4283925f, 32'hc21ed597, 32'hc290dc78, 32'hc2b21824};
test_bias[3058:3058] = '{32'h42907a3f};
test_output[3058:3058] = '{32'hc48bcd0f};
test_input[24472:24479] = '{32'h428215a6, 32'h41428457, 32'h42ad63db, 32'hc290aea4, 32'hc1b37539, 32'h406f107d, 32'hc189bbf9, 32'h429ee6b2};
test_weights[24472:24479] = '{32'h410ac317, 32'h4296dfed, 32'hc1744254, 32'h41614e49, 32'h42387138, 32'h428bc5fd, 32'hc2a0cf72, 32'hc26a7bc8};
test_bias[3059:3059] = '{32'h4276fb89};
test_output[3059:3059] = '{32'hc5976d81};
test_input[24480:24487] = '{32'h424ad533, 32'hc28e362a, 32'hc28e7d13, 32'h413cd73f, 32'h42830b33, 32'h42400ff0, 32'hc1f0880b, 32'h40db338a};
test_weights[24480:24487] = '{32'hc2672c7c, 32'h41a222a3, 32'h4265ed78, 32'h4285a402, 32'h41d2260d, 32'hc252f63e, 32'h4259235a, 32'h42b71851};
test_bias[3060:3060] = '{32'hc1a0c1bb};
test_output[3060:3060] = '{32'hc614aa88};
test_input[24488:24495] = '{32'hc242d822, 32'hc22250c5, 32'hc25ef1b4, 32'h4298340a, 32'h422e6f50, 32'h428b8b43, 32'h421023fe, 32'h4256f993};
test_weights[24488:24495] = '{32'hc22ac313, 32'h4198598b, 32'hc2c696e3, 32'h42993e53, 32'hc162301e, 32'hc2a3c60b, 32'h42421207, 32'h42a16216};
test_bias[3061:3061] = '{32'h4282e3e5};
test_output[3061:3061] = '{32'h46433279};
test_input[24496:24503] = '{32'hc244535b, 32'h42198d62, 32'hc1e9ff32, 32'hc24a2af4, 32'h426ffc88, 32'h410c4f08, 32'hc2ae3647, 32'hc10e4731};
test_weights[24496:24503] = '{32'h4222ebd0, 32'hbffdab04, 32'h412cd2cb, 32'hc2bb9dab, 32'hc225ba1f, 32'hc2bcbdec, 32'hc1d93fe4, 32'hc22ad6a2};
test_bias[3062:3062] = '{32'h42ae5ca3};
test_output[3062:3062] = '{32'h44e9a74d};
test_input[24504:24511] = '{32'h4272bd54, 32'h416db6f5, 32'hc0d2e405, 32'h42a2a16a, 32'h4294bca1, 32'h418e03b3, 32'h42accedd, 32'h42b253a6};
test_weights[24504:24511] = '{32'h4241c2d7, 32'h42a83432, 32'h41a69d04, 32'hc1272e03, 32'hc1d30c0a, 32'h424d3573, 32'h42bfde96, 32'h42bfea33};
test_bias[3063:3063] = '{32'hc19ada07};
test_output[3063:3063] = '{32'h46944164};
test_input[24512:24519] = '{32'h4024c2ff, 32'hc248f557, 32'hc241f6bd, 32'h426c24a1, 32'hc29f4eba, 32'hc2b62509, 32'h415591c7, 32'h4181a39b};
test_weights[24512:24519] = '{32'h42af9b3d, 32'hc297f159, 32'hc29df4f3, 32'hc2bb62c4, 32'h403af18f, 32'hbea54764, 32'h415ec891, 32'h42909ad9};
test_bias[3064:3064] = '{32'h40a4edb1};
test_output[3064:3064] = '{32'h455acb6b};
test_input[24520:24527] = '{32'hc22939c4, 32'h4245e83b, 32'hc1a7c6fe, 32'hc1749ec7, 32'h42a8f709, 32'h42874e6f, 32'hc28d309a, 32'h42a5cf9b};
test_weights[24520:24527] = '{32'h422b8cda, 32'hc2848881, 32'h4236759c, 32'hc16d42cf, 32'hc1974227, 32'h4098ae49, 32'hc289f5d3, 32'h428e1df3};
test_bias[3065:3065] = '{32'hc2108556};
test_output[3065:3065] = '{32'h4562b1b3};
test_input[24528:24535] = '{32'h40b92e62, 32'hc1777f4b, 32'hc2922f89, 32'hc298cc52, 32'hc2182f49, 32'hc2a82e53, 32'hc254c0c2, 32'hc2851cb3};
test_weights[24528:24535] = '{32'h42c42e0c, 32'h42a2c155, 32'h42adce45, 32'hc2c738bd, 32'h41a78b4f, 32'h40f51bb1, 32'h427f143b, 32'h421c4b41};
test_bias[3066:3066] = '{32'hc0ba37bd};
test_output[3066:3066] = '{32'hc5d6c084};
test_input[24536:24543] = '{32'hc2823428, 32'hc2753f7e, 32'hc149bc33, 32'hc2480b20, 32'hc280e443, 32'h41eaa48d, 32'hc2b65ca4, 32'hc2415e9e};
test_weights[24536:24543] = '{32'h4200b498, 32'hc28de3ca, 32'h42294ec2, 32'h427f6ecb, 32'h4233d512, 32'h42a35c88, 32'h424af5ac, 32'hc25804ba};
test_bias[3067:3067] = '{32'h42807ad5};
test_output[3067:3067] = '{32'hc575571b};
test_input[24544:24551] = '{32'hc28d2f45, 32'hc24a8f3d, 32'hc2a9f867, 32'h4272fd4c, 32'hc13066f1, 32'hc204816c, 32'h420c4e06, 32'h427e388a};
test_weights[24544:24551] = '{32'h428de962, 32'hc27db637, 32'hc1890c90, 32'h427713b7, 32'hc2b4567e, 32'h4213b942, 32'hc236013b, 32'h426c79be};
test_bias[3068:3068] = '{32'h411dd8ae};
test_output[3068:3068] = '{32'h45a74952};
test_input[24552:24559] = '{32'h42820b18, 32'h42babb55, 32'h42a38dc0, 32'h42b561ea, 32'hc28249a1, 32'hc1676418, 32'h4222d9f7, 32'hc2a1e23e};
test_weights[24552:24559] = '{32'h3ff6862b, 32'hc289c261, 32'hc298d8ee, 32'h428373a8, 32'hc0aea7e0, 32'hc26cf91c, 32'h422adc1f, 32'h42354a9c};
test_bias[3069:3069] = '{32'hc260d4bf};
test_output[3069:3069] = '{32'hc5e64072};
test_input[24560:24567] = '{32'h429ba59b, 32'hc26046db, 32'hc28040a5, 32'hc2489067, 32'h42b64db3, 32'h4293c2d9, 32'hc1bf64f6, 32'hbeaddabb};
test_weights[24560:24567] = '{32'hc2a9cb6e, 32'hc1d8efca, 32'h42977a12, 32'hc21bcb1b, 32'h3f51ddf4, 32'hc29c2ea6, 32'h426d9a61, 32'hc18f1b38};
test_bias[3070:3070] = '{32'hc207a018};
test_output[3070:3070] = '{32'hc66c7880};
test_input[24568:24575] = '{32'h42962525, 32'h42151cb0, 32'h41f77979, 32'hc2bf2644, 32'hc29dc77a, 32'hc23a7954, 32'hc1969511, 32'h422289f3};
test_weights[24568:24575] = '{32'hc2300aca, 32'hc24fc548, 32'h429ecdc8, 32'hc1cbfd84, 32'h42c19758, 32'h42c0cb25, 32'h429f3532, 32'hc09b911e};
test_bias[3071:3071] = '{32'h42b67e2e};
test_output[3071:3071] = '{32'hc65c06e1};
test_input[24576:24583] = '{32'hc20fb748, 32'hc1960fd2, 32'h4284f648, 32'h420b2993, 32'hc25646f5, 32'h4229425b, 32'h42953d64, 32'h41f1ef67};
test_weights[24576:24583] = '{32'h425141c1, 32'hc283b33f, 32'h42c4037f, 32'hc285be28, 32'h41508676, 32'h42a72ec9, 32'hc19fb877, 32'h42a600c8};
test_bias[3072:3072] = '{32'h4184c450};
test_output[3072:3072] = '{32'h45e7e4f5};
test_input[24584:24591] = '{32'h41c82ddd, 32'h42befd67, 32'h428a01e8, 32'hc2629386, 32'h420bc0e9, 32'hc2c387ca, 32'hc1aa07df, 32'h42c1eeda};
test_weights[24584:24591] = '{32'h418ecae5, 32'h42660cf2, 32'h414a812c, 32'h428fd41e, 32'h429341b9, 32'hc1aab88d, 32'h42932644, 32'hc2c43aca};
test_bias[3073:3073] = '{32'h4182c809};
test_output[3073:3073] = '{32'hc564fd9b};
test_input[24592:24599] = '{32'hc0741a39, 32'h423e3ec7, 32'hc1a2eec9, 32'h421a44e1, 32'hc1444a23, 32'hc28f3a2a, 32'hc2aba687, 32'h3ef0acb2};
test_weights[24592:24599] = '{32'hc2b55f37, 32'h4270a280, 32'hc204effd, 32'h4282f16b, 32'hc1fba6f2, 32'h429e98de, 32'h426a1a8d, 32'hc2c6a7d3};
test_bias[3074:3074] = '{32'hc2b4fa08};
test_output[3074:3074] = '{32'hc57cc163};
test_input[24600:24607] = '{32'hc2a76270, 32'hc2923c18, 32'hc0e0e3c6, 32'h42c7d742, 32'hc292df9b, 32'hc2c015f3, 32'h42a56637, 32'hc185271d};
test_weights[24600:24607] = '{32'h42abdcde, 32'h41912f7f, 32'hc2c5f27a, 32'h41cf0db9, 32'h42bf226e, 32'h42382cb1, 32'h42b62a45, 32'hc2c46456};
test_bias[3075:3075] = '{32'hc29495bc};
test_output[3075:3075] = '{32'hc5ed0649};
test_input[24608:24615] = '{32'hc16a5790, 32'hc12b667e, 32'h42a7e3d6, 32'h42a5eee4, 32'hc171e0ba, 32'h42210aa7, 32'hc2113f6f, 32'h427d678e};
test_weights[24608:24615] = '{32'h42a5a8b0, 32'h42a71b4f, 32'h4242384a, 32'h42c50462, 32'h427f7c05, 32'hc0bc2f7b, 32'h428d952c, 32'h42408d1f};
test_bias[3076:3076] = '{32'hc274f1e2};
test_output[3076:3076] = '{32'h46123063};
test_input[24616:24623] = '{32'hc25ff051, 32'h422c48cd, 32'hc2962fbe, 32'hc1b591d7, 32'hc1e26ae8, 32'h40ada1e1, 32'h4259932f, 32'h424ae2a1};
test_weights[24616:24623] = '{32'h4064eadf, 32'h424030c5, 32'hc2ad5204, 32'h42823ede, 32'h4289b509, 32'hc2321c62, 32'h42b39e29, 32'h42472350};
test_bias[3077:3077] = '{32'h4161ec7c};
test_output[3077:3077] = '{32'h463d9301};
test_input[24624:24631] = '{32'hc1868897, 32'h42aa44b9, 32'h402b1c96, 32'hc2b58f45, 32'hc1c92e7d, 32'hc2745d26, 32'h42c7583b, 32'hc17d0b4d};
test_weights[24624:24631] = '{32'hc22c6869, 32'hc276a34e, 32'hc2153863, 32'h4214a1bf, 32'h41709d05, 32'h40e0bb9c, 32'h42b4b76c, 32'hc292220a};
test_bias[3078:3078] = '{32'hc253cf95};
test_output[3078:3078] = '{32'h44a305d8};
test_input[24632:24639] = '{32'hc2aa51b5, 32'hc24a9a6b, 32'h419eb964, 32'h4297044e, 32'hc238b8e7, 32'hc22e61af, 32'hc28043a0, 32'h4295809d};
test_weights[24632:24639] = '{32'h41c62607, 32'h422c4637, 32'h426a7a70, 32'h42a1215c, 32'hc2a00d05, 32'hc20c6074, 32'hc27e6259, 32'h425715d1};
test_bias[3079:3079] = '{32'hc094ebb5};
test_output[3079:3079] = '{32'h467e4a50};
test_input[24640:24647] = '{32'hc2509a45, 32'hc093f59b, 32'hc0731428, 32'hc287c9ec, 32'hc229fcfb, 32'h42ac00ef, 32'hc220e4cf, 32'hc245cd8f};
test_weights[24640:24647] = '{32'hc14ebbd7, 32'h42c5d1b2, 32'h42177fd4, 32'h429dc906, 32'h41b2f14e, 32'h427b4489, 32'hc2c38e6f, 32'hc259c1d9};
test_bias[3080:3080] = '{32'h42b58b17};
test_output[3080:3080] = '{32'h45b7df2b};
test_input[24648:24655] = '{32'h4222f053, 32'h423df6d7, 32'hc2a88671, 32'h426e3b20, 32'hc1f2baf3, 32'h41db3612, 32'hc290a9a5, 32'h4276797f};
test_weights[24648:24655] = '{32'h4244f5e9, 32'h427e217c, 32'h42083b8d, 32'h4291ce22, 32'hc284509b, 32'hc1e4b100, 32'h42926ded, 32'h4214801e};
test_bias[3081:3081] = '{32'h41b71da3};
test_output[3081:3081] = '{32'h4593eef2};
test_input[24656:24663] = '{32'h4135816e, 32'h42b1f16b, 32'hc28a78cf, 32'hc288719b, 32'hc2532e39, 32'hc1c3af6a, 32'hc2a575bf, 32'hc2a134f3};
test_weights[24656:24663] = '{32'h41b1ed73, 32'h4242322f, 32'hc039565f, 32'hc231951b, 32'hc1f143a9, 32'hc28ecdf1, 32'hc27fb174, 32'hc1e8323e};
test_bias[3082:3082] = '{32'hc2a957a6};
test_output[3082:3082] = '{32'h4691f5e9};
test_input[24664:24671] = '{32'h429fdfd0, 32'h412639e8, 32'h42aed89f, 32'h40d9c919, 32'hc1c591e6, 32'hc11a4095, 32'h42b6990e, 32'h425ab2e4};
test_weights[24664:24671] = '{32'hc28664a9, 32'hc29ed829, 32'h41f0a19c, 32'hc2ad25ed, 32'hc258b4ae, 32'hc12a5ffb, 32'hc2af9eb7, 32'h42101136};
test_bias[3083:3083] = '{32'hc28379b1};
test_output[3083:3083] = '{32'hc609f47c};
test_input[24672:24679] = '{32'h4212f3d7, 32'h42bc7cb6, 32'h422a7efd, 32'hc17ae95b, 32'hc1d35675, 32'hc2b6c12c, 32'h422fd3a4, 32'hc2a038ca};
test_weights[24672:24679] = '{32'hc26bf19a, 32'hc1a93879, 32'h42bef130, 32'h41ca122b, 32'hc22d17d8, 32'h42a4137d, 32'hc2bc07c7, 32'h42299de2};
test_bias[3084:3084] = '{32'h42859d04};
test_output[3084:3084] = '{32'hc65f7d70};
test_input[24680:24687] = '{32'h42535548, 32'hc2ad3a3a, 32'h40fcd024, 32'hc2946a29, 32'h416837c3, 32'hc269db0e, 32'hc2c27356, 32'h42039434};
test_weights[24680:24687] = '{32'hc238e59d, 32'hc2c732ac, 32'hc198fd34, 32'h40ae9877, 32'h42210e70, 32'h42836bcb, 32'h422c9800, 32'hc18b6729};
test_bias[3085:3085] = '{32'h422fd0aa};
test_output[3085:3085] = '{32'hc5131318};
test_input[24688:24695] = '{32'h42961a89, 32'hc222a661, 32'h4244fb59, 32'hc28da6ef, 32'hc2b54ba5, 32'h40a1568d, 32'h418a3761, 32'h42123474};
test_weights[24688:24695] = '{32'hc2b028e8, 32'hc226ce07, 32'h4222448e, 32'h4092386e, 32'hc20eb9fa, 32'hc1b79fc4, 32'h42b27f9d, 32'h421aaae0};
test_bias[3086:3086] = '{32'hc247deca};
test_output[3086:3086] = '{32'h452df461};
test_input[24696:24703] = '{32'h425b6c61, 32'hc2c75ec1, 32'hc25fe065, 32'hc261cd5f, 32'h424e050d, 32'hbfe3eee3, 32'h41d54cc9, 32'h419fd0f7};
test_weights[24696:24703] = '{32'hc2ac22ba, 32'hc21c18e6, 32'h42a02acb, 32'hc2181c05, 32'h42b3a26a, 32'h42b92b7f, 32'h41fd4dfe, 32'hc28a21aa};
test_bias[3087:3087] = '{32'hc0b8c14d};
test_output[3087:3087] = '{32'h443c49a7};
test_input[24704:24711] = '{32'hc245675c, 32'h41d2db11, 32'hc146d85f, 32'hc29c40d1, 32'hc1ccd505, 32'hc23e4db8, 32'h423de449, 32'h41a4b40f};
test_weights[24704:24711] = '{32'hc22fa7a1, 32'h42016980, 32'h42354663, 32'hc24212ef, 32'hc281e18b, 32'hc2a019c2, 32'h4238fc9a, 32'hc10d00f0};
test_bias[3088:3088] = '{32'h4286c891};
test_output[3088:3088] = '{32'h46579f9f};
test_input[24712:24719] = '{32'hc0ea2495, 32'hc2b553fd, 32'hc2557766, 32'h4220cea5, 32'h41efd426, 32'hc221d2de, 32'hc1afa41b, 32'h42a211fd};
test_weights[24712:24719] = '{32'h428b0757, 32'h4249a92c, 32'h42a435a7, 32'hc1c40621, 32'h42be6295, 32'h42095b78, 32'h42bc147b, 32'h42b761ea};
test_bias[3089:3089] = '{32'h4298dd74};
test_output[3089:3089] = '{32'hc55d3b47};
test_input[24720:24727] = '{32'hc2c292bf, 32'hc2a319a3, 32'h42ae7505, 32'hc2a6e958, 32'hc1689196, 32'h4246ac9f, 32'hc21b9da1, 32'hc2174030};
test_weights[24720:24727] = '{32'h428e5ac8, 32'h428677ee, 32'h429ad0c7, 32'hc231df86, 32'hc156554f, 32'h4016f510, 32'h429ae084, 32'hc2ab565d};
test_bias[3090:3090] = '{32'h429f8378};
test_output[3090:3090] = '{32'hc4a5bdb2};
test_input[24728:24735] = '{32'h42c6bab7, 32'hc2a9fce7, 32'hc2a2fd03, 32'hc11558e7, 32'hc20f02b0, 32'h4250f0bf, 32'hc2ac9d76, 32'hc21af302};
test_weights[24728:24735] = '{32'hc2180633, 32'hc2b5e496, 32'h4276ddcb, 32'hc29538d8, 32'hc2502cda, 32'h429fe448, 32'hc18a4391, 32'h4217d8da};
test_bias[3091:3091] = '{32'h42273da6};
test_output[3091:3091] = '{32'h45b2bf85};
test_input[24736:24743] = '{32'hc21039c8, 32'h421528dd, 32'hc2878826, 32'hc07b983f, 32'h429f5366, 32'h428b9b9b, 32'h4247814a, 32'h4274d648};
test_weights[24736:24743] = '{32'h4287ae1f, 32'hc2a7774a, 32'h3fe4c999, 32'hc0fae0d2, 32'hc1517a2a, 32'hc262195f, 32'hc2020747, 32'h421d8fec};
test_bias[3092:3092] = '{32'hc28811bb};
test_output[3092:3092] = '{32'hc61b16c8};
test_input[24744:24751] = '{32'h4135d9ec, 32'hc2a1cf3e, 32'h41ad71e6, 32'hc2a8d51b, 32'hc28cb05b, 32'h428e676d, 32'h42bb76c0, 32'hc2b9d2c6};
test_weights[24744:24751] = '{32'hc261c540, 32'hc212b42f, 32'h42229cfb, 32'h419e6986, 32'h41d0cdd0, 32'h42c34081, 32'hc103a7ac, 32'h41f074fe};
test_bias[3093:3093] = '{32'hc23e1717};
test_output[3093:3093] = '{32'h453df434};
test_input[24752:24759] = '{32'hc20b1b34, 32'hc29f008c, 32'h41dfdffa, 32'hc24277f9, 32'h42b6ae53, 32'h41575770, 32'h4282d90b, 32'hc1c7eca9};
test_weights[24752:24759] = '{32'h41867197, 32'hc228e73f, 32'h41577532, 32'h40b69f31, 32'hc2c129fe, 32'hc089b049, 32'h420405a9, 32'hc2a85eac};
test_bias[3094:3094] = '{32'hc29daa53};
test_output[3094:3094] = '{32'hc4e3eee0};
test_input[24760:24767] = '{32'hc1ab1371, 32'hc29947e7, 32'hc266fa32, 32'hc2af3e35, 32'hc2b6d3d1, 32'h427a148c, 32'h41ed20e5, 32'hc2990223};
test_weights[24760:24767] = '{32'hc1fb9cac, 32'h42b7c981, 32'h42aed2a1, 32'h42a8d7ec, 32'hc260e814, 32'hc29840e5, 32'h42c13ea4, 32'h4281e8ba};
test_bias[3095:3095] = '{32'h41d5d897};
test_output[3095:3095] = '{32'hc6a041fe};
test_input[24768:24775] = '{32'h429c5fb4, 32'h4298ccb3, 32'hc188ac9d, 32'hc239c0f0, 32'h428c7d8b, 32'hc2264dc5, 32'hc1b92463, 32'h424f6611};
test_weights[24768:24775] = '{32'h4291bb3c, 32'h42b18698, 32'hc23db528, 32'hbfc103df, 32'h41596336, 32'h42b60b6f, 32'hc1ffde89, 32'hc120a219};
test_bias[3096:3096] = '{32'h4179df95};
test_output[3096:3096] = '{32'h462830d9};
test_input[24776:24783] = '{32'hc0dfda21, 32'h41c1f83a, 32'h427adaf9, 32'h4104cb2a, 32'h420825eb, 32'hc1ce405a, 32'hc2439465, 32'h4248d5e7};
test_weights[24776:24783] = '{32'h42b6d49a, 32'h41303aee, 32'hc2bc1076, 32'h416ceaf0, 32'hc111d60f, 32'h423d8dc7, 32'h42802611, 32'h417cce33};
test_bias[3097:3097] = '{32'hc1c0ab7e};
test_output[3097:3097] = '{32'hc61ce93a};
test_input[24784:24791] = '{32'hc2126f29, 32'h4270797c, 32'h42380b68, 32'hc292040f, 32'hc19b22a6, 32'h42bbef8e, 32'hc23fd4df, 32'h409c4dd0};
test_weights[24784:24791] = '{32'hc25af561, 32'h415119af, 32'h42ac84dd, 32'hc25f176f, 32'h427f5f39, 32'hc2864244, 32'hc1c32373, 32'h428fda16};
test_bias[3098:3098] = '{32'h429f99d5};
test_output[3098:3098] = '{32'h4598aa08};
test_input[24792:24799] = '{32'h4273880e, 32'hc2c3c51e, 32'hc2536d9e, 32'hc29f68c2, 32'h40910f14, 32'h42aa5787, 32'h42a8743c, 32'hc1d4b77e};
test_weights[24792:24799] = '{32'hc2177bb6, 32'hc28da481, 32'h40e1a0e0, 32'hc202320a, 32'hc2324418, 32'hc2b7a2b5, 32'h41ce57b6, 32'h410bfa55};
test_bias[3099:3099] = '{32'h42c2d367};
test_output[3099:3099] = '{32'h4457d1a2};
test_input[24800:24807] = '{32'h42afdc38, 32'hc1df90c0, 32'hc2634269, 32'hc2b9f457, 32'h418c4a1c, 32'hc1684188, 32'hc2bbf171, 32'hc2692e76};
test_weights[24800:24807] = '{32'h41273675, 32'h42a232e9, 32'hc14f483b, 32'h420a87c2, 32'h41e19fc7, 32'h412d3ea0, 32'hc2341bfd, 32'hc24e1a49};
test_bias[3100:3100] = '{32'h420c1928};
test_output[3100:3100] = '{32'h456bffba};
test_input[24808:24815] = '{32'h4180676a, 32'h41038f1c, 32'h41d8f447, 32'hc288aa92, 32'h4216a7e5, 32'hc131cc68, 32'h418d1445, 32'h419e7edf};
test_weights[24808:24815] = '{32'h427112a9, 32'h42b76621, 32'hc245ee8f, 32'hc1c2e6ce, 32'hc2715c73, 32'hc26309e3, 32'hc2a69cb9, 32'hc26397e9};
test_bias[3101:3101] = '{32'h419d303e};
test_output[3101:3101] = '{32'hc507e772};
test_input[24816:24823] = '{32'hc2206c1e, 32'h424d9485, 32'hc2bc0566, 32'hc1824bdf, 32'hc279f482, 32'hc0bb548c, 32'h429fbb95, 32'hc2b44824};
test_weights[24816:24823] = '{32'hc2253941, 32'h429e261b, 32'h42931b79, 32'hc2645921, 32'h418eb237, 32'h42c2858b, 32'h42b7694c, 32'h41272df2};
test_bias[3102:3102] = '{32'hc184fa69};
test_output[3102:3102] = '{32'h458a0a99};
test_input[24824:24831] = '{32'h42245168, 32'hc27878bd, 32'h418c3db5, 32'hc2b98b21, 32'hc1a2f375, 32'h418951c1, 32'hc1c35e63, 32'hc00d62af};
test_weights[24824:24831] = '{32'hc1c9568a, 32'h41af5a2e, 32'h42b8c86d, 32'h42954d64, 32'h419203ee, 32'hc25a331d, 32'hc2950770, 32'h427fcd4c};
test_bias[3103:3103] = '{32'h409d60d1};
test_output[3103:3103] = '{32'hc5e4f06e};
test_input[24832:24839] = '{32'hc15d55b0, 32'h4202060a, 32'hc1067fe6, 32'h41e60f12, 32'h3fa49975, 32'hc0c44764, 32'hc22f62f2, 32'hc010a512};
test_weights[24832:24839] = '{32'h3fe2060c, 32'hc188a768, 32'h421afde1, 32'hc251188c, 32'h427e340d, 32'hbe32cdcc, 32'hc24e47ac, 32'h42bcb906};
test_bias[3104:3104] = '{32'h418b1ed8};
test_output[3104:3104] = '{32'hc3824a3e};
test_input[24840:24847] = '{32'hc18da96c, 32'h4277a9c4, 32'hc13aaff6, 32'hc0f00e6b, 32'h429f0658, 32'hc175a2ed, 32'h41fed667, 32'h4197d51a};
test_weights[24840:24847] = '{32'hc22f68d2, 32'h420c8aa0, 32'hc2a6dd3a, 32'h4276781b, 32'hc2b8e06e, 32'h42ac59c5, 32'hc24409bc, 32'hc1f58e87};
test_bias[3105:3105] = '{32'h41512454};
test_output[3105:3105] = '{32'hc5e5638a};
test_input[24848:24855] = '{32'h42921165, 32'hc260b31f, 32'hc214b729, 32'h42430831, 32'hc2b3860f, 32'h4130c201, 32'hbf9689da, 32'hc1bd3ea5};
test_weights[24848:24855] = '{32'h424084f0, 32'h42599ce4, 32'h427a9257, 32'hc2c40668, 32'h42a2cd0f, 32'h429718e6, 32'hc19b8b8a, 32'h41e19c75};
test_bias[3106:3106] = '{32'h41bdadff};
test_output[3106:3106] = '{32'hc656b5d7};
test_input[24856:24863] = '{32'h3f867f05, 32'h424faa20, 32'hc2b7d8cc, 32'h424b74b7, 32'hc29603d3, 32'hc2a60394, 32'hc22d6e19, 32'h429e7a36};
test_weights[24856:24863] = '{32'h4218a234, 32'hc20aace1, 32'h42ae8a8d, 32'hc25c6867, 32'hc22cd590, 32'h412ac0d9, 32'h4167f996, 32'h4231b37d};
test_bias[3107:3107] = '{32'h4292e778};
test_output[3107:3107] = '{32'hc5e30469};
test_input[24864:24871] = '{32'hc29d9a7f, 32'hc2ae7c8f, 32'hc07a3e85, 32'hc2447d24, 32'h42b54101, 32'h423c91d4, 32'hc128c26f, 32'hc2a8bbb6};
test_weights[24864:24871] = '{32'h42bc9649, 32'h42676216, 32'hc260e0ea, 32'h42998e88, 32'h42c47a8d, 32'hbf078a20, 32'hc2032cb3, 32'h42bdfa54};
test_bias[3108:3108] = '{32'hc299ef75};
test_output[3108:3108] = '{32'hc668be98};
test_input[24872:24879] = '{32'h40ba88c8, 32'hc2afd8ba, 32'hc0b50626, 32'hc17d22e9, 32'hc20682e6, 32'h428a0d91, 32'h416234db, 32'h429f81fa};
test_weights[24872:24879] = '{32'h42138fdb, 32'h422b6a34, 32'h3e1a80c7, 32'hc110ed7d, 32'h42a8d0d0, 32'hc299aa71, 32'hc1d48025, 32'h4074610a};
test_bias[3109:3109] = '{32'hc2bb26f5};
test_output[3109:3109] = '{32'hc6371389};
test_input[24880:24887] = '{32'h41ced14b, 32'h42212998, 32'hc2187294, 32'hc09095d1, 32'h407afaf1, 32'hc00849f9, 32'h41d8bd0a, 32'h42c126cd};
test_weights[24880:24887] = '{32'h42ae33fe, 32'h408de8d9, 32'h416945c9, 32'h42288fd8, 32'hc23f6c07, 32'hc10babb3, 32'h4203ae2c, 32'hc2931e2d};
test_bias[3110:3110] = '{32'h41d910da};
test_output[3110:3110] = '{32'hc591ed88};
test_input[24888:24895] = '{32'hc21357f8, 32'h4299a711, 32'h4121a728, 32'h422ae4a3, 32'hc1cf6f80, 32'hc06ea75f, 32'h4180422a, 32'h4246dd7f};
test_weights[24888:24895] = '{32'h3f9e36cb, 32'hc243f8a1, 32'h4252315f, 32'hc24f04fa, 32'h42492cc7, 32'hc22b7b8d, 32'h42becec6, 32'hc198c249};
test_bias[3111:3111] = '{32'h411e00f2};
test_output[3111:3111] = '{32'hc5bcde9a};
test_input[24896:24903] = '{32'h4289ea75, 32'hc16f4371, 32'h419ae0f2, 32'hc25fa0e5, 32'h42b5b3d7, 32'h41d45eee, 32'h41fdcdb2, 32'hc24265d5};
test_weights[24896:24903] = '{32'h419bd80f, 32'hc2846d4a, 32'h42788927, 32'hc2ba8fb5, 32'hc25c0fb3, 32'hc2566455, 32'h42b103b6, 32'h42c37ad9};
test_bias[3112:3112] = '{32'h42be2879};
test_output[3112:3112] = '{32'h43f1a73e};
test_input[24904:24911] = '{32'hc2c2ceba, 32'h41d9f2c8, 32'h418329b8, 32'hc1cca44d, 32'h429103d2, 32'hc14d8807, 32'hc118fa79, 32'hc1168033};
test_weights[24904:24911] = '{32'hc248e0f1, 32'hc2c3fdb3, 32'hc22dedf1, 32'h42a226de, 32'hc202b1cc, 32'h4204a504, 32'h413c94c0, 32'hc24cd8ba};
test_bias[3113:3113] = '{32'hc1055a57};
test_output[3113:3113] = '{32'hc53b7622};
test_input[24912:24919] = '{32'hc2c5384e, 32'hc241e41f, 32'hc2341053, 32'h41d62f53, 32'h4138c0b0, 32'hc2b18aee, 32'hc0bc43c2, 32'hc2bd5145};
test_weights[24912:24919] = '{32'h4219afce, 32'hc1dc8e32, 32'h423637c6, 32'hc1febdbf, 32'hc21d135b, 32'hc1222870, 32'hc070f4ce, 32'hc0d93420};
test_bias[3114:3114] = '{32'hc2a280be};
test_output[3114:3114] = '{32'hc5872f92};
test_input[24920:24927] = '{32'h42627709, 32'hc13eed7f, 32'hc1309762, 32'hc2c0287a, 32'hc226903a, 32'hc1ecf0d4, 32'hc24c36bc, 32'hc29762ab};
test_weights[24920:24927] = '{32'hc23bee33, 32'h429374e4, 32'h411ae380, 32'hc25964d7, 32'hc2771c13, 32'hc2487d26, 32'h42b2894e, 32'h41ef82e4};
test_bias[3115:3115] = '{32'hc27ea968};
test_output[3115:3115] = '{32'hc49ce5b9};
test_input[24928:24935] = '{32'hc2c7aece, 32'hc2a19f65, 32'h4219fa6f, 32'hc059396a, 32'hc2790971, 32'h4220e971, 32'hc1fa3cb3, 32'h42829450};
test_weights[24928:24935] = '{32'h426595f3, 32'hc2304a8d, 32'hc0c19fae, 32'hc19014a7, 32'hc27cbf02, 32'hc2020432, 32'h42bac947, 32'h41ac184e};
test_bias[3116:3116] = '{32'h427b22ec};
test_output[3116:3116] = '{32'hc4920cb9};
test_input[24936:24943] = '{32'h427e2124, 32'hc204d185, 32'h4213912f, 32'h41f0be73, 32'h428805c4, 32'h4284929e, 32'h423f87df, 32'hc2a19c7a};
test_weights[24936:24943] = '{32'h42891907, 32'h42b49351, 32'hc1b86821, 32'h3f4d877c, 32'hc228b5e4, 32'h41b077f8, 32'h402a7db8, 32'hc1a67d6a};
test_bias[3117:3117] = '{32'hc2340dc4};
test_output[3117:3117] = '{32'h445e2dac};
test_input[24944:24951] = '{32'h42897875, 32'hc21d5a2f, 32'h41a00028, 32'hc2a5eba2, 32'h41cdda83, 32'hc243ef02, 32'hc2b7b31a, 32'hc293e653};
test_weights[24944:24951] = '{32'hc155ccef, 32'h410b3a46, 32'h42a228fc, 32'hc23a4bcf, 32'hc2b450cc, 32'h423e9bfd, 32'hc2822743, 32'h42813efb};
test_bias[3118:3118] = '{32'hc0d0a3b7};
test_output[3118:3118] = '{32'h443e9b2b};
test_input[24952:24959] = '{32'hc19813ee, 32'hc285b7a7, 32'h42023b60, 32'h4238e464, 32'hc264450f, 32'hc25eed50, 32'h422c086a, 32'h42a35f96};
test_weights[24952:24959] = '{32'hc28a4f43, 32'h42343a4c, 32'hc2588fe4, 32'hc009a55c, 32'h425358aa, 32'hc27b5d3f, 32'hc113f281, 32'h40fb4e7d};
test_bias[3119:3119] = '{32'hc25eff43};
test_output[3119:3119] = '{32'hc5344e12};
test_input[24960:24967] = '{32'h40b79a18, 32'h41a26566, 32'hc2b5b6e3, 32'h42b7e6a5, 32'h42a13481, 32'hc1c0d454, 32'hc18bfa65, 32'h405d03dc};
test_weights[24960:24967] = '{32'h429050ea, 32'h42a43bfd, 32'hc29ec6c4, 32'h4282ff6c, 32'h41956a91, 32'hc206c554, 32'hc11712a5, 32'hc1b57b53};
test_bias[3120:3120] = '{32'h42841b54};
test_output[3120:3120] = '{32'h468af61a};
test_input[24968:24975] = '{32'hc2b31605, 32'h42aebc99, 32'hc2026629, 32'hc1d817c4, 32'hc28daca5, 32'hc217b3cb, 32'hc28abc73, 32'h4126b5b8};
test_weights[24968:24975] = '{32'hc22180e3, 32'hc26bd7ec, 32'h42313c6e, 32'h40a60c1e, 32'hc1403958, 32'h42baf3b0, 32'h4222c3ee, 32'h428ca51b};
test_bias[3121:3121] = '{32'hc2306f2f};
test_output[3121:3121] = '{32'hc5f865d1};
test_input[24976:24983] = '{32'h425acb5c, 32'hc2aee3b2, 32'hc1e826f3, 32'hc2a6f209, 32'hc2b26d1f, 32'h42a974bf, 32'hc2452aec, 32'hc1afb04a};
test_weights[24976:24983] = '{32'h4148939e, 32'hc08f7e75, 32'h4295be13, 32'h42a6db3a, 32'hbff5554c, 32'hc2444c91, 32'h41d15c63, 32'h4208d959};
test_bias[3122:3122] = '{32'h4221fc97};
test_output[3122:3122] = '{32'hc65b7ab6};
test_input[24984:24991] = '{32'h4293661c, 32'hc10a89b2, 32'h421c2c73, 32'h42b8cf74, 32'hc2649233, 32'h40a0ecd9, 32'hc182dfc0, 32'hc25d428a};
test_weights[24984:24991] = '{32'h42736814, 32'hc25ee683, 32'h42b425c8, 32'hc1bb1197, 32'hc2843e5a, 32'hc287e16d, 32'h4184b868, 32'hc295b875};
test_bias[3123:3123] = '{32'h421f3262};
test_output[3123:3123] = '{32'h46559510};
test_input[24992:24999] = '{32'hc25c5148, 32'hc25c47ac, 32'h3f4632df, 32'hc2962e4f, 32'hc19f325b, 32'h429857b8, 32'hc0bbdacf, 32'h41f7ad82};
test_weights[24992:24999] = '{32'h42b81104, 32'hc2764086, 32'h417f43a6, 32'hc10282ca, 32'h42b2cf13, 32'h426786de, 32'hc21648f5, 32'h42759d56};
test_bias[3124:3124] = '{32'h41b38389};
test_output[3124:3124] = '{32'h45687daf};
test_input[25000:25007] = '{32'h414b9532, 32'hc2be898f, 32'h42c0ab21, 32'h42b56c5b, 32'h42adabc7, 32'h425aa388, 32'hc27d4230, 32'h42a603a3};
test_weights[25000:25007] = '{32'hc15f7a13, 32'hc278fdcc, 32'hc1ee65b2, 32'hc2afa7e0, 32'h4282e264, 32'h42b1e557, 32'hc207da23, 32'hc21bae13};
test_bias[3125:3125] = '{32'hc2c015f1};
test_output[3125:3125] = '{32'h4585d87c};
test_input[25008:25015] = '{32'h4188780d, 32'h4000952f, 32'h4233dd4e, 32'hc2069d3b, 32'h4261e4a8, 32'h41ab4189, 32'hc19dc372, 32'h421516ee};
test_weights[25008:25015] = '{32'hc2786d70, 32'h42a690ec, 32'h411bb8f3, 32'hc289ebeb, 32'h42a68ed2, 32'hc03ce0f3, 32'hc225ab70, 32'hc218df4e};
test_bias[3126:3126] = '{32'hc2642a6e};
test_output[3126:3126] = '{32'h45b68b1e};
test_input[25016:25023] = '{32'h427de832, 32'h41aeb875, 32'hc29a7e57, 32'hc2412f43, 32'hc25c8da7, 32'h416b8264, 32'hc2233019, 32'hc26d2485};
test_weights[25016:25023] = '{32'hc29a983c, 32'h41cb5b8c, 32'h42b8785c, 32'h41bef5bd, 32'h3f37106d, 32'h42899427, 32'hc23fd67f, 32'hc0cb0993};
test_bias[3127:3127] = '{32'hc2c297ca};
test_output[3127:3127] = '{32'hc6133222};
test_input[25024:25031] = '{32'hc2bfe24c, 32'h4280936a, 32'hc28c93ba, 32'h412a544a, 32'hc2aa142f, 32'hc282e1bd, 32'h4290090c, 32'hc29f7007};
test_weights[25024:25031] = '{32'h41e5e2c9, 32'h4082b3a6, 32'hc2c10833, 32'h42b8da54, 32'h42c0b14b, 32'h4288aca3, 32'h41dfd203, 32'hc17380b3};
test_bias[3128:3128] = '{32'h425010e4};
test_output[3128:3128] = '{32'hc5807d0e};
test_input[25032:25039] = '{32'h4113bd63, 32'hc2a0a04b, 32'hc2c4127a, 32'hc28d6514, 32'hc1fc90f6, 32'h41e758d4, 32'h41060879, 32'hc0f30ee4};
test_weights[25032:25039] = '{32'hc15fd599, 32'h42567af6, 32'hc243d294, 32'h428a21ec, 32'h419f7586, 32'h429a78b9, 32'h3f181a04, 32'h410fb03e};
test_bias[3129:3129] = '{32'hc2b3de6d};
test_output[3129:3129] = '{32'hc53fbdf9};
test_input[25040:25047] = '{32'hc168125b, 32'h428f59ab, 32'hbfc6bc4a, 32'h4169541c, 32'h41c81816, 32'h418a460e, 32'hc293714e, 32'hc20c2430};
test_weights[25040:25047] = '{32'h42adaf78, 32'h42a11be4, 32'hc29a4c2b, 32'h423099db, 32'h408f8b05, 32'h4242533d, 32'hc22981c3, 32'hc28641bb};
test_bias[3130:3130] = '{32'hc1f43467};
test_output[3130:3130] = '{32'h46366c41};
test_input[25048:25055] = '{32'h4081545f, 32'hc0f29c50, 32'hc24cd37f, 32'h41e46765, 32'h42a041d0, 32'hc0ca3bdb, 32'h428f42e3, 32'h42abca21};
test_weights[25048:25055] = '{32'hc23df3d4, 32'h4250452a, 32'h407bba02, 32'h41e7d339, 32'hc1c602c3, 32'h428187b5, 32'h420e3550, 32'h4254792d};
test_bias[3131:3131] = '{32'hc0ccf855};
test_output[3131:3131] = '{32'h45946baf};
test_input[25056:25063] = '{32'h422900d9, 32'h42be6d7e, 32'hc2bdd54f, 32'hc23c6656, 32'h41f59046, 32'hc2637a3c, 32'hc06552fc, 32'hc0eb973d};
test_weights[25056:25063] = '{32'hc18cf68d, 32'h41b9353c, 32'hc2121678, 32'hc27160cd, 32'hc251b605, 32'h4208f61c, 32'hc1d7851b, 32'hc1546bd1};
test_bias[3132:3132] = '{32'hc2b6df6c};
test_output[3132:3132] = '{32'h4586d733};
test_input[25064:25071] = '{32'hc20b2ae3, 32'h42641bdb, 32'hc299005a, 32'h4209f0a2, 32'h4294b648, 32'hc27bb126, 32'hc24fb11f, 32'hc26fec4f};
test_weights[25064:25071] = '{32'h421e53b5, 32'h413ca3b5, 32'h427e606a, 32'h42c0681e, 32'hc1061809, 32'h423fc827, 32'h3fd771f3, 32'hc21cd82f};
test_bias[3133:3133] = '{32'h42994d00};
test_output[3133:3133] = '{32'hc55df122};
test_input[25072:25079] = '{32'h41e19903, 32'h41f281a5, 32'h41842a96, 32'h42822702, 32'h421a8ff9, 32'h42b89d57, 32'h42a0037b, 32'hc24e9ad7};
test_weights[25072:25079] = '{32'hc2996905, 32'h40325b45, 32'hc1e543ef, 32'hc28c6d29, 32'h41a218d4, 32'hc1b4a5fa, 32'h42bc88ae, 32'h42570ff4};
test_bias[3134:3134] = '{32'h4295d3ab};
test_output[3134:3134] = '{32'hc55fed97};
test_input[25080:25087] = '{32'h42bcf981, 32'h42c5dcc6, 32'h41d123cf, 32'h41bbb61f, 32'hc2a7542a, 32'h42b797f1, 32'hc294d008, 32'hc22c06d9};
test_weights[25080:25087] = '{32'hc2a31c86, 32'hc2a0d16d, 32'h41f48bac, 32'h429f3eb4, 32'hc1f488fa, 32'hc1c3adfa, 32'hc2567bf9, 32'hbfdffbc2};
test_bias[3135:3135] = '{32'hc2845849};
test_output[3135:3135] = '{32'hc607aadb};
test_input[25088:25095] = '{32'h4005fd3a, 32'h4225287f, 32'h41e82faa, 32'h424df355, 32'h42c4191b, 32'h424cf239, 32'hc2c4d6b0, 32'hc21d6eb0};
test_weights[25088:25095] = '{32'hc1dbb141, 32'h428eb2ae, 32'hc2af18a2, 32'hc2212a5b, 32'h420ad54b, 32'hc23cbb66, 32'h429c5f6a, 32'h40f1a34b};
test_bias[3136:3136] = '{32'h41951b51};
test_output[3136:3136] = '{32'hc6082bd1};
test_input[25096:25103] = '{32'hc2af8b39, 32'h41232115, 32'hc09bcc49, 32'hc28d83dc, 32'h4281cc29, 32'hc21672b6, 32'hc2b319cb, 32'h423fdd81};
test_weights[25096:25103] = '{32'hc2c79e4e, 32'h42860ac5, 32'hc17fefbf, 32'hc14fb45c, 32'h429ab104, 32'hc282626b, 32'hc242f3eb, 32'h4116eb0c};
test_bias[3137:3137] = '{32'h41edf2e6};
test_output[3137:3137] = '{32'h46b1cd15};
test_input[25104:25111] = '{32'h4185c083, 32'hc2403de2, 32'h4110a818, 32'h42c75706, 32'hc288c083, 32'hc23f8e48, 32'h41afde60, 32'hc1e16af6};
test_weights[25104:25111] = '{32'hc197cd35, 32'hc2a84d33, 32'h420ab63e, 32'h420810a5, 32'hc2bc4326, 32'hc2b74c9b, 32'hc2b37512, 32'h4240e24c};
test_bias[3138:3138] = '{32'h4219b731};
test_output[3138:3138] = '{32'h4669cdd1};
test_input[25112:25119] = '{32'hc1784ed6, 32'hc1fb880e, 32'h42acdec4, 32'h419f90a6, 32'hc2348d5f, 32'h41a4d615, 32'hc064c245, 32'h420bb1cf};
test_weights[25112:25119] = '{32'h429934fb, 32'h4247241d, 32'h3f1fb975, 32'hc29f0ef0, 32'h41bb944a, 32'h42576391, 32'h427c1e47, 32'hc197bc09};
test_bias[3139:3139] = '{32'h42ad6929};
test_output[3139:3139] = '{32'hc59d629e};
test_input[25120:25127] = '{32'h42ae5801, 32'hc2b1da2f, 32'hc20f5204, 32'hc0751d15, 32'hc2500c99, 32'hc292936d, 32'hc2b02d04, 32'h42c5dc60};
test_weights[25120:25127] = '{32'h41f53540, 32'h428c9434, 32'h4266825c, 32'hc212cb94, 32'hc28c327f, 32'hc22a7619, 32'h4291df84, 32'hc11f1350};
test_bias[3140:3140] = '{32'hc294b2f9};
test_output[3140:3140] = '{32'hc5c243eb};
test_input[25128:25135] = '{32'h42a6e364, 32'h42c44a10, 32'h42bf1811, 32'h4250a04c, 32'hc2584c8d, 32'h41ea9b25, 32'h41ac2d48, 32'hc24e7757};
test_weights[25128:25135] = '{32'hc285bc1d, 32'h42a395bf, 32'h42c5d282, 32'hc26fda6e, 32'hc0b18896, 32'h4293b607, 32'h4274fa26, 32'hc0d6af30};
test_bias[3141:3141] = '{32'h41f010d1};
test_output[3141:3141] = '{32'h464a0d0d};
test_input[25136:25143] = '{32'hc210a110, 32'h410af5a2, 32'h4130f9ef, 32'h428074a2, 32'hc28d1160, 32'hc22b131e, 32'h42ba05f4, 32'h42ad7e2b};
test_weights[25136:25143] = '{32'hc250bdc6, 32'h42531fc4, 32'h42c22ac6, 32'h41c49d83, 32'hc2a53f26, 32'hc1f31b4b, 32'hc22923a8, 32'h4269671c};
test_bias[3142:3142] = '{32'hbd8cf523};
test_output[3142:3142] = '{32'h464f16e9};
test_input[25144:25151] = '{32'h41018efa, 32'hc0f35157, 32'hc2a36811, 32'hc29e0849, 32'hc2a8b402, 32'h4260291e, 32'hc1d32d6f, 32'hc26171f5};
test_weights[25144:25151] = '{32'h413cbd64, 32'hc2a8fd67, 32'hc20bb5cb, 32'hc21c9e29, 32'h42299f94, 32'hc2c78305, 32'hc2c70869, 32'hc23d2b40};
test_bias[3143:3143] = '{32'hc1cf38ca};
test_output[3143:3143] = '{32'h452e0afd};
test_input[25152:25159] = '{32'h419523fe, 32'h422b9c2f, 32'h42286de1, 32'hc28277d5, 32'hc2c6d538, 32'hc2ada074, 32'h42125086, 32'h3f17a6e1};
test_weights[25152:25159] = '{32'h4245eca8, 32'h42bd1035, 32'hc18ac2c2, 32'h42c432b0, 32'hc1c21d00, 32'hc191ef20, 32'h41945114, 32'h4287730a};
test_bias[3144:3144] = '{32'hc1f92043};
test_output[3144:3144] = '{32'h451e35e8};
test_input[25160:25167] = '{32'hc26c9a1d, 32'hc2116f3b, 32'h41a90905, 32'h41daadf4, 32'hc2860bd9, 32'hc225270a, 32'h4250a958, 32'hbf430105};
test_weights[25160:25167] = '{32'h42985b49, 32'hc29c765e, 32'h429f3dc8, 32'hc1e417f4, 32'hc2a8cdf7, 32'h42b77b13, 32'hc19d394a, 32'hbf47c48a};
test_bias[3145:3145] = '{32'hc1b36634};
test_output[3145:3145] = '{32'h427dcb67};
test_input[25168:25175] = '{32'h42a06883, 32'h429a948a, 32'hc1bd3b00, 32'h421b206c, 32'hc1d3b147, 32'hc25ca8b1, 32'hc2c69048, 32'hc2b93338};
test_weights[25168:25175] = '{32'h422b4702, 32'h42700662, 32'hc2922874, 32'hc2b142aa, 32'h42275132, 32'h42022bf9, 32'h42acbfb0, 32'hc16f8da5};
test_bias[3146:3146] = '{32'h429b0282};
test_output[3146:3146] = '{32'hc5642077};
test_input[25176:25183] = '{32'h4277a6ab, 32'h423f24d5, 32'hc1c05df3, 32'hc2673900, 32'h4110656c, 32'h4257c2fd, 32'hc1e4e3c0, 32'h427a5fd6};
test_weights[25176:25183] = '{32'h42c4600c, 32'h421b4d81, 32'hbfe5539f, 32'h4264536b, 32'h42794c36, 32'hc2290143, 32'hc1fef20a, 32'hc1f22aa1};
test_bias[3147:3147] = '{32'hc26423b2};
test_output[3147:3147] = '{32'h44f027d4};
test_input[25184:25191] = '{32'hc265f082, 32'h429bdd19, 32'h4255ab99, 32'hc25d57f7, 32'hc19dee3b, 32'h42082f8a, 32'h423472c1, 32'hc236291b};
test_weights[25184:25191] = '{32'hc219f789, 32'h42a369c2, 32'hc2992410, 32'h4272b312, 32'hc191050d, 32'hc2b80ff1, 32'hc2bf0120, 32'h428039af};
test_bias[3148:3148] = '{32'h4226b83b};
test_output[3148:3148] = '{32'hc609f50f};
test_input[25192:25199] = '{32'h41cbcf12, 32'hc1029efe, 32'hc28750bc, 32'hc22bc809, 32'h423d7b88, 32'hbf1168f0, 32'hc2b3e0b0, 32'hc2536de4};
test_weights[25192:25199] = '{32'hc2a96d2b, 32'h40c96846, 32'hc254881d, 32'h415a1bdb, 32'hc23bf490, 32'h411ef6cd, 32'h41eab553, 32'hc2ab44e1};
test_bias[3149:3149] = '{32'hc10203da};
test_output[3149:3149] = '{32'h43dffac4};
test_input[25200:25207] = '{32'hc229fe94, 32'h424cb7f2, 32'h41019bcb, 32'hc1ab44a1, 32'hc2b958bb, 32'h428e50e2, 32'hc2539a04, 32'hc2a58b29};
test_weights[25200:25207] = '{32'hc2a1e7d8, 32'h41346758, 32'hc2a52fdb, 32'h413c801d, 32'h4201be74, 32'hc12e1f9c, 32'hc199d213, 32'hc290b1eb};
test_bias[3150:3150] = '{32'h4199ebc9};
test_output[3150:3150] = '{32'h45c62468};
test_input[25208:25215] = '{32'hc14820a3, 32'h42956472, 32'hc1710fe9, 32'hc2ad43a0, 32'h4295d91a, 32'hc168a88e, 32'hc250a9a9, 32'h401cc879};
test_weights[25208:25215] = '{32'hc243d9b5, 32'hc28f3dcd, 32'hc2216a38, 32'hc21d54e0, 32'h42b54ecb, 32'h42785fc9, 32'hc1970cab, 32'h427ba849};
test_bias[3151:3151] = '{32'hbfc28783};
test_output[3151:3151] = '{32'h45c50735};
test_input[25216:25223] = '{32'h4289dc9f, 32'h418109d8, 32'h427b450f, 32'hc2bad9ba, 32'hc27eba30, 32'hc185d63c, 32'h429d6de5, 32'hc11c7325};
test_weights[25216:25223] = '{32'h425043d4, 32'hc1ca5a25, 32'h41e61143, 32'hc1da47b3, 32'h42a54e6d, 32'h4296e934, 32'h42b8ef76, 32'h42871f2a};
test_bias[3152:3152] = '{32'hc1193f43};
test_output[3152:3152] = '{32'h45ee192a};
test_input[25224:25231] = '{32'hc21a7267, 32'h423fe2a7, 32'h42831895, 32'hc23aadde, 32'h42bbb141, 32'h424fb040, 32'hc29bf991, 32'hc2994dbf};
test_weights[25224:25231] = '{32'hc100bfb2, 32'h429740f5, 32'hc289b560, 32'h426c7dff, 32'hc26fa973, 32'hc2a58fd1, 32'h42525744, 32'h428bc319};
test_bias[3153:3153] = '{32'h41136b34};
test_output[3153:3153] = '{32'hc6b15e5c};
test_input[25232:25239] = '{32'hc2ac2761, 32'hc2a491b2, 32'h424b8ba2, 32'h42bd4b80, 32'h42aaf459, 32'h4289c33f, 32'h42a6aaa5, 32'hc26cdcc9};
test_weights[25232:25239] = '{32'h4267484e, 32'h4290ff4b, 32'h428fcf69, 32'h420d49fb, 32'hc202e204, 32'h4299a80d, 32'h42704dd0, 32'h42bd77e8};
test_bias[3154:3154] = '{32'hc1c8d87a};
test_output[3154:3154] = '{32'hc5019c0b};
test_input[25240:25247] = '{32'hc2800e05, 32'h4281b251, 32'hc2a08cc2, 32'h41ba30ac, 32'h42c5798f, 32'h42b1c800, 32'hc2329e00, 32'h428a4e69};
test_weights[25240:25247] = '{32'hc287c5ec, 32'hc02cf7ec, 32'hc2c5c735, 32'h426721c8, 32'h4286e571, 32'hc2a26315, 32'h42a60532, 32'hc1195ff9};
test_bias[3155:3155] = '{32'h42771e5f};
test_output[3155:3155] = '{32'h460633a7};
test_input[25248:25255] = '{32'hc1184d94, 32'h428c633f, 32'h423cc42a, 32'hc28ba56d, 32'hc2c09a58, 32'hc09431e1, 32'h4199df3c, 32'hc26d3c0c};
test_weights[25248:25255] = '{32'h42988445, 32'h41ab8a30, 32'h42c6ab0e, 32'h42c67ebf, 32'h42a3f880, 32'h41b4a8d2, 32'h3da68119, 32'h42986224};
test_bias[3156:3156] = '{32'hc2849024};
test_output[3156:3156] = '{32'hc65b78f7};
test_input[25256:25263] = '{32'h427b9633, 32'hc20da98b, 32'h4269ea72, 32'h417274d7, 32'h42994964, 32'h428a7286, 32'hc253eeb5, 32'h421d09fb};
test_weights[25256:25263] = '{32'hc18df118, 32'hc282f394, 32'h41d5d556, 32'hc2452c7e, 32'hc2aed805, 32'h4237f27f, 32'h42976f60, 32'h41d1a5aa};
test_bias[3157:3157] = '{32'hc236d35b};
test_output[3157:3157] = '{32'hc58d7433};
test_input[25264:25271] = '{32'h422f6a81, 32'h42c6df3c, 32'hc2c4bb5e, 32'hc25f882a, 32'hc2c6c86e, 32'h428ea952, 32'hc229dce2, 32'hc108f613};
test_weights[25264:25271] = '{32'h42992c81, 32'h418483fa, 32'h428aa1fa, 32'hc28edb70, 32'hc2b1f4b5, 32'hc2974aa5, 32'hc1a89b99, 32'hc1ad0d79};
test_bias[3158:3158] = '{32'h42a38e29};
test_output[3158:3158] = '{32'h45d42600};
test_input[25272:25279] = '{32'h418d25b6, 32'hc255c3a1, 32'hc226e09e, 32'hc1ee59c4, 32'hc2ab1951, 32'hc20486ed, 32'h4179a70a, 32'h4275829c};
test_weights[25272:25279] = '{32'hc238567b, 32'h41dff1d5, 32'h42be9207, 32'hc1a35b47, 32'h42a34aeb, 32'hc2ae495a, 32'h42bf0592, 32'hc2b7e070};
test_bias[3159:3159] = '{32'h4244a621};
test_output[3159:3159] = '{32'hc658d415};
test_input[25280:25287] = '{32'hc2a1ea2a, 32'h42868665, 32'hc0e76e1f, 32'hc2a5f7fa, 32'hc28dd453, 32'h4298c8b5, 32'hc2a69cbc, 32'h42286242};
test_weights[25280:25287] = '{32'h422656d5, 32'hc261d436, 32'h42bfbf51, 32'hc255e37b, 32'h42ad5992, 32'h4290297b, 32'hc2937b8c, 32'h42525747};
test_bias[3160:3160] = '{32'hc2c483bf};
test_output[3160:3160] = '{32'h4583323f};
test_input[25288:25295] = '{32'h41b0e5a1, 32'h419773f9, 32'hc2a2a6f7, 32'h42a1ce69, 32'hc1ff7874, 32'h41bf4857, 32'h428784f0, 32'h42c177cd};
test_weights[25288:25295] = '{32'h4288b537, 32'h4245c60e, 32'hc1cf6ecd, 32'h400b9133, 32'hc10f9517, 32'h42a299a0, 32'hc0ba3a5d, 32'h42baae65};
test_bias[3161:3161] = '{32'h42afc927};
test_output[3161:3161] = '{32'h4675178a};
test_input[25296:25303] = '{32'hc2ae2253, 32'h425560d0, 32'h418aac4a, 32'hc2239bf7, 32'hc23d3dc0, 32'h423ec822, 32'hc2284561, 32'h42c0d364};
test_weights[25296:25303] = '{32'h42c7a2e9, 32'h411ac7c8, 32'hc26a2734, 32'h42bb17fb, 32'h42ade7c7, 32'hc2bb7005, 32'h42123090, 32'h417e5b70};
test_bias[3162:3162] = '{32'h42904786};
test_output[3162:3162] = '{32'hc6a83852};
test_input[25304:25311] = '{32'hc119e878, 32'h42a754d5, 32'h425285be, 32'hc261e315, 32'hc15d1491, 32'h414641db, 32'h41b0ecc7, 32'h420fda40};
test_weights[25304:25311] = '{32'h40426c8c, 32'hc2c07354, 32'h400bcc53, 32'hc295e9cd, 32'h3e8ccd32, 32'h4273bbb3, 32'hc2775607, 32'h41480c7b};
test_bias[3163:3163] = '{32'h417a66d7};
test_output[3163:3163] = '{32'hc572b0bb};
test_input[25312:25319] = '{32'hc2c01f56, 32'h422a5e32, 32'hc1b93fb7, 32'h42c0071c, 32'h42589d01, 32'hc08552cf, 32'h42b287af, 32'h42488346};
test_weights[25312:25319] = '{32'hc2a920e3, 32'hc238942c, 32'hc2c39305, 32'h42997ae3, 32'h42bb52b9, 32'hc20429d1, 32'h4235bc61, 32'hc179e60a};
test_bias[3164:3164] = '{32'hc2a86b0a};
test_output[3164:3164] = '{32'h46bcf960};
test_input[25320:25327] = '{32'hc29f57b4, 32'h4042a313, 32'hc225384e, 32'hc29942ac, 32'h428c9ae5, 32'hc22ac59b, 32'h42a3545f, 32'hc0c66c65};
test_weights[25320:25327] = '{32'h42a5dc8a, 32'hc220ffc1, 32'hc20fb7f7, 32'h42628c56, 32'h42242010, 32'h42a8d870, 32'h42819950, 32'hc2bc3f48};
test_bias[3165:3165] = '{32'h3eaf3eed};
test_output[3165:3165] = '{32'hc58a6be3};
test_input[25328:25335] = '{32'hc28cecd1, 32'hc291a087, 32'h3f89d3dc, 32'h41f82110, 32'h4240a0b8, 32'h428ec7ca, 32'hc2396934, 32'hc287f21e};
test_weights[25328:25335] = '{32'hc2a98141, 32'hc06163b6, 32'h426c3a42, 32'h40063b9a, 32'h40c426c6, 32'hc21ea18b, 32'hbec38afe, 32'h41e028a2};
test_bias[3166:3166] = '{32'hc195cd2e};
test_output[3166:3166] = '{32'h44ef6b17};
test_input[25336:25343] = '{32'hc28bf8b1, 32'hc2873849, 32'h40d2177d, 32'h4201bfe2, 32'hc19cd099, 32'hc1ade178, 32'h421e1e3a, 32'h42a1ae42};
test_weights[25336:25343] = '{32'hc1918d28, 32'h420316da, 32'h425d5496, 32'hc2259839, 32'h42951f0a, 32'hc260011d, 32'hc19a7138, 32'hc2a84672};
test_bias[3167:3167] = '{32'hc2bf3561};
test_output[3167:3167] = '{32'hc6198b25};
test_input[25344:25351] = '{32'hc2c3a0e3, 32'h425cd53f, 32'hc0a19450, 32'h3f858ea0, 32'hc2893772, 32'h4186dd1c, 32'h4290dd61, 32'h4298c8dc};
test_weights[25344:25351] = '{32'h42807ac4, 32'h41d5da9b, 32'hc2024f7a, 32'hc21ef6bb, 32'hc12269e4, 32'h41275d62, 32'h42ae348f, 32'h411b7807};
test_bias[3168:3168] = '{32'h426957b6};
test_output[3168:3168] = '{32'h454e1ba1};
test_input[25352:25359] = '{32'hc2521dac, 32'hc25d417b, 32'h41c04a69, 32'h422aa873, 32'h429efb57, 32'h42b849f7, 32'hc2c66369, 32'h4218a859};
test_weights[25352:25359] = '{32'h42a9babb, 32'hc08f7b5b, 32'hbe91023d, 32'h4199cc7c, 32'hc297d9b6, 32'h424f650a, 32'hc16a89bb, 32'h428887d5};
test_bias[3169:3169] = '{32'h418842f2};
test_output[3169:3169] = '{32'hc4107583};
test_input[25360:25367] = '{32'h42319abe, 32'h424982f0, 32'h42107d52, 32'h429a7d2b, 32'h40d71dd0, 32'h42a40a89, 32'h41f86d00, 32'hc2436d0c};
test_weights[25360:25367] = '{32'h42abd97f, 32'h41efefd0, 32'hc20a2421, 32'h42610869, 32'h41880e57, 32'h42563eec, 32'h41cf8c26, 32'h42564770};
test_bias[3170:3170] = '{32'h425df13a};
test_output[3170:3170] = '{32'h462e9e56};
test_input[25368:25375] = '{32'h425fd2b8, 32'hc1def832, 32'h4295cb7e, 32'hc148817c, 32'hc2b801c5, 32'h42bca2d6, 32'h3fd00a77, 32'hc21b2fad};
test_weights[25368:25375] = '{32'hc24d9ab1, 32'hc2146c6b, 32'h40bf6b5f, 32'hc204c6b1, 32'h41f6e386, 32'hc1a76c3b, 32'h4298c877, 32'hc25c2bf2};
test_bias[3171:3171] = '{32'h42b1a936};
test_output[3171:3171] = '{32'hc5572bc4};
test_input[25376:25383] = '{32'hc2c0f48a, 32'h42b67fc6, 32'h42af2b4c, 32'h4248d98d, 32'h428f0496, 32'h4122624c, 32'h4266a3e7, 32'hc2a9a0df};
test_weights[25376:25383] = '{32'hc2b5f109, 32'h4298e3c1, 32'h422a0efa, 32'h42717d57, 32'hc0701a23, 32'hc2c71a34, 32'hc1ba6b4d, 32'h41c5a4d5};
test_bias[3172:3172] = '{32'h4281bb1e};
test_output[3172:3172] = '{32'h468b7d0e};
test_input[25384:25391] = '{32'h4235b68c, 32'hc1c1228b, 32'hc2b42e56, 32'hc2704152, 32'h42ad6d5b, 32'hc2ba788a, 32'hc23c6cf2, 32'hc2164fbd};
test_weights[25384:25391] = '{32'h42780087, 32'h4286692a, 32'h419049bb, 32'h41baad4e, 32'hc2978168, 32'h42696047, 32'hc20572c2, 32'h427b07ac};
test_bias[3173:3173] = '{32'h42580d2d};
test_output[3173:3173] = '{32'hc663b63f};
test_input[25392:25399] = '{32'h4259c87b, 32'h4261cc3c, 32'hc2839818, 32'h4259f418, 32'h42a1db5d, 32'hc193d19a, 32'hc232755a, 32'h428f9c4a};
test_weights[25392:25399] = '{32'hc256ec18, 32'h424b286d, 32'h42c0bc01, 32'hc16fd719, 32'h40a1bec3, 32'hc2301db8, 32'hc1cff2a5, 32'hc2939d50};
test_bias[3174:3174] = '{32'hc00d5f57};
test_output[3174:3174] = '{32'hc61e5dfd};
test_input[25400:25407] = '{32'hc1a93937, 32'hc208a36a, 32'h4275089c, 32'h41ffbc82, 32'h422d1257, 32'h419d45e4, 32'hc27776a4, 32'hc0ff17f1};
test_weights[25400:25407] = '{32'h42520d23, 32'h42bd0329, 32'h42b1be8e, 32'hc20315c8, 32'h41009d2f, 32'hc2c68e1b, 32'hc100b0b1, 32'h4201626d};
test_bias[3175:3175] = '{32'hc210449e};
test_output[3175:3175] = '{32'hc4a7d82c};
test_input[25408:25415] = '{32'h422d1d47, 32'h42c3a102, 32'h421e399f, 32'h419233c3, 32'h41bd15a7, 32'hc1b4dc12, 32'h3ca492b3, 32'h42722ef7};
test_weights[25408:25415] = '{32'h41f9d938, 32'hc2a7c04b, 32'hc2abb4b8, 32'h42a0e771, 32'h42425392, 32'h4106fe1c, 32'h428f0cea, 32'h42bff35c};
test_bias[3176:3176] = '{32'hc08567c6};
test_output[3176:3176] = '{32'hc4fb950b};
test_input[25416:25423] = '{32'hc1c846da, 32'hc2875bdf, 32'hc2b848d5, 32'h4208c552, 32'hc261b065, 32'hc24c54a6, 32'h4282d649, 32'hc2131b42};
test_weights[25416:25423] = '{32'h40c0d1a9, 32'hc284e597, 32'h4252a1d8, 32'h428e4dc0, 32'hc28366bc, 32'hc2832742, 32'hc1ad6946, 32'hc2a1ae3f};
test_bias[3177:3177] = '{32'hc24e6536};
test_output[3177:3177] = '{32'h4623dd92};
test_input[25424:25431] = '{32'h426569a9, 32'hc29c08a2, 32'hc29770b7, 32'hc1b1fb4a, 32'h429965c3, 32'h42949995, 32'h41b2cb8a, 32'hc18995de};
test_weights[25424:25431] = '{32'h41407491, 32'hc2be5afc, 32'h418473b8, 32'h427019d3, 32'hc2af29df, 32'hc08fee15, 32'hc1dfe318, 32'hc11066ae};
test_bias[3178:3178] = '{32'h428c8fb6};
test_output[3178:3178] = '{32'hc4f0aa3a};
test_input[25432:25439] = '{32'hc2585629, 32'hc29c3f88, 32'hc28b97f1, 32'hc27d7b5e, 32'hc2342a85, 32'h429fc3f4, 32'hc2863078, 32'hc2babda4};
test_weights[25432:25439] = '{32'hc204a2d1, 32'hc25f57ec, 32'h41b813c3, 32'h41d9e6c8, 32'h42909678, 32'hc2be0706, 32'hc0ecaca9, 32'h418839a0};
test_bias[3179:3179] = '{32'h424006fc};
test_output[3179:3179] = '{32'hc60db1b1};
test_input[25440:25447] = '{32'hc0f563c2, 32'h41828115, 32'h4186b96a, 32'h402d11c1, 32'hc29a36da, 32'h424f43d0, 32'hc2573612, 32'hc2affdf6};
test_weights[25440:25447] = '{32'hc28588cb, 32'hc2bcf5f5, 32'h42799b37, 32'hc1c3d9c2, 32'hc1ccc182, 32'h3fc1ba81, 32'hc244827e, 32'h42466f9b};
test_bias[3180:3180] = '{32'hc127ef68};
test_output[3180:3180] = '{32'h43895414};
test_input[25448:25455] = '{32'hc23bbf88, 32'h422a1bde, 32'hc2b0812c, 32'h42500b36, 32'h428554cc, 32'h42323a9b, 32'hc2a8fd15, 32'hc232fc92};
test_weights[25448:25455] = '{32'hc1b89d1f, 32'h426ff558, 32'h42b85d77, 32'h42ad8a0b, 32'h42b86362, 32'hc2b8f810, 32'hc2c0878f, 32'hc19e7151};
test_bias[3181:3181] = '{32'hc288cabf};
test_output[3181:3181] = '{32'h462bb3de};
test_input[25456:25463] = '{32'hc2238f9e, 32'h423a21fa, 32'h4297615f, 32'h42b9ff00, 32'hc23ad6d7, 32'h41b00c82, 32'hc20b1086, 32'h42ada4cc};
test_weights[25456:25463] = '{32'h40fbcd29, 32'hc2a7ef25, 32'h42c1221f, 32'h42314046, 32'h4272b167, 32'h4288363e, 32'h42c434ef, 32'h41a44a0b};
test_bias[3182:3182] = '{32'h418e875a};
test_output[3182:3182] = '{32'h4584ffcb};
test_input[25464:25471] = '{32'h4278b8f1, 32'h42c73701, 32'hc25bab77, 32'hc2389ca9, 32'h428a2db9, 32'h42abadd7, 32'h425fb46e, 32'hc2873091};
test_weights[25464:25471] = '{32'hc1050023, 32'h427800a7, 32'hc1243adf, 32'h424da4f8, 32'hc284adff, 32'h420a7f59, 32'hc17030ef, 32'h429da5d1};
test_bias[3183:3183] = '{32'h41899943};
test_output[3183:3183] = '{32'hc5747eb8};
test_input[25472:25479] = '{32'hc26a6291, 32'hc0b58fa9, 32'h4244e5ba, 32'h422ebfaf, 32'h42870166, 32'hc2659cb1, 32'hc272a54c, 32'hc207e3d1};
test_weights[25472:25479] = '{32'hc2c12923, 32'h40a5d563, 32'hc29d6a30, 32'hc2ad1540, 32'hbfd7f7f7, 32'hc29ca68b, 32'h4297bc73, 32'hc2940f90};
test_bias[3184:3184] = '{32'hc1b158dd};
test_output[3184:3184] = '{32'h43778b61};
test_input[25480:25487] = '{32'hc26384d2, 32'hc2b9f640, 32'hc1937873, 32'h4225dc3c, 32'h428bdbd2, 32'h425c92c5, 32'hc106e30d, 32'hc1834bd8};
test_weights[25480:25487] = '{32'h429c965f, 32'h4295f336, 32'hc299be6a, 32'hc28f6127, 32'h42767110, 32'hc0367c33, 32'h42bc2278, 32'hc23a9c98};
test_bias[3185:3185] = '{32'h426eda54};
test_output[3185:3185] = '{32'hc609729c};
test_input[25488:25495] = '{32'h41ab41c9, 32'h4223297f, 32'hc2c4e9a3, 32'hc274640e, 32'h42b2e6d0, 32'hc282b971, 32'h428a26fb, 32'hc2964c0d};
test_weights[25488:25495] = '{32'hc240d01c, 32'h424363f9, 32'hc19d11c9, 32'hc2b8ab3e, 32'h4295a729, 32'hc10b529f, 32'hc196fd1e, 32'h42b80b36};
test_bias[3186:3186] = '{32'h3f0ca9b2};
test_output[3186:3186] = '{32'h45ecd8a0};
test_input[25496:25503] = '{32'h428f08cb, 32'hc2898e4f, 32'h42ad448a, 32'h428f54d4, 32'hc2b2db82, 32'hc20c940d, 32'hc1fc1faf, 32'hc287908b};
test_weights[25496:25503] = '{32'hc176f41c, 32'h422378a0, 32'hc152ee6f, 32'h42a54e98, 32'hc2bd9866, 32'hc23dc14b, 32'h42690dab, 32'hc199117c};
test_bias[3187:3187] = '{32'hc29347b5};
test_output[3187:3187] = '{32'h46227a5f};
test_input[25504:25511] = '{32'hc1bd3338, 32'h420b41ab, 32'hc2961398, 32'hc283bd78, 32'hc2c5cb32, 32'hc26c6d1c, 32'hc2ad186d, 32'h425357ec};
test_weights[25504:25511] = '{32'hc2bfb867, 32'hc22ee65f, 32'hc244a8d4, 32'hc0b189fb, 32'h4275a02e, 32'h4249b305, 32'hc2b785e2, 32'hc1a694a4};
test_bias[3188:3188] = '{32'hc2a17dff};
test_output[3188:3188] = '{32'h451cb073};
test_input[25512:25519] = '{32'hc279ae76, 32'h4201efd7, 32'h4297751c, 32'hc2a20f5a, 32'h41ad2d90, 32'hc1cfcad1, 32'hc1243865, 32'hc2073c59};
test_weights[25512:25519] = '{32'h42c0a188, 32'h42255fe2, 32'h425888a8, 32'h42a4069a, 32'hc114ee64, 32'h42a593af, 32'hc15befc0, 32'h425a91e7};
test_bias[3189:3189] = '{32'hc242fcd7};
test_output[3189:3189] = '{32'hc630e7f5};
test_input[25520:25527] = '{32'h421c99e1, 32'h418c8bf7, 32'hc1c3415d, 32'hc285a1b5, 32'h42a8311f, 32'hc2148c39, 32'hc22c9605, 32'h429e1894};
test_weights[25520:25527] = '{32'hc232f446, 32'hc22c9d79, 32'hc2b4f21d, 32'hc288f310, 32'hc2411717, 32'h42064aa6, 32'h3fcdef9d, 32'hc24d553c};
test_bias[3190:3190] = '{32'hc2988ea0};
test_output[3190:3190] = '{32'hc5a3a0e7};
test_input[25528:25535] = '{32'h4243e1bb, 32'hc0c51a07, 32'h42a24ae5, 32'hc26a30e8, 32'h423fd370, 32'hc11f9707, 32'h42b8f4b4, 32'hc29962df};
test_weights[25528:25535] = '{32'h41ab13c1, 32'h42b4cbfb, 32'h423ee482, 32'hc29724f7, 32'h421bfef7, 32'hc1eabf72, 32'h415a687f, 32'h423998c8};
test_bias[3191:3191] = '{32'hc292361d};
test_output[3191:3191] = '{32'h46061506};
test_input[25536:25543] = '{32'h417d69bc, 32'hc16be6a9, 32'hc1bd208f, 32'h421b3d17, 32'h42ba0ddd, 32'h42a1b87f, 32'hc2ba7743, 32'h42aa5c9f};
test_weights[25536:25543] = '{32'hc269500a, 32'hc29307dd, 32'hc21483d2, 32'hc0f58274, 32'h4236c779, 32'hc28d9aa0, 32'h4203b24b, 32'hc1de7f39};
test_bias[3192:3192] = '{32'hc2871318};
test_output[3192:3192] = '{32'hc5c302d1};
test_input[25544:25551] = '{32'h421a8ce0, 32'hc2384833, 32'h4196226e, 32'h429fc73b, 32'hc2b8be06, 32'hc2559973, 32'hc0f7d6e6, 32'h42ab35d9};
test_weights[25544:25551] = '{32'hc24f2594, 32'h42026d4e, 32'h423513c7, 32'hc2142ce8, 32'h3fc710d1, 32'h4285d1d0, 32'h428b4f7d, 32'h42c6357a};
test_bias[3193:3193] = '{32'hc2bd3c01};
test_output[3193:3193] = '{32'hc4b8faa8};
test_input[25552:25559] = '{32'h42644fed, 32'h4251aeb2, 32'hc2951e7c, 32'h41f9950e, 32'hc2a11a93, 32'hc18c7390, 32'h427bfdf6, 32'hc2a63d6b};
test_weights[25552:25559] = '{32'hc2a225c6, 32'hc2b1602e, 32'h3f23adfb, 32'h3d26b160, 32'h42ac6409, 32'h418d5a81, 32'h423d4eb8, 32'h420a5920};
test_bias[3194:3194] = '{32'h42335633};
test_output[3194:3194] = '{32'hc68051e9};
test_input[25560:25567] = '{32'hc2837e44, 32'hc2893dd8, 32'hc140a3c4, 32'hbfcb2f1a, 32'hc157b5b5, 32'h42c0393a, 32'h42729ce2, 32'hc27cadc5};
test_weights[25560:25567] = '{32'h4265b674, 32'hc28dad69, 32'hc2ab134b, 32'h41cc78b3, 32'hc0163b9c, 32'hc2a8d402, 32'hc1d4d8e7, 32'hc18efd0f};
test_bias[3195:3195] = '{32'h4200d6cb};
test_output[3195:3195] = '{32'hc5c9db2c};
test_input[25568:25575] = '{32'h424c5a29, 32'h428244ca, 32'h4151e2c9, 32'hc205badb, 32'h4208381e, 32'hc20fc5b3, 32'h42a5e5c9, 32'hc210c0bd};
test_weights[25568:25575] = '{32'h405e922d, 32'hc265f417, 32'hc1b81c74, 32'h41b065dd, 32'hc22601b9, 32'hc299b1a7, 32'h41408d75, 32'h42382ba6};
test_bias[3196:3196] = '{32'h427d849c};
test_output[3196:3196] = '{32'hc5715a85};
test_input[25576:25583] = '{32'h41f7a926, 32'hc2be4b76, 32'h42589c94, 32'h42b9cf96, 32'h42acbe9e, 32'hc288a238, 32'hc2249d62, 32'h3fb00355};
test_weights[25576:25583] = '{32'hc21ade2b, 32'hc2a7ef4e, 32'hc26bd40d, 32'hc2bb3176, 32'hc2c1ff9e, 32'h41202f1d, 32'hc1eade2c, 32'h42a9a6e4};
test_bias[3197:3197] = '{32'h40c881f2};
test_output[3197:3197] = '{32'hc6487214};
test_input[25584:25591] = '{32'hc077a682, 32'h418c74cd, 32'h4295935e, 32'hc2b32060, 32'hc2b37adc, 32'h4254b615, 32'hc1dba75f, 32'hc10a22e6};
test_weights[25584:25591] = '{32'h4211e68d, 32'hc2132565, 32'h4226de2f, 32'hc24daf39, 32'h41c96da8, 32'h41923bcd, 32'hc2bab123, 32'h4161b272};
test_bias[3198:3198] = '{32'hc13d6eae};
test_output[3198:3198] = '{32'h45fc81e4};
test_input[25592:25599] = '{32'h42afbe62, 32'h429a6bc3, 32'hc2602b81, 32'h42be3c94, 32'hc2871066, 32'h4101339c, 32'h424ad2b7, 32'hc2b24e6c};
test_weights[25592:25599] = '{32'hc08dba30, 32'hc277de8e, 32'hc2a6dfa7, 32'h428b4cf5, 32'h41333276, 32'hc2b8b9a1, 32'hc232f362, 32'hc2867576};
test_bias[3199:3199] = '{32'h417b33be};
test_output[3199:3199] = '{32'h4602b85d};
test_input[25600:25607] = '{32'h429fe72f, 32'h422df715, 32'hc2265c53, 32'hc285504a, 32'hc1443561, 32'hc24bf87f, 32'h4299dc94, 32'h4191bc4b};
test_weights[25600:25607] = '{32'h4129dae0, 32'h4270ea67, 32'hc1af2d97, 32'hc2c1769c, 32'h421b0d50, 32'h4241e6b8, 32'h4192abbd, 32'hc26d1284};
test_bias[3200:3200] = '{32'hc27f8916};
test_output[3200:3200] = '{32'h45fe92e6};
test_input[25608:25615] = '{32'hc2beffec, 32'h42af7675, 32'hc1c8e97b, 32'hc2126f6b, 32'hc22a670c, 32'hc24b8fcd, 32'hc28cf119, 32'hc2350cfc};
test_weights[25608:25615] = '{32'h41f9040a, 32'h4232829f, 32'h42b8da0e, 32'hc273d558, 32'h423fe222, 32'h4115af8f, 32'h42a7b1b1, 32'hc1cf868b};
test_bias[3201:3201] = '{32'h428f9fa0};
test_output[3201:3201] = '{32'hc5c5cbb3};
test_input[25616:25623] = '{32'hc2abd529, 32'h41c07c3f, 32'hc228b84b, 32'hc27e3fa8, 32'h426f816d, 32'hc282f962, 32'hc2bf2149, 32'h428526be};
test_weights[25616:25623] = '{32'hc28440bc, 32'hc12afcfe, 32'hc15322ec, 32'hc13cd5cf, 32'hc0b5af3d, 32'hc2558337, 32'h410c198b, 32'h42347b90};
test_bias[3202:3202] = '{32'h42516494};
test_output[3202:3202] = '{32'h463d2870};
test_input[25624:25631] = '{32'h421a02f5, 32'hc1c8f4c7, 32'h41e5f1b2, 32'h42c253b0, 32'hc280a438, 32'h4298e1d4, 32'hc14273d7, 32'h40004fdc};
test_weights[25624:25631] = '{32'h424f61ff, 32'hc1fe4170, 32'h4126823c, 32'h42b70201, 32'h42bbdbde, 32'hc253d17e, 32'hc28925f9, 32'h421681ec};
test_bias[3203:3203] = '{32'h42ae0d0e};
test_output[3203:3203] = '{32'h4534add3};
test_input[25632:25639] = '{32'h41adb092, 32'hc248e2f0, 32'h42021ed4, 32'h420f232e, 32'h41f8dd89, 32'hc2aee81b, 32'hc2468ee1, 32'h426e11cb};
test_weights[25632:25639] = '{32'hc282bc8c, 32'h41e9c88b, 32'h4247bf09, 32'h41ed4143, 32'h4283ffe5, 32'h42bd1412, 32'hc1ae1805, 32'h429668e4};
test_bias[3204:3204] = '{32'hc1e11bf2};
test_output[3204:3204] = '{32'hc45dec16};
test_input[25640:25647] = '{32'hc12c359e, 32'hc19df6cd, 32'hc22437ef, 32'h42be30e9, 32'hc287464a, 32'hc20f51c3, 32'hc1f47915, 32'h42a35780};
test_weights[25640:25647] = '{32'hc1c495aa, 32'h4236a4af, 32'hc259077f, 32'hc28ecc01, 32'hc2a3dacf, 32'h42226ed5, 32'h426a53e7, 32'h4288ae7b};
test_bias[3205:3205] = '{32'h422d1944};
test_output[3205:3205] = '{32'h452a199b};
test_input[25648:25655] = '{32'hc2c02e90, 32'h4289e436, 32'hc13066f2, 32'hc2802c59, 32'h421cad3f, 32'hc239b776, 32'h42757894, 32'hc2c6bfd6};
test_weights[25648:25655] = '{32'hc21b956f, 32'hc1ac7530, 32'hc1ef0dba, 32'h4296a86d, 32'hc1e71460, 32'hc1ba3be1, 32'h42061f99, 32'hc29807da};
test_bias[3206:3206] = '{32'h42599228};
test_output[3206:3206] = '{32'h45e64573};
test_input[25656:25663] = '{32'hc2b86b45, 32'h4279a2a7, 32'h42b05b2e, 32'h41a3d96a, 32'hc1d317cc, 32'h42b57be1, 32'h429c2e50, 32'hc227f02f};
test_weights[25656:25663] = '{32'h419bee4e, 32'h42a8b57d, 32'h421787c5, 32'h41904cd2, 32'h40e01777, 32'h42a762c4, 32'hc284cf2b, 32'hc2a81beb};
test_bias[3207:3207] = '{32'hc21d205b};
test_output[3207:3207] = '{32'h46496b5a};
test_input[25664:25671] = '{32'h40b07a7a, 32'h41d549ae, 32'h42a4f805, 32'hc2005d18, 32'h418a0290, 32'hc2795624, 32'h42469610, 32'hc26864cd};
test_weights[25664:25671] = '{32'hc23b543b, 32'h42b68dac, 32'hc25a3918, 32'hc28948ce, 32'hc2050b35, 32'h42325df5, 32'h429186eb, 32'hc1494175};
test_bias[3208:3208] = '{32'h4170f1de};
test_output[3208:3208] = '{32'h445cbdc2};
test_input[25672:25679] = '{32'h42922c83, 32'hc263a057, 32'h427be5b8, 32'h42755ead, 32'hc29e8d9c, 32'hc2ba8b81, 32'hc2b1dfc8, 32'hc0b40c69};
test_weights[25672:25679] = '{32'hc2a1e676, 32'hc23d8348, 32'hc19cc6c2, 32'hc2b4e020, 32'h42bf03ed, 32'hc089fbd3, 32'hc1d72c87, 32'hc19c68b0};
test_bias[3209:3209] = '{32'h414b6f26};
test_output[3209:3209] = '{32'hc665022c};
test_input[25680:25687] = '{32'h42a5c079, 32'hc237a23a, 32'h4251b047, 32'hc2bbc61e, 32'hc2b01aaf, 32'hc2c113b1, 32'h415e07a6, 32'hc29b6b7a};
test_weights[25680:25687] = '{32'h42270e27, 32'h420203e5, 32'h4027a488, 32'hc1ae5e95, 32'h4291d63a, 32'hc260dcb6, 32'hc287f3b7, 32'hc135ad95};
test_bias[3210:3210] = '{32'hc1c76c07};
test_output[3210:3210] = '{32'h45401372};
test_input[25688:25695] = '{32'h418077db, 32'hc1fd643e, 32'hc29e62af, 32'h42483c36, 32'hc24a9e22, 32'hc1b28ec1, 32'hc2bc5274, 32'h42405216};
test_weights[25688:25695] = '{32'h420f5a2e, 32'h42094a04, 32'hc1d980bd, 32'h415644e9, 32'hc0815bd3, 32'hc273c8cc, 32'hc2a8f935, 32'hc1d8106f};
test_bias[3211:3211] = '{32'h422eafed};
test_output[3211:3211] = '{32'h46254591};
test_input[25696:25703] = '{32'hc2c4cb6d, 32'hc19b5385, 32'hc2b1fba1, 32'hc2065997, 32'h42adb7b7, 32'hc0cc3c9a, 32'hc219c348, 32'h42c067ad};
test_weights[25696:25703] = '{32'h4275f73e, 32'h422d7a6a, 32'h4286c3cc, 32'h42b43c0b, 32'h4290f7ed, 32'hc11d2dcd, 32'hc29f13a0, 32'hc13fa06c};
test_bias[3212:3212] = '{32'hc2567ac4};
test_output[3212:3212] = '{32'hc5f0ccfa};
test_input[25704:25711] = '{32'h4260316d, 32'h41d6245e, 32'h42b73e77, 32'h42a04484, 32'h41b04583, 32'hc25bee0f, 32'h409d6d64, 32'h427979d3};
test_weights[25704:25711] = '{32'h42023814, 32'h425da4fc, 32'h3fad50ff, 32'hc235335d, 32'hc24f7110, 32'hc2b01d14, 32'hc1d5e20b, 32'hc18ae5b6};
test_bias[3213:3213] = '{32'h40d9daea};
test_output[3213:3213] = '{32'h450f52a5};
test_input[25712:25719] = '{32'hc22945a3, 32'h407d485d, 32'hc25919d2, 32'hc29f9fe2, 32'hbfbfff68, 32'h4120538a, 32'hc231df9c, 32'hc2c3bff6};
test_weights[25712:25719] = '{32'hc1ba2bf4, 32'hc28a019b, 32'h42845c38, 32'hc1bb6153, 32'h41f25245, 32'h427d1f24, 32'hc212d2ef, 32'h408957ff};
test_bias[3214:3214] = '{32'hc2339317};
test_output[3214:3214] = '{32'h443a4823};
test_input[25720:25727] = '{32'hc113090c, 32'hc0efef95, 32'h429f9721, 32'hc29a8d08, 32'hc12bec59, 32'hc2bcaf4e, 32'hc27a8532, 32'h42b61e2c};
test_weights[25720:25727] = '{32'hc2bf68c2, 32'hc1f97e4e, 32'hc1c3aa3c, 32'h42a5384d, 32'h42c5c147, 32'h41e04274, 32'h42bf7be5, 32'hc2693948};
test_bias[3215:3215] = '{32'hc25d4b58};
test_output[3215:3215] = '{32'hc6ae2420};
test_input[25728:25735] = '{32'hc26e08d0, 32'hc22de288, 32'h41c2a062, 32'h428edace, 32'hc24cf688, 32'h42addf9a, 32'hc01690b7, 32'hc2151dcd};
test_weights[25728:25735] = '{32'hc2a7fb3a, 32'h423d0b32, 32'h4278d22c, 32'h42999af7, 32'hc23a043c, 32'hc0b6f27b, 32'hc28407aa, 32'h4225f033};
test_bias[3216:3216] = '{32'h42923e12};
test_output[3216:3216] = '{32'h46243a8d};
test_input[25736:25743] = '{32'hc1ad0877, 32'hc297759c, 32'hc2c4c5e5, 32'h42672d8d, 32'hc2b9f3bc, 32'hc19b6393, 32'hc28caedd, 32'hc27c02a6};
test_weights[25736:25743] = '{32'hc1133e71, 32'h41f80722, 32'h4139b386, 32'h42bd03af, 32'h42a59434, 32'h40088f7b, 32'hc061947a, 32'hc2c317f5};
test_bias[3217:3217] = '{32'h421b80f8};
test_output[3217:3217] = '{32'h4458382e};
test_input[25744:25751] = '{32'hc24fa05d, 32'hc251ac9f, 32'h41f97283, 32'h429b238a, 32'hc1cac656, 32'hc251428c, 32'hc228c833, 32'h42c45f8a};
test_weights[25744:25751] = '{32'h42031a58, 32'hc2642df1, 32'hc2c5d593, 32'hc20b650a, 32'hc29f38c0, 32'h40f59f56, 32'h42a9c40c, 32'h4287f82a};
test_bias[3218:3218] = '{32'h40130457};
test_output[3218:3218] = '{32'h43558d45};
test_input[25752:25759] = '{32'hc0d84d8b, 32'h428d680d, 32'h4243ca25, 32'h427f7fd0, 32'hc0fefd76, 32'hc285225a, 32'h42c0eb1d, 32'h42712387};
test_weights[25752:25759] = '{32'hc289f5bd, 32'hc1ccd653, 32'hbf03e738, 32'hc1730740, 32'hc17f1043, 32'h407878c2, 32'h42a62220, 32'h4288c74a};
test_bias[3219:3219] = '{32'h4295be8e};
test_output[3219:3219] = '{32'h46182d57};
test_input[25760:25767] = '{32'hc26e2246, 32'hc28638e5, 32'h42c0f092, 32'h4227cf3b, 32'h41d90e15, 32'h41439cb6, 32'hc202e1d1, 32'h421b8a3e};
test_weights[25760:25767] = '{32'h4239c51c, 32'hc21642b4, 32'h427413c1, 32'hc2b1a300, 32'hc25506aa, 32'hc24df9d3, 32'h42c7d6e5, 32'h40ce2eb9};
test_bias[3220:3220] = '{32'hc1209354};
test_output[3220:3220] = '{32'hc5472e1a};
test_input[25768:25775] = '{32'h42780794, 32'h4202ac6c, 32'h42027802, 32'h415d4c05, 32'hc244aea7, 32'h4133a4cf, 32'hc0920272, 32'h421949b6};
test_weights[25768:25775] = '{32'hc18ab334, 32'h42c7a407, 32'hc273b096, 32'h4190939b, 32'h42b08530, 32'hc2a610fb, 32'h42951769, 32'h40e847b6};
test_bias[3221:3221] = '{32'hc25cb1d5};
test_output[3221:3221] = '{32'hc59a63b4};
test_input[25776:25783] = '{32'hc2b3f3a9, 32'hc2ae3fc6, 32'hc1dc49e7, 32'hc182f8c8, 32'hc1b0c6e9, 32'h41ac1e4a, 32'h4278e97e, 32'hc2a8ffb1};
test_weights[25776:25783] = '{32'hc1bc2008, 32'hc2336936, 32'hc21105a1, 32'h4205266e, 32'h429d1fd1, 32'h424e7616, 32'hc228186c, 32'hc12ea825};
test_bias[3222:3222] = '{32'hc2823a6d};
test_output[3222:3222] = '{32'h457fdb47};
test_input[25784:25791] = '{32'hc1b738c4, 32'h40968e1d, 32'h42524b6c, 32'h4246999d, 32'h42b3870e, 32'hc24864a7, 32'hc19756eb, 32'h41ac673d};
test_weights[25784:25791] = '{32'hc2a2cc4a, 32'hc1b2e43b, 32'hc23cb7b7, 32'h4232bef2, 32'hc2bb73fc, 32'h41c318af, 32'h4261f296, 32'hc11f4cae};
test_bias[3223:3223] = '{32'hc29ef944};
test_output[3223:3223] = '{32'hc614712a};
test_input[25792:25799] = '{32'h42b56623, 32'h412e0827, 32'hc20712a6, 32'hc2925e1a, 32'hc1fc188b, 32'hc0dd176c, 32'h429ee211, 32'h423fe997};
test_weights[25792:25799] = '{32'h41e61431, 32'hc1f1a9f9, 32'hc1f346c9, 32'h428989fc, 32'h42771bad, 32'hc239ad73, 32'h405e234b, 32'h41c9f831};
test_bias[3224:3224] = '{32'h4219bbd9};
test_output[3224:3224] = '{32'hc4e4524f};
test_input[25800:25807] = '{32'h42b37e36, 32'hc2300c94, 32'hc2a34a9e, 32'hc27a5239, 32'hc28a268c, 32'hc146a737, 32'hc2a5f715, 32'h41850c4f};
test_weights[25800:25807] = '{32'h42c5a3cf, 32'hc236e5fe, 32'hc259da4d, 32'hc2c7f994, 32'h42b6d7f5, 32'hc2a6cae9, 32'h42bf910a, 32'h42bc3dfd};
test_bias[3225:3225] = '{32'h42135e3c};
test_output[3225:3225] = '{32'h461b9d93};
test_input[25808:25815] = '{32'hc0837b27, 32'h42935394, 32'h42adad9c, 32'hc26822d3, 32'hc20cfeb4, 32'h4202fc47, 32'hc2555654, 32'hc2323090};
test_weights[25808:25815] = '{32'h4292e7e0, 32'hc28e0969, 32'h422825d7, 32'hc23d7a6a, 32'hc1519e55, 32'hc21f9623, 32'h42b4f340, 32'hbef9f351};
test_bias[3226:3226] = '{32'h40ee8331};
test_output[3226:3226] = '{32'hc595352d};
test_input[25816:25823] = '{32'hc26e9c7f, 32'hc244f21a, 32'hc2bbbe58, 32'h420eb3f1, 32'hc1aaab33, 32'hc2c1cfb1, 32'h4017eab0, 32'h42230f43};
test_weights[25816:25823] = '{32'hc27067ae, 32'h41e0af96, 32'hc2a631d9, 32'h428cb594, 32'h42b45415, 32'hc28cebfd, 32'hc1dec90a, 32'h41cd167e};
test_bias[3227:3227] = '{32'hc2929634};
test_output[3227:3227] = '{32'h468f2601};
test_input[25824:25831] = '{32'h42c35148, 32'h420a3aa7, 32'h410674ad, 32'hc05a03ac, 32'h42659bc8, 32'h42a3d6ae, 32'h42c6c6c0, 32'hc24beb3a};
test_weights[25824:25831] = '{32'hc08acf87, 32'h429eb16b, 32'hc212019d, 32'hc186dcc8, 32'h423a6666, 32'h41b32f74, 32'h4259bba2, 32'hc2a840ea};
test_bias[3228:3228] = '{32'h3fb5221c};
test_output[3228:3228] = '{32'h467e5c23};
test_input[25832:25839] = '{32'hc2587e76, 32'h4263c084, 32'h42962a2f, 32'hc09d3e9b, 32'hc2570a58, 32'hc2bc70c2, 32'hc2162da3, 32'h42b3418d};
test_weights[25832:25839] = '{32'h41c4cc6a, 32'h424d642f, 32'hc207eead, 32'hc10f4086, 32'h42acf896, 32'hc230233d, 32'hc27282de, 32'h41b9970e};
test_bias[3229:3229] = '{32'h42a7fa19};
test_output[3229:3229] = '{32'h453cfa24};
test_input[25840:25847] = '{32'h42906d4a, 32'hc25e55bf, 32'h42019ef0, 32'hc1c2f320, 32'hc29f3a98, 32'hc28e5b06, 32'h42aaf358, 32'hc21bf172};
test_weights[25840:25847] = '{32'hc2a24ddd, 32'h419a32d6, 32'h429b8bf6, 32'h42051f9c, 32'hc161df29, 32'hc2a02527, 32'hc13fa85f, 32'hc249b831};
test_bias[3230:3230] = '{32'h42c6df8c};
test_output[3230:3230] = '{32'h45252867};
test_input[25848:25855] = '{32'hc289ffbe, 32'hc2921781, 32'hc1e5a58e, 32'h42401286, 32'hc248cdad, 32'h42808dd7, 32'h428767ab, 32'hc26645a0};
test_weights[25848:25855] = '{32'hc2738afb, 32'hc19dea5c, 32'hc12d3db2, 32'h4296dbfe, 32'h42657047, 32'hc2803517, 32'hc23fd198, 32'h42640215};
test_bias[3231:3231] = '{32'h424bc03b};
test_output[3231:3231] = '{32'hc573d550};
test_input[25856:25863] = '{32'hc2b252f4, 32'hc293b5ce, 32'h42a227f5, 32'hc2b1ca8b, 32'h4232172a, 32'hc0fcdaa0, 32'h42c0e544, 32'hc2b0db69};
test_weights[25856:25863] = '{32'h42c7d60f, 32'h425963d6, 32'h42835e9f, 32'hc1dc0899, 32'hc2b6819d, 32'h41a1467b, 32'h40b18197, 32'hc220bec0};
test_bias[3232:3232] = '{32'h41ad68a1};
test_output[3232:3232] = '{32'hc5a47fc3};
test_input[25864:25871] = '{32'h426f6159, 32'hc2916d07, 32'hc2ae70c5, 32'hc20ea2de, 32'hc27dc7a8, 32'h421c040a, 32'hc28f24ed, 32'h4291a222};
test_weights[25864:25871] = '{32'hc0caa018, 32'h40769ee2, 32'h426d4412, 32'hc2426a3c, 32'h41c38a7d, 32'hc2478f22, 32'h425a5515, 32'hc262812e};
test_bias[3233:3233] = '{32'h420e35f6};
test_output[3233:3233] = '{32'hc6739a89};
test_input[25872:25879] = '{32'hc0f0fc65, 32'h41078e25, 32'hc0105bda, 32'hc24e8ff3, 32'hc27314b2, 32'hc265a91e, 32'hc1538c84, 32'h42b93c38};
test_weights[25872:25879] = '{32'hc2bb3611, 32'h42a2de33, 32'h42860e99, 32'h42c002d2, 32'h42c7d8c7, 32'hc2a5fa46, 32'hc2a5d930, 32'hc166831e};
test_bias[3234:3234] = '{32'h42107fb9};
test_output[3234:3234] = '{32'hc5a33bd5};
test_input[25880:25887] = '{32'h4214b9fe, 32'h410445db, 32'hbf6cb861, 32'h42b369dc, 32'h42af9fa7, 32'h42779863, 32'hc2324c68, 32'hc26cd6b8};
test_weights[25880:25887] = '{32'hc1b006c9, 32'h42a744e1, 32'h428030e8, 32'h40a00577, 32'hc003a10f, 32'hc29169c3, 32'hc14f2240, 32'hc21abbf1};
test_bias[3235:3235] = '{32'h427ca9b2};
test_output[3235:3235] = '{32'hc4b9f8be};
test_input[25888:25895] = '{32'h42a694c2, 32'hc203ed26, 32'h42b80176, 32'hc200efb7, 32'hc00c80e8, 32'h414ae625, 32'h41534935, 32'h41f3d1ce};
test_weights[25888:25895] = '{32'h40cd28c7, 32'h41fe4dc7, 32'h41db08c5, 32'h42a51702, 32'h41b3046e, 32'hc2b863fa, 32'h42c30229, 32'hc28b428c};
test_bias[3236:3236] = '{32'hbfa49862};
test_output[3236:3236] = '{32'hc5296559};
test_input[25896:25903] = '{32'h4221b7f4, 32'h42996ea4, 32'h41e61326, 32'h4281a77e, 32'hc23b2eda, 32'hc0832752, 32'h42c5a6ed, 32'h400bb991};
test_weights[25896:25903] = '{32'hc0a05510, 32'h42a40479, 32'hc286f064, 32'h41304220, 32'h4257fbab, 32'h426aeb48, 32'h41b48ff1, 32'hc1954460};
test_bias[3237:3237] = '{32'hc2c68451};
test_output[3237:3237] = '{32'h4582cd2b};
test_input[25904:25911] = '{32'h414110fe, 32'hc18763aa, 32'h42c345e9, 32'h41250f7f, 32'h40125dad, 32'h4258fbbc, 32'h410ce393, 32'hc2131866};
test_weights[25904:25911] = '{32'hc2605ba3, 32'hc24e2dc3, 32'hc2911f36, 32'h42a66998, 32'hc29738be, 32'h42385fe3, 32'h429b3f95, 32'h42238681};
test_bias[3238:3238] = '{32'h429774df};
test_output[3238:3238] = '{32'hc58afad0};
test_input[25912:25919] = '{32'h419f4204, 32'h42574d9e, 32'h42c6abb1, 32'h415432ec, 32'h4252ebcf, 32'hc24f7361, 32'h42a6177f, 32'h42a0bf62};
test_weights[25912:25919] = '{32'hc2922d7b, 32'hc1c17a3c, 32'hbcbd7da1, 32'h42a09734, 32'hc1dfa655, 32'hc2c63d0a, 32'hc243afeb, 32'hc29c803b};
test_bias[3239:3239] = '{32'hc2108ac6};
test_output[3239:3239] = '{32'hc6037f7b};
test_input[25920:25927] = '{32'hc2658e63, 32'h42ad9032, 32'h42a6db72, 32'hc2ba2c36, 32'h420ea98d, 32'hc2713c6b, 32'hc1f20d73, 32'h427c158e};
test_weights[25920:25927] = '{32'h42969874, 32'hc259be3c, 32'h428ebe6f, 32'h423f96f3, 32'h421d41e5, 32'hc2951282, 32'h42b6d45a, 32'h42b0a611};
test_bias[3240:3240] = '{32'h42917e8a};
test_output[3240:3240] = '{32'h4498a2ce};
test_input[25928:25935] = '{32'h428f0aec, 32'hc2adfd39, 32'hc2b2e517, 32'hc1f932bf, 32'h41074cb9, 32'h427aadf4, 32'h422f7e59, 32'hc26a9199};
test_weights[25928:25935] = '{32'h41d317df, 32'hc292fe13, 32'h42215df9, 32'hc200e8f7, 32'h413ef427, 32'hc290b0d0, 32'h42b65955, 32'hc2b12d07};
test_bias[3241:3241] = '{32'h42480ee4};
test_output[3241:3241] = '{32'h4623e253};
test_input[25936:25943] = '{32'h421aee68, 32'hc2c3d47a, 32'h42b8a428, 32'h40475a8b, 32'hc2a2e224, 32'hc13d56f0, 32'h427ad807, 32'h3fbe485b};
test_weights[25936:25943] = '{32'hc1212123, 32'hc1f551b2, 32'hc2a8189d, 32'hc29f429d, 32'hc289d78d, 32'h429f1194, 32'hc26a13c2, 32'h429c75fc};
test_bias[3242:3242] = '{32'hc2440e2d};
test_output[3242:3242] = '{32'hc5872cad};
test_input[25944:25951] = '{32'h42494570, 32'h4249b094, 32'hc0f556de, 32'hc1d77365, 32'hbfd9221f, 32'h42c39c89, 32'h3f766024, 32'hc1b18a37};
test_weights[25944:25951] = '{32'hc2712a9d, 32'h421a19f2, 32'h42c6289f, 32'hc17d6e1b, 32'h42a64435, 32'h41669dad, 32'h4268792b, 32'h429a7c3a};
test_bias[3243:3243] = '{32'hc23e55fd};
test_output[3243:3243] = '{32'hc4e8ad18};
test_input[25952:25959] = '{32'h4271e560, 32'hc2b04d0c, 32'h420ec18f, 32'hc29d60ff, 32'h42c16e60, 32'hc2862c94, 32'h42a0c749, 32'h42bb7672};
test_weights[25952:25959] = '{32'h42397c0f, 32'hc14e88e0, 32'hc291b3a8, 32'hc22cbacb, 32'h41ab2d9e, 32'h429461de, 32'hc2644749, 32'hc2abea52};
test_bias[3244:3244] = '{32'hc26c5539};
test_output[3244:3244] = '{32'hc629ddd0};
test_input[25960:25967] = '{32'hc01c2cb9, 32'h42a06d38, 32'hc27c0c16, 32'hc22d155e, 32'h42a53ef2, 32'h428f2566, 32'h428bc04c, 32'hc28e81f3};
test_weights[25960:25967] = '{32'hc29ea659, 32'h4291921d, 32'hc2c7bf4d, 32'h40299bb3, 32'h4059166e, 32'h40dbffe6, 32'hc0fb40eb, 32'h40c674ac};
test_bias[3245:3245] = '{32'h41bbac60};
test_output[3245:3245] = '{32'h463bbeda};
test_input[25968:25975] = '{32'hc29c6010, 32'h42136e3b, 32'hc218ba96, 32'hc2693aa8, 32'hc27e6710, 32'h4268add4, 32'h426a8846, 32'h41cbaa38};
test_weights[25968:25975] = '{32'h423f7ac7, 32'h4198facf, 32'h42123ad5, 32'hc21bd740, 32'hc220a322, 32'hc1207c32, 32'hc14ede01, 32'hc1e2e906};
test_bias[3246:3246] = '{32'h41bd53c5};
test_output[3246:3246] = '{32'hc4ce0051};
test_input[25976:25983] = '{32'hc235359d, 32'hc238ef1c, 32'hc2a13cc4, 32'h424d331d, 32'h42306c65, 32'h427d308c, 32'h42b24779, 32'hc21f3bd8};
test_weights[25976:25983] = '{32'h427115b8, 32'hc11aa11e, 32'h410f2536, 32'h41abdd22, 32'h41c849a3, 32'h42bbd442, 32'h41eaedcd, 32'hc1b493a4};
test_bias[3247:3247] = '{32'h414f7525};
test_output[3247:3247] = '{32'h46078cc4};
test_input[25984:25991] = '{32'h42c25a14, 32'h41e51ebf, 32'h41dcdb54, 32'hc2be9c75, 32'h41b4d81b, 32'h4116d4a5, 32'h42c0d130, 32'h4289788d};
test_weights[25984:25991] = '{32'hc2bd2ca1, 32'h42a64acd, 32'hc23bf65f, 32'hc26b5ad7, 32'hc22befdb, 32'h4230531b, 32'h42a2eca1, 32'h41ac7da2};
test_bias[3248:3248] = '{32'h429f5ffa};
test_output[3248:3248] = '{32'h45c6ba9f};
test_input[25992:25999] = '{32'h41dd6592, 32'h428a5d3d, 32'hc25d9f34, 32'h429c4856, 32'hc28bc53b, 32'h3fa5d23d, 32'hc1d62ad6, 32'h41c139e7};
test_weights[25992:25999] = '{32'h42785050, 32'h42595f85, 32'h423235e1, 32'h4114bd32, 32'hc1b8b296, 32'hc1cebe6b, 32'h429f55e1, 32'hc2a2d550};
test_bias[3249:3249] = '{32'h4215c9e9};
test_output[3249:3249] = '{32'h449cb675};
test_input[26000:26007] = '{32'h42c3984e, 32'hc16e87f3, 32'hc281702c, 32'h42310cc8, 32'h4288b018, 32'h419902ca, 32'h4204623f, 32'hc1808b33};
test_weights[26000:26007] = '{32'hc2c07ea7, 32'hc1e3949a, 32'h41a76e26, 32'h42b43b33, 32'hc10c7011, 32'h425e1ef9, 32'hc2bbff59, 32'hc18dcc98};
test_bias[3250:3250] = '{32'h42c1d5c3};
test_output[3250:3250] = '{32'hc606b5c4};
test_input[26008:26015] = '{32'h41974761, 32'h42c5140b, 32'h429be4a8, 32'h42486592, 32'h42acc175, 32'hc2812d69, 32'hc1a73de7, 32'hc1268a2d};
test_weights[26008:26015] = '{32'h422b1d05, 32'h422cd838, 32'hc28e1ebb, 32'h42170bec, 32'h426843fd, 32'h42ac528c, 32'h42c56250, 32'hc28bf2ce};
test_bias[3251:3251] = '{32'h4242b397};
test_output[3251:3251] = '{32'hc3cfd831};
test_input[26016:26023] = '{32'hc14edf68, 32'h42196ee5, 32'h413fc6d5, 32'hc1f05714, 32'h4285cd72, 32'h4197bd5e, 32'hc21a9f51, 32'hc2717a3a};
test_weights[26016:26023] = '{32'hc1bb496d, 32'hc128b7dd, 32'h425ce2e1, 32'hc29b9ff0, 32'hc2af5a83, 32'hc237334a, 32'hc29293b2, 32'hc28c76a4};
test_bias[3252:3252] = '{32'h423293cb};
test_output[3252:3252] = '{32'h454d0dfa};
test_input[26024:26031] = '{32'hc19ae31a, 32'hc1bcce37, 32'h40562cae, 32'h41358e0f, 32'hc23511f3, 32'hc203ffb4, 32'h416a83b3, 32'hc0a178bd};
test_weights[26024:26031] = '{32'h428512ff, 32'h408e90fd, 32'h405f3a61, 32'h4287ea23, 32'h418d18f2, 32'h41ec130d, 32'h428d33ac, 32'hc21f7366};
test_bias[3253:3253] = '{32'hc2a9037d};
test_output[3253:3253] = '{32'hc499e9e1};
test_input[26032:26039] = '{32'h421c4755, 32'hc2ac99aa, 32'hc20d4809, 32'h41b32d4f, 32'hc23a44aa, 32'h41f3b86a, 32'hc264be17, 32'hc29fd324};
test_weights[26032:26039] = '{32'h42b8d903, 32'h428c7d3f, 32'h40c48439, 32'h429c4a88, 32'hc2a76185, 32'h42088bbf, 32'hc17cb96e, 32'h416c318f};
test_bias[3254:3254] = '{32'h429d93ad};
test_output[3254:3254] = '{32'h456edbdc};
test_input[26040:26047] = '{32'hc237be48, 32'hc2025f08, 32'h421e2750, 32'h42275473, 32'hc25d3a93, 32'hc1f66129, 32'h419bd8a9, 32'h429cb97d};
test_weights[26040:26047] = '{32'h42238797, 32'hc20c0818, 32'hc160379f, 32'h418e78fb, 32'h41aa0fe8, 32'hc28e0259, 32'hc15a7681, 32'hc276241e};
test_bias[3255:3255] = '{32'hc2c7d0ee};
test_output[3255:3255] = '{32'hc593976d};
test_input[26048:26055] = '{32'hc29c8cb1, 32'hc2735aa6, 32'h4217832c, 32'hc2ba48e9, 32'hc215b46a, 32'hc0db5fb8, 32'h417351a8, 32'h42995261};
test_weights[26048:26055] = '{32'h40ced1e3, 32'hc1b71304, 32'h3fc83cb9, 32'hc27369c3, 32'h4213fd74, 32'hc0f2ce6e, 32'hc126c83c, 32'h42c741f5};
test_bias[3256:3256] = '{32'hc1e42529};
test_output[3256:3256] = '{32'h4646ee3d};
test_input[26056:26063] = '{32'hc2a062eb, 32'hc2b7cdda, 32'h41be460c, 32'h42a70dcc, 32'hc2689561, 32'hc1a0faa4, 32'h41e605ea, 32'h4280efb7};
test_weights[26056:26063] = '{32'hc132ea71, 32'hc27bd707, 32'h42bb5f9c, 32'h41f380ba, 32'h3fea0315, 32'hc169559e, 32'hc28afd1d, 32'h41d89508};
test_bias[3257:3257] = '{32'hc1aeccc8};
test_output[3257:3257] = '{32'h46319806};
test_input[26064:26071] = '{32'hc2bc557e, 32'h41c850e2, 32'hc296e61c, 32'h40a8f90f, 32'hc1fe7ad6, 32'hc2a318ec, 32'hc0ca090d, 32'h4202c6a8};
test_weights[26064:26071] = '{32'h42815bda, 32'hc0e2e7c3, 32'hc26cf20a, 32'hc18767b1, 32'h42b3b093, 32'hc2a94f63, 32'hc2922cf6, 32'hc2a2a220};
test_bias[3258:3258] = '{32'h429ecf57};
test_output[3258:3258] = '{32'h421e5f25};
test_input[26072:26079] = '{32'hc29cb755, 32'h41ca0fb7, 32'h42605906, 32'hc211b793, 32'hc2a5aaf4, 32'h41eaa8b3, 32'h42c65da8, 32'hc25db520};
test_weights[26072:26079] = '{32'hc2c1c682, 32'hc1851c8f, 32'hc29d0720, 32'h42a0236e, 32'hc2b43306, 32'h426df866, 32'hc2714073, 32'hc28524b5};
test_bias[3259:3259] = '{32'hc239bf29};
test_output[3259:3259] = '{32'h45d207d6};
test_input[26080:26087] = '{32'h42640776, 32'h4269cb09, 32'hbf828973, 32'h3fdac1f1, 32'h41411653, 32'h4267f74c, 32'h414b7223, 32'h41dd9055};
test_weights[26080:26087] = '{32'hc293e8e0, 32'h4274ef2e, 32'hc102bbfd, 32'h421d05be, 32'h41b19e54, 32'h4282ce61, 32'h41edbe4f, 32'hc293a15d};
test_bias[3260:3260] = '{32'hc194d75d};
test_output[3260:3260] = '{32'h44e2c465};
test_input[26088:26095] = '{32'h42816bc9, 32'h42ac1bdc, 32'hc29a02d5, 32'hc244e6e4, 32'h429ef749, 32'h4243e5ad, 32'h41b97e4c, 32'h42094e48};
test_weights[26088:26095] = '{32'hc2171e51, 32'hc261dac0, 32'h42aad997, 32'h429758f8, 32'h4297b519, 32'h420748ca, 32'hc19eeda1, 32'hc1d63415};
test_bias[3261:3261] = '{32'hc196bd36};
test_output[3261:3261] = '{32'hc630e05a};
test_input[26096:26103] = '{32'h409a5a1e, 32'h425637b6, 32'h41d3d5de, 32'h42b3a0ba, 32'hc2a8c14a, 32'hc294b88d, 32'hc2810407, 32'h425b71de};
test_weights[26096:26103] = '{32'hc2bf6a69, 32'h410b7c35, 32'h41c76ff2, 32'h4284ffdf, 32'h42ae25e5, 32'h419e78e7, 32'h40d7ff01, 32'h42ad0070};
test_bias[3262:3262] = '{32'h42add21c};
test_output[3262:3262] = '{32'h450a6e3c};
test_input[26104:26111] = '{32'hbe6400fb, 32'hc2ad84dc, 32'hc2a14fb1, 32'h42b09829, 32'hc1651300, 32'h420be56d, 32'hc2a55e0b, 32'hc26aeeb9};
test_weights[26104:26111] = '{32'h422c620e, 32'hc220afeb, 32'h42c7df0d, 32'h424db61e, 32'hc2af3c67, 32'h4284bc54, 32'h423ba048, 32'h4296b21e};
test_bias[3263:3263] = '{32'h426e5ac2};
test_output[3263:3263] = '{32'hc5934326};
test_input[26112:26119] = '{32'h4212ad35, 32'h409b745f, 32'hc2a0d5c2, 32'hc2bc4b43, 32'h41e02962, 32'hc2bc7f93, 32'hc2b87d95, 32'hc1e69796};
test_weights[26112:26119] = '{32'h421fd766, 32'h420b105c, 32'hc2c38a5d, 32'h42bb6c42, 32'h424342b9, 32'h41ea6cfb, 32'hc237bbce, 32'h4230dd97};
test_bias[3264:3264] = '{32'h4169c973};
test_output[3264:3264] = '{32'h450d1415};
test_input[26120:26127] = '{32'hc2664fb7, 32'hc2a2764b, 32'hc0961e89, 32'h42b4d8d0, 32'h423bc006, 32'h4284d507, 32'h4291b4fd, 32'h41bba89d};
test_weights[26120:26127] = '{32'hc24156fa, 32'h4249278f, 32'hc26dde16, 32'h429d1a3f, 32'hc29b04b2, 32'hc0f55bdd, 32'hc2669733, 32'h4233d9f2};
test_bias[3265:3265] = '{32'hc27a75ad};
test_output[3265:3265] = '{32'hc49f6652};
test_input[26128:26135] = '{32'h4289f667, 32'hc28057dc, 32'hc2c305c4, 32'hc1f379eb, 32'h4237ac57, 32'h4270ebcb, 32'h42734b2e, 32'hc2af7980};
test_weights[26128:26135] = '{32'hc205bd17, 32'h426f7402, 32'h419c73d4, 32'hc2574e9d, 32'hc2506bbe, 32'hc20fb9eb, 32'hc28cac2c, 32'hc25e211f};
test_bias[3266:3266] = '{32'hc14fe47d};
test_output[3266:3266] = '{32'hc6226108};
test_input[26136:26143] = '{32'h42c6f803, 32'h42a86645, 32'hc2bdd5b8, 32'hc26e40f4, 32'h41dffd41, 32'h41e82686, 32'hc28b1d0e, 32'h42a3432c};
test_weights[26136:26143] = '{32'h4262a43b, 32'hc1ed8fe9, 32'h422b0d5c, 32'h42113a2f, 32'hc11686ee, 32'hc28bc745, 32'hc2a023c8, 32'h42b8fa5f};
test_bias[3267:3267] = '{32'hc22a860d};
test_output[3267:3267] = '{32'h45f0a1c4};
test_input[26144:26151] = '{32'h4231ad65, 32'h419eda88, 32'h40d83570, 32'hc2a2a8f6, 32'h41b9f5fe, 32'h4126bf93, 32'h40ee13dc, 32'h42123acc};
test_weights[26144:26151] = '{32'hc29def73, 32'hc120a4d8, 32'hc1092c24, 32'h4285664c, 32'h4234b731, 32'hc1e172f1, 32'h40f4acf8, 32'h41b76548};
test_bias[3268:3268] = '{32'hc2ad1c95};
test_output[3268:3268] = '{32'hc5ee4660};
test_input[26152:26159] = '{32'hc2a7ced7, 32'hc29489f0, 32'h42c56ba0, 32'h42ba0a25, 32'hc2116b6b, 32'h42ba0dd9, 32'hc29d53f9, 32'hc0b65922};
test_weights[26152:26159] = '{32'h42c1d199, 32'hc233b264, 32'h429b4458, 32'hc1e949cf, 32'hc2262933, 32'h418ca4df, 32'hc2922e60, 32'h42105c0b};
test_bias[3269:3269] = '{32'h42bd4c6e};
test_output[3269:3269] = '{32'h460bb149};
test_input[26160:26167] = '{32'h4209e267, 32'h42aa1d1b, 32'hc176ae60, 32'hc2bccda8, 32'h42aa5318, 32'hc299b838, 32'hc0ecfa6e, 32'h41c9d60f};
test_weights[26160:26167] = '{32'h424def61, 32'h42486f7b, 32'h42058583, 32'hc0fcc5b0, 32'hc18daf94, 32'h42845452, 32'hc1a52a15, 32'hc20274f0};
test_bias[3270:3270] = '{32'hc2a71341};
test_output[3270:3270] = '{32'hc486ea76};
test_input[26168:26175] = '{32'h41461138, 32'hc2b5dfbf, 32'h42c72c20, 32'h40ab3040, 32'h41c0a743, 32'h412196aa, 32'hc28bf3d6, 32'hc2acc339};
test_weights[26168:26175] = '{32'h4214de2a, 32'h4253981f, 32'hc1a53053, 32'hc12a2a80, 32'h421d79f3, 32'h42994148, 32'h41a28141, 32'hc20b2df3};
test_bias[3271:3271] = '{32'h42a822c0};
test_output[3271:3271] = '{32'hc5400b70};
test_input[26176:26183] = '{32'h42883782, 32'h4268de38, 32'hc2227101, 32'h40434c0c, 32'hc260a14c, 32'h423b5ad8, 32'h421636b7, 32'h42320d65};
test_weights[26176:26183] = '{32'h429132ff, 32'hc2a574ef, 32'h42b4d907, 32'h429d91a1, 32'h4215269d, 32'hc28aa0b7, 32'h4217e538, 32'hc2918f06};
test_bias[3272:3272] = '{32'h42b8be5c};
test_output[3272:3272] = '{32'hc621f43e};
test_input[26184:26191] = '{32'hc21efaa6, 32'h423531cf, 32'h420484e3, 32'hc28c1712, 32'hc26ee527, 32'h42462ad8, 32'hc29704bb, 32'hc2c62ce1};
test_weights[26184:26191] = '{32'h4241c3a2, 32'hc223cfd4, 32'h4245a82a, 32'h4177e700, 32'hc19ba8a3, 32'h42a02b0d, 32'h427329a4, 32'hc2c0f90c};
test_bias[3273:3273] = '{32'h429a6d41};
test_output[3273:3273] = '{32'h45d9248b};
test_input[26192:26199] = '{32'h42c3a0e5, 32'hc1161c50, 32'h42ab3c16, 32'h429b643f, 32'h426073c8, 32'h42259966, 32'h423a07bf, 32'h42343871};
test_weights[26192:26199] = '{32'h421af36d, 32'hc22a5471, 32'hbd826670, 32'h41baf0cf, 32'hc1c9a7ce, 32'hc28b8593, 32'hc263c5a8, 32'hc2b629c7};
test_bias[3274:3274] = '{32'hbf03bbbf};
test_output[3274:3274] = '{32'hc59e025f};
test_input[26200:26207] = '{32'h41c1e2a5, 32'hc1c03868, 32'h4294bd89, 32'h419b1fb4, 32'hc1ef0b6b, 32'hc2b23980, 32'hc2b7d718, 32'hc0857bda};
test_weights[26200:26207] = '{32'hc24e8f59, 32'h42563897, 32'h426c3af6, 32'h42b6cec8, 32'h42289aad, 32'hc029826e, 32'h41c74da8, 32'h424cf599};
test_bias[3275:3275] = '{32'hc1c4acf4};
test_output[3275:3275] = '{32'h4294b795};
test_input[26208:26215] = '{32'hc26802ef, 32'hc14a5f97, 32'hc1a5df18, 32'h426214aa, 32'h427dc4eb, 32'hc1eed1f8, 32'h422ac42f, 32'hc27ef25f};
test_weights[26208:26215] = '{32'h4297854f, 32'hc2119da1, 32'hc2c3355a, 32'h428e8f9d, 32'h4279ad04, 32'hc2c49bb3, 32'h3c7f4a29, 32'h423316ec};
test_bias[3276:3276] = '{32'hc1fe6d74};
test_output[3276:3276] = '{32'h45bf83dc};
test_input[26216:26223] = '{32'hc2578196, 32'h4193ebab, 32'hc152f68a, 32'hc15687ea, 32'hc1870ffb, 32'h42581ea0, 32'hc28a7968, 32'h4241476e};
test_weights[26216:26223] = '{32'h412ac472, 32'h4144db16, 32'hc23b2d42, 32'h42ad3e1a, 32'h42878133, 32'h41c92731, 32'hbfa8b354, 32'h421d4178};
test_bias[3277:3277] = '{32'h4256ace2};
test_output[3277:3277] = '{32'h44aae8c1};
test_input[26224:26231] = '{32'h428b99af, 32'h42a88fa2, 32'hc1a51228, 32'hc194ba04, 32'h41d20f8c, 32'hc279489f, 32'h404a47ea, 32'hc29a1e36};
test_weights[26224:26231] = '{32'hc2a50ef8, 32'h42170b6a, 32'h424df171, 32'hc248a80d, 32'h40c94ab5, 32'hc1001d37, 32'hc0ec43c6, 32'hc2623737};
test_bias[3278:3278] = '{32'hc24d5422};
test_output[3278:3278] = '{32'h450bfb81};
test_input[26232:26239] = '{32'h42a6bcc4, 32'hc23bf0ed, 32'hc0478e3e, 32'hc2240b93, 32'hc2c065d8, 32'hc2c0b8d4, 32'h41d8c6bd, 32'hc253a2fe};
test_weights[26232:26239] = '{32'h423ac852, 32'hc2458657, 32'h427dc671, 32'hc22a5ff4, 32'h428e5fae, 32'hc25c9092, 32'h4183e903, 32'h42c11a83};
test_bias[3279:3279] = '{32'h401cadf3};
test_output[3279:3279] = '{32'h44c408bc};
test_input[26240:26247] = '{32'h40acf10e, 32'hc0674714, 32'h42176297, 32'h42c53b9d, 32'hc2a1c0c8, 32'h42585180, 32'h425caee9, 32'h41492c5d};
test_weights[26240:26247] = '{32'h41ee59a0, 32'h40ab8ef7, 32'h42902764, 32'h4198147b, 32'hc2250f1e, 32'hc2730e0b, 32'hc19fb583, 32'h42913314};
test_bias[3280:3280] = '{32'h420c3a6d};
test_output[3280:3280] = '{32'h45910f6e};
test_input[26248:26255] = '{32'h42201769, 32'h4277218e, 32'h424b6478, 32'h42825607, 32'h4182f716, 32'hc03a5b92, 32'h4225c4f2, 32'hc183d931};
test_weights[26248:26255] = '{32'h42949500, 32'h428a9615, 32'hc25ace43, 32'h4192bc26, 32'h42b192e8, 32'h408991a5, 32'hc2b46779, 32'h4191cb7a};
test_bias[3281:3281] = '{32'h41df89a7};
test_output[3281:3281] = '{32'h4541aae6};
test_input[26256:26263] = '{32'hc2536a25, 32'hc2a1de6c, 32'h406728da, 32'hc2a842f2, 32'hc22f3a42, 32'hc19f873f, 32'h428efe83, 32'h42808458};
test_weights[26256:26263] = '{32'h421b6bd2, 32'hc12c3a06, 32'hc281125b, 32'h42a285de, 32'h4118a544, 32'h42860496, 32'hc202d354, 32'hc200ca73};
test_bias[3282:3282] = '{32'hc257e562};
test_output[3282:3282] = '{32'hc6620ea1};
test_input[26264:26271] = '{32'hc2c10acb, 32'hc2c6a320, 32'h41cfb251, 32'hc23cb4ea, 32'h40b1a721, 32'hc2aa52de, 32'hc24c14a8, 32'h41ce0127};
test_weights[26264:26271] = '{32'h4237951d, 32'h419c13ab, 32'h42890c1b, 32'hc1a0de76, 32'h424b26dd, 32'hc2a188ec, 32'h425d9c4d, 32'h42558748};
test_bias[3283:3283] = '{32'hc268af8b};
test_output[3283:3283] = '{32'h44fb4563};
test_input[26272:26279] = '{32'hc21f9a46, 32'h429a2634, 32'h420b123c, 32'hc2a8e254, 32'h41c9ba17, 32'hc2205e5c, 32'h42b9e0db, 32'h4218f087};
test_weights[26272:26279] = '{32'h3f0f0fd4, 32'h42996986, 32'h421d915d, 32'h42c78935, 32'h428f2b0d, 32'hc26dae0c, 32'h4190507b, 32'h4078742e};
test_bias[3284:3284] = '{32'h42bd1117};
test_output[3284:3284] = '{32'h459a6cd8};
test_input[26280:26287] = '{32'hc1cd478d, 32'h4214b3f7, 32'hbff94901, 32'hc24198c6, 32'h42961931, 32'h40b4ceae, 32'hc1c18bc0, 32'hc2299920};
test_weights[26280:26287] = '{32'h420b454f, 32'h42b3c6e9, 32'h42361df9, 32'h423c7737, 32'h41c06b35, 32'h42c74dd6, 32'hc2a69335, 32'hc29ead6b};
test_bias[3285:3285] = '{32'hc1c07293};
test_output[3285:3285] = '{32'h45f3d1b8};
test_input[26288:26295] = '{32'hc2296c78, 32'hc2b95d3a, 32'h42a9e558, 32'hc19282cc, 32'h42ba2201, 32'hc2a4a8a9, 32'hc2878fd0, 32'h4230cf71};
test_weights[26288:26295] = '{32'h412ffb86, 32'hc29a9ce8, 32'h41ab5e0d, 32'h4218848f, 32'h429135c2, 32'hc24db58c, 32'h413b77db, 32'h40bf6480};
test_bias[3286:3286] = '{32'h428c7ce0};
test_output[3286:3286] = '{32'h468f5fde};
test_input[26296:26303] = '{32'h428b6f8e, 32'hc1ef115a, 32'h423532c6, 32'hc2922b88, 32'hbef6a517, 32'hc2c43cd3, 32'hc28f5df1, 32'hc273d477};
test_weights[26296:26303] = '{32'h42a1fcdc, 32'hc29ffc3b, 32'hc2ab995c, 32'hc29c655c, 32'hc2b0985e, 32'h41a96735, 32'hc0b7ce01, 32'h427491d4};
test_bias[3287:3287] = '{32'h4196ae6d};
test_output[3287:3287] = '{32'h458daf58};
test_input[26304:26311] = '{32'hc1122cb6, 32'h425a922a, 32'hc26b6f1d, 32'h42b8cb22, 32'h423e9ce5, 32'hc11c4eb4, 32'hc2ae4fd4, 32'h42a49c55};
test_weights[26304:26311] = '{32'h41eb9a1b, 32'hc291995e, 32'hc23e7341, 32'h410c9408, 32'h4218b730, 32'h41ca4fe8, 32'h429fdd27, 32'hc235286e};
test_bias[3288:3288] = '{32'hbf9b8489};
test_output[3288:3288] = '{32'hc6186f58};
test_input[26312:26319] = '{32'h41a21bf8, 32'hc284b282, 32'h40dbb579, 32'h419d6e10, 32'hc25c42f0, 32'hc16e07d4, 32'h3f1909b3, 32'hc23cc9b5};
test_weights[26312:26319] = '{32'h410d7ff1, 32'h428e69ec, 32'hc234d21f, 32'hc2bdc78b, 32'hc2af2af8, 32'hc203ac23, 32'h40addf80, 32'hc1ec2e2b};
test_bias[3289:3289] = '{32'hc26d9eb1};
test_output[3289:3289] = '{32'hc2925bde};
test_input[26320:26327] = '{32'hc215894e, 32'hc21fdae5, 32'hc2b99f75, 32'h424ffec9, 32'hc25fa26d, 32'hc27ecb96, 32'h42a8f7ea, 32'hc245c169};
test_weights[26320:26327] = '{32'hc186a151, 32'h418681ea, 32'hc289b52a, 32'hc20989a5, 32'h425a7b54, 32'hc2095826, 32'hc25e9d63, 32'hc2721eb0};
test_bias[3290:3290] = '{32'hc2a62d00};
test_output[3290:3290] = '{32'h44ed959d};
test_input[26328:26335] = '{32'h40d062d1, 32'h42729e69, 32'h41941825, 32'hc29da99b, 32'h42117486, 32'h42aa9b8c, 32'hc29de1b8, 32'hc2a15df7};
test_weights[26328:26335] = '{32'hc0962e15, 32'h4285d9a6, 32'h428825b5, 32'hc2c61f80, 32'hc2c53be6, 32'hc2aa8aa3, 32'hc2ba6472, 32'hc207e423};
test_bias[3291:3291] = '{32'hc210bfad};
test_output[3291:3291] = '{32'h46402f9e};
test_input[26336:26343] = '{32'hc27fd4fe, 32'h4235234c, 32'h42a41020, 32'h4253d28a, 32'h42a7547e, 32'hc298eb33, 32'hc2c02c2a, 32'h423aaf59};
test_weights[26336:26343] = '{32'hc228832e, 32'hc2b544d2, 32'h41f44446, 32'hc28575d2, 32'hc26c6fd3, 32'hc1e29c44, 32'hc1fb15b5, 32'hc1599f3d};
test_bias[3292:3292] = '{32'hc1f6355c};
test_output[3292:3292] = '{32'hc533458a};
test_input[26344:26351] = '{32'h422366a7, 32'h41246abe, 32'hc0531b03, 32'hc01c5d90, 32'h4128a006, 32'h42993be3, 32'hc29e53e7, 32'h4246205f};
test_weights[26344:26351] = '{32'h41a9637b, 32'h42188ff6, 32'h4084cae2, 32'hc28dacc3, 32'h41ed3189, 32'h420f1d7c, 32'h42669d85, 32'h4290aa36};
test_bias[3293:3293] = '{32'h429d787f};
test_output[3293:3293] = '{32'h455ef60e};
test_input[26352:26359] = '{32'h4231bff8, 32'hc287a9b9, 32'h4208acb7, 32'h421e5969, 32'h42a3d73f, 32'h420d9234, 32'h426a79ac, 32'h420e524a};
test_weights[26352:26359] = '{32'h42144578, 32'h4155ebbb, 32'hc1c833b6, 32'h40883862, 32'h3f91dfdc, 32'h425770c7, 32'h41ea617a, 32'h42767090};
test_bias[3294:3294] = '{32'h428a38e2};
test_output[3294:3294] = '{32'h45bc7fa3};
test_input[26360:26367] = '{32'h42854be2, 32'h42be76d7, 32'h41411a5f, 32'h424a0f4b, 32'hc2c7e8a6, 32'h4246fc6e, 32'hc20048f0, 32'hc21024fc};
test_weights[26360:26367] = '{32'h42bd3326, 32'h429f2ab7, 32'h412e181a, 32'hc10cde67, 32'hc28834f8, 32'h425c502e, 32'h410b25df, 32'h41db86e3};
test_bias[3295:3295] = '{32'hc120ca1e};
test_output[3295:3295] = '{32'h46aa9f80};
test_input[26368:26375] = '{32'h42913f42, 32'h420bf3b8, 32'h42056711, 32'h41b3c7ce, 32'hc1287ab9, 32'h42b41c03, 32'hc1620492, 32'hc1c211ec};
test_weights[26368:26375] = '{32'hc1516f07, 32'h4276c768, 32'hc130fac7, 32'hc29c0892, 32'h42b35270, 32'h42160cdc, 32'h428c012a, 32'hc291068e};
test_bias[3296:3296] = '{32'h423de08a};
test_output[3296:3296] = '{32'h451218fd};
test_input[26376:26383] = '{32'h41c24406, 32'h41d762c5, 32'h42aa5025, 32'hc201ac42, 32'h421a6105, 32'hc1c44c42, 32'h42bf7a4c, 32'hc08da6e9};
test_weights[26376:26383] = '{32'hc287fa32, 32'h422e2996, 32'h42931f3d, 32'hc21eec21, 32'h42653d3a, 32'h42bd5584, 32'hc21c332c, 32'h427afb5e};
test_bias[3297:3297] = '{32'hc1f124de};
test_output[3297:3297] = '{32'h45363f66};
test_input[26384:26391] = '{32'h4258eddf, 32'h4271b06b, 32'hc0ab4191, 32'hc1eea557, 32'h42ab3424, 32'hc21d74b7, 32'h42853e2d, 32'hc24d48d3};
test_weights[26384:26391] = '{32'h419fec38, 32'h42a8e25a, 32'h4277f1f3, 32'hc2a0ab55, 32'hc10abbf4, 32'h40987dda, 32'h42460e8c, 32'hc259fea6};
test_bias[3298:3298] = '{32'h4297c95b};
test_output[3298:3298] = '{32'h4652d2e0};
test_input[26392:26399] = '{32'h4229240c, 32'hc2661e6c, 32'h42a31bab, 32'h414346e4, 32'hc2ad9737, 32'hc25d08b4, 32'hc0acb25f, 32'h42c5ce04};
test_weights[26392:26399] = '{32'h424eb61f, 32'hc2bd6185, 32'h423c634b, 32'hbf495292, 32'h42146d43, 32'hc184dc11, 32'h42be1694, 32'h42923e1c};
test_bias[3299:3299] = '{32'hc2c73214};
test_output[3299:3299] = '{32'h467691b7};
test_input[26400:26407] = '{32'h42665127, 32'hc28cbe6b, 32'hc2992b7b, 32'h4194c8f7, 32'h42079075, 32'h41309832, 32'hc29d815b, 32'hc261512d};
test_weights[26400:26407] = '{32'hc1ba18e7, 32'h407aa7a4, 32'h423f9737, 32'hc261e31d, 32'hc260d6b5, 32'hc28aee4f, 32'hc13e5dbf, 32'hc006c5ed};
test_bias[3300:3300] = '{32'hc2b8d3b7};
test_output[3300:3300] = '{32'hc5fb5061};
test_input[26408:26415] = '{32'h4225925b, 32'h41a27f98, 32'h421963fa, 32'h422fa936, 32'h42839f08, 32'h411c5797, 32'hc2c1d32a, 32'hc2843ad6};
test_weights[26408:26415] = '{32'hc1091771, 32'h424227de, 32'hc2c182f7, 32'h42983158, 32'hc0c87f38, 32'hc26494e1, 32'h4282c283, 32'hc11d42dc};
test_bias[3301:3301] = '{32'hc0766209};
test_output[3301:3301] = '{32'hc5c7f14c};
test_input[26416:26423] = '{32'hc129a6fc, 32'h40854c7e, 32'hc19722fd, 32'hc28944d9, 32'hc226b7f5, 32'hc1f2ec19, 32'h42b4f960, 32'h42206ad8};
test_weights[26416:26423] = '{32'h3dd18f4e, 32'hc25ef7bd, 32'hc20699e1, 32'hc2748226, 32'hc07d905b, 32'hc2425437, 32'h41500d50, 32'h41533a68};
test_bias[3302:3302] = '{32'h427c7f26};
test_output[3302:3302] = '{32'h45fa3b48};
test_input[26424:26431] = '{32'h41258e43, 32'h42874acf, 32'h42775a21, 32'h42a0e822, 32'h427fe92d, 32'hc23f9c9b, 32'hc2630ad1, 32'h424cc66b};
test_weights[26424:26431] = '{32'hc2a41038, 32'hc2981c20, 32'h427ae4c8, 32'hc2bc2b90, 32'hc228c30e, 32'hc2928cb7, 32'hc013c974, 32'h41f21472};
test_bias[3303:3303] = '{32'h421b8420};
test_output[3303:3303] = '{32'hc5df93ef};
test_input[26432:26439] = '{32'h41b28cd6, 32'hc1452161, 32'hc289a04d, 32'h41099312, 32'hc1d36bbd, 32'h41a9a279, 32'h42b6fc52, 32'h42a97c8a};
test_weights[26432:26439] = '{32'h424dc8ab, 32'hc2906ddb, 32'hc28dfeee, 32'h4192139d, 32'h42a8593b, 32'hc1a58a49, 32'h41ebfa89, 32'h429768e3};
test_bias[3304:3304] = '{32'hc2a45de4};
test_output[3304:3304] = '{32'h46522546};
test_input[26440:26447] = '{32'hc24113af, 32'h4251fefc, 32'h4094de2d, 32'h422d5056, 32'hc2310561, 32'hc212b47a, 32'hc2aa785b, 32'hc15c7d7f};
test_weights[26440:26447] = '{32'h409484e3, 32'h42a12ead, 32'hc2904ab2, 32'h4259909b, 32'h42b5591c, 32'h4264ff41, 32'hc2c77036, 32'h4182d039};
test_bias[3305:3305] = '{32'h42aa6d36};
test_output[3305:3305] = '{32'h46014bc1};
test_input[26448:26455] = '{32'h42c7ba10, 32'h41b9b6f6, 32'hc2490e50, 32'h42b21b2c, 32'h42a9f2b4, 32'h42b64c1b, 32'h4291ab25, 32'hc26f3461};
test_weights[26448:26455] = '{32'hc24f831e, 32'hc20094d3, 32'hc284cfc5, 32'h427a192d, 32'h422e45ea, 32'hc26f4823, 32'hc1bc36b6, 32'h41a0c507};
test_bias[3306:3306] = '{32'hc2a60263};
test_output[3306:3306] = '{32'hc4dd3ac9};
test_input[26456:26463] = '{32'h4164b6fc, 32'h429a8237, 32'h427ddaa5, 32'hc20b2025, 32'h429b9c3e, 32'hc2b3a897, 32'hc1b67644, 32'h419a1b75};
test_weights[26456:26463] = '{32'hc289efbb, 32'h422b27ee, 32'h428bf5f7, 32'h42c139ae, 32'h42712125, 32'h3f3142f1, 32'hc28c2497, 32'hc015f5d5};
test_bias[3307:3307] = '{32'hc2bf943a};
test_output[3307:3307] = '{32'h461437d9};
test_input[26464:26471] = '{32'h4202c86d, 32'hc2c52536, 32'h42ae23f3, 32'h4280fa26, 32'h424c2cb4, 32'h41e27c2b, 32'hc2b188fa, 32'h42bb9d83};
test_weights[26464:26471] = '{32'hc2a71e3e, 32'hc2becce8, 32'hc28c1766, 32'h3f09ef8f, 32'hc1d3a6a8, 32'hc2a24343, 32'h429773ed, 32'h4156b499};
test_bias[3308:3308] = '{32'h41803433};
test_output[3308:3308] = '{32'hc6049b58};
test_input[26472:26479] = '{32'h42a87964, 32'hc1cb9cd8, 32'hc1ef14de, 32'h4298b1db, 32'h4277de2a, 32'h41861943, 32'h41bd3c82, 32'hc1cfe799};
test_weights[26472:26479] = '{32'h4293ad7f, 32'hc1502dbc, 32'hc11472cb, 32'h42c2afad, 32'hc1283b26, 32'hc0d0db88, 32'h418a35be, 32'hc136fc89};
test_bias[3309:3309] = '{32'hc20fa3db};
test_output[3309:3309] = '{32'h465d653c};
test_input[26480:26487] = '{32'hc209fdff, 32'hc2721d1e, 32'hc29deaa2, 32'hc142e81a, 32'hc2874d0f, 32'h42ac4add, 32'hc2991dd8, 32'h42a195ae};
test_weights[26480:26487] = '{32'hc2838dae, 32'h421f915d, 32'hc08eb824, 32'hc28d0316, 32'hc2936a5e, 32'hc2a278c0, 32'h42b8284a, 32'h42169b29};
test_bias[3310:3310] = '{32'h424ff4c0};
test_output[3310:3310] = '{32'hc5992d10};
test_input[26488:26495] = '{32'hc24df619, 32'h42823f54, 32'hc2bbdea6, 32'h42be206a, 32'h42bdfa55, 32'hc2974d3a, 32'h421941e5, 32'hc0d4d995};
test_weights[26488:26495] = '{32'hc0e8d10f, 32'hc1b8f772, 32'h41b89119, 32'hc2a9e733, 32'h423c0aae, 32'hc2882168, 32'hc1a7b85a, 32'hc26d00e9};
test_bias[3311:3311] = '{32'hc1fb3291};
test_output[3311:3311] = '{32'hc5097ea1};
test_input[26496:26503] = '{32'h4293f218, 32'h4202976f, 32'hc21caba9, 32'hc17c8c11, 32'hc147a923, 32'hc265bf54, 32'hc2b5bf6f, 32'h42a2239e};
test_weights[26496:26503] = '{32'hc2c4c304, 32'hc2c2e5dc, 32'hc1588dce, 32'hc2bdc6a5, 32'h421c1e31, 32'h42b207a3, 32'hc27bc0e3, 32'hc238c396};
test_bias[3312:3312] = '{32'hc1800f1c};
test_output[3312:3312] = '{32'hc63ca0b9};
test_input[26504:26511] = '{32'hc097acb1, 32'hc20b94be, 32'h42a9f9f4, 32'hc122db70, 32'h4203290f, 32'h426dd1f0, 32'h42c1ecef, 32'hc1b74eb0};
test_weights[26504:26511] = '{32'hc280c542, 32'h42a37dd6, 32'h4251468e, 32'h42b2861b, 32'h424d1a77, 32'h42809fba, 32'hc1c61150, 32'h40eb76c4};
test_bias[3313:3313] = '{32'h42c45742};
test_output[3313:3313] = '{32'h457b87e6};
test_input[26512:26519] = '{32'hc1266d0d, 32'h42ae8370, 32'hc0d7b6b5, 32'hc19e6cca, 32'hc1ab1a31, 32'h42b23a59, 32'h42258db1, 32'h41e266ca};
test_weights[26512:26519] = '{32'hc198555a, 32'h421a8c00, 32'h41c43fb1, 32'hc2189187, 32'hc2917462, 32'hc2a1e408, 32'h422a8b42, 32'h42556bb7};
test_bias[3314:3314] = '{32'hc2883d89};
test_output[3314:3314] = '{32'h44d57de7};
test_input[26520:26527] = '{32'hc2bc6f4f, 32'hc213d8c0, 32'h41914eae, 32'h424be470, 32'h40fcd65b, 32'hc1cb01ec, 32'hc2275e16, 32'hc292fd88};
test_weights[26520:26527] = '{32'hc003ad8a, 32'h42c7f7b1, 32'hc2ac378a, 32'hc2c026c2, 32'h42a5113d, 32'hc1b39386, 32'hc2be3334, 32'hc2998396};
test_bias[3315:3315] = '{32'h41502547};
test_output[3315:3315] = '{32'h445f09b4};
test_input[26528:26535] = '{32'hc29908f0, 32'h4155239c, 32'hc21ead92, 32'hc0a67c13, 32'h42b1f242, 32'hc1ffee38, 32'h40c59a9b, 32'h42056a3b};
test_weights[26528:26535] = '{32'h4279696f, 32'h42c46e43, 32'h42b5a81c, 32'h4286d1ea, 32'hc1eea253, 32'hc19ded3d, 32'h42c7c400, 32'hc2600810};
test_bias[3316:3316] = '{32'h42844969};
test_output[3316:3316] = '{32'hc62600b6};
test_input[26536:26543] = '{32'hc2b4c507, 32'h4257c701, 32'hc2c5c887, 32'hc275d5e3, 32'h41100f3a, 32'hc2bba4ed, 32'hc107e2bb, 32'hc23cfd79};
test_weights[26536:26543] = '{32'hc2750001, 32'hbf131287, 32'h42bacad5, 32'hc1aac2af, 32'hc2a9bd5e, 32'h4199e240, 32'h427d5797, 32'h419d62e1};
test_bias[3317:3317] = '{32'h42917d2a};
test_output[3317:3317] = '{32'hc5c775a2};
test_input[26544:26551] = '{32'hc20e2cd4, 32'hc2af4da4, 32'h424150cc, 32'hc0b59f47, 32'h426feb33, 32'hc19a5722, 32'hc0053a8f, 32'hc1d12610};
test_weights[26544:26551] = '{32'hc2b75863, 32'hc21e97ad, 32'hc20ae634, 32'hc2a4aee3, 32'hc1955158, 32'h412684da, 32'h42030be1, 32'hc0b98231};
test_bias[3318:3318] = '{32'h42afe798};
test_output[3318:3318] = '{32'h4588ae27};
test_input[26552:26559] = '{32'hc1d9c09d, 32'h41aaa83e, 32'hc28832ba, 32'hc19e7aa6, 32'hc1fc87e3, 32'hc2874177, 32'h42adfcd2, 32'hc281562f};
test_weights[26552:26559] = '{32'hc2ad452c, 32'hc2099bd7, 32'hc28b71fd, 32'h42b904b8, 32'h42aa754a, 32'hc2a1fd7a, 32'h4115f34d, 32'h422bbc93};
test_bias[3319:3319] = '{32'h403366eb};
test_output[3319:3319] = '{32'h45a7c3cd};
test_input[26560:26567] = '{32'hc2c386ad, 32'hc1ff0cc0, 32'hc1a9202f, 32'hc0d767e3, 32'hc21935a6, 32'h42b4f8f9, 32'h4250c93d, 32'hc011eee3};
test_weights[26560:26567] = '{32'hc253532d, 32'hc25b1c13, 32'hc2bdf53f, 32'h42baab9e, 32'hc09ec48e, 32'h42a8b95c, 32'h4268dc1a, 32'h42a04b69};
test_bias[3320:3320] = '{32'h418d7ae1};
test_output[3320:3320] = '{32'h4694584d};
test_input[26568:26575] = '{32'hc18f46a5, 32'h4294c31b, 32'h4238fa63, 32'h427372fb, 32'hc2ab46c9, 32'h426694b9, 32'h415fb920, 32'h41b99454};
test_weights[26568:26575] = '{32'h420f3021, 32'hc0d399dd, 32'hc2af42e9, 32'h4246f14e, 32'hc03004b4, 32'h4262fcb9, 32'h42b9c975, 32'hc203c3e3};
test_bias[3321:3321] = '{32'hc237447d};
test_output[3321:3321] = '{32'h44e5a8db};
test_input[26576:26583] = '{32'h40435e55, 32'hc2954441, 32'h428b6c2f, 32'hc28a5c32, 32'h428b77e5, 32'hc1c6bbe0, 32'hc0b921f6, 32'hc2ab4372};
test_weights[26576:26583] = '{32'hc2ba2333, 32'h41854d4e, 32'hc24bde0f, 32'hc1e61618, 32'hc22c87e9, 32'hc2b1afc2, 32'h423dc20d, 32'hc180a79e};
test_bias[3322:3322] = '{32'hc1a064aa};
test_output[3322:3322] = '{32'hc52f92f9};
test_input[26584:26591] = '{32'hc2a89a82, 32'hc2584b5d, 32'h42c63946, 32'hc249e25a, 32'hc2305107, 32'hc2bceeac, 32'h42b9da3f, 32'hc256bad5};
test_weights[26584:26591] = '{32'hc15464bc, 32'h412cfa06, 32'h419c8ed2, 32'h42998330, 32'hc0c45c7c, 32'hc23185c2, 32'hc2834834, 32'hc24ca08b};
test_bias[3323:3323] = '{32'hc2875349};
test_output[3323:3323] = '{32'hc3b31494};
test_input[26592:26599] = '{32'hc0de8a4a, 32'h42af1e29, 32'h4161ad33, 32'h42b49a1d, 32'h41cfcf8e, 32'hc28fee9f, 32'h4234560f, 32'hc2bdb2f4};
test_weights[26592:26599] = '{32'h42a8001d, 32'h42675936, 32'h42b51857, 32'h41b1504a, 32'hc2c7322f, 32'h42734e53, 32'hc21c214f, 32'hc23ab95c};
test_bias[3324:3324] = '{32'h41ae312a};
test_output[3324:3324] = '{32'h4559ba7d};
test_input[26600:26607] = '{32'hc182dad4, 32'hc292fa36, 32'h3e73d35a, 32'h42ac26d9, 32'h42b1c829, 32'hc1fe7ba3, 32'hc26d7ed5, 32'h42bf91ca};
test_weights[26600:26607] = '{32'hc2264c4a, 32'hc2571f22, 32'h42b5a36b, 32'hc17c6b26, 32'h41ac6f88, 32'h42b6e1f7, 32'hc2513e4f, 32'h42c0da0d};
test_bias[3325:3325] = '{32'h424594cd};
test_output[3325:3325] = '{32'h46659a5e};
test_input[26608:26615] = '{32'hc1c48881, 32'h42887961, 32'h42c048b0, 32'h42b8f9d5, 32'hc240eb99, 32'h40526e45, 32'hc1f20526, 32'h427dc47d};
test_weights[26608:26615] = '{32'hc22e83b0, 32'hc1fd64df, 32'hc2aea08a, 32'h422f57e0, 32'hc01f50f2, 32'h42bafa42, 32'hc25fd7b3, 32'h414166ae};
test_bias[3326:3326] = '{32'h42c14523};
test_output[3326:3326] = '{32'hc518ddeb};
test_input[26616:26623] = '{32'hbfcf051b, 32'h4295bcca, 32'h42b2cb35, 32'hc151dd48, 32'hc2838033, 32'h42b4d81b, 32'h427a0f78, 32'h418cf3e6};
test_weights[26616:26623] = '{32'hc1dac495, 32'hc1f2a650, 32'hc283c89e, 32'h41a5f5c4, 32'h42681999, 32'h42191f3d, 32'hc1c6391e, 32'h428f43cd};
test_bias[3327:3327] = '{32'hc2677aa2};
test_output[3327:3327] = '{32'hc60dff24};
test_input[26624:26631] = '{32'h42490208, 32'h3ed14162, 32'h40b65132, 32'h429deb90, 32'hc2b6ab2c, 32'h42816668, 32'hc2aef367, 32'hc2b62df6};
test_weights[26624:26631] = '{32'h423a6860, 32'h42c2caa3, 32'h429ca6d0, 32'hc2b38f7e, 32'h42a1ab35, 32'h4245618d, 32'hc09786dd, 32'h41e7e9df};
test_bias[3328:3328] = '{32'hc164b7c7};
test_output[3328:3328] = '{32'hc62710af};
test_input[26632:26639] = '{32'hc2113c87, 32'hc21f7727, 32'hc2c0e412, 32'hc1f71ac9, 32'hc2a315f7, 32'h4221a5a8, 32'hc2457c04, 32'h42bfeb0b};
test_weights[26632:26639] = '{32'h4244b12f, 32'hc2b02310, 32'h42986974, 32'h429c2831, 32'h41350771, 32'hc19fab7f, 32'h42706f16, 32'h42b74ba3};
test_bias[3329:3329] = '{32'h4257e387};
test_output[3329:3329] = '{32'hc572c432};
test_input[26640:26647] = '{32'hc2a81441, 32'hbe4757d0, 32'h42a7d650, 32'h41db42b7, 32'h418ab756, 32'h42a3b724, 32'h42100376, 32'h42938c52};
test_weights[26640:26647] = '{32'hc229f24b, 32'h42373ec7, 32'hbf352c6d, 32'h42c6868a, 32'hc2a4f0b4, 32'h42253603, 32'h41b376eb, 32'h3faf2940};
test_bias[3330:3330] = '{32'h4235a787};
test_output[3330:3330] = '{32'h460e9f2a};
test_input[26648:26655] = '{32'hc0ff9e98, 32'h40c653c6, 32'h428c1633, 32'hc23ec277, 32'h4243b715, 32'h42a15b31, 32'h42bc0e6b, 32'hc211c86e};
test_weights[26648:26655] = '{32'h41ddb530, 32'h42493e08, 32'h3f2372fc, 32'hc2c6ed2b, 32'h4186fcc2, 32'hc23fcc51, 32'h428ff572, 32'hc08e96ab};
test_bias[3331:3331] = '{32'hc1e4136f};
test_output[3331:3331] = '{32'h46088691};
test_input[26656:26663] = '{32'hc223a5db, 32'h4250b3e6, 32'h42310166, 32'hc2853883, 32'hc29e3a61, 32'hc2ba8fa0, 32'h409f9f6f, 32'h42155b88};
test_weights[26656:26663] = '{32'hc26c3380, 32'h4284ff16, 32'h41aa034e, 32'hc1b6ef95, 32'h41575c7a, 32'h42881540, 32'h3f9ce2af, 32'h420786ca};
test_bias[3332:3332] = '{32'hc20a0e11};
test_output[3332:3332] = '{32'h4507defc};
test_input[26664:26671] = '{32'hc19c8f1c, 32'h429875f8, 32'hc2737dae, 32'h4136c9b5, 32'hc24bede8, 32'hc23818f1, 32'hc27aef07, 32'hc2678040};
test_weights[26664:26671] = '{32'h4280d9c9, 32'h4299a27d, 32'hc2616b0f, 32'h42b924e9, 32'h4284376d, 32'h427fc9b4, 32'h42884faf, 32'hc2b13d19};
test_bias[3333:3333] = '{32'h425589e5};
test_output[3333:3333] = '{32'h4565c2fc};
test_input[26672:26679] = '{32'hc2a2568a, 32'h41d66e55, 32'hc26cc8bb, 32'h42911a28, 32'h42bfa3a2, 32'hc113f30a, 32'h419312b9, 32'hc15ed896};
test_weights[26672:26679] = '{32'hc23bc160, 32'h422ef16c, 32'h428eb4d0, 32'hc2bbb5f9, 32'hc2ac9ec9, 32'h42a0188a, 32'hc26e823b, 32'hc106b4ec};
test_bias[3334:3334] = '{32'h41dec312};
test_output[3334:3334] = '{32'hc67a3164};
test_input[26680:26687] = '{32'hc11e3eb4, 32'hc2b1b164, 32'hc261cc15, 32'hc1639888, 32'hc19b899d, 32'h42c00cb4, 32'hc18c5af1, 32'hc200ff5b};
test_weights[26680:26687] = '{32'h429321c8, 32'h42351c51, 32'hc1cc18cc, 32'h428866b2, 32'h42aac26f, 32'hc29a780c, 32'hc210e855, 32'h4229d2bb};
test_bias[3335:3335] = '{32'hc01e3ab7};
test_output[3335:3335] = '{32'hc65c3338};
test_input[26688:26695] = '{32'h4283db10, 32'h41dba9d2, 32'hc132d3a9, 32'hc2aa6987, 32'hc1881279, 32'h4229f9e3, 32'h41601048, 32'h428aa651};
test_weights[26688:26695] = '{32'h42491de3, 32'hc21ef230, 32'hc27f1167, 32'hc2699aad, 32'h41f668a2, 32'h4261f706, 32'h41275f2d, 32'h418e157e};
test_bias[3336:3336] = '{32'h426b32ab};
test_output[3336:3336] = '{32'h462f66e6};
test_input[26696:26703] = '{32'h41d101de, 32'h427c05ae, 32'h42301f75, 32'h42961035, 32'h40fb9f54, 32'h425f30a7, 32'h42179042, 32'hc16c84c6};
test_weights[26696:26703] = '{32'h423acebc, 32'h41a665ae, 32'h42af8dd7, 32'hc2aeaa45, 32'hc2587c55, 32'hc10df09b, 32'hc2979050, 32'hc0a21937};
test_bias[3337:3337] = '{32'h42166e1c};
test_output[3337:3337] = '{32'hc56fcb5e};
test_input[26704:26711] = '{32'h41a302c1, 32'h423cc46d, 32'h42b6b8b6, 32'h41806a46, 32'hc2a446fa, 32'h428984f0, 32'hc1023be9, 32'hc10d35bc};
test_weights[26704:26711] = '{32'hbf4ae540, 32'hc243fbe4, 32'h409ee05f, 32'hc2ac7c3b, 32'h42a8ef5e, 32'hc2a705a0, 32'hc21f00f1, 32'hc2129386};
test_bias[3338:3338] = '{32'h419877bc};
test_output[3338:3338] = '{32'hc66ea551};
test_input[26712:26719] = '{32'h42a002e2, 32'h42885203, 32'h428b65f7, 32'hc0838e47, 32'hc2b5d0ad, 32'hc2acf157, 32'hc165169b, 32'h42637778};
test_weights[26712:26719] = '{32'h42925ea9, 32'h41a0b1f7, 32'h42267c4e, 32'h411c854c, 32'h42a57c70, 32'hc261d12c, 32'h41909209, 32'h41354a84};
test_bias[3339:3339] = '{32'h42bde986};
test_output[3339:3339] = '{32'h45f7aac4};
test_input[26720:26727] = '{32'hc24ca425, 32'h421b33ac, 32'h424cba89, 32'h42b89886, 32'hc2b57b8d, 32'hc235970f, 32'h42878bda, 32'h428083d1};
test_weights[26720:26727] = '{32'hc2b687dd, 32'h42290eb4, 32'h429e5a83, 32'h42b56421, 32'h42196e5b, 32'h3d6365de, 32'h427eb8e7, 32'hc2a7d4ce};
test_bias[3340:3340] = '{32'hc2c7d3d0};
test_output[3340:3340] = '{32'h465be431};
test_input[26728:26735] = '{32'h4295f6fe, 32'h3c4033bb, 32'h42232a17, 32'hc2560769, 32'hc2925dff, 32'hc19a4e1a, 32'h408cfe03, 32'hc2b919cd};
test_weights[26728:26735] = '{32'hc28ab114, 32'hc28022c4, 32'hc276c315, 32'hc2651790, 32'h4230d2a5, 32'h3fac14d8, 32'h4276ce9e, 32'hc1e2398a};
test_bias[3341:3341] = '{32'h426d5d87};
test_output[3341:3341] = '{32'hc59b28b6};
test_input[26736:26743] = '{32'h41d73a53, 32'hc1059f22, 32'h41b02b0c, 32'hc2a80011, 32'hc268ae59, 32'hc2867400, 32'hc0a187ef, 32'h42c60227};
test_weights[26736:26743] = '{32'h4278577f, 32'hc228c7af, 32'hc22c3195, 32'hc22ddded, 32'hc20d9de8, 32'h4286ab37, 32'h429b3573, 32'hc29c19e9};
test_bias[3342:3342] = '{32'hc2832b6e};
test_output[3342:3342] = '{32'hc5b92f40};
test_input[26744:26751] = '{32'hc26cc02c, 32'h424f6323, 32'hc1e2c9cc, 32'h416db115, 32'h417d0284, 32'h4151100d, 32'hc29e95cb, 32'hc1b4fa37};
test_weights[26744:26751] = '{32'h41e4ebc8, 32'h4205b416, 32'h4297223c, 32'hc0cfb044, 32'hc235c0e3, 32'h41bf91c4, 32'hc298fc0c, 32'h429b8843};
test_bias[3343:3343] = '{32'h4073f53a};
test_output[3343:3343] = '{32'h44d51e3b};
test_input[26752:26759] = '{32'hc159510f, 32'hc1d9012c, 32'h42b34e81, 32'hc2a076fe, 32'hc2145315, 32'hc0d9e9d5, 32'h4267fea7, 32'hc2c0877f};
test_weights[26752:26759] = '{32'hc2425e6b, 32'hc21ddbff, 32'h42b5cb32, 32'hc290600f, 32'hc258ea8d, 32'hc17eb42a, 32'h426ae81e, 32'hc269ec51};
test_bias[3344:3344] = '{32'hc2a94fd2};
test_output[3344:3344] = '{32'h46d0eba3};
test_input[26760:26767] = '{32'hc25688c6, 32'h426e2713, 32'h423f1c8b, 32'h422651d3, 32'hc28188b0, 32'h411053af, 32'hc2861fcc, 32'h40f69087};
test_weights[26760:26767] = '{32'hc23ffe33, 32'hc1b2a75b, 32'h42119daf, 32'h4221494e, 32'h428d1ddd, 32'h429b1174, 32'hc2af2190, 32'h41be2f69};
test_bias[3345:3345] = '{32'hc0239449};
test_output[3345:3345] = '{32'h45d5d8bd};
test_input[26768:26775] = '{32'hc249605d, 32'h3fdf2f8a, 32'hc00e772c, 32'hc2bd0ef9, 32'h42a1129c, 32'hc2c2acab, 32'hc254e694, 32'h42186846};
test_weights[26768:26775] = '{32'hc2aa27e7, 32'hc1ae6096, 32'h428ec46a, 32'h4179be5f, 32'hc220e5b0, 32'h42815dea, 32'hc2c6bf2d, 32'h40498586};
test_bias[3346:3346] = '{32'hc299571d};
test_output[3346:3346] = '{32'hc4c70ca6};
test_input[26776:26783] = '{32'h428b1c3f, 32'h42b35e6a, 32'hc19da750, 32'h3f219e6f, 32'hc1ee432c, 32'hc1661d32, 32'h425fcd88, 32'hc104cf27};
test_weights[26776:26783] = '{32'h41f27fc0, 32'hc21bb26e, 32'hc1879f43, 32'h42a64a27, 32'hc1e6d393, 32'hc20601e8, 32'h42a28b2a, 32'h41ef3560};
test_bias[3347:3347] = '{32'hc2bab85f};
test_output[3347:3347] = '{32'h458e3707};
test_input[26784:26791] = '{32'h411ec58a, 32'hc2a2f470, 32'hc2b2cb57, 32'hc2700000, 32'hc281761e, 32'h428352ea, 32'hc055fccf, 32'h42b2ef63};
test_weights[26784:26791] = '{32'hc2b649c4, 32'h42ad31f6, 32'hc2aa68ef, 32'h41b5657f, 32'h42767a38, 32'hc2b97714, 32'hc2998aa2, 32'hc2603243};
test_bias[3348:3348] = '{32'h424974cb};
test_output[3348:3348] = '{32'hc680d18b};
test_input[26792:26799] = '{32'hc28a1571, 32'h41f7f62a, 32'hc2650a69, 32'h42c7f9a7, 32'h42666632, 32'h42453397, 32'h42929421, 32'hc1bc911a};
test_weights[26792:26799] = '{32'h40ad1500, 32'hc280f443, 32'h41cd1d4e, 32'hc1e28269, 32'hc26d0b79, 32'h40418ded, 32'h414a42e6, 32'h4209d6a3};
test_bias[3349:3349] = '{32'h42775517};
test_output[3349:3349] = '{32'hc6187d3f};
test_input[26800:26807] = '{32'hc22678f9, 32'h41d08554, 32'hc1c65dca, 32'hc2ae2569, 32'hc154248d, 32'hc2c4ded1, 32'h41dcf87c, 32'h42562d3b};
test_weights[26800:26807] = '{32'h420bfa28, 32'hc2603cbc, 32'h41323a58, 32'hc2369afd, 32'h42af7ef7, 32'h422d098f, 32'h41b42b6b, 32'h4286269c};
test_bias[3350:3350] = '{32'h3fa38b74};
test_output[3350:3350] = '{32'hc3d4d160};
test_input[26808:26815] = '{32'h42616155, 32'hc0bdda6a, 32'h42ba1aca, 32'h4133ddb9, 32'h418eb4a9, 32'h42366a02, 32'hc05a68d6, 32'hc2969584};
test_weights[26808:26815] = '{32'h41f670eb, 32'h41c22d43, 32'h40dd2995, 32'hc1e27dca, 32'h4254c239, 32'hc1b3f708, 32'hc2400852, 32'h427d9ac7};
test_bias[3351:3351] = '{32'hc225f47e};
test_output[3351:3351] = '{32'hc52fbc3c};
test_input[26816:26823] = '{32'h42b2e53a, 32'h41ca478e, 32'hc27b4159, 32'h41704e46, 32'h4288e594, 32'hc29780fc, 32'hc1e8af4c, 32'hc2bff953};
test_weights[26816:26823] = '{32'hc26ac227, 32'h4222a91d, 32'h42b143ee, 32'h42833a43, 32'h4241d40d, 32'h42316fb0, 32'h41fffe19, 32'h41408f70};
test_bias[3352:3352] = '{32'h40761576};
test_output[3352:3352] = '{32'hc62ac382};
test_input[26824:26831] = '{32'h424c2850, 32'hc290e2d4, 32'h42a95ff4, 32'hc2954f3e, 32'hc2854720, 32'h421b52a3, 32'h422ff0ef, 32'hc24ea3a3};
test_weights[26824:26831] = '{32'hc2994235, 32'hc23a5ebe, 32'hc25ac56d, 32'hc22ac457, 32'h42c256a3, 32'hc263da42, 32'hc2b42b7b, 32'hc245bf3e};
test_bias[3353:3353] = '{32'hc0bd9db3};
test_output[3353:3353] = '{32'hc63cc849};
test_input[26832:26839] = '{32'hc24cb002, 32'h4203cb04, 32'hc1a88d28, 32'h41c15b4f, 32'hc25d1a54, 32'h41bc4030, 32'hc20c9db3, 32'h4285d966};
test_weights[26832:26839] = '{32'hc2a5a1ad, 32'hc2b43c37, 32'h42ad46e0, 32'hc2a3aa94, 32'hc28e86d6, 32'hc1fd1fd7, 32'hc2834a41, 32'h429776c2};
test_bias[3354:3354] = '{32'hc236089d};
test_output[3354:3354] = '{32'h45f9b3b8};
test_input[26840:26847] = '{32'hc19a525f, 32'hc2654b3d, 32'h4183fe82, 32'hc2700de3, 32'hc17629c8, 32'hc2bf33f0, 32'hc286dd13, 32'h41ca9b49};
test_weights[26840:26847] = '{32'hc18906d7, 32'hc2c49d33, 32'h41ad0b92, 32'hc27287e4, 32'h41cc76d8, 32'h428231f2, 32'h414722ed, 32'h3e071ce6};
test_bias[3355:3355] = '{32'h42bcdd7c};
test_output[3355:3355] = '{32'h4522b442};
test_input[26848:26855] = '{32'h42c55aff, 32'h42a4477a, 32'h4064a740, 32'hc2b81b9b, 32'hc24aa3eb, 32'h4290b8fa, 32'hc2bc39ec, 32'h42ac82aa};
test_weights[26848:26855] = '{32'hbfe37984, 32'h4212e412, 32'h42348249, 32'hc1d6772c, 32'hc1ef9b80, 32'hc2475946, 32'hc294500c, 32'h42a38935};
test_bias[3356:3356] = '{32'h41fb431a};
test_output[3356:3356] = '{32'h468848fc};
test_input[26856:26863] = '{32'h3f2e7824, 32'h40a5d432, 32'hc2a0c94d, 32'hc21e230e, 32'h426e7a75, 32'hc1a6be5a, 32'hc29b7211, 32'h41d3ee10};
test_weights[26856:26863] = '{32'hc0a98196, 32'hc1f0212e, 32'h412b96ed, 32'h42c301b0, 32'hc1cc30a6, 32'hc187a8f9, 32'hbeaa4f25, 32'hc29cdd1b};
test_bias[3357:3357] = '{32'h4226aa89};
test_output[3357:3357] = '{32'hc5fbb465};
test_input[26864:26871] = '{32'hc20f79ce, 32'h415fa862, 32'hc25a9022, 32'h421c62b7, 32'hc12cd96c, 32'h42bd755e, 32'hc29419d3, 32'hc2654785};
test_weights[26864:26871] = '{32'hc0f08d64, 32'h409ab2bc, 32'h428b29a3, 32'h414a776e, 32'h42013827, 32'hc299c2b7, 32'hc2bb4a22, 32'hc23c1b74};
test_bias[3358:3358] = '{32'h408edc15};
test_output[3358:3358] = '{32'hc471d73d};
test_input[26872:26879] = '{32'h41f939c0, 32'hc1b678b7, 32'h423f7bc5, 32'h42b0146d, 32'h4268602a, 32'h4123cb14, 32'h42a16d7f, 32'h428d3e7d};
test_weights[26872:26879] = '{32'h419e66b5, 32'hc202f54c, 32'h42be9620, 32'hc0e654ed, 32'h42bf71c9, 32'hc248a2bf, 32'h42951fa2, 32'hc2b4cace};
test_bias[3359:3359] = '{32'hc2638feb};
test_output[3359:3359] = '{32'h461af185};
test_input[26880:26887] = '{32'hc215f5ca, 32'hc0e02942, 32'hc21bd026, 32'hc28e1fbb, 32'h41ec4a86, 32'h42c29ed5, 32'h415b2584, 32'hc1ac747d};
test_weights[26880:26887] = '{32'h42227769, 32'h40dade39, 32'h4258e708, 32'h42043473, 32'h40e65817, 32'h42516419, 32'h42c57723, 32'h4221c3e3};
test_bias[3360:3360] = '{32'hc10149e5};
test_output[3360:3360] = '{32'hc37c8f1d};
test_input[26888:26895] = '{32'hc2af1768, 32'hc2a24ef1, 32'hc2bc3a99, 32'h41bb1844, 32'h41dfd600, 32'hc28f8718, 32'hc1bc1fac, 32'h425d703d};
test_weights[26888:26895] = '{32'hc2a59fcc, 32'hc124ae99, 32'hc21e0d06, 32'hc2502a0e, 32'h426113cb, 32'hc1e83190, 32'h42b117af, 32'h429df040};
test_bias[3361:3361] = '{32'hc242335a};
test_output[3361:3361] = '{32'h4680ca01};
test_input[26896:26903] = '{32'h41dbcdce, 32'hc2a38db4, 32'hc2602c26, 32'h4280b5fa, 32'hc1517f52, 32'h42652de1, 32'hc245f298, 32'h4293787d};
test_weights[26896:26903] = '{32'h40997c07, 32'hc29e9763, 32'hc25c4418, 32'hc29f18a1, 32'h42af53ff, 32'hc2b614a0, 32'hc0d523b1, 32'hc22d0cb0};
test_bias[3362:3362] = '{32'hc285b857};
test_output[3362:3362] = '{32'hc59320e7};
test_input[26904:26911] = '{32'h41c6a2dd, 32'hc1a6ed05, 32'hc19fa7f1, 32'h420bb94d, 32'hc2854ba4, 32'hc209646e, 32'h427fc605, 32'hc288ea7e};
test_weights[26904:26911] = '{32'hc1d91e58, 32'hc03e3b75, 32'hc1fe6440, 32'h41a5de07, 32'h41dcc86e, 32'h4125b8a4, 32'h4233e3c8, 32'h4200294f};
test_bias[3363:3363] = '{32'hc054c4eb};
test_output[3363:3363] = '{32'hc440497c};
test_input[26912:26919] = '{32'h42aea20f, 32'hc25b57a8, 32'hc2ae3a28, 32'hc16ab6e9, 32'hc22bfbe7, 32'hc253c95b, 32'h42befcb5, 32'hc29fd2c7};
test_weights[26912:26919] = '{32'hc214ba7c, 32'h429fefcc, 32'h41bce719, 32'hc228f1dd, 32'hbf0c5dea, 32'hc1da5fd4, 32'h41aaa165, 32'h42948bd3};
test_bias[3364:3364] = '{32'hc189aa96};
test_output[3364:3364] = '{32'hc633f012};
test_input[26920:26927] = '{32'hc233d99c, 32'h4235c1bc, 32'hc20ef3da, 32'h40fa35f5, 32'hc1781725, 32'h42aaba0f, 32'hc219ee96, 32'h42936297};
test_weights[26920:26927] = '{32'hc2a3b3ee, 32'hc2b64a5c, 32'h42914c37, 32'h42b05ba1, 32'hc29b0201, 32'h42453b4b, 32'h4289aa54, 32'h428f514f};
test_bias[3365:3365] = '{32'hc0ec82fd};
test_output[3365:3365] = '{32'h45b118d6};
test_input[26928:26935] = '{32'h41326c7f, 32'h42945b5c, 32'hc23d03be, 32'h414cf1bb, 32'hc28248f8, 32'h41512611, 32'h426388bf, 32'h42c0d609};
test_weights[26928:26935] = '{32'h425e98b4, 32'hc2211585, 32'h42c5d68e, 32'hc18ad932, 32'hc295f9c7, 32'hc11142f1, 32'h4218e293, 32'hc216bed1};
test_bias[3366:3366] = '{32'hc1d8d9d7};
test_output[3366:3366] = '{32'hc578fa3e};
test_input[26936:26943] = '{32'hc0e22809, 32'h428041fc, 32'h42104c20, 32'h422d4dab, 32'hc269d004, 32'h424ae509, 32'hc2031122, 32'h41f5a868};
test_weights[26936:26943] = '{32'h42a56d73, 32'hc29e01e6, 32'hc0fac12f, 32'hc2bc4cd9, 32'hc274618e, 32'hc139b361, 32'h42046dff, 32'h4298f916};
test_bias[3367:3367] = '{32'h412b288a};
test_output[3367:3367] = '{32'hc5b3ddf1};
test_input[26944:26951] = '{32'hc0598b0e, 32'h408cdf7b, 32'h41f11fed, 32'h42715f62, 32'hc27ed985, 32'hc29d5cde, 32'hc22c0717, 32'h41747a23};
test_weights[26944:26951] = '{32'h420dd9b7, 32'hc15f0a19, 32'hc13a74dc, 32'hc187f211, 32'h42650234, 32'h4208ba5f, 32'h416bac79, 32'hc19e34b6};
test_bias[3368:3368] = '{32'h426834af};
test_output[3368:3368] = '{32'hc6091552};
test_input[26952:26959] = '{32'hc2afceab, 32'hc2be08e4, 32'h4230c65f, 32'h42881669, 32'h42b54907, 32'h4227809e, 32'h42a11ab0, 32'hc1d372b9};
test_weights[26952:26959] = '{32'hc29a3456, 32'h42808573, 32'h42794bf2, 32'hbf2d1014, 32'hc15922eb, 32'hc1c7ef17, 32'h42c68dcc, 32'hc14d3ff9};
test_bias[3369:3369] = '{32'hc1d1ff5b};
test_output[3369:3369] = '{32'h46131498};
test_input[26960:26967] = '{32'hc23aaa66, 32'h42039c7e, 32'h4226b03c, 32'hc1a301a9, 32'h428512df, 32'hc2c12c30, 32'hc17494ae, 32'hc28c97da};
test_weights[26960:26967] = '{32'h41be487f, 32'hc2c48522, 32'h423ce375, 32'h4257fcee, 32'h42627474, 32'hc2a9d1dd, 32'hc1393b2e, 32'h4236d156};
test_bias[3370:3370] = '{32'h4297efe3};
test_output[3370:3370] = '{32'h45ace5a3};
test_input[26968:26975] = '{32'hc2829a38, 32'h4184af94, 32'h42a180e6, 32'h4179e2db, 32'h410945db, 32'h42565663, 32'h42699961, 32'hc2a414c4};
test_weights[26968:26975] = '{32'h42a9ae44, 32'h4223443d, 32'hc278ed92, 32'hc1064a33, 32'hc13d635f, 32'hc2b1b2dc, 32'hc2849c59, 32'hc0866f7b};
test_bias[3371:3371] = '{32'h42583c22};
test_output[3371:3371] = '{32'hc68f673d};
test_input[26976:26983] = '{32'h4172399e, 32'hc2785728, 32'hc13956b3, 32'h42c14b6e, 32'h427346dc, 32'h41e0e29b, 32'hc2877c61, 32'hc2679d8b};
test_weights[26976:26983] = '{32'hc2196fe5, 32'h41a32e12, 32'h42644299, 32'h41566d87, 32'hc2bb2446, 32'h428898e1, 32'hbe0e287a, 32'hc1bb2f16};
test_bias[3372:3372] = '{32'h429b9bd9};
test_output[3372:3372] = '{32'hc55d5d41};
test_input[26984:26991] = '{32'h41fb3851, 32'h4273818c, 32'h41f5bc10, 32'h42c72ee6, 32'h426d1621, 32'hc28d80db, 32'hc21765d9, 32'hc2b4ed8b};
test_weights[26984:26991] = '{32'hc1adbfce, 32'hc2c0aee0, 32'hc120df2e, 32'hc2167e81, 32'h42c0550f, 32'h427b8a80, 32'h42377e39, 32'h428a22a4};
test_bias[3373:3373] = '{32'h42510e2d};
test_output[3373:3373] = '{32'hc6870881};
test_input[26992:26999] = '{32'hc0c5beb1, 32'hc225823b, 32'h4196d9d1, 32'h422f84e4, 32'h423b3575, 32'hc2a0f306, 32'hc2649cd5, 32'hc1ced3a3};
test_weights[26992:26999] = '{32'hc28cf80a, 32'hc256ecd0, 32'h4105b8b3, 32'h41e2d945, 32'h417542dc, 32'h4227392e, 32'hc1b38550, 32'h428883b4};
test_bias[3374:3374] = '{32'hc177c79c};
test_output[3374:3374] = '{32'h44650871};
test_input[27000:27007] = '{32'hc28ccffa, 32'h428c665b, 32'h4179e0bf, 32'h426d252d, 32'hc18e179f, 32'hc29fe521, 32'h42be1789, 32'h4216394a};
test_weights[27000:27007] = '{32'hc266ead5, 32'h427f6b2a, 32'h428b0669, 32'hc21f5497, 32'h42985d14, 32'h41885faf, 32'h42bad4e8, 32'hc295b268};
test_bias[3375:3375] = '{32'h42a54101};
test_output[3375:3375] = '{32'h46274690};
test_input[27008:27015] = '{32'h419f2af7, 32'hc03ff1cf, 32'hc2876a6f, 32'hc0d2ccff, 32'hc229d857, 32'hc21eca04, 32'h42c70209, 32'h415929eb};
test_weights[27008:27015] = '{32'hc2938004, 32'hc0a33dc3, 32'h42156769, 32'hc2a54907, 32'hbea06fad, 32'hc0175799, 32'hc2af07ae, 32'h412eb66b};
test_bias[3376:3376] = '{32'hc27cbeef};
test_output[3376:3376] = '{32'hc63ac1dd};
test_input[27016:27023] = '{32'h421ee180, 32'hc2ad4e3c, 32'hc14c6726, 32'h42362765, 32'h42a004fd, 32'h428f327f, 32'hc2645bf6, 32'h42ad1131};
test_weights[27016:27023] = '{32'h4273e38c, 32'hc2478646, 32'h426fb313, 32'hc2a49d87, 32'h4105a6d7, 32'h405167fb, 32'hc2a7ce0a, 32'hc15f82d4};
test_bias[3377:3377] = '{32'h4258b805};
test_output[3377:3377] = '{32'h45d3831b};
test_input[27024:27031] = '{32'h42a6fb5c, 32'hc17981dd, 32'hc29bb6d2, 32'hc0cabe4e, 32'h429d587e, 32'h41b33a58, 32'h4291dca1, 32'hc12488df};
test_weights[27024:27031] = '{32'h428c5acc, 32'hc2b4a367, 32'hc28f624a, 32'h429e4604, 32'hc20f1922, 32'h426ca73a, 32'hc2539ec4, 32'hc1cefece};
test_bias[3378:3378] = '{32'hc01a4375};
test_output[3378:3378] = '{32'h45e30194};
test_input[27032:27039] = '{32'hc2a8b0e4, 32'hc10c2758, 32'h426fc079, 32'h42b9f23a, 32'hc2b487cd, 32'h4220f37d, 32'hc15ef83f, 32'hc2bfc141};
test_weights[27032:27039] = '{32'h42a2087f, 32'hc2ba021f, 32'hc20d182a, 32'h425e5e02, 32'h42c19b61, 32'hc27efe99, 32'h428367aa, 32'hc2860813};
test_bias[3379:3379] = '{32'h4215e955};
test_output[3379:3379] = '{32'hc608413a};
test_input[27040:27047] = '{32'h41de91de, 32'h4223f28e, 32'hbe7ee1a3, 32'hc2b42e29, 32'hc26abe64, 32'h425ed10d, 32'hbf841a4f, 32'hc1a75de2};
test_weights[27040:27047] = '{32'hc237aa0b, 32'h429cebf5, 32'hc26b03b2, 32'hc040d17b, 32'hc230f2ac, 32'h42c197c8, 32'hc29e0e11, 32'hc2a29575};
test_bias[3380:3380] = '{32'h40bfa7c5};
test_output[3380:3380] = '{32'h463b8312};
test_input[27048:27055] = '{32'hc086428f, 32'h427c1c63, 32'hc2798f26, 32'h41290399, 32'h424917df, 32'hc2a35c3d, 32'h41c65797, 32'hc252d086};
test_weights[27048:27055] = '{32'hc1bd1859, 32'hc19ed5dc, 32'hc27c5972, 32'hc192282b, 32'hc25a8954, 32'hc17fc3bb, 32'h416fb3e5, 32'h42a062bb};
test_bias[3381:3381] = '{32'h42897273};
test_output[3381:3381] = '{32'hc524c724};
test_input[27056:27063] = '{32'hc2431b36, 32'h42c742be, 32'hc183b344, 32'hc1665c17, 32'h4207afcc, 32'hc185f689, 32'hc18a6066, 32'hc28a4d28};
test_weights[27056:27063] = '{32'h42458104, 32'hc2053653, 32'hc2c25b91, 32'h418c0ee6, 32'hc28d3ba1, 32'h41de2b21, 32'h40c7d43a, 32'hc23cc42d};
test_bias[3382:3382] = '{32'hc28e7735};
test_output[3382:3382] = '{32'hc581d828};
test_input[27064:27071] = '{32'hc27fff31, 32'h427edad3, 32'hc2c4dff6, 32'h41f932d7, 32'h41919dbb, 32'hc1e3297c, 32'h41ab07b0, 32'hc2c37c8f};
test_weights[27064:27071] = '{32'hc130e2cc, 32'h4238a591, 32'hc2867613, 32'hc0fe663c, 32'h4289a4a6, 32'hc28b819a, 32'h425bac22, 32'hc2bead90};
test_bias[3383:3383] = '{32'h42c48594};
test_output[3383:3383] = '{32'h46ba46f1};
test_input[27072:27079] = '{32'h421777d2, 32'h4199efb1, 32'h425ad045, 32'h421b91dd, 32'h42c7c7d7, 32'h41900c4d, 32'h4296c024, 32'h42886dca};
test_weights[27072:27079] = '{32'hc14eee53, 32'hc11a2193, 32'h42bd6ccb, 32'h41f6a0f9, 32'h4266443a, 32'h426c62f3, 32'hc236d147, 32'h420fb9c4};
test_bias[3384:3384] = '{32'h41b00f94};
test_output[3384:3384] = '{32'h46346e01};
test_input[27080:27087] = '{32'h42153aab, 32'hc1c4bc9b, 32'hc268f382, 32'hc250a29f, 32'h428ded3e, 32'hc24ce24d, 32'hc29f689a, 32'hc1b5b761};
test_weights[27080:27087] = '{32'hc27ff3ba, 32'hc2061df9, 32'h409da93d, 32'h428f7c75, 32'hc1be576b, 32'h42b88868, 32'hc1b74b1e, 32'hc2b09cea};
test_bias[3385:3385] = '{32'hc21266c7};
test_output[3385:3385] = '{32'hc6004a78};
test_input[27088:27095] = '{32'hc2c63dda, 32'hc20be630, 32'hc16b190a, 32'h423c1113, 32'h42945666, 32'h411b2bbe, 32'hc2711803, 32'h41193e45};
test_weights[27088:27095] = '{32'hc1c1c80e, 32'hc22f0263, 32'hc19d0538, 32'h41a5f9a2, 32'h429be7c6, 32'h42a8713d, 32'hc28b18cb, 32'h41515be9};
test_bias[3386:3386] = '{32'hc2b7e1f3};
test_output[3386:3386] = '{32'h467a4b33};
test_input[27096:27103] = '{32'hc295d967, 32'h42c474f1, 32'h428acadc, 32'h42aa935f, 32'hc1e34d37, 32'h42b28bae, 32'h40f7f8b0, 32'h42a4f344};
test_weights[27096:27103] = '{32'h42b74f54, 32'hc27ca8c9, 32'h42a9c328, 32'hc2288dd6, 32'h428d579f, 32'h425362e8, 32'hc240e8d0, 32'hc2434598};
test_bias[3387:3387] = '{32'hc2b0ae83};
test_output[3387:3387] = '{32'hc6442722};
test_input[27104:27111] = '{32'hc11ab13b, 32'hc2b8e018, 32'hc2618224, 32'h4223cd40, 32'h425771bb, 32'hc0c71d8f, 32'hc17a49b2, 32'h4247b1bc};
test_weights[27104:27111] = '{32'hc00f4901, 32'hc29f8a7a, 32'h424246e2, 32'h418a543e, 32'h40754ab7, 32'hc29ce888, 32'h42a0dcc9, 32'h42485cb6};
test_bias[3388:3388] = '{32'hc2b90087};
test_output[3388:3388] = '{32'h45e14f90};
test_input[27112:27119] = '{32'h4264efd1, 32'h429f126d, 32'h427ec99f, 32'hc28191f4, 32'hc2131ae7, 32'hc22a3847, 32'h42bdae3b, 32'h421c43d8};
test_weights[27112:27119] = '{32'hc10a2d5f, 32'hc0c78eec, 32'hc28ea685, 32'hc25d6688, 32'hc205b813, 32'hc24d43f3, 32'hc23e173a, 32'hc2b85052};
test_bias[3389:3389] = '{32'hc28e2e09};
test_output[3389:3389] = '{32'hc5d1c674};
test_input[27120:27127] = '{32'h42489187, 32'h424dc115, 32'h41b8ecea, 32'h42b52343, 32'h3f56e8eb, 32'h40935750, 32'hc28c3b40, 32'hc22c6004};
test_weights[27120:27127] = '{32'hc16e70f0, 32'h414c1286, 32'hc23b87dd, 32'hc23e793a, 32'hc2b60069, 32'hc0fd1b82, 32'h41a44ae7, 32'h42c4c64b};
test_bias[3390:3390] = '{32'h40938544};
test_output[3390:3390] = '{32'hc6302ea3};
test_input[27128:27135] = '{32'hc2986a56, 32'hc1d269bb, 32'hc1b59009, 32'h4239abf4, 32'hc28e3ff2, 32'hc265dd31, 32'h429bc441, 32'hc29134eb};
test_weights[27128:27135] = '{32'h42bcc09e, 32'h424175aa, 32'hc1a6b239, 32'hc14ff9f0, 32'h429ad474, 32'h41472170, 32'hc211ce99, 32'h42a0fae6};
test_bias[3391:3391] = '{32'hbf22b9b4};
test_output[3391:3391] = '{32'hc6b7970e};
test_input[27136:27143] = '{32'h414c9668, 32'h3ee099ca, 32'hc281d762, 32'h4288e11c, 32'h42041e96, 32'h425126a5, 32'hc22af637, 32'h418399a2};
test_weights[27136:27143] = '{32'h42850769, 32'hc2665027, 32'hc22d07e7, 32'hc1d5360e, 32'h42a0f40d, 32'h4272e52b, 32'h424c949c, 32'h41ba501a};
test_bias[3392:3392] = '{32'hc1d9c147};
test_output[3392:3392] = '{32'h45b5a5bb};
test_input[27144:27151] = '{32'h40bfe141, 32'hc1e9d693, 32'hc2901e97, 32'hc255bf39, 32'h4152cc99, 32'h41a274c0, 32'h4216fa5a, 32'hc1b57efd};
test_weights[27144:27151] = '{32'h42c50738, 32'hc25b4be9, 32'hc288854b, 32'hc2bbd4fe, 32'h4281084f, 32'h41f6af7d, 32'hc22780ca, 32'h41b3a0e7};
test_bias[3393:3393] = '{32'h42c173cb};
test_output[3393:3393] = '{32'h46357615};
test_input[27152:27159] = '{32'hc2183420, 32'h419c7e07, 32'h41be972a, 32'hc1a3ea76, 32'hc23c72d4, 32'h42789c3a, 32'h41c3904e, 32'hc28f942b};
test_weights[27152:27159] = '{32'h426f1b68, 32'hc2705e18, 32'hc2c6d15b, 32'hc0db6c7c, 32'h40877290, 32'hc27edf5d, 32'hc22f3e8f, 32'h42adf638};
test_bias[3394:3394] = '{32'h42b115a2};
test_output[3394:3394] = '{32'hc6855083};
test_input[27160:27167] = '{32'hc0fd8c53, 32'h42890522, 32'hc1c3be96, 32'hc2818ecd, 32'h42808fd9, 32'h425215e1, 32'hc2870702, 32'h428c7e59};
test_weights[27160:27167] = '{32'hc2068315, 32'hc1d7fc55, 32'h41dc2e0a, 32'h424b7726, 32'h423820ba, 32'h4296ca60, 32'hc1438d2b, 32'hc2bfd291};
test_bias[3395:3395] = '{32'h42290743};
test_output[3395:3395] = '{32'hc58cb72f};
test_input[27168:27175] = '{32'h42b529ed, 32'hc2944959, 32'hc29d13e3, 32'h41ea34a5, 32'hc20fa123, 32'h42a3437c, 32'h424b7c39, 32'h42826e5f};
test_weights[27168:27175] = '{32'hc2a2cdfc, 32'hc22257fc, 32'h421c85f2, 32'h42546ccb, 32'hc1b7f97f, 32'hc275feb2, 32'hc2bdfffc, 32'hc1df57bb};
test_bias[3396:3396] = '{32'h42a0ee12};
test_output[3396:3396] = '{32'hc68214e7};
test_input[27176:27183] = '{32'h42b658e6, 32'hc24d0a7c, 32'h40c1d1cf, 32'hc2a9d764, 32'h402d81dc, 32'hc1f6615f, 32'hc2b81d29, 32'hc097a5e9};
test_weights[27176:27183] = '{32'hc2a7d990, 32'h428e0364, 32'hc18d527a, 32'h41de3126, 32'h41f6cfc9, 32'hc2a95841, 32'h42119cf7, 32'h4212e640};
test_bias[3397:3397] = '{32'hc2a5b640};
test_output[3397:3397] = '{32'hc665477a};
test_input[27184:27191] = '{32'h423927e6, 32'hc2975283, 32'h4026761c, 32'hc270869e, 32'hc284833d, 32'hc2a22998, 32'hc1ea236b, 32'hc2c31d4a};
test_weights[27184:27191] = '{32'hc2876b76, 32'h41cbe561, 32'hc2b64006, 32'hc2050c6d, 32'hc1933499, 32'h429e5f3d, 32'hc2a4351c, 32'h429c18b7};
test_bias[3398:3398] = '{32'h4286987a};
test_output[3398:3398] = '{32'hc6553310};
test_input[27192:27199] = '{32'hc27dffa4, 32'hc26a4f07, 32'h425865a7, 32'hc2b0fe25, 32'hc2a5a48c, 32'h41ae2d55, 32'h42b9751b, 32'hc2596d71};
test_weights[27192:27199] = '{32'hc0600976, 32'h41354642, 32'h41a49537, 32'hc28e6b99, 32'hc2391f7e, 32'h42885ade, 32'h4232590b, 32'hc2140b2f};
test_bias[3399:3399] = '{32'h41c90fda};
test_output[3399:3399] = '{32'h46903c8b};
test_input[27200:27207] = '{32'h42547c13, 32'h429b9e19, 32'h41a5f262, 32'hc018d4c4, 32'hc240a9ba, 32'hc228cd03, 32'hc25bf2a0, 32'hc2932ca0};
test_weights[27200:27207] = '{32'hc2ae77a3, 32'hc21cc6fa, 32'hc24df3e3, 32'hc233cd36, 32'h42432332, 32'hc1abd5d3, 32'hc2bdff01, 32'hc2922ae6};
test_bias[3400:3400] = '{32'h4188f69e};
test_output[3400:3400] = '{32'h4404cc16};
test_input[27208:27215] = '{32'hc2abf119, 32'h42a40de5, 32'h40510add, 32'h42ad4df7, 32'hc2677c10, 32'hc26f8a21, 32'hc268affa, 32'h42bf7775};
test_weights[27208:27215] = '{32'hc0e449b1, 32'h4249a7c5, 32'hc290eb7f, 32'hc1e55912, 32'h41ed7524, 32'hc1262879, 32'h42428a77, 32'hc2ad9cba};
test_bias[3401:3401] = '{32'hc24b4050};
test_output[3401:3401] = '{32'hc620495e};
test_input[27216:27223] = '{32'h429d4d4f, 32'hc2b83ab2, 32'h42970b2f, 32'hbff4bb1c, 32'hc272974e, 32'hc2c6a4b1, 32'hc296bc93, 32'h422fe9bc};
test_weights[27216:27223] = '{32'hc203ff12, 32'h41d3ebc2, 32'hc1701d5a, 32'h420f1965, 32'h42a21923, 32'hc2a684b2, 32'hc28b8177, 32'hc1203035};
test_bias[3402:3402] = '{32'h4186f477};
test_output[3402:3402] = '{32'h44f3cd1f};
test_input[27224:27231] = '{32'h40d1a711, 32'h4259f83d, 32'hc2506592, 32'hc23afc3c, 32'hc1e10032, 32'hbe8fef8c, 32'h420f1bb4, 32'hc21463f4};
test_weights[27224:27231] = '{32'h4207a9ef, 32'hc283d8f6, 32'hc27bddfc, 32'hc2a44d66, 32'h415197ad, 32'h42571f20, 32'h40b8f7ad, 32'h4197fe31};
test_bias[3403:3403] = '{32'hc286e8dc};
test_output[3403:3403] = '{32'h452f19f5};
test_input[27232:27239] = '{32'h42ad2943, 32'h41f40dc6, 32'h424f44c9, 32'h42c686a6, 32'hc21e5468, 32'hc25a62cc, 32'hbf3dc54e, 32'h41b8c3b9};
test_weights[27232:27239] = '{32'h41c4cafb, 32'h3f1b08fc, 32'hc200f791, 32'h42aa11c2, 32'hc12de884, 32'h41d5a58c, 32'hc2a058b8, 32'hc19db273};
test_bias[3404:3404] = '{32'hc2149b16};
test_output[3404:3404] = '{32'h45e90cd8};
test_input[27240:27247] = '{32'h42446b03, 32'hc2ac2a16, 32'hc242cc86, 32'hc2930460, 32'h40d7aa29, 32'h426974b6, 32'h4254684b, 32'h42acb61c};
test_weights[27240:27247] = '{32'hc2485bc0, 32'h3fc0a82f, 32'h42be8616, 32'hc2c5a5c4, 32'hc26cd2e4, 32'hc2aaf423, 32'h423d71da, 32'h42c09e47};
test_bias[3405:3405] = '{32'hc20bcaea};
test_output[3405:3405] = '{32'h45aa285c};
test_input[27248:27255] = '{32'h403cb56d, 32'hc106035a, 32'h4029eaa2, 32'hc20875d6, 32'hc1557f73, 32'hc2a9a149, 32'hc16ee57f, 32'hc24561a0};
test_weights[27248:27255] = '{32'hc19ad423, 32'hc2c13f77, 32'hc27ddd22, 32'hc2acc589, 32'h418f4f0e, 32'hc298c95e, 32'h42bfac17, 32'hc18d8ed1};
test_bias[3406:3406] = '{32'h42564a37};
test_output[3406:3406] = '{32'h4610cb6f};
test_input[27256:27263] = '{32'h4208e3d8, 32'hc13060ce, 32'h425581e7, 32'h424e9af5, 32'hc202fb00, 32'h41d075ff, 32'hc29b6798, 32'hc208051c};
test_weights[27256:27263] = '{32'h4287e1fa, 32'hc29a128f, 32'hc0a063ba, 32'h4169240d, 32'hc03afec1, 32'h41e2ac2e, 32'hc2c13495, 32'hc2aa6513};
test_bias[3407:3407] = '{32'h42999636};
test_output[3407:3407] = '{32'h4669f675};
test_input[27264:27271] = '{32'h4252ddc0, 32'h42bdbf25, 32'h42a11001, 32'hc26a1749, 32'h4201b005, 32'h3f8b8426, 32'h429c8415, 32'h42b2a26a};
test_weights[27264:27271] = '{32'hc152849c, 32'h42928504, 32'hc2550e10, 32'hc1bb8677, 32'h42ae6f84, 32'h41b82bdd, 32'hbdeebbdf, 32'h3f08fb81};
test_bias[3408:3408] = '{32'h400489ab};
test_output[3408:3408] = '{32'h45c2c671};
test_input[27272:27279] = '{32'hc28c8e31, 32'hc287fe85, 32'hc2537aa3, 32'hc26c74f3, 32'h4288a198, 32'hc0ae574a, 32'hc2900556, 32'hc2ba1906};
test_weights[27272:27279] = '{32'hc16f02ff, 32'hc254a6c0, 32'h42770dbb, 32'h41800fd5, 32'hc29a670d, 32'hc0e9abf5, 32'h42823461, 32'hc239b760};
test_bias[3409:3409] = '{32'hc09c95f8};
test_output[3409:3409] = '{32'hc5a10fec};
test_input[27280:27287] = '{32'hc287e735, 32'h428d7cac, 32'hc27f0cae, 32'h41ac73cd, 32'h4176f6a1, 32'h42053d15, 32'h42671d55, 32'hc1b4baf9};
test_weights[27280:27287] = '{32'h425452bd, 32'h42bc9d8e, 32'hc290f479, 32'hc29a0dd2, 32'hc1686d86, 32'h4229e2d4, 32'h41158b6d, 32'hc2780280};
test_bias[3410:3410] = '{32'h42c26290};
test_output[3410:3410] = '{32'h46109840};
test_input[27288:27295] = '{32'h427f522a, 32'hc25340e2, 32'h422d3678, 32'hc233bd1f, 32'h42355fc2, 32'h42c0b031, 32'h40ac4a86, 32'h423f3c7d};
test_weights[27288:27295] = '{32'hc2249a2e, 32'hc29248db, 32'h421d6085, 32'hc22027c3, 32'hc19ee1e8, 32'hc22deeb6, 32'h425ac82a, 32'h420375bc};
test_bias[3411:3411] = '{32'hc201f797};
test_output[3411:3411] = '{32'h44b94ed6};
test_input[27296:27303] = '{32'h4229199c, 32'h40e56e52, 32'hc2555443, 32'h4288f444, 32'hc26c8c34, 32'hc271ff91, 32'hc24836df, 32'hc1f3f461};
test_weights[27296:27303] = '{32'hc0ac262d, 32'h405f71ec, 32'h42a68140, 32'h424c0231, 32'h41dbcb9d, 32'hc149a281, 32'hc2733cdd, 32'h4296b1d0};
test_bias[3412:3412] = '{32'h41a7d58a};
test_output[3412:3412] = '{32'hc49ba7b0};
test_input[27304:27311] = '{32'hc2a2d69e, 32'h42288cdd, 32'hc27197e4, 32'hc2490201, 32'h428aeb9f, 32'h422ba718, 32'h426545ac, 32'hc1e6125c};
test_weights[27304:27311] = '{32'hbfd428ff, 32'hc28ef70e, 32'h427d9075, 32'h421e2147, 32'h4203e3af, 32'hc25a531b, 32'h41dc5300, 32'h42947eee};
test_bias[3413:3413] = '{32'hc11277a5};
test_output[3413:3413] = '{32'hc611793e};
test_input[27312:27319] = '{32'h41967685, 32'hc25841ab, 32'h42ba608b, 32'hc296a5b3, 32'h41f1e73d, 32'hc2c31dae, 32'hc2128694, 32'hc2b3c431};
test_weights[27312:27319] = '{32'hc1cabb78, 32'h421987c4, 32'h409432eb, 32'hc21be0f5, 32'hc17fe354, 32'h4186014c, 32'hc249bfbb, 32'h40fa31a3};
test_bias[3414:3414] = '{32'hc11ef216};
test_output[3414:3414] = '{32'hc327aedc};
test_input[27320:27327] = '{32'h42965622, 32'h429ff9ad, 32'h418dfcf4, 32'hc2ba3b19, 32'h422f26a8, 32'hc2560755, 32'h428c5bae, 32'hc2873a31};
test_weights[27320:27327] = '{32'h42a0596e, 32'h424fc52c, 32'hc25b3d51, 32'h402c61d7, 32'h42679baa, 32'hc292f796, 32'hc006b5f1, 32'h42314415};
test_bias[3415:3415] = '{32'h429de64e};
test_output[3415:3415] = '{32'h46411f88};
test_input[27328:27335] = '{32'hc22bfe8c, 32'h41d84bf8, 32'hc16563a2, 32'hc27a5b7f, 32'h4248d949, 32'h413d8733, 32'h42b933f0, 32'hc296b717};
test_weights[27328:27335] = '{32'h41237a9f, 32'h429f8c8f, 32'hc194f0ff, 32'hc2901d15, 32'h42882c97, 32'h425fa8b6, 32'h417cee8f, 32'h4214e17b};
test_bias[3416:3416] = '{32'h41d06136};
test_output[3416:3416] = '{32'h4610b2b0};
test_input[27336:27343] = '{32'h42426b85, 32'h425399b0, 32'hc256bd8d, 32'hc1212241, 32'hc2a2bdd9, 32'h42c286d1, 32'hc29fa04f, 32'hc20a0152};
test_weights[27336:27343] = '{32'hc1a9a261, 32'h42ac1430, 32'hc2c75bca, 32'hc2b4c5ab, 32'h42c32783, 32'hc2bbb10d, 32'hc25ff22d, 32'h42c1bb7a};
test_bias[3417:3417] = '{32'hc1e7a51a};
test_output[3417:3417] = '{32'hc5c15e35};
test_input[27344:27351] = '{32'h4298d476, 32'h41123983, 32'h42924a93, 32'h42a784a9, 32'h41cedec2, 32'h42bf8441, 32'h41953595, 32'h420b5b2d};
test_weights[27344:27351] = '{32'h4254a7d6, 32'h428686a3, 32'hc23f6be7, 32'hc285ddb1, 32'h42bbdfbf, 32'h42413596, 32'hbf7ca11a, 32'hc2b0154c};
test_bias[3418:3418] = '{32'h42773af7};
test_output[3418:3418] = '{32'hc3c76e41};
test_input[27352:27359] = '{32'h42b9a5f5, 32'hc1463d52, 32'hc2bac8b2, 32'hc2056c66, 32'hc23d8d23, 32'h41ac8cb8, 32'h4262bd3c, 32'h4187d0d8};
test_weights[27352:27359] = '{32'hc198c1db, 32'hc267554d, 32'h42afa6b9, 32'hc2950b40, 32'h425eead2, 32'h428239d5, 32'h42470a17, 32'hc282c33d};
test_bias[3419:3419] = '{32'h427948ab};
test_output[3419:3419] = '{32'hc5c2df02};
test_input[27360:27367] = '{32'h4287c4ef, 32'hc2595962, 32'h3fd0b291, 32'h4200bba3, 32'hc1d5b776, 32'h42aa457f, 32'h421e7dad, 32'h41405162};
test_weights[27360:27367] = '{32'hc221fca1, 32'hc143e458, 32'h42bcc72a, 32'h42b8d302, 32'h423553a7, 32'hc208696b, 32'h42a7f7aa, 32'h4282aef4};
test_bias[3420:3420] = '{32'hc14e711c};
test_output[3420:3420] = '{32'h4480be27};
test_input[27368:27375] = '{32'h419c884d, 32'h423e062f, 32'hc2a891a9, 32'h426e8c41, 32'hc0c56d16, 32'hc261f32a, 32'h421dc428, 32'h417d6370};
test_weights[27368:27375] = '{32'h420b95b6, 32'hc254b01d, 32'h429affb8, 32'hc1a67217, 32'h42c7e04d, 32'h425a6a2a, 32'h41a9f296, 32'hc23ff28e};
test_bias[3421:3421] = '{32'h41caf1ae};
test_output[3421:3421] = '{32'hc64e76c8};
test_input[27376:27383] = '{32'h4218f775, 32'h42a39d1b, 32'hc169d8e1, 32'h42af662a, 32'h42433e5d, 32'hc2282051, 32'h4192db00, 32'h428e33c3};
test_weights[27376:27383] = '{32'h426f9ff9, 32'h41b30cfe, 32'h42c07a5a, 32'h42b55e3b, 32'hc1a53850, 32'h41d0ab86, 32'hc08a282d, 32'h42aad8e6};
test_bias[3422:3422] = '{32'h4071fe27};
test_output[3422:3422] = '{32'h46638844};
test_input[27384:27391] = '{32'hc2aa6a49, 32'hc2977dcb, 32'h41eae466, 32'h42b2de22, 32'hc2bf5e29, 32'h417147ff, 32'hc25b8e09, 32'hc0ff10bc};
test_weights[27384:27391] = '{32'hc17ba266, 32'h428c25d3, 32'h423e90c9, 32'hc26fcf82, 32'hc2bab71e, 32'h429f4aaa, 32'h4120b1dc, 32'h42563eb1};
test_bias[3423:3423] = '{32'h42863714};
test_output[3423:3423] = '{32'h44a18372};
test_input[27392:27399] = '{32'h4291241e, 32'h427b4b53, 32'h42434de9, 32'h41e0d83d, 32'h429cc1cc, 32'hc223890d, 32'h42a7ffee, 32'hc1589b8c};
test_weights[27392:27399] = '{32'h42aa73f0, 32'h4210a5af, 32'h42ac52c7, 32'hc2c77d79, 32'hc2bfeaa9, 32'h428e33f0, 32'h420b284e, 32'h42587666};
test_bias[3424:3424] = '{32'h41c81c63};
test_output[3424:3424] = '{32'h44cde080};
test_input[27400:27407] = '{32'hc2208efd, 32'hc274c7c8, 32'h416bb900, 32'h428837d8, 32'h4271e70f, 32'h421939f9, 32'h4251b0c7, 32'h418ae5fa};
test_weights[27400:27407] = '{32'hc2b6bd62, 32'h424f1fe9, 32'hc2af7a98, 32'hc0bfc5af, 32'hbfe2af94, 32'hc2106b7e, 32'h419043aa, 32'h41acc188};
test_bias[3425:3425] = '{32'hc2615e07};
test_output[3425:3425] = '{32'hc4b2879c};
test_input[27408:27415] = '{32'h4116561f, 32'hc2b07702, 32'h4128d1a5, 32'h4294d6b8, 32'h428e50df, 32'h42a2c217, 32'hc298c63a, 32'h42c42ae9};
test_weights[27408:27415] = '{32'h42706b66, 32'hc2be53f5, 32'h428c3556, 32'hc2b1005e, 32'h42151882, 32'hc123b282, 32'h42166f54, 32'h4080b489};
test_bias[3426:3426] = '{32'h426ac05b};
test_output[3426:3426] = '{32'h451d2e9a};
test_input[27416:27423] = '{32'hc0569bcb, 32'h42a595cc, 32'h4237eae7, 32'hc1cffbb1, 32'hc2c6e7b8, 32'h42ba6c20, 32'h427a820f, 32'h426cf97d};
test_weights[27416:27423] = '{32'hc230726f, 32'hc1a1f7d1, 32'h429d928d, 32'hc2866abc, 32'hc11fcf44, 32'hbfa193b4, 32'h4280a147, 32'h41bd13af};
test_bias[3427:3427] = '{32'h4286f5f9};
test_output[3427:3427] = '{32'h461f92f4};
test_input[27424:27431] = '{32'h4085bb05, 32'h424f86e6, 32'h426479da, 32'hc27f4c60, 32'hc2af770b, 32'h41c98a74, 32'hc257ae4f, 32'h40a912e0};
test_weights[27424:27431] = '{32'hc1f42413, 32'h41c4d92b, 32'h42b16e93, 32'hc002c412, 32'hc2242432, 32'hc182f52c, 32'hc235b761, 32'hc19096a9};
test_bias[3428:3428] = '{32'h42aeff0c};
test_output[3428:3428] = '{32'h463b2088};
test_input[27432:27439] = '{32'h427e8895, 32'h427911ea, 32'h424bc756, 32'hc1839ff8, 32'h41f9921e, 32'hc253109f, 32'hc29f5d9a, 32'h4179432e};
test_weights[27432:27439] = '{32'h4287e426, 32'h429ec9c4, 32'h429b4b4b, 32'h4214f6d4, 32'h41bb5f84, 32'h425310c3, 32'h41f81977, 32'h4225e046};
test_bias[3429:3429] = '{32'h429e4d99};
test_output[3429:3429] = '{32'h4609aab1};
test_input[27440:27447] = '{32'hc20d8062, 32'hc2b47520, 32'hc2c04a81, 32'h416180a1, 32'hc2224736, 32'h428c724e, 32'h4275894a, 32'h42167f7f};
test_weights[27440:27447] = '{32'hc27aa8e6, 32'hc1e73a92, 32'h42c01a2b, 32'h427ec5d1, 32'hc1f8ba28, 32'hc2829b96, 32'h42625f49, 32'h42b0e3ea};
test_bias[3430:3430] = '{32'hc18020cd};
test_output[3430:3430] = '{32'hc24d7ce3};
test_input[27448:27455] = '{32'hc2600b56, 32'h42c088d1, 32'hc1e868ee, 32'h42b1a783, 32'hc225079c, 32'h424d9eeb, 32'hc2b6d4d8, 32'hc25c4c78};
test_weights[27448:27455] = '{32'h42868df9, 32'hc2ba6f69, 32'h42408dcb, 32'hc100636b, 32'h41b31794, 32'h4242523a, 32'h416ea7d3, 32'h424c4227};
test_bias[3431:3431] = '{32'h41e3f1eb};
test_output[3431:3431] = '{32'hc688262b};
test_input[27456:27463] = '{32'hc2c3c7a8, 32'h42c0934e, 32'hc2818455, 32'hc2baca88, 32'h42051e66, 32'hc299bb4f, 32'hc214634e, 32'hc28a8458};
test_weights[27456:27463] = '{32'h42b20ec4, 32'hc190d3ea, 32'hc0bfa62a, 32'hc2c288ed, 32'hc235f988, 32'hc29fe53e, 32'hc267b5dc, 32'hc2a01db2};
test_bias[3432:3432] = '{32'hc0c3ca08};
test_output[3432:3432] = '{32'h46311312};
test_input[27464:27471] = '{32'h4204e042, 32'h3ee5c9d7, 32'hc1e0efa5, 32'h4286d13a, 32'hc181e06d, 32'hc2b116a9, 32'hc2bde859, 32'h42207ac7};
test_weights[27464:27471] = '{32'h42c22bf4, 32'hc28891f0, 32'h426f52db, 32'hc0aee637, 32'h4284b0db, 32'hc242a6b8, 32'hc1a5b881, 32'h42602f9c};
test_bias[3433:3433] = '{32'hc10620cf};
test_output[3433:3433] = '{32'h46061a98};
test_input[27472:27479] = '{32'hbdcd7972, 32'hc294feb0, 32'h4298b178, 32'h4289e15a, 32'hc1963b28, 32'hc20d236b, 32'h42555b0f, 32'hc29d903e};
test_weights[27472:27479] = '{32'hc1042c8c, 32'h3f95f1dc, 32'h42c34c45, 32'hc2977628, 32'h4282cdd5, 32'hc0dfcd48, 32'h41a1b4f3, 32'h422aafe7};
test_bias[3434:3434] = '{32'hc13d3d1e};
test_output[3434:3434] = '{32'hc48d1fb8};
test_input[27480:27487] = '{32'hc1389a0d, 32'h4241eb5f, 32'h40880e59, 32'h429a3ab0, 32'h410d0e29, 32'hbff62afd, 32'hc27396c4, 32'h41c08801};
test_weights[27480:27487] = '{32'hc22972a6, 32'h42b1dc2e, 32'hc0b8a7c5, 32'h429d273d, 32'h42ad6cce, 32'hc24a3095, 32'h427b802b, 32'h3fb7afc7};
test_bias[3435:3435] = '{32'hbf93de85};
test_output[3435:3435] = '{32'h45f6e88b};
test_input[27488:27495] = '{32'h4121fa6c, 32'h41dd4b03, 32'hc1230f22, 32'hc24e0c9a, 32'h42b22c2b, 32'hc09a1d2d, 32'hc26f00e0, 32'h4205bf73};
test_weights[27488:27495] = '{32'hc2c093cf, 32'h424356c0, 32'hc19d5ef0, 32'h42c50077, 32'h425ede51, 32'h40fc997f, 32'hc245c14b, 32'h410137aa};
test_bias[3436:3436] = '{32'hc28a002b};
test_output[3436:3436] = '{32'h455ff2e8};
test_input[27496:27503] = '{32'hc27c3245, 32'hc2ac68cd, 32'hc2610e1a, 32'h422c58ed, 32'hc292ea85, 32'h42abf946, 32'hc255d4ed, 32'h42147db5};
test_weights[27496:27503] = '{32'h4126ebff, 32'hc0e90284, 32'hc1bed2c1, 32'hc1ef810f, 32'hc203d827, 32'h41a80b7b, 32'h4253f3eb, 32'h429b1664};
test_bias[3437:3437] = '{32'hbfb414ef};
test_output[3437:3437] = '{32'h458630e4};
test_input[27504:27511] = '{32'h4250b411, 32'hc2399f6a, 32'h4278cee4, 32'hc22e37da, 32'h42ab1ac8, 32'hc2b6e806, 32'hc2c5488c, 32'hc1b49f04};
test_weights[27504:27511] = '{32'hc254aae3, 32'hc221195a, 32'hc1efe841, 32'hc1825f35, 32'h4293e781, 32'h428066f0, 32'hc24be8f0, 32'h42bb05c0};
test_bias[3438:3438] = '{32'hc2c2adc5};
test_output[3438:3438] = '{32'h4497d5fa};
test_input[27512:27519] = '{32'h4275f2f3, 32'h422ef827, 32'hc23645f7, 32'h428f555d, 32'hc2b02dbb, 32'hc22f7209, 32'h41fdced1, 32'hc2a730fe};
test_weights[27512:27519] = '{32'h42b458b2, 32'h416663fc, 32'hc23d465f, 32'h40fb6217, 32'hc2a9a830, 32'hc241a677, 32'h4270d1ac, 32'h420c42d5};
test_bias[3439:3439] = '{32'hc2a27256};
test_output[3439:3439] = '{32'h4687d61a};
test_input[27520:27527] = '{32'hc08b45f2, 32'hc17929d9, 32'hc2a2976b, 32'h42addf59, 32'hc1f45426, 32'h421ba436, 32'hc1f1b7c0, 32'h425ed0e4};
test_weights[27520:27527] = '{32'hc24c6ea7, 32'hc2a40918, 32'h42210881, 32'hc24fc613, 32'h41efb32b, 32'hc2b9cd1c, 32'hc2a4dff9, 32'h421b12d4};
test_bias[3440:3440] = '{32'h41c0d952};
test_output[3440:3440] = '{32'hc5c00288};
test_input[27528:27535] = '{32'h4282cc6b, 32'hc191c0cd, 32'h426c0c3e, 32'h4125ae83, 32'h42a29792, 32'hc1f57e6f, 32'h4274c426, 32'hc286293a};
test_weights[27528:27535] = '{32'hc2145dac, 32'h4234b7d4, 32'h4283b776, 32'h42a10560, 32'hc2a9d92f, 32'hc1d5a4bd, 32'hc2c34fe5, 32'h42b4dfd7};
test_bias[3441:3441] = '{32'hc1db8e5f};
test_output[3441:3441] = '{32'hc6825602};
test_input[27536:27543] = '{32'h40017fbc, 32'hc2c67e54, 32'h41954783, 32'hc23b42d7, 32'h4252773d, 32'h41e204e0, 32'hc294361e, 32'hc29abde7};
test_weights[27536:27543] = '{32'h40dfaabb, 32'hc24ca65b, 32'hc2a91c6f, 32'h420e77a6, 32'h42b839af, 32'h4204f453, 32'hc28ff758, 32'hc18100ed};
test_bias[3442:3442] = '{32'hc0a5b321};
test_output[3442:3442] = '{32'h465e04ad};
test_input[27544:27551] = '{32'h419a67ba, 32'hc2a94a9a, 32'h42c3bfb5, 32'hc22ce018, 32'hc1e851d7, 32'h41f221c2, 32'h429d6873, 32'h40eb0086};
test_weights[27544:27551] = '{32'h4261d0f5, 32'h411669af, 32'h41c48d1c, 32'hc2952fd4, 32'hc0f50f68, 32'h42c7fba1, 32'h408e695c, 32'hc227e8e1};
test_bias[3443:3443] = '{32'h42513bd6};
test_output[3443:3443] = '{32'h4610c5ca};
test_input[27552:27559] = '{32'hc10afc12, 32'h424382ed, 32'h4294a4d7, 32'h42a71e7c, 32'h422a7b1c, 32'h41898d3a, 32'hc2708e49, 32'hc2987a31};
test_weights[27552:27559] = '{32'hc1c7a3d8, 32'hc27bcdd9, 32'h424a55dd, 32'h41aead19, 32'h41bace07, 32'hc2bcccf9, 32'h41be79d2, 32'hc2106398};
test_bias[3444:3444] = '{32'hc04a266c};
test_output[3444:3444] = '{32'h45554e5d};
test_input[27560:27567] = '{32'h422936ff, 32'hc225c76b, 32'h424193f9, 32'h412ada11, 32'h42218121, 32'h41f997ea, 32'hc2846e92, 32'hc25489cd};
test_weights[27560:27567] = '{32'hc26ce2ab, 32'h42524682, 32'h3e4875b5, 32'hc2171230, 32'h4095dbef, 32'h4285a389, 32'h42b10baf, 32'h4277a390};
test_bias[3445:3445] = '{32'h4283f9ac};
test_output[3445:3445] = '{32'hc639c4c5};
test_input[27568:27575] = '{32'h42a62053, 32'h428a0211, 32'h415d02f1, 32'hc287067c, 32'h4234a4dc, 32'h42bfdfd1, 32'hc278d8bb, 32'h422a1b2e};
test_weights[27568:27575] = '{32'hc2b0e603, 32'h420124b0, 32'h426aee56, 32'h427c112d, 32'h42c3c843, 32'h420ff2b0, 32'h42aafe85, 32'h42be39c4};
test_bias[3446:3446] = '{32'hc1524750};
test_output[3446:3446] = '{32'hc4f70195};
test_input[27576:27583] = '{32'h41cfa796, 32'h426b9e47, 32'h42a95725, 32'h4281eb7d, 32'h4189b4d5, 32'h427d37c6, 32'hc259d784, 32'h40c900ba};
test_weights[27576:27583] = '{32'hc286eb62, 32'hc1bf88f4, 32'hc2a3d800, 32'h42448148, 32'hc2b75225, 32'hc24dddbd, 32'hc1202b2b, 32'hbfb05e63};
test_bias[3447:3447] = '{32'h42bb0627};
test_output[3447:3447] = '{32'hc62da0f0};
test_input[27584:27591] = '{32'h40efc245, 32'hc2b4b336, 32'hc126ccba, 32'h42289d4f, 32'hc28df045, 32'hc2a39136, 32'h42b06e3a, 32'hc2935190};
test_weights[27584:27591] = '{32'h42b01db3, 32'h41cdc8b0, 32'h4293dd29, 32'h411762a2, 32'h42567cbd, 32'hc1ae3413, 32'h425a9b58, 32'h41f1c446};
test_bias[3448:3448] = '{32'h42a76920};
test_output[3448:3448] = '{32'hc4acc1bd};
test_input[27592:27599] = '{32'hc1a654b4, 32'hc1e464ec, 32'h42a9445a, 32'hc26d964d, 32'h42a822eb, 32'hc1a98883, 32'h426f7ea2, 32'h42580339};
test_weights[27592:27599] = '{32'hc27675fa, 32'h42b05412, 32'h42414adb, 32'h41ce89c9, 32'hc143a57c, 32'hc1ad2c16, 32'hc23e6d1d, 32'h41bad4cd};
test_bias[3449:3449] = '{32'hc1d250bf};
test_output[3449:3449] = '{32'hc45819fe};
test_input[27600:27607] = '{32'h4283e974, 32'hc285eb13, 32'h424b1971, 32'hc141901a, 32'hc1973fff, 32'hc2835c88, 32'hbff086c0, 32'h4100c240};
test_weights[27600:27607] = '{32'hc272e632, 32'hc16665f8, 32'hc108c652, 32'hc263f92c, 32'h429e568b, 32'h42b0303f, 32'hc1122ff9, 32'hc22b7912};
test_bias[3450:3450] = '{32'h42c5e1fe};
test_output[3450:3450] = '{32'hc620e511};
test_input[27608:27615] = '{32'h42bb911e, 32'hbefc350b, 32'h41a471a4, 32'hc14ce0cf, 32'hc2a42ec2, 32'hc128860c, 32'hc09918bf, 32'h41a5140e};
test_weights[27608:27615] = '{32'h425c1f66, 32'h412dd246, 32'h42a7c4d1, 32'h4280b06a, 32'hc22e9ec7, 32'hc21e6eb9, 32'hc2ac6678, 32'h42ac8267};
test_bias[3451:3451] = '{32'h429cf9d3};
test_output[3451:3451] = '{32'h46409e63};
test_input[27616:27623] = '{32'hc28a5384, 32'hc1ef4f4f, 32'h42996eeb, 32'h420b00c4, 32'hc2a90ec2, 32'hc23e1812, 32'hc2a05e41, 32'hc21d7d8f};
test_weights[27616:27623] = '{32'h4298dfb7, 32'h412c7f28, 32'h42a237c0, 32'hc28046de, 32'h42803d6e, 32'h4276b64e, 32'hc244e274, 32'hc2bdf823};
test_bias[3452:3452] = '{32'hc292adc2};
test_output[3452:3452] = '{32'hc513182c};
test_input[27624:27631] = '{32'hc2b932bb, 32'hc18f40e0, 32'h4258da54, 32'hc245f561, 32'hc0e91f8e, 32'hc276cbe7, 32'hc2a9041c, 32'hc218255b};
test_weights[27624:27631] = '{32'h42b56d2d, 32'hc12d3507, 32'hc2522f00, 32'h423c4e67, 32'h429d45e3, 32'h429472e2, 32'hc2a77520, 32'hc23bd88c};
test_bias[3453:3453] = '{32'hc2b3ab05};
test_output[3453:3453] = '{32'hc618938a};
test_input[27632:27639] = '{32'hc191ed3b, 32'hc2794d84, 32'hc1e27108, 32'hc2adeddf, 32'h41a039ac, 32'hc261bbdb, 32'h3f37481e, 32'h428ed5f2};
test_weights[27632:27639] = '{32'h42a7e16b, 32'h42b8134a, 32'h42668538, 32'h4285ba80, 32'h428a46e8, 32'h41e0b44b, 32'hc1fbb67b, 32'hc1e5aa8e};
test_bias[3454:3454] = '{32'hbf1598ea};
test_output[3454:3454] = '{32'hc684b694};
test_input[27640:27647] = '{32'hc23e77ac, 32'h40e230f2, 32'hc2bd94b4, 32'hc2c3b20d, 32'hc22a528f, 32'h429e1fd2, 32'hc2bb5c1b, 32'hc1bd9b95};
test_weights[27640:27647] = '{32'h421ceaac, 32'hbf11527c, 32'h421e6949, 32'h42337969, 32'h42937d07, 32'h428b0100, 32'h4162ff60, 32'h42b82cdf};
test_bias[3455:3455] = '{32'hc1fde4ec};
test_output[3455:3455] = '{32'hc62f12d9};
test_input[27648:27655] = '{32'h41a89d13, 32'h42158eb3, 32'hc29ddb69, 32'hc2a74c13, 32'h426a840c, 32'hc2a2e5df, 32'h424d2e78, 32'hc23b09ae};
test_weights[27648:27655] = '{32'hc2222865, 32'h419efe2e, 32'hc2bb9e96, 32'hc13baab9, 32'hc2940b40, 32'h4291950f, 32'hc2733bb0, 32'h4244a5f5};
test_bias[3456:3456] = '{32'h419ea0ed};
test_output[3456:3456] = '{32'hc5e705a1};
test_input[27656:27663] = '{32'h428302fc, 32'hc21cdd6b, 32'hc247dc09, 32'h4210595f, 32'h40bed5f2, 32'hc2b49004, 32'h4279aea1, 32'hc248d7c6};
test_weights[27656:27663] = '{32'h42be5b82, 32'h42a9a18c, 32'hc1cd63fd, 32'h42b1ff80, 32'h4283a3db, 32'h42ac18d1, 32'hc2a977d7, 32'h42307345};
test_bias[3457:3457] = '{32'hc1c62731};
test_output[3457:3457] = '{32'hc5ea6dec};
test_input[27664:27671] = '{32'hc2b4ce89, 32'h4279afb1, 32'hc2456c74, 32'hc28cde8a, 32'hc28204f4, 32'h42845d43, 32'hc25c9a0e, 32'hc044b7ab};
test_weights[27664:27671] = '{32'h42ba8a86, 32'h41405236, 32'h4287ee8a, 32'hc24ea35b, 32'h4238cad0, 32'h425135d6, 32'h420b0991, 32'h427cb396};
test_bias[3458:3458] = '{32'hc2aa78ed};
test_output[3458:3458] = '{32'hc60ebf30};
test_input[27672:27679] = '{32'hc281d1f0, 32'h41e33e31, 32'hc28c68d6, 32'hc1fb743e, 32'hc20554ce, 32'hc2b2bcb1, 32'h410d2a9b, 32'h41c37e96};
test_weights[27672:27679] = '{32'h42a82dfd, 32'h41c8a034, 32'hc1bc6e03, 32'hc2beb3d9, 32'h4194e523, 32'h4212e27a, 32'h410facf4, 32'hc16bfbf5};
test_bias[3459:3459] = '{32'h41dd860d};
test_output[3459:3459] = '{32'hc584d70c};
test_input[27680:27687] = '{32'hc150a51c, 32'hc2920027, 32'h41f05b65, 32'hc207479e, 32'hc28f10c7, 32'hc278af2b, 32'h42742f7a, 32'hc2992585};
test_weights[27680:27687] = '{32'h410baf55, 32'hc2c75228, 32'h41b7764f, 32'hc1a7d05c, 32'hc29198c3, 32'h42a1f11b, 32'h422046a9, 32'hc1ec4aa9};
test_bias[3460:3460] = '{32'h40dd62c6};
test_output[3460:3460] = '{32'h46521fc8};
test_input[27688:27695] = '{32'hc118981e, 32'h42a37539, 32'hc28e469b, 32'hc275cc4c, 32'h41cbb1ee, 32'hc2b0b3da, 32'h4225051d, 32'h40d11df0};
test_weights[27688:27695] = '{32'hc292c042, 32'h429b45bc, 32'hc26aeefa, 32'hc2b3ffc8, 32'h4174e95f, 32'h40777af3, 32'hc1df2cba, 32'h4280879f};
test_bias[3461:3461] = '{32'hc2194519};
test_output[3461:3461] = '{32'h467a8186};
test_input[27696:27703] = '{32'h4273ac69, 32'h42b51922, 32'h41e69835, 32'hc21e2fc3, 32'hc1aae089, 32'hc2b482fd, 32'h41962e05, 32'h4290b3d4};
test_weights[27696:27703] = '{32'h429ea97a, 32'h42035cd0, 32'h42c44d8d, 32'h42bea898, 32'h42acf0c4, 32'h42b404cc, 32'h418bef69, 32'hc1b7f9c8};
test_bias[3462:3462] = '{32'h419af016};
test_output[3462:3462] = '{32'hc58a2af0};
test_input[27704:27711] = '{32'hc2321f44, 32'h42b18f8c, 32'h42a2a05e, 32'hc1ca2650, 32'hc26ed9b7, 32'hc27ae15b, 32'h41a9a669, 32'h411582f8};
test_weights[27704:27711] = '{32'h424d9070, 32'hc2c11de6, 32'hc29dd91f, 32'hc214af4a, 32'hc29006f9, 32'h4262cd2f, 32'h42056f9e, 32'h418449af};
test_bias[3463:3463] = '{32'hc2b017b0};
test_output[3463:3463] = '{32'hc6679600};
test_input[27712:27719] = '{32'h42b2f7e8, 32'hc29fde0b, 32'hc27d975a, 32'h428c21df, 32'hc2b38d1d, 32'hc2986eb5, 32'h424b2922, 32'h428fce65};
test_weights[27712:27719] = '{32'h41468ed7, 32'hbf8e4a42, 32'hc21990db, 32'h4297f99c, 32'h42705c50, 32'hc2a3e666, 32'hc2ad34d2, 32'h4208d97b};
test_bias[3464:3464] = '{32'h42abb941};
test_output[3464:3464] = '{32'h45f89fc6};
test_input[27720:27727] = '{32'hc261a237, 32'h42982db0, 32'hbfa21244, 32'h42050b49, 32'hc14ff568, 32'h42ae634f, 32'h424688e8, 32'h42ac7ea7};
test_weights[27720:27727] = '{32'h42b374dc, 32'hc1c959f9, 32'h42a48c75, 32'h426b0039, 32'hc2b6e0e6, 32'hc2a81dcc, 32'hc1fb7523, 32'h4227a289};
test_bias[3465:3465] = '{32'h423ab336};
test_output[3465:3465] = '{32'hc60f3990};
test_input[27728:27735] = '{32'hc1df5f35, 32'hc25fc7e9, 32'h41ef4ad8, 32'hc2632db0, 32'hc17fa41e, 32'h42644133, 32'h4259be02, 32'h41b52e1d};
test_weights[27728:27735] = '{32'h3f109035, 32'h424c3554, 32'hc21e188d, 32'h42652aab, 32'hc27e4ad6, 32'h41bf4107, 32'hc0b4f33f, 32'hc21ea0a9};
test_bias[3466:3466] = '{32'h42875eb8};
test_output[3466:3466] = '{32'hc5bd923e};
test_input[27736:27743] = '{32'h42aea63c, 32'h41403881, 32'hc023435f, 32'h42373efc, 32'h424aa0c8, 32'hc26f74af, 32'h42409a07, 32'h42963ada};
test_weights[27736:27743] = '{32'hc16b82e3, 32'hc2c6e182, 32'hc2550ee3, 32'hc1a8c877, 32'hc25dc85f, 32'hc2bd500c, 32'hc25aa0c0, 32'h428eb42a};
test_bias[3467:3467] = '{32'hc256bde1};
test_output[3467:3467] = '{32'h450ad43b};
test_input[27744:27751] = '{32'hc1573831, 32'h42a93113, 32'h42b1ec43, 32'h4283d1ff, 32'h421c06e5, 32'hc0847971, 32'hc2412f1c, 32'h41ba7348};
test_weights[27744:27751] = '{32'hc2c43d82, 32'hc1b53c64, 32'hc2c32c47, 32'h41d7858d, 32'hc2800c6a, 32'h428ce122, 32'h42911f2f, 32'hc28a938e};
test_bias[3468:3468] = '{32'hc101d14b};
test_output[3468:3468] = '{32'hc670eb2c};
test_input[27752:27759] = '{32'h41e982e7, 32'h42a85853, 32'h41098329, 32'h4105966f, 32'h41a9eee9, 32'h42aca678, 32'h424e473c, 32'h41edb9ed};
test_weights[27752:27759] = '{32'h41603812, 32'h426529d1, 32'h42b6dc4d, 32'h41dc865c, 32'h424e08ec, 32'hc2777d41, 32'h3feeba75, 32'h42a8c071};
test_bias[3469:3469] = '{32'h42a9deee};
test_output[3469:3469] = '{32'h459285b6};
test_input[27760:27767] = '{32'h42aceba4, 32'hc2c098c6, 32'h4270e178, 32'hc15f2147, 32'h42be4cc7, 32'hc1ba7f6e, 32'h425973c7, 32'h42290ccc};
test_weights[27760:27767] = '{32'h41f09e4e, 32'h426058d7, 32'hc29c0dcf, 32'hc1650475, 32'h401e069d, 32'hc230bb49, 32'h421fda63, 32'hc2122cb4};
test_bias[3470:3470] = '{32'h411f6811};
test_output[3470:3470] = '{32'hc5a8a60f};
test_input[27768:27775] = '{32'h422043d3, 32'hc1152237, 32'h424c54e7, 32'hc2affd27, 32'h4183b7df, 32'h40c9f16b, 32'h41d1f661, 32'h425c0d9b};
test_weights[27768:27775] = '{32'h428c0a01, 32'hc21c71df, 32'hc210650b, 32'h41a723f9, 32'h426fa712, 32'h4279f2b7, 32'hc28bb2a2, 32'h4290ce10};
test_bias[3471:3471] = '{32'hc2b45d62};
test_output[3471:3471] = '{32'h4537004e};
test_input[27776:27783] = '{32'h429d3c6f, 32'hc2ac8392, 32'h42814b0c, 32'h424be2b1, 32'hc11d7bae, 32'h404d8484, 32'hc2664a3c, 32'h425630ab};
test_weights[27776:27783] = '{32'hbe5b9940, 32'hc1aed1e7, 32'hc22fbc38, 32'h429e1734, 32'hc2b990dd, 32'hc26e44fd, 32'h42879c31, 32'h42850e46};
test_bias[3472:3472] = '{32'hc1e4e8f2};
test_output[3472:3472] = '{32'h45550fba};
test_input[27784:27791] = '{32'h4287610a, 32'h424d1a9d, 32'hc0ee86fc, 32'hc1e4abf4, 32'h42c1c5aa, 32'h3f8117d5, 32'hc17cb094, 32'h42a46863};
test_weights[27784:27791] = '{32'h42b3cce0, 32'hc28d3823, 32'h41a61cd1, 32'hc250132e, 32'hc247392d, 32'hc245c131, 32'h42a667c2, 32'h42650ed3};
test_bias[3473:3473] = '{32'h427557d2};
test_output[3473:3473] = '{32'h4514829a};
test_input[27792:27799] = '{32'hc21644e8, 32'h420c2b28, 32'h424a81d6, 32'h41c2c1c6, 32'h42a3846f, 32'hc27b9f21, 32'hc0df7b7b, 32'h423d4279};
test_weights[27792:27799] = '{32'hc285e91f, 32'h41bfe31a, 32'h4282e2e3, 32'hc106f052, 32'h42af74fe, 32'h416c9673, 32'hc0b17b08, 32'hc2242039};
test_bias[3474:3474] = '{32'h42a47f37};
test_output[3474:3474] = '{32'h462a16c2};
test_input[27800:27807] = '{32'hc2809ddd, 32'h418caa69, 32'h4212dd0a, 32'h427047ee, 32'hc22d1ba5, 32'hc204f5e6, 32'hc2b097ec, 32'h413cb65e};
test_weights[27800:27807] = '{32'h4238e6b7, 32'hc23dc01f, 32'hc111218e, 32'hc1da4dfb, 32'hc251f2fa, 32'hc13e6b84, 32'hc27cca34, 32'h429a7b51};
test_bias[3475:3475] = '{32'h423947de};
test_output[3475:3475] = '{32'h455618ab};
test_input[27808:27815] = '{32'hc229f590, 32'h4141c0df, 32'hc10afa0b, 32'hc288f7fb, 32'hc295e661, 32'hc2b626a2, 32'h428aa965, 32'h42b1ca15};
test_weights[27808:27815] = '{32'h421142ed, 32'h42391b92, 32'hc2468f5c, 32'h428abbf7, 32'hc2b54594, 32'hbf0810fd, 32'h428a185f, 32'h40d32b42};
test_bias[3476:3476] = '{32'hc1641d32};
test_output[3476:3476] = '{32'h45d7983f};
test_input[27816:27823] = '{32'h4113d46a, 32'h429e94db, 32'h42b3dc6d, 32'h4041cd21, 32'h41c74753, 32'h42186048, 32'hc2539c74, 32'h4137849e};
test_weights[27816:27823] = '{32'h42b7d386, 32'hc2ad64fc, 32'h40c015b8, 32'hc2c0e1e7, 32'hc22fcf25, 32'hc23d7648, 32'hc1ec8d80, 32'h428c12a0};
test_bias[3477:3477] = '{32'hc24b2065};
test_output[3477:3477] = '{32'hc5c6bd44};
test_input[27824:27831] = '{32'hc2785c90, 32'h42b5b15c, 32'h41e64fc3, 32'h419526eb, 32'hc2b763f5, 32'h429f73af, 32'h409fa441, 32'hc280c1a4};
test_weights[27824:27831] = '{32'hc24eeb8f, 32'h4203d42d, 32'hc2671461, 32'h42a2298b, 32'h4227ed42, 32'hbfae6c9b, 32'h423740d6, 32'h42a1821f};
test_bias[3478:3478] = '{32'hc2c4983d};
test_output[3478:3478] = '{32'hc539c307};
test_input[27832:27839] = '{32'hc2a95f80, 32'hc1980293, 32'hc29991f7, 32'hc274b1fc, 32'h42702b17, 32'h4244e7dd, 32'h42364b4a, 32'h42a128d3};
test_weights[27832:27839] = '{32'h423825c6, 32'h4298bb1b, 32'hc297d8b7, 32'hc2bf7da3, 32'h4238bb22, 32'h41b1b73f, 32'hc2749bbd, 32'h4285b4d8};
test_bias[3479:3479] = '{32'hc27271df};
test_output[3479:3479] = '{32'h46471c4d};
test_input[27840:27847] = '{32'h422f7848, 32'hc2912289, 32'hc2b9bebd, 32'hc2840536, 32'h3f4ca0ef, 32'hc1f99e2e, 32'h42a4d14a, 32'hc276cf72};
test_weights[27840:27847] = '{32'hc103002e, 32'hc26c01c2, 32'h421cf4c4, 32'hc264d223, 32'h42c08057, 32'hc214cd25, 32'hc212d1d5, 32'h41743a6c};
test_bias[3480:3480] = '{32'h41c341cd};
test_output[3480:3480] = '{32'h44a8b858};
test_input[27848:27855] = '{32'hc2bec4f7, 32'h422b0837, 32'hc25c510a, 32'h41505973, 32'hc105b561, 32'hc1ac026d, 32'h427fd215, 32'hc2410609};
test_weights[27848:27855] = '{32'hc2afb868, 32'h42823b21, 32'hc27ab64c, 32'h4222dd55, 32'hc2647b56, 32'h409ecd73, 32'hc19a9f96, 32'hc2c742de};
test_bias[3481:3481] = '{32'hc29fc44b};
test_output[3481:3481] = '{32'h46948328};
test_input[27856:27863] = '{32'h427e0cc1, 32'hc0ef6289, 32'h42b8aa36, 32'hc20039ac, 32'h4280bba2, 32'hc2111060, 32'h42bb1297, 32'hc28b95f6};
test_weights[27856:27863] = '{32'h42b92c4c, 32'h42aa8f7e, 32'hc1ccb1ea, 32'hc293da65, 32'h42391314, 32'h429d4b5c, 32'hc24a6be7, 32'h42b33845};
test_bias[3482:3482] = '{32'h41b86f28};
test_output[3482:3482] = '{32'hc5aea6b9};
test_input[27864:27871] = '{32'h41d46b77, 32'hc286ee7e, 32'hc2487a86, 32'hc179d415, 32'hc00d8979, 32'h42af6a9e, 32'hc2b4c2d7, 32'hc15cf5f0};
test_weights[27864:27871] = '{32'hc27faef8, 32'h42152a31, 32'hc22c734c, 32'h42751703, 32'hc2644f1c, 32'hc018e8ba, 32'hc2954b7c, 32'h3f015a76};
test_bias[3483:3483] = '{32'hc1adc354};
test_output[3483:3483] = '{32'h45629938};
test_input[27872:27879] = '{32'h420c73d3, 32'hc194cc69, 32'hc2b168af, 32'hc205c3d6, 32'hc281ab5d, 32'hc24c7d5b, 32'h4203e467, 32'hc2064b17};
test_weights[27872:27879] = '{32'h427d7425, 32'h41acf549, 32'hc2914a73, 32'hc22b48f0, 32'h418624d2, 32'h422fd83b, 32'hc22e9f14, 32'h421af5e8};
test_bias[3484:3484] = '{32'hc16dddda};
test_output[3484:3484] = '{32'h456193b1};
test_input[27880:27887] = '{32'h42c6debc, 32'hc2a7db44, 32'h429450e1, 32'hc1567000, 32'hc23ac316, 32'h42b6dd30, 32'hbffd7e4e, 32'h42426d72};
test_weights[27880:27887] = '{32'h4240a9d5, 32'h418f442c, 32'h4244301b, 32'h4248e454, 32'hc28eaf99, 32'hc183d4f8, 32'h428d1570, 32'hc25b6e38};
test_bias[3485:3485] = '{32'h42b1df4b};
test_output[3485:3485] = '{32'h45a76cb4};
test_input[27888:27895] = '{32'hc1bce62d, 32'h428ee83e, 32'h424c96fc, 32'hc2abc6d0, 32'h40a88bb1, 32'hc25d520e, 32'hc1870f32, 32'h412970c5};
test_weights[27888:27895] = '{32'hc24cea14, 32'h42c26737, 32'hc2629cee, 32'hc1b3a4f1, 32'hc1a89f15, 32'hc1c17af8, 32'hc19f4449, 32'h423aa85b};
test_bias[3486:3486] = '{32'hc29d8cfc};
test_output[3486:3486] = '{32'h460f32b7};
test_input[27896:27903] = '{32'h4126ab37, 32'hc29c59cc, 32'h4219eb89, 32'h429b6541, 32'h3fd908a2, 32'h426327bc, 32'hc26862ee, 32'hc22e6fde};
test_weights[27896:27903] = '{32'h4274f45a, 32'hc25b7ad2, 32'h41b5dd8c, 32'h424bde41, 32'hc286211e, 32'h42c65f99, 32'h42c78e49, 32'hc07a83c7};
test_bias[3487:3487] = '{32'hc2849c7a};
test_output[3487:3487] = '{32'h4615d338};
test_input[27904:27911] = '{32'h422b2ee2, 32'hc1e4664c, 32'h41a16d19, 32'hc1840507, 32'hc20a5c1d, 32'h42b27ec6, 32'hc1b7a4c6, 32'h41ffecc2};
test_weights[27904:27911] = '{32'h41da5a21, 32'h42b22827, 32'h4160ff3f, 32'hc2843e01, 32'h41676412, 32'hc2b405ca, 32'h42afac75, 32'h429b20c2};
test_bias[3488:3488] = '{32'hc29c2460};
test_output[3488:3488] = '{32'hc5fe9690};
test_input[27912:27919] = '{32'h424ddc37, 32'hc26a9df9, 32'hc2a92e7e, 32'h41a65043, 32'h4254a2d3, 32'hc2c05197, 32'hc05497f6, 32'h417b11b7};
test_weights[27912:27919] = '{32'hc1384ee4, 32'h413b0ec0, 32'h42c34984, 32'hc1dc0a16, 32'h41345d69, 32'hc1379aae, 32'hc294bdda, 32'h42b1727a};
test_bias[3489:3489] = '{32'h42204f6a};
test_output[3489:3489] = '{32'hc5d24087};
test_input[27920:27927] = '{32'h429bd144, 32'h42bbb020, 32'hc20fecb5, 32'h423894c0, 32'hc2694cf7, 32'h4241fd4d, 32'h41ea1d99, 32'h42aa5204};
test_weights[27920:27927] = '{32'h41ace562, 32'h42a9458e, 32'h42a715af, 32'hc20a5f8f, 32'h41b9982b, 32'hc2ae1d8d, 32'hc2aec400, 32'h42243cba};
test_bias[3490:3490] = '{32'h42bae447};
test_output[3490:3490] = '{32'h43f0df02};
test_input[27928:27935] = '{32'hc1010cd2, 32'hc10ccc0f, 32'h4214528b, 32'h403dce13, 32'h41c46809, 32'hc2c7974c, 32'hc25577d2, 32'h42af8458};
test_weights[27928:27935] = '{32'h42729ac2, 32'hc1e27d04, 32'h4280b6d7, 32'hc228ee90, 32'hc2621226, 32'hc0c566b8, 32'hc0217362, 32'hc2b3079e};
test_bias[3491:3491] = '{32'h40dae697};
test_output[3491:3491] = '{32'hc5ca0889};
test_input[27936:27943] = '{32'h42c0ee4f, 32'h4295b872, 32'h41a16369, 32'h41713187, 32'h42c0829b, 32'h42aacc9a, 32'h42457406, 32'hc2abfe2f};
test_weights[27936:27943] = '{32'h42ab3620, 32'hc200621d, 32'hc22be5af, 32'hc07d4609, 32'h429c2c71, 32'h4185b81c, 32'hc2b3c927, 32'h42361575};
test_bias[3492:3492] = '{32'hc1f0c68a};
test_output[3492:3492] = '{32'h45ab91f3};
test_input[27944:27951] = '{32'h42467287, 32'hc1ee771f, 32'h4228a780, 32'hc200b53c, 32'h4245ca52, 32'hc225f457, 32'h42b132cd, 32'h426d8886};
test_weights[27944:27951] = '{32'hc1db8646, 32'hc224e38c, 32'h418c336b, 32'hc2490ed5, 32'h429232f8, 32'h42acf439, 32'h429e57db, 32'hc241862f};
test_bias[3493:3493] = '{32'hc2165cca};
test_output[3493:3493] = '{32'h45c692f9};
test_input[27952:27959] = '{32'h421f29b8, 32'hc0e88ce8, 32'h42875834, 32'h428ff37c, 32'h4239ed3f, 32'h413c1903, 32'hc2c68b04, 32'h429270ec};
test_weights[27952:27959] = '{32'hc28fdca2, 32'h41d2a215, 32'h42237bfb, 32'h422c9b4a, 32'h42a8d65b, 32'h4283bd97, 32'h42960e71, 32'h42a698cc};
test_bias[3494:3494] = '{32'h419a0ea5};
test_output[3494:3494] = '{32'h45c155d5};
test_input[27960:27967] = '{32'h419b5f42, 32'hc22524af, 32'hc2752544, 32'h42876297, 32'hc174f11a, 32'h42b3ce12, 32'hc274a38f, 32'h424c0008};
test_weights[27960:27967] = '{32'hc051945e, 32'h42b75123, 32'h42ab0910, 32'hc27fa9c8, 32'h4240d778, 32'hc2a60da7, 32'h4280f815, 32'hc25a3901};
test_bias[3495:3495] = '{32'hc2b4b1c7};
test_output[3495:3495] = '{32'hc6de24c5};
test_input[27968:27975] = '{32'hc17fdc51, 32'h42b4e954, 32'hc2849824, 32'h4234891f, 32'h4216e265, 32'hc0dae4e5, 32'hc14a886c, 32'hc2339fcc};
test_weights[27968:27975] = '{32'hc2c2aa42, 32'hc212c088, 32'hc1a7e8e3, 32'hc2941882, 32'hc2705e42, 32'hc22c8d09, 32'hc272bbc7, 32'h423224ff};
test_bias[3496:3496] = '{32'h4209a8df};
test_output[3496:3496] = '{32'hc5d70e3e};
test_input[27976:27983] = '{32'h42861fe9, 32'h429ad074, 32'h42aa6bd2, 32'hc2bf4703, 32'hc28830b8, 32'h42b5ecd9, 32'h42424021, 32'h40dacbc2};
test_weights[27976:27983] = '{32'h42134b0e, 32'h41c89393, 32'h42c324ec, 32'hc284309b, 32'hc181a1e0, 32'h42a05012, 32'h42af67c2, 32'h42b15d3f};
test_bias[3497:3497] = '{32'h41e35f64};
test_output[3497:3497] = '{32'h46fc9c3c};
test_input[27984:27991] = '{32'hc158907c, 32'hc2564e08, 32'hc2aab25a, 32'h425efa0e, 32'hc1eda26b, 32'hc23aefe7, 32'h42ad7ec6, 32'hc276abd5};
test_weights[27984:27991] = '{32'hc1979a43, 32'h42407307, 32'hc291860c, 32'h420ece2e, 32'hc2a35f56, 32'hc21b552d, 32'h42bd8444, 32'h429c0509};
test_bias[3498:3498] = '{32'h429100bc};
test_output[3498:3498] = '{32'h465488ce};
test_input[27992:27999] = '{32'h42256963, 32'hc2413d42, 32'hc2c20caf, 32'hc29ac741, 32'h41c40292, 32'h42963aae, 32'h423d8596, 32'h429889cf};
test_weights[27992:27999] = '{32'hc20bdf47, 32'h40abec69, 32'h422a8cbf, 32'h42775a20, 32'h428e93f0, 32'h414cf808, 32'hc2c01247, 32'hc1c7e176};
test_bias[3499:3499] = '{32'hc225baf4};
test_output[3499:3499] = '{32'hc661417d};
test_input[28000:28007] = '{32'h40805ed6, 32'hc2254d55, 32'h42556e4d, 32'hc0c2938d, 32'hc2c15986, 32'hc29b9e18, 32'h3fb7b7b6, 32'hc16049ce};
test_weights[28000:28007] = '{32'h42342367, 32'h41a1da37, 32'hc26a498e, 32'h42ae49a9, 32'hc0e68147, 32'hc1b842a2, 32'h41f2b1ab, 32'hc283c045};
test_bias[3500:3500] = '{32'hc2b1f952};
test_output[3500:3500] = '{32'hc46c0324};
test_input[28008:28015] = '{32'hc1ae7bde, 32'hc235aa49, 32'h42c0bc3d, 32'h426da40d, 32'h40d44985, 32'hc2be301d, 32'h42bbac8c, 32'hc2bb5976};
test_weights[28008:28015] = '{32'hc22c4485, 32'hc20da498, 32'hc299523b, 32'hc27b31fa, 32'h40f36cdb, 32'h42775e72, 32'hc28459ca, 32'hc23ec1fe};
test_bias[3501:3501] = '{32'hc2891d93};
test_output[3501:3501] = '{32'hc67d511c};
test_input[28016:28023] = '{32'hc28fc624, 32'hc2086266, 32'hc1d7b39d, 32'hc1a2fcf2, 32'hc2623fac, 32'hc27b3287, 32'h41c558e7, 32'h42963831};
test_weights[28016:28023] = '{32'h40ae4404, 32'h420690c8, 32'hc2a4e663, 32'hc02478e7, 32'hc20e5280, 32'h40e05b52, 32'hc25225e4, 32'hc1a73dd6};
test_bias[3502:3502] = '{32'hc1d493c8};
test_output[3502:3502] = '{32'hc411e871};
test_input[28024:28031] = '{32'h429c308f, 32'hc280db89, 32'h4284afcd, 32'hc1f1b149, 32'hc19bda8b, 32'hc2c18c32, 32'hc223afcb, 32'h42a25f30};
test_weights[28024:28031] = '{32'h4216cb7c, 32'hc24514d1, 32'hc231c550, 32'hc1a05e45, 32'h41b95241, 32'hc2ab47d4, 32'hc295f872, 32'h41f97938};
test_bias[3503:3503] = '{32'hc18a9a05};
test_output[3503:3503] = '{32'h46865601};
test_input[28032:28039] = '{32'h428631be, 32'hc2af9218, 32'h425ce05f, 32'h427cd224, 32'h41c2e5c8, 32'hc239070a, 32'h40e18631, 32'h42819af8};
test_weights[28032:28039] = '{32'hc1faff66, 32'hc29da60b, 32'h4126c100, 32'h41a1f447, 32'h40271a9a, 32'h42639553, 32'h41a14e97, 32'hc292149f};
test_bias[3504:3504] = '{32'hc2b8f038};
test_output[3504:3504] = '{32'hc4119193};
test_input[28040:28047] = '{32'hc236ce57, 32'hc2aec102, 32'hc2963724, 32'hc1eb6388, 32'hc2c6a52c, 32'h3f9aaec8, 32'h42a862fe, 32'h407429df};
test_weights[28040:28047] = '{32'h42bb25e3, 32'hc2a3e971, 32'hc1d1f374, 32'h42b8cd82, 32'h422eac0a, 32'h418a9837, 32'h428dc039, 32'hc203f5c9};
test_bias[3505:3505] = '{32'h421d490c};
test_output[3505:3505] = '{32'h4567557c};
test_input[28048:28055] = '{32'h41dcdff7, 32'hc29c7325, 32'hc29c83dd, 32'h40d8c060, 32'h4270dd69, 32'hc26e0075, 32'hc20eb66e, 32'hc1beb88b};
test_weights[28048:28055] = '{32'hc23627c5, 32'hc1b03f77, 32'h42626ac0, 32'hc2bcd5cb, 32'h4236bafc, 32'h42644fca, 32'hc2c0ee1f, 32'hc263e704};
test_bias[3506:3506] = '{32'h4266ef32};
test_output[3506:3506] = '{32'hc3c36202};
test_input[28056:28063] = '{32'h42c1d583, 32'h42b04a01, 32'h42ba142d, 32'h42381cde, 32'hc2951e0a, 32'h42b6a6a6, 32'h423c3081, 32'hc158690d};
test_weights[28056:28063] = '{32'h42b70489, 32'h42624279, 32'h42697313, 32'h41f7ca82, 32'h3f847f59, 32'h41cf1506, 32'h42222392, 32'hc26adb7e};
test_bias[3507:3507] = '{32'h42a14e96};
test_output[3507:3507] = '{32'h46c965fa};
test_input[28064:28071] = '{32'h42a7525d, 32'hc2afc0ec, 32'hc239b2fe, 32'h428bc909, 32'h428ebe66, 32'hc21a8e15, 32'h42a6e8e9, 32'h40e4a838};
test_weights[28064:28071] = '{32'hc1f6a61e, 32'h41f556d1, 32'hc2c39010, 32'hc18ca561, 32'hc2c228bd, 32'hc2b86c7b, 32'hc289b39f, 32'hc2107d67};
test_bias[3508:3508] = '{32'hc23b6911};
test_output[3508:3508] = '{32'hc631d132};
test_input[28072:28079] = '{32'hc2ac274a, 32'hc263f2f3, 32'h414ef379, 32'hc1cddf5a, 32'h421bbbaf, 32'h4283a2d8, 32'hc2129047, 32'h42b9a59a};
test_weights[28072:28079] = '{32'h4287586b, 32'h41971fb5, 32'h41c61bc3, 32'hc2b30c82, 32'h42a9f142, 32'h42909fe4, 32'h4225b2d0, 32'hc2278e08};
test_bias[3509:3509] = '{32'h42b2540a};
test_output[3509:3509] = '{32'hc4bed62c};
test_input[28080:28087] = '{32'hc2302182, 32'hc10f6591, 32'h4205142f, 32'h4176e404, 32'hc18006a6, 32'hc2c47230, 32'hc2b207e5, 32'hc2041912};
test_weights[28080:28087] = '{32'h41cb1c42, 32'h42c0dc28, 32'hc15225a0, 32'h42321643, 32'h41482dca, 32'h42102b9f, 32'hc21227af, 32'hc2044fbf};
test_bias[3510:3510] = '{32'hc201ee2f};
test_output[3510:3510] = '{32'hc4910549};
test_input[28088:28095] = '{32'hc28e2210, 32'hc2843b0e, 32'hc29ab933, 32'h42b4c067, 32'h413e96ff, 32'hc27e83fd, 32'h42aa70e5, 32'hc196e5f0};
test_weights[28088:28095] = '{32'h420368e9, 32'h421100fa, 32'h41ebe25a, 32'hc2a1a3ac, 32'hc282feda, 32'h42b2360e, 32'hc1b6d67c, 32'h4200bf8b};
test_bias[3511:3511] = '{32'h4263202d};
test_output[3511:3511] = '{32'hc6b5c122};
test_input[28096:28103] = '{32'hc1b2d08b, 32'h42444248, 32'hc2a78dc1, 32'h429b3999, 32'hc2be2f0f, 32'h41f9b523, 32'h428ab1ac, 32'h421a1f5d};
test_weights[28096:28103] = '{32'h42b49b3c, 32'h412aa99c, 32'hc23f1d25, 32'h42be08bb, 32'hc183201e, 32'hc25d180f, 32'h401187bb, 32'h420fc181};
test_bias[3512:3512] = '{32'hc29c9b55};
test_output[3512:3512] = '{32'h462eae80};
test_input[28104:28111] = '{32'hc2394756, 32'hc20925f6, 32'h428276a5, 32'h3fd7cf49, 32'hc2486a0e, 32'h429babbd, 32'hc2869416, 32'hc2a6e172};
test_weights[28104:28111] = '{32'h420651d6, 32'hc096dee0, 32'h429b3594, 32'hc1d4530e, 32'hc25c0ccb, 32'hc2132619, 32'h4232208c, 32'h4291eb64};
test_bias[3513:3513] = '{32'hc2858920};
test_output[3513:3513] = '{32'hc5b01275};
test_input[28112:28119] = '{32'h41d0d5f8, 32'h420d4f0c, 32'hc2810ce3, 32'hc274f837, 32'hc1ed64ce, 32'hc2b5de8b, 32'h41dc436f, 32'hc2bb8a5a};
test_weights[28112:28119] = '{32'h41f103ca, 32'h4207ad92, 32'h411fb438, 32'h41e721d1, 32'h420ca903, 32'hc1b0d006, 32'h42151e18, 32'h4237eb85};
test_bias[3514:3514] = '{32'h41f52199};
test_output[3514:3514] = '{32'hc529cea7};
test_input[28120:28127] = '{32'hc196c27f, 32'h3f87dbc7, 32'hc264bcbd, 32'hc2c69775, 32'h42883acb, 32'h4273014c, 32'hc296dd88, 32'h42b19876};
test_weights[28120:28127] = '{32'h423687df, 32'h3f3e0ad1, 32'hc239b172, 32'h42b7ad13, 32'h420a0ad2, 32'h424393d1, 32'h424c5a58, 32'hc2af858e};
test_bias[3515:3515] = '{32'h42133e15};
test_output[3515:3515] = '{32'hc654b1a5};
test_input[28128:28135] = '{32'hc2941172, 32'h421f6e52, 32'hc2a579a5, 32'hc132ee69, 32'hc26eae11, 32'h42a2df89, 32'hc282aaf9, 32'h42a1421c};
test_weights[28128:28135] = '{32'h42b2aada, 32'h4127034f, 32'h41f66f31, 32'hc1938c87, 32'h423fd838, 32'h42bcda3c, 32'hc2405f76, 32'h423ee5ce};
test_bias[3516:3516] = '{32'hc2a4ed9d};
test_output[3516:3516] = '{32'h4547b705};
test_input[28136:28143] = '{32'hc1837edf, 32'h42b80ae6, 32'h428cac92, 32'h42519767, 32'h4212368f, 32'h41c0f949, 32'hc2ab30ea, 32'hc2a07454};
test_weights[28136:28143] = '{32'hc2696d54, 32'hc22ecde6, 32'hc288419a, 32'h414a2534, 32'hc27f86d4, 32'h4205f427, 32'hc1caf6fe, 32'hc2756ddc};
test_bias[3517:3517] = '{32'hc2a57b14};
test_output[3517:3517] = '{32'hc4d58182};
test_input[28144:28151] = '{32'hc2c6e67a, 32'hc0f12f3e, 32'h41b790fc, 32'h41e96757, 32'h4292548c, 32'h4235e1aa, 32'h41c212e4, 32'hc2a2d967};
test_weights[28144:28151] = '{32'hc2902c0f, 32'hc29dab4c, 32'hc1c37083, 32'h41adda80, 32'h3f98d794, 32'hc18b9518, 32'hc2c71fa2, 32'hbf5e8ff6};
test_bias[3518:3518] = '{32'h42905731};
test_output[3518:3518] = '{32'h4597d24f};
test_input[28152:28159] = '{32'hc2055491, 32'hc1523940, 32'h426fe45a, 32'hc25905d5, 32'hc2a81cd4, 32'hc2ad8c0c, 32'h41b53b8a, 32'h41960d52};
test_weights[28152:28159] = '{32'hc2c225f5, 32'h42983e41, 32'hc2899945, 32'hbfe5776d, 32'h41c9e423, 32'hc2b5abea, 32'h4224f9ed, 32'h42c77837};
test_bias[3519:3519] = '{32'h42c22915};
test_output[3519:3519] = '{32'h45d6ad94};
test_input[28160:28167] = '{32'h429396ad, 32'hc2455724, 32'hc1308d8d, 32'hc2a04554, 32'h42c6d6b8, 32'h41d6885e, 32'hc2856653, 32'hc2b1ceba};
test_weights[28160:28167] = '{32'hc23f4413, 32'hc2b8f06b, 32'hc0c9b82a, 32'h42acbaba, 32'h42a900d5, 32'hc2c6244e, 32'h4113d564, 32'hc2812624};
test_bias[3520:3520] = '{32'hc24fcd74};
test_output[3520:3520] = '{32'h459c391f};
test_input[28168:28175] = '{32'hc27be745, 32'h42c0d5af, 32'h42b4ef79, 32'hc21bed29, 32'hc2235524, 32'h425edbc7, 32'h429a53d4, 32'h425c5db9};
test_weights[28168:28175] = '{32'hc20cbcca, 32'hc2af8951, 32'hc26d8571, 32'hc2529e4e, 32'hc2a5c15b, 32'h42b87e74, 32'hc23e2d1f, 32'h41b2b2e2};
test_bias[3521:3521] = '{32'h40bbbc8a};
test_output[3521:3521] = '{32'hc55929ac};
test_input[28176:28183] = '{32'h41a37290, 32'hc222adef, 32'h42362f1c, 32'h428e6bd3, 32'h428b11db, 32'h4277eb0a, 32'h4292ca51, 32'hbff60659};
test_weights[28176:28183] = '{32'h42afdeb5, 32'h42248fab, 32'h41d557c5, 32'hc27f1b7a, 32'hc12164be, 32'h410a28c0, 32'h427a632a, 32'h4038cb46};
test_bias[3522:3522] = '{32'h42253ab4};
test_output[3522:3522] = '{32'h449d8993};
test_input[28184:28191] = '{32'hc1cb2912, 32'hc2ac8ac1, 32'h41d57c23, 32'hc192845a, 32'hc18dca1c, 32'hc14c0f3f, 32'h42b6973f, 32'h41b24272};
test_weights[28184:28191] = '{32'h42780d0b, 32'h41650a47, 32'hc1781c2b, 32'hc193ac03, 32'h4263de67, 32'h42a56436, 32'h42702d22, 32'h4189f540};
test_bias[3523:3523] = '{32'h41bbeb13};
test_output[3523:3523] = '{32'h446ae78e};
test_input[28192:28199] = '{32'hc1374adb, 32'hc2a37861, 32'h423d967c, 32'h3f64c699, 32'h42088aaa, 32'h41612f6a, 32'hc253487f, 32'h426a62bc};
test_weights[28192:28199] = '{32'hc2bd54a0, 32'h4269b2b5, 32'h4296ea32, 32'hc1062d21, 32'h4245fea5, 32'h41b3d5ff, 32'h42995987, 32'h426b91c8};
test_bias[3524:3524] = '{32'h422a08a1};
test_output[3524:3524] = '{32'h44a5ef8c};
test_input[28200:28207] = '{32'hc2bcc976, 32'hc2b92f6a, 32'hc1451789, 32'h42280961, 32'h4284d3c6, 32'hc2c17d73, 32'h42992c9d, 32'h4204f1bc};
test_weights[28200:28207] = '{32'h41f5bbf3, 32'h41cff12b, 32'hc1f4b478, 32'h42021cea, 32'hc0d050fc, 32'h41d3afbd, 32'h42008d9a, 32'h4249df5b};
test_bias[3525:3525] = '{32'h422d4d74};
test_output[3525:3525] = '{32'hc5145278};
test_input[28208:28215] = '{32'hc22f10a6, 32'h4155de9f, 32'h42b8b3bd, 32'hc28eefb5, 32'hc2493b23, 32'hc1f09e08, 32'hc191f26a, 32'hc1a5922f};
test_weights[28208:28215] = '{32'hc26d6c61, 32'h42925754, 32'h42674ffa, 32'h42ad8659, 32'h422e31b6, 32'hc0f4772e, 32'h4211d145, 32'h42909bcb};
test_bias[3526:3526] = '{32'hc1bcd317};
test_output[3526:3526] = '{32'hc4b2d218};
test_input[28216:28223] = '{32'hc191a180, 32'hc2a38e93, 32'h41eb282a, 32'h4254aa20, 32'hc2b92841, 32'hc29e26ee, 32'h422297c2, 32'hc29333d9};
test_weights[28216:28223] = '{32'hc2b3149a, 32'hc2bfc4d2, 32'h42024e47, 32'hc2b5c127, 32'hc1bf4d0f, 32'hc2a25475, 32'hc26faa12, 32'hc1668806};
test_bias[3527:3527] = '{32'hc179a3fb};
test_output[3527:3527] = '{32'h46489a78};
test_input[28224:28231] = '{32'hc247e640, 32'h42983cb2, 32'hc2893938, 32'h410f93cc, 32'h419b6bf5, 32'h42c0d56d, 32'h41ca0bff, 32'hc189d407};
test_weights[28224:28231] = '{32'hc103d91d, 32'h4200bfe2, 32'hc2b290bb, 32'h419a7cb7, 32'hc2a69509, 32'h4291e350, 32'h41817363, 32'h41c196e2};
test_bias[3528:3528] = '{32'hc055bb08};
test_output[3528:3528] = '{32'h46639136};
test_input[28232:28239] = '{32'hc1c14dac, 32'hc12965c9, 32'hc257eea1, 32'h41f186f4, 32'hc292c441, 32'h427d7e00, 32'hc2c0c516, 32'hc1d3bcee};
test_weights[28232:28239] = '{32'h428ea34f, 32'hc294afaf, 32'hc2af586b, 32'hc26e5b02, 32'hc29fa01e, 32'h42ae6640, 32'h42a326dd, 32'hc1aa583e};
test_bias[3529:3529] = '{32'hc220aafa};
test_output[3529:3529] = '{32'h45bccaee};
test_input[28240:28247] = '{32'h40efaf15, 32'hc152ee3b, 32'h42a5facd, 32'h41c9fea0, 32'hc1b3a198, 32'h4295661c, 32'hc1cbfe9e, 32'hc21490c2};
test_weights[28240:28247] = '{32'h428d1e1e, 32'hc2878bc5, 32'h4277cf68, 32'h4289cb80, 32'hc1c6d63b, 32'h427c3d62, 32'h42b905a0, 32'h41ed303f};
test_bias[3530:3530] = '{32'h417e6184};
test_output[3530:3530] = '{32'h461e3d7c};
test_input[28248:28255] = '{32'h423b65d2, 32'h42a22aa0, 32'hc2270d13, 32'hc25315d2, 32'hc21d19ed, 32'hc1d7f3b4, 32'h41a174e7, 32'hc22785d3};
test_weights[28248:28255] = '{32'hc28a579c, 32'hc2ab9dda, 32'h423ebcb8, 32'hc2b808db, 32'hc0852892, 32'hc2b8b7f7, 32'hc19c9d3c, 32'hc2a80b5a};
test_bias[3531:3531] = '{32'h428e7e7b};
test_output[3531:3531] = '{32'hc4b94550};
test_input[28256:28263] = '{32'h41cfbdc1, 32'hc2561db4, 32'h42166d2e, 32'hc2862584, 32'hc16660bb, 32'h421be750, 32'h41b44639, 32'hc2ad4ce6};
test_weights[28256:28263] = '{32'h412a7895, 32'h427add51, 32'h42111fba, 32'hc2a8d789, 32'h42855a90, 32'hc276023a, 32'h428fef50, 32'hc298ec76};
test_bias[3532:3532] = '{32'hc2b0bdc6};
test_output[3532:3532] = '{32'h4608afe6};
test_input[28264:28271] = '{32'h429fbaf9, 32'h42b9f0bd, 32'h423b65d1, 32'hc1a22deb, 32'h4253bc1c, 32'hc2127368, 32'h4241c6fd, 32'h416524e6};
test_weights[28264:28271] = '{32'hc2bcbba3, 32'hc18db787, 32'hc29612b9, 32'hc2be77a0, 32'hc1e236f5, 32'h42bb4656, 32'h4216e36c, 32'h41949286};
test_bias[3533:3533] = '{32'hc20dd8ef};
test_output[3533:3533] = '{32'hc6550e0e};
test_input[28272:28279] = '{32'hc2bdf995, 32'h42213267, 32'hc21bf244, 32'h40207877, 32'hc1cc5108, 32'h423156e3, 32'h426054c0, 32'h41756153};
test_weights[28272:28279] = '{32'h4248b6c3, 32'h422dcc2e, 32'hc1fae523, 32'h426eaae1, 32'h426fe6e1, 32'h426b0c5a, 32'h40eedd92, 32'hc25f08ce};
test_bias[3534:3534] = '{32'hc2a47c7c};
test_output[3534:3534] = '{32'hc4880a91};
test_input[28280:28287] = '{32'h42c5b8d4, 32'hc2a3b0f8, 32'hc1b507a5, 32'h423d34b5, 32'hc287a7e9, 32'h42369bdd, 32'h42ba439f, 32'hc1ac94fb};
test_weights[28280:28287] = '{32'hc24792cf, 32'h4243b0e5, 32'h42b9e92a, 32'hc1cebc15, 32'hc18283ed, 32'h4230c1f9, 32'h423585ad, 32'h4278a515};
test_bias[3535:3535] = '{32'h41245118};
test_output[3535:3535] = '{32'hc5c316db};
test_input[28288:28295] = '{32'h429ade86, 32'hc1e1f22e, 32'hc252c058, 32'hc28e9f36, 32'h42c04c17, 32'h42597822, 32'hc215df5c, 32'h42915767};
test_weights[28288:28295] = '{32'h42beee38, 32'h416938e6, 32'hc18e90a7, 32'hc2c57825, 32'h42b4919a, 32'hc20b74e0, 32'hc2970a9e, 32'h3ff4df05};
test_bias[3536:3536] = '{32'hc27fcdf0};
test_output[3536:3536] = '{32'h46c094bc};
test_input[28296:28303] = '{32'h42a1c96d, 32'hc2aec5cb, 32'h41a3a924, 32'hc28c8cca, 32'h42bc0220, 32'h4289b6a2, 32'h40cd6edb, 32'hc2755fef};
test_weights[28296:28303] = '{32'h42222222, 32'hc12f0c38, 32'hc221d15a, 32'h423f0ffe, 32'hc19aca79, 32'h41827f14, 32'hc1be2325, 32'hc1fa331b};
test_bias[3537:3537] = '{32'hc284ee43};
test_output[3537:3537] = '{32'h4483ccad};
test_input[28304:28311] = '{32'h42ac51c3, 32'h42861400, 32'hc2b017fb, 32'h3f6b773a, 32'h4200889b, 32'hc2460c6f, 32'h42268cb2, 32'h41f8acc7};
test_weights[28304:28311] = '{32'h420a1ac8, 32'hc2bd65f9, 32'hc2acda01, 32'hc29bcdc5, 32'h42a96feb, 32'h4259e13b, 32'hc167dc56, 32'h42c008e1};
test_bias[3538:3538] = '{32'h41dc26d3};
test_output[3538:3538] = '{32'h45ce31dd};
test_input[28312:28319] = '{32'h41e1b6f9, 32'h41c93947, 32'h420168b4, 32'h41cf0f77, 32'hc2ae1d8d, 32'hc2bb5966, 32'h428b5372, 32'hc211cde2};
test_weights[28312:28319] = '{32'hc22abc7b, 32'hc218eedf, 32'h41305ca0, 32'h42b8356a, 32'hc28154c7, 32'hc1b138fd, 32'hc2b9ff99, 32'hc19837e8};
test_bias[3539:3539] = '{32'hc1026f19};
test_output[3539:3539] = '{32'h451b61fb};
test_input[28320:28327] = '{32'h425f6d61, 32'hc23c1f87, 32'hc24e65d1, 32'h42705842, 32'hc2c460a4, 32'hc296edfb, 32'h4281902a, 32'h42777413};
test_weights[28320:28327] = '{32'h41d08b28, 32'h41d9c5ef, 32'h42aea503, 32'hc2657ce7, 32'hc19aa59d, 32'h421379d8, 32'h42919928, 32'h421c013e};
test_bias[3540:3540] = '{32'h42432d10};
test_output[3540:3540] = '{32'hc4b97c3b};
test_input[28328:28335] = '{32'hc2b8f06c, 32'hc28058ca, 32'hc2a03be4, 32'hc145d585, 32'hc251ae42, 32'hc2632246, 32'hc0ef6ada, 32'hc2959656};
test_weights[28328:28335] = '{32'h418ef333, 32'h427897b9, 32'h4284b11a, 32'hc1d20e99, 32'hc2baae60, 32'h41ab0a22, 32'hc2bcb7a5, 32'hc2bdd4a4};
test_bias[3541:3541] = '{32'h42c0b566};
test_output[3541:3541] = '{32'h446d3c22};
test_input[28336:28343] = '{32'h423b9579, 32'h42bd3c8c, 32'hbfe7d99c, 32'hc2795f8c, 32'hc2a18fa1, 32'hc212466a, 32'h427d3272, 32'hc23d2745};
test_weights[28336:28343] = '{32'hc281d694, 32'h4144bb4b, 32'hc2677a32, 32'hc2a9b379, 32'h42a15c82, 32'hc2a5f053, 32'hc215441c, 32'hc19e1180};
test_bias[3542:3542] = '{32'h427076fe};
test_output[3542:3542] = '{32'hc4a72afb};
test_input[28344:28351] = '{32'h428f8f6a, 32'h4290c9b1, 32'hc2a1c213, 32'hc1d6243d, 32'h419dde1f, 32'hc27af387, 32'hc1aab274, 32'hc22913c1};
test_weights[28344:28351] = '{32'h427a7c6d, 32'hc11db67b, 32'h4258e3db, 32'hc20b7ed4, 32'hc1cdf885, 32'h41bb71dd, 32'hc211c3f7, 32'h42c053de};
test_bias[3543:3543] = '{32'hc2419033};
test_output[3543:3543] = '{32'hc59bc1f7};
test_input[28352:28359] = '{32'h42055e58, 32'hc29ff5ef, 32'h41550360, 32'h41aac349, 32'h429c08c6, 32'h4210cf38, 32'h4229fa3f, 32'hc23a8172};
test_weights[28352:28359] = '{32'h420e8161, 32'hc2bbc081, 32'h42b52d6a, 32'h41a9966b, 32'hc29360bc, 32'h41451f60, 32'h428f6b29, 32'hc28574a8};
test_bias[3544:3544] = '{32'hc2c0112b};
test_output[3544:3544] = '{32'h462da87f};
test_input[28360:28367] = '{32'h42c6dbf2, 32'hc222bfa3, 32'hc2bd2006, 32'hc223697b, 32'hc198aeda, 32'hc261db5d, 32'h421fb11e, 32'h40d7102f};
test_weights[28360:28367] = '{32'h42a6d976, 32'hc2bc1adc, 32'hc2952449, 32'hc2b67a8b, 32'h42b24e20, 32'h425c9355, 32'h415d5930, 32'h4256bfb7};
test_bias[3545:3545] = '{32'h429494ba};
test_output[3545:3545] = '{32'h469501be};
test_input[28368:28375] = '{32'hc05fc1bd, 32'h4212c634, 32'hc2896165, 32'hc25a0a35, 32'h42c0d207, 32'hc282a85a, 32'hc21dfa0c, 32'h4272723c};
test_weights[28368:28375] = '{32'h41683413, 32'h4211850f, 32'h42636099, 32'hc2b845c6, 32'h419bdd0b, 32'h428c58e3, 32'hc2b8e99c, 32'h42a76a69};
test_bias[3546:3546] = '{32'h41b8453e};
test_output[3546:3546] = '{32'h4603f02b};
test_input[28376:28383] = '{32'hc19424aa, 32'h42c67e0f, 32'hc28a0747, 32'h42700262, 32'h42553ba6, 32'hc20145f7, 32'h42b84455, 32'h41c7ee8c};
test_weights[28376:28383] = '{32'h428c393f, 32'hc1cacc35, 32'h4091e0d4, 32'h420d88d6, 32'h429f8e0a, 32'h41538801, 32'h41ac7864, 32'h420b13aa};
test_bias[3547:3547] = '{32'h4246a8b6};
test_output[3547:3547] = '{32'h4593a5a7};
test_input[28384:28391] = '{32'hc2923031, 32'hc26be95a, 32'hc0c04c46, 32'hc2300aa6, 32'hc13c9441, 32'h41bd5324, 32'hc27616ec, 32'hbf984e3b};
test_weights[28384:28391] = '{32'h42680f5d, 32'hc0da281a, 32'h4091e618, 32'h41a62c37, 32'h42ae5fb2, 32'h4189bea9, 32'h41d6d502, 32'hc14114f5};
test_bias[3548:3548] = '{32'h41a5a000};
test_output[3548:3548] = '{32'hc5db49d7};
test_input[28392:28399] = '{32'hc2a5e762, 32'h42b40cbd, 32'h4234c042, 32'h426e878e, 32'hc24f0c49, 32'hc24660c7, 32'h42b35580, 32'hc2a5437e};
test_weights[28392:28399] = '{32'h429faf93, 32'hc1ba99cf, 32'hc29bedff, 32'hc2825fc6, 32'h42c6ce77, 32'h420c6b64, 32'h41e08ce2, 32'hc0a4b0a4};
test_bias[3549:3549] = '{32'h42b3e17a};
test_output[3549:3549] = '{32'hc69c2716};
test_input[28400:28407] = '{32'hbfbf2bde, 32'h42c5507c, 32'hc22d77d4, 32'h423df8bb, 32'h42025d87, 32'hc176dcb3, 32'h42a99cc3, 32'h4207e129};
test_weights[28400:28407] = '{32'h41b44997, 32'h42385fd9, 32'hc13bc3de, 32'hc2b32e68, 32'hc272fc7c, 32'hc20886fa, 32'h41b22bbc, 32'h42894886};
test_bias[3550:3550] = '{32'hc087dadd};
test_output[3550:3550] = '{32'h455cadeb};
test_input[28408:28415] = '{32'h4294099e, 32'hc1ca4c6b, 32'hc2865afb, 32'h41ce5754, 32'hc292e341, 32'h42186ca8, 32'hc1e115c6, 32'hc1e567bb};
test_weights[28408:28415] = '{32'hc2999049, 32'h4205c0b3, 32'h4293408e, 32'hc22faa85, 32'hc2adfa50, 32'hc1c39b93, 32'h42280b65, 32'h425eaf8a};
test_bias[3551:3551] = '{32'h40091756};
test_output[3551:3551] = '{32'hc61b1b4d};
test_input[28416:28423] = '{32'hc29474ed, 32'hc209960d, 32'hc2abff43, 32'h419cb8b1, 32'h418c568a, 32'hc18fc2f2, 32'hc2446c72, 32'hc2493c2d};
test_weights[28416:28423] = '{32'hc2a87192, 32'h4190985e, 32'h42ac1145, 32'hc223f8fe, 32'h40c34a7e, 32'h40a7d1bd, 32'hc1211b2f, 32'hc2b683e7};
test_bias[3552:3552] = '{32'hc12be1c8};
test_output[3552:3552] = '{32'h451d3b27};
test_input[28424:28431] = '{32'h429d347d, 32'h42a7fe16, 32'hc2b7ee51, 32'hc25176a3, 32'h423b303d, 32'h42a4f489, 32'h4227b9e0, 32'hc1e89a2a};
test_weights[28424:28431] = '{32'hbf16c3bc, 32'hc2697067, 32'hc0601e43, 32'h421b7baf, 32'h428dac18, 32'h4194efb8, 32'h4284f778, 32'h42824945};
test_bias[3553:3553] = '{32'hc297e09b};
test_output[3553:3553] = '{32'hc47864dd};
test_input[28432:28439] = '{32'h42184cb3, 32'h4265a46a, 32'hc2618299, 32'h41929ece, 32'h42893f50, 32'h42a980cc, 32'h42b89f31, 32'h41e32afa};
test_weights[28432:28439] = '{32'hc10a99be, 32'hc26aea45, 32'hc1f77a6d, 32'hc2623d4c, 32'h41700bf0, 32'hc1aa3c54, 32'hc21fda70, 32'h410a4251};
test_bias[3554:3554] = '{32'hc2040801};
test_output[3554:3554] = '{32'hc5e26533};
test_input[28440:28447] = '{32'hc2676c68, 32'h4232ac68, 32'h3f737659, 32'h41e32291, 32'hc2c44b61, 32'hc2abfea4, 32'hc2492928, 32'h42af2236};
test_weights[28440:28447] = '{32'h41f5e0cc, 32'hc2bd8e79, 32'hc28061b5, 32'h4284979b, 32'h42284fb5, 32'hc2b0b00f, 32'h41a64053, 32'hc2843d8e};
test_bias[3555:3555] = '{32'hc2be6da7};
test_output[3555:3555] = '{32'hc5ef2a53};
test_input[28448:28455] = '{32'h41519030, 32'hc0a6e3a9, 32'h429a8601, 32'h41252cab, 32'hc1c3d351, 32'h42297309, 32'hc2c62f18, 32'h42474754};
test_weights[28448:28455] = '{32'hc2be424b, 32'hc22f7d98, 32'h4117201f, 32'h42c47b41, 32'hc1a12c6d, 32'h426ef641, 32'hc2000edc, 32'h413a8a58};
test_bias[3556:3556] = '{32'hc22782cb};
test_output[3556:3556] = '{32'h45e9301d};
test_input[28456:28463] = '{32'h4241590d, 32'h41e73434, 32'h42b19b90, 32'h4129002b, 32'h421828fe, 32'hc2375dc2, 32'hc25c0c1c, 32'h423f80be};
test_weights[28456:28463] = '{32'hc16fb86b, 32'hc24dd592, 32'h4275f6ae, 32'h4260d05e, 32'h428656a3, 32'h41e1593f, 32'h421a60d7, 32'h40a807e5};
test_bias[3557:3557] = '{32'h425451a3};
test_output[3557:3557] = '{32'h454d808f};
test_input[28464:28471] = '{32'hc0f2fafa, 32'h41b1e3e3, 32'h4244fdac, 32'hc2212e48, 32'h42b14663, 32'hc2c6c21f, 32'h42845746, 32'hc0034cfe};
test_weights[28464:28471] = '{32'h42500d60, 32'hc2563059, 32'hc11ada95, 32'hc299b499, 32'h41b2ee3c, 32'h4103ff3a, 32'hc2b2a090, 32'h4177eaa4};
test_bias[3558:3558] = '{32'hc1b2036c};
test_output[3558:3558] = '{32'hc56b6cd0};
test_input[28472:28479] = '{32'hc25ffc33, 32'h42bcd5e5, 32'hc2bb2d2f, 32'h41a60f12, 32'h4118fbc6, 32'h41831391, 32'hc2827953, 32'hc2b5da0d};
test_weights[28472:28479] = '{32'h418a76f3, 32'h42a5f987, 32'hc26c35bd, 32'h41a08801, 32'h405c69a5, 32'hc1800858, 32'h42a7864c, 32'hc1080aff};
test_bias[3559:3559] = '{32'hc26d62ca};
test_output[3559:3559] = '{32'h45f4ac22};
test_input[28480:28487] = '{32'hc215b1f8, 32'hc2bbfd04, 32'hc2c4a42c, 32'h41b280bb, 32'hc25169b5, 32'h42b20cc7, 32'h41f822de, 32'h42260bd3};
test_weights[28480:28487] = '{32'hc293fd2b, 32'h421bc9f6, 32'hc2c0a300, 32'h40be4ee3, 32'h42857821, 32'hc291c821, 32'h41ee887b, 32'h421b80d6};
test_bias[3560:3560] = '{32'h40e4ec1c};
test_output[3560:3560] = '{32'h449f4080};
test_input[28488:28495] = '{32'hc2ae3269, 32'h42adb9fa, 32'h41a59ad8, 32'h42affa18, 32'h42bf9248, 32'hc2be7495, 32'h40d34811, 32'hc1e2938f};
test_weights[28488:28495] = '{32'h418cd592, 32'hc17a1572, 32'h42bd503d, 32'h4287567a, 32'h42bf26a5, 32'hc23bf7da, 32'h4299f220, 32'hc22cbe4a};
test_bias[3561:3561] = '{32'h415d6c2a};
test_output[3561:3561] = '{32'h469f5ad3};
test_input[28496:28503] = '{32'h412f2719, 32'hc14aa0ec, 32'h415a798e, 32'h42044696, 32'h41ae0561, 32'h410ccca1, 32'h41c0d2cd, 32'h42bafe9a};
test_weights[28496:28503] = '{32'h41beeca5, 32'hc28a41c8, 32'h4222bb4d, 32'hc253d161, 32'h4289d667, 32'h42503923, 32'hc289e0cc, 32'h41e61c9c};
test_bias[3562:3562] = '{32'h42ba92f6};
test_output[3562:3562] = '{32'h453cb57f};
test_input[28504:28511] = '{32'hc1ac593e, 32'hc1e48860, 32'h3fc17039, 32'h42415428, 32'hc273c94a, 32'hbf52dc21, 32'h41d2dde4, 32'h42b4bc67};
test_weights[28504:28511] = '{32'h416be435, 32'hc268197b, 32'h41458499, 32'hc124041f, 32'h3f09d15e, 32'h4279a1af, 32'hc225a585, 32'hc299601a};
test_bias[3563:3563] = '{32'h42b304e3};
test_output[3563:3563] = '{32'hc5df89a2};
test_input[28512:28519] = '{32'h42430f1d, 32'h41f18ef0, 32'hc27582dd, 32'hc2b6cbcd, 32'hc24cd8f4, 32'h423146c6, 32'h429e5e20, 32'h418a2d8a};
test_weights[28512:28519] = '{32'hc1a971ef, 32'h42a317b3, 32'h42992e2e, 32'h4016f19e, 32'hc2099176, 32'hc1d34ef1, 32'h42a721b9, 32'h42c71184};
test_bias[3564:3564] = '{32'hc2931560};
test_output[3564:3564] = '{32'h45a7b21d};
test_input[28520:28527] = '{32'h42921c33, 32'hc2428f99, 32'h42828207, 32'h425789f9, 32'hc227537a, 32'hc21d5b04, 32'hc2590115, 32'hc218576a};
test_weights[28520:28527] = '{32'hc2c37bcb, 32'hc1c83c1a, 32'hc1746d1f, 32'hc24c9765, 32'h42bb881f, 32'hc198b43b, 32'h423f6589, 32'h423371f8};
test_bias[3565:3565] = '{32'hc185b14a};
test_output[3565:3565] = '{32'hc6862150};
test_input[28528:28535] = '{32'hbfd0d5a1, 32'h427b5292, 32'hc294d59d, 32'h41aa3387, 32'h425c6ada, 32'h41b5328e, 32'hc2bfd6f2, 32'hc238a693};
test_weights[28528:28535] = '{32'hc28b5f56, 32'hc286abf3, 32'h426ad994, 32'h42a2a809, 32'h421f2e1a, 32'h41b9e302, 32'hc2c3232b, 32'h40f712da};
test_bias[3566:3566] = '{32'h420c4eec};
test_output[3566:3566] = '{32'h459c44a3};
test_input[28536:28543] = '{32'h40ccb3e2, 32'hc2521524, 32'hc085fdac, 32'hc2860702, 32'hc0817787, 32'hc2136d83, 32'h4267e219, 32'h3f303092};
test_weights[28536:28543] = '{32'h42b3c3d2, 32'h429792da, 32'h41491542, 32'h42ae7ded, 32'h42b04ff0, 32'hc1e3e6f8, 32'h42872779, 32'h40b12b23};
test_bias[3567:3567] = '{32'hc290598b};
test_output[3567:3567] = '{32'hc594d208};
test_input[28544:28551] = '{32'hc20b2e92, 32'hc29d94b9, 32'hc262f50c, 32'hc2530720, 32'hc28c09bd, 32'hc26c0e39, 32'h428a1189, 32'h422516c6};
test_weights[28544:28551] = '{32'hc2ac72c6, 32'h42648b5a, 32'h42bddf4e, 32'hc1275f5b, 32'h42b9ca18, 32'h421ab1f0, 32'h3fbecfd3, 32'hc2a17735};
test_bias[3568:3568] = '{32'hc2354903};
test_output[3568:3568] = '{32'hc68fbad8};
test_input[28552:28559] = '{32'hc2aa8b31, 32'h3f9555c1, 32'hc28ae129, 32'hc190db04, 32'hc19066de, 32'hc29bb332, 32'hc2a71eb4, 32'hc1454e00};
test_weights[28552:28559] = '{32'h41ec1af7, 32'h41aeb040, 32'h4169972e, 32'h40b38b7b, 32'h418318e6, 32'h41b8d273, 32'hc1a25615, 32'hc13f0304};
test_bias[3569:3569] = '{32'hc2815f14};
test_output[3569:3569] = '{32'hc5752bfc};
test_input[28560:28567] = '{32'hc1823994, 32'h42975c1e, 32'h429799fc, 32'h417b4600, 32'h429218c8, 32'h42b7c5df, 32'hc26bedd4, 32'hbfa3b7ea};
test_weights[28560:28567] = '{32'hc2c0121b, 32'hc240b74c, 32'hbfdc06fd, 32'h429ccc8c, 32'h42a47d68, 32'hc296c1d8, 32'h427a0104, 32'h424caa24};
test_bias[3570:3570] = '{32'h42aed75e};
test_output[3570:3570] = '{32'hc5ade6e1};
test_input[28568:28575] = '{32'hc28a5d88, 32'h406d4f69, 32'hc10459a9, 32'hc1f6cd0b, 32'h429a0a5a, 32'hc244f6bf, 32'h4283824d, 32'hc28413ed};
test_weights[28568:28575] = '{32'h4089039b, 32'hc205eb44, 32'hc2883dbe, 32'h428560d1, 32'hc2bb94bc, 32'h42badae6, 32'hc22a5bbf, 32'hc298e269};
test_bias[3571:3571] = '{32'hc1fa98cb};
test_output[3571:3571] = '{32'hc634085b};
test_input[28576:28583] = '{32'h42accf5b, 32'h421f1e60, 32'h42c611c4, 32'hc2b6d4d7, 32'hc29ae383, 32'h42b8d96d, 32'h42925ede, 32'hc2a7d5e7};
test_weights[28576:28583] = '{32'hc267aeb0, 32'hc1227c49, 32'hc1432e74, 32'hc2937089, 32'h427278de, 32'hbf775415, 32'h42c233e7, 32'hc14086bd};
test_bias[3572:3572] = '{32'hc1252d48};
test_output[3572:3572] = '{32'h45574750};
test_input[28584:28591] = '{32'h410fd6f0, 32'h3ed34728, 32'hc2113d2b, 32'h428313d8, 32'hc282585d, 32'h423b6a52, 32'h4297a401, 32'hc296d57e};
test_weights[28584:28591] = '{32'hc1158b47, 32'h423de275, 32'hc243decf, 32'hc26d5254, 32'h4254687c, 32'h423bbced, 32'h426181d7, 32'hc25e5393};
test_bias[3573:3573] = '{32'h4191d926};
test_output[3573:3573] = '{32'h459dbf63};
test_input[28592:28599] = '{32'hc1213487, 32'h4278763c, 32'hc2b0c5ef, 32'hc2915648, 32'hc21874d2, 32'hc1f93b92, 32'hc2c166ff, 32'hc1e34a24};
test_weights[28592:28599] = '{32'hc292f7de, 32'hc28d5e0c, 32'h421ceeee, 32'hc2a15417, 32'hc1866d13, 32'h42460581, 32'hc1edc1a5, 32'h415a577f};
test_bias[3574:3574] = '{32'h4100cac0};
test_output[3574:3574] = '{32'h43a82396};
test_input[28600:28607] = '{32'hc190cbe0, 32'hc18b8780, 32'hc2653902, 32'h41915b8e, 32'hc2bbaaab, 32'h42221989, 32'hbf3999ad, 32'h4244959e};
test_weights[28600:28607] = '{32'hc2b1c761, 32'h427e23f9, 32'h42881e02, 32'hc2be23cd, 32'hc21e6e03, 32'hc1e6508b, 32'hc2b8075f, 32'h4251702c};
test_bias[3575:3575] = '{32'h4247ae43};
test_output[3575:3575] = '{32'h42e1cfc4};
test_input[28608:28615] = '{32'hc269daac, 32'hc21a6000, 32'hc2b5b7e9, 32'hc283d997, 32'hc10094e5, 32'hc2002a20, 32'hc23cb1df, 32'hc216f58f};
test_weights[28608:28615] = '{32'hc2ae972f, 32'hc052ed88, 32'h42c690d7, 32'h41fe54fd, 32'hc2399f84, 32'h429e20c1, 32'hc1a462dd, 32'h424e8635};
test_bias[3576:3576] = '{32'h419ef2a6};
test_output[3576:3576] = '{32'hc60cb625};
test_input[28616:28623] = '{32'h42a19a39, 32'hc155f3a3, 32'h41e69a5a, 32'h4203438d, 32'h42b43700, 32'hc2b2f6b5, 32'hc2802457, 32'h41a2ab38};
test_weights[28616:28623] = '{32'hc29d7deb, 32'hc240f57b, 32'h42a7086d, 32'h42bbdc9c, 32'h42892cd5, 32'hc1467377, 32'hc2961ed0, 32'hc26b000d};
test_bias[3577:3577] = '{32'hc2611071};
test_output[3577:3577] = '{32'h4625f229};
test_input[28624:28631] = '{32'hc1fd42e3, 32'hc28cbe0b, 32'h42abdd7d, 32'hc1aa1c51, 32'h423a1100, 32'h41dc20d7, 32'h42c23054, 32'hc2ad0d52};
test_weights[28624:28631] = '{32'hc23859f3, 32'hc298af17, 32'hc214206c, 32'hc21d7696, 32'h3f7dc679, 32'h40372c24, 32'hc12465bb, 32'hc22ab52e};
test_bias[3578:3578] = '{32'h41bb4956};
test_output[3578:3578] = '{32'h45e50baf};
test_input[28632:28639] = '{32'hc1201899, 32'hc29b974a, 32'h41deea0e, 32'h4115be06, 32'hc207c680, 32'h3f9955fd, 32'h41850d5a, 32'h429b2bb4};
test_weights[28632:28639] = '{32'hc1822092, 32'hc1ffcb53, 32'hc1f4e86a, 32'h40f3942d, 32'h41e272a2, 32'h418b289f, 32'h421dd165, 32'hc2912a1f};
test_bias[3579:3579] = '{32'h427ad508};
test_output[3579:3579] = '{32'hc578ff95};
test_input[28640:28647] = '{32'hc19edeb8, 32'hc206671c, 32'h4205d2b5, 32'hc2a46fc7, 32'hc28626dc, 32'hc02e4d94, 32'h42427762, 32'hc28717ac};
test_weights[28640:28647] = '{32'h42abe189, 32'h4186104a, 32'h42478cda, 32'hc23730a1, 32'hc2b2b9f6, 32'hc289a629, 32'h41643780, 32'hc2ae9de8};
test_bias[3580:3580] = '{32'h4096dd9d};
test_output[3580:3580] = '{32'h467916f8};
test_input[28648:28655] = '{32'h422e9d87, 32'h42794770, 32'hc21f7fa4, 32'h409bf7f9, 32'h4293f553, 32'h40664830, 32'hc29faae0, 32'hc1d37a1a};
test_weights[28648:28655] = '{32'hc2c4c68e, 32'hc27f64b2, 32'hc2c24531, 32'hc1398ef7, 32'h41ef21bf, 32'h417b6429, 32'h42bb34df, 32'h418f2be4};
test_bias[3581:3581] = '{32'hc16995a8};
test_output[3581:3581] = '{32'hc61e9745};
test_input[28656:28663] = '{32'hc2168de4, 32'hc1fb8024, 32'hc1a9958b, 32'hc290e905, 32'hc2af0296, 32'h42c6432f, 32'hc23e9f82, 32'h42a8cb43};
test_weights[28656:28663] = '{32'hc1a35649, 32'hc2aa0dac, 32'hc24b0a80, 32'hc2899362, 32'h41aa64f0, 32'h41ea9918, 32'h4296b637, 32'hc25fcec2};
test_bias[3582:3582] = '{32'hc1c5e64d};
test_output[3582:3582] = '{32'h4509eb3f};
test_input[28664:28671] = '{32'h4291aa82, 32'hc28e9968, 32'hc1c3e892, 32'h40928ccd, 32'hc2042b5f, 32'h42320e6c, 32'hc0518691, 32'hc1bee993};
test_weights[28664:28671] = '{32'h4198f2e9, 32'hc260529c, 32'h414ac149, 32'h42376632, 32'hc2c51944, 32'h4292b855, 32'h426b9552, 32'hc1d2eec0};
test_bias[3583:3583] = '{32'hc2c20adf};
test_output[3583:3583] = '{32'h463ddf8a};
test_input[28672:28679] = '{32'h42510772, 32'h42909f84, 32'hc269aecd, 32'h42057a82, 32'h4215cd3f, 32'h4206560d, 32'hc220b5b2, 32'hc26e5480};
test_weights[28672:28679] = '{32'hc27b3950, 32'hc1616fb0, 32'h423b797a, 32'h428ee1bb, 32'hc2b029dc, 32'hc18a4673, 32'h411fcfdc, 32'h4254d7d7};
test_bias[3584:3584] = '{32'h41342620};
test_output[3584:3584] = '{32'hc63cfae0};
test_input[28680:28687] = '{32'hc13f9cb6, 32'h41c556e7, 32'hc2abee1d, 32'h41468a40, 32'hc250cd65, 32'h42548b95, 32'hc24fcbc9, 32'h42517987};
test_weights[28680:28687] = '{32'hc180ebb2, 32'h41e5afb5, 32'h42150721, 32'hc2b551de, 32'h4283b99f, 32'h42779b7f, 32'h424eeac6, 32'h3f9cac6a};
test_bias[3585:3585] = '{32'hc15fe5a1};
test_output[3585:3585] = '{32'hc5c22488};
test_input[28688:28695] = '{32'hc2a387cb, 32'h42c6cc40, 32'h42a5fce7, 32'h4285ff43, 32'hc1963614, 32'hc1e03290, 32'hc1cd8802, 32'h422f6a0a};
test_weights[28688:28695] = '{32'h427bd992, 32'hc29659a5, 32'h4277cb15, 32'hc20ebebf, 32'h42bc2391, 32'hc2acce3b, 32'hc28a2ee7, 32'h41ec0890};
test_bias[3586:3586] = '{32'h41d1add8};
test_output[3586:3586] = '{32'hc5bf3e61};
test_input[28696:28703] = '{32'hc28885f3, 32'hc2a68520, 32'h427d48d4, 32'hc2b09059, 32'hc2a5a7d8, 32'h42219b2f, 32'h42a9a236, 32'hc0e82a5a};
test_weights[28696:28703] = '{32'hc2b6dd19, 32'hc289f2de, 32'h404bc63b, 32'hc289a338, 32'hc13a341c, 32'h42a108a2, 32'hc2889b10, 32'h420fc7e6};
test_bias[3587:3587] = '{32'h42b4e43c};
test_output[3587:3587] = '{32'h46810509};
test_input[28704:28711] = '{32'hc286ceeb, 32'h42b2c704, 32'hc187fd7c, 32'h408f5d83, 32'h42c4b6c4, 32'hc226b68f, 32'h42a91554, 32'hc294ff98};
test_weights[28704:28711] = '{32'hc2c0a964, 32'h42a69182, 32'hc2a471fd, 32'h41d3092b, 32'h42ac62b0, 32'h411cd384, 32'h42949714, 32'hc280df9c};
test_bias[3588:3588] = '{32'hc2ba9a6a};
test_output[3588:3588] = '{32'h4706cefc};
test_input[28712:28719] = '{32'hc25bfc07, 32'h42b00d6d, 32'hc2877553, 32'hc29bed66, 32'h41753b37, 32'h429bccd3, 32'h4292006f, 32'h4296a4d7};
test_weights[28712:28719] = '{32'h4276f908, 32'h427c5895, 32'hc24f8417, 32'h41b2d616, 32'hc296fd35, 32'hc1b0764f, 32'hc25f5d5e, 32'hc29ffc3f};
test_bias[3589:3589] = '{32'h428ff22e};
test_output[3589:3589] = '{32'hc60c4250};
test_input[28720:28727] = '{32'hc2a903c6, 32'hbfdadaf9, 32'hc204ba0d, 32'hc25b2b83, 32'hc2869ddc, 32'hc188cff9, 32'hc0fff7a4, 32'hc2918cd4};
test_weights[28720:28727] = '{32'hc2b6d6f6, 32'h425bc18b, 32'h41750a31, 32'hc2825f3a, 32'h41d8be65, 32'hc2389678, 32'hc1ecfd88, 32'h40bea64c};
test_bias[3590:3590] = '{32'h42a59246};
test_output[3590:3590] = '{32'h46152c0b};
test_input[28728:28735] = '{32'h428691ba, 32'h4272443b, 32'h41b2e71a, 32'hc2bff335, 32'hc2be5fd4, 32'hc29b47a6, 32'hc29df336, 32'h42649d9e};
test_weights[28728:28735] = '{32'hc1969df6, 32'hc2a0373e, 32'h429e9150, 32'hc222a5af, 32'h41d65b1a, 32'h423ac910, 32'h423ff025, 32'h423429ab};
test_bias[3591:3591] = '{32'hc26c0485};
test_output[3591:3591] = '{32'hc5f6ab7f};
test_input[28736:28743] = '{32'hc174b549, 32'h42a13ee0, 32'h4267ac06, 32'h41a35226, 32'hc10e5916, 32'h42a2df8e, 32'h428d2c4c, 32'h424eec1c};
test_weights[28736:28743] = '{32'hc29f9c09, 32'h4208be4f, 32'h425ebc3b, 32'hc24718ab, 32'hc1b001e2, 32'h412974ae, 32'h42b28117, 32'hc2973ab0};
test_bias[3592:3592] = '{32'h424178e5};
test_output[3592:3592] = '{32'h461742b1};
test_input[28744:28751] = '{32'h41b6a123, 32'h40b23759, 32'h41836c23, 32'h407c7f23, 32'h428ca396, 32'h41dfdc57, 32'hc2b252cb, 32'hc25a37f3};
test_weights[28744:28751] = '{32'h41f28fc7, 32'hc23e9d1e, 32'hc2849d67, 32'hc284e553, 32'hc267b5a7, 32'h42a8b14d, 32'h428073ce, 32'hc2779c7c};
test_bias[3593:3593] = '{32'h41859bc4};
test_output[3593:3593] = '{32'hc59b54b9};
test_input[28752:28759] = '{32'h42b05461, 32'h41e8c041, 32'h413a45e1, 32'hc2abb61c, 32'hc0c83731, 32'hc28eb643, 32'h413ded22, 32'h423e10af};
test_weights[28752:28759] = '{32'h419376d1, 32'h426a6901, 32'hc1e5ba68, 32'hc23a93ad, 32'hc29ae6a9, 32'hc237fa93, 32'hc2794677, 32'h41461138};
test_bias[3594:3594] = '{32'hc285149e};
test_output[3594:3594] = '{32'h4624d3f0};
test_input[28760:28767] = '{32'h4268b1d3, 32'h422fe0e2, 32'h421f3094, 32'h413a2692, 32'hc232fb5a, 32'hc2996327, 32'h4194b555, 32'hc189b4fe};
test_weights[28760:28767] = '{32'hc261ce74, 32'h41f24c35, 32'hc242fecc, 32'hc2a8b1ab, 32'hc2668778, 32'h40f121a7, 32'h42075136, 32'h423dc483};
test_bias[3595:3595] = '{32'h419faa50};
test_output[3595:3595] = '{32'hc53e0a83};
test_input[28768:28775] = '{32'hc0a096b0, 32'hbfcf5680, 32'hc01e392f, 32'hc2747947, 32'h40f98192, 32'hc20bde3b, 32'hc1c4b48c, 32'hbe99fec4};
test_weights[28768:28775] = '{32'h423f7680, 32'h42746d9a, 32'hc1c851a5, 32'hc24c782f, 32'h429474f9, 32'hc1fbc0cd, 32'hc2943058, 32'h41c150df};
test_bias[3596:3596] = '{32'h429c1a9a};
test_output[3596:3596] = '{32'h45c8959d};
test_input[28776:28783] = '{32'h41eb9690, 32'h428c5637, 32'hc1b0ffa4, 32'h42bdd588, 32'h428c8143, 32'hc2823c62, 32'h42bec7fb, 32'hc113dad3};
test_weights[28776:28783] = '{32'h410afaaa, 32'hc200341b, 32'hc270c28f, 32'h422ba45c, 32'hc2bd5680, 32'hc094781a, 32'hc1cefede, 32'hc2540a93};
test_bias[3597:3597] = '{32'hc20aa07c};
test_output[3597:3597] = '{32'hc59ab0d5};
test_input[28784:28791] = '{32'hc296a1b9, 32'h4198b093, 32'h42a7a20c, 32'hc200cd17, 32'h420bcef8, 32'hc18b7458, 32'hc28978f3, 32'h41598c9b};
test_weights[28784:28791] = '{32'hc28c652e, 32'hc1c2aee3, 32'h42bdf083, 32'hc22a6d59, 32'hc13962e7, 32'h41975bb3, 32'hc2817d5f, 32'h42aab7fd};
test_bias[3598:3598] = '{32'h42588267};
test_output[3598:3598] = '{32'h46951991};
test_input[28792:28799] = '{32'hc206bcaa, 32'hc27fd7ad, 32'h41396512, 32'h428d90ce, 32'hc2659f6e, 32'hc1021d70, 32'hc0a796a7, 32'h42160f75};
test_weights[28792:28799] = '{32'hc28134d9, 32'h423633d6, 32'hc1c549d6, 32'hc136c0df, 32'h42932e3c, 32'hc19d31f9, 32'hc2933683, 32'h429be387};
test_bias[3599:3599] = '{32'hc289cf24};
test_output[3599:3599] = '{32'hc525f9c6};
test_input[28800:28807] = '{32'h42210b2b, 32'hc1a928e8, 32'hc2bd8e88, 32'hc0e07aa0, 32'h4276bbf6, 32'hc2ab82c2, 32'hc2962635, 32'h42167ef2};
test_weights[28800:28807] = '{32'h42a56d59, 32'hc2ac3481, 32'h429cb725, 32'h41713f93, 32'hc2c64a89, 32'h421d174b, 32'h420d3dde, 32'hc23e957a};
test_bias[3600:3600] = '{32'h42193c55};
test_output[3600:3600] = '{32'hc67e3979};
test_input[28808:28815] = '{32'hc2b8bcd4, 32'hc1ec6d9a, 32'hc1caf0e5, 32'hc1c93cf2, 32'h42168355, 32'h429dddf8, 32'h42ab9b11, 32'h41ca650b};
test_weights[28808:28815] = '{32'hc1a80952, 32'hc235344e, 32'h421ab474, 32'h426accde, 32'h41e03c6e, 32'h42c6ce79, 32'hc26f99a9, 32'h420c968c};
test_bias[3601:3601] = '{32'h4215f80e};
test_output[3601:3601] = '{32'h45ac2a73};
test_input[28816:28823] = '{32'hc186cf33, 32'hc2006b88, 32'hc289930d, 32'h42ad5711, 32'hc1776976, 32'hc253ec09, 32'hc2abe254, 32'hc2a20865};
test_weights[28816:28823] = '{32'h4274e7cf, 32'hc2bb1537, 32'hc1f3124b, 32'h42746ffe, 32'h423d6289, 32'hc2a3f0e8, 32'h425845ef, 32'hc2958c2b};
test_bias[3602:3602] = '{32'h4214c2e9};
test_output[3602:3602] = '{32'h4661436c};
test_input[28824:28831] = '{32'hc2975e29, 32'h42b832b2, 32'hc2b43975, 32'h419fcddd, 32'h42b739e1, 32'h4287942c, 32'hc2217d15, 32'hc2757af7};
test_weights[28824:28831] = '{32'h41ac6668, 32'h4157d173, 32'h42128678, 32'h418da0c6, 32'h41b3ddc4, 32'hc25af09b, 32'hc0f7cedd, 32'h42a8773c};
test_bias[3603:3603] = '{32'h429fc097};
test_output[3603:3603] = '{32'hc6188e29};
test_input[28832:28839] = '{32'hc284b9cb, 32'hc200d143, 32'h427f03d5, 32'h42961bb2, 32'h423aad60, 32'h41b7c560, 32'hc2a06661, 32'h42a0b0b3};
test_weights[28832:28839] = '{32'h41c3fb37, 32'h426fd773, 32'h425eff09, 32'h42b4f2ce, 32'hc29285a0, 32'h401deb1b, 32'hc1d0978f, 32'hc281d54b};
test_bias[3604:3604] = '{32'h42ab63fe};
test_output[3604:3604] = '{32'h43c1585e};
test_input[28840:28847] = '{32'hc282dc92, 32'h41ca4d45, 32'h41b30d18, 32'hc13bb2d3, 32'hc13080f5, 32'hc0d06ddf, 32'h42ac31fb, 32'hc2bcdce1};
test_weights[28840:28847] = '{32'h426e01d4, 32'hc226527c, 32'hc22d609c, 32'hc0435ad9, 32'h4181b1a8, 32'hc2c5c8a1, 32'h427e8f69, 32'h423bc03c};
test_bias[3605:3605] = '{32'hc1f4aa0e};
test_output[3605:3605] = '{32'hc5896bb6};
test_input[28848:28855] = '{32'h42a589fc, 32'hc22939eb, 32'hbfa3ae7f, 32'hc191ebe2, 32'hc25f3d5b, 32'hc21c2d4a, 32'hc2c4dda6, 32'h42563de8};
test_weights[28848:28855] = '{32'hc2a2c95e, 32'h42b08e0d, 32'hc2615414, 32'h4264ba93, 32'hc23c5e8d, 32'hc2c69b92, 32'hc21876a9, 32'h42c50384};
test_bias[3606:3606] = '{32'hc121dbd6};
test_output[3606:3606] = '{32'h457f0b31};
test_input[28856:28863] = '{32'hc2acdf2f, 32'hc251ccec, 32'hc2bd6677, 32'hc2c33203, 32'h41d20562, 32'hc220d54c, 32'hc21bdf3d, 32'hc2630c98};
test_weights[28856:28863] = '{32'h4204f034, 32'hc0e544fd, 32'hc2045985, 32'h42b3392a, 32'hc23dd01e, 32'hc293f22e, 32'h42b559c4, 32'h42a000ae};
test_bias[3607:3607] = '{32'hc16c5aed};
test_output[3607:3607] = '{32'hc662185c};
test_input[28864:28871] = '{32'h42b4ed6f, 32'hc1107456, 32'h41c8274e, 32'h429c2e4f, 32'h4106bfc2, 32'h41f7f639, 32'h4167eb8a, 32'h423a917b};
test_weights[28864:28871] = '{32'h42b23b67, 32'hc240a3b1, 32'hc2c07726, 32'hc269557c, 32'hc1db779c, 32'h4227808e, 32'hc2903a28, 32'hc2a02935};
test_bias[3608:3608] = '{32'hc260bc06};
test_output[3608:3608] = '{32'hc50bc108};
test_input[28872:28879] = '{32'h42baf190, 32'h41e61faf, 32'hc295ca8a, 32'hc28d3398, 32'hc11b51f8, 32'hc234bad0, 32'hc23fca53, 32'hc2baf3cc};
test_weights[28872:28879] = '{32'hc2ae061e, 32'hc2500a26, 32'hc1858048, 32'hc25845d1, 32'hc0f08fb3, 32'h426dd4aa, 32'h42bcbd41, 32'h42a51b38};
test_bias[3609:3609] = '{32'hc25225c7};
test_output[3609:3609] = '{32'hc6981b71};
test_input[28880:28887] = '{32'hc29009d8, 32'h42c5b45d, 32'h4249a794, 32'hc2a5a3b0, 32'hc27b7e8d, 32'hc25986ae, 32'h417642e4, 32'hc27b6889};
test_weights[28880:28887] = '{32'hc25701eb, 32'h42bb3f64, 32'h42410b3f, 32'hc23e2a85, 32'h41bb2ea8, 32'hc1c3db4e, 32'h4229745a, 32'h4254deb7};
test_bias[3610:3610] = '{32'h42962ea1};
test_output[3610:3610] = '{32'h4682c617};
test_input[28888:28895] = '{32'h42752137, 32'hc219dc80, 32'h41c9ccbe, 32'h42727d79, 32'h4211287b, 32'hc232e17c, 32'h41cfce3f, 32'h412a482d};
test_weights[28888:28895] = '{32'h420eab18, 32'hc21619ec, 32'h41299306, 32'h42058863, 32'hc23dc8b4, 32'hc2a35674, 32'hc1932303, 32'h4296bb8e};
test_bias[3611:3611] = '{32'h42a264e9};
test_output[3611:3611] = '{32'h46010139};
test_input[28896:28903] = '{32'hc0d553d2, 32'hc28726b0, 32'h42812881, 32'h41b95613, 32'h42c7aa7a, 32'h41d283f9, 32'hc2be8876, 32'hc2a64d98};
test_weights[28896:28903] = '{32'h42c05ab2, 32'hc2a682f4, 32'h42b53f58, 32'h41b6c951, 32'h42816b99, 32'h4273a2ca, 32'hc27c06e8, 32'hc2879e46};
test_bias[3612:3612] = '{32'hc2a62297};
test_output[3612:3612] = '{32'h46f216d2};
test_input[28904:28911] = '{32'h417bb38e, 32'hc1ea69d1, 32'hc25a925d, 32'hc2514bee, 32'hc2b1dd39, 32'hc2576f74, 32'hc1bcb741, 32'hc22e24f7};
test_weights[28904:28911] = '{32'h420620d4, 32'h423e1325, 32'h409f9abd, 32'h425a66ee, 32'h4288baf9, 32'hbf95ea24, 32'hc28be637, 32'h427d8131};
test_bias[3613:3613] = '{32'h4200df4b};
test_output[3613:3613] = '{32'hc62d3fe4};
test_input[28912:28919] = '{32'hc23c58b8, 32'h42c7a168, 32'h41385141, 32'hc2866ad4, 32'hc2c2986c, 32'hc04c059f, 32'h422f01f2, 32'h42986a53};
test_weights[28912:28919] = '{32'hc21dc68a, 32'h429c1a93, 32'h42c552cf, 32'h427f205d, 32'hc294239e, 32'hc180c18c, 32'h425ac8ce, 32'hc01b90cd};
test_bias[3614:3614] = '{32'h4271ee1a};
test_output[3614:3614] = '{32'h467a6165};
test_input[28920:28927] = '{32'hc1e847a9, 32'h428b9a41, 32'hc2b8d985, 32'hc2ad17d0, 32'h422fc193, 32'hc252ac0a, 32'h40c7de8f, 32'h429ff821};
test_weights[28920:28927] = '{32'hc2a2a044, 32'h40ca5174, 32'h4283b0c6, 32'hc24415a4, 32'hc196c8b9, 32'h41cdd7c3, 32'h429996ef, 32'hc1becbbc};
test_bias[3615:3615] = '{32'hc2a0fcf9};
test_output[3615:3615] = '{32'hc52aca77};
test_input[28928:28935] = '{32'h42661192, 32'h4199f918, 32'h42c14408, 32'h42ad0fbf, 32'hc186742a, 32'h42b0f594, 32'hc27bee0f, 32'h42281f0d};
test_weights[28928:28935] = '{32'h4234723a, 32'hbe953949, 32'h42771dd1, 32'h41acfb3c, 32'h429da2d1, 32'h422a101d, 32'hc2aadbbf, 32'h4255a5de};
test_bias[3616:3616] = '{32'h42505a2d};
test_output[3616:3616] = '{32'h46a08150};
test_input[28936:28943] = '{32'hc2943eb4, 32'h42a49b1b, 32'hc2c73d52, 32'h3e4069ec, 32'hc184860f, 32'hc216befc, 32'h41e32393, 32'hc2a9ffac};
test_weights[28936:28943] = '{32'h413ed9e9, 32'hc26c704c, 32'h429bb479, 32'hc2c5993b, 32'hc2aa3ca6, 32'hc2190728, 32'hc1e8eeb6, 32'hc2390427};
test_bias[3617:3617] = '{32'hc2ac4b72};
test_output[3617:3617] = '{32'hc5ef25d7};
test_input[28944:28951] = '{32'hc19b2d2e, 32'h42724de6, 32'h42548296, 32'hc27af76e, 32'hc2c1ffec, 32'h4215b537, 32'hc262fba2, 32'h40d8e562};
test_weights[28944:28951] = '{32'hc2522aa2, 32'h4293e2b1, 32'h4282fd63, 32'hc26720b3, 32'h41919b5f, 32'hc285bf48, 32'h415b4b64, 32'h4211c57a};
test_bias[3618:3618] = '{32'hc290da25};
test_output[3618:3618] = '{32'h45f19da3};
test_input[28952:28959] = '{32'hc29e6b02, 32'h4278d69f, 32'h4283fa69, 32'h422c8f54, 32'h41555ce0, 32'hc2c366ad, 32'hc2a9e287, 32'hc29315e9};
test_weights[28952:28959] = '{32'hc1e56925, 32'h42b0c670, 32'hc15ed6fe, 32'hc0cf49eb, 32'h42bf39f6, 32'h4140c080, 32'hc2883e47, 32'h41ff0d88};
test_bias[3619:3619] = '{32'h424632c2};
test_output[3619:3619] = '{32'h461ec32a};
test_input[28960:28967] = '{32'h427448af, 32'hc28350b6, 32'hc18f0c55, 32'hc253a720, 32'hc29f97c0, 32'h42c6e1b9, 32'h42b2dd77, 32'h4243ea8d};
test_weights[28960:28967] = '{32'hc2a7f40c, 32'hc2190a2a, 32'hc1b15b0e, 32'hc1c5093d, 32'hc17265ba, 32'hc1f308d0, 32'hc215fd6b, 32'h420ce4fa};
test_bias[3620:3620] = '{32'hc2a9984b};
test_output[3620:3620] = '{32'hc58acfa8};
test_input[28968:28975] = '{32'h420d85be, 32'h402c3d09, 32'hc2477148, 32'h421d9488, 32'hc22a464f, 32'hc1e083cd, 32'hc2b9f99d, 32'h41318592};
test_weights[28968:28975] = '{32'h40f38d8e, 32'hc25e8714, 32'hc261d852, 32'h423a5639, 32'hc235e267, 32'hc2a9ae62, 32'h42015d65, 32'hc1fa9ee9};
test_bias[3621:3621] = '{32'hc2997d40};
test_output[3621:3621] = '{32'h45b0b76e};
test_input[28976:28983] = '{32'h4217ab11, 32'hc2865817, 32'hc28eeff6, 32'h42a0689c, 32'hc278d741, 32'hc14813f0, 32'h40ac6209, 32'h4256042e};
test_weights[28976:28983] = '{32'h4201ed6c, 32'hc26b7aa8, 32'h42044c0b, 32'h42ad254d, 32'hc291bb3c, 32'h42b854cb, 32'hc272bf06, 32'h413e2f9f};
test_bias[3622:3622] = '{32'hc27ab22c};
test_output[3622:3622] = '{32'h46514282};
test_input[28984:28991] = '{32'hc124263c, 32'hc25aaab1, 32'hc26e98e5, 32'hc0babc25, 32'h41928898, 32'hc2a6492c, 32'hc1fd0ffb, 32'h41f9b431};
test_weights[28984:28991] = '{32'h41cc8f51, 32'hc1c0ced7, 32'hc2001ff1, 32'hbfa2fa4c, 32'hc179fbef, 32'hc2a4458a, 32'hbf803cc0, 32'hc29cf61a};
test_bias[3623:3623] = '{32'hc1561145};
test_output[3623:3623] = '{32'h45dd664b};
test_input[28992:28999] = '{32'hc15aa78c, 32'h41c6d2a9, 32'hc29a8170, 32'hc2b1d227, 32'hc29fb86b, 32'h427d3cf9, 32'h421c1d4f, 32'h41b8c68f};
test_weights[28992:28999] = '{32'h42c58629, 32'hc2bf3ef4, 32'hc0e23447, 32'h415c0419, 32'h42a77fcc, 32'hc27d0155, 32'hc1a355c4, 32'h42a32137};
test_bias[3624:3624] = '{32'hc28d2de9};
test_output[3624:3624] = '{32'hc65bfb95};
test_input[29000:29007] = '{32'h41936a70, 32'hc17af13a, 32'h424a8cd3, 32'h424eec05, 32'hc2c42044, 32'h41a83901, 32'hc213f62b, 32'hc2ae462c};
test_weights[29000:29007] = '{32'hbfb227b7, 32'h41a32132, 32'h4299ab6f, 32'hc28b226d, 32'h42a79ba5, 32'hc1ff56aa, 32'h4206aec2, 32'h414d4ffd};
test_bias[3625:3625] = '{32'hc280370e};
test_output[3625:3625] = '{32'hc631a9cd};
test_input[29008:29015] = '{32'h418cbe0c, 32'hc1ab9496, 32'h427ed3e0, 32'h42c59695, 32'h428914e6, 32'hc2096c84, 32'hc2230c3f, 32'h420cbaa4};
test_weights[29008:29015] = '{32'hc21511be, 32'h42bee340, 32'h4187aa20, 32'hc241ecd1, 32'hc14fac52, 32'h41b7bb53, 32'h41f73bf1, 32'h4256d3d8};
test_bias[3626:3626] = '{32'hc2a47abb};
test_output[3626:3626] = '{32'hc5ebb8ad};
test_input[29016:29023] = '{32'h42b39a47, 32'h42ba1901, 32'h413a5f5c, 32'h41efa6c6, 32'h41878c5f, 32'h428d181b, 32'hc216eebc, 32'h421310c6};
test_weights[29016:29023] = '{32'hc25df0ef, 32'h4258d859, 32'h42217fe1, 32'h42819a05, 32'hc095fc3d, 32'hc0766532, 32'h41fa43e4, 32'hbfb1c242};
test_bias[3627:3627] = '{32'hc20c5841};
test_output[3627:3627] = '{32'h4455e482};
test_input[29024:29031] = '{32'hc2759c82, 32'h428dab61, 32'h41e3592e, 32'hc26d1917, 32'hc2ac5de3, 32'h4124bd1c, 32'h42a2be13, 32'hc28cb572};
test_weights[29024:29031] = '{32'hc293e8ca, 32'h420529b3, 32'h40c79fdc, 32'hc122bc1e, 32'hc2b42a3f, 32'hc29b90e4, 32'h42837654, 32'h4284eab1};
test_bias[3628:3628] = '{32'hc2839e83};
test_output[3628:3628] = '{32'h466e44fc};
test_input[29032:29039] = '{32'h42c5fec4, 32'hc202ff58, 32'h426b1d7e, 32'hc143ddb3, 32'h4152ef91, 32'h42a42f5c, 32'hc2a144d9, 32'h41c1f332};
test_weights[29032:29039] = '{32'hc29cf387, 32'hc1ccabc0, 32'h3f5b5033, 32'hc27fdc90, 32'hc28308eb, 32'hc29c1881, 32'hc1e051a9, 32'hc28c14bd};
test_bias[3629:3629] = '{32'hc262bd76};
test_output[3629:3629] = '{32'hc648f928};
test_input[29040:29047] = '{32'hc2b27e28, 32'h4292572c, 32'hc132b683, 32'h405772d6, 32'h42a25cd9, 32'h41bf009e, 32'h41a945e9, 32'h40f21b58};
test_weights[29040:29047] = '{32'hc2ad55ef, 32'h42b707d7, 32'hc1b3fcc1, 32'h4239cb17, 32'hc223c542, 32'hc2ba1c09, 32'h4286e672, 32'hc2a373aa};
test_bias[3630:3630] = '{32'h4250846f};
test_output[3630:3630] = '{32'h461ea89d};
test_input[29048:29055] = '{32'h42c65864, 32'h414e0288, 32'hc267a4e4, 32'h41a6042f, 32'h41bcaf63, 32'h4132e0d5, 32'h4225c5d3, 32'h429dff06};
test_weights[29048:29055] = '{32'h42bee607, 32'h41de2df5, 32'hc0b5d5ed, 32'hc299b5c0, 32'h4295f409, 32'hc20cf2ac, 32'hc2bba41f, 32'hc2304d56};
test_bias[3631:3631] = '{32'hc24edad8};
test_output[3631:3631] = '{32'h451ce532};
test_input[29056:29063] = '{32'hc142bbf8, 32'h42807841, 32'hc0f92bff, 32'h42c2f9c5, 32'hc0328b97, 32'h42a94aad, 32'hc28ea118, 32'h3f907afa};
test_weights[29056:29063] = '{32'h424326b7, 32'h40cfec79, 32'hc27f0ea4, 32'h421ec69b, 32'hc27c2b6e, 32'h427f32ef, 32'h41ab154d, 32'hc11f1122};
test_bias[3632:3632] = '{32'hc22b03dc};
test_output[3632:3632] = '{32'h45ffd7a8};
test_input[29064:29071] = '{32'hc1fa6600, 32'hc1c3ca99, 32'h42235e99, 32'hc24b5725, 32'hc2aeac2e, 32'h41f3ef6f, 32'h4287553b, 32'h41c7f466};
test_weights[29064:29071] = '{32'hc1fada54, 32'hc2981fd5, 32'hc150d61a, 32'h41fac746, 32'hc29a6554, 32'hc2a86365, 32'h41e00282, 32'h400e3052};
test_bias[3633:3633] = '{32'h4105f171};
test_output[3633:3633] = '{32'h45d60f9a};
test_input[29072:29079] = '{32'hc2b3c246, 32'h41a348ec, 32'h42936143, 32'h4298d32a, 32'hc191d5e8, 32'h426b71a2, 32'h427949f6, 32'hc10a59ff};
test_weights[29072:29079] = '{32'hc0f25c01, 32'hc2b9ae21, 32'h4235400e, 32'hc2bff2ed, 32'h42c18731, 32'h4204d597, 32'hc1fde1ed, 32'hc27a6d36};
test_bias[3634:3634] = '{32'hc20706b6};
test_output[3634:3634] = '{32'hc5cac1ee};
test_input[29080:29087] = '{32'hc2aecb0b, 32'h4296d205, 32'hc23f2c6d, 32'hc18520ef, 32'h42a4dbf3, 32'h422c7b9f, 32'hc21a307c, 32'hc25b0725};
test_weights[29080:29087] = '{32'h4284074d, 32'hc18d2761, 32'h40d5a05e, 32'h429d3b94, 32'h42047474, 32'hc2c289bd, 32'h413f70a0, 32'hc2c6e3e7};
test_bias[3635:3635] = '{32'h41b0cf1a};
test_output[3635:3635] = '{32'hc5a20ee0};
test_input[29088:29095] = '{32'h4244abd9, 32'hc1c8193f, 32'hc29966f4, 32'hc2659c80, 32'h422e264e, 32'hc19d7c42, 32'h423245ca, 32'hc2614f75};
test_weights[29088:29095] = '{32'hc2aab74c, 32'h42a2dc42, 32'hc1d4a8f1, 32'h41177cf1, 32'hc265755c, 32'hc0542b33, 32'h423fc782, 32'h4228e6ba};
test_bias[3636:3636] = '{32'hc2c14845};
test_output[3636:3636] = '{32'hc5eaa5e0};
test_input[29096:29103] = '{32'hc20265a2, 32'hc2481b64, 32'h4223d3b2, 32'hc25aeb82, 32'hc28090fb, 32'hc24709e1, 32'h423a7ec7, 32'h42137a7b};
test_weights[29096:29103] = '{32'h41b345e6, 32'h42ae519a, 32'h429c547a, 32'h421f8202, 32'hc2acba84, 32'h4240dcc7, 32'h413753c2, 32'h4243a05c};
test_bias[3637:3637] = '{32'hc2b16f42};
test_output[3637:3637] = '{32'h44a62acf};
test_input[29104:29111] = '{32'h42892c31, 32'h42054a09, 32'h42646b6f, 32'h41d80d75, 32'hc2c3e51b, 32'h42aeede2, 32'h42a6e84e, 32'h41daf590};
test_weights[29104:29111] = '{32'h411538d0, 32'hc2c39ed5, 32'hc1a4d545, 32'h417d256a, 32'hc233a322, 32'hc251db68, 32'h4153e78c, 32'hc08fa1ae};
test_bias[3638:3638] = '{32'hc1697e0c};
test_output[3638:3638] = '{32'hc521f1a1};
test_input[29112:29119] = '{32'hc22c1348, 32'hc2b8b1ca, 32'hc2b73e91, 32'hc1f7ca56, 32'h4294ef96, 32'hc1048be5, 32'hc2246a1f, 32'hc26d7874};
test_weights[29112:29119] = '{32'h4240921a, 32'hc2912e92, 32'hc1e103be, 32'h428e7bb2, 32'h4113810c, 32'hc1c96ff1, 32'h42b8d0d7, 32'hc28db855};
test_bias[3639:3639] = '{32'h420f78fe};
test_output[3639:3639] = '{32'h45c63367};
test_input[29120:29127] = '{32'hc12fc11c, 32'h4229416b, 32'hc1a2e301, 32'hc2640961, 32'h42802429, 32'h410221b2, 32'hc2ad4c16, 32'hc19a8e6d};
test_weights[29120:29127] = '{32'h420e18fb, 32'hc213eff1, 32'h426fd18e, 32'hc2bc6da4, 32'hc22e5030, 32'hc2b30466, 32'h42b82831, 32'hc1da6946};
test_bias[3640:3640] = '{32'hc1ece787};
test_output[3640:3640] = '{32'hc6099633};
test_input[29128:29135] = '{32'hc260ed33, 32'h42b67b5e, 32'hc1ce89e6, 32'h42941fdf, 32'hc204c63f, 32'h42850c67, 32'h42b60044, 32'h41153053};
test_weights[29128:29135] = '{32'h42bfc725, 32'hc22dc7bb, 32'hc223f6cb, 32'h42a9ea4e, 32'h427f8fdc, 32'hc0aedc44, 32'hc2bda0ee, 32'hc276f4d6};
test_bias[3641:3641] = '{32'hc2a9d504};
test_output[3641:3641] = '{32'hc6574a29};
test_input[29136:29143] = '{32'h42bdd7bd, 32'h40975824, 32'h422c5627, 32'hc27cc0a0, 32'h42aee1c2, 32'h42a4ca61, 32'h41501220, 32'hc294a7a0};
test_weights[29136:29143] = '{32'h42c691b7, 32'hc29073eb, 32'h428b79dd, 32'hc26c2119, 32'h41e4c72f, 32'hc28ebcc2, 32'h42976284, 32'hc15ce98d};
test_bias[3642:3642] = '{32'h426eb1d2};
test_output[3642:3642] = '{32'h4662af07};
test_input[29144:29151] = '{32'h41d93844, 32'h41d47e80, 32'h429ff7c4, 32'h42196872, 32'hc26b2770, 32'hc203640d, 32'hc1d1f3bb, 32'h423f6dfd};
test_weights[29144:29151] = '{32'hc19c7565, 32'hc29aaa19, 32'h42b4f575, 32'hc0d29fed, 32'h41051de0, 32'hbef62a3e, 32'h41baea4e, 32'h42279300};
test_bias[3643:3643] = '{32'hc1f3afeb};
test_output[3643:3643] = '{32'h45a53a8d};
test_input[29152:29159] = '{32'hc1154b89, 32'h429d67d2, 32'hc2574483, 32'h42b05e88, 32'h413e723f, 32'h4126b7ab, 32'hc2bca4fd, 32'hc216f611};
test_weights[29152:29159] = '{32'h422305bd, 32'h42437a13, 32'h418d5573, 32'h428a0704, 32'hc21a90ab, 32'h426a9dcd, 32'h4140fb08, 32'h426b676e};
test_bias[3644:3644] = '{32'h427371f7};
test_output[3644:3644] = '{32'h45aa7354};
test_input[29160:29167] = '{32'h42c740ce, 32'hc221a420, 32'hc2632182, 32'hc0756716, 32'hc1c14dd9, 32'hc042bee0, 32'h42a85122, 32'hc1aaf8fd};
test_weights[29160:29167] = '{32'h42a73702, 32'hc2afe760, 32'h4272c720, 32'h40c46132, 32'hc29895d3, 32'h42c7599b, 32'h40be397e, 32'h41dab33e};
test_bias[3645:3645] = '{32'h42bf3f59};
test_output[3645:3645] = '{32'h461bb64b};
test_input[29168:29175] = '{32'hc1c814c1, 32'hc070a17e, 32'h41c2f10b, 32'hc07db624, 32'hc21157f9, 32'hc2a15513, 32'h41b017ae, 32'h423d090c};
test_weights[29168:29175] = '{32'h42bdac2c, 32'h42465242, 32'h42bc0b0e, 32'hc253f668, 32'hc2872f9c, 32'hc22d29f6, 32'h4204df16, 32'hc28b356d};
test_bias[3646:3646] = '{32'h426be013};
test_output[3646:3646] = '{32'h4553fc50};
test_input[29176:29183] = '{32'hc2634690, 32'h41da33bf, 32'hc1e2b48b, 32'h422dfc35, 32'h4123c522, 32'hc0034ff6, 32'h427483b1, 32'hc197344e};
test_weights[29176:29183] = '{32'h42a04fdf, 32'h41836324, 32'hc07c42d3, 32'hc0879956, 32'hc2b4cdfa, 32'hc1b9f800, 32'hc248e65a, 32'h42308947};
test_bias[3647:3647] = '{32'h42b467ba};
test_output[3647:3647] = '{32'hc60a9b39};
test_input[29184:29191] = '{32'h41a67e41, 32'hc0bbceec, 32'h42bd6b29, 32'h41253e02, 32'h42929ce7, 32'hc2291b9a, 32'hc297ce69, 32'h428c012d};
test_weights[29184:29191] = '{32'h42c37648, 32'hc2bb475a, 32'h4253c5c1, 32'hc23782bf, 32'h417a6840, 32'h4268f8e7, 32'h4230f529, 32'h42a85794};
test_bias[3648:3648] = '{32'hc14a2f59};
test_output[3648:3648] = '{32'h460229e2};
test_input[29192:29199] = '{32'h42900e30, 32'hc222b260, 32'h422f9c45, 32'hc1e38c26, 32'hc194aeb9, 32'hc25dd32d, 32'h4274b87f, 32'hbf357016};
test_weights[29192:29199] = '{32'hc29e84a3, 32'h429188a6, 32'hc0ebd995, 32'hc28ad4f7, 32'h4111be3e, 32'h42a2821f, 32'hc26dcfc6, 32'hc1155325};
test_bias[3649:3649] = '{32'h429f29ff};
test_output[3649:3649] = '{32'hc66e30db};
test_input[29200:29207] = '{32'h40be910a, 32'h42bb8ded, 32'hc19a9c9e, 32'hc2417eed, 32'hc1712315, 32'h4201a76d, 32'hc217a816, 32'h42ac1efd};
test_weights[29200:29207] = '{32'hc206eef8, 32'h4263b70f, 32'h42b2afe3, 32'hc0612b46, 32'hc2a682e2, 32'hc144b4fd, 32'hc220bb18, 32'h3fc8db0c};
test_bias[3650:3650] = '{32'h427a332a};
test_output[3650:3650] = '{32'h45c07490};
test_input[29208:29215] = '{32'h42bd8a4f, 32'h421deede, 32'hc2489233, 32'hc19fd76b, 32'h42a6ff26, 32'h428696db, 32'h42944998, 32'hc24273be};
test_weights[29208:29215] = '{32'h4246413a, 32'hc219a70a, 32'h421d1ad4, 32'hc1a7e2e4, 32'hc26af7b5, 32'h42b9f852, 32'hc0e8ebaa, 32'h41bb09bc};
test_bias[3651:3651] = '{32'hc2c54ba9};
test_output[3651:3651] = '{32'h449700ba};
test_input[29216:29223] = '{32'hc24ad053, 32'hc1df2f5c, 32'hc24a14cc, 32'h42718352, 32'h41e4ca89, 32'hc186b650, 32'h423e12a3, 32'h425b3e9e};
test_weights[29216:29223] = '{32'hc2787b0b, 32'h42a17ee5, 32'hc24de0e0, 32'hc19f2975, 32'h42a34af4, 32'hc21092c7, 32'hbeecb5ce, 32'h427b32a4};
test_bias[3652:3652] = '{32'h412f4327};
test_output[3652:3652] = '{32'h46077ae5};
test_input[29224:29231] = '{32'h429290d2, 32'hc2927b6e, 32'h421f2d44, 32'hc2b0e0ac, 32'hc243f521, 32'hc1b7c11d, 32'h421a4e36, 32'hc236e881};
test_weights[29224:29231] = '{32'hc1528a98, 32'h41c095db, 32'hc10bf314, 32'hc290821d, 32'hc1ff2249, 32'h40afb759, 32'hc2b92f8e, 32'hc1efb040};
test_bias[3653:3653] = '{32'hc042ef1a};
test_output[3653:3653] = '{32'h451f1d9b};
test_input[29232:29239] = '{32'h42706162, 32'hc142e144, 32'hc22e7e6a, 32'h4224880e, 32'h42b16c91, 32'hc2b8606d, 32'h40bdc8c7, 32'hc1be727f};
test_weights[29232:29239] = '{32'hc262e099, 32'h42a61b67, 32'hc25cc0e6, 32'hc0cec4fd, 32'hc29151d7, 32'hc28a7c78, 32'h425e98bc, 32'h421a37b5};
test_bias[3654:3654] = '{32'hc29a9428};
test_output[3654:3654] = '{32'hc53bde31};
test_input[29240:29247] = '{32'h4275ba44, 32'h41bf5dea, 32'hc2837f4b, 32'h428065cf, 32'hc1246a3e, 32'h4252621f, 32'h42be3847, 32'hc1a2d59c};
test_weights[29240:29247] = '{32'hc2a66370, 32'hc23808ab, 32'hc1c9258a, 32'hc2a1bab5, 32'hc2b32cfc, 32'hc1e96e7b, 32'hc2c15eeb, 32'hc11893b1};
test_bias[3655:3655] = '{32'h4197ca6a};
test_output[3655:3655] = '{32'hc69724c0};
test_input[29248:29255] = '{32'hc283c376, 32'h42351288, 32'h420b4ac2, 32'hbf0da61e, 32'h42a704bd, 32'hc26727f5, 32'hc2919695, 32'h4189e993};
test_weights[29248:29255] = '{32'h42b7c196, 32'h41dac885, 32'hc2962600, 32'hc29ef106, 32'h428bc8bc, 32'hc29da07f, 32'hc1062868, 32'h42c10a35};
test_bias[3656:3656] = '{32'h418cb6bb};
test_output[3656:3656] = '{32'h45a58cee};
test_input[29256:29263] = '{32'h41fb3920, 32'hc2bc3529, 32'h41684f07, 32'h4228be48, 32'hc22429fd, 32'h40b68877, 32'hc2953e93, 32'h42c5e835};
test_weights[29256:29263] = '{32'h426052c4, 32'hc24a34de, 32'h42a8514e, 32'h426d2b9d, 32'h4188206d, 32'hc21e39da, 32'h42bad328, 32'hc24a467d};
test_bias[3657:3657] = '{32'h42a5748e};
test_output[3657:3657] = '{32'hc520e6d5};
test_input[29264:29271] = '{32'hc28d94b5, 32'h4280e28b, 32'h42563ed9, 32'h41cde42b, 32'h420224d9, 32'hc2ac0fe3, 32'hc1efc083, 32'h4034406f};
test_weights[29264:29271] = '{32'hc26f072c, 32'h4214c154, 32'h416bdc94, 32'h42c7e037, 32'h41653fbf, 32'hc2957a82, 32'hc1a157ea, 32'h40ef1b7b};
test_bias[3658:3658] = '{32'h4191eac8};
test_output[3658:3658] = '{32'h4688f04a};
test_input[29272:29279] = '{32'hc2393f2d, 32'hc2293605, 32'hc104dbbf, 32'hc20b6f81, 32'h428fb19d, 32'h42008320, 32'h423b8c89, 32'h428bc6ab};
test_weights[29272:29279] = '{32'hc264f97f, 32'hc208c0da, 32'h42266bd1, 32'hc24d05a8, 32'hc2b3e400, 32'h422f05cd, 32'hc257afdf, 32'h426ac3a0};
test_bias[3659:3659] = '{32'hc24f1f92};
test_output[3659:3659] = '{32'h44fa7a20};
test_input[29280:29287] = '{32'hc1387cae, 32'hc28d076a, 32'hc281d9c2, 32'hc29d0bb6, 32'h425ad35d, 32'hc1be05c3, 32'hc22c2584, 32'h4207c8bb};
test_weights[29280:29287] = '{32'h42bf9f75, 32'h424940b0, 32'h428ac2e7, 32'hc122aaa9, 32'h42891cae, 32'h426807bd, 32'hc205ff06, 32'hc189e2db};
test_bias[3660:3660] = '{32'hc26ddb03};
test_output[3660:3660] = '{32'hc5a2286d};
test_input[29288:29295] = '{32'h424f0284, 32'h41c47a88, 32'hc2ac3b8e, 32'hc28479ff, 32'hc230f7ab, 32'h42ba5184, 32'hc287c33b, 32'h423691ba};
test_weights[29288:29295] = '{32'h42931e07, 32'hc1bad6f0, 32'h42bea8c3, 32'hc28be569, 32'h428ae38e, 32'hc22cd863, 32'h4236b626, 32'hc1df4fab};
test_bias[3661:3661] = '{32'h40960a2a};
test_output[3661:3661] = '{32'hc6388b7e};
test_input[29296:29303] = '{32'hc23e1ac2, 32'hc15077e7, 32'h3f37c277, 32'hc0f4c3f5, 32'hc0220085, 32'hc2a93691, 32'h421f54bf, 32'hc20d0bef};
test_weights[29296:29303] = '{32'h4296ed29, 32'h42679ff7, 32'h42b343eb, 32'h41928263, 32'hbf01f27b, 32'h411a2006, 32'hc2bc9cbe, 32'h425af6f7};
test_bias[3662:3662] = '{32'hc2a95aca};
test_output[3662:3662] = '{32'hc62be748};
test_input[29304:29311] = '{32'hc165f0f5, 32'h41c0b452, 32'hc2b6574c, 32'h41a75f19, 32'h41e22477, 32'h42ba7f88, 32'hc15fc2c0, 32'h429f284f};
test_weights[29304:29311] = '{32'hc2782b8f, 32'hc0b76699, 32'h41bb1f4f, 32'h4227dcae, 32'hc2800dd9, 32'hc205c385, 32'h42873a14, 32'hc28ef267};
test_bias[3663:3663] = '{32'hc283d57b};
test_output[3663:3663] = '{32'hc63d81ca};
test_input[29312:29319] = '{32'hc256a04c, 32'hc143c183, 32'hc2a0859b, 32'hc24349a8, 32'h41eb185b, 32'hc108b094, 32'hc1edb274, 32'h4274974d};
test_weights[29312:29319] = '{32'hc21fa0af, 32'h421027a2, 32'hc26b2c2a, 32'h42b1dfc9, 32'hc1ccac4a, 32'h4212369c, 32'hc289682a, 32'hc2c6f96b};
test_bias[3664:3664] = '{32'hc24c0e20};
test_output[3664:3664] = '{32'hc54082a5};
test_input[29320:29327] = '{32'hc26a884d, 32'h416bc4dc, 32'hc262351a, 32'hc287b155, 32'h409b154c, 32'h4290d92d, 32'hc2562411, 32'hc2c6ea9d};
test_weights[29320:29327] = '{32'hc29d7c81, 32'hc1d44a9b, 32'h4296a390, 32'h42ba4775, 32'h42ac2cef, 32'h42c6f12f, 32'hc2a9abd7, 32'h428ffc9e};
test_bias[3665:3665] = '{32'h41d05d13};
test_output[3665:3665] = '{32'hc4a57f73};
test_input[29328:29335] = '{32'h41a3f335, 32'h429378a1, 32'hc2a64963, 32'h426558cc, 32'h417bd80b, 32'h420cf99f, 32'hc2b57b0b, 32'h428d6583};
test_weights[29328:29335] = '{32'hc22cc19b, 32'h427d3ee7, 32'hc001d8d0, 32'hc2373d39, 32'hc29c587d, 32'h427f7eac, 32'hc25645d6, 32'hc29cf7d1};
test_bias[3666:3666] = '{32'hc21ba380};
test_output[3666:3666] = '{32'h44ca6649};
test_input[29336:29343] = '{32'h42a1b8c7, 32'hc293c124, 32'hc29af947, 32'hc23e6907, 32'hc24d8dff, 32'h428435e2, 32'hc2c738f6, 32'h426d668d};
test_weights[29336:29343] = '{32'hc20be931, 32'h423339dd, 32'h42488b45, 32'hc2beb630, 32'hc1f6caf7, 32'hc232f55d, 32'hc2892ce9, 32'hc153e4e0};
test_bias[3667:3667] = '{32'hc2983a23};
test_output[3667:3667] = '{32'hc45d9c38};
test_input[29344:29351] = '{32'hc1b8334e, 32'hc1e5bc4b, 32'hc2848367, 32'hc1966fac, 32'hc10f9845, 32'h41629190, 32'h429ad089, 32'hc2a45e20};
test_weights[29344:29351] = '{32'hc2a1bf3c, 32'hc2438ced, 32'h406828ae, 32'h42bef395, 32'hbe74a2f9, 32'hc0e32fae, 32'h42176a40, 32'hc24146e1};
test_bias[3668:3668] = '{32'h427cb864};
test_output[3668:3668] = '{32'h45fd0271};
test_input[29352:29359] = '{32'hc2ac139f, 32'hc1aebeac, 32'h4136395b, 32'hc27d16f6, 32'hc2667d3b, 32'h426b8599, 32'h425880cb, 32'hc1925bc5};
test_weights[29352:29359] = '{32'hc21d8a21, 32'h42664a44, 32'h414961d3, 32'h420c1b12, 32'h4181b11b, 32'hc2702475, 32'h42936e33, 32'hc07bb2d5};
test_bias[3669:3669] = '{32'hc0d050d3};
test_output[3669:3669] = '{32'hc3b1c5f6};
test_input[29360:29367] = '{32'hc28b4410, 32'h426a4aa6, 32'h41b83047, 32'h41f7eb07, 32'hc1837caa, 32'h421a2f5e, 32'hc2a82275, 32'h42a0646d};
test_weights[29360:29367] = '{32'h425892c4, 32'hc29eb20f, 32'hc102ba31, 32'h4149bb62, 32'hc26e511e, 32'hc138d253, 32'h424f07d4, 32'h421812ed};
test_bias[3670:3670] = '{32'h420e694c};
test_output[3670:3670] = '{32'hc60bcf25};
test_input[29368:29375] = '{32'h41d77e11, 32'hc1a5e0b9, 32'h428559f9, 32'h42a61014, 32'hc0a2ee03, 32'hc2c366e2, 32'h42b04f6c, 32'hc1268f18};
test_weights[29368:29375] = '{32'hc28c5b65, 32'hc29baeb7, 32'h422847dc, 32'h42420b60, 32'hc20f2c4c, 32'h428e06f5, 32'h419f6772, 32'hc2bdaa9c};
test_bias[3671:3671] = '{32'h427deaab};
test_output[3671:3671] = '{32'h45230069};
test_input[29376:29383] = '{32'h427a4b2a, 32'h41978b94, 32'hc2123fbb, 32'hc1b4cde3, 32'hc1f64a11, 32'hc13f8efd, 32'h42299e2a, 32'h4283587c};
test_weights[29376:29383] = '{32'hc28a8953, 32'h429c10b9, 32'hc28706d3, 32'h4088836c, 32'hc23acb28, 32'hc2b159a1, 32'hc29b25af, 32'hc16740d4};
test_bias[3672:3672] = '{32'h4281df90};
test_output[3672:3672] = '{32'hc506e8aa};
test_input[29384:29391] = '{32'hc2809719, 32'hc22fe41b, 32'h42009423, 32'hc1e56738, 32'hc2bdf146, 32'hc2286269, 32'hbf161a49, 32'h40900e1f};
test_weights[29384:29391] = '{32'h4189ce87, 32'hc186fd97, 32'hc0c518d2, 32'h42507a2d, 32'h4258889a, 32'h4229e9f3, 32'hc270f765, 32'hc265df52};
test_bias[3673:3673] = '{32'h4183007b};
test_output[3673:3673] = '{32'hc60fa987};
test_input[29392:29399] = '{32'hc204c3db, 32'h421980b4, 32'h416c699a, 32'hc2a8e4b7, 32'h42abaf98, 32'h41e4c4e2, 32'hc2b40112, 32'hc2a6ea93};
test_weights[29392:29399] = '{32'hc15317cf, 32'hc2ab50d0, 32'h42ad11b6, 32'hc2b7288d, 32'hc2b6f3b5, 32'h4299126b, 32'hc28808a2, 32'h410ca9ce};
test_bias[3674:3674] = '{32'hbfbf5246};
test_output[3674:3674] = '{32'h45b7eb4d};
test_input[29400:29407] = '{32'h42453a37, 32'hc2151e33, 32'hc2837385, 32'h423b668d, 32'hc22fa805, 32'h418c166c, 32'hc2949a4f, 32'h42ba1796};
test_weights[29400:29407] = '{32'h40ed4199, 32'hc20323b6, 32'h420dff32, 32'h42c2bf45, 32'h420a0692, 32'hc2931ea0, 32'h42776a1a, 32'hc28a061e};
test_bias[3675:3675] = '{32'hc243ee1a};
test_output[3675:3675] = '{32'hc61d13de};
test_input[29408:29415] = '{32'hc207b11b, 32'h423ea59e, 32'hc24b7427, 32'h42845f73, 32'hc206ee42, 32'h41389028, 32'hc112cdd1, 32'h40a72817};
test_weights[29408:29415] = '{32'hc16ca5dc, 32'hc29f4618, 32'hc2ac147d, 32'hc2a71a79, 32'hc289e55b, 32'hc249310a, 32'h427f175e, 32'hc2bed648};
test_bias[3676:3676] = '{32'hc293d82c};
test_output[3676:3676] = '{32'hc57137a3};
test_input[29416:29423] = '{32'h419c5c04, 32'h412e88a3, 32'h42ac660c, 32'h427403d4, 32'h41d98677, 32'h42416d8d, 32'hc2b573e4, 32'h42170c5f};
test_weights[29416:29423] = '{32'h42b7cb2b, 32'hc262d338, 32'hc0eec4df, 32'hc2581f46, 32'hc1f22490, 32'hc150b2ca, 32'h42a4aa5b, 32'hc133d4b3};
test_bias[3677:3677] = '{32'h41ff88d0};
test_output[3677:3677] = '{32'hc63cb6bd};
test_input[29424:29431] = '{32'h42c1b7b6, 32'hc29d8e37, 32'hc1922c4f, 32'hc28848cc, 32'h428dc233, 32'hc21e1bf6, 32'hc1d45b0a, 32'h4224e597};
test_weights[29424:29431] = '{32'h420f0e7b, 32'hc2234e16, 32'h426a2b69, 32'hc18fb1f8, 32'h42038287, 32'h41804de9, 32'hc26da843, 32'hc2958ce7};
test_bias[3678:3678] = '{32'h429b3954};
test_output[3678:3678] = '{32'h45ddf92d};
test_input[29432:29439] = '{32'h40ae3de1, 32'hc1efbe97, 32'h4163d34a, 32'h420f7b54, 32'h4258ba7f, 32'hc13178cd, 32'hc1f10495, 32'h423c9414};
test_weights[29432:29439] = '{32'hc28c9770, 32'h41ae05a6, 32'h42c3ae15, 32'hc1f74fff, 32'hc1a2def5, 32'h42bbf51a, 32'h42061e2d, 32'hc2b630e7};
test_bias[3679:3679] = '{32'hc2176d37};
test_output[3679:3679] = '{32'hc600ba46};
test_input[29440:29447] = '{32'hc200ebde, 32'h4289c98e, 32'h41eef011, 32'h426e675a, 32'hc2492ecd, 32'h425a33d1, 32'h426a4a94, 32'h42b65375};
test_weights[29440:29447] = '{32'hc2b9f2f7, 32'h429fd742, 32'h4277f9b3, 32'hc1e76466, 32'hc113e0e0, 32'h4199f4f9, 32'hc293c4fa, 32'h42b8da90};
test_bias[3680:3680] = '{32'hc1c7e3f8};
test_output[3680:3680] = '{32'h465e28fa};
test_input[29448:29455] = '{32'h42c0def7, 32'h4088a520, 32'h420dbc43, 32'h428a4d94, 32'h42598883, 32'hc2753140, 32'hc2193ec8, 32'hc23a4e94};
test_weights[29448:29455] = '{32'h4255670e, 32'hc12053fb, 32'hc2a94565, 32'h4138fd54, 32'h418a0b7d, 32'hc2891515, 32'h42934f5e, 32'hc0073e61};
test_bias[3681:3681] = '{32'hc2823997};
test_output[3681:3681] = '{32'h45a43020};
test_input[29456:29463] = '{32'h41d74b8a, 32'h42b8e3f9, 32'hc1aa76d8, 32'h4290304b, 32'h420d3b5a, 32'h42c140db, 32'h421dadd4, 32'hc2c15c58};
test_weights[29456:29463] = '{32'hc27c0966, 32'h42242beb, 32'h42822105, 32'h4178991d, 32'h428aeb54, 32'h42808518, 32'h40a248cb, 32'h42983220};
test_bias[3682:3682] = '{32'hc2c1ffbb};
test_output[3682:3682] = '{32'h454a7bab};
test_input[29464:29471] = '{32'hc229b66e, 32'h4299af27, 32'hc1e8969a, 32'hc2a57210, 32'hc1920f15, 32'h4283ced7, 32'hc0e93c7c, 32'hc201e807};
test_weights[29464:29471] = '{32'h425d4a90, 32'hc26b9b6d, 32'hc29c7230, 32'h41af87cc, 32'hc16ed4bc, 32'h42c5a640, 32'h420f0afa, 32'h429b0074};
test_bias[3683:3683] = '{32'h42c6d7cc};
test_output[3683:3683] = '{32'hc5102eda};
test_input[29472:29479] = '{32'h3fe442e6, 32'hc1f4adb3, 32'hc2364f33, 32'hc20303f0, 32'h3fdf863e, 32'h429ff48d, 32'hc28c17a9, 32'h429b58a1};
test_weights[29472:29479] = '{32'hc1fe95c6, 32'hc2aca55e, 32'hc221a32d, 32'h428a8fac, 32'h42a526b2, 32'hc1ff8f10, 32'h41efdb57, 32'hc280bc70};
test_bias[3684:3684] = '{32'h4278f26b};
test_output[3684:3684] = '{32'hc5e3e225};
test_input[29480:29487] = '{32'hc2aacde7, 32'hc22c6a25, 32'h42b57f3b, 32'h4213ba9f, 32'h42b562a0, 32'h41a597af, 32'hc284306a, 32'h4297a856};
test_weights[29480:29487] = '{32'hc29e9bdf, 32'h4161b6da, 32'hc2a927a3, 32'hc27ae9bb, 32'hc131b28f, 32'hc1bc732b, 32'h42c63f7d, 32'h41d685b6};
test_bias[3685:3685] = '{32'hc290efae};
test_output[3685:3685] = '{32'hc61ae305};
test_input[29488:29495] = '{32'hc2565c1d, 32'h410bfb1f, 32'hc224159f, 32'h42b7d329, 32'h41ffacae, 32'h4272d042, 32'h4295b97b, 32'hc1be8d03};
test_weights[29488:29495] = '{32'hc05cb15a, 32'hc28fe7ba, 32'h42ae9d12, 32'hc209dc5f, 32'h42aaedf4, 32'h428558d1, 32'hc2ad05bd, 32'h42a8e6ae};
test_bias[3686:3686] = '{32'h425a909b};
test_output[3686:3686] = '{32'hc60a4205};
test_input[29496:29503] = '{32'h4276e519, 32'h42373701, 32'hc2861db7, 32'h410d7693, 32'hc2c7b91e, 32'h416627c7, 32'hc0f88e01, 32'hc280ff5a};
test_weights[29496:29503] = '{32'hc2243688, 32'h4118e100, 32'h413d726c, 32'hc24d1d14, 32'h42c63574, 32'hc238001f, 32'hc2c773cf, 32'hc1674e1e};
test_bias[3687:3687] = '{32'h41e7b4e1};
test_output[3687:3687] = '{32'hc63e1864};
test_input[29504:29511] = '{32'h42968271, 32'h42c6e7ae, 32'h429925ec, 32'h42afcddb, 32'h426059cf, 32'hc249efb3, 32'hc1e98bb0, 32'h41cb04c9};
test_weights[29504:29511] = '{32'h42506eef, 32'h421c562e, 32'h4199c8f3, 32'h42a67135, 32'h40f26ebd, 32'h426b7365, 32'hc2aacd36, 32'hc2a317da};
test_bias[3688:3688] = '{32'hc1df6328};
test_output[3688:3688] = '{32'h4661b31a};
test_input[29512:29519] = '{32'h421ad62d, 32'hc09be177, 32'h418d7076, 32'h42899a05, 32'h41ad7b91, 32'h423ad6f5, 32'h410c8d01, 32'hc23a5d59};
test_weights[29512:29519] = '{32'h4188ce9c, 32'h422c2b72, 32'hc1d116a1, 32'hc1e97d98, 32'h3f872a91, 32'hc26f892a, 32'hc1a257fc, 32'h42b1bc48};
test_bias[3689:3689] = '{32'hc27f2c9a};
test_output[3689:3689] = '{32'hc60f5a79};
test_input[29520:29527] = '{32'hc132bfb2, 32'hc1c98a6e, 32'hc1541616, 32'hc2ac410c, 32'hc2791802, 32'hc1bed355, 32'hc263c723, 32'hc1a48ca4};
test_weights[29520:29527] = '{32'h429ff603, 32'hc0dcef8c, 32'h428da728, 32'h42b43146, 32'hc2225495, 32'h40717b19, 32'h4218a698, 32'hc0b50817};
test_bias[3690:3690] = '{32'hc29545c7};
test_output[3690:3690] = '{32'hc60e616e};
test_input[29528:29535] = '{32'hc2188813, 32'h4281c7b5, 32'h425248c8, 32'h42c2d59b, 32'h41318e2c, 32'hc27c1f4f, 32'hc29b01a6, 32'h41efde14};
test_weights[29528:29535] = '{32'hc28deeb1, 32'hc2996110, 32'hc291ae37, 32'hc289bf0d, 32'hbf590e2a, 32'hc177fd5b, 32'hc2547ad1, 32'hc2baae53};
test_bias[3691:3691] = '{32'h423cda2a};
test_output[3691:3691] = '{32'hc623afb8};
test_input[29536:29543] = '{32'h41220527, 32'hc164013e, 32'h42a104a1, 32'hc0860510, 32'hc24f7bd0, 32'h425d75bc, 32'h42829c86, 32'h4224c6ee};
test_weights[29536:29543] = '{32'hc252d753, 32'hc1d54851, 32'h41a21416, 32'h4290ecaf, 32'h42542e3b, 32'h42b5c37f, 32'h42a0867a, 32'h42240edd};
test_bias[3692:3692] = '{32'hc2a35885};
test_output[3692:3692] = '{32'h4620fdc9};
test_input[29544:29551] = '{32'h4275f810, 32'h42196db5, 32'h42b80b5e, 32'h41eb49bf, 32'hc291c149, 32'h4294e731, 32'h42c1cc58, 32'h4257d6e0};
test_weights[29544:29551] = '{32'h42af7462, 32'h42a5cc87, 32'hc20b420f, 32'hc2b5e9c8, 32'h42a2209f, 32'hc1fdef24, 32'h429d981a, 32'h42678236};
test_bias[3693:3693] = '{32'h421b3946};
test_output[3693:3693] = '{32'h45a32e29};
test_input[29552:29559] = '{32'h42c2cdda, 32'hc2450514, 32'h4212491f, 32'hc1a4d89f, 32'h42b04750, 32'h42c475fe, 32'hc2662936, 32'h42bf10da};
test_weights[29552:29559] = '{32'hc23ea314, 32'hc237071a, 32'h41a89040, 32'h42124437, 32'hc265a331, 32'hc1d8a7d6, 32'h428e0228, 32'h42a540d3};
test_bias[3694:3694] = '{32'h4285e255};
test_output[3694:3694] = '{32'hc5c24535};
test_input[29560:29567] = '{32'hc23d2327, 32'h420a4c78, 32'h41da1891, 32'hc1917139, 32'h42b04eb2, 32'hc0a0e17d, 32'hc2ac232a, 32'hc1ab9e20};
test_weights[29560:29567] = '{32'hc24ebf2c, 32'h4273e9b6, 32'h42832399, 32'hc2638624, 32'h42bde426, 32'h42885b5f, 32'hc1e69c15, 32'hc20a3e27};
test_bias[3695:3695] = '{32'h42b0abaa};
test_output[3695:3695] = '{32'h46922f81};
test_input[29568:29575] = '{32'h4295a184, 32'h428af42b, 32'h423246e5, 32'hc2a38446, 32'hc23c1340, 32'h3efe99e5, 32'hc20ff29a, 32'h42baf78c};
test_weights[29568:29575] = '{32'h4133a859, 32'hc108aa11, 32'h42a8b158, 32'hc18d9de7, 32'hc1fa108a, 32'hc26ba63c, 32'h42b78eb1, 32'h4260de52};
test_bias[3696:3696] = '{32'hc007ebe9};
test_output[3696:3696] = '{32'h460a3015};
test_input[29576:29583] = '{32'h41ff640e, 32'hc2ab0310, 32'hc258aa3d, 32'hc18b95f0, 32'hc29982ff, 32'hc1c9a7c0, 32'hc0ac317d, 32'h428fee0d};
test_weights[29576:29583] = '{32'h429c227b, 32'hc1e1d1d8, 32'hc217a23b, 32'h415f643a, 32'h3fed273a, 32'hc22802e0, 32'h4094bcd7, 32'h429500d0};
test_bias[3697:3697] = '{32'h429113fc};
test_output[3697:3697] = '{32'h464bc49e};
test_input[29584:29591] = '{32'hc2a4cc36, 32'hc17e07d7, 32'hc1acb07f, 32'h4290c051, 32'hc1a9d5cc, 32'hc2930ce9, 32'h4154c01d, 32'hc1dd6805};
test_weights[29584:29591] = '{32'h42b31624, 32'hc24bbc1e, 32'hc2b3d8fa, 32'h42536f78, 32'hc2a08dc8, 32'hc2a1f7cd, 32'hc2b2827c, 32'h419e98c3};
test_bias[3698:3698] = '{32'h420ddd8a};
test_output[3698:3698] = '{32'h45a11e67};
test_input[29592:29599] = '{32'h41892d96, 32'hc0e0b2a1, 32'h42970d2a, 32'hc0c79e5f, 32'h42ab9e5f, 32'hc201da39, 32'hc26aab6a, 32'h40acc3a7};
test_weights[29592:29599] = '{32'hc12695de, 32'hc19fef5b, 32'h42826cbe, 32'h41b55d2a, 32'hc2a0c31c, 32'h42557925, 32'hc202127e, 32'h3f15ae5e};
test_bias[3699:3699] = '{32'hc2b98dad};
test_output[3699:3699] = '{32'hc50122d0};
test_input[29600:29607] = '{32'hc0bb110a, 32'hc2923f3b, 32'h42b9bf84, 32'h42b91540, 32'h41a87c20, 32'hc222b154, 32'hc203258a, 32'hc279ca9c};
test_weights[29600:29607] = '{32'hc295af6e, 32'h42c3b856, 32'hc23cc9ac, 32'h42c55c08, 32'h41c7565f, 32'hc2588f92, 32'h42ab963e, 32'h421ffff5};
test_bias[3700:3700] = '{32'h42b8cda9};
test_output[3700:3700] = '{32'hc58b6a85};
test_input[29608:29615] = '{32'h41774e83, 32'hc1d88e67, 32'hc2a7f896, 32'h427d9edf, 32'hc2bcf525, 32'hc29a95d4, 32'hc135ec7f, 32'hc2bd2b9e};
test_weights[29608:29615] = '{32'hc1bae119, 32'h42075f70, 32'hc23ae82e, 32'h425d4006, 32'h4047bd51, 32'h428b6aed, 32'h42522b3b, 32'h4292ada9};
test_bias[3701:3701] = '{32'hc2477bb4};
test_output[3701:3701] = '{32'hc5de452e};
test_input[29616:29623] = '{32'h42033071, 32'h41f9470c, 32'hc28e2747, 32'h42c40ea2, 32'hc194ccda, 32'hc0c33df5, 32'h414080ca, 32'hc2911bb8};
test_weights[29616:29623] = '{32'hc0da3f4e, 32'hc2a4052f, 32'hc26dcc5b, 32'h42474d80, 32'hc25b37c7, 32'h422334ba, 32'h4145b834, 32'h425d5220};
test_bias[3702:3702] = '{32'hc1331270};
test_output[3702:3702] = '{32'h4549832d};
test_input[29624:29631] = '{32'h421a931e, 32'h41034048, 32'hc1ef9746, 32'hc271c627, 32'h4291c442, 32'h42633bef, 32'hc28c7b57, 32'h41a81175};
test_weights[29624:29631] = '{32'hc2a97518, 32'hc2714a52, 32'h422750e2, 32'hc2371add, 32'h426c37af, 32'h4170efd6, 32'h40a04590, 32'h412015c8};
test_bias[3703:3703] = '{32'h428558fb};
test_output[3703:3703] = '{32'h4530daed};
test_input[29632:29639] = '{32'h421a909b, 32'hc28042bd, 32'hc2547a3b, 32'h42b6abed, 32'h4136e16a, 32'hc2894cba, 32'h4157c845, 32'h42b285bb};
test_weights[29632:29639] = '{32'hc2a4b4d3, 32'hc2661e13, 32'h4278d0ec, 32'h41dcbc0e, 32'hc0648732, 32'h428a91b1, 32'hc1a8cdc8, 32'hc0b155b9};
test_bias[3704:3704] = '{32'h42280b89};
test_output[3704:3704] = '{32'hc5b59afb};
test_input[29640:29647] = '{32'h41c0b2a3, 32'h4286f37c, 32'hc21e693a, 32'hc2c22daf, 32'h42219175, 32'h428857aa, 32'h4289bd6f, 32'hc1fff2ef};
test_weights[29640:29647] = '{32'hc22134e8, 32'h40e7ec58, 32'h41d62415, 32'h42b3788d, 32'hc1a1b08e, 32'hc256586a, 32'h4189cdb6, 32'h4286871c};
test_bias[3705:3705] = '{32'hc2a287d4};
test_output[3705:3705] = '{32'hc6766a14};
test_input[29648:29655] = '{32'hc27a4a6d, 32'hc2239245, 32'hc2521c0d, 32'hc20ec536, 32'h418c9321, 32'h42569410, 32'h411d5327, 32'h42830fdb};
test_weights[29648:29655] = '{32'h41519b87, 32'hc20fcdc7, 32'h415527ec, 32'h42494c05, 32'hc2861989, 32'h41934f61, 32'hc2a60d2c, 32'hc2890929};
test_bias[3706:3706] = '{32'hc1cb9e1a};
test_output[3706:3706] = '{32'hc5e63ebe};
test_input[29656:29663] = '{32'hc28d6352, 32'h408ea9b4, 32'hbf4138aa, 32'hc2862b12, 32'h41f3a0dc, 32'h42187e32, 32'hc19b1ff3, 32'h42be6a02};
test_weights[29656:29663] = '{32'h42a1e94d, 32'h423d644b, 32'h41e69563, 32'hc299e3b8, 32'hc2b47851, 32'h426e4df6, 32'hc1b5fb89, 32'h4187ea04};
test_bias[3707:3707] = '{32'h42c6f628};
test_output[3707:3707] = '{32'h44a3ab77};
test_input[29664:29671] = '{32'hc120ea09, 32'hc2a35de9, 32'h41bace88, 32'hc26c0aa0, 32'hc2bcf9b3, 32'h42214ebb, 32'h422fde9a, 32'hc29c2c94};
test_weights[29664:29671] = '{32'hc2402b3d, 32'h4291dded, 32'hc14fb51b, 32'hc2958b31, 32'h4290f160, 32'hc1dc8f50, 32'h427d66ff, 32'hc2b69935};
test_bias[3708:3708] = '{32'hc2896f6a};
test_output[3708:3708] = '{32'h440256cd};
test_input[29672:29679] = '{32'h420b6c31, 32'h42a7956f, 32'hc2ac24b0, 32'h42c15c43, 32'hc2b23b7c, 32'h424f54c4, 32'h41a51145, 32'hc111f0b2};
test_weights[29672:29679] = '{32'h42c16dc6, 32'h42216b62, 32'hc25343bd, 32'hc0fb34c5, 32'hc22d1ad7, 32'h4297e82e, 32'hc23e1a92, 32'h42c4569a};
test_bias[3709:3709] = '{32'hc2050a8a};
test_output[3709:3709] = '{32'h46804f4c};
test_input[29680:29687] = '{32'h419f8831, 32'h419dfe4b, 32'h41d6796a, 32'hc2a8b366, 32'hc154fb5c, 32'hc28f9412, 32'h41613657, 32'hc2855b40};
test_weights[29680:29687] = '{32'h42a6c6ba, 32'h41a408ca, 32'hc231c83f, 32'h42ab0b62, 32'h42c6e7d7, 32'hc1de0621, 32'h41b53622, 32'h428bb6f3};
test_bias[3710:3710] = '{32'h429035c1};
test_output[3710:3710] = '{32'hc61b4046};
test_input[29688:29695] = '{32'hc26b29b4, 32'hbe7ec86c, 32'hc2a92fc4, 32'hc2855259, 32'h42220d35, 32'hc225023b, 32'h42be9440, 32'hc093e92c};
test_weights[29688:29695] = '{32'hc2ae35c8, 32'h429151f4, 32'h41b2856d, 32'h428d45b4, 32'h414d7785, 32'hc2b07b0a, 32'h4219a58d, 32'hc2017d35};
test_bias[3711:3711] = '{32'h4248518b};
test_output[3711:3711] = '{32'h45cbf684};
test_input[29696:29703] = '{32'h41b4c0ef, 32'h4239ae1d, 32'hc20080d2, 32'h41589704, 32'h4282e24d, 32'hc1f7acf9, 32'hc21b4310, 32'h42890843};
test_weights[29696:29703] = '{32'h4092f398, 32'h42c412ac, 32'hc182a9b1, 32'hc2947273, 32'hc2c5254c, 32'h42207e01, 32'hc192f37f, 32'hc1a01616};
test_bias[3712:3712] = '{32'h423b3f8d};
test_output[3712:3712] = '{32'hc5810d6d};
test_input[29704:29711] = '{32'h4251db27, 32'h422110c4, 32'hc14f2f2f, 32'h4184da33, 32'h3fc3ce4e, 32'hc2992893, 32'h42c5a1e8, 32'hc228fbaa};
test_weights[29704:29711] = '{32'h4187f640, 32'h42744e66, 32'hc26ce123, 32'hc2b0cb24, 32'hc27b493b, 32'h4209bc54, 32'hc2b5f4eb, 32'hc27394fa};
test_bias[3713:3713] = '{32'hc209cda8};
test_output[3713:3713] = '{32'hc5cc3986};
test_input[29712:29719] = '{32'h4239fa77, 32'h42385a43, 32'hc00fab05, 32'h41a39331, 32'h42b4b79e, 32'hc190ffc5, 32'h42b67c3f, 32'h42b4f52a};
test_weights[29712:29719] = '{32'h42a650eb, 32'h42589b02, 32'hc2ba388e, 32'hc2c01379, 32'hc25605db, 32'hc2943f33, 32'hc2879e0b, 32'hc21d8e86};
test_bias[3714:3714] = '{32'hc279c7dc};
test_output[3714:3714] = '{32'hc607e482};
test_input[29720:29727] = '{32'hc293418f, 32'h42a94d5d, 32'h4230fedf, 32'hc2bff069, 32'h42c4168c, 32'h416679f8, 32'hc2675526, 32'h41eff86a};
test_weights[29720:29727] = '{32'h42c4bcc4, 32'h427892e0, 32'hc2c265f2, 32'hc28fb345, 32'h408564fa, 32'hc1807bac, 32'h425be6cf, 32'h428ad3f9};
test_bias[3715:3715] = '{32'h417648d1};
test_output[3715:3715] = '{32'hc392196b};
test_input[29728:29735] = '{32'h42781d7a, 32'hc191d269, 32'hc22a58b2, 32'hc2892752, 32'hc253b9bb, 32'hc234d3ef, 32'hc29d714b, 32'h42187618};
test_weights[29728:29735] = '{32'hc2b6489b, 32'hc22118da, 32'h408f0978, 32'h411bc875, 32'h42573444, 32'hc23d0f30, 32'hc0038687, 32'h42abb97a};
test_bias[3716:3716] = '{32'hc2a5ce1a};
test_output[3716:3716] = '{32'hc5440e0b};
test_input[29736:29743] = '{32'h4279f57a, 32'hc28c3d67, 32'h42861170, 32'hc293ee99, 32'hc29eb2f9, 32'hbf11d066, 32'hc26f73fe, 32'hc227dc86};
test_weights[29736:29743] = '{32'hc28a3a3b, 32'h426031af, 32'hc0dfb88b, 32'h42c433c0, 32'hc25bb111, 32'h42c039b7, 32'hc0ba1175, 32'h4261e558};
test_bias[3717:3717] = '{32'hc106813b};
test_output[3717:3717] = '{32'hc65612e5};
test_input[29744:29751] = '{32'hc2b24de5, 32'hc1de73d1, 32'hc0b72949, 32'h429ea0e5, 32'hc28ac398, 32'hc1b52979, 32'hc26b1377, 32'hc1d0a277};
test_weights[29744:29751] = '{32'hc11037df, 32'h42bf5bab, 32'hc23f9c64, 32'h4274fd42, 32'hc262ebca, 32'h426b28e3, 32'hc2068bbc, 32'h3e02c3ad};
test_bias[3718:3718] = '{32'hc01f6ca1};
test_output[3718:3718] = '{32'h45f55612};
test_input[29752:29759] = '{32'hc2248bae, 32'h41b52658, 32'h4279fe24, 32'h4196116f, 32'hc20d8103, 32'hc2475f1b, 32'hc20d27b3, 32'h4236da9d};
test_weights[29752:29759] = '{32'hc2637f38, 32'h416dcf2d, 32'h4245d3ac, 32'h429303f8, 32'hc2369218, 32'hc24d3174, 32'hc2ac3417, 32'h427d2258};
test_bias[3719:3719] = '{32'hc22b925b};
test_output[3719:3719] = '{32'h46866beb};
test_input[29760:29767] = '{32'h4219ce66, 32'hc2a7d152, 32'h428d7373, 32'hc2c72b8e, 32'hc1d9cfed, 32'h42388f29, 32'h4245b508, 32'h41a92662};
test_weights[29760:29767] = '{32'hc10331cc, 32'hc11a996a, 32'h427aec37, 32'h42391f3c, 32'h4260033e, 32'hbff2715d, 32'hc265dee0, 32'hc1e8f7e4};
test_bias[3720:3720] = '{32'hc28fd61c};
test_output[3720:3720] = '{32'hc59687b9};
test_input[29768:29775] = '{32'hc1d7c12e, 32'h42972203, 32'hc2b40db0, 32'hc0d65399, 32'h422ee08b, 32'h4049d9f6, 32'hc150c703, 32'hc22dbfc2};
test_weights[29768:29775] = '{32'hc2924216, 32'h4233f323, 32'h4139a2c1, 32'h426874c9, 32'hc15d8c27, 32'hc1d0170f, 32'hc24ed941, 32'hc297bde3};
test_bias[3721:3721] = '{32'h4109f9c2};
test_output[3721:3721] = '{32'h45e1ed35};
test_input[29776:29783] = '{32'hc1efbe5e, 32'hc29835a3, 32'h413e6f6a, 32'h424dd2db, 32'h41c2e156, 32'hc23b7663, 32'hc280afac, 32'h42ad2925};
test_weights[29776:29783] = '{32'h42be657e, 32'hc23e2b03, 32'hc11f232e, 32'h41092852, 32'h4265be42, 32'h429121f3, 32'hc01ef867, 32'hc231d319};
test_bias[3722:3722] = '{32'hc194395d};
test_output[3722:3722] = '{32'hc5906bbd};
test_input[29784:29791] = '{32'h4284ea12, 32'hc1b32e4e, 32'hc299b970, 32'hc2a348c7, 32'hc181eb1a, 32'hc28dc7f1, 32'h40d6dd2d, 32'h41b3ddd6};
test_weights[29784:29791] = '{32'h4158c611, 32'hc2bc842a, 32'h4207c89d, 32'hc291c539, 32'hc2004ddd, 32'hc2727824, 32'h421b2906, 32'hc291dd35};
test_bias[3723:3723] = '{32'hc2305007};
test_output[3723:3723] = '{32'h46184e75};
test_input[29792:29799] = '{32'hc268e2e5, 32'h42b4f3b3, 32'hc2ba0292, 32'h41cea2ae, 32'h42284c20, 32'h42434928, 32'hbd062bf5, 32'hc22209fc};
test_weights[29792:29799] = '{32'hc1c79bc4, 32'h42a5320a, 32'hc18fc77b, 32'hc2c4f5e0, 32'hc2836138, 32'hc25a3ca3, 32'h42b0f12b, 32'h42890832};
test_bias[3724:3724] = '{32'h428b89b5};
test_output[3724:3724] = '{32'hc2a527eb};
test_input[29800:29807] = '{32'hc1d14b0d, 32'hc0cbbd32, 32'hc1ffd223, 32'hc23f1e39, 32'hc1f159c9, 32'h42b98d61, 32'h42a20830, 32'h428430fb};
test_weights[29800:29807] = '{32'hc2bcaa37, 32'h4180d169, 32'h42be3822, 32'hc27d8391, 32'h4041497b, 32'hc2a37f2d, 32'h426b1452, 32'h41f8c45d};
test_bias[3725:3725] = '{32'hc2583f63};
test_output[3725:3725] = '{32'h44b3e9fb};
test_input[29808:29815] = '{32'h42957316, 32'hc2163ba3, 32'hc18701c5, 32'hc2b8e0f8, 32'hc28a03b8, 32'hc1fb02af, 32'h41eb4589, 32'h409bb469};
test_weights[29808:29815] = '{32'hc2bf88b8, 32'h42b72a9b, 32'hc2b5e3b2, 32'hc1b7ad54, 32'h40a8f718, 32'h42bf2349, 32'hc293f6fb, 32'hc2537445};
test_bias[3726:3726] = '{32'hc2c3dc59};
test_output[3726:3726] = '{32'hc6488262};
test_input[29816:29823] = '{32'h42beaef9, 32'h429c8bf8, 32'hc248a134, 32'hc2364274, 32'h42555834, 32'h41b49576, 32'hc2c5144b, 32'hc287f762};
test_weights[29816:29823] = '{32'h422608e1, 32'h42a8b282, 32'hc2c3caf7, 32'h422c28ed, 32'h42870ca7, 32'h42a51db1, 32'hc13869f0, 32'hc27315b5};
test_bias[3727:3727] = '{32'hc226c7bf};
test_output[3727:3727] = '{32'h46bd0ee5};
test_input[29824:29831] = '{32'hc24314c6, 32'h429c817c, 32'hc22d35fa, 32'h41bb30d3, 32'hc2c1c54d, 32'h425831da, 32'hc21852f4, 32'hc07fa62a};
test_weights[29824:29831] = '{32'h42a9a3cc, 32'h417dcceb, 32'h419863db, 32'h42940e2a, 32'h423ab2d5, 32'hc239fb64, 32'hc1c72a32, 32'hc2465697};
test_bias[3728:3728] = '{32'hc2a35dff};
test_output[3728:3728] = '{32'hc5f8b63f};
test_input[29832:29839] = '{32'h42a59ab0, 32'hc23dcb9d, 32'h4127a17a, 32'h425fc82d, 32'h42157a2f, 32'hc280e540, 32'h42ae0e95, 32'hc2ae26ea};
test_weights[29832:29839] = '{32'h42b72149, 32'h419b9afd, 32'hc1fcee53, 32'h4172ae76, 32'hc2915dde, 32'hc27a42b2, 32'hc2a180b2, 32'h42af8095};
test_bias[3729:3729] = '{32'h41b0b70a};
test_output[3729:3729] = '{32'hc5c052e1};
test_input[29840:29847] = '{32'h42829a1f, 32'hc1b491fa, 32'h42a99f56, 32'h40a7f01a, 32'hc1b63818, 32'hc1cc18b6, 32'h42723010, 32'hc235cb58};
test_weights[29840:29847] = '{32'hc2b43ecf, 32'h41ae6b4c, 32'hc285a138, 32'h4205150f, 32'h40ac8d6c, 32'hc2ad59ee, 32'h41ae464a, 32'hc20724b6};
test_bias[3730:3730] = '{32'h42a4bee5};
test_output[3730:3730] = '{32'hc5d5df7d};
test_input[29848:29855] = '{32'hc2c25f79, 32'hc1c45a86, 32'hc298459b, 32'h42775536, 32'h419f89de, 32'h3ed71176, 32'hc250ad43, 32'h42ae18d8};
test_weights[29848:29855] = '{32'hc29f192f, 32'h4140f7a1, 32'h4208041d, 32'hc1898850, 32'hc1af1581, 32'h3f0c98f1, 32'hc29ac73f, 32'h428a7cca};
test_bias[3731:3731] = '{32'hc22bc2f5};
test_output[3731:3731] = '{32'h4650e38f};
test_input[29856:29863] = '{32'h4165529a, 32'hc1e553b2, 32'h428358b9, 32'h418fae3a, 32'hc2834612, 32'hc26c35be, 32'hc021cb5f, 32'hc2678cc5};
test_weights[29856:29863] = '{32'h420c0e9f, 32'hc2b11b2b, 32'h414d4573, 32'hc2c6442c, 32'hc23fd2b2, 32'h427608cd, 32'h421fa27d, 32'h40fbb4cf};
test_bias[3732:3732] = '{32'h42328fbe};
test_output[3732:3732] = '{32'h448a484d};
test_input[29864:29871] = '{32'h4145deee, 32'hc2aeeb74, 32'h429edc2d, 32'h42ac84f1, 32'h4244e7d6, 32'h41f4fca5, 32'hc2189508, 32'hc23bb9ff};
test_weights[29864:29871] = '{32'hc2bb1da9, 32'hc2c1ddce, 32'h41616211, 32'hc147471b, 32'hc289c30e, 32'h424bcc41, 32'hc2a3de3c, 32'hc2660c8d};
test_bias[3733:3733] = '{32'h40afafac};
test_output[3733:3733] = '{32'h4631933f};
test_input[29872:29879] = '{32'hc21426ab, 32'h4280653d, 32'h42023ea2, 32'hc255221c, 32'hc1a633fe, 32'hc17ae634, 32'hc0d4748a, 32'h40a7857e};
test_weights[29872:29879] = '{32'h426a29f6, 32'hc2c20b79, 32'hc14c52e5, 32'h429309f3, 32'hc2a7b8bf, 32'hc2bdcbb6, 32'hc2a12e09, 32'hc1355751};
test_bias[3734:3734] = '{32'hc094a894};
test_output[3734:3734] = '{32'hc60d125a};
test_input[29880:29887] = '{32'hc1cd6d9b, 32'hc235acab, 32'hc2adddbc, 32'h4294f8cf, 32'hc117b3f5, 32'hc2813a30, 32'h4267d2ef, 32'hc2c5d899};
test_weights[29880:29887] = '{32'h415ff203, 32'h429d858d, 32'hc2837a2b, 32'h41a88195, 32'hc2a91514, 32'h428b7f4d, 32'hc2b1bb23, 32'hc1e26f21};
test_bias[3735:3735] = '{32'h424c030d};
test_output[3735:3735] = '{32'hc5261538};
test_input[29888:29895] = '{32'h42497100, 32'hc2409513, 32'h42ac422e, 32'h4212f100, 32'hc2c36739, 32'h4001afcd, 32'hc2a5733c, 32'h424fa6b7};
test_weights[29888:29895] = '{32'hc1746e10, 32'h4287a6a0, 32'h42503d62, 32'h4219c57a, 32'hc13401df, 32'h4232142e, 32'h41cd8040, 32'hc2b20dcb};
test_bias[3736:3736] = '{32'h42a2349b};
test_output[3736:3736] = '{32'hc561ee4c};
test_input[29896:29903] = '{32'h420f60ef, 32'hc2943b34, 32'h41bf78b3, 32'h427c4a28, 32'h412a303f, 32'h42096a2b, 32'hc1b7bee6, 32'hc26b36cd};
test_weights[29896:29903] = '{32'hc27870e7, 32'hc25a35da, 32'hc27c6b26, 32'hc2a7c3f7, 32'hc21ab653, 32'hc0a7b55f, 32'h42289481, 32'hc2acfebe};
test_bias[3737:3737] = '{32'hc2b1f6aa};
test_output[3737:3737] = '{32'hc4c14720};
test_input[29904:29911] = '{32'h42c21fbd, 32'h41e4a0e4, 32'hc06dee5b, 32'hc0115ff9, 32'h417ea337, 32'h4211bfdb, 32'h41025a05, 32'hc12e2c77};
test_weights[29904:29911] = '{32'hc27a3c1c, 32'h42af2f4e, 32'h426ba113, 32'hc2b469c6, 32'h42b19ffa, 32'h42275d61, 32'hc2b2dea2, 32'h41ec53de};
test_bias[3738:3738] = '{32'hc19fa58b};
test_output[3738:3738] = '{32'hc4d66157};
test_input[29912:29919] = '{32'h42a74537, 32'h424a0b0c, 32'h42a2290d, 32'hc0802035, 32'h419fbaaf, 32'h427d2865, 32'h41f17c3b, 32'hc2acfb98};
test_weights[29912:29919] = '{32'hc21d3b3d, 32'hc20dee3b, 32'hc1706ceb, 32'hc0bc8e52, 32'h41d4a9a8, 32'hc17fbf49, 32'h42b85be3, 32'hc2c4b8db};
test_bias[3739:3739] = '{32'hc22fa083};
test_output[3739:3739] = '{32'h458c547a};
test_input[29920:29927] = '{32'h4285d937, 32'hc00ab757, 32'h421dfbf4, 32'hc26f96ae, 32'hc28b7ecb, 32'hc254f924, 32'h423428be, 32'hc267a4dc};
test_weights[29920:29927] = '{32'hc1f53f78, 32'hc121e434, 32'hc2626911, 32'h42b12879, 32'hc28dc756, 32'h4210a759, 32'hc2810f04, 32'h416d8fd4};
test_bias[3740:3740] = '{32'hc1b2baf6};
test_output[3740:3740] = '{32'hc621924d};
test_input[29928:29935] = '{32'hc229ce5d, 32'hc2c19f19, 32'h41e3ec5c, 32'h42821510, 32'h420a69ed, 32'hc01eec1d, 32'h42210a65, 32'h41c01cb2};
test_weights[29928:29935] = '{32'hc0d8c18a, 32'h4279af8f, 32'h428b95f1, 32'h429fdb32, 32'h412de049, 32'hc2997931, 32'hc288c3ea, 32'h42431838};
test_bias[3741:3741] = '{32'h41d90c10};
test_output[3741:3741] = '{32'h43ddb429};
test_input[29936:29943] = '{32'hc09f208f, 32'h4296ab9a, 32'hc218fdfe, 32'hc261a193, 32'h429e561c, 32'hc295efeb, 32'h41bc8593, 32'hc2c7af07};
test_weights[29936:29943] = '{32'h41e7a93c, 32'h417e9fee, 32'h42abdf38, 32'h42b99022, 32'hc25b599d, 32'hc14aaae9, 32'h42136677, 32'hc2804d30};
test_bias[3742:3742] = '{32'h426926d5};
test_output[3742:3742] = '{32'hc55c5c63};
test_input[29944:29951] = '{32'h41b506d6, 32'hc22f03f6, 32'h40f1fc13, 32'h412db70e, 32'hc297dbd6, 32'hc173078a, 32'h42bfb517, 32'hc2a1a315};
test_weights[29944:29951] = '{32'hc1d211e3, 32'hc0d6b202, 32'h41de4e05, 32'h42a6abf3, 32'hc1ca532d, 32'hc29a1ea9, 32'hc1b51637, 32'h4223c333};
test_bias[3743:3743] = '{32'h4280a1e6};
test_output[3743:3743] = '{32'hc4bca304};
test_input[29952:29959] = '{32'h42a0b072, 32'hc1d9ef78, 32'h42416132, 32'h42a4c525, 32'hc230b338, 32'hc1f9359d, 32'hc13bb438, 32'h41aa7f51};
test_weights[29952:29959] = '{32'h42146dcc, 32'h4295d189, 32'hc2bf5494, 32'h4279afec, 32'hc2c143b0, 32'h425b113d, 32'hc24ce1cd, 32'h4166bc46};
test_bias[3744:3744] = '{32'h4198ca04};
test_output[3744:3744] = '{32'h459aa339};
test_input[29960:29967] = '{32'hc23a0dd9, 32'hc2820cc7, 32'hc25a8fd7, 32'h42853e3d, 32'h42979d74, 32'h42995679, 32'h420f2236, 32'hc1212014};
test_weights[29960:29967] = '{32'h4213eefe, 32'h4287b80b, 32'h428e6d61, 32'h42a2c68f, 32'hc2bba7e9, 32'h4147c908, 32'h42b6f238, 32'hc2ace374};
test_bias[3745:3745] = '{32'hc1e54798};
test_output[3745:3745] = '{32'hc5cf919b};
test_input[29968:29975] = '{32'h3f2504bd, 32'hc28764da, 32'hc28c4997, 32'h428d53c0, 32'h41bae33d, 32'h4293645e, 32'hc2a6b35e, 32'hc28edeb2};
test_weights[29968:29975] = '{32'hc1238cf6, 32'h42140123, 32'h404d0a71, 32'h410d50cb, 32'h41a695b6, 32'h429f53e0, 32'h4213121c, 32'hc28befe8};
test_bias[3746:3746] = '{32'hc29b9382};
test_output[3746:3746] = '{32'h45bea8df};
test_input[29976:29983] = '{32'hc2a88228, 32'h42a09cd9, 32'hc26d6c5f, 32'hc29b3748, 32'h417b90d9, 32'hc28f0c91, 32'h42603ec1, 32'h4136c844};
test_weights[29976:29983] = '{32'hc1f2b5f1, 32'h41a9e521, 32'h41f7f922, 32'h41ce4f7f, 32'h429d068c, 32'hc1e0cacd, 32'h42a6f335, 32'hc25210e6};
test_bias[3747:3747] = '{32'hc297289a};
test_output[3747:3747] = '{32'h45efa655};
test_input[29984:29991] = '{32'hc1936853, 32'hc2009ef1, 32'h414cc88b, 32'hc23e3ba2, 32'h42b0ab88, 32'hc2bd82e3, 32'h428a5334, 32'hc1e30b82};
test_weights[29984:29991] = '{32'h420f3c37, 32'h426fc235, 32'hc1e63f49, 32'hc23ff2ad, 32'h423f4ad7, 32'hc28aa9a9, 32'h41f2fb59, 32'h41686916};
test_bias[3748:3748] = '{32'h42a3672b};
test_output[3748:3748] = '{32'h4639cae8};
test_input[29992:29999] = '{32'hc023138e, 32'hc180f0a0, 32'hc282c496, 32'hc2671dc9, 32'h428b6a1b, 32'h425723c3, 32'hc222b976, 32'h420013e7};
test_weights[29992:29999] = '{32'h412a787b, 32'h428600bf, 32'h41b6b915, 32'hc18bba2f, 32'hc1f8aec5, 32'hc20c9fc3, 32'h419b2a2c, 32'hc2c2c76c};
test_bias[3749:3749] = '{32'h422ad8b2};
test_output[3749:3749] = '{32'hc614a6c2};
test_input[30000:30007] = '{32'h4288f8c8, 32'h4208d554, 32'hc29233df, 32'h42ae633c, 32'h41974949, 32'hc2ad69f5, 32'h42670ebd, 32'hc298dfd4};
test_weights[30000:30007] = '{32'hc1e3d1da, 32'hc1fd1f7a, 32'h417419a3, 32'hc1296094, 32'hc1d6210a, 32'h427f7dfc, 32'h42c22f80, 32'hc296e06e};
test_bias[3750:3750] = '{32'hc29c2a4e};
test_output[3750:3750] = '{32'h43355920};
test_input[30008:30015] = '{32'hc2bc5bce, 32'h426da749, 32'h421cc8ea, 32'h42b2d4e4, 32'h419f545d, 32'h428afc32, 32'hc0958b7b, 32'hbfa47eee};
test_weights[30008:30015] = '{32'h42b30dc8, 32'h424ad420, 32'hc230125f, 32'hc227314e, 32'hc23589a2, 32'hbf82adb4, 32'hc2246a14, 32'hc2a686f8};
test_bias[3751:3751] = '{32'h42226b94};
test_output[3751:3751] = '{32'hc633f324};
test_input[30016:30023] = '{32'h42876613, 32'hc2b62b5a, 32'hc2ace5cf, 32'h429262a0, 32'hc24322b7, 32'hc28f56cf, 32'hc2a237f7, 32'hc1fee06d};
test_weights[30016:30023] = '{32'h42b34d3b, 32'h4201e741, 32'h42259731, 32'hbf499ea5, 32'h42b94e8b, 32'h4214c1e1, 32'h418e66e2, 32'hc285d545};
test_bias[3752:3752] = '{32'h42a0e2bc};
test_output[3752:3752] = '{32'hc5d8ef2a};
test_input[30024:30031] = '{32'h4229ed5d, 32'hc0d5beef, 32'hc2272141, 32'hc2a023b2, 32'h42bbb7f0, 32'h425b8dac, 32'h4172a1c7, 32'h429a006b};
test_weights[30024:30031] = '{32'h42a704e0, 32'hc11a2d1c, 32'h409df511, 32'hc24ff488, 32'h42255e33, 32'hc2913041, 32'h429cddac, 32'h42870154};
test_bias[3753:3753] = '{32'h4248bb08};
test_output[3753:3753] = '{32'h46593643};
test_input[30032:30039] = '{32'hc2117d52, 32'h4217a2ab, 32'h42a0a358, 32'h42a7fcba, 32'hc1f15c42, 32'hc2b6f5d6, 32'hc28a3006, 32'hc2a88a4d};
test_weights[30032:30039] = '{32'hc20900bd, 32'hc2ad3a62, 32'h42621b32, 32'h41379983, 32'hc200c578, 32'hc20adac3, 32'hc1306714, 32'hc2822c74};
test_bias[3754:3754] = '{32'h4207b40f};
test_output[3754:3754] = '{32'h4659170e};
test_input[30040:30047] = '{32'h40cb62c9, 32'h42c7b278, 32'h4285cccc, 32'h424547e1, 32'h41938717, 32'h4202938f, 32'h42c3a35a, 32'hc22ac708};
test_weights[30040:30047] = '{32'h40660a6b, 32'h41b2b1b8, 32'h42b3f23a, 32'hc20767d8, 32'h42875202, 32'h42aa22ad, 32'hc286876f, 32'h423ffbc3};
test_bias[3755:3755] = '{32'h429ecb4c};
test_output[3755:3755] = '{32'h4501df3e};
test_input[30048:30055] = '{32'h41f55669, 32'h429837d3, 32'hc21ebd5e, 32'h429d530a, 32'h4242e1e8, 32'hc202710d, 32'hc224ef1f, 32'hc2c63989};
test_weights[30048:30055] = '{32'h41ef0dbf, 32'hc160f1d2, 32'h416cf34d, 32'hc28ead65, 32'hc2305f37, 32'hc2ae18d1, 32'hc2b0db30, 32'h42976b45};
test_bias[3756:3756] = '{32'h42ae26e1};
test_output[3756:3756] = '{32'hc6136414};
test_input[30056:30063] = '{32'h4243f72f, 32'h426a14c1, 32'hc0cc29a0, 32'hc2553385, 32'h42837780, 32'h42824d44, 32'h42c0419d, 32'hc201386f};
test_weights[30056:30063] = '{32'hc207e180, 32'h4284b18b, 32'h427cc9e1, 32'h42009fe7, 32'h420e8d4d, 32'hc275cdde, 32'h3fae8d2e, 32'h4271abd6};
test_bias[3757:3757] = '{32'h402b80ab};
test_output[3757:3757] = '{32'hc5531c65};
test_input[30064:30071] = '{32'h42ac9724, 32'h404f5e1a, 32'hc029b494, 32'hc249c8a8, 32'hc2bc56e5, 32'hc1f3c013, 32'h42083192, 32'h42a7da75};
test_weights[30064:30071] = '{32'h400adc52, 32'hc2c68ed3, 32'hc1d9373a, 32'hc250a332, 32'h4223fd2d, 32'h400f5e92, 32'hc2032910, 32'hc19ea73b};
test_bias[3758:3758] = '{32'h413dceec};
test_output[3758:3758] = '{32'hc5810948};
test_input[30072:30079] = '{32'h427af057, 32'h42597ba8, 32'hc2a077e2, 32'hc28401fb, 32'hc25489cf, 32'h42958e25, 32'hc28168a0, 32'hc111055b};
test_weights[30072:30079] = '{32'hc286c75d, 32'h428a6471, 32'hc19fea1e, 32'hc27e6a87, 32'hc24614b5, 32'hc298259a, 32'hc1f7b5c7, 32'h42559539};
test_bias[3759:3759] = '{32'h4269f0de};
test_output[3759:3759] = '{32'h457112f0};
test_input[30080:30087] = '{32'hc2789327, 32'hc2bedd68, 32'h4265082d, 32'h41877c6f, 32'h42961033, 32'hc1ac8b9a, 32'h422822e4, 32'h42c03d37};
test_weights[30080:30087] = '{32'h423b9888, 32'hc27a952e, 32'hc1f23526, 32'h42bbb08a, 32'h42317879, 32'hc1a0d198, 32'hc28ba1e4, 32'hc290787c};
test_bias[3760:3760] = '{32'h42423652};
test_output[3760:3760] = '{32'hc544b097};
test_input[30088:30095] = '{32'h40ba7e72, 32'hc10b4722, 32'hc297034b, 32'h414f3919, 32'hc204a291, 32'hc20ba1ed, 32'h42baed78, 32'hbf32cb19};
test_weights[30088:30095] = '{32'h42750f92, 32'h418c1458, 32'hc192af80, 32'h4199476d, 32'h428185d1, 32'h42912fcf, 32'h423d019b, 32'hc280ffd7};
test_bias[3761:3761] = '{32'hc265e90d};
test_output[3761:3761] = '{32'h44c2f3a9};
test_input[30096:30103] = '{32'h41806759, 32'h415cd2b2, 32'hc1ae2756, 32'hc2808b75, 32'hc2181dd2, 32'hc25ab1a5, 32'h42b6a0c0, 32'h42ba966e};
test_weights[30096:30103] = '{32'hc2601acc, 32'h425fbe75, 32'hc1b0bd82, 32'hc27a60eb, 32'hc1c1c9ee, 32'h426c68bd, 32'hc28f665e, 32'h42796851};
test_bias[3762:3762] = '{32'h429e78bd};
test_output[3762:3762] = '{32'h44b0f7c8};
test_input[30104:30111] = '{32'hc190ae41, 32'h413c77cb, 32'h42445d60, 32'hc288dc49, 32'h42435fc4, 32'hc1c396ae, 32'hc20a464d, 32'h42b5bc8a};
test_weights[30104:30111] = '{32'hc1cc5420, 32'h4210b1a1, 32'hc2afa845, 32'h423f6d95, 32'hc2953b4d, 32'hc2174a41, 32'h418eef88, 32'hc2b5ad54};
test_bias[3763:3763] = '{32'hc1a3b2a3};
test_output[3763:3763] = '{32'hc68f0d66};
test_input[30112:30119] = '{32'h41f82b38, 32'hc1d3570f, 32'hc1e730ca, 32'h42bb2f3c, 32'hc269071e, 32'hc17aaf5f, 32'h4173930e, 32'h42aa757d};
test_weights[30112:30119] = '{32'hc2584822, 32'h42a87bbd, 32'h416c30da, 32'hc20cd9b5, 32'h42ae1f99, 32'hc297fe85, 32'h420f6aae, 32'hc06eaea8};
test_bias[3764:3764] = '{32'h42a3998f};
test_output[3764:3764] = '{32'hc62ef1f0};
test_input[30120:30127] = '{32'h4193da4d, 32'h412dc543, 32'h4222c7c1, 32'hc2737983, 32'h420b532a, 32'h42462402, 32'h425d6e5d, 32'h4100ca4a};
test_weights[30120:30127] = '{32'h41ef587a, 32'hc2724c7d, 32'hc257623f, 32'h4286b85a, 32'h4214243b, 32'hc288b533, 32'h4291e179, 32'h4291f70c};
test_bias[3765:3765] = '{32'h42af0f02};
test_output[3765:3765] = '{32'hc56c3736};
test_input[30128:30135] = '{32'hc227f4e5, 32'h42a1e95d, 32'hc1f76116, 32'h420208ea, 32'hc2afd6e4, 32'hc066c612, 32'h420e95f8, 32'h42b25cc2};
test_weights[30128:30135] = '{32'hc26680ec, 32'h40a0ae8f, 32'hc21f309b, 32'hc21508f8, 32'h414af379, 32'h3ff6096f, 32'h429759e2, 32'hc299dfd9};
test_bias[3766:3766] = '{32'hc15dd8cb};
test_output[3766:3766] = '{32'hc51963a3};
test_input[30136:30143] = '{32'h41c1be1d, 32'hc2995ba8, 32'h42a85e10, 32'hc0a9c9d6, 32'hc216a53e, 32'h41d2528f, 32'hc231c11a, 32'hc26cf981};
test_weights[30136:30143] = '{32'h429e9c8b, 32'hc21a4528, 32'h422be2e9, 32'h407ea611, 32'hc29251c4, 32'hc27025aa, 32'hc22752f1, 32'hc24ba8c1};
test_bias[3767:3767] = '{32'h41bda78e};
test_output[3767:3767] = '{32'h466358f1};
test_input[30144:30151] = '{32'hc0e7ac0d, 32'h429e6133, 32'hc2858270, 32'hc20e0951, 32'hc2409636, 32'hc28fe1cc, 32'h41ee6d9e, 32'h42a5d425};
test_weights[30144:30151] = '{32'hc2a3f842, 32'hc2c35a54, 32'hc2264bbc, 32'hc27772a9, 32'hc0e8f44c, 32'hc2518605, 32'h41d4fc37, 32'hc2afef77};
test_bias[3768:3768] = '{32'h4295b1a6};
test_output[3768:3768] = '{32'hc58be130};
test_input[30152:30159] = '{32'hc05e44fe, 32'h3f1b9181, 32'h429709f0, 32'hc29cfcc5, 32'hc287586f, 32'hc2b10996, 32'h4297728e, 32'hc274d9fe};
test_weights[30152:30159] = '{32'hc19a451d, 32'hc1a5153e, 32'hc2c427d8, 32'hc2953251, 32'h42a6c0e4, 32'h42af5c33, 32'hc23d4f9b, 32'h4204b61a};
test_bias[3769:3769] = '{32'h42a59512};
test_output[3769:3769] = '{32'hc69fa0ee};
test_input[30160:30167] = '{32'hc2acc511, 32'h4280b763, 32'hc2c0d140, 32'hc2423408, 32'hc2a25315, 32'h411007d1, 32'h421ffff6, 32'h417059be};
test_weights[30160:30167] = '{32'h3f3f13b1, 32'hc2bda256, 32'h429c51bd, 32'h423a50b3, 32'hc2a0424d, 32'h41f1e6c9, 32'hc2790479, 32'hc17b61d8};
test_bias[3770:3770] = '{32'hc28ec98b};
test_output[3770:3770] = '{32'hc63b4554};
test_input[30168:30175] = '{32'hc1743544, 32'h421f1868, 32'hc2200e06, 32'h42bb0a6a, 32'hc265722e, 32'hc1fe89dd, 32'h4221bca4, 32'h41bc22b2};
test_weights[30168:30175] = '{32'h40103bf3, 32'h42b31d73, 32'hc2709f22, 32'h3fb539e4, 32'h414611d2, 32'h404be342, 32'h41ce7222, 32'h420d1662};
test_bias[3771:3771] = '{32'hc2ade58b};
test_output[3771:3771] = '{32'h45dc0ce0};
test_input[30176:30183] = '{32'h42235af9, 32'h4105374d, 32'hc288e83a, 32'h41d359f0, 32'hc29c4fc8, 32'h42b5cec5, 32'h40b8a676, 32'hc1068149};
test_weights[30176:30183] = '{32'h4130a912, 32'hc19414a7, 32'h417615ae, 32'h4201a29e, 32'h42b72e1a, 32'h42526df3, 32'h42718bd9, 32'h41e8f820};
test_bias[3772:3772] = '{32'h3e512ebb};
test_output[3772:3772] = '{32'hc507c11d};
test_input[30184:30191] = '{32'hc244b0e8, 32'h41dc209d, 32'h4204a0e7, 32'h42acc4d2, 32'hc26ebcf9, 32'hc2737c4b, 32'h427cdd64, 32'hc200d3cf};
test_weights[30184:30191] = '{32'h42c7fe21, 32'hc283e1ac, 32'h42be7fcc, 32'hc286b9a2, 32'hc2a2ee38, 32'h428b8ab1, 32'hc22ce633, 32'hc16f187d};
test_bias[3773:3773] = '{32'h4224aeb1};
test_output[3773:3773] = '{32'hc62bad1b};
test_input[30192:30199] = '{32'h429a435c, 32'hc274db4c, 32'hc201e09a, 32'hc279057d, 32'hc2a9d030, 32'h415badf8, 32'h42099abe, 32'hc2619edf};
test_weights[30192:30199] = '{32'hc2b7befe, 32'h41b32913, 32'hc248ca07, 32'h424f2af3, 32'h41f50a0e, 32'h42657071, 32'h428672de, 32'hc2be5b46};
test_bias[3774:3774] = '{32'hc1142bed};
test_output[3774:3774] = '{32'hc5830752};
test_input[30200:30207] = '{32'h426e4f70, 32'h4203d38c, 32'hc2c7016c, 32'hc027815e, 32'h4283b000, 32'hc2a0cd50, 32'h4104f7f8, 32'hc0b72186};
test_weights[30200:30207] = '{32'h42bf2198, 32'h428010a2, 32'h42c7d647, 32'hc1cd9dcd, 32'hc2b57de0, 32'hc2ab2295, 32'hc0ac4c5f, 32'h42961f10};
test_bias[3775:3775] = '{32'hc1e73181};
test_output[3775:3775] = '{32'hc4d0b27a};
test_input[30208:30215] = '{32'hc2899993, 32'h42309dc4, 32'h42b2a23f, 32'hc22b0a71, 32'hc2923c50, 32'hc20c6b6f, 32'h42924c49, 32'hc2a93092};
test_weights[30208:30215] = '{32'hc0cbf8c1, 32'hc170154c, 32'h4287eb8e, 32'h41ff8f52, 32'h417010f7, 32'h42b9e23b, 32'hc2b0108d, 32'h42b10279};
test_bias[3776:3776] = '{32'hc282c84c};
test_output[3776:3776] = '{32'hc658bece};
test_input[30216:30223] = '{32'hc09aa218, 32'h429c22b3, 32'h42580d79, 32'hc2a88d7f, 32'hc1bd6bda, 32'h42afbbbb, 32'hc0c256b6, 32'h42c570db};
test_weights[30216:30223] = '{32'h42c2dec0, 32'h42447494, 32'hbfba0457, 32'hc2b5deb4, 32'hc2a47b53, 32'h40c4c71f, 32'hc1d5f559, 32'hc2c39071};
test_bias[3777:3777] = '{32'h42b53d79};
test_output[3777:3777] = '{32'h457c4171};
test_input[30224:30231] = '{32'h41de5c3a, 32'h428ac95f, 32'hc1aa76f7, 32'h3fa99bce, 32'hc2359cbd, 32'h42b084d0, 32'h41466eee, 32'hc2bf3c38};
test_weights[30224:30231] = '{32'hc20f9faf, 32'hc2c17ba0, 32'hc2bdabbd, 32'h4290a55a, 32'h422ba755, 32'h4265c810, 32'h41625941, 32'hbeff07e8};
test_bias[3778:3778] = '{32'h41ed2082};
test_output[3778:3778] = '{32'hc50ac35a};
test_input[30232:30239] = '{32'hc291f6c2, 32'hc29bc9de, 32'h4241561c, 32'h429edb6e, 32'hc1db8bbf, 32'hc271d7ac, 32'h418f48b2, 32'h42504fac};
test_weights[30232:30239] = '{32'hc28cbc1e, 32'hc17e80ce, 32'h425d9fbc, 32'hc284bc77, 32'h424a3850, 32'h42158d43, 32'hc046798f, 32'hc282b14d};
test_bias[3779:3779] = '{32'h42593867};
test_output[3779:3779] = '{32'hc54c72c7};
test_input[30240:30247] = '{32'hc00d7320, 32'hc2b0eff5, 32'h42aa9071, 32'h42a409b7, 32'hc24bff53, 32'hc24ae244, 32'h40d9a2f2, 32'h4083f414};
test_weights[30240:30247] = '{32'hc1d3f645, 32'hc27045f4, 32'h428bbb17, 32'h4284cf66, 32'h42182827, 32'h42366f3f, 32'h42661a86, 32'h42143aad};
test_bias[3780:3780] = '{32'h4198e47c};
test_output[3780:3780] = '{32'h464c7d5d};
test_input[30248:30255] = '{32'hc2421e7e, 32'h422709df, 32'hc2629e60, 32'h42a377e4, 32'hc2bf9837, 32'hc1fda769, 32'hc2278ca1, 32'hc2b46b98};
test_weights[30248:30255] = '{32'h42ba5a7b, 32'h426b5d7c, 32'hc203b729, 32'hc29638d7, 32'hc280b251, 32'h41b9d79d, 32'h428de8cd, 32'hc2ac35ee};
test_bias[3781:3781] = '{32'hc25b40fb};
test_output[3781:3781] = '{32'h456f6469};
test_input[30256:30263] = '{32'h429d8396, 32'h4218ffb9, 32'hc2a90021, 32'h42861825, 32'hc2abf1f8, 32'h418a8596, 32'h42b5c98f, 32'hc20511ae};
test_weights[30256:30263] = '{32'h424a5212, 32'hc2b98546, 32'h4257eb23, 32'h425550eb, 32'hc1ea55ef, 32'hc1734eb6, 32'h4128f6ca, 32'hc214fa43};
test_bias[3782:3782] = '{32'h41e735b4};
test_output[3782:3782] = '{32'h4575c87e};
test_input[30264:30271] = '{32'hc2150750, 32'hc2c64c5c, 32'hc1c909b6, 32'h4157898c, 32'h425e726d, 32'h423d6005, 32'h42a84436, 32'hc2a7d5eb};
test_weights[30264:30271] = '{32'hc1d8a186, 32'h41e788a4, 32'h426409b4, 32'h4114bb10, 32'hc2949995, 32'h411d39a6, 32'hc2711160, 32'hc22f4960};
test_bias[3783:3783] = '{32'h429198ff};
test_output[3783:3783] = '{32'hc5fed84d};
test_input[30272:30279] = '{32'h4081760a, 32'h4190824d, 32'hc28ae85a, 32'h42bb9430, 32'h42adf69c, 32'hc2bef1cd, 32'h42a53e26, 32'h420fbe37};
test_weights[30272:30279] = '{32'h42a07019, 32'h413b3df5, 32'hc1655776, 32'h428dd085, 32'hc1fb6b82, 32'h427475bb, 32'hc1cd00f3, 32'hc152c4d1};
test_bias[3784:3784] = '{32'h4118fd3b};
test_output[3784:3784] = '{32'hc53979c4};
test_input[30280:30287] = '{32'hc28e8890, 32'hc17f2f45, 32'h42b0c6b8, 32'h42bba8ab, 32'hc2c3856a, 32'h421cee83, 32'h4270aab5, 32'h42bc13c9};
test_weights[30280:30287] = '{32'hc246c057, 32'hc2b7329d, 32'hc2ae398d, 32'hc23b515e, 32'hc232b28c, 32'h4172cfdd, 32'hc2419412, 32'h42373456};
test_bias[3785:3785] = '{32'hc2895789};
test_output[3785:3785] = '{32'hc4488f72};
test_input[30288:30295] = '{32'hc22be0db, 32'h42158cc9, 32'h41546f4a, 32'hbf2cc9f6, 32'hc29c7b47, 32'hc26937f2, 32'h4273ac9c, 32'hc2b75ecd};
test_weights[30288:30295] = '{32'hc23cfcc4, 32'hc240d0a8, 32'hc0a9e726, 32'h420f017d, 32'hc29fb9d5, 32'h42a7da6e, 32'h428c80b3, 32'h41844294};
test_bias[3786:3786] = '{32'h42b59cb6};
test_output[3786:3786] = '{32'h4587b991};
test_input[30296:30303] = '{32'h428d0e46, 32'h426a21a4, 32'hc2170736, 32'h42489e38, 32'h42bb2f7e, 32'h42943192, 32'h42a2b8d6, 32'h42a49b12};
test_weights[30296:30303] = '{32'hc270ee2c, 32'h424e9f99, 32'hc250cfca, 32'hc21f95ea, 32'hbe8eda48, 32'hbf2a6da8, 32'hc17f2830, 32'hc2c4f0ac};
test_bias[3787:3787] = '{32'hc24c6e0a};
test_output[3787:3787] = '{32'hc6287b81};
test_input[30304:30311] = '{32'h4274412b, 32'h41abd5f2, 32'h422ade00, 32'h42745d99, 32'hc17da712, 32'h42c1b3bc, 32'hc12dd8bf, 32'hc202ad03};
test_weights[30304:30311] = '{32'h42990405, 32'h425c35fb, 32'hbdb98ad2, 32'h4207e1af, 32'h42655ccf, 32'h4226b6f6, 32'hc2b7e047, 32'hc2737bf2};
test_bias[3788:3788] = '{32'hc227f81d};
test_output[3788:3788] = '{32'h465abba5};
test_input[30312:30319] = '{32'h3ff2e3dc, 32'h423b5841, 32'hc2867612, 32'hc208e5c1, 32'h42af7aea, 32'hc29a8334, 32'h427ab98d, 32'h424876b9};
test_weights[30312:30319] = '{32'hc09b0552, 32'h418f0960, 32'h429917d5, 32'hc2223726, 32'h42aad2d8, 32'hc2036874, 32'hc2947fc0, 32'h42b0c5a3};
test_bias[3789:3789] = '{32'h4203ce39};
test_output[3789:3789] = '{32'h45d7f31e};
test_input[30320:30327] = '{32'hc20160ba, 32'h427c7a47, 32'h4205f28f, 32'hc1ef9304, 32'h42476a5d, 32'hc286d892, 32'h4283cd79, 32'hc2682669};
test_weights[30320:30327] = '{32'hc2557a73, 32'hc11f521c, 32'h42449698, 32'h42457372, 32'h3ee6c779, 32'h41913274, 32'h40888c73, 32'h4299ed09};
test_bias[3790:3790] = '{32'h4280b3b4};
test_output[3790:3790] = '{32'hc57d92fc};
test_input[30328:30335] = '{32'hc23f726f, 32'hc1bf78a0, 32'hc0c0fe2f, 32'h4204185c, 32'h42c51be8, 32'h42a2b778, 32'h42944308, 32'hc29ab538};
test_weights[30328:30335] = '{32'hc2427f68, 32'hc2b0ce00, 32'hc2526752, 32'hc29875ef, 32'h42c5e9f2, 32'h41c39218, 32'h425f6260, 32'h3f7f7fbc};
test_bias[3791:3791] = '{32'hc29c1c31};
test_output[3791:3791] = '{32'h468c623a};
test_input[30336:30343] = '{32'h42062bb1, 32'h415c84f9, 32'h422ee1cb, 32'h428edbfb, 32'hc27cf1d8, 32'h41f46183, 32'h4202a583, 32'h4293ca86};
test_weights[30336:30343] = '{32'hc1fb1a80, 32'h424b6254, 32'hc1f6b82e, 32'hc2bd2bee, 32'h4224d338, 32'h42a34672, 32'hc2387a88, 32'hc265246c};
test_bias[3792:3792] = '{32'h42b22437};
test_output[3792:3792] = '{32'hc65e2bbd};
test_input[30344:30351] = '{32'h408e5ea9, 32'h4280d76b, 32'h426b402d, 32'hc2c5fd16, 32'h42605525, 32'h4222027d, 32'h4097a44e, 32'hc1b34431};
test_weights[30344:30351] = '{32'hc27ca4b2, 32'h42ab26b3, 32'hc1cbaa5a, 32'h41b718ec, 32'hc23db795, 32'hc1f7546c, 32'h42a31cd1, 32'hc28712fa};
test_bias[3793:3793] = '{32'hc1b0038c};
test_output[3793:3793] = '{32'hc40d5b23};
test_input[30352:30359] = '{32'h429fa2f0, 32'h42394d3e, 32'h42330969, 32'hc03a2a00, 32'hc26cdec5, 32'hbfbb55e6, 32'h42ab4aea, 32'h421314d5};
test_weights[30352:30359] = '{32'h42127c96, 32'hc2985a75, 32'h4196b592, 32'hc1964af4, 32'h429b39fa, 32'h42872ccb, 32'h42a5d995, 32'hc1a48a42};
test_bias[3794:3794] = '{32'hbe2a62a0};
test_output[3794:3794] = '{32'h44f2d9b0};
test_input[30360:30367] = '{32'hc15d5d45, 32'h42b0c251, 32'h41666e4d, 32'hc1a87340, 32'h40626d6d, 32'hc2700891, 32'h424ab581, 32'h4162570f};
test_weights[30360:30367] = '{32'h41326932, 32'h40f8fcc4, 32'h42751ca7, 32'hc1771e25, 32'h42c68663, 32'hc18f35f3, 32'hc29b79df, 32'h424386fe};
test_bias[3795:3795] = '{32'h428a192d};
test_output[3795:3795] = '{32'hc1476ce0};
test_input[30368:30375] = '{32'h40d2270d, 32'hc29a88bb, 32'hc20b0901, 32'h42a61578, 32'h424cc314, 32'h41804acd, 32'hbed01e2a, 32'hc2b8b636};
test_weights[30368:30375] = '{32'h4268470e, 32'hc186ca93, 32'h428fa712, 32'hc227e438, 32'h42a19b16, 32'h4272feed, 32'h42639deb, 32'h41c3a480};
test_bias[3796:3796] = '{32'hc12ab2bd};
test_output[3796:3796] = '{32'hc4b91755};
test_input[30376:30383] = '{32'hc1b50de3, 32'h429f5535, 32'h41eb0f10, 32'hc2075be5, 32'h423fb865, 32'hc261bc0b, 32'hc288afcb, 32'h42c572db};
test_weights[30376:30383] = '{32'h42c3a73b, 32'h42a08f23, 32'h4248348c, 32'hc2b61459, 32'h3fe49d43, 32'hc243992b, 32'h42992a90, 32'hc2a9422f};
test_bias[3797:3797] = '{32'h41d50f3e};
test_output[3797:3797] = '{32'hc4f803a8};
test_input[30384:30391] = '{32'h421267a3, 32'hc1e4b5fb, 32'hc18fd3b6, 32'h41a230c5, 32'hc23c3b6d, 32'h422e0075, 32'hc2ba92c0, 32'h42ab7bff};
test_weights[30384:30391] = '{32'h41fd335e, 32'hc235d20a, 32'h428c038e, 32'h4281d674, 32'h418856ee, 32'hc28de164, 32'hc2a959dc, 32'h42430fba};
test_bias[3798:3798] = '{32'hc243f5f6};
test_output[3798:3798] = '{32'h46268bac};
test_input[30392:30399] = '{32'h41a6823f, 32'hc0b266ac, 32'hc2b6c20c, 32'hc22a0bf3, 32'h421fde8c, 32'h40c8a654, 32'hbf6047b9, 32'h41f4e31c};
test_weights[30392:30399] = '{32'h423aed01, 32'h4177b67b, 32'h42ac203b, 32'hc2746c51, 32'hc22cab9f, 32'h42665d0c, 32'h429f1791, 32'h41ba0875};
test_bias[3799:3799] = '{32'hc27a9cd8};
test_output[3799:3799] = '{32'hc5a167f8};
test_input[30400:30407] = '{32'h412c58b3, 32'hc26e966e, 32'hc168710d, 32'hc2a1b916, 32'h425cbe4f, 32'h41d6eb95, 32'h42bbcb59, 32'h429b0fc1};
test_weights[30400:30407] = '{32'h40f4a97f, 32'hc2beae56, 32'hc261f8bb, 32'hc2bf74c8, 32'h41bd46be, 32'hc2940694, 32'hc1cd14ba, 32'hbfa5bc27};
test_bias[3800:3800] = '{32'h41a59f4e};
test_output[3800:3800] = '{32'h462e6471};
test_input[30408:30415] = '{32'h422aaa0b, 32'hc2376b86, 32'h426280ca, 32'hc25fd0f1, 32'hc21bd581, 32'h42bdc6d3, 32'h4239837c, 32'h42727c74};
test_weights[30408:30415] = '{32'hc26303b2, 32'hc275543f, 32'h42906c5e, 32'hc2a3c66f, 32'hc163725a, 32'h40c16937, 32'h41bf9fbe, 32'hc2a9d7f2};
test_bias[3801:3801] = '{32'hc19fd459};
test_output[3801:3801] = '{32'h45bfa0a4};
test_input[30416:30423] = '{32'h41c26308, 32'hc2124941, 32'h42187ba9, 32'hc109e6f2, 32'hc286dbd9, 32'h4164cd83, 32'h41bbc00b, 32'hc2bcbebc};
test_weights[30416:30423] = '{32'hc1e8226b, 32'hc1c51a08, 32'hc2695066, 32'h42a91df6, 32'hc20530e0, 32'hc202ba2e, 32'hc29b2bd0, 32'h42bcce1e};
test_bias[3802:3802] = '{32'hc29c8723};
test_output[3802:3802] = '{32'hc6382a48};
test_input[30424:30431] = '{32'hc1b0db30, 32'h42c74a21, 32'hc1288703, 32'hc2a3b3d6, 32'h40dd1298, 32'h42c71a60, 32'hc26cc13c, 32'h426c3f2b};
test_weights[30424:30431] = '{32'hc28a8fca, 32'h428c3d6e, 32'h4232aea6, 32'h42ae216f, 32'h42079525, 32'hc2948e00, 32'hc2c14a5b, 32'hc27b5507};
test_bias[3803:3803] = '{32'h42523b82};
test_output[3803:3803] = '{32'hc582852f};
test_input[30432:30439] = '{32'hc283c767, 32'h42384c37, 32'h41bdc7d7, 32'h420b3be9, 32'h40415dae, 32'h428f74eb, 32'h421ba4af, 32'h423393ba};
test_weights[30432:30439] = '{32'hc1cd15fb, 32'h42a3a039, 32'h4221efcf, 32'h42abd89f, 32'h3fd53416, 32'hc209aa12, 32'h3ecbdad8, 32'h4285ad5b};
test_bias[3804:3804] = '{32'h41269419};
test_output[3804:3804] = '{32'h461bd365};
test_input[30440:30447] = '{32'hc2c44102, 32'hc1b4292b, 32'h423d783e, 32'h4201ba8e, 32'hc288f060, 32'hc2aacbee, 32'h4285db75, 32'h4206191d};
test_weights[30440:30447] = '{32'hc25cd87d, 32'h42915573, 32'hc25d7238, 32'hc299e83d, 32'h4025af8f, 32'hc24bc998, 32'h413a6bd0, 32'h40a947f1};
test_bias[3805:3805] = '{32'hc297f06b};
test_output[3805:3805] = '{32'h45685dbf};
test_input[30448:30455] = '{32'hc0827746, 32'hc0cad619, 32'hc2c2bf40, 32'hc230dace, 32'hc2c0f52a, 32'hc2a734c2, 32'h42aae063, 32'hc137c882};
test_weights[30448:30455] = '{32'h42c09491, 32'hc2999de8, 32'hc20df110, 32'hc27d8361, 32'h41c43a5c, 32'h429a7ad6, 32'h40ae991c, 32'h42655a3e};
test_bias[3806:3806] = '{32'h4250f533};
test_output[3806:3806] = '{32'hc52345eb};
test_input[30456:30463] = '{32'h42c1d93a, 32'h428ad5b9, 32'h422c7ed1, 32'h4238d6e3, 32'h42499365, 32'h429d496e, 32'h41b67889, 32'h42ab697a};
test_weights[30456:30463] = '{32'h4264b917, 32'h422c45b6, 32'hc1a7f4fd, 32'h42038261, 32'hc251d617, 32'hc2052d87, 32'hc2a434db, 32'hc127c206};
test_bias[3807:3807] = '{32'h423e2d80};
test_output[3807:3807] = '{32'h44910018};
test_input[30464:30471] = '{32'hc1ecf677, 32'h42c36474, 32'h42ac3aaf, 32'h42c0df95, 32'hc2b0131f, 32'h42aa52bc, 32'hc08f2a07, 32'hc2b0f556};
test_weights[30464:30471] = '{32'h41f156c4, 32'h421dbe0b, 32'h426587ce, 32'h3fc8e9e7, 32'h4260dc8f, 32'h42a819dc, 32'hc230d236, 32'hc22d8239};
test_bias[3808:3808] = '{32'hc2346de0};
test_output[3808:3808] = '{32'h465eadce};
test_input[30472:30479] = '{32'hc28570b6, 32'h426a52ba, 32'h428b9b4a, 32'h40bb433f, 32'h42b4e1cc, 32'hc27f8533, 32'hc2aa7a12, 32'h4268a23a};
test_weights[30472:30479] = '{32'h427405e5, 32'hc24013a0, 32'h42a25483, 32'h425112ac, 32'hc1293f4d, 32'h4281f588, 32'hc29f2678, 32'h42844933};
test_bias[3809:3809] = '{32'hc1ce2cac};
test_output[3809:3809] = '{32'h458f4367};
test_input[30480:30487] = '{32'hc23df77f, 32'hc263eeac, 32'h41048c58, 32'h42103678, 32'hc2487d1d, 32'h41f23681, 32'h415ae11e, 32'hc2617a76};
test_weights[30480:30487] = '{32'hc27b2acc, 32'h41cc5f25, 32'hc1ca4ecd, 32'hc1069a72, 32'h4277289a, 32'h42697e33, 32'h40602337, 32'h425d8399};
test_bias[3810:3810] = '{32'hc2afea82};
test_output[3810:3810] = '{32'hc5595d45};
test_input[30488:30495] = '{32'hc264a9c4, 32'h4059cc1d, 32'hc1256476, 32'h42b1bf98, 32'hc15aa0e8, 32'hc24840b9, 32'hc23be695, 32'h425598cb};
test_weights[30488:30495] = '{32'h41dbabbc, 32'hc16457ae, 32'h42acde2e, 32'h40f8b7f3, 32'h40081f5a, 32'h42b48ae4, 32'h41b8c8ec, 32'hc1f8629e};
test_bias[3811:3811] = '{32'h420ae2d8};
test_output[3811:3811] = '{32'hc60dd646};
test_input[30496:30503] = '{32'hc28f94cc, 32'hc1ccb813, 32'h41aa2147, 32'hc2a23dfa, 32'hc2477318, 32'hc24c5e8e, 32'h42a7161d, 32'h41c83429};
test_weights[30496:30503] = '{32'hc1ba5fd5, 32'h42ab8382, 32'h42b618c7, 32'hc0ed0be9, 32'hc0bfa348, 32'h3e887b37, 32'hc22c6c4f, 32'hc241a4e5};
test_bias[3812:3812] = '{32'h41be0dfd};
test_output[3812:3812] = '{32'hc51b8caf};
test_input[30504:30511] = '{32'h40b2491d, 32'hc0a32a31, 32'hc192c50f, 32'hc258182f, 32'hc1273b57, 32'hc024fdf9, 32'hc2bf3be5, 32'hc2af8f01};
test_weights[30504:30511] = '{32'h40c7faa1, 32'hc0a77f84, 32'h41a2a4f0, 32'h42b9a648, 32'h4125bae9, 32'hc1abfb1e, 32'hc218ff37, 32'h4209c961};
test_bias[3813:3813] = '{32'hc2bbcbd8};
test_output[3813:3813] = '{32'hc5973b09};
test_input[30512:30519] = '{32'hc2bfb965, 32'h4118ecf6, 32'h425002ba, 32'h3e017314, 32'hc22472e4, 32'hc2be5b98, 32'hc1b5599a, 32'h420ef045};
test_weights[30512:30519] = '{32'h42ae5f74, 32'hc1cb8d27, 32'h42c79977, 32'h4294ec6c, 32'h4243f79c, 32'hc2506ad9, 32'h42b23965, 32'h424dc019};
test_bias[3814:3814] = '{32'hc0c5beba};
test_output[3814:3814] = '{32'hc421371c};
test_input[30520:30527] = '{32'h428a0aaf, 32'h41f3b568, 32'h42b66a79, 32'hc293efec, 32'h41aab51c, 32'h42879ac3, 32'hc1cbe33b, 32'hc28142e2};
test_weights[30520:30527] = '{32'h42c3dd92, 32'h42adf2a8, 32'h4288701a, 32'h42beaaec, 32'h428bb4f2, 32'hc29ca95a, 32'h41c53bdf, 32'hc1311d80};
test_bias[3815:3815] = '{32'hc2391a20};
test_output[3815:3815] = '{32'h4595fdd8};
test_input[30528:30535] = '{32'hc263a409, 32'h3ed6c261, 32'h423d34b0, 32'hc2c48ce2, 32'h41f5839a, 32'h429d326d, 32'hc27be5e0, 32'h41c186dd};
test_weights[30528:30535] = '{32'hc25352af, 32'h419e7d71, 32'hc209c54a, 32'hc27c7bd8, 32'h3fe924e4, 32'hc1e86cae, 32'hc2721718, 32'hc0a0d167};
test_bias[3816:3816] = '{32'hc20edb2b};
test_output[3816:3816] = '{32'h460cdda6};
test_input[30536:30543] = '{32'h4244b745, 32'h412be891, 32'h4032103c, 32'h3f580d19, 32'hc28e2495, 32'hc2b80af8, 32'hc245ec25, 32'hc20f0c29};
test_weights[30536:30543] = '{32'hc292cae5, 32'h41c3c982, 32'h426d353f, 32'hc18f8b7f, 32'h4125fccd, 32'h4233c019, 32'hc2c3155d, 32'hc2c3ace8};
test_bias[3817:3817] = '{32'hc2853036};
test_output[3817:3817] = '{32'h433d66e2};
test_input[30544:30551] = '{32'h428c2e75, 32'h41df9379, 32'h419a6dcb, 32'hc2ab1787, 32'h41ce6431, 32'h420a9da6, 32'hc2b016e4, 32'hc1899ceb};
test_weights[30544:30551] = '{32'hc28a8940, 32'h420f65c7, 32'h422833cd, 32'h40bc3bb4, 32'hc2a64d93, 32'hc23b9c1b, 32'h42aa70a7, 32'hc1cba107};
test_bias[3818:3818] = '{32'hc2913165};
test_output[3818:3818] = '{32'hc661d494};
test_input[30552:30559] = '{32'h41df19e6, 32'h428a1e1a, 32'h41f82e6b, 32'h408325f4, 32'h4156535d, 32'hc2ae3a1e, 32'h425a55dc, 32'hc26dad99};
test_weights[30552:30559] = '{32'hc04ce7a2, 32'h4290ace0, 32'hc25f633d, 32'h42c48222, 32'hc2b099f6, 32'hc238b50b, 32'hc2a1b7c9, 32'h42b01d6c};
test_bias[3819:3819] = '{32'hc298f53c};
test_output[3819:3819] = '{32'hc54ea2c6};
test_input[30560:30567] = '{32'hc29da5cc, 32'h4264985d, 32'hc2997b2e, 32'h41d174c3, 32'hc24cae5c, 32'h4296c556, 32'h429a0d0b, 32'hc1a5716d};
test_weights[30560:30567] = '{32'hc2a06159, 32'h427c2dbc, 32'hc269e607, 32'hc298c712, 32'h426d77b9, 32'hc1a0728e, 32'h4257ee82, 32'hc26ec482};
test_bias[3820:3820] = '{32'hc1d41b95};
test_output[3820:3820] = '{32'h464eadbe};
test_input[30568:30575] = '{32'hc2881fee, 32'h429420c3, 32'hc2022d78, 32'h42b89632, 32'h425f9609, 32'h428bf7a3, 32'hc11b7c95, 32'hc23949ee};
test_weights[30568:30575] = '{32'h42314f90, 32'h4250f37f, 32'hc0b16770, 32'hc2860d0e, 32'h426e889b, 32'hc1d6987b, 32'h4279ef4e, 32'hc28ab875};
test_bias[3821:3821] = '{32'hc19e2959};
test_output[3821:3821] = '{32'hc48af75c};
test_input[30576:30583] = '{32'hc284daf6, 32'hc219acae, 32'hc24788ef, 32'hc228c413, 32'hc1bdca26, 32'h4286aa72, 32'h42a9a2b1, 32'hc1d7edb3};
test_weights[30576:30583] = '{32'h421ca573, 32'hc1d098a6, 32'hc18c8ee5, 32'h42880526, 32'hc09ac866, 32'hc1ded210, 32'h428360bc, 32'h42a74a29};
test_bias[3822:3822] = '{32'hc20ba47a};
test_output[3822:3822] = '{32'hc501a4ab};
test_input[30584:30591] = '{32'h4055f0cd, 32'h416362bb, 32'hc1ef11ae, 32'h42086c50, 32'hc2123018, 32'h4282263a, 32'h413131ae, 32'h428c0ee3};
test_weights[30584:30591] = '{32'h42640f7b, 32'hc1541bb4, 32'h41201684, 32'hc2a788ec, 32'hc2a88ad6, 32'h4255875c, 32'hc1f08655, 32'hc1a56e5c};
test_bias[3823:3823] = '{32'hc2c7e5e6};
test_output[3823:3823] = '{32'h44bddc47};
test_input[30592:30599] = '{32'hc2b5d8b8, 32'h42a7c9bf, 32'hc2918c97, 32'h429f5a04, 32'hc2bf6ee6, 32'hc2adb70c, 32'hc1e84f2b, 32'hc2633404};
test_weights[30592:30599] = '{32'hc2c06251, 32'hc28c9c97, 32'hc2432ded, 32'hc28e95de, 32'h42411aa5, 32'h4287f134, 32'h41112960, 32'h42b07bab};
test_bias[3824:3824] = '{32'hc2308f2c};
test_output[3824:3824] = '{32'hc66c5751};
test_input[30600:30607] = '{32'hc19ae76a, 32'hc2c51ee3, 32'h42bdde50, 32'h41b8f128, 32'h41f28631, 32'hc27eac45, 32'hc187ba0c, 32'h42b28095};
test_weights[30600:30607] = '{32'hc277136a, 32'hc24deb33, 32'hc1c56b17, 32'h4285060e, 32'hc128a369, 32'hc2c2bc48, 32'h428a12b5, 32'h40d9b76e};
test_bias[3825:3825] = '{32'h421f1b5e};
test_output[3825:3825] = '{32'h462910e9};
test_input[30608:30615] = '{32'h3f8f7af4, 32'hc294291d, 32'hc2b37e3f, 32'hc1d31a83, 32'hc2374d93, 32'h3f76c724, 32'hc1f85c4b, 32'h41ec4fae};
test_weights[30608:30615] = '{32'h418f3392, 32'h425135b6, 32'hc2292da6, 32'h428b3d09, 32'h41c78564, 32'hc17d8339, 32'h419d135d, 32'h419005ba};
test_bias[3826:3826] = '{32'hc26a3179};
test_output[3826:3826] = '{32'hc547652b};
test_input[30616:30623] = '{32'hc2c4e384, 32'h42af64c6, 32'hc2b38b91, 32'h42bf5d2e, 32'hc221b352, 32'hc22ff408, 32'h42b79f43, 32'hc26913c5};
test_weights[30616:30623] = '{32'h4231c625, 32'h420039bc, 32'hc2330368, 32'h422ca9b5, 32'h42587ba0, 32'hc29027d6, 32'h4254cc4f, 32'hc2882434};
test_bias[3827:3827] = '{32'hc1eec048};
test_output[3827:3827] = '{32'h468006f2};
test_input[30624:30631] = '{32'hc262b22e, 32'hc27fec82, 32'hc256be16, 32'h42073982, 32'h40f254fc, 32'hc240df35, 32'h4291ca04, 32'h427dc344};
test_weights[30624:30631] = '{32'hc1e6f7de, 32'h42ad54c1, 32'h42889c50, 32'hc2bea635, 32'h41b96336, 32'hc2a9b355, 32'hc1e43603, 32'hc28b48f6};
test_bias[3828:3828] = '{32'hc229b0f1};
test_output[3828:3828] = '{32'hc64c3df8};
test_input[30632:30639] = '{32'hc290b04f, 32'hc29f29b7, 32'hc225a5ce, 32'h42a6d8db, 32'hc1c6c7ea, 32'hc2c2a949, 32'h428c50e5, 32'hc23a70c0};
test_weights[30632:30639] = '{32'hc1ea03ee, 32'h4200c162, 32'hc2066d11, 32'hc100b3a6, 32'h421c2d0a, 32'hc285dbf6, 32'hc27fb7c0, 32'hc217b381};
test_bias[3829:3829] = '{32'hc25479fb};
test_output[3829:3829] = '{32'h453e8cfb};
test_input[30640:30647] = '{32'hc29fd9f3, 32'hc29d1e50, 32'hc2996ab1, 32'h4255a775, 32'h41bc3332, 32'h42adc580, 32'h4272229e, 32'h42a014d7};
test_weights[30640:30647] = '{32'hc289efff, 32'hc2889308, 32'h42c328e2, 32'h42aa22eb, 32'hc20f21d2, 32'hc12811cc, 32'h4237b361, 32'hc18b7490};
test_bias[3830:3830] = '{32'hc13081b5};
test_output[3830:3830] = '{32'h45ec168b};
test_input[30648:30655] = '{32'h429a2b22, 32'hc2ae5452, 32'hc221c833, 32'h42a065f1, 32'hc281623b, 32'h42824fc5, 32'hc1b0afdb, 32'hc150073b};
test_weights[30648:30655] = '{32'hc295730f, 32'hc277c0cb, 32'h41bbcb1a, 32'hc282ffc2, 32'hc1814a67, 32'h4289e06d, 32'hc20a8912, 32'h424ce71a};
test_bias[3831:3831] = '{32'h429b8082};
test_output[3831:3831] = '{32'hc454740f};
test_input[30656:30663] = '{32'h424a186a, 32'h4290c234, 32'hc27e2c42, 32'hc181c95f, 32'h4289e8ce, 32'h41aa3ba1, 32'hc2a103d7, 32'h41ff32af};
test_weights[30656:30663] = '{32'hc25aa481, 32'hc29fa460, 32'hc26c8c1e, 32'hc2b0780d, 32'h4200876d, 32'h4228a425, 32'hc2920863, 32'h42accd39};
test_bias[3832:3832] = '{32'h429aa714};
test_output[3832:3832] = '{32'h46046b38};
test_input[30664:30671] = '{32'h41ee8e63, 32'hc188d0f6, 32'hc259c528, 32'h4089db84, 32'hc04dcc17, 32'hc29d3b04, 32'hc24aee78, 32'h42af8cd1};
test_weights[30664:30671] = '{32'h42a4d995, 32'hc11a9c99, 32'h409f7281, 32'h41a1aa2e, 32'h426ea4df, 32'h42a116d6, 32'h423b1be2, 32'h42a2da49};
test_bias[3833:3833] = '{32'h42af2225};
test_output[3833:3833] = '{32'h44422a58};
test_input[30672:30679] = '{32'h427007e8, 32'h42966196, 32'hc04991a9, 32'h41caac99, 32'h41f45539, 32'h41539b18, 32'hc25aa9ca, 32'hc21d4805};
test_weights[30672:30679] = '{32'hc1e79921, 32'hc1287334, 32'hc2360d89, 32'hc174e111, 32'h42615484, 32'hc1f19cb8, 32'hc12e4eaa, 32'h42394f6f};
test_bias[3834:3834] = '{32'h424df3aa};
test_output[3834:3834] = '{32'hc5242bf7};
test_input[30680:30687] = '{32'hc2bb9924, 32'hc2b847d0, 32'hc18b5565, 32'h41b21c85, 32'hc20438ac, 32'hc2002881, 32'h41ee73df, 32'h428d1362};
test_weights[30680:30687] = '{32'h428cfe93, 32'hc256b5f3, 32'hc1e9ef3b, 32'hc299bb07, 32'hc21ef791, 32'hc1a090b8, 32'h42153430, 32'hc2b4a1f0};
test_bias[3835:3835] = '{32'hc2836a1b};
test_output[3835:3835] = '{32'hc5c2e4d7};
test_input[30688:30695] = '{32'hc246e6a3, 32'hc255db14, 32'h42b5c5ff, 32'hc2102641, 32'h42adaa02, 32'h42287fe4, 32'h42359162, 32'hc12746ab};
test_weights[30688:30695] = '{32'hc2894b94, 32'hc2a4df56, 32'hc28d88e7, 32'hc10c6c43, 32'h42c22341, 32'hc29b81f0, 32'hc1daf9c8, 32'hc298db39};
test_bias[3836:3836] = '{32'hc2c72189};
test_output[3836:3836] = '{32'h45c55d5c};
test_input[30696:30703] = '{32'hc29ef818, 32'hc2b62d74, 32'hc2259248, 32'hc2717ae2, 32'h42608ba3, 32'hc0d89fd6, 32'h411a0a8d, 32'h42144733};
test_weights[30696:30703] = '{32'hc09be050, 32'hc2567783, 32'hc2b88aba, 32'hc28bbfd7, 32'hc23ed81b, 32'h427c5ed8, 32'h41cf182d, 32'h42aadbe0};
test_bias[3837:3837] = '{32'h4219c6ab};
test_output[3837:3837] = '{32'h4655674b};
test_input[30704:30711] = '{32'h42b4245b, 32'h41daba41, 32'hc2541295, 32'hc252c2eb, 32'hc22919c2, 32'h42adbda3, 32'hc1aba8a1, 32'h4181546e};
test_weights[30704:30711] = '{32'h411af0d9, 32'hc21272a4, 32'h42b1b69d, 32'hc26c60b9, 32'h4282d001, 32'h426f4256, 32'hc26c5f14, 32'h42be19eb};
test_bias[3838:3838] = '{32'hc265a1a6};
test_output[3838:3838] = '{32'h4557c2a9};
test_input[30712:30719] = '{32'h42989818, 32'hc265ef1c, 32'hc10ed690, 32'hc27fcbc3, 32'hc28d167a, 32'hc1a380ad, 32'hc29648df, 32'hc25fde71};
test_weights[30712:30719] = '{32'h4226f5a4, 32'hc21ef106, 32'hc25093fa, 32'hc164526c, 32'hc1cbf0ce, 32'hc095ccdf, 32'h42488b74, 32'h402da7f4};
test_bias[3839:3839] = '{32'hc09e623e};
test_output[3839:3839] = '{32'h4596858e};
test_input[30720:30727] = '{32'h42b43e98, 32'h425c92f6, 32'h42842d4f, 32'hc1f46697, 32'h42b7616d, 32'h3fc3b142, 32'h42069e0d, 32'hc2bd46b2};
test_weights[30720:30727] = '{32'h4234dbc7, 32'h41a0f783, 32'hc00f53c3, 32'hc2a4d229, 32'hc16ee8d7, 32'hc1a654c2, 32'hc25ba623, 32'h42aa8763};
test_bias[3840:3840] = '{32'h42546d39};
test_output[3840:3840] = '{32'hc567f0f8};
test_input[30728:30735] = '{32'hc27ca95f, 32'hc2b3ac51, 32'h42245b4c, 32'h42b8a42b, 32'hc1a4200b, 32'h3f6b17b1, 32'h4255fc11, 32'hc086fa88};
test_weights[30728:30735] = '{32'hc201db5d, 32'h429cd593, 32'h42b5734c, 32'hc2929ca1, 32'hc2ac9088, 32'hbffb6b0f, 32'h421c4f7b, 32'hc2b19d00};
test_bias[3841:3841] = '{32'h42635178};
test_output[3841:3841] = '{32'hc569fadd};
test_input[30736:30743] = '{32'hc2aeb46e, 32'hc2678d0b, 32'h4246dedc, 32'h427acced, 32'h425c0a53, 32'h42a94f8f, 32'hc1a0bb4f, 32'h422691cc};
test_weights[30736:30743] = '{32'hc2bf8d12, 32'hc27ac7e9, 32'h410bd21f, 32'hc23f1319, 32'h42bbced7, 32'hc10b754a, 32'h42bf36e3, 32'hc218e3d8};
test_bias[3842:3842] = '{32'h423bb0c0};
test_output[3842:3842] = '{32'h46227424};
test_input[30744:30751] = '{32'hc2778a71, 32'h42a52d80, 32'hc0a51a69, 32'hc0a798d4, 32'h42c23dee, 32'h428f87ea, 32'hc24b2343, 32'h42347abe};
test_weights[30744:30751] = '{32'h4284426f, 32'hc29fb520, 32'h41c71c02, 32'hc2b537ba, 32'h40cd918e, 32'hc25a00a6, 32'hc2b80fba, 32'hc12d5423};
test_bias[3843:3843] = '{32'h41812cc5};
test_output[3843:3843] = '{32'hc6134e6f};
test_input[30752:30759] = '{32'hc20e3c37, 32'hc24731a5, 32'hc02520bb, 32'h40934275, 32'h42a81d4d, 32'h4280aa52, 32'h4253b0ca, 32'hc22f35ff};
test_weights[30752:30759] = '{32'hc2097d79, 32'h4143a0fe, 32'hc288d28d, 32'h407b9d9d, 32'hc29f40c0, 32'hc2630b46, 32'h41953867, 32'h41fb21bb};
test_bias[3844:3844] = '{32'hc0bcd4c2};
test_output[3844:3844] = '{32'hc61b2a59};
test_input[30760:30767] = '{32'h425557de, 32'hc2818d8a, 32'h41e7f837, 32'h414c0bcf, 32'hc20a11d1, 32'hc19c2b5c, 32'h40fed101, 32'hc09f96e2};
test_weights[30760:30767] = '{32'hc1ada1e1, 32'hc23c1df0, 32'h41e89c97, 32'hc2c74325, 32'hc246ca26, 32'hc2c5c1ff, 32'h41c96c30, 32'h429acb9e};
test_bias[3845:3845] = '{32'h41efc3f2};
test_output[3845:3845] = '{32'h459abb72};
test_input[30768:30775] = '{32'h40e5afac, 32'h42a0abaf, 32'h41c29b2c, 32'h4154dae6, 32'h41e4a6dd, 32'h42b3e152, 32'hc257211f, 32'hc0bc05ee};
test_weights[30768:30775] = '{32'h419a5788, 32'h42494f7b, 32'hc2893b14, 32'hc2a49680, 32'hc280bdd8, 32'hc1de4817, 32'hbffc352f, 32'hc1b31bd3};
test_bias[3846:3846] = '{32'hc284f76b};
test_output[3846:3846] = '{32'hc52be215};
test_input[30776:30783] = '{32'h4231a160, 32'h427f55e0, 32'h420af8b1, 32'h4235b5db, 32'hc25a7def, 32'h42b76695, 32'h4144f989, 32'hc24fb645};
test_weights[30776:30783] = '{32'h422d88fd, 32'hc28ba4f8, 32'hc2387c2e, 32'h427d6423, 32'hc2a64a45, 32'h4237d826, 32'hc1559d55, 32'hc0de5f54};
test_bias[3847:3847] = '{32'h42ba3591};
test_output[3847:3847] = '{32'h45f37637};
test_input[30784:30791] = '{32'hc2b0842a, 32'hc2b9c932, 32'h426c577f, 32'hc1b59bac, 32'h426807c0, 32'h41e1f301, 32'hc0f5b8bb, 32'h41c56880};
test_weights[30784:30791] = '{32'h4248dcf7, 32'h428a0c70, 32'h423da78d, 32'hc207edc2, 32'h41416a66, 32'h41da652b, 32'hc0f8c9ac, 32'h429e8764};
test_bias[3848:3848] = '{32'h42be473a};
test_output[3848:3848] = '{32'hc5667e8c};
test_input[30792:30799] = '{32'h4248425d, 32'h4241fdc5, 32'hc19ca27b, 32'hc2689377, 32'h42813083, 32'hc253d381, 32'hc1175e25, 32'hc1cf0e4c};
test_weights[30792:30799] = '{32'h429e8930, 32'h4291f8dd, 32'h42c3be59, 32'hc175e703, 32'h408b1283, 32'h40e9dd70, 32'h408ccc39, 32'hc2a30787};
test_bias[3849:3849] = '{32'h42954d8b};
test_output[3849:3849] = '{32'h4605282a};
test_input[30800:30807] = '{32'h40dd50a8, 32'hc18ccf5d, 32'hc04a17f2, 32'hc2547b50, 32'h4278ef9d, 32'h41826002, 32'h42035ff9, 32'hc286caae};
test_weights[30800:30807] = '{32'hc1bb0cfa, 32'h4257cefe, 32'hc0ae7cea, 32'hc29816c9, 32'hc2c14ca8, 32'h42280442, 32'hc2b17b7c, 32'h41c6ebcf};
test_bias[3850:3850] = '{32'hc2ada569};
test_output[3850:3850] = '{32'hc5dcb174};
test_input[30808:30815] = '{32'hc281cc74, 32'h42b9449d, 32'h42bc508c, 32'h423e6f33, 32'hc2c38bc8, 32'h42ba43f5, 32'hc2b593af, 32'h42bda0b4};
test_weights[30808:30815] = '{32'h4267a25a, 32'hc0d92ae0, 32'h41c646ba, 32'h42c023f9, 32'h41423069, 32'hc2b4210b, 32'hc11f18cf, 32'h422945bb};
test_bias[3851:3851] = '{32'hc18b06cb};
test_output[3851:3851] = '{32'hc506c5ab};
test_input[30816:30823] = '{32'h4161ecd4, 32'h41552b12, 32'h4220d6a2, 32'h4244644b, 32'hc15d2174, 32'hc29453ea, 32'hc2aeed34, 32'hc2ac9ad6};
test_weights[30816:30823] = '{32'h42462b31, 32'h42998e82, 32'h4210f24a, 32'hc2101cd9, 32'hc2af110e, 32'hc29f272b, 32'h42c07ddc, 32'hc0dd2469};
test_bias[3852:3852] = '{32'hc21529a3};
test_output[3852:3852] = '{32'h4425cf1e};
test_input[30824:30831] = '{32'h41ff93c1, 32'h42b4882a, 32'hc20525ee, 32'h4016f399, 32'h414c35ef, 32'h429d1a54, 32'hc1510a7c, 32'hc2b1a5c9};
test_weights[30824:30831] = '{32'h427b5258, 32'hc25622a7, 32'hc23440e4, 32'hc2b22afe, 32'h41d3c45a, 32'h42392ec1, 32'h42abcc82, 32'hc205d8a0};
test_bias[3853:3853] = '{32'hc12c4424};
test_output[3853:3853] = '{32'h4585b3a7};
test_input[30832:30839] = '{32'hc1075530, 32'hc27be757, 32'h422c316d, 32'hc29ce39e, 32'h4138a01d, 32'h41f62413, 32'hc2c488ef, 32'hc1a65805};
test_weights[30832:30839] = '{32'hc28b1b9d, 32'hc20a37df, 32'hc2b8a403, 32'hc184f0a1, 32'hc2555436, 32'hc2ae365c, 32'h42a98d5d, 32'h428aab4c};
test_bias[3854:3854] = '{32'hc2bee61d};
test_output[3854:3854] = '{32'hc64c364a};
test_input[30840:30847] = '{32'hc2372f9e, 32'h41c4f5bc, 32'h40d1fbd3, 32'h419b0d21, 32'h428ea1f1, 32'h41141be7, 32'hc1ecabe8, 32'h414ba1e0};
test_weights[30840:30847] = '{32'h429d4824, 32'hc28a9455, 32'h425ced66, 32'hc284bc54, 32'hc2ba95b5, 32'h41d2e064, 32'h42878cfa, 32'h41fdf2bf};
test_bias[3855:3855] = '{32'hc1f141d6};
test_output[3855:3855] = '{32'hc65efef7};
test_input[30848:30855] = '{32'hc20e478e, 32'hc1066b3e, 32'h429d0bc8, 32'h427eaa32, 32'h4237be84, 32'h40dfa764, 32'hc24867af, 32'hc2b5577a};
test_weights[30848:30855] = '{32'hc2bee9c0, 32'h42c662d2, 32'h4287fa44, 32'h42c1b339, 32'h42bdc8a4, 32'h42a4bcc5, 32'hc117d34e, 32'hc13ddf59};
test_bias[3856:3856] = '{32'h429ba1dd};
test_output[3856:3856] = '{32'h46a12d58};
test_input[30856:30863] = '{32'hc270de84, 32'h4261de21, 32'hc287c37f, 32'hc0aa4e34, 32'hc2b2b10c, 32'hc1d5a0da, 32'h422bbcb3, 32'hc27ee41d};
test_weights[30856:30863] = '{32'hc225b982, 32'h42a34853, 32'h42aa7dc2, 32'h4203fb0a, 32'h42c0644a, 32'h41c3e8a2, 32'h427d76d8, 32'h4228556e};
test_bias[3857:3857] = '{32'h41d6aee7};
test_output[3857:3857] = '{32'hc5fb41be};
test_input[30864:30871] = '{32'h41865027, 32'h41fc19a4, 32'h4299962e, 32'h41e4633e, 32'h421fd7d8, 32'h4238701a, 32'hc1f945da, 32'hc28bf5ab};
test_weights[30864:30871] = '{32'hc28ce0dc, 32'hc2ac6d8a, 32'hc2800652, 32'hc1885f51, 32'h40f55630, 32'hc15b803e, 32'h3fdf15d2, 32'hc239a2ed};
test_bias[3858:3858] = '{32'h4203ae06};
test_output[3858:3858] = '{32'hc5c80d7d};
test_input[30872:30879] = '{32'hc21ea78b, 32'h41e9196f, 32'h4229de70, 32'hc1e0fdbe, 32'h42108031, 32'hc2054d86, 32'hc1365ead, 32'h3f798241};
test_weights[30872:30879] = '{32'h41b4cd2f, 32'hc146fe31, 32'hc28d9c58, 32'h427d5966, 32'hc240a3d5, 32'h428a69d5, 32'h40002726, 32'h416f755d};
test_bias[3859:3859] = '{32'hc2820530};
test_output[3859:3859] = '{32'hc61ed98b};
test_input[30880:30887] = '{32'h42bb32ee, 32'h42a00561, 32'hc2b97768, 32'h4293b9e9, 32'hc1c123ba, 32'hc2611a7c, 32'h4294c1f9, 32'h411b2166};
test_weights[30880:30887] = '{32'hc1c57e3c, 32'h42bd00d6, 32'h40dd925d, 32'h42c699f2, 32'h429cb944, 32'h42299706, 32'h41f8e1ad, 32'hc218e306};
test_bias[3860:3860] = '{32'h421e100f};
test_output[3860:3860] = '{32'h4616c065};
test_input[30888:30895] = '{32'h428818d6, 32'h4243fcfd, 32'h41bfe92d, 32'h40e66700, 32'h40e4c666, 32'h42004567, 32'hc193bb9d, 32'hc1cf2005};
test_weights[30888:30895] = '{32'h42a7994e, 32'h42be257e, 32'h426861ce, 32'hc0c486f6, 32'h4107e737, 32'hc130eb00, 32'hc23073cc, 32'hc0716d6e};
test_bias[3861:3861] = '{32'h41d8db5c};
test_output[3861:3861] = '{32'h46410ec5};
test_input[30896:30903] = '{32'h41ee4658, 32'h42a3ec42, 32'hc1b60578, 32'hc2b6cf3d, 32'h42866ebb, 32'hc2b2e7c9, 32'h42be99ba, 32'hc289543d};
test_weights[30896:30903] = '{32'h4203b8b7, 32'hc21f9ff3, 32'h42b26e60, 32'hc29e134f, 32'h42c140c6, 32'h423fa8d6, 32'h41ab75de, 32'hc268f872};
test_bias[3862:3862] = '{32'hc27a4084};
test_output[3862:3862] = '{32'h462d51fc};
test_input[30904:30911] = '{32'h41d98cb7, 32'hc26214a1, 32'h41b6b999, 32'hc293c445, 32'h420cf8ac, 32'h42c64b7f, 32'hc2a9aa74, 32'hc2b720e6};
test_weights[30904:30911] = '{32'hc2157516, 32'hc28d05bd, 32'h41789545, 32'hc28d0728, 32'h42c147ea, 32'h42827935, 32'h42bc9ec3, 32'hc1e2935e};
test_bias[3863:3863] = '{32'h41ad7d5d};
test_output[3863:3863] = '{32'h464b78d2};
test_input[30912:30919] = '{32'hc21684a2, 32'h414529de, 32'h416ba19a, 32'h41cd969a, 32'hc2716795, 32'hc049c564, 32'h429b32b8, 32'h424812b2};
test_weights[30912:30919] = '{32'h4274ad1e, 32'h40d5883a, 32'hc22a4d5c, 32'hc2680652, 32'hc0df75e9, 32'hc2c70882, 32'h4106e3ab, 32'hc2176f6a};
test_bias[3864:3864] = '{32'h40d68790};
test_output[3864:3864] = '{32'hc5971608};
test_input[30920:30927] = '{32'hc2c4f907, 32'h415a41a2, 32'hc2281726, 32'hc1cfa84d, 32'hc14d33a1, 32'hc2757773, 32'hc236139d, 32'hc2a001ee};
test_weights[30920:30927] = '{32'hc29a3529, 32'h41104a58, 32'hc23a113b, 32'hc2afd75f, 32'h4217adf4, 32'h426c879b, 32'h42a63339, 32'hc25132dc};
test_bias[3865:3865] = '{32'h42b508bf};
test_output[3865:3865] = '{32'h46022a55};
test_input[30928:30935] = '{32'hc28446d1, 32'h41ba74e9, 32'hc183d487, 32'hc2c326ee, 32'h417877cc, 32'hc204e007, 32'hc2bccc2d, 32'h41c4f5b8};
test_weights[30928:30935] = '{32'hc2a6443e, 32'hc12fd15e, 32'hc215df40, 32'h42929db4, 32'h3e357f81, 32'h420793f0, 32'h4190d78d, 32'h4185b007};
test_bias[3866:3866] = '{32'hc2b4853c};
test_output[3866:3866] = '{32'hc56dca04};
test_input[30936:30943] = '{32'h4281b506, 32'h42a8405e, 32'h429014c2, 32'hc2b78732, 32'hc29fb107, 32'h428cc269, 32'hc25ccceb, 32'hc23210a1};
test_weights[30936:30943] = '{32'hc2afa324, 32'hc262b02f, 32'h41b99193, 32'hc23030bb, 32'hc2399551, 32'h42332834, 32'h42157b74, 32'h42bd4e59};
test_bias[3867:3867] = '{32'hc267f8a4};
test_output[3867:3867] = '{32'hc5841c8d};
test_input[30944:30951] = '{32'hc1fd2570, 32'hc1100eb7, 32'h427bc457, 32'hc092f6ff, 32'h42920c56, 32'hc1869cf6, 32'hc18a1206, 32'h41acdaab};
test_weights[30944:30951] = '{32'hc2279319, 32'h4215382b, 32'hc25f96d8, 32'h421a02fb, 32'hc2890c1b, 32'h42b47073, 32'hc2a9ef19, 32'hc2295556};
test_bias[3868:3868] = '{32'hc234f89a};
test_output[3868:3868] = '{32'hc6084334};
test_input[30952:30959] = '{32'h4106e2ca, 32'hc25a9d99, 32'hc2c5cab1, 32'h41955338, 32'h42853952, 32'h3fe9efe2, 32'hc2ad2e12, 32'h416ae277};
test_weights[30952:30959] = '{32'hc28e06c3, 32'hc232ded3, 32'h40aa18ee, 32'hc21d441b, 32'hc0ceb5fd, 32'h42021cc9, 32'h41a41568, 32'h4248b6f6};
test_bias[3869:3869] = '{32'hc1dfb098};
test_output[3869:3869] = '{32'hc455196d};
test_input[30960:30967] = '{32'hc0f76e2e, 32'hc28e435e, 32'hc22bf07a, 32'hc22d8c80, 32'hc1c9ed83, 32'h426f37b4, 32'h40e8f2ca, 32'h420b0af3};
test_weights[30960:30967] = '{32'hc2456876, 32'h42a7d2f0, 32'hc2983bcc, 32'hc27a047e, 32'hc262ea6d, 32'h42be2f3a, 32'h42040dd9, 32'h42161916};
test_bias[3870:3870] = '{32'hc1ce8f56};
test_output[3870:3870] = '{32'h460d291c};
test_input[30968:30975] = '{32'hc2156422, 32'h41e3e970, 32'h425690ed, 32'hc232b637, 32'hc224c503, 32'hc21e48a0, 32'h4268d9ca, 32'h411869d3};
test_weights[30968:30975] = '{32'h426839f5, 32'h42c520a8, 32'hc107b07b, 32'h42bdb6f6, 32'hc1ae2b30, 32'hc291f886, 32'h416ce7b8, 32'h42a75e96};
test_bias[3871:3871] = '{32'hc0ec28a5};
test_output[3871:3871] = '{32'h44acebf6};
test_input[30976:30983] = '{32'hc2b76c0b, 32'hc27ade1e, 32'h42a3abcc, 32'hc0e3179d, 32'h42be1a92, 32'hc220d029, 32'hc1d31d2b, 32'h41bf9e6d};
test_weights[30976:30983] = '{32'hc2438b71, 32'h421c17c8, 32'hc258c2e8, 32'hc294b32f, 32'hc29ef1dd, 32'hc21214d9, 32'hc2bc8b17, 32'hc20eda16};
test_bias[3872:3872] = '{32'h408798aa};
test_output[3872:3872] = '{32'hc5c58208};
test_input[30984:30991] = '{32'h40af6017, 32'h41b444ef, 32'h42a67758, 32'h42addc8e, 32'h41b1949b, 32'h4248dbc8, 32'hc2ab50d0, 32'h42a75ace};
test_weights[30984:30991] = '{32'hc2278b07, 32'h41c2a6eb, 32'h41a05649, 32'h429e9437, 32'h429e7da5, 32'hc18497f5, 32'hc20b149b, 32'h42bd96fc};
test_bias[3873:3873] = '{32'h42b4c8fc};
test_output[3873:3873] = '{32'h46a28e93};
test_input[30992:30999] = '{32'h426932fc, 32'h42a708c8, 32'h429c3830, 32'hc238feef, 32'h4231488a, 32'h41729f58, 32'h427b107d, 32'h424c726c};
test_weights[30992:30999] = '{32'h427a412e, 32'h4201ce56, 32'hc2baff59, 32'h422e9cb3, 32'h4239aa71, 32'hc10cec63, 32'h42acc5fe, 32'h424c598e};
test_bias[3874:3874] = '{32'h42c3ebde};
test_output[3874:3874] = '{32'h45dd94a1};
test_input[31000:31007] = '{32'hc21692e0, 32'hc24f18b6, 32'hc2ad4647, 32'hc210d7d3, 32'h40052e03, 32'hc29ab4bb, 32'h41be180a, 32'hc1a5bc8e};
test_weights[31000:31007] = '{32'hc1373a71, 32'hc244143d, 32'hbf5c6687, 32'h4151d156, 32'hc1451916, 32'h42abe9f3, 32'h423dce58, 32'h42b5aa0f};
test_bias[3875:3875] = '{32'h42b1655c};
test_output[3875:3875] = '{32'hc5951b74};
test_input[31008:31015] = '{32'h41fcdff3, 32'hc2419f03, 32'h40b41fbe, 32'h42a1dbcc, 32'h424e02d4, 32'hc20e8849, 32'h424e4544, 32'hc25f68fb};
test_weights[31008:31015] = '{32'hc0c1cd92, 32'h40a612a6, 32'h42a10b81, 32'hc170cbb6, 32'h40bca736, 32'h3e2ba52f, 32'hc1a56231, 32'h41b1150f};
test_bias[3876:3876] = '{32'hc27ec3c5};
test_output[3876:3876] = '{32'hc54cbc37};
test_input[31016:31023] = '{32'hc1a982c8, 32'hc1fcc246, 32'h4284c8cb, 32'h4255cc0e, 32'hc214f28f, 32'hc10b83e6, 32'h42492ba4, 32'hc145c929};
test_weights[31016:31023] = '{32'h41c9c1c6, 32'h42ac168a, 32'h42511037, 32'hc23b1f87, 32'h428d764b, 32'h42783c32, 32'h421e3b11, 32'h429ea766};
test_bias[3877:3877] = '{32'h420efa78};
test_output[3877:3877] = '{32'hc589ecfa};
test_input[31024:31031] = '{32'hc1bda850, 32'hc238d48e, 32'h3f91b807, 32'hc0050a7b, 32'h416fc3d8, 32'h422d0203, 32'h42425a3b, 32'h42914f2c};
test_weights[31024:31031] = '{32'h42c16958, 32'hc2af902d, 32'h42b51747, 32'hc1f813f5, 32'h42a8ecde, 32'h403b0d3a, 32'h42a907ff, 32'h429c5edb};
test_bias[3878:3878] = '{32'hc2b031f8};
test_output[3878:3878] = '{32'h464b7856};
test_input[31032:31039] = '{32'h4291bcbd, 32'h3f9ca83b, 32'hc2c7f6b1, 32'hc2c2cf68, 32'h40516b00, 32'hc2932a35, 32'hc242336a, 32'h42a0761b};
test_weights[31032:31039] = '{32'hc2a75246, 32'h421c7502, 32'hc2c09b56, 32'h429afad0, 32'h3f54e24e, 32'hc181ec4b, 32'h429644ba, 32'h424dd2b8};
test_bias[3879:3879] = '{32'hc2bba467};
test_output[3879:3879] = '{32'hc514f3b6};
test_input[31040:31047] = '{32'hc2b369ab, 32'hc2af3e11, 32'h4182e89f, 32'h4205e035, 32'hc1502a99, 32'h42a1eddb, 32'h4134f146, 32'h42c56efd};
test_weights[31040:31047] = '{32'hc281b9a2, 32'h422e6113, 32'h42a74804, 32'hc0b34cd3, 32'hc22cbe95, 32'hc1fb18d7, 32'h418c0d45, 32'h421dd852};
test_bias[3880:3880] = '{32'h41eb7b4b};
test_output[3880:3880] = '{32'h45a65b4c};
test_input[31048:31055] = '{32'h40f493ad, 32'h42a31dff, 32'h42370a6c, 32'h411f4e37, 32'hc232705b, 32'h423e9463, 32'hc0e1c5ec, 32'hc2b5736e};
test_weights[31048:31055] = '{32'hc21a7f89, 32'hc2beb048, 32'h42c00f3a, 32'h41bcdb4d, 32'h42063310, 32'hc1a0ad76, 32'hc2c71a7c, 32'h429e2806};
test_bias[3881:3881] = '{32'h422bc6b8};
test_output[3881:3881] = '{32'hc640928b};
test_input[31056:31063] = '{32'hc25762f3, 32'hc2840c8c, 32'hc22ae4e9, 32'hc183f4a7, 32'h42908927, 32'hc29061e8, 32'h429a74d4, 32'hc1c04238};
test_weights[31056:31063] = '{32'h42c73a35, 32'hc1d857e0, 32'hc1adb3d0, 32'hc2a1709c, 32'h41ab237a, 32'h423d0ca1, 32'h4007f553, 32'h4293e148};
test_bias[3882:3882] = '{32'h4200f914};
test_output[3882:3882] = '{32'hc594ef11};
test_input[31064:31071] = '{32'hc03dabd6, 32'hc1d031a1, 32'h416ff325, 32'h42283047, 32'h427ba9cc, 32'hc100f962, 32'h42bcff9a, 32'hc216b06f};
test_weights[31064:31071] = '{32'h41d8f33e, 32'h42b881f8, 32'h42c6a7e6, 32'hc278a82c, 32'h4182b2bb, 32'h42368759, 32'hc1a63cbc, 32'hc10f55e6};
test_bias[3883:3883] = '{32'h41893b20};
test_output[3883:3883] = '{32'hc58e5349};
test_input[31072:31079] = '{32'h3f68c077, 32'h41bee407, 32'hc01ac7cc, 32'hc1837372, 32'h427a0214, 32'h42bf26e6, 32'h4230300f, 32'h4290a3fb};
test_weights[31072:31079] = '{32'hc1e996cd, 32'h42b1db7c, 32'hc2523261, 32'hc1599057, 32'hbfecf070, 32'h41f7ba54, 32'hc21ba4fa, 32'h4003116d};
test_bias[3884:3884] = '{32'hc0e8be7a};
test_output[3884:3884] = '{32'h45684c0f};
test_input[31080:31087] = '{32'h42ae36aa, 32'hc280c287, 32'h41ccae12, 32'h426cd631, 32'h42b3720d, 32'h4134de43, 32'hc2a5927d, 32'hc11fcbc1};
test_weights[31080:31087] = '{32'hc2a7a3a0, 32'hc1f5f58c, 32'h42677f7c, 32'h42a98f8f, 32'h429eee5d, 32'hc2c72f65, 32'hc29a155e, 32'h42926160};
test_bias[3885:3885] = '{32'hc10f3d06};
test_output[3885:3885] = '{32'h464852d7};
test_input[31088:31095] = '{32'hc164b405, 32'h3f88b3ca, 32'h41196253, 32'h42965493, 32'hc276f466, 32'h42399f80, 32'h425bf29d, 32'h42a7f2c6};
test_weights[31088:31095] = '{32'hc22eeabe, 32'hc2aa8c03, 32'hc2852bd3, 32'hc2c47129, 32'hc28eaf7f, 32'hc2c5b647, 32'hc209c7c1, 32'hc12df168};
test_bias[3886:3886] = '{32'h42334c6c};
test_output[3886:3886] = '{32'hc623008b};
test_input[31096:31103] = '{32'hc2b930ca, 32'hc2053b68, 32'hc18c2035, 32'hc17b3722, 32'h41da7b35, 32'h42c135aa, 32'h3f1730a2, 32'hc296debc};
test_weights[31096:31103] = '{32'h42af8008, 32'hc1e83363, 32'h42a0cc01, 32'h4243c33b, 32'h42494e59, 32'hbfd4414c, 32'hc15e9661, 32'h42944c18};
test_bias[3887:3887] = '{32'hc2c391bb};
test_output[3887:3887] = '{32'hc657f132};
test_input[31104:31111] = '{32'hc10f009b, 32'h423ab137, 32'h423e688f, 32'hc24c9314, 32'h42402244, 32'hc2a40e90, 32'hc2b5eee9, 32'h422faae1};
test_weights[31104:31111] = '{32'h41aae0e8, 32'hc28e0d8e, 32'h4111c950, 32'hc23fa94e, 32'hc229201c, 32'hc29a5dd5, 32'h424281e3, 32'h415a3d24};
test_bias[3888:3888] = '{32'h421b7bcd};
test_output[3888:3888] = '{32'hc2d5b542};
test_input[31112:31119] = '{32'hc2707072, 32'h41822746, 32'hc107d963, 32'h421ef7af, 32'hc1eac4e1, 32'h4293a574, 32'h4212c991, 32'h4197688a};
test_weights[31112:31119] = '{32'h4285d51b, 32'h41e9d87a, 32'hc1be99c9, 32'hc220844e, 32'h41824274, 32'hc171b579, 32'hc10435ee, 32'h420fb3d5};
test_bias[3889:3889] = '{32'h42bccf75};
test_output[3889:3889] = '{32'hc5bd69ea};
test_input[31120:31127] = '{32'hc29a7956, 32'hc2b98d97, 32'hc1168f98, 32'h410b7af0, 32'hc2bd9379, 32'hc2a16063, 32'hc28bede4, 32'h42b29d8a};
test_weights[31120:31127] = '{32'h42b09b5d, 32'h41abbafb, 32'hc1da1cfd, 32'hc283db78, 32'hc2aaaa8d, 32'hc098f126, 32'h4159c889, 32'h428b8772};
test_bias[3890:3890] = '{32'h42502adc};
test_output[3890:3890] = '{32'h4592132a};
test_input[31128:31135] = '{32'hc2846a31, 32'hc23524af, 32'h420eceb5, 32'h42a0a396, 32'h42aa9b30, 32'h4244c16d, 32'hc288e431, 32'h419d3c41};
test_weights[31128:31135] = '{32'hc2b4ef9e, 32'h4243eb85, 32'h429c20b7, 32'h420be3c4, 32'hc284db16, 32'h410f6188, 32'hc0baca79, 32'h418a0108};
test_bias[3891:3891] = '{32'hc1a86e29};
test_output[3891:3891] = '{32'h4597daeb};
test_input[31136:31143] = '{32'hc23d39e4, 32'h42a0a1bc, 32'h416aec7f, 32'hc2895141, 32'h41c5ad8d, 32'h4206e0cb, 32'h41889250, 32'h41b42b18};
test_weights[31136:31143] = '{32'hc2a25adf, 32'h40e0529c, 32'hc27e402a, 32'h40d20233, 32'hc2221d2d, 32'h424f8cbe, 32'h42159562, 32'hc09757a8};
test_bias[3892:3892] = '{32'hc20f7976};
test_output[3892:3892] = '{32'h45853c96};
test_input[31144:31151] = '{32'h3fbb1c6c, 32'h410a1704, 32'hc24a20cc, 32'h42bb69ee, 32'h42571581, 32'hc0c96ea2, 32'h3e99820c, 32'h42977afd};
test_weights[31144:31151] = '{32'hc0e8dfea, 32'hc168b885, 32'h42810a68, 32'hc292bd07, 32'h4234cf5d, 32'hc29b604d, 32'hc1147510, 32'h42569491};
test_bias[3893:3893] = '{32'hc2121d46};
test_output[3893:3893] = '{32'hc5500529};
test_input[31152:31159] = '{32'h429a39eb, 32'hc293b004, 32'h42c2602f, 32'hc287242c, 32'h426a26b1, 32'hc2848ec2, 32'hc2a315fb, 32'hc29dc709};
test_weights[31152:31159] = '{32'h41dc83b9, 32'h42508c17, 32'hc24db593, 32'hc151bed7, 32'hc159a26e, 32'hc26d2e20, 32'h4221d820, 32'hc2bd0992};
test_bias[3894:3894] = '{32'h42b35890};
test_output[3894:3894] = '{32'h44c0fb61};
test_input[31160:31167] = '{32'h4286a7c2, 32'h41a1d1b0, 32'h4277d8d3, 32'hc24f6471, 32'h42c66a52, 32'h40e9f4d0, 32'h421f0223, 32'hc2954040};
test_weights[31160:31167] = '{32'h42733b9c, 32'h4277ccd9, 32'h42714620, 32'h418092ca, 32'hc2c543b2, 32'h4296a30a, 32'hc0008ba5, 32'h42313fde};
test_bias[3895:3895] = '{32'h42a6d106};
test_output[3895:3895] = '{32'hc585f2e4};
test_input[31168:31175] = '{32'hc24b3149, 32'h422a8226, 32'hc20fa8d4, 32'h421193a3, 32'h427feddb, 32'h42c781a3, 32'h418673f7, 32'hc23e8c2b};
test_weights[31168:31175] = '{32'hc1e16e6a, 32'hc1c78864, 32'h41be3ac7, 32'h4216becf, 32'h4218fa55, 32'h423687df, 32'hc2196774, 32'hc29d4924};
test_bias[3896:3896] = '{32'hc280656c};
test_output[3896:3896] = '{32'h462aa950};
test_input[31176:31183] = '{32'h4283abb1, 32'hc2b1f356, 32'h42ab44de, 32'hc2066a2e, 32'h42192142, 32'hc2626062, 32'h4187c775, 32'hc29de844};
test_weights[31176:31183] = '{32'hc266010c, 32'h4251cf2d, 32'h42c674a1, 32'h4214679b, 32'hc16e4302, 32'hc2a8b732, 32'hc2c29d23, 32'h425a4639};
test_bias[3897:3897] = '{32'hc02e70d0};
test_output[3897:3897] = '{32'hc539089d};
test_input[31184:31191] = '{32'h428c5051, 32'hc2baa7c1, 32'hc184c139, 32'hc1fa1486, 32'hc2aeb21a, 32'h41bf36cc, 32'h41e2d409, 32'h4088bc6b};
test_weights[31184:31191] = '{32'hc1f69fbd, 32'hc2a56a8b, 32'h42acf9af, 32'hc2aaed34, 32'h4221a25a, 32'h4241948e, 32'hc2a99ce0, 32'hc2ab8b2f};
test_bias[3898:3898] = '{32'hc1ed0065};
test_output[3898:3898] = '{32'h44ca5f16};
test_input[31192:31199] = '{32'h41f02a9f, 32'h426f5825, 32'h424f62c1, 32'hc1d9ee16, 32'hc2c4fc72, 32'hc227a5ef, 32'h42a5a4a6, 32'h4274cf5e};
test_weights[31192:31199] = '{32'hc2be3d56, 32'h40480abe, 32'hc2a36745, 32'hc26c8c73, 32'h4182ef6a, 32'h41cbef4a, 32'h419bf823, 32'hc20c23c1};
test_bias[3899:3899] = '{32'h421b2cf2};
test_output[3899:3899] = '{32'hc60442c0};
test_input[31200:31207] = '{32'h41b51e9a, 32'h4285a702, 32'hc0d496ec, 32'hc046c8c1, 32'h40987bc1, 32'hc1063793, 32'hc29163b4, 32'hc2b0eb3a};
test_weights[31200:31207] = '{32'h408204fa, 32'hc1964c6a, 32'hc0959b84, 32'hc2baa4e8, 32'hc24706ad, 32'hc299c13f, 32'hc2bf944e, 32'h425e150d};
test_bias[3900:3900] = '{32'h42b43b88};
test_output[3900:3900] = '{32'h44d56d80};
test_input[31208:31215] = '{32'h42bdcfb6, 32'hc1315b71, 32'h41af5b72, 32'h42796a6d, 32'hc0df4966, 32'h4267998b, 32'hc2b7911b, 32'h4240e6f8};
test_weights[31208:31215] = '{32'hc2b46b01, 32'h42a5d904, 32'hbfda6e38, 32'hc2127a3c, 32'hc26e81da, 32'h428d265b, 32'h416751b0, 32'hc2b7a01e};
test_bias[3901:3901] = '{32'h42806af3};
test_output[3901:3901] = '{32'hc64af5ba};
test_input[31216:31223] = '{32'hc042ce11, 32'h4236d8ed, 32'h4108fdbc, 32'hc18525f4, 32'h428a8118, 32'h42ac6211, 32'h41dc2112, 32'h42344107};
test_weights[31216:31223] = '{32'h419d50f3, 32'hc218c40f, 32'h42b1f655, 32'hc1dd0e91, 32'hc2326691, 32'hc26f1533, 32'hc226d343, 32'h42516857};
test_bias[3902:3902] = '{32'h4286367d};
test_output[3902:3902] = '{32'hc5ebcd02};
test_input[31224:31231] = '{32'h41de512a, 32'h42a081d7, 32'hc256bfdc, 32'hc2afc201, 32'h4261fa53, 32'h42a5f792, 32'h42c775d0, 32'hc2717fd6};
test_weights[31224:31231] = '{32'hc25609e0, 32'hc28c78ea, 32'h416ca257, 32'hc2a97660, 32'h42640af9, 32'hc1bd152e, 32'h42aecd87, 32'h41c3faa9};
test_bias[3903:3903] = '{32'hc2c732d7};
test_output[3903:3903] = '{32'h45f7adcb};
test_input[31232:31239] = '{32'h424fb11c, 32'h42575e7e, 32'hc2ba4f12, 32'h419d504a, 32'h42b8b84f, 32'h41587906, 32'h416060a9, 32'hc252dad2};
test_weights[31232:31239] = '{32'h42896f1a, 32'hc233ce57, 32'hc25e29fc, 32'h42a2a118, 32'hc19dad52, 32'h422c9f46, 32'hc207a16b, 32'hc214b140};
test_bias[3904:3904] = '{32'h42a67d02};
test_output[3904:3904] = '{32'h4600ed5a};
test_input[31240:31247] = '{32'h4270efa1, 32'h41bd9694, 32'hc254eaa4, 32'h42a824df, 32'hc1bf50ef, 32'hc210322a, 32'h42555121, 32'hc2b88eca};
test_weights[31240:31247] = '{32'hc01f1379, 32'h42c026a4, 32'h42a45930, 32'hc28559d1, 32'hc2215970, 32'h41c30bc5, 32'h42a84f64, 32'h42a24fad};
test_bias[3905:3905] = '{32'hc150f0bd};
test_output[3905:3905] = '{32'hc6287338};
test_input[31248:31255] = '{32'h414ada64, 32'hc1c0addb, 32'h425cfae2, 32'h42895a21, 32'h41ff721d, 32'h42852366, 32'hc206f7aa, 32'h4197896c};
test_weights[31248:31255] = '{32'h4217aa54, 32'hc227837c, 32'h4218f2c7, 32'hc2863a77, 32'hc29e2209, 32'h425f3f2d, 32'h42b672c5, 32'hc201bc8a};
test_bias[3906:3906] = '{32'h41e0d58e};
test_output[3906:3906] = '{32'hc5599075};
test_input[31256:31263] = '{32'h4209201f, 32'hc2a2fa7d, 32'hc1db5ff7, 32'hc2a52cb9, 32'h41d6dfcc, 32'h42a72f55, 32'h42c05570, 32'h42a633ce};
test_weights[31256:31263] = '{32'hc151b400, 32'h42af9d80, 32'hc29eeb89, 32'h41a5d3c0, 32'hc1309f73, 32'hc2b2e16f, 32'h425c77c5, 32'h41fd5631};
test_bias[3907:3907] = '{32'h42b249c9};
test_output[3907:3907] = '{32'hc5d74c43};
test_input[31264:31271] = '{32'hc233ad0e, 32'hc211fd56, 32'h429359b2, 32'hc1a8368a, 32'h4291fd49, 32'h42c2689c, 32'hc220cfa8, 32'hc1e830b0};
test_weights[31264:31271] = '{32'hc2909a48, 32'hc2286767, 32'hc1993d3d, 32'h4280ce11, 32'hc28ae773, 32'hc26c4f42, 32'hc2147a77, 32'h429e9f47};
test_bias[3908:3908] = '{32'hc29dde53};
test_output[3908:3908] = '{32'hc6174779};
test_input[31272:31279] = '{32'hc225ffe5, 32'hc1518b22, 32'hc1aee4cb, 32'h4245341e, 32'h4104fb22, 32'h4274569a, 32'h4210c8db, 32'hc2adad71};
test_weights[31272:31279] = '{32'hc236addf, 32'h42541d23, 32'h41d237a5, 32'h4204f0ec, 32'hc2024ec6, 32'h414abfbd, 32'hc2432ff7, 32'h415dd30c};
test_bias[3909:3909] = '{32'h42762404};
test_output[3909:3909] = '{32'hc30c7d86};
test_input[31280:31287] = '{32'h4296afa0, 32'hc2853e69, 32'hc261eda3, 32'h429651e2, 32'hc285d4c4, 32'h41bb0c72, 32'hc26ff0e8, 32'hc228f4ad};
test_weights[31280:31287] = '{32'h42511122, 32'hc25ad7b6, 32'hc1885a9f, 32'hc1bb5264, 32'hc2916ed7, 32'h422f2c6f, 32'h428635ad, 32'h42b17a64};
test_bias[3910:3910] = '{32'h4219be22};
test_output[3910:3910] = '{32'h459a62e2};
test_input[31288:31295] = '{32'hc2a8839e, 32'hc257d0d2, 32'hc185ad1f, 32'hc2bd3ba6, 32'h40ea9474, 32'hc063b958, 32'h42c1bdfa, 32'h41d1b544};
test_weights[31288:31295] = '{32'h42346684, 32'h421bdac4, 32'hc2622839, 32'hc29a7ed6, 32'h422c3465, 32'h4183b599, 32'hc27beb15, 32'h42175510};
test_bias[3911:3911] = '{32'h4232712d};
test_output[3911:3911] = '{32'hc519820d};
test_input[31296:31303] = '{32'h41780313, 32'h4219a4f8, 32'h42782061, 32'hc13a8424, 32'h42026bd1, 32'h42aad6cd, 32'h427d0daa, 32'hc1198a9e};
test_weights[31296:31303] = '{32'hc16f2ee4, 32'h40818c97, 32'hc2266218, 32'hc24dcd7b, 32'h42318358, 32'hc28476aa, 32'h420f436b, 32'h429d1d4c};
test_bias[3912:3912] = '{32'h4223dc2b};
test_output[3912:3912] = '{32'hc5935246};
test_input[31304:31311] = '{32'h4247d57c, 32'hc295cd53, 32'hc0f73058, 32'h425f7ea6, 32'hc2bb051e, 32'hc2ae0f7f, 32'h42a346fe, 32'hc2b48026};
test_weights[31304:31311] = '{32'hc1b73917, 32'hc23adcd4, 32'h429fa1a8, 32'h422a994c, 32'hc257328b, 32'hc2412782, 32'h4132af3a, 32'hc2839f31};
test_bias[3913:3913] = '{32'h40bf4587};
test_output[3913:3913] = '{32'h469de79c};
test_input[31312:31319] = '{32'hc2a766a6, 32'hc2a7da30, 32'h4255fb18, 32'hc2695ba3, 32'h42a04f04, 32'hc2a44a23, 32'hc285da64, 32'h428704a4};
test_weights[31312:31319] = '{32'h42995561, 32'hc20811de, 32'h42958db1, 32'h42508f88, 32'hc1961714, 32'h41901fa6, 32'hc2b0f988, 32'hc2b4412a};
test_bias[3914:3914] = '{32'h41888aca};
test_output[3914:3914] = '{32'hc5b324ab};
test_input[31320:31327] = '{32'hc2566208, 32'h42b18f92, 32'h428bdd97, 32'hc26668bb, 32'h42b4d68c, 32'hc2a0f592, 32'h42a4740a, 32'hc2a7a6ab};
test_weights[31320:31327] = '{32'hc0c17bff, 32'h418d14fb, 32'h41ddbac5, 32'h4293d69d, 32'h42a1d783, 32'hc2915155, 32'hc22b69a9, 32'hc29bb841};
test_bias[3915:3915] = '{32'hc2081dfd};
test_output[3915:3915] = '{32'h46755d80};
test_input[31328:31335] = '{32'h42bb8a89, 32'h4279c465, 32'hc16b5916, 32'hc283f6b0, 32'h41a48abb, 32'h42984499, 32'hc2c1f8c7, 32'h42b2630e};
test_weights[31328:31335] = '{32'hc2a8e4b2, 32'h425bcae3, 32'hc1e8394a, 32'hc2b907a9, 32'h42855b78, 32'hc2b84ac3, 32'h411f53a9, 32'hc0e006a0};
test_bias[3916:3916] = '{32'hc1a8381a};
test_output[3916:3916] = '{32'hc5a2dc20};
test_input[31336:31343] = '{32'hc21be40b, 32'h42bf3a8d, 32'h41fc17b8, 32'hc2afc0dc, 32'h428c4952, 32'h4287770a, 32'h42890f0f, 32'hc1ce9317};
test_weights[31336:31343] = '{32'h410083aa, 32'h423b7986, 32'hc25b88d3, 32'h420bdf40, 32'h4016bde3, 32'h42973584, 32'hc241e8e8, 32'h42a0ed8e};
test_bias[3917:3917] = '{32'hc2a71f71};
test_output[3917:3917] = '{32'hc44fd884};
test_input[31344:31351] = '{32'hc027cceb, 32'h42b12787, 32'h42a1aa67, 32'h410859c0, 32'hc248ae04, 32'h4201080c, 32'hc263753f, 32'hc221497c};
test_weights[31344:31351] = '{32'hc19e8da6, 32'hc29ec9f7, 32'hc1624458, 32'hc276718e, 32'hc1afd0e8, 32'h429ebfad, 32'h428cddaa, 32'h42a82271};
test_bias[3918:3918] = '{32'h42b5a46c};
test_output[3918:3918] = '{32'hc6400702};
test_input[31352:31359] = '{32'h42b06374, 32'hc2b1b479, 32'hc2835c27, 32'h42c285c1, 32'h41fe3e4c, 32'hc28ed576, 32'hc1b1a9b8, 32'hc24ef1bb};
test_weights[31352:31359] = '{32'hc2a997ff, 32'hc142a698, 32'hc06aa1f3, 32'h421cd5dc, 32'hc01e7ffc, 32'h427de8a4, 32'hc2a8fc73, 32'h424dd28d};
test_bias[3919:3919] = '{32'hc2c50882};
test_output[3919:3919] = '{32'hc5f4fcf6};
test_input[31360:31367] = '{32'h42b7bcd6, 32'hc0b3cc90, 32'h429e9c8f, 32'h4263eaa6, 32'hc1e5294c, 32'hc2be3b95, 32'h41acb34f, 32'h412a323f};
test_weights[31360:31367] = '{32'hc19543ff, 32'hc0a7dd63, 32'hc2b61237, 32'h42586e39, 32'h42955f9f, 32'hc201bba2, 32'h42c771ef, 32'h42a75232};
test_bias[3920:3920] = '{32'hc1cb7a95};
test_output[3920:3920] = '{32'hc4e85027};
test_input[31368:31375] = '{32'hc28b4163, 32'h42c3fd2c, 32'hc2b43991, 32'h428f5fdb, 32'hc27335e1, 32'hc10a5768, 32'h42971651, 32'hc288183f};
test_weights[31368:31375] = '{32'hc1c3967b, 32'h40b2154d, 32'h4204bfb2, 32'h3fa8b763, 32'hc1d320d7, 32'h4290cfb3, 32'h42c4e718, 32'h42bf6f3d};
test_bias[3921:3921] = '{32'hc192d1c6};
test_output[3921:3921] = '{32'h449a7b8d};
test_input[31376:31383] = '{32'h428c8c9e, 32'h41c0ccc0, 32'h41ce7d61, 32'h42b34355, 32'h4225d1ab, 32'hc1b25756, 32'hc2bb60b8, 32'h422a1bad};
test_weights[31376:31383] = '{32'hc1f57a3a, 32'hc2370ece, 32'h412e63b4, 32'h41a9c45f, 32'hc1e3ad2a, 32'hc17b5550, 32'hc2aae7fd, 32'h4299d50d};
test_bias[3922:3922] = '{32'h4125c9f7};
test_output[3922:3922] = '{32'h4612978c};
test_input[31384:31391] = '{32'h422e1aac, 32'h41ba2ae0, 32'h41df6adb, 32'hc2935d87, 32'hc0e2bf7b, 32'hc2944689, 32'h429ffdbd, 32'h42907ece};
test_weights[31384:31391] = '{32'hc2a7c9a3, 32'hc1e6d2ae, 32'h4271ce4f, 32'hc2b0e797, 32'hc23ff049, 32'h41d25607, 32'hc2aa9659, 32'h420b7bb6};
test_bias[3923:3923] = '{32'hc1a3e5f0};
test_output[3923:3923] = '{32'hc5002d7a};
test_input[31392:31399] = '{32'h42a9e70b, 32'h423c8715, 32'hc2a495c7, 32'hc0291de5, 32'hc29bf032, 32'h424de85f, 32'hc083cfb2, 32'hc211cb46};
test_weights[31392:31399] = '{32'h41baf632, 32'h425c5a19, 32'hc2c22c34, 32'hc2bf3c33, 32'hc2442fa2, 32'h423df0c2, 32'hc285efd6, 32'hc2516f77};
test_bias[3924:3924] = '{32'hc29ae257};
test_output[3924:3924] = '{32'h46a59e60};
test_input[31400:31407] = '{32'h4120a581, 32'hc27653fd, 32'h42423bb7, 32'h4287cbf9, 32'hc246b42d, 32'hc2b19a65, 32'h42b1744a, 32'hc15e1434};
test_weights[31400:31407] = '{32'hc26a4af4, 32'h42b94271, 32'hc20cad7f, 32'hc1087754, 32'h42b7f92c, 32'hc259b216, 32'hc28b77f4, 32'hc1ca5f96};
test_bias[3925:3925] = '{32'hc1dcd550};
test_output[3925:3925] = '{32'hc65d8ede};
test_input[31408:31415] = '{32'hc2be3287, 32'h42a85cc6, 32'hc2c473de, 32'h427c9670, 32'hc28a4ddd, 32'h41e05ec8, 32'h4234b723, 32'h42387975};
test_weights[31408:31415] = '{32'hc29b90e7, 32'hc2aa210d, 32'hc1644547, 32'h42763949, 32'hc1e845c8, 32'h429f8e90, 32'hc24f92f2, 32'hc241da8e};
test_bias[3926:3926] = '{32'hc2948ced};
test_output[3926:3926] = '{32'h459fe0d9};
test_input[31416:31423] = '{32'h41c92618, 32'hc248223f, 32'hc2be2b6e, 32'h4200f60e, 32'h428c1676, 32'h410e74c7, 32'hc28d12c6, 32'h428d9052};
test_weights[31416:31423] = '{32'hc2adae82, 32'hc2a80ab6, 32'h41ddadcc, 32'h4290a6b9, 32'hc284a20c, 32'hc2c6aaf6, 32'hc29d87b0, 32'hc10c7b7b};
test_bias[3927:3927] = '{32'h42501ffa};
test_output[3927:3927] = '{32'h4492c8a4};
test_input[31424:31431] = '{32'hc24b9cb5, 32'hc25791cb, 32'h4242e439, 32'h424a3bb6, 32'h416e23c0, 32'h3f7d4292, 32'h413b265c, 32'hc29798ae};
test_weights[31424:31431] = '{32'hc2c732b2, 32'hc2873ce9, 32'hc1ea8c4c, 32'h3f6d7db0, 32'hc283abbb, 32'hc2105359, 32'hc229a0d1, 32'h423beb34};
test_bias[3928:3928] = '{32'h4288c0a0};
test_output[3928:3928] = '{32'h45118425};
test_input[31432:31439] = '{32'h41cc1d14, 32'hc1f9aa50, 32'h423c53b5, 32'hc27bdb67, 32'h423a043d, 32'h4209eecf, 32'hc2abed70, 32'hc28ecb66};
test_weights[31432:31439] = '{32'h40dcec4f, 32'hc29b819c, 32'hc2a6c012, 32'h4103e8fa, 32'h4297def0, 32'h42375444, 32'hc2c71c07, 32'h42c64d64};
test_bias[3929:3929] = '{32'h422f304f};
test_output[3929:3929] = '{32'h4595c54b};
test_input[31440:31447] = '{32'hc16b0314, 32'hc20bce73, 32'h426b218b, 32'h422c42f9, 32'h416e26df, 32'h4255b4ed, 32'h41d841c2, 32'hc1912cf0};
test_weights[31440:31447] = '{32'hc11c4cdc, 32'h42a2466a, 32'h41897099, 32'hc20ecc72, 32'hc235dc42, 32'hc28f9560, 32'hc29769fc, 32'h40448a47};
test_bias[3930:3930] = '{32'h42b26ee6};
test_output[3930:3930] = '{32'hc6184525};
test_input[31448:31455] = '{32'h4285b638, 32'hc288c6bb, 32'hc1e58dea, 32'h4219577c, 32'hc0ed4bf5, 32'hc125b1e3, 32'h410a8b00, 32'h424e2793};
test_weights[31448:31455] = '{32'hc2c3d5ba, 32'hc106bc85, 32'hc28e55d0, 32'hc298ad05, 32'hc0d25b96, 32'h41dff6b4, 32'h425ee68c, 32'h423b0dcf};
test_bias[3931:3931] = '{32'hc26c169d};
test_output[3931:3931] = '{32'hc58532cc};
test_input[31456:31463] = '{32'h4214853b, 32'h42b80396, 32'hc20abd8d, 32'hc2c0d75a, 32'h41c9207c, 32'hc27420e3, 32'hc137c013, 32'hc256144d};
test_weights[31456:31463] = '{32'h426c3649, 32'hc133df78, 32'hc2101e15, 32'hc2168946, 32'hc09370a7, 32'h42bf09df, 32'h41802b75, 32'h41a6ecde};
test_bias[3932:3932] = '{32'h41c709e3};
test_output[3932:3932] = '{32'hc49417c4};
test_input[31464:31471] = '{32'h41462d1e, 32'hc2633835, 32'hc2921327, 32'h42c37ed9, 32'h4258444f, 32'hc292240d, 32'h41fbffd7, 32'h42ab0ba8};
test_weights[31464:31471] = '{32'hc242db4a, 32'h418321f2, 32'hc10a19a2, 32'h424270ee, 32'hc208e90e, 32'h42823d64, 32'hc28affb5, 32'hc251cb9d};
test_bias[3933:3933] = '{32'h429facb8};
test_output[3933:3933] = '{32'hc61231aa};
test_input[31472:31479] = '{32'hc2531694, 32'h42901f09, 32'hc2c34a05, 32'h4233b06a, 32'h4260ee32, 32'h419e9c89, 32'hc26f1af2, 32'hc2343b77};
test_weights[31472:31479] = '{32'hc25d04c3, 32'hc2903262, 32'h40f42238, 32'h42ba06f9, 32'hc14246c7, 32'h4286d0f3, 32'hc2010ca2, 32'h41ceb4b4};
test_bias[3934:3934] = '{32'hc2b67c99};
test_output[3934:3934] = '{32'h451b09c8};
test_input[31480:31487] = '{32'hc2b9d709, 32'h413e621d, 32'h41e5a605, 32'hc26af2ee, 32'hc1b6a218, 32'hc210ffed, 32'h41daa290, 32'hc2ac2595};
test_weights[31480:31487] = '{32'h4204ad8e, 32'hc25216ab, 32'h428d018d, 32'hbead7348, 32'hc23ca984, 32'hc2958898, 32'h4274ba68, 32'hc2318c0a};
test_bias[3935:3935] = '{32'hc277e411};
test_output[3935:3935] = '{32'h45ec12cb};
test_input[31488:31495] = '{32'hc2bfcb3a, 32'hc2bc76f3, 32'h41bf7969, 32'h41826f0e, 32'hc17f8971, 32'h418299b5, 32'hc28781f2, 32'hc118db0c};
test_weights[31488:31495] = '{32'hc13bc7e4, 32'h426285d2, 32'h41848a55, 32'h42437fb1, 32'h4288b8dc, 32'h42bb8f3f, 32'hc2bc3444, 32'hbf6a0623};
test_bias[3936:3936] = '{32'hc2af06f8};
test_output[3936:3936] = '{32'h4568695f};
test_input[31496:31503] = '{32'hc2652778, 32'h42abc3d2, 32'h418cc2fc, 32'hc2904f3c, 32'h412cd359, 32'h42a8e1be, 32'hc2ba9767, 32'h418906ac};
test_weights[31496:31503] = '{32'h4215285d, 32'hc29697a2, 32'h42b2e598, 32'hc291ebe7, 32'h42021d9b, 32'h4101df11, 32'h41d103ac, 32'hbebdddda};
test_bias[3937:3937] = '{32'h4293b2a7};
test_output[3937:3937] = '{32'hc5419ccd};
test_input[31504:31511] = '{32'hc2b5f972, 32'hc28607f9, 32'h41bb1835, 32'hc24a65ee, 32'hc2aacb78, 32'hc27a7d26, 32'hc2a6e32b, 32'hc2917146};
test_weights[31504:31511] = '{32'hc29133ec, 32'hc1ecd66c, 32'h421a1473, 32'hc260141e, 32'hc0b8cea7, 32'h42261401, 32'hc1eb1dd6, 32'h41ea5a42};
test_bias[3938:3938] = '{32'h424c5ccb};
test_output[3938:3938] = '{32'h46257e0a};
test_input[31512:31519] = '{32'h42075b0e, 32'hc03e90d3, 32'hc20ae86f, 32'h42a2bd7d, 32'hc2003cc6, 32'hc1ac2dc5, 32'h429215eb, 32'hc089e3b3};
test_weights[31512:31519] = '{32'h4213e7ce, 32'h420a1222, 32'hc1ca1d17, 32'hc235cabf, 32'h4294142f, 32'hc23456cb, 32'hbffbc8ec, 32'hc29fae04};
test_bias[3939:3939] = '{32'h42483589};
test_output[3939:3939] = '{32'hc530937b};
test_input[31520:31527] = '{32'h42327639, 32'h4234ec28, 32'h423d5c88, 32'h42aa04ed, 32'hc2b01c2f, 32'hc1cea0e7, 32'h4260b5d6, 32'h4162289a};
test_weights[31520:31527] = '{32'hc23e67ed, 32'hc0a58c16, 32'h42170401, 32'hc2b4ce14, 32'hc2bee62d, 32'h3fccd490, 32'h414f3090, 32'h42b64266};
test_bias[3940:3940] = '{32'hc1aa76ff};
test_output[3940:3940] = '{32'h4503631f};
test_input[31528:31535] = '{32'hc21799f9, 32'hc1f9e09a, 32'h41e035ef, 32'h42b7f2ed, 32'hc2b30cd7, 32'hc22f50c1, 32'hc173a505, 32'hc1985301};
test_weights[31528:31535] = '{32'h428bcacf, 32'h42a6db20, 32'hc264353c, 32'hc283a652, 32'hc186a632, 32'h42839a33, 32'hc1c14565, 32'h4248ae7e};
test_bias[3941:3941] = '{32'h41ff4e20};
test_output[3941:3941] = '{32'hc667e2ff};
test_input[31536:31543] = '{32'hc1bc020f, 32'h41240cd4, 32'hc2875c22, 32'h425aaa13, 32'h424e685e, 32'hc2b0b635, 32'hc1d30535, 32'hc2a66885};
test_weights[31536:31543] = '{32'hc2038a62, 32'hc294fc11, 32'h418b7272, 32'h42afaf9d, 32'h42a7e57a, 32'h419decb0, 32'h41f262d4, 32'hc247ad99};
test_bias[3942:3942] = '{32'hc223d4c1};
test_output[3942:3942] = '{32'h4614f1ad};
test_input[31544:31551] = '{32'h4273d224, 32'h41d85e31, 32'hc2b7a48d, 32'hbe916d4c, 32'hc2b9608e, 32'hc2c62fc6, 32'hc23d5985, 32'h427a8a3b};
test_weights[31544:31551] = '{32'hc149738c, 32'hc1fdf617, 32'hc1df2853, 32'h42b75adc, 32'hc2aaf284, 32'hc227da16, 32'hc22f7451, 32'hc1c4098c};
test_bias[3943:3943] = '{32'h422d8593};
test_output[3943:3943] = '{32'h46541b60};
test_input[31552:31559] = '{32'h41b6e107, 32'h4281702a, 32'hc1d66ef5, 32'hc2826a67, 32'hc1a86b26, 32'h42a7712f, 32'h42c0e26f, 32'h42b9013f};
test_weights[31552:31559] = '{32'h41510e00, 32'h425098c4, 32'hc2143a22, 32'h427fce2f, 32'h4289fe22, 32'h3e95a622, 32'hc28be9e2, 32'h402068a8};
test_bias[3944:3944] = '{32'h4246eb0b};
test_output[3944:3944] = '{32'hc5e7232f};
test_input[31560:31567] = '{32'hc227cbe1, 32'hc23313d2, 32'hc28ccd15, 32'hc259ced1, 32'h42b117e2, 32'hc0c85925, 32'h427657b1, 32'h42842ca0};
test_weights[31560:31567] = '{32'hc217f327, 32'h421ddc6f, 32'h42798703, 32'h42b4867e, 32'hc21e0d4c, 32'hc0e2830b, 32'h428e78c6, 32'hc236ee7b};
test_bias[3945:3945] = '{32'h419251e7};
test_output[3945:3945] = '{32'hc6347d81};
test_input[31568:31575] = '{32'hc2793d08, 32'h4117081d, 32'h40ad8c76, 32'h4080bdfd, 32'hc2971480, 32'hc20d9469, 32'h424ae842, 32'h4196ae35};
test_weights[31568:31575] = '{32'h429ae327, 32'h421e4a44, 32'h42bbc88b, 32'h4285490c, 32'h422fec9b, 32'h418f8bac, 32'hc1df3d3d, 32'hc25ed21b};
test_bias[3946:3946] = '{32'hc0b4324d};
test_output[3946:3946] = '{32'hc61dd9a3};
test_input[31576:31583] = '{32'hbdb2d4a4, 32'h41215f1e, 32'h40ce7e88, 32'h42a70ca3, 32'hc22ee1e1, 32'h41289ecf, 32'hc2a8325a, 32'h42226d6f};
test_weights[31576:31583] = '{32'hc2b9be80, 32'h42802c00, 32'h40c28dfd, 32'hc15bdaba, 32'hc0c24a38, 32'h41e84237, 32'h42aee33b, 32'h42c39246};
test_bias[3947:3947] = '{32'h42b9bf61};
test_output[3947:3947] = '{32'hc5464d3a};
test_input[31584:31591] = '{32'h42b08a2f, 32'h41dfc8a5, 32'hc20f1f6b, 32'hc2bd916d, 32'h4251cc73, 32'hc2ab4300, 32'h4240830d, 32'hc256dae4};
test_weights[31584:31591] = '{32'hbfe13ac7, 32'h42b9ce0c, 32'h42a20e14, 32'h40cbad19, 32'h428250ec, 32'h4271cc6b, 32'h4276f32b, 32'hc24ed5ef};
test_bias[3948:3948] = '{32'hc29a7a5c};
test_output[3948:3948] = '{32'h45325a24};
test_input[31592:31599] = '{32'hc261ffc6, 32'hc2b4a0ff, 32'h412f7f6d, 32'hc2c60388, 32'hc195436a, 32'h4234377c, 32'h42ae6e1b, 32'hc14df68b};
test_weights[31592:31599] = '{32'hc1a4813c, 32'hc0d12135, 32'hc2be3bf3, 32'h422a4a59, 32'hc2ad331b, 32'h4227cfb3, 32'h429e8065, 32'h4256de97};
test_bias[3949:3949] = '{32'h42aacced};
test_output[3949:3949] = '{32'h45c50ba5};
test_input[31600:31607] = '{32'hc29fc61e, 32'hc21b8865, 32'h42c17f91, 32'h42abfc2c, 32'hc2a7fec8, 32'h428d9b66, 32'hc1de4a98, 32'hc0abc86e};
test_weights[31600:31607] = '{32'h4107607d, 32'h42c7a034, 32'hc1f182fa, 32'hc2927bb5, 32'h4219ed65, 32'h4286076c, 32'hc17e8064, 32'h429a1279};
test_bias[3950:3950] = '{32'hc27ea55e};
test_output[3950:3950] = '{32'hc6402ad4};
test_input[31608:31615] = '{32'h418b2ed0, 32'h42875003, 32'h4227544e, 32'h422a8a6c, 32'hc26baa27, 32'hc2b7c8e2, 32'hc22fafc2, 32'hc2ae5dd1};
test_weights[31608:31615] = '{32'hc28198d0, 32'h42c4d290, 32'hc2ba20ca, 32'h42adb048, 32'hc20edd11, 32'h41614368, 32'h41d87ebc, 32'hc1c5e5e9};
test_bias[3951:3951] = '{32'hc252293d};
test_output[3951:3951] = '{32'h45dcd2c6};
test_input[31616:31623] = '{32'h4240d20e, 32'h42b06091, 32'h42731ebe, 32'hc28ae041, 32'hc1abd3a5, 32'hc2c14728, 32'h427fc264, 32'h4264902c};
test_weights[31616:31623] = '{32'h42288447, 32'h41fb9456, 32'h4207f60c, 32'hc157dc4b, 32'h4213efea, 32'hc2908a92, 32'h42b02b08, 32'hc2bb3554};
test_bias[3952:3952] = '{32'hc0f950be};
test_output[3952:3952] = '{32'h465f016e};
test_input[31624:31631] = '{32'h4248afd6, 32'hc1d40392, 32'h408d1066, 32'hc217f5b4, 32'hc2a92d33, 32'hc2448c87, 32'h4295bc21, 32'hc242f4a3};
test_weights[31624:31631] = '{32'hc2ba96a3, 32'hc2c574ec, 32'hc2231568, 32'hc25f1a43, 32'h42c38fe8, 32'hc1360897, 32'hc2bde8be, 32'hc21b5843};
test_bias[3953:3953] = '{32'h42c7d64f};
test_output[3953:3953] = '{32'hc64a65ac};
test_input[31632:31639] = '{32'h41d2c568, 32'h42a8d262, 32'hc2499eb7, 32'h42872a12, 32'h42b69547, 32'h42458e0c, 32'h42878dac, 32'h4201fb9e};
test_weights[31632:31639] = '{32'h4287bc3b, 32'hc2421ce2, 32'h3fdc4ec8, 32'hc2940e53, 32'hc18ca630, 32'hc27d5e51, 32'h412ea9c9, 32'h42aaab9d};
test_bias[3954:3954] = '{32'h4246676f};
test_output[3954:3954] = '{32'hc605e36b};
test_input[31640:31647] = '{32'h4220d7c9, 32'hc2a6c67b, 32'hc22e5836, 32'hc1e4e78b, 32'hc240c94e, 32'h400d04f5, 32'hc27fc615, 32'h42a3c114};
test_weights[31640:31647] = '{32'hc23d51d1, 32'h420525c9, 32'hc2756970, 32'hc0da1d66, 32'h4200c514, 32'h40368d68, 32'hc095823d, 32'h42bd23b1};
test_bias[3955:3955] = '{32'h42a64c63};
test_output[3955:3955] = '{32'h45950ffb};
test_input[31648:31655] = '{32'h4206ae46, 32'h42649781, 32'h424705e3, 32'h411ddca0, 32'hc28635f3, 32'hc1656ff6, 32'hc1171ac4, 32'h41ea07c1};
test_weights[31648:31655] = '{32'hc257c37d, 32'h403f7d65, 32'h424a6210, 32'hc1a8d465, 32'h420a15d3, 32'h42ace835, 32'hbfa114aa, 32'h4292c0b2};
test_bias[3956:3956] = '{32'hc201d98f};
test_output[3956:3956] = '{32'hc43f9574};
test_input[31656:31663] = '{32'h42169d74, 32'h427e2711, 32'hc2427aaa, 32'h41f7edc0, 32'h426ea035, 32'hc165b0ec, 32'h421719c0, 32'h41a452f0};
test_weights[31656:31663] = '{32'h4183b5f8, 32'hc2a53b91, 32'h42651c6e, 32'hc23daf08, 32'hc2a31c6a, 32'hc2891dbd, 32'h42adb4bc, 32'hc2848d1a};
test_bias[3957:3957] = '{32'h41331f30};
test_output[3957:3957] = '{32'hc62948c2};
test_input[31664:31671] = '{32'hc2834968, 32'hc1322f27, 32'hc2af450d, 32'hc2704739, 32'h41bcf9ee, 32'hc260e5e3, 32'h429eb2db, 32'hc2a6df5e};
test_weights[31664:31671] = '{32'hc289798f, 32'hc2a378b1, 32'h41205c6f, 32'h42787ac9, 32'hc0b9a393, 32'h421e5a54, 32'h4105f50b, 32'h4261c804};
test_bias[3958:3958] = '{32'hc1d207aa};
test_output[3958:3958] = '{32'hc5afae69};
test_input[31672:31679] = '{32'h423d6326, 32'hc23590db, 32'h4262babb, 32'h42b4a58e, 32'hc2898f64, 32'h405cb3b5, 32'h423a7cb0, 32'h42856099};
test_weights[31672:31679] = '{32'h41fb29a0, 32'hc2966314, 32'h42b594a9, 32'h423e21cf, 32'hc2384a9f, 32'hc1c94095, 32'hc2833d5c, 32'hc127b424};
test_bias[3959:3959] = '{32'h40844d2f};
test_output[3959:3959] = '{32'h46558c89};
test_input[31680:31687] = '{32'hc2853110, 32'hc266f992, 32'h41a9b0bf, 32'h41d52856, 32'h4177a2d3, 32'h4241e33d, 32'hc0cf4f0b, 32'h428fb931};
test_weights[31680:31687] = '{32'hc2a645e0, 32'h41de1250, 32'hc28eb1a0, 32'h4231cf6e, 32'h42a0a257, 32'h41b55adb, 32'h4246ea21, 32'hc26328fb};
test_bias[3960:3960] = '{32'h42338de7};
test_output[3960:3960] = '{32'h44c68a17};
test_input[31688:31695] = '{32'hc292d40f, 32'hc23fc98d, 32'hc2156cfa, 32'hc299a981, 32'h412ae9b1, 32'hc2a5c875, 32'h40ad7cd1, 32'hc205af0a};
test_weights[31688:31695] = '{32'hc1b1d17b, 32'h4282695a, 32'hc0679b6c, 32'hc255516d, 32'hc23f6970, 32'hc2ac8cc7, 32'h42a5265e, 32'hc24269b7};
test_bias[3961:3961] = '{32'hc1cb001a};
test_output[3961:3961] = '{32'h4632839d};
test_input[31696:31703] = '{32'hc27e57a6, 32'hc27f75f1, 32'hc1ccb0a8, 32'h4209e112, 32'h42b5452d, 32'hc20b57c3, 32'hc1e94a60, 32'hc2089a50};
test_weights[31696:31703] = '{32'hc2abcf2d, 32'hc199a77b, 32'hbf637400, 32'hc21a30d4, 32'h4048dc86, 32'h42a24655, 32'hc281502b, 32'h41b0b376};
test_bias[3962:3962] = '{32'hc2c5151e};
test_output[3962:3962] = '{32'h457218b2};
test_input[31704:31711] = '{32'h40c50efe, 32'hc279cbfb, 32'hc14d891e, 32'h42a76490, 32'hc2b0bb67, 32'hc29fb20b, 32'hc18b5cb2, 32'h42135dfc};
test_weights[31704:31711] = '{32'h429812c8, 32'h41b2e1b6, 32'hc2a6edb1, 32'hc11f5c98, 32'hbffb837f, 32'h4222d40e, 32'hc2902805, 32'hc28433ed};
test_bias[3963:3963] = '{32'h4290e990};
test_output[3963:3963] = '{32'hc5984c46};
test_input[31712:31719] = '{32'hc2a9ff16, 32'h42018944, 32'h418cb850, 32'h42b730cb, 32'hbe7966e5, 32'hc2b413d1, 32'h429e1b60, 32'hc2810a09};
test_weights[31712:31719] = '{32'hc19d8756, 32'hc21acabe, 32'h422bdea9, 32'hc1ae006f, 32'hc286b874, 32'hc27d0a77, 32'hc292f786, 32'hc286ca13};
test_bias[3964:3964] = '{32'hc2577682};
test_output[3964:3964] = '{32'h45535a76};
test_input[31720:31727] = '{32'h41e7c1d5, 32'hc28578b5, 32'hc2182137, 32'h4279ae0c, 32'h422f9185, 32'h41b50b05, 32'h426a151f, 32'h41c3bacf};
test_weights[31720:31727] = '{32'hc25f463b, 32'h41df93c5, 32'hc1f30ed1, 32'h4252722e, 32'h413a7557, 32'hc1e1ec8f, 32'h4130d4d3, 32'h42a097ab};
test_bias[3965:3965] = '{32'hc2c0617e};
test_output[3965:3965] = '{32'h45510ee7};
test_input[31728:31735] = '{32'h428538b3, 32'hc1902837, 32'h42a988a0, 32'hc258c2df, 32'h42bfa5c5, 32'hc2a65812, 32'h423b03a9, 32'hc2905e9a};
test_weights[31728:31735] = '{32'h4286a01e, 32'h42a0200f, 32'hc2447179, 32'h41b9b47a, 32'hc154962e, 32'hc2c2f08d, 32'h42624175, 32'h426abf85};
test_bias[3966:3966] = '{32'hc2c4435b};
test_output[3966:3966] = '{32'h452cbdd4};
test_input[31736:31743] = '{32'h425c8cdf, 32'h41506691, 32'h420e954a, 32'hc2a8f16c, 32'h42c09e1f, 32'h41f4553a, 32'h41d51829, 32'hc27d92df};
test_weights[31736:31743] = '{32'hc1f40f70, 32'h4201e205, 32'hc274bd0e, 32'h4293d52a, 32'h42763bc3, 32'hc2930a66, 32'h40b878f6, 32'h4233054e};
test_bias[3967:3967] = '{32'hc2026ef1};
test_output[3967:3967] = '{32'hc6083421};
test_input[31744:31751] = '{32'h42874b7e, 32'h42b6a2f6, 32'hc280ac13, 32'hc22fcafb, 32'h4213d8b6, 32'h42c3d709, 32'hc282c1ce, 32'hc1d7776a};
test_weights[31744:31751] = '{32'h40f8d683, 32'hc2b90981, 32'h42833d95, 32'hc298f164, 32'h4232c9ad, 32'hc2c28bc1, 32'hc256120a, 32'h41f9dead};
test_bias[3968:3968] = '{32'h429fa67a};
test_output[3968:3968] = '{32'hc6597bd6};
test_input[31752:31759] = '{32'hc2919a3f, 32'h422ce17e, 32'hc0cce565, 32'h42866564, 32'h42ab6231, 32'h427193f6, 32'hc1730919, 32'hc24a6933};
test_weights[31752:31759] = '{32'hc1c10fbd, 32'hc2a6ce58, 32'h42b5b786, 32'h42532894, 32'h42a5ae27, 32'h42adcebd, 32'hc095249d, 32'hc2838c5c};
test_bias[3969:3969] = '{32'hc2b336c7};
test_output[3969:3969] = '{32'h46830d1d};
test_input[31760:31767] = '{32'hc28ad999, 32'hc2b70e51, 32'hc1b0923b, 32'hc25ee5f6, 32'hc1f8bb90, 32'h42b2e8b5, 32'h423d7c37, 32'hc1ffdbde};
test_weights[31760:31767] = '{32'h42881d35, 32'hc2a451cd, 32'hc1bec83d, 32'h418302e7, 32'h42961b88, 32'h42915e41, 32'h42b2ebdd, 32'h42a7e591};
test_bias[3970:3970] = '{32'h42b0433e};
test_output[3970:3970] = '{32'h4600696a};
test_input[31768:31775] = '{32'h42bbb43b, 32'h429a12c5, 32'hc2af8f8e, 32'h427ed69e, 32'h4231e433, 32'h41996ec3, 32'h41bb901b, 32'h4221ec0f};
test_weights[31768:31775] = '{32'hc09fd64d, 32'h422a7968, 32'hbf4a4c9d, 32'hc2a7432c, 32'hc267c55c, 32'h42ac6bcb, 32'h424f1d23, 32'hc23b2696};
test_bias[3971:3971] = '{32'h428a41de};
test_output[3971:3971] = '{32'hc578aab5};
test_input[31776:31783] = '{32'h42a81be3, 32'h418e826d, 32'h42b65738, 32'h41bc8502, 32'hc25fbd7e, 32'hc25d9964, 32'h42c1de10, 32'hc2059b76};
test_weights[31776:31783] = '{32'hc1b725a4, 32'hc2aa342b, 32'h41a4b990, 32'h42146652, 32'h42c367d2, 32'h42965569, 32'hc13774c5, 32'hc29e13a0};
test_bias[3972:3972] = '{32'hc2b59d3c};
test_output[3972:3972] = '{32'hc60ac0e2};
test_input[31784:31791] = '{32'h42289d16, 32'h40ba3c50, 32'h42472df6, 32'hc29151eb, 32'hc2b5fca9, 32'hc1026f92, 32'h414f942a, 32'hc2c0be5f};
test_weights[31784:31791] = '{32'hc2b26f1c, 32'hc2044c63, 32'hc21bdf94, 32'h419f1e1d, 32'hc24c0f7c, 32'hc27ed03c, 32'hc20bbac0, 32'hc2653d7b};
test_bias[3973:3973] = '{32'hc2265a0e};
test_output[3973:3973] = '{32'h45322c07};
test_input[31792:31799] = '{32'h422782d4, 32'h4238b82b, 32'hc25d37c6, 32'hc15a6206, 32'hc2a7c653, 32'hc19bc37b, 32'h42839796, 32'hc116c8fb};
test_weights[31792:31799] = '{32'hc2a9fc62, 32'h41564c48, 32'hc20bfa01, 32'h42ac939c, 32'h428c64b5, 32'h42aa55e9, 32'hc210b3e8, 32'hc2840214};
test_bias[3974:3974] = '{32'h3ef22ee8};
test_output[3974:3974] = '{32'hc6337f30};
test_input[31800:31807] = '{32'hc2ad9c51, 32'hc2044e88, 32'h41332bcb, 32'h417106cf, 32'hc2750915, 32'h405c0d8d, 32'hc28d6add, 32'hc23aa651};
test_weights[31800:31807] = '{32'h42a20217, 32'hc20d8b79, 32'hc2a856a7, 32'h41c96a73, 32'hc2b6a1fc, 32'hc0bca614, 32'h4282919a, 32'hc1723c96};
test_bias[3975:3975] = '{32'hbd77751a};
test_output[3975:3975] = '{32'hc594c40e};
test_input[31808:31815] = '{32'h428bb76c, 32'hc2b27f8f, 32'h41959b0c, 32'h4229de23, 32'hc266e37b, 32'h426f2e85, 32'hc29d0fb3, 32'hc2462342};
test_weights[31808:31815] = '{32'hc2b0430c, 32'h4288ac40, 32'hc1d12098, 32'hc2af0615, 32'hc1a04d9f, 32'h41fa821e, 32'h42466922, 32'h41c7f900};
test_bias[3976:3976] = '{32'h4190d62f};
test_output[3976:3976] = '{32'hc690e678};
test_input[31816:31823] = '{32'hc21381ab, 32'h41f25851, 32'hc2b6edcf, 32'hc23392ce, 32'h42162c11, 32'h42a25704, 32'hc2b625a9, 32'h428a42f1};
test_weights[31816:31823] = '{32'hc2294244, 32'h42b64020, 32'hc19bbdbe, 32'hc273e5cd, 32'hc20029f9, 32'h4221d008, 32'hc229dca9, 32'h42b671e7};
test_bias[3977:3977] = '{32'h4134214a};
test_output[3977:3977] = '{32'h46a4e10a};
test_input[31824:31831] = '{32'hc2a8fc44, 32'h41cf5a68, 32'h4269aff3, 32'h41bf4993, 32'h423f78cd, 32'hc290b2ff, 32'h42c7e86d, 32'h42adf342};
test_weights[31824:31831] = '{32'h428c80df, 32'h42bb174a, 32'hbccfd010, 32'hc12f1335, 32'h41bf76d8, 32'h422894f8, 32'h42aff441, 32'hc0ac45d0};
test_bias[3978:3978] = '{32'hc2acc22c};
test_output[3978:3978] = '{32'h4520133f};
test_input[31832:31839] = '{32'h42ac57aa, 32'hc27b6380, 32'h42a5f2fc, 32'hc278b29f, 32'hc2be9586, 32'h41e4d60d, 32'h42bbeb91, 32'h402ef99a};
test_weights[31832:31839] = '{32'hc230749f, 32'h41705541, 32'hc2c74581, 32'h42058914, 32'h42ba8271, 32'hc10fe43c, 32'h41e18f37, 32'hc234ef08};
test_bias[3979:3979] = '{32'h410a62f1};
test_output[3979:3979] = '{32'hc6a98373};
test_input[31840:31847] = '{32'h429aea1d, 32'h422fb86a, 32'hc2a8b098, 32'hc17066e1, 32'h41d621f3, 32'h403b0705, 32'h4252cea6, 32'hc26e7cd0};
test_weights[31840:31847] = '{32'h42978322, 32'hc0aee426, 32'hc1ccf257, 32'h417cf20c, 32'h4216fc5a, 32'h41b421b4, 32'hc256512f, 32'hc1d1f747};
test_bias[3980:3980] = '{32'hc2b14553};
test_output[3980:3980] = '{32'h45e37ce8};
test_input[31848:31855] = '{32'hc2a01474, 32'hc27d2b84, 32'hc1ca89a8, 32'hc2b0a63b, 32'h428081ec, 32'h412847d8, 32'hc23c6daa, 32'h4268a767};
test_weights[31848:31855] = '{32'hc256a013, 32'h423f8bd2, 32'hc2ae83f3, 32'h4283e83c, 32'hc25e5eb7, 32'hc1ccd40c, 32'hc28de008, 32'h42bfe197};
test_bias[3981:3981] = '{32'hc1b0fd0a};
test_output[3981:3981] = '{32'h452920cb};
test_input[31856:31863] = '{32'h41eb2afc, 32'h41b8f93e, 32'hc14c587d, 32'hc1942087, 32'hc1e1891c, 32'h4025e005, 32'h4244e8c0, 32'hc26a4b4b};
test_weights[31856:31863] = '{32'hc1fbf7ae, 32'hc186ba94, 32'hc254e15a, 32'hc2973a13, 32'hc2b921ef, 32'h419402ad, 32'hc280e095, 32'hc1f6df2a};
test_bias[3982:3982] = '{32'h4224ef99};
test_output[3982:3982] = '{32'h45032b1a};
test_input[31864:31871] = '{32'h4202e260, 32'h423f1f16, 32'hc1c12bd1, 32'h42aad7c0, 32'h42581627, 32'hc244e552, 32'h419a042f, 32'hc28574e2};
test_weights[31864:31871] = '{32'h42c4574d, 32'h42a25f85, 32'h4283085d, 32'hc19b950d, 32'h425a96a2, 32'h40de9b97, 32'hc28eb845, 32'hc20ac036};
test_bias[3983:3983] = '{32'h425e350c};
test_output[3983:3983] = '{32'h45e8f1a6};
test_input[31872:31879] = '{32'hc2c4824d, 32'h42791bf5, 32'h42b46840, 32'h41c80fc9, 32'hc28e2b9b, 32'hc28af1cf, 32'h422c624a, 32'hc2bfe5da};
test_weights[31872:31879] = '{32'h428f1975, 32'hc1ac05b9, 32'h4195792c, 32'h4221567f, 32'h42a725f0, 32'hc2be761e, 32'h42940730, 32'h424a59d6};
test_bias[3984:3984] = '{32'h422dd5f5};
test_output[3984:3984] = '{32'hc5cee693};
test_input[31880:31887] = '{32'h427da271, 32'h429c770d, 32'hc26c5a1f, 32'h42b661e2, 32'h42c37561, 32'h429be5c3, 32'hc2c785d4, 32'h423edfc0};
test_weights[31880:31887] = '{32'hc24aab3f, 32'h4207dfd9, 32'h4291bbe0, 32'h42b8f197, 32'hc1b3910e, 32'hc200fe44, 32'h42893b73, 32'hc11099c3};
test_bias[3985:3985] = '{32'h42725c45};
test_output[3985:3985] = '{32'hc6027de2};
test_input[31888:31895] = '{32'h428ca3a0, 32'h4242c763, 32'hc284d141, 32'hc23f3636, 32'h42075fa8, 32'hc2986ced, 32'hc270aa9b, 32'h421d2b78};
test_weights[31888:31895] = '{32'hc2369499, 32'hc2315d4a, 32'hc2974468, 32'h4249ccaf, 32'hc29f4dbe, 32'h42aa85be, 32'h4218dfa0, 32'hc2ae2b93};
test_bias[3986:3986] = '{32'hc1c1902c};
test_output[3986:3986] = '{32'hc68a41f6};
test_input[31896:31903] = '{32'h429e4818, 32'h42984106, 32'h40b30c8e, 32'h42843453, 32'h4223743a, 32'hc1d7acd7, 32'h42363da2, 32'hc28eb4cb};
test_weights[31896:31903] = '{32'h41e8ade0, 32'h429d0c82, 32'hc1b04aed, 32'hc29c368c, 32'h410383aa, 32'hc2b14f42, 32'h400ad599, 32'h428e420e};
test_bias[3987:3987] = '{32'hc2a80360};
test_output[3987:3987] = '{32'h4424b523};
test_input[31904:31911] = '{32'h4287f724, 32'h428e8313, 32'h42885ce9, 32'h41c55b75, 32'h4293e829, 32'hc25c5843, 32'h42401397, 32'hc233f351};
test_weights[31904:31911] = '{32'h425655bf, 32'hc1c37c8a, 32'hc29ecbd7, 32'h422c250a, 32'hc292319d, 32'hc1a26f3f, 32'hc287881f, 32'hc1ab9fc4};
test_bias[3988:3988] = '{32'hc1b8fe26};
test_output[3988:3988] = '{32'hc60d6644};
test_input[31912:31919] = '{32'h42c7d20d, 32'hc02fed66, 32'hc2aedd18, 32'hc196c042, 32'hc238e002, 32'hc23974ee, 32'h426d19a3, 32'hc2ae8ca7};
test_weights[31912:31919] = '{32'h4264268f, 32'hc1e4ba52, 32'hc24b3b47, 32'h4193a6c7, 32'h4269871f, 32'hc22aa905, 32'hc17dc5c3, 32'hc19d3ded};
test_bias[3989:3989] = '{32'hc289ba2d};
test_output[3989:3989] = '{32'h461a076e};
test_input[31920:31927] = '{32'h4131e583, 32'h41eae038, 32'hc240d6ae, 32'h42824e6c, 32'hc26e7a76, 32'hc2b94c09, 32'h42b7c380, 32'h42c06a3c};
test_weights[31920:31927] = '{32'h427dc9b8, 32'hc2359f02, 32'hc2598f62, 32'hc2aab4d5, 32'hc208ee24, 32'h41fd6ea7, 32'h428f8434, 32'hc2b07c51};
test_bias[3990:3990] = '{32'h41d7f789};
test_output[3990:3990] = '{32'hc5c5cfce};
test_input[31928:31935] = '{32'h40982120, 32'hc251ddaf, 32'hc14a39d1, 32'h42b5960b, 32'h423bb425, 32'h41d9585c, 32'hc27ba6fa, 32'hc25c2298};
test_weights[31928:31935] = '{32'h429a6f19, 32'hc295153e, 32'h429609a7, 32'h420f737a, 32'h407ad99c, 32'hc24592a5, 32'h429aa663, 32'h429fe538};
test_bias[3991:3991] = '{32'h4247768b};
test_output[3991:3991] = '{32'hc56cac30};
test_input[31936:31943] = '{32'h42959885, 32'hc28d5f9e, 32'hc17d10ac, 32'hc19a511b, 32'h42062dca, 32'hc234333b, 32'hc25fe42a, 32'hc2a9f7a9};
test_weights[31936:31943] = '{32'h429d2bfc, 32'hbec6bd1e, 32'h41d511c9, 32'hc1c6d4fa, 32'hc18bab4b, 32'h42c23d57, 32'h418fecec, 32'hc2359066};
test_bias[3992:3992] = '{32'h42b1f620};
test_output[3992:3992] = '{32'h45766430};
test_input[31944:31951] = '{32'h41592251, 32'hc2480037, 32'hc2acca13, 32'hc208c5f1, 32'h42164b09, 32'h42467f19, 32'h42130a38, 32'hc18fa75e};
test_weights[31944:31951] = '{32'hc151514f, 32'hc2b42fcb, 32'h4246c40e, 32'h4255bcac, 32'h41df1dc7, 32'hc29c7836, 32'hc1fb325f, 32'hc2a3c232};
test_bias[3993:3993] = '{32'h41f2cf38};
test_output[3993:3993] = '{32'hc585c88c};
test_input[31952:31959] = '{32'h41e2d083, 32'hc28f3156, 32'hc24209ca, 32'hc25c262d, 32'h41b6290d, 32'h4071d1fe, 32'h42a6795f, 32'hc1f5ca00};
test_weights[31952:31959] = '{32'hc23cda37, 32'hc28425cf, 32'hc28abef8, 32'hc2bb7153, 32'h408ae2a2, 32'hc12ea71c, 32'h4133dd4a, 32'hc2c38a6f};
test_bias[3994:3994] = '{32'h426cc4dd};
test_output[3994:3994] = '{32'h46798f59};
test_input[31960:31967] = '{32'h42a2f385, 32'h42b9d1e6, 32'h41769b53, 32'hc2b2b012, 32'h4278e195, 32'h42628bfc, 32'h42956e3a, 32'h420736ed};
test_weights[31960:31967] = '{32'hc17b2e7a, 32'h41b318eb, 32'hc2a2499e, 32'hc24f3387, 32'hc2be84c3, 32'hc26cf666, 32'hc2a44a58, 32'hc29f503a};
test_bias[3995:3995] = '{32'hc21f9ae5};
test_output[3995:3995] = '{32'hc65a5831};
test_input[31968:31975] = '{32'h41b7d3b1, 32'h428ca355, 32'hc24a4ffd, 32'hc0fb0a1e, 32'hc2c6f687, 32'hc287dea0, 32'h42009772, 32'hc2ba7028};
test_weights[31968:31975] = '{32'h42c2b2d5, 32'hc0e267ff, 32'h42b964e1, 32'h42472e16, 32'hc291a3d8, 32'hc29de82b, 32'h424473cf, 32'h425b443c};
test_bias[3996:3996] = '{32'hc2bb51db};
test_output[3996:3996] = '{32'h45b05c32};
test_input[31976:31983] = '{32'h40b08092, 32'h4251f765, 32'hc213cc79, 32'hc290d2dc, 32'hc2882a09, 32'h42b8fe1f, 32'h429f06bc, 32'hc2c68d68};
test_weights[31976:31983] = '{32'h42c3d3de, 32'h4245c82f, 32'h41fd33b7, 32'hc2b8fc41, 32'hc1decf95, 32'hc274d8c3, 32'hc1b5e2c7, 32'hbfaaa443};
test_bias[3997:3997] = '{32'hc10f6e70};
test_output[3997:3997] = '{32'h4548d8d1};
test_input[31984:31991] = '{32'h4130003d, 32'hc2254756, 32'h40f33f46, 32'h41c01497, 32'hc1c89cbe, 32'h42b7ed4f, 32'h415221fc, 32'hc266da2d};
test_weights[31984:31991] = '{32'h42a97831, 32'hc1dab351, 32'hc2138581, 32'h41c14c0e, 32'h425e3d92, 32'h42b70fbf, 32'h405aca93, 32'h429f5851};
test_bias[3998:3998] = '{32'h42a17b97};
test_output[3998:3998] = '{32'h45998975};
test_input[31992:31999] = '{32'h420107b7, 32'hc23904b7, 32'h4180c9d3, 32'h42ab3857, 32'h42bcf065, 32'h42c0f9b1, 32'hc1cf7acd, 32'hc28b2089};
test_weights[31992:31999] = '{32'hc251acc5, 32'hc0f3bdce, 32'h41aa1e5b, 32'hc1d18a5e, 32'hc2c1f020, 32'h406c3993, 32'h423f48f1, 32'h42b27a94};
test_bias[3999:3999] = '{32'hc251e8db};
test_output[3999:3999] = '{32'hc698af34};
end
`endif
