`timescale 1ns/1ns

module conv_forward_layer();

	parameter CYCLE = 2;
    parameter MULT_DELAY = 5;
	 parameter ADD_DELAY = 7;
    parameter WIDTH = 4;
	 
	 parameter NUM_TESTS 	= 10000;
	 parameter NUM_COLS 		= (WIDTH*2) +2;
	 parameter MEM_SIZE		= NUM_TESTS*NUM_COLS; 

    reg clk, reset, enable;
    reg [31:0] in_vec [WIDTH-1:0];
    reg [31:0] weight_vec [WIDTH-1:0];
	 reg [31:0] out;
    reg [31:0] mem [MEM_SIZE];
	 
	    //forever cycle the clk
    always begin
        #(CYCLE) clk = 0;
        #(CYCLE) clk = 1;
    end
	 
	conv_forward 	#(.WIDTH(WIDTH))
						conv_forward_inst(
							.clk(clk),
							.reset(reset),
							.enable(enable),
							.in_data(in_vec),
							.weights(weight_vec),
							.out_data(out)
						);
							
	 
	int i, j;
    initial begin
        reset = 0;
		  enable = 1;
		  //read the test data generated by Python into memory
		  $readmemh("/home/b/FPGA-CNN/test/test_data/conv_forward_test_data.hex", mem);
		  //for all test cases
		  for (i = 0; i < MEM_SIZE; i=i) begin
				//copy input to register
				for (j = 0; j < WIDTH; j++, i++) begin
					in_vec[j] = mem[i];
				end
				//copy weight vector to register
				for (j = 0; j < WIDTH; j++, i++) begin
					weight_vec[j] = mem[i];
				end
				//TODO: read bias term 
				
				//wait for it...
				#(CYCLE*(MULT_DELAY + ADD_DELAY*WIDTH))
				
				//check output
				assert( out == mem[i+1] );
				//increment twice to skip output val and bias_term, once to move pointer
				i = i + 3;
			end
        $display("############################################\n");
        $display("All tests passed!\n");
        $display("############################################\n");
    end

endmodule

module conv_forward #(parameter WIDTH = 8)
									(
										input logic					clk,
										input logic					reset,
										input logic					enable,
										input logic		[31:0] 	in_data 	[WIDTH-1:0],
										input logic		[31:0]	weights	[WIDTH-1:0],
										output logic	[31:0] 	out_data
									);
										
	wire connections [2*WIDTH-1] ;
	
	genvar i, j;
	generate 
		//create float_mult blocks to multiply WIDTH number 
		//of inputs with weights
		for (i = 0; i < WIDTH; i++) begin : GEN_MULTS
			wire [31:0] result;
			float_mult float_mult_inst(
												.clk_en(!reset),
												.clock(clk),
												.dataa(in_data[i]),
												.datab(weights[i]),
												.result(result)
												);
		end 
		//need input from 2 previous blocks so number of 
		//blocks in each next layer is half of previous
		for (i = WIDTH/2; i > 1; i = i/2) begin : SUM_MULTS
			wire [31:0] results [i];
			//for each block in new layer, connect to 2 prev 
			for (j = 0; j < i; j++) begin : REDUCE_SUMS
				float_add float_add_inst(
												 .aclr(!reset),
												 .clock(clk),
												 .dataa(GEN_MULTS[j].result),
												 .datab(GEN_MULTS[j+i].result),
												 .result(results[j])
												 );
			end
		end
	endgenerate
	
										
endmodule 