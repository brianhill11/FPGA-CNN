`ifndef CONV_FORWARD_TEST_H
`define CONV_FORWARD_TEST_H
reg [31:0] test_input [40000];
reg [31:0] test_weights [40000];
reg [31:0] test_bias [5000];
reg [31:0] test_output [5000];
initial begin
test_input[0:7] = '{32'h3f37dfe9, 32'h42b39c76, 32'hc2584a42, 32'h42882ccc, 32'h4299ec61, 32'hc1dcf953, 32'h42421267, 32'h429b7cf2};
test_weights[0:7] = '{32'hc13021fd, 32'h4250693c, 32'h41aa96c6, 32'h41ff7772, 32'h40abf4c8, 32'hc0c58b7f, 32'hc2167ea2, 32'hc2940472};
test_bias[0:0] = '{32'hc2acac35};
test_output[0:0] = '{32'hc4ad9ec9};
test_input[8:15] = '{32'h42712075, 32'h42c7482c, 32'h40abf39f, 32'h41e188f5, 32'hc2a82b8c, 32'hc2ac054b, 32'h41aecdb5, 32'hc0b02186};
test_weights[8:15] = '{32'h41854fb4, 32'hc292f2f3, 32'h41403a4c, 32'hbf9b2f56, 32'hc19dd782, 32'h404bc8df, 32'hc2b95004, 32'h42ae0ef8};
test_bias[1:1] = '{32'hc2129c60};
test_output[1:1] = '{32'hc5e88a1d};
test_input[16:23] = '{32'h41f047ff, 32'hc2a970d6, 32'hc24c5d5c, 32'h41c830e3, 32'h41d3590b, 32'hc299f0ae, 32'h42ac459a, 32'h41a6bfd3};
test_weights[16:23] = '{32'hc29bdb75, 32'h42c609fe, 32'hc14651bb, 32'hc1aa2aed, 32'h42c39799, 32'hc2378e09, 32'hc18c736d, 32'hc23e65d3};
test_bias[2:2] = '{32'hc2aee04f};
test_output[2:2] = '{32'hc5de05bb};
test_input[24:31] = '{32'h41dabd48, 32'hc2c1bbe6, 32'hc1d1eba6, 32'h42048f3f, 32'h42b2a752, 32'hc2a7373f, 32'h42acedf5, 32'h424974a2};
test_weights[24:31] = '{32'hc11aef4c, 32'h42acea7d, 32'hc26009b2, 32'h4250759f, 32'hc2bf996c, 32'hc2929a30, 32'h3df72912, 32'h4161a8df};
test_bias[3:3] = '{32'hc252aa78};
test_output[3:3] = '{32'hc5e11e09};
test_input[32:39] = '{32'hc28e3876, 32'h41f6d004, 32'hc2889b7e, 32'hc28b3642, 32'h42b95cd2, 32'h42a86af0, 32'hc1a5764e, 32'hc289525a};
test_weights[32:39] = '{32'h42a9e1b6, 32'hc22041f0, 32'h425c1589, 32'h413cb045, 32'hc24e7d91, 32'h42aebb59, 32'h41e7835e, 32'h42bf50a6};
test_bias[4:4] = '{32'hc27fba74};
test_output[4:4] = '{32'hc681022d};
test_input[40:47] = '{32'h41a68624, 32'h42af4f40, 32'hc12e791e, 32'hc29d79ed, 32'h423921c7, 32'hc158d8b9, 32'h42157c42, 32'h3f71b215};
test_weights[40:47] = '{32'hc290fe82, 32'hc285afbd, 32'h419d5ea5, 32'h42a9ae53, 32'h426d3a29, 32'hc23ace30, 32'hc299e4d4, 32'hc1cac0f4};
test_bias[5:5] = '{32'h42951474};
test_output[5:5] = '{32'hc656382c};
test_input[48:55] = '{32'h421631a6, 32'hc2b8bddb, 32'hc1397a06, 32'h409c0d2a, 32'hc294a47d, 32'hc1a8ca27, 32'h42769414, 32'h423c715d};
test_weights[48:55] = '{32'h41822238, 32'h42956143, 32'h42bfc9fa, 32'h4118b30f, 32'h41b0dc5d, 32'h41956e27, 32'h409c259a, 32'hc2ba7046};
test_bias[6:6] = '{32'hc2ae3b56};
test_output[6:6] = '{32'hc6540256};
test_input[56:63] = '{32'hc20e6a99, 32'h42b1d713, 32'h429432cd, 32'hc2abc17a, 32'h42c6e092, 32'h3fd38271, 32'h42889263, 32'h42653dc1};
test_weights[56:63] = '{32'h413fc333, 32'h426a1409, 32'h40ee3f12, 32'hc2732196, 32'hc247f20f, 32'hc1457816, 32'h41c0af44, 32'h42a4c658};
test_bias[7:7] = '{32'hc2aff013};
test_output[7:7] = '{32'h4638ef5a};
test_input[64:71] = '{32'hc2af6f2d, 32'hc039b4cc, 32'hc277934c, 32'h42c453dd, 32'hc2001029, 32'h42aec559, 32'hc2992a8e, 32'hc28fb832};
test_weights[64:71] = '{32'h421dda73, 32'hc2b78b99, 32'h41c2604a, 32'h40ea90fc, 32'hc0a408ad, 32'h41cd662e, 32'h41af8416, 32'hc1bb8729};
test_bias[8:8] = '{32'h42579315};
test_output[8:8] = '{32'hc4bd3683};
test_input[72:79] = '{32'h40d31ac9, 32'h4255fe69, 32'hc2814401, 32'h419985a9, 32'hc091560d, 32'h42bc5195, 32'h42a9ca7f, 32'hc29b883c};
test_weights[72:79] = '{32'hc2ba3d6b, 32'hc1bbb517, 32'h42ba4d94, 32'h42bfb755, 32'hc2ae16eb, 32'h422e06ca, 32'hc23d2cae, 32'hc2bfaf1f};
test_bias[9:9] = '{32'hc218c3a6};
test_output[9:9] = '{32'h44e62899};
test_input[80:87] = '{32'hc2604ce9, 32'h3f37ad2a, 32'hc2aee47a, 32'hc17e6e94, 32'h42526d4e, 32'h4182c45a, 32'hc29e1ba8, 32'h4196f73e};
test_weights[80:87] = '{32'hc00b87f9, 32'hc2aea105, 32'hc1c50e01, 32'hc208612a, 32'h42671c43, 32'hc0c137c9, 32'hc2c30a4d, 32'hc1703b8d};
test_bias[10:10] = '{32'h41ebcb86};
test_output[10:10] = '{32'h464d8024};
test_input[88:95] = '{32'h427e1322, 32'h42593ac6, 32'hc0ac8260, 32'h41a2b109, 32'h42899263, 32'h42a6b6f7, 32'hc25e32f0, 32'h4211b373};
test_weights[88:95] = '{32'h42b22a9a, 32'h42b2a609, 32'hc29ed8a2, 32'h426333f6, 32'h4209f5d0, 32'hc20c610b, 32'hc2be682c, 32'h3f7077aa};
test_bias[11:11] = '{32'hc2b0e499};
test_output[11:11] = '{32'h46830c0d};
test_input[96:103] = '{32'hc1865a00, 32'h421d9662, 32'h4031d8ab, 32'h412ee968, 32'hc29a8c27, 32'h408ac255, 32'h4213487e, 32'h4285c339};
test_weights[96:103] = '{32'h410b3aa4, 32'h429e2459, 32'hc130a170, 32'h4294ef15, 32'h422f7f0f, 32'h426304ee, 32'hc1c5824c, 32'hc299c088};
test_bias[12:12] = '{32'h42760074};
test_output[12:12] = '{32'hc5a82771};
test_input[104:111] = '{32'h414aa088, 32'hc226bb93, 32'hc13f8a31, 32'hc0a9d5bd, 32'hc1b8cb6e, 32'hc1d75e6e, 32'hc24dfe62, 32'h41f175ae};
test_weights[104:111] = '{32'h42ad9043, 32'h42ba9563, 32'hc255bb6f, 32'hc20ab513, 32'hc28f3ac1, 32'hc1ee7b2f, 32'h428d3f13, 32'hc257cdd4};
test_bias[13:13] = '{32'hc2690d26};
test_output[13:13] = '{32'hc597068f};
test_input[112:119] = '{32'hc220cd59, 32'h41ad378c, 32'h41bbde8e, 32'h3f8cc4b1, 32'hc19d8f17, 32'h42a6c218, 32'h4030652c, 32'hc1652012};
test_weights[112:119] = '{32'h41d0f063, 32'hc28e6dd1, 32'h4092b124, 32'h42a7575e, 32'hc22bfa40, 32'h424b4576, 32'h42781a68, 32'h41e9df06};
test_bias[14:14] = '{32'hc18488b6};
test_output[14:14] = '{32'h4517b741};
test_input[120:127] = '{32'hc2c7ab36, 32'hc259331f, 32'hc2a7c7a7, 32'h42353cb7, 32'h42833d0d, 32'h42926d47, 32'hc2bb3d01, 32'hc28ad82d};
test_weights[120:127] = '{32'hc1634f2b, 32'h41eb7e56, 32'hc2782763, 32'h4244b2bf, 32'hc166a63b, 32'h419a6aa8, 32'hc29e5ee0, 32'hc1dc578d};
test_bias[15:15] = '{32'hc1a4ddbd};
test_output[15:15] = '{32'h468500b4};
test_input[128:135] = '{32'hc1e5bece, 32'h425f1d1a, 32'hc1c0caa5, 32'h427a06bb, 32'hc2152af9, 32'hc27071a1, 32'h42a9cd7b, 32'h4184a222};
test_weights[128:135] = '{32'h428c3172, 32'h4212a375, 32'hc2bbe021, 32'h423361b5, 32'hc1dc36bc, 32'hc272a4b1, 32'hc1d79b6e, 32'hc20ecd1a};
test_bias[16:16] = '{32'hc2a59551};
test_output[16:16] = '{32'h45d4c62e};
test_input[136:143] = '{32'h41a16e21, 32'h42c77357, 32'h414a32a7, 32'h42318ea1, 32'hc0e87958, 32'h42a33fc5, 32'h41e7f619, 32'h4219187e};
test_weights[136:143] = '{32'hbd83f272, 32'hc23974b0, 32'h41339d63, 32'h428cb8fd, 32'h4198b9fc, 32'h4216462c, 32'h425ceed8, 32'h42b0663b};
test_bias[17:17] = '{32'h429c2ae6};
test_output[17:17] = '{32'h45cefac7};
test_input[144:151] = '{32'h41753263, 32'hc2968b60, 32'hc228e0f3, 32'hc2403101, 32'h42bb8f03, 32'h4227c741, 32'h41b0b4f7, 32'hc29e2931};
test_weights[144:151] = '{32'h3f4adc7c, 32'h407d0f1f, 32'hc2864e94, 32'hc02de79d, 32'hc1984cc5, 32'h42538a58, 32'h41a61895, 32'hc0ff5c13};
test_bias[18:18] = '{32'hc23063dd};
test_output[18:18] = '{32'h4581f607};
test_input[152:159] = '{32'h42b2632a, 32'h428a1ba6, 32'h42981700, 32'hc283024e, 32'hc2ab7d27, 32'h40c35c18, 32'h42aa34fc, 32'h41ab47c0};
test_weights[152:159] = '{32'hc1b94a1b, 32'h429ac289, 32'hc2a98ce8, 32'hc170762a, 32'h4274c41a, 32'h429d7ea3, 32'hc2582b52, 32'hc2c23ad9};
test_bias[19:19] = '{32'hc28fdc2e};
test_output[19:19] = '{32'hc656148a};
test_input[160:167] = '{32'h423755bd, 32'h425511e6, 32'hc2816d8f, 32'hbdbdffda, 32'h42ae35da, 32'h3ff139b8, 32'h428b8553, 32'h42aaff56};
test_weights[160:167] = '{32'hc2303125, 32'h42b1400d, 32'hc11e6e83, 32'h4298a494, 32'hc1de7ed7, 32'h4247826d, 32'h4285cec4, 32'hc2b7a8c3};
test_bias[20:20] = '{32'h4222f2ec};
test_output[20:20] = '{32'hc50583c4};
test_input[168:175] = '{32'h4091f361, 32'hc20ec974, 32'hc2b930b9, 32'h40645590, 32'h4266ff26, 32'hc10181d0, 32'h422610f8, 32'h419a6e78};
test_weights[168:175] = '{32'h40ab4c65, 32'h418128fe, 32'h4215d5b5, 32'h413e173e, 32'hc16f1a86, 32'h420f5f07, 32'h41bbcc8d, 32'h4200a303};
test_bias[21:21] = '{32'hbf9f57db};
test_output[21:21] = '{32'hc55d0fc8};
test_input[176:183] = '{32'h41f420ff, 32'hc0949906, 32'h3ecfe94f, 32'hc1cf8bf3, 32'h42bc4e5d, 32'hc2886478, 32'hc0e1f8cf, 32'hc260181e};
test_weights[176:183] = '{32'h41813716, 32'hc2630abe, 32'hc1a37e68, 32'hc06f7122, 32'hc28abe8b, 32'h4194d8cb, 32'hc281f0fd, 32'h42978c85};
test_bias[22:22] = '{32'hc223151b};
test_output[22:22] = '{32'hc628795f};
test_input[184:191] = '{32'h429787dc, 32'h42c6e00a, 32'h419dc9c1, 32'hc2a0c1d6, 32'h429255f7, 32'h4177ce3c, 32'h4287eab3, 32'h41e4058a};
test_weights[184:191] = '{32'hc190b092, 32'hc2b962c4, 32'h42244794, 32'hc2044abd, 32'hbf8d75f7, 32'h419b15cd, 32'h42784116, 32'hc288537a};
test_bias[23:23] = '{32'h415a5875};
test_output[23:23] = '{32'hc5901906};
test_input[192:199] = '{32'hc2149f3c, 32'hc133868a, 32'hc216974f, 32'hc261b8b0, 32'hc28e9472, 32'hc17c8ceb, 32'h4290a157, 32'hc22111d2};
test_weights[192:199] = '{32'hc1736c72, 32'hc2c76258, 32'hc281e634, 32'h422d0db3, 32'h412ef419, 32'h42b8a740, 32'h42518790, 32'h42a01b98};
test_bias[24:24] = '{32'h40f09e5f};
test_output[24:24] = '{32'h41b6cbbc};
test_input[200:207] = '{32'hc28d3ca8, 32'h4283e63c, 32'hc273bb2c, 32'hc219f65f, 32'h41bc9648, 32'hc2af9624, 32'h42965480, 32'hc21772c9};
test_weights[200:207] = '{32'h428345e0, 32'h429adc3b, 32'h427e3a23, 32'h40ec3e1d, 32'h42408fe5, 32'h42bf7781, 32'hc114f7b0, 32'h42b75d11};
test_bias[25:25] = '{32'hc2a7fc67};
test_output[25:25] = '{32'hc66da9fc};
test_input[208:215] = '{32'h417fcc7e, 32'hc282a72a, 32'h4283c046, 32'hc27955e9, 32'h41d53a5f, 32'h4224e699, 32'h429af453, 32'h41b6eb98};
test_weights[208:215] = '{32'hc1e8430e, 32'h42489c78, 32'hc27bf359, 32'hc160a2fc, 32'h428460b2, 32'hc21a4a8e, 32'h4145c8ae, 32'hc20d82a5};
test_bias[26:26] = '{32'h417ef7fa};
test_output[26:26] = '{32'hc5d09f38};
test_input[216:223] = '{32'h429ccc36, 32'h4221b71b, 32'hc1c4ee24, 32'hc28e1e65, 32'hc2406214, 32'h402d76dd, 32'h41c5a3d4, 32'h42c7fdb3};
test_weights[216:223] = '{32'h4110d388, 32'hc24cb602, 32'hc2aed141, 32'hc22209be, 32'hc29f0b16, 32'hc224b33d, 32'h4224d0fd, 32'hc22420b4};
test_bias[27:27] = '{32'hc13665c5};
test_output[27:27] = '{32'h4585fb79};
test_input[224:231] = '{32'hc2b64d43, 32'hc1a2b29a, 32'hc1aac4b8, 32'hc2c37c11, 32'h41b709b8, 32'h41e5be2f, 32'hc1698bb5, 32'hbdaeb726};
test_weights[224:231] = '{32'hc2444721, 32'h41a7de36, 32'h41852696, 32'hc2132621, 32'hc1bfdcee, 32'hc26ebfb6, 32'h4203820e, 32'h429e0a04};
test_bias[28:28] = '{32'hc2129c2d};
test_output[28:28] = '{32'h458ca22b};
test_input[232:239] = '{32'hc2990ac1, 32'hc2bb4aa6, 32'hc2c13d1d, 32'hc1c09abf, 32'hc2affc3d, 32'hbf5a193e, 32'hc01047a9, 32'h42166a80};
test_weights[232:239] = '{32'hc1a60083, 32'hc205da73, 32'hc2972c90, 32'h41e587d4, 32'h4233615c, 32'hc18a8636, 32'hc2242b70, 32'h410be833};
test_bias[29:29] = '{32'h4289a9c6};
test_output[29:29] = '{32'h45f6a6a2};
test_input[240:247] = '{32'h418d02f5, 32'h42497c6d, 32'hc198a151, 32'hc05778cd, 32'h4290c178, 32'hc2b17fbc, 32'hc2a04e7a, 32'hc11baaa5};
test_weights[240:247] = '{32'hc210fe92, 32'h42a100d6, 32'hc29fffdc, 32'hc1e481a5, 32'hc29f31d9, 32'h42207a54, 32'h407880f4, 32'hc289aa68};
test_bias[30:30] = '{32'hc2b20705};
test_output[30:30] = '{32'hc57adb47};
test_input[248:255] = '{32'hc19c3ceb, 32'h426fcfaf, 32'h41e0b3e5, 32'h423d32b0, 32'h409c6d41, 32'h41cec464, 32'hc2499235, 32'h42ac2e5e};
test_weights[248:255] = '{32'hbec84be5, 32'hc29071a0, 32'h42898213, 32'h4187129f, 32'hc227d9f4, 32'hc21b00f6, 32'hc2c0f4b1, 32'h41c5ca79};
test_bias[31:31] = '{32'h428320a8};
test_output[31:31] = '{32'h45850545};
test_input[256:263] = '{32'h42c365d7, 32'h42b0eb69, 32'h419ef684, 32'hc2941921, 32'h4255b1da, 32'h41e465eb, 32'hc1d77d66, 32'h425c659a};
test_weights[256:263] = '{32'h41fc1f6b, 32'h4085e07e, 32'h417b2484, 32'hc186d013, 32'hc2c6de32, 32'hc25597ec, 32'h42ae82e8, 32'hc2a6f8e5};
test_bias[32:32] = '{32'h416a91a9};
test_output[32:32] = '{32'hc608ee00};
test_input[264:271] = '{32'hc20b2241, 32'h414fb297, 32'hc275d483, 32'h426c19fa, 32'h427cf77d, 32'h4215e244, 32'hc08027ba, 32'h409692ed};
test_weights[264:271] = '{32'hc12c6785, 32'h4245eda2, 32'hc1ae3999, 32'h41bf46d7, 32'h422b3939, 32'hc2c402ca, 32'hc2bdaa32, 32'hc28bce99};
test_bias[33:33] = '{32'hc231eb7b};
test_output[33:33] = '{32'h452f7f9c};
test_input[272:279] = '{32'h42810fb1, 32'hc28848d6, 32'hc201c6a8, 32'h420c1c05, 32'hc1f9106c, 32'hc2a1f339, 32'h429e12e4, 32'h424d35c9};
test_weights[272:279] = '{32'h42a24bd8, 32'h40c21aa9, 32'h41c795f4, 32'hc28f66b7, 32'hc1f9817e, 32'h41cfb5d4, 32'h4284e85c, 32'h42368b3b};
test_bias[34:34] = '{32'h418ea0bb};
test_output[34:34] = '{32'h45f971f0};
test_input[280:287] = '{32'h3f190494, 32'hc1940709, 32'h4207198c, 32'h42978fe8, 32'hc29d4209, 32'hc2b81ea5, 32'h429e7fbd, 32'hc1bf9dff};
test_weights[280:287] = '{32'h425cde09, 32'h4216ecfe, 32'h42098398, 32'h4236a1f0, 32'h4290b9b0, 32'h427b2717, 32'hc2c791de, 32'hc1d833dc};
test_bias[35:35] = '{32'hc2626dfc};
test_output[35:35] = '{32'hc667bd13};
test_input[288:295] = '{32'hc2505a3c, 32'h42a2c7e8, 32'h41e912ab, 32'h427cd62d, 32'hc180b994, 32'h42713899, 32'hc2ad990c, 32'h42b9fc8c};
test_weights[288:295] = '{32'h42297ce7, 32'hc2371978, 32'hc0736ea4, 32'h426b9049, 32'h42a8b84e, 32'h427eb873, 32'hc296fa05, 32'h42830c6a};
test_bias[36:36] = '{32'hc2a4affa};
test_output[36:36] = '{32'h4646d422};
test_input[296:303] = '{32'hc23ac27c, 32'hc28e01c2, 32'h42c23c73, 32'h42a33ca0, 32'hc29a133d, 32'h42c7e90e, 32'h421f4799, 32'hc216576e};
test_weights[296:303] = '{32'hc1a5bbad, 32'h4065c655, 32'hc2a1d702, 32'hc2c26ed4, 32'h4262a0dd, 32'h42b06dfb, 32'hc1c5a30a, 32'hc28cc4bf};
test_bias[37:37] = '{32'h42a97075};
test_output[37:37] = '{32'hc60ac795};
test_input[304:311] = '{32'hc201a4b8, 32'hc29ae1aa, 32'hc0695a44, 32'h41864beb, 32'h426e79ee, 32'hc22775e4, 32'h428a9b91, 32'hc2281bab};
test_weights[304:311] = '{32'h41ecf63b, 32'hc29c65b4, 32'h4259f34b, 32'h42b74f53, 32'hc242ff65, 32'h4208325c, 32'hc2bb1732, 32'h4190960f};
test_bias[38:38] = '{32'h420fc82f};
test_output[38:38] = '{32'hc59f76c1};
test_input[312:319] = '{32'hc1f790eb, 32'h41713b6a, 32'h41800230, 32'hc294bb55, 32'hc18505c6, 32'hc2344ff2, 32'hc10c705b, 32'hbfba498b};
test_weights[312:319] = '{32'hc28a042c, 32'h423d2695, 32'hc2c7487b, 32'h42737862, 32'hc259416f, 32'h4206d953, 32'h42971652, 32'hc25639d8};
test_bias[39:39] = '{32'h4287b2b9};
test_output[39:39] = '{32'hc589b1c5};
test_input[320:327] = '{32'hc10c5a5d, 32'h414922d5, 32'h41c57d6f, 32'hc00955d7, 32'h42a6ed86, 32'h422bad23, 32'h414736a3, 32'hc28b9fca};
test_weights[320:327] = '{32'h418e0438, 32'h4157e90d, 32'hc2a96059, 32'h42abab71, 32'h41329748, 32'h42081c21, 32'h4218323c, 32'h42bfd8ac};
test_bias[40:40] = '{32'h42933837};
test_output[40:40] = '{32'hc5bc10da};
test_input[328:335] = '{32'hc1b3709a, 32'hc19fa618, 32'hc2a361c5, 32'hc23b1d60, 32'hc2c1e478, 32'h422face0, 32'hc26f7775, 32'h4049b90c};
test_weights[328:335] = '{32'hc0a4b429, 32'h402efa4e, 32'h428dbf1c, 32'hc2351afb, 32'hc292b0aa, 32'h41a2e7d3, 32'h41beab4b, 32'hc1e267f7};
test_bias[41:41] = '{32'h41da6049};
test_output[41:41] = '{32'h45359422};
test_input[336:343] = '{32'h417fe8a3, 32'h42ae5aa8, 32'h42376ec9, 32'h41a8f2b7, 32'hbba1d646, 32'hc2adf6a5, 32'hc24d521a, 32'hc2c5aafc};
test_weights[336:343] = '{32'hc2bee9c6, 32'hc26afea5, 32'h42112728, 32'hc20ed8e1, 32'hc29efda8, 32'hc286b09a, 32'h42bfa4f8, 32'hc2c28c0c};
test_bias[42:42] = '{32'h422bbce9};
test_output[42:42] = '{32'h4597d0c5};
test_input[344:351] = '{32'h42521db0, 32'h425c510d, 32'h42314cce, 32'hc24b4289, 32'hc2490304, 32'h42c5cf68, 32'h420514da, 32'hc12f6177};
test_weights[344:351] = '{32'h42a7ab77, 32'hc20141fa, 32'h416d6bd1, 32'hc291c63d, 32'hc1d65ba0, 32'hc2973f13, 32'hc290f9c3, 32'hc1494003};
test_bias[43:43] = '{32'hc1c65d8a};
test_output[43:43] = '{32'hc4b4c70e};
test_input[352:359] = '{32'h41be7a80, 32'hc2193cbc, 32'hc1ed6c73, 32'h429b6dc5, 32'hc0e29644, 32'h4118b836, 32'h422d8f7b, 32'hc2817b96};
test_weights[352:359] = '{32'h42ac8829, 32'h417404bd, 32'h421be029, 32'h42829a71, 32'h42a545ae, 32'hc2b8b6ca, 32'hc2913360, 32'hc2ab1731};
test_bias[44:44] = '{32'hbeab8080};
test_output[44:44] = '{32'h45c529f6};
test_input[360:367] = '{32'h40b79fd3, 32'h42a9728f, 32'h40bbdd14, 32'h420a8751, 32'h41b31357, 32'h4283b433, 32'hc1e82090, 32'hc02f4044};
test_weights[360:367] = '{32'h42aa8f4a, 32'h429e4739, 32'hc26ee055, 32'h41edc35b, 32'h4197b3b5, 32'hc2830dde, 32'h42be2eb4, 32'h40b398a6};
test_bias[45:45] = '{32'hc28e907a};
test_output[45:45] = '{32'h448e129a};
test_input[368:375] = '{32'h42b9d32c, 32'h41667d52, 32'hc19f6b50, 32'h42b47de5, 32'h4246e218, 32'hc24b0caf, 32'hc29f595d, 32'hc2444dd2};
test_weights[368:375] = '{32'h41ac2e30, 32'h41a5226f, 32'hc2c41c2a, 32'h42694f22, 32'hc2a40a89, 32'h4248d591, 32'hc0cdfc08, 32'hc1d4b874};
test_bias[46:46] = '{32'h41d9dc00};
test_output[46:46] = '{32'h4593e860};
test_input[376:383] = '{32'hc2752127, 32'h4185a38d, 32'hc1dfeee5, 32'hc122a04a, 32'hc1ddcc21, 32'h4239b72d, 32'h41587b9b, 32'h411ed9bf};
test_weights[376:383] = '{32'hc22e1fa3, 32'hc20478a8, 32'h42834fd2, 32'hc1176801, 32'h41981024, 32'h423169bf, 32'h42bde3b5, 32'hc29d7d4b};
test_bias[47:47] = '{32'h41cabbee};
test_output[47:47] = '{32'h4518144f};
test_input[384:391] = '{32'hc26bcddf, 32'hc239aa16, 32'hc205f63f, 32'hc29e90f4, 32'h42a779d4, 32'h42845e5c, 32'hc235a70d, 32'h42a09ad4};
test_weights[384:391] = '{32'h4220b6be, 32'hc2894bb9, 32'h42a192ad, 32'hc09324ce, 32'h429f3fad, 32'hc1ab6e77, 32'hc246056f, 32'h4263b98b};
test_bias[48:48] = '{32'hc2794ee9};
test_output[48:48] = '{32'h4623cec1};
test_input[392:399] = '{32'h426b3b13, 32'hc151e4d3, 32'h42245496, 32'h4217d7a9, 32'hc0a0495a, 32'hc289a265, 32'h4108906a, 32'hc23e087d};
test_weights[392:399] = '{32'h413f2bda, 32'hc180fa7e, 32'h405ff0a3, 32'hc131737c, 32'h4292de8f, 32'hc22f719d, 32'hc299f314, 32'h421bc790};
test_bias[49:49] = '{32'hc27ddd23};
test_output[49:49] = '{32'h4433315b};
test_input[400:407] = '{32'h428deba3, 32'hc219042b, 32'hc1dd9a09, 32'h42b014e1, 32'h42c0b0cf, 32'hc2183540, 32'hc2305ee3, 32'h429cfae5};
test_weights[400:407] = '{32'hc200392e, 32'h418a1a02, 32'hc1e298e0, 32'hc29ddcaa, 32'hc2c1c536, 32'h41ba2f88, 32'h42a74060, 32'hc2863e4d};
test_bias[50:50] = '{32'hc02f24f4};
test_output[50:50] = '{32'hc6dcec10};
test_input[408:415] = '{32'hc282456a, 32'hc29e6804, 32'hc15bf4cb, 32'h42435460, 32'hc1479414, 32'hc294468f, 32'hc2a42d67, 32'hc2272436};
test_weights[408:415] = '{32'h42620948, 32'h42b6e402, 32'hc1ea6186, 32'hc2b18377, 32'h42a7a566, 32'h42abda4d, 32'h42a3e5e0, 32'h42acecfd};
test_bias[51:51] = '{32'hc24a8eb2};
test_output[51:51] = '{32'hc6ff2b0f};
test_input[416:423] = '{32'hc2519b77, 32'hc08747a2, 32'hc2902bec, 32'h42b5bca9, 32'hc127f18d, 32'h428cec0a, 32'h422a6ed2, 32'hc15e764a};
test_weights[416:423] = '{32'h42b789b1, 32'hc271b320, 32'hc2a0b65f, 32'h42005872, 32'h428fbabf, 32'h4247285f, 32'h4291a8de, 32'h427ab692};
test_bias[52:52] = '{32'h428c3b21};
test_output[52:52] = '{32'h460fe9c9};
test_input[424:431] = '{32'hc19dbc28, 32'h422a784d, 32'hc1f4467e, 32'hc1cb7fc6, 32'h41c5691e, 32'h42426c62, 32'hc198e5c2, 32'h42a1f8b8};
test_weights[424:431] = '{32'hc2aad61b, 32'h41a13ed3, 32'h42b5b7f9, 32'h42a8bec7, 32'hc20a16ea, 32'h41251725, 32'hc280f1b2, 32'hc2a48ca4};
test_bias[53:53] = '{32'h4105d84d};
test_output[53:53] = '{32'hc5feb225};
test_input[432:439] = '{32'h428e025c, 32'h423c8eef, 32'hc2056f52, 32'h423d8ff5, 32'h4262bc6a, 32'hc2166f11, 32'hc2b42a39, 32'h42299b3b};
test_weights[432:439] = '{32'hc2b7091e, 32'hc22bf1d6, 32'hc24501c2, 32'h4284e18f, 32'hc28ed455, 32'hc24464f1, 32'h42c3c1f1, 32'h42a19abf};
test_bias[54:54] = '{32'hc1f61541};
test_output[54:54] = '{32'hc63170f1};
test_input[440:447] = '{32'h4165c6b9, 32'hc2134d9d, 32'hc21c656f, 32'h429fab4d, 32'hc23e3754, 32'h42b10aac, 32'h418dcb3c, 32'h40a6226c};
test_weights[440:447] = '{32'h4287676c, 32'hc1715955, 32'h428fb018, 32'h417970d9, 32'hc24555b7, 32'hc256f0ce, 32'hc248f09f, 32'hc2a8bf47};
test_bias[55:55] = '{32'hc149dfda};
test_output[55:55] = '{32'hc56cc585};
test_input[448:455] = '{32'hc2a69ddc, 32'h422349fb, 32'hc206f77b, 32'hc2b35676, 32'hc1555068, 32'hc2b4c050, 32'hc2b94f5f, 32'h421ca267};
test_weights[448:455] = '{32'hc22c19a2, 32'hc21d34aa, 32'h4292049d, 32'hc241c344, 32'hc023f2b7, 32'hc0c1de88, 32'hc1d9857c, 32'h42b439c6};
test_bias[56:56] = '{32'hc08bba08};
test_output[56:56] = '{32'h4623d5db};
test_input[456:463] = '{32'hc1f5f99e, 32'hc2ab4df1, 32'hc11dcf00, 32'hc23b6207, 32'hc16d9016, 32'hc19abed5, 32'h4234c19d, 32'h41cecbc8};
test_weights[456:463] = '{32'h429f79f1, 32'hc29d06d1, 32'hc259d626, 32'hc28d2e57, 32'h428c0546, 32'h4283f65a, 32'h41fa5f51, 32'hc282ef6f};
test_bias[57:57] = '{32'hc04d6631};
test_output[57:57] = '{32'h45ac80dc};
test_input[464:471] = '{32'hc275f280, 32'hc21c2639, 32'hc1a10ac0, 32'hc24f53a3, 32'hc20345f5, 32'h40e29064, 32'h42a42b02, 32'hc1dcf9d6};
test_weights[464:471] = '{32'hc0dd61c4, 32'h41a7485e, 32'h428ef38b, 32'h42457528, 32'h42b5fdb7, 32'hc265e464, 32'hc2c549ce, 32'hc29c3fa9};
test_bias[58:58] = '{32'hc12c4037};
test_output[58:58] = '{32'hc6568e1e};
test_input[472:479] = '{32'h428b7ad0, 32'hc28c57fd, 32'h42218ef7, 32'h4230a927, 32'h41c10e72, 32'h429b6471, 32'h42c3312f, 32'hc246f350};
test_weights[472:479] = '{32'hc29a1d8c, 32'h42309c5a, 32'hc276379a, 32'hc265e82d, 32'hc2945dec, 32'hc28e5440, 32'hc0d1c15f, 32'hc2922dfb};
test_bias[59:59] = '{32'hc25aba7a};
test_output[59:59] = '{32'hc68ba6cf};
test_input[480:487] = '{32'hc206d336, 32'hc2134551, 32'h426ce68b, 32'h41f420f5, 32'h42b5cee2, 32'hc211b7e5, 32'h427d5d83, 32'h4185b432};
test_weights[480:487] = '{32'h424d734d, 32'h41de073a, 32'h42a3ad13, 32'h42316785, 32'h417919e0, 32'hc1a1b4d3, 32'h415f7dff, 32'h42bd38fa};
test_bias[60:60] = '{32'h427d784e};
test_output[60:60] = '{32'h45fe01dc};
test_input[488:495] = '{32'hc1fab2dd, 32'h4297fb79, 32'hc2c40ac8, 32'hc295dbc0, 32'h414fb7e0, 32'h425cea3e, 32'hc230e956, 32'h420b02e5};
test_weights[488:495] = '{32'hc272eab9, 32'hc22b35a7, 32'h428ddf82, 32'h42c5387c, 32'hc158d45a, 32'h42b59c52, 32'h428a0727, 32'h41f2989c};
test_bias[61:61] = '{32'h4101aeb8};
test_output[61:61] = '{32'hc648ab4b};
test_input[496:503] = '{32'h422bc725, 32'hc102f62b, 32'hc29950bb, 32'hc29b6b12, 32'h4281c819, 32'hc2369d90, 32'hc28568f7, 32'hc0c796e6};
test_weights[496:503] = '{32'h42b0c8fc, 32'hc2a492b6, 32'h42a155fa, 32'h4168d805, 32'h42a2a2f9, 32'h4287ddcb, 32'hc1af98fa, 32'h425a53ca};
test_bias[62:62] = '{32'h42ba94aa};
test_output[62:62] = '{32'h4408cd3a};
test_input[504:511] = '{32'hc11159cf, 32'hc0c65750, 32'h42bce477, 32'hc2b89600, 32'hc294d25f, 32'h42952493, 32'hc248673f, 32'h42762d39};
test_weights[504:511] = '{32'h42be4abe, 32'h426c0fb5, 32'h421cc915, 32'hc2901347, 32'hc22b124f, 32'h42b6e429, 32'h4154dc27, 32'hc222d0a1};
test_bias[63:63] = '{32'h42b92e1b};
test_output[63:63] = '{32'h467aabfb};
test_input[512:519] = '{32'hc2c40ba9, 32'h429c72b0, 32'hc262a7d7, 32'h4285af44, 32'h417f55e3, 32'h411f24b1, 32'hc2811928, 32'h4202c841};
test_weights[512:519] = '{32'hc2821bfd, 32'hc0bb4274, 32'hc289c5b7, 32'hc2b85276, 32'hc1d4557a, 32'hc2923397, 32'h42b2b681, 32'hc2b5dbef};
test_bias[64:64] = '{32'h41668058};
test_output[64:64] = '{32'hc5c2378d};
test_input[520:527] = '{32'h42600355, 32'h42ba37d3, 32'hbecd51b4, 32'hc27d6c71, 32'h42060265, 32'hc286259c, 32'h428f57dd, 32'hc2b8f2cc};
test_weights[520:527] = '{32'hc0ed50c2, 32'h42aa8785, 32'h42285a83, 32'hc25f2218, 32'hc028c4c1, 32'hbf16b28c, 32'h42c5a453, 32'hc1de1dcb};
test_bias[65:65] = '{32'hc252b9ee};
test_output[65:65] = '{32'h46a0db0e};
test_input[528:535] = '{32'h41886277, 32'hc1296568, 32'hc1d3546c, 32'hc1be6bd1, 32'hc25ef30a, 32'hc284be3a, 32'hc2297089, 32'hc14d8054};
test_weights[528:535] = '{32'hc0e77925, 32'hc2a62483, 32'h42949b62, 32'h41779599, 32'hc266545a, 32'h41e8cfc8, 32'hc2136ab8, 32'hc284fc75};
test_bias[66:66] = '{32'hc2b2b952};
test_output[66:66] = '{32'h44fd9a64};
test_input[536:543] = '{32'h4239777b, 32'hc2b0854c, 32'h42c4c983, 32'h42acea13, 32'h420bffb3, 32'h4051439d, 32'h422afc81, 32'hc288e79e};
test_weights[536:543] = '{32'hc20ee10c, 32'h423576cd, 32'h42ac1eac, 32'hc17e249f, 32'hc2a75eda, 32'hc2862645, 32'h42349a95, 32'hc0c2ee74};
test_bias[67:67] = '{32'h429ae3f6};
test_output[67:67] = '{32'h44319be0};
test_input[544:551] = '{32'hc2506e6e, 32'h428b612b, 32'hc1684642, 32'hc2b0a186, 32'h42bb1cec, 32'hc2aed11f, 32'h41c30461, 32'h42184e2d};
test_weights[544:551] = '{32'h42a46f2b, 32'h4295a207, 32'h41d02da5, 32'hc21704dc, 32'h40b81587, 32'hc231b55f, 32'hc293e5a2, 32'hc29de573};
test_bias[68:68] = '{32'hc13b8718};
test_output[68:68] = '{32'h4559f6a5};
test_input[552:559] = '{32'hc28ed442, 32'h4226a75c, 32'h421090af, 32'hc2af039a, 32'h42add2d7, 32'h426fdae3, 32'hc29c6bf9, 32'hc17e5183};
test_weights[552:559] = '{32'hbec0bc06, 32'hc212cdce, 32'h42479f3f, 32'h4220a2af, 32'h42b37583, 32'h40e2cfca, 32'h42189898, 32'h42026bae};
test_bias[69:69] = '{32'hc2a66bfb};
test_output[69:69] = '{32'h44b2362d};
test_input[560:567] = '{32'h4278c751, 32'h4290b18d, 32'hc1b70f8d, 32'h42965c2b, 32'hc2955ed1, 32'hbee6c4e7, 32'h415b75e1, 32'h42176f9d};
test_weights[560:567] = '{32'hc211a746, 32'hc2938c2f, 32'hc249fd1d, 32'h42bc56f4, 32'h41d912ec, 32'h42ac15e2, 32'hc1949371, 32'h419ba4ec};
test_bias[70:70] = '{32'h428bb46e};
test_output[70:70] = '{32'hc45c1c56};
test_input[568:575] = '{32'hc2badaaa, 32'h415e8cdf, 32'hc12edb55, 32'hc2418dc0, 32'h417d3ab1, 32'h42946363, 32'h429ae47a, 32'hc18cde01};
test_weights[568:575] = '{32'hc2bbe832, 32'h42bcfb4c, 32'h41f52a64, 32'hc288f3a9, 32'hc1f5f074, 32'hc2480f9b, 32'hc2225610, 32'hc256abd3};
test_bias[71:71] = '{32'h429d4bff};
test_output[71:71] = '{32'h45d30e8d};
test_input[576:583] = '{32'hc283b592, 32'hc1a232b0, 32'h42582030, 32'hc2aeba9d, 32'hc2113b12, 32'hc2882370, 32'h42853244, 32'h42959288};
test_weights[576:583] = '{32'h4249ceb9, 32'h40fb8bb4, 32'h42c40f9a, 32'h41a3311a, 32'h4286a7a5, 32'h42828533, 32'hc1503d6a, 32'h40da8c4c};
test_bias[72:72] = '{32'h421ca300};
test_output[72:72] = '{32'hc5e016ca};
test_input[584:591] = '{32'h4272eea0, 32'h41dd850c, 32'hc1e72550, 32'hc284cb92, 32'hc2b2f8b2, 32'h41ec8b8d, 32'hc2628a8f, 32'hc298b195};
test_weights[584:591] = '{32'hc23c4e9b, 32'h42b0d1db, 32'hc2017ae8, 32'hc2b43543, 32'h3fa7cc40, 32'hbf9cd313, 32'hc2370e81, 32'hc1e43ff4};
test_bias[73:73] = '{32'hc2c4415c};
test_output[73:73] = '{32'h462c4590};
test_input[592:599] = '{32'h421e3b8c, 32'hc19c1916, 32'h42189841, 32'hc120e752, 32'h41011664, 32'hc21da6bd, 32'hc0909c1e, 32'h41c2b242};
test_weights[592:599] = '{32'h42a9c1b5, 32'hc2a19d78, 32'h426403b0, 32'h427f12f2, 32'hc1b74c35, 32'h427dbaba, 32'h42b5136c, 32'hc2a4c221};
test_bias[74:74] = '{32'hc206f191};
test_output[74:74] = '{32'h44a6e162};
test_input[600:607] = '{32'h42a25fdc, 32'h42924c6f, 32'h4267d782, 32'hc0ec1857, 32'h413d508a, 32'hc29485d7, 32'hc27b779f, 32'hc28ea175};
test_weights[600:607] = '{32'hc1aa65bc, 32'hc25e9456, 32'h427c8efc, 32'h4262489d, 32'h41ba5e99, 32'hc15ecb45, 32'h420b3ce1, 32'h4230bbac};
test_bias[75:75] = '{32'hc1b75481};
test_output[75:75] = '{32'hc5ce8f79};
test_input[608:615] = '{32'hc2b083fe, 32'hc29ad884, 32'hc2528c22, 32'h4135c5db, 32'hc286dfcd, 32'h41980c76, 32'hc2c1b852, 32'h429afcf2};
test_weights[608:615] = '{32'h42005980, 32'hc0fe0c7b, 32'hc299ca07, 32'hc2950b52, 32'hc29b8319, 32'h423d89ee, 32'hc2b8cf0c, 32'hc21593cd};
test_bias[76:76] = '{32'h429d04d7};
test_output[76:76] = '{32'h464f2b07};
test_input[616:623] = '{32'hc1538dde, 32'hc1220fe9, 32'h41a1b594, 32'hc2ba05d8, 32'h42534d09, 32'hc1871e51, 32'hc2b2c972, 32'h41f92822};
test_weights[616:623] = '{32'h428a9901, 32'h4256b72f, 32'h411f44c0, 32'hc29b39a0, 32'h41c90b9f, 32'h416aa8dd, 32'h42b0d073, 32'hc2a4838e};
test_bias[77:77] = '{32'hc17156a9};
test_output[77:77] = '{32'hc55700eb};
test_input[624:631] = '{32'h423bc89e, 32'hc259e49e, 32'h41b7f42e, 32'hc26f6c9e, 32'h420e146f, 32'hc2922fe1, 32'hc26bfab6, 32'hc19f285c};
test_weights[624:631] = '{32'hc22d278d, 32'hc2109b6b, 32'h42174c93, 32'h41f9d060, 32'hc21784a9, 32'h427cd9b5, 32'hc20af743, 32'hc28316bf};
test_bias[78:78] = '{32'hc21cdcc9};
test_output[78:78] = '{32'hc5681d9b};
test_input[632:639] = '{32'h4203682c, 32'h42588475, 32'h418d93e6, 32'hc008b6a6, 32'hc15d7f99, 32'hc1fd9465, 32'h42b477f6, 32'hc2c7ea83};
test_weights[632:639] = '{32'hc1fc1ea1, 32'h42679fef, 32'h412ed62a, 32'h42a5b515, 32'hc217d6d4, 32'hbf61e433, 32'hc2c308c7, 32'h417ae557};
test_bias[79:79] = '{32'hc210a372};
test_output[79:79] = '{32'hc5f1b02d};
test_input[640:647] = '{32'h41dc0ce7, 32'h41669479, 32'h42bfc482, 32'hc197a3cb, 32'hc2b84f95, 32'h41f1eb16, 32'hc258f737, 32'h42b6cbdc};
test_weights[640:647] = '{32'h415a3e07, 32'hc2b766f8, 32'hc2825a06, 32'hc2a0a2cf, 32'hc285bdef, 32'hc2c16de5, 32'h4265d0b2, 32'hc18094dd};
test_bias[80:80] = '{32'hc2b78190};
test_output[80:80] = '{32'hc5de43c0};
test_input[648:655] = '{32'hc25bb01b, 32'h42409666, 32'h4243f3e4, 32'hc2a14986, 32'h425971ca, 32'hc2536010, 32'h428b416f, 32'h42307490};
test_weights[648:655] = '{32'hc13e1e93, 32'h4291426f, 32'h41fae33f, 32'hc0b40697, 32'hc1179948, 32'hc1ba2f49, 32'h4204f94e, 32'hc260d425};
test_bias[81:81] = '{32'h421d75fc};
test_output[81:81] = '{32'h45d24660};
test_input[656:663] = '{32'h416b912e, 32'h42949553, 32'hc2bb3ef0, 32'hc203e189, 32'h42c54832, 32'h41dfb929, 32'hc288a67d, 32'hc2b48513};
test_weights[656:663] = '{32'hc255af6b, 32'hc1c2326e, 32'h424dd910, 32'hc20db0d7, 32'h42ada67e, 32'hc2bb2f81, 32'h4118ea39, 32'h42c395b4};
test_bias[82:82] = '{32'h41e7673b};
test_output[82:82] = '{32'hc6183ebf};
test_input[664:671] = '{32'h42b8ce38, 32'hc1de97b2, 32'h42aca2ea, 32'h42681993, 32'h42aa7207, 32'h428ae8cb, 32'h414bd18b, 32'hc182d951};
test_weights[664:671] = '{32'hc2722621, 32'h4219bf7d, 32'hc08243e6, 32'h427f920c, 32'hc18c33a6, 32'h429b9d8a, 32'hc2730829, 32'h42a7c7d4};
test_bias[83:83] = '{32'hc18ec479};
test_output[83:83] = '{32'hc4c315a3};
test_input[672:679] = '{32'hc2962938, 32'h4213483c, 32'hc1dd0f37, 32'h41c6f507, 32'hc22fd131, 32'hc1a3b4c6, 32'hc25e88f9, 32'hc2b857be};
test_weights[672:679] = '{32'h42305cb4, 32'hc1906ade, 32'h414910ff, 32'hc29c5faa, 32'hc1c70604, 32'h4201f82b, 32'h4195d4e2, 32'hc13b80c8};
test_bias[84:84] = '{32'h42c7ae5b};
test_output[84:84] = '{32'hc5b22113};
test_input[680:687] = '{32'hc1170336, 32'h4277e7cd, 32'hc295a76c, 32'hc26725b2, 32'h429428f9, 32'hc1c5e3a6, 32'h41e3d7d5, 32'h429a393d};
test_weights[680:687] = '{32'hc25f1b33, 32'h4210dc84, 32'h429447bb, 32'hc22d2334, 32'h418a8c55, 32'h429e85c2, 32'hc2af4577, 32'h427224fc};
test_bias[85:85] = '{32'h42b17b31};
test_output[85:85] = '{32'h44a377d3};
test_input[688:695] = '{32'h422a7b9c, 32'hc20445c7, 32'hc2becfe3, 32'h423a1c0b, 32'h42a829c6, 32'h42b28b27, 32'hc288247b, 32'h41fc8ed5};
test_weights[688:695] = '{32'h4242ef38, 32'h3f03932c, 32'h429a09ef, 32'h420799db, 32'h42b6b54c, 32'hc2862d06, 32'h4212db95, 32'h4114df12};
test_bias[86:86] = '{32'h40b21cb4};
test_output[86:86] = '{32'hc583d41e};
test_input[696:703] = '{32'h42693d4b, 32'h4286e202, 32'hc20c01cb, 32'hc115924b, 32'hc289e243, 32'h4193b617, 32'hc2afd6a6, 32'h4272f43a};
test_weights[696:703] = '{32'h42b03b66, 32'h42813d88, 32'h423fdc07, 32'h429e12f8, 32'h4205d269, 32'hc22b3b3c, 32'h4158197a, 32'hc186d830};
test_bias[87:87] = '{32'hc138a882};
test_output[87:87] = '{32'h44dbd781};
test_input[704:711] = '{32'hc29218b5, 32'h42c56a21, 32'hc28d0447, 32'hc111d727, 32'hc2b5b0bf, 32'h42a868a4, 32'h40fb0a28, 32'hc287c582};
test_weights[704:711] = '{32'hc08ea487, 32'h42238f46, 32'hc2a5047d, 32'h428dcb3f, 32'hc07466e8, 32'h429bb7f9, 32'hc2228116, 32'hc2b16bb8};
test_bias[88:88] = '{32'hc26cbddd};
test_output[88:88] = '{32'h46ac80bd};
test_input[712:719] = '{32'hc274c04c, 32'h411e031f, 32'hc2c5c59c, 32'h42677b41, 32'hc2b63113, 32'hc26a1fa1, 32'hc2a862a1, 32'h41505b0e};
test_weights[712:719] = '{32'h42779ab6, 32'hc1b88e5e, 32'h4299a40a, 32'h4229da71, 32'hc258b2fc, 32'hc0ba0681, 32'h418dae92, 32'hc192da87};
test_bias[89:89] = '{32'h42085f32};
test_output[89:89] = '{32'hc5ae396c};
test_input[720:727] = '{32'h420b4284, 32'hc196f60b, 32'h4082dea3, 32'h4227518b, 32'h4257875b, 32'h4284dae1, 32'hc215e972, 32'h421d3594};
test_weights[720:727] = '{32'hc2c7ad82, 32'hc28348f7, 32'hc2833fbf, 32'h4032afb0, 32'hc08b8feb, 32'hc283c2cb, 32'h4299d0d7, 32'hc1dd9c80};
test_bias[90:90] = '{32'hc0cd2342};
test_output[90:90] = '{32'hc62b8640};
test_input[728:735] = '{32'h429ba58f, 32'h42bb684a, 32'hc294fb8b, 32'hc210dc0f, 32'hc14d965e, 32'h41e92e0a, 32'h41c1edf9, 32'hc1cb8606};
test_weights[728:735] = '{32'h426bde18, 32'hc20df7b7, 32'h42837d2b, 32'h41a1debb, 32'hc29a105f, 32'hc1f023c1, 32'h42804bcf, 32'hc1ac1b44};
test_bias[91:91] = '{32'hc2062117};
test_output[91:91] = '{32'hc5087352};
test_input[736:743] = '{32'hc2a998f3, 32'h42c5c045, 32'hc27017b8, 32'h4283947f, 32'h41a3bb09, 32'h4225377e, 32'hc2893715, 32'hc0c7c32a};
test_weights[736:743] = '{32'hc2a3262f, 32'h418aed59, 32'h427714d2, 32'hc298f68e, 32'hc21e5208, 32'hc1a3ca55, 32'h41ee76f8, 32'h42706238};
test_bias[92:92] = '{32'h41d02cc6};
test_output[92:92] = '{32'hc581d662};
test_input[744:751] = '{32'hc249e23d, 32'h419aa7f3, 32'h418aaab1, 32'hc1772ec4, 32'hc1d69c89, 32'h42b02921, 32'hc1633237, 32'hc2b09435};
test_weights[744:751] = '{32'hc2659e8e, 32'hc22311d0, 32'hc2bca4ec, 32'h423115dc, 32'hc02372cb, 32'h42828a89, 32'h42a80bd7, 32'hc09f37d0};
test_bias[93:93] = '{32'h42b4a7ff};
test_output[93:93] = '{32'h459a82fd};
test_input[752:759] = '{32'hc25b2004, 32'hc2544b43, 32'hc18fe134, 32'h4234a983, 32'h42c591d6, 32'hc0423f2c, 32'hc26c52e9, 32'h41bb0d3e};
test_weights[752:759] = '{32'hc2af318e, 32'hc26b81cf, 32'hc089a7d3, 32'hc2165a77, 32'hc1428a63, 32'hc27bda5c, 32'hc202a30f, 32'h428ccab2};
test_bias[94:94] = '{32'h42826059};
test_output[94:94] = '{32'h460b973f};
test_input[760:767] = '{32'hc21eabfa, 32'hc29e3297, 32'hc27c66b9, 32'h420b9468, 32'hc2a67a2f, 32'h41eeb71b, 32'h4296ae06, 32'h40bb0c99};
test_weights[760:767] = '{32'hc16a0250, 32'h4242879f, 32'hc107ad19, 32'h40044eb1, 32'hc2535b45, 32'hc2271861, 32'hc297196a, 32'h40367fbb};
test_bias[95:95] = '{32'hc211285d};
test_output[95:95] = '{32'hc5a31945};
test_input[768:775] = '{32'hc26d2fac, 32'hc0eecc83, 32'hc2ae92ba, 32'hc25a9872, 32'hc0f060ca, 32'hc2502268, 32'hc284be07, 32'hc2c1dd63};
test_weights[768:775] = '{32'hc2852846, 32'h41b3a013, 32'hc29c6893, 32'h428f6366, 32'h42113af0, 32'hc2b73509, 32'hc2c2f2f2, 32'hc2ac0fad};
test_bias[96:96] = '{32'h425b06a4};
test_output[96:96] = '{32'h46cb7b47};
test_input[776:783] = '{32'hc25a86bc, 32'h42ab31d0, 32'h42a6197d, 32'hc186ae17, 32'hc28c0560, 32'h42930fa6, 32'hc278e49b, 32'hc29ea53b};
test_weights[776:783] = '{32'hc12c31a9, 32'h40f1c1ec, 32'h41943422, 32'h42627dec, 32'hc2b70d45, 32'hc279050c, 32'h41ad0dc9, 32'hc234f38b};
test_bias[97:97] = '{32'h3e8c6c80};
test_output[97:97] = '{32'h45b825c3};
test_input[784:791] = '{32'hc25e9608, 32'h4238e092, 32'hc1af1c34, 32'h42381735, 32'hc194ed8e, 32'h42b4dee2, 32'h4201bf4c, 32'hc23decd3};
test_weights[784:791] = '{32'hc22d06e9, 32'hc24446bf, 32'hc2a4d1b1, 32'hc0d4703f, 32'hc1917324, 32'h428a4cde, 32'hbc9cc3cf, 32'h42671dd9};
test_bias[98:98] = '{32'hc280173a};
test_output[98:98] = '{32'h45a96b8c};
test_input[792:799] = '{32'h42902638, 32'h428048f9, 32'h41984a1c, 32'hc2837a73, 32'h424a48d5, 32'h40a19704, 32'hc20a6df9, 32'hc2b220d3};
test_weights[792:799] = '{32'hc2c35600, 32'hc2091c1d, 32'hc2c4204f, 32'hc28e6273, 32'hc1263261, 32'hc239d1aa, 32'hc184b8c9, 32'hc06c78e0};
test_bias[99:99] = '{32'hc1f20131};
test_output[99:99] = '{32'hc5c53c77};
test_input[800:807] = '{32'hc20d5305, 32'hc1ab7c19, 32'hc2064cbe, 32'hc2748453, 32'h41ee8714, 32'hc2b355f8, 32'h4259ebb6, 32'h41a54730};
test_weights[800:807] = '{32'h42602273, 32'h41e8ddc6, 32'hc2b14a5b, 32'h42b0429a, 32'hc291318f, 32'h42463a68, 32'h42758375, 32'hc2c0caa6};
test_bias[100:100] = '{32'hc26231fc};
test_output[100:100] = '{32'hc6215c7d};
test_input[808:815] = '{32'hc0a25310, 32'h42129c25, 32'h4293a850, 32'h41e1b346, 32'h4292728b, 32'h42b55d3e, 32'hc29d871c, 32'h4153f353};
test_weights[808:815] = '{32'hc2052cb5, 32'hc2b365f9, 32'h42b15df8, 32'h4160ea39, 32'hc299ec0f, 32'h42908fbe, 32'hc28a7441, 32'hc286a405};
test_bias[101:101] = '{32'h4196d0cd};
test_output[101:101] = '{32'h4611b01a};
test_input[816:823] = '{32'h42628d10, 32'h41d1791d, 32'hc242b324, 32'h410feb30, 32'h41a1faf6, 32'h4240e34a, 32'hc28e4764, 32'h429ae717};
test_weights[816:823] = '{32'hc2994662, 32'h4181d37f, 32'hc08d06c8, 32'hbfc72f0f, 32'hc2c08c34, 32'h425add7e, 32'hc29685d3, 32'hc2bfb6a6};
test_bias[102:102] = '{32'h42c1b00e};
test_output[102:102] = '{32'hc59c3a04};
test_input[824:831] = '{32'h411cc09e, 32'h42c26f98, 32'h41ff544e, 32'h421804b4, 32'h42ab29cd, 32'h424b809e, 32'hc14aae64, 32'hc24eceaa};
test_weights[824:831] = '{32'h424af505, 32'hc2c4f64a, 32'h40e4dabf, 32'hc264454a, 32'h42c2d52f, 32'h429a6d14, 32'h4198575f, 32'hc2bce218};
test_bias[103:103] = '{32'hc15da7ee};
test_output[103:103] = '{32'h45b79b6d};
test_input[832:839] = '{32'hc2998d8a, 32'h4271590c, 32'h42591155, 32'hc2921241, 32'h41f73761, 32'hc1db2413, 32'hc1fc8dec, 32'h41c4aed9};
test_weights[832:839] = '{32'hc235cb5a, 32'h426bf29a, 32'hc2151ebc, 32'h41b18a09, 32'hc2552869, 32'hc26c46ea, 32'hc224316e, 32'h42b70416};
test_bias[104:104] = '{32'h3f81c83d};
test_output[104:104] = '{32'h45d85412};
test_input[840:847] = '{32'hc0c4a84e, 32'h428bce25, 32'hc2a674b4, 32'hbf9275c6, 32'hc2b48f20, 32'h42399ffd, 32'hc28529e8, 32'h42592abf};
test_weights[840:847] = '{32'h41a1fb90, 32'h428a8fe0, 32'h4132af29, 32'hc2ba5e25, 32'h428e5bd4, 32'hc2c2412f, 32'hc00715a6, 32'h42a5f703};
test_bias[105:105] = '{32'h41ce7b9b};
test_output[105:105] = '{32'hc513e1a8};
test_input[848:855] = '{32'h416aeb0d, 32'hc2add7dc, 32'h42c3848e, 32'hc2157421, 32'h41b2147a, 32'hc28979c8, 32'hc2224a8e, 32'h424f34e7};
test_weights[848:855] = '{32'h429ee5aa, 32'hc23058d8, 32'h42c70c21, 32'h418234e7, 32'h42904368, 32'hc2028020, 32'hc27e34c7, 32'h4225d5af};
test_bias[106:106] = '{32'h429c924b};
test_output[106:106] = '{32'h46b1e8ce};
test_input[856:863] = '{32'h4283c2b3, 32'hc298d7f0, 32'h4209111b, 32'h42a6ebb8, 32'hc2bcc86f, 32'hc2837ea6, 32'hc1a16fbd, 32'h4295af3e};
test_weights[856:863] = '{32'hc2a5a9c6, 32'hc23b8342, 32'hc1d23b2d, 32'h4210c645, 32'h409a48aa, 32'h421454c1, 32'hc21c1a3a, 32'hc1c01fcf};
test_bias[107:107] = '{32'hc223bd0d};
test_output[107:107] = '{32'hc567231a};
test_input[864:871] = '{32'h42aa48bc, 32'hc1e30015, 32'h428e698a, 32'hc2517e41, 32'hc2951c40, 32'h42aaa127, 32'h42a537a5, 32'hc2a6f5ed};
test_weights[864:871] = '{32'h42b61192, 32'hc211852a, 32'hc25ac5d1, 32'h421c4083, 32'h42b36983, 32'h40cc42bc, 32'hc2c00185, 32'hc2907cc9};
test_bias[108:108] = '{32'hc258bcda};
test_output[108:108] = '{32'hc5a434fa};
test_input[872:879] = '{32'h4272ed41, 32'h42c21891, 32'hc0cf0502, 32'h42a184be, 32'h42a3f6be, 32'h42a16c49, 32'hc1c119b2, 32'hc28ed88a};
test_weights[872:879] = '{32'hc16875c2, 32'h4280a374, 32'h41cec9eb, 32'h4286bdea, 32'h4193b8bd, 32'h42734e3b, 32'h40843a9e, 32'hc08a8592};
test_bias[109:109] = '{32'hc2bc7050};
test_output[109:109] = '{32'h46862770};
test_input[880:887] = '{32'hc26fc4c2, 32'h428c5d7b, 32'hc29bbc6b, 32'h422f4170, 32'h427f4390, 32'h42ac89d6, 32'h429d0b4f, 32'hc19a4bea};
test_weights[880:887] = '{32'h42a7a3d6, 32'h42439415, 32'hc19f0c75, 32'h427abaa4, 32'hc2a4a0b7, 32'hc238d17a, 32'hc219f208, 32'hc28c1427};
test_bias[110:110] = '{32'hc2c5f295};
test_output[110:110] = '{32'hc601cde0};
test_input[888:895] = '{32'h42c5e3fe, 32'h42a2feae, 32'h411754bb, 32'h422d3a8f, 32'hc2bb7d1c, 32'hc2af81ee, 32'h425df1fd, 32'hc2ab1811};
test_weights[888:895] = '{32'h42b7ddb6, 32'hc2354e72, 32'h4291c16b, 32'h42042a69, 32'h4276305b, 32'h42b815c6, 32'hc26a3454, 32'h425e1b1e};
test_bias[111:111] = '{32'h423d400c};
test_output[111:111] = '{32'hc65f0f45};
test_input[896:903] = '{32'h4277cadf, 32'h4266eed3, 32'hc277341b, 32'hc2454db0, 32'h40cb0ae3, 32'h42a2be03, 32'h42964c96, 32'h427136a1};
test_weights[896:903] = '{32'h4229e852, 32'hc23d27aa, 32'hc2be67df, 32'hc24e8a63, 32'hc25c40cd, 32'h424e248d, 32'hc263c840, 32'h42967850};
test_bias[112:112] = '{32'hc1d79cc4};
test_output[112:112] = '{32'h4641d9e4};
test_input[904:911] = '{32'h42b91eea, 32'hc281be08, 32'h42b34052, 32'h420f37b5, 32'h41e8891e, 32'hc166384d, 32'h41d8b594, 32'hc0a4f9e7};
test_weights[904:911] = '{32'hc2b5eb6d, 32'hc1fc4b73, 32'h415a8cf6, 32'hbf87573c, 32'h41b2d3a9, 32'hc2c092bc, 32'h42b6687f, 32'h4139bc10};
test_bias[113:113] = '{32'hc19152f8};
test_output[113:113] = '{32'hc43dd2ff};
test_input[912:919] = '{32'hc0b5e466, 32'h4287c9c1, 32'h420c596f, 32'hc24831be, 32'hc1717af3, 32'hc27e876b, 32'hc29fdbf6, 32'hc2b5fdce};
test_weights[912:919] = '{32'h42ab3dc0, 32'h42475e21, 32'h42ac4a22, 32'h428e5d97, 32'hc22be501, 32'h41b22210, 32'hc2141761, 32'h4244cbb3};
test_bias[114:114] = '{32'hc171d4b4};
test_output[114:114] = '{32'h4260d11c};
test_input[920:927] = '{32'h42652c6b, 32'h427952ff, 32'hc2868ed9, 32'hc247127d, 32'hbfb89345, 32'h41dca41d, 32'hc2275917, 32'h42479630};
test_weights[920:927] = '{32'hc2782bed, 32'hc1c4c348, 32'hc2b9ba98, 32'h40216932, 32'hc1b30706, 32'hc20696f7, 32'h41fa9990, 32'hc15587ed};
test_bias[115:115] = '{32'hc2b2c806};
test_output[115:115] = '{32'hc4f0dec7};
test_input[928:935] = '{32'hc2a4297d, 32'hc2bbcc8b, 32'h4299f5ef, 32'hc2984ae9, 32'hc11a554c, 32'hc1794ae3, 32'h422ee4e8, 32'h411b4a3c};
test_weights[928:935] = '{32'hc2c241f9, 32'hc2105bb9, 32'hc26f7c8f, 32'hc28d5a26, 32'hc03ada1a, 32'h427d70e0, 32'hc265ac42, 32'hc2c45d5f};
test_bias[116:116] = '{32'hc2107a2e};
test_output[116:116] = '{32'h45efdb3a};
test_input[936:943] = '{32'h423a4722, 32'h4287578b, 32'hc29f790b, 32'hc2307ad2, 32'hc29437db, 32'hc29622f2, 32'hc10ee823, 32'h415aca5b};
test_weights[936:943] = '{32'hc03f3c65, 32'hc2b2b42f, 32'hc29bdc64, 32'hc26464cf, 32'h42734304, 32'h41b87b70, 32'hc032fb2c, 32'hc2a2ebfe};
test_bias[117:117] = '{32'hc23ec6ce};
test_output[117:117] = '{32'hc596daa0};
test_input[944:951] = '{32'hc14db8da, 32'h424dedd4, 32'h4299780c, 32'h4290b934, 32'hc2430c4d, 32'h4232acec, 32'hc2a71e9c, 32'h4253f2fb};
test_weights[944:951] = '{32'hc2986fd2, 32'h4113dbd5, 32'hc2bc1b82, 32'h428917e7, 32'hc1c08849, 32'hc2695195, 32'h42731dc9, 32'h41a6d52b};
test_bias[118:118] = '{32'h4209506c};
test_output[118:118] = '{32'hc5c0e4db};
test_input[952:959] = '{32'hc2a07334, 32'hc2614fa2, 32'h41affa14, 32'hc1ea6829, 32'h4159c190, 32'h4212b358, 32'h42984080, 32'h41e3f00c};
test_weights[952:959] = '{32'h41492918, 32'hc2afe44b, 32'h42b956dd, 32'h413930a2, 32'h4157ef68, 32'hc1295215, 32'hc293e0d0, 32'h42057c4b};
test_bias[119:119] = '{32'h42991daf};
test_output[119:119] = '{32'h4451afc4};
test_input[960:967] = '{32'hc2a14d87, 32'h4141fcee, 32'h427c742b, 32'h41851b77, 32'h428c9d9e, 32'hc2a7109f, 32'h428b0bfa, 32'h42bbdc18};
test_weights[960:967] = '{32'hc1b0060f, 32'hc21fb21b, 32'h428597e8, 32'h420655b4, 32'hc081fabe, 32'h4135a4a0, 32'h41f4fee6, 32'hc2650369};
test_bias[120:120] = '{32'hc173a2d8};
test_output[120:120] = '{32'h44c3e870};
test_input[968:975] = '{32'hc180c782, 32'h41d302dd, 32'h41cec7a1, 32'h42b8fad7, 32'hbf8c8aaf, 32'h42b89aa1, 32'h421af6dd, 32'hc2c0f7ce};
test_weights[968:975] = '{32'h4242a75e, 32'h42ae4bf4, 32'hc23af76d, 32'hc283cb48, 32'hc1a8b504, 32'hc2782686, 32'h42bb185d, 32'h429c723c};
test_bias[121:121] = '{32'h4253fd23};
test_output[121:121] = '{32'hc6700367};
test_input[976:983] = '{32'h4259dc4c, 32'h4234057b, 32'h42c43723, 32'hc1c623ae, 32'h429abee5, 32'h41e6e0f2, 32'hc191a280, 32'hc205c789};
test_weights[976:983] = '{32'hc27c9db7, 32'hc1d1518d, 32'h42afff55, 32'hc1e89456, 32'hc237b0aa, 32'h40fb6516, 32'h41b52301, 32'h41474bd1};
test_bias[122:122] = '{32'hc28472f4};
test_output[122:122] = '{32'h4400ae17};
test_input[984:991] = '{32'hbe0750af, 32'hc1f1d799, 32'hc2054554, 32'hc186b939, 32'hc26937f9, 32'h402de397, 32'h42c52193, 32'hc2142141};
test_weights[984:991] = '{32'h428b57bd, 32'hc2880274, 32'h41c66731, 32'h428cd92f, 32'hc290af84, 32'hc221f29d, 32'hc2444bd9, 32'h42bfe318};
test_bias[123:123] = '{32'h424523b7};
test_output[123:123] = '{32'hc583340d};
test_input[992:999] = '{32'h42b781be, 32'h4255dad4, 32'hc29a86f7, 32'h41bfed09, 32'hc1eb3598, 32'hc1db9665, 32'h41e92f63, 32'hc2b19e3b};
test_weights[992:999] = '{32'h4178adb5, 32'hc2b9a975, 32'h423bd9ae, 32'hc28824dc, 32'hc299af6a, 32'h429c8497, 32'h420c5158, 32'hc26a7fcc};
test_bias[124:124] = '{32'h4232001d};
test_output[124:124] = '{32'hc516e067};
test_input[1000:1007] = '{32'h41e57d3c, 32'h429cafe1, 32'hc292d700, 32'hc2428afd, 32'h42b0ae2e, 32'hc2022c94, 32'hc28f218c, 32'h428cbedb};
test_weights[1000:1007] = '{32'h42783eeb, 32'hc2388652, 32'hc2839193, 32'hc297c2cc, 32'hc1372ef6, 32'hc202766f, 32'h428e99d6, 32'hc25bbc42};
test_bias[125:125] = '{32'h4197a0ec};
test_output[125:125] = '{32'hc50a4ea1};
test_input[1008:1015] = '{32'hc0861fb8, 32'hc2849759, 32'hc22a2079, 32'hc11146c1, 32'h42380611, 32'hc1ec24c0, 32'h4145d9df, 32'h4296f45a};
test_weights[1008:1015] = '{32'h419393d3, 32'h42b3cd06, 32'hc1611f9a, 32'h41e30641, 32'hc2017652, 32'h3eef9a78, 32'h42284bbe, 32'hc25cbdf1};
test_bias[126:126] = '{32'hc1d2dd4d};
test_output[126:126] = '{32'hc629dad9};
test_input[1016:1023] = '{32'h42b37877, 32'hc23f70c3, 32'h421b2ea4, 32'hc28fe97f, 32'hc1a5e511, 32'hc1e9dba2, 32'h42810969, 32'hc1241434};
test_weights[1016:1023] = '{32'h41baafb9, 32'h4219e91b, 32'h422a5da1, 32'h40ca14ec, 32'h41a44c5e, 32'h42b3211d, 32'hc208f1b9, 32'h423008f6};
test_bias[127:127] = '{32'hc25c611e};
test_output[127:127] = '{32'hc586a6e0};
test_input[1024:1031] = '{32'hc1598379, 32'hc22502c1, 32'hc1992891, 32'hc2aa33bf, 32'h424eb3a3, 32'hc2820320, 32'h42ad5ae5, 32'hc27c3a54};
test_weights[1024:1031] = '{32'h412f6ef0, 32'h40f1b963, 32'hc1a2dadd, 32'hc22a76fc, 32'h4126557d, 32'h4219792f, 32'h4217c8ec, 32'h42179523};
test_bias[128:128] = '{32'hc2709be5};
test_output[128:128] = '{32'h451861e0};
test_input[1032:1039] = '{32'hc18b267e, 32'h421addb7, 32'h41f28139, 32'h41ea93d7, 32'h3fdcad50, 32'hbea66003, 32'h4250c491, 32'hc10e715c};
test_weights[1032:1039] = '{32'h405959da, 32'h42820109, 32'h40bd50fc, 32'hc21b32e0, 32'hc282f926, 32'hc29656b2, 32'h418dd61e, 32'hc1802d6b};
test_bias[129:129] = '{32'hc264c955};
test_output[129:129] = '{32'h4517588c};
test_input[1040:1047] = '{32'hc0df610d, 32'h427d66eb, 32'hc228edaa, 32'h41d22838, 32'hc2b4a755, 32'h429a73d2, 32'h4213d139, 32'hc28ba816};
test_weights[1040:1047] = '{32'h410added, 32'h42443146, 32'h413edb5e, 32'h421fe68e, 32'h41969e91, 32'hc0710098, 32'hc09f92dc, 32'h427d344c};
test_bias[130:130] = '{32'h42c2ff7c};
test_output[130:130] = '{32'hc535969a};
test_input[1048:1055] = '{32'hc22e802e, 32'hc2b7dbdd, 32'h426f7b8b, 32'hc1edcd5b, 32'h42aebbcd, 32'hc298401b, 32'hc1a64904, 32'h42a48b49};
test_weights[1048:1055] = '{32'h3e815a77, 32'hc267e093, 32'h4168c682, 32'hc21299a9, 32'h40b063f4, 32'hc2159a71, 32'h40a53aec, 32'hc1c40989};
test_bias[131:131] = '{32'h42b9290c};
test_output[131:131] = '{32'h460601d5};
test_input[1056:1063] = '{32'hc2c40029, 32'h42b46c88, 32'hc1a4beb8, 32'hc246cd62, 32'hc22c2322, 32'hc105ab26, 32'hbfccccf7, 32'hc1dfada7};
test_weights[1056:1063] = '{32'h42b72637, 32'h42b8d102, 32'h420c7ba6, 32'hc2382324, 32'h426bdfe2, 32'hc2aa2a6e, 32'hc2352200, 32'h40b3046e};
test_bias[132:132] = '{32'hc1ce453b};
test_output[132:132] = '{32'hc47c7c5d};
test_input[1064:1071] = '{32'hc1b7ed03, 32'hc1f29316, 32'h42c0c5a8, 32'h41dc08c1, 32'h42c21a1f, 32'h42bae9d2, 32'h3f4c5f4c, 32'hc194fcb4};
test_weights[1064:1071] = '{32'h41520572, 32'hbfa44dde, 32'h42075af3, 32'hc297d958, 32'hc1cd5475, 32'hc29d9842, 32'h423aa7ea, 32'h42400d8f};
test_bias[133:133] = '{32'h42ac293f};
test_output[133:133] = '{32'hc617cdba};
test_input[1072:1079] = '{32'h428e3bdd, 32'hc138fcc3, 32'hc2c5fc6d, 32'h42a360d0, 32'hc28d4d8e, 32'h429e2963, 32'h42c4f900, 32'hc23365fa};
test_weights[1072:1079] = '{32'h42813426, 32'h422d1a22, 32'hc149b42a, 32'h426f7976, 32'h42377a1d, 32'hc25fcc23, 32'hc241a6a6, 32'hc2113b6b};
test_bias[134:134] = '{32'h4153d09f};
test_output[134:134] = '{32'hc40bc603};
test_input[1080:1087] = '{32'hc2a8b190, 32'h429ae882, 32'hc18566c3, 32'h4281fe06, 32'hc2b108fe, 32'hc22e4b74, 32'h4295f43b, 32'hc2a8188a};
test_weights[1080:1087] = '{32'hc22f3079, 32'h41fab71b, 32'h427f673e, 32'h4265cdea, 32'h4293cbe8, 32'h3f5bf197, 32'hc2c0937e, 32'h422edbc0};
test_bias[135:135] = '{32'h420a4773};
test_output[135:135] = '{32'hc6071b12};
test_input[1088:1095] = '{32'h4285bd1f, 32'hc28e37c8, 32'h427c4c87, 32'hc1ee50c7, 32'hc2179b66, 32'h424ea108, 32'hc2508c80, 32'hc20aae0d};
test_weights[1088:1095] = '{32'hc1df8885, 32'hc296e5db, 32'hc1cc7c90, 32'hbfa1b6d7, 32'h41908b74, 32'h411ac9cb, 32'hc25c03ed, 32'h428d4b9e};
test_bias[136:136] = '{32'hc1931de4};
test_output[136:136] = '{32'h45058fbf};
test_input[1096:1103] = '{32'hc1f39182, 32'hc272c9c9, 32'h3f0ff8e8, 32'h42afbf2d, 32'hc219e718, 32'hc229093a, 32'hc232bed9, 32'hc29cf8dd};
test_weights[1096:1103] = '{32'hc2ad0931, 32'hc2b12e3c, 32'hbf876f14, 32'hc2c42151, 32'h42c12f8e, 32'hc1c84c41, 32'h412316f1, 32'hc297dd51};
test_bias[137:137] = '{32'h42a64ac0};
test_output[137:137] = '{32'h451123ea};
test_input[1104:1111] = '{32'hc21f1ca9, 32'h40893ac5, 32'hc289da91, 32'h40e196e7, 32'hc175f0a4, 32'hc0afe8d2, 32'hc2aab8eb, 32'hc14b5a8f};
test_weights[1104:1111] = '{32'hc26ec6ad, 32'h42613a5d, 32'h3f5b64a1, 32'h42c19021, 32'hc2b0e9de, 32'h428cc873, 32'h42b6d522, 32'hc25b18f7};
test_bias[138:138] = '{32'hc282c235};
test_output[138:138] = '{32'hc5390b28};
test_input[1112:1119] = '{32'hc2a35179, 32'hc00c353e, 32'hc1ab8b19, 32'h42c61387, 32'h42a5677c, 32'hc262e4cc, 32'hc296f82a, 32'hc1eb09e4};
test_weights[1112:1119] = '{32'h423f2374, 32'hc299b643, 32'h41a71146, 32'hc2a189b7, 32'h42940d2a, 32'hc1fd1059, 32'hc26bc621, 32'h42c18b51};
test_bias[139:139] = '{32'hc19f272d};
test_output[139:139] = '{32'hc5275fc6};
test_input[1120:1127] = '{32'hc121e056, 32'h425819fe, 32'h41a68119, 32'h42540121, 32'hc28dcabf, 32'hc243ed59, 32'h4271c802, 32'hc26a5f7f};
test_weights[1120:1127] = '{32'hc2876921, 32'hc201f343, 32'hc2af3277, 32'hc08d3306, 32'h41bb0d55, 32'h425aaa73, 32'hc0e172d5, 32'h410a05fa};
test_bias[140:140] = '{32'h42b09b9e};
test_output[140:140] = '{32'hc601c625};
test_input[1128:1135] = '{32'h409fccde, 32'hc252c72e, 32'h42a2dab8, 32'hc2bef552, 32'h4290d7cb, 32'h418ff509, 32'hc2814747, 32'h42c04050};
test_weights[1128:1135] = '{32'h419a0fd4, 32'hc29c15ce, 32'hc2a81e0c, 32'hc2805add, 32'h42031554, 32'hc2c64c0d, 32'hc258f056, 32'hc2c01399};
test_bias[141:141] = '{32'hc2a34743};
test_output[141:141] = '{32'hc4d7df9d};
test_input[1136:1143] = '{32'hc18601fe, 32'h40c945f4, 32'hc0fb5660, 32'h42b8b4a2, 32'h428ee456, 32'h420c2303, 32'hc2458539, 32'h41c304ab};
test_weights[1136:1143] = '{32'hc19b82a9, 32'h42519720, 32'h4226810f, 32'h4270ec4e, 32'hc2c2b930, 32'hc17c4368, 32'hc1abee03, 32'h4285e9c0};
test_bias[142:142] = '{32'hc28057c4};
test_output[142:142] = '{32'h447ce2e7};
test_input[1144:1151] = '{32'hc212c929, 32'hc22fc960, 32'h41028284, 32'hc19fa4be, 32'h42a6d821, 32'h42c6c70e, 32'hc222ba81, 32'h429dc683};
test_weights[1144:1151] = '{32'h42a83629, 32'h41d90fa0, 32'hc04fd9de, 32'hc2978fbc, 32'hc2c41a4b, 32'hc1d2881f, 32'hc27e87f1, 32'hc1d5b1d6};
test_bias[143:143] = '{32'hc2945b78};
test_output[143:143] = '{32'hc64df3bf};
test_input[1152:1159] = '{32'h41cf0001, 32'hc250fe68, 32'hc18b0ea1, 32'hc1a3031b, 32'hc0f07ad8, 32'h41ae3593, 32'h42be7cb9, 32'hc188ae36};
test_weights[1152:1159] = '{32'h425cecd9, 32'h42b4d2cb, 32'h42a1c1bf, 32'hc26f0c92, 32'hc1be7dcf, 32'hc26f9821, 32'hc2b00f30, 32'h42b3a004};
test_bias[144:144] = '{32'h42856f18};
test_output[144:144] = '{32'hc661f114};
test_input[1160:1167] = '{32'hc2b5e600, 32'hbf81db1c, 32'hc1247a4e, 32'h428ba945, 32'h421e733b, 32'h4283c197, 32'hc1fb22e9, 32'h4228b305};
test_weights[1160:1167] = '{32'hc2457933, 32'hc28d8018, 32'hc254fac3, 32'hc2bafe84, 32'hc16bef40, 32'hc2993b1c, 32'h425766de, 32'h40ae3508};
test_bias[145:145] = '{32'h41c95a58};
test_output[145:145] = '{32'hc6049bba};
test_input[1168:1175] = '{32'h40e995a4, 32'h41ca1eed, 32'hc2ac9ab8, 32'hc1ec2654, 32'hc1dc34d7, 32'h425046e5, 32'hc2bcaf54, 32'h42b3e88c};
test_weights[1168:1175] = '{32'h42529567, 32'hc2b92d72, 32'hc1b36b00, 32'h41d32ae0, 32'h42bcd5dd, 32'h42905d75, 32'hc248b626, 32'hc2bf2b25};
test_bias[146:146] = '{32'hc0fb2332};
test_output[146:146] = '{32'hc55b7364};
test_input[1176:1183] = '{32'h41cb1829, 32'h421d6f37, 32'h42aa4e2d, 32'h424963f9, 32'h415740dc, 32'h42b01434, 32'hc2b6ea58, 32'hc25f5ec1};
test_weights[1176:1183] = '{32'h421f25ce, 32'hc25e0bd5, 32'h42bce7cc, 32'hc29b55f5, 32'hc2974091, 32'hc281778b, 32'hc19d6d9b, 32'hc299fb60};
test_bias[147:147] = '{32'h428fde16};
test_output[147:147] = '{32'h4516c3f2};
test_input[1184:1191] = '{32'h420f1d0a, 32'h429c11a2, 32'h423582bb, 32'hc2a88670, 32'hc2ad256f, 32'hc178c965, 32'h428b905a, 32'hc2081477};
test_weights[1184:1191] = '{32'h41e3848e, 32'hc2393342, 32'hc29e8206, 32'h424f8a17, 32'hc2b54128, 32'hc2932a3c, 32'h424fcbe4, 32'hc2a75588};
test_bias[148:148] = '{32'hc1e92f7e};
test_output[148:148] = '{32'h4598247d};
test_input[1192:1199] = '{32'h426d6710, 32'hc0a92d64, 32'hc29ae568, 32'hc2bc9fc0, 32'h42362a77, 32'hc101e653, 32'h4223b5cf, 32'h42987520};
test_weights[1192:1199] = '{32'h423f3c4f, 32'h40ea8f34, 32'hc20c32d3, 32'hc19e35fc, 32'h41478416, 32'h42385d37, 32'h4227f1af, 32'h428c0222};
test_bias[149:149] = '{32'hc283bcc8};
test_output[149:149] = '{32'h466383ca};
test_input[1200:1207] = '{32'h42b3ecdc, 32'h42bd7881, 32'hc20f7f3b, 32'hc1a4a72c, 32'hc190364e, 32'hc28edbaa, 32'h42431b4b, 32'h416ca619};
test_weights[1200:1207] = '{32'hc262d533, 32'hbfad1e9b, 32'hc2025a94, 32'h40f2d246, 32'hbf699002, 32'hc202d492, 32'hc2a54983, 32'h411fede5};
test_bias[150:150] = '{32'h41bbf3a3};
test_output[150:150] = '{32'hc5b2dee7};
test_input[1208:1215] = '{32'hc289820b, 32'hc1b61a04, 32'hc2aabdc0, 32'h3f8af707, 32'h42a3fc9b, 32'h422519f5, 32'hc0876afc, 32'hc1b02be3};
test_weights[1208:1215] = '{32'hc0a0e228, 32'hc29526c2, 32'hc1897bb3, 32'h41e09b4b, 32'hc2874317, 32'h4227d595, 32'hc25a4af6, 32'hc299d06f};
test_bias[151:151] = '{32'hc28bc41d};
test_output[151:151] = '{32'h44c5c16e};
test_input[1216:1223] = '{32'hc1b2f2bb, 32'h424a7b2f, 32'hc1dccd81, 32'hc28207dd, 32'hc23df7f7, 32'h42aef5cf, 32'hc1db8b31, 32'h42a886ac};
test_weights[1216:1223] = '{32'h4295ded2, 32'hc23003ff, 32'h42512420, 32'h423c8cd7, 32'h42227632, 32'h40ad51dc, 32'h423acd54, 32'hc2583b68};
test_bias[152:152] = '{32'hc2978734};
test_output[152:152] = '{32'hc6768bf9};
test_input[1224:1231] = '{32'hc2883e1a, 32'hc2ba712c, 32'hc28519f8, 32'hc2a37249, 32'h4254d24e, 32'h422778fd, 32'h429d3850, 32'h42a56629};
test_weights[1224:1231] = '{32'hc2a52321, 32'h41703d3d, 32'h411ee2c1, 32'hc2bc57e7, 32'h427cbcbc, 32'h4162b42c, 32'h420fbf97, 32'h4283f2cb};
test_bias[153:153] = '{32'hc2a7243c};
test_output[153:153] = '{32'h46b6e922};
test_input[1232:1239] = '{32'hc2a3bfe1, 32'hc19971cd, 32'hc2ae2aff, 32'h4200fa23, 32'h42afea75, 32'h42a1aec7, 32'h41881bf1, 32'hc1f091b0};
test_weights[1232:1239] = '{32'hc2c3bbb8, 32'h422c4de9, 32'hc2920e17, 32'h418f7a68, 32'hc23de7c9, 32'hc2797ec9, 32'hc2afb75d, 32'hc1926176};
test_bias[154:154] = '{32'h3f47cff8};
test_output[154:154] = '{32'h4577a524};
test_input[1240:1247] = '{32'h41173a8e, 32'h428c2d6b, 32'hc10fcd00, 32'hc2930494, 32'hc29c9d12, 32'h41adf02b, 32'hc1eddb1b, 32'hc1e0760e};
test_weights[1240:1247] = '{32'h41aa6dad, 32'hc0d5e3c3, 32'h42884f61, 32'hc1e75409, 32'h42b14e92, 32'hc28b0ac2, 32'hc28d9fde, 32'h4276a42a};
test_bias[155:155] = '{32'hc2b760ea};
test_output[155:155] = '{32'hc5d86114};
test_input[1248:1255] = '{32'hc16ea3df, 32'h42ba0b98, 32'h4208a784, 32'h42b18442, 32'hc0e606a0, 32'hc225a0ce, 32'h42bc058d, 32'h42538106};
test_weights[1248:1255] = '{32'hc1c94029, 32'hc12ef833, 32'hc113d337, 32'h42b87304, 32'h422b5141, 32'hc0c4d6aa, 32'h4233d1f8, 32'hc1242068};
test_bias[156:156] = '{32'hc0251f9a};
test_output[156:156] = '{32'h4629a085};
test_input[1256:1263] = '{32'h42a0431c, 32'hc27ed679, 32'h427b81ed, 32'h419d2abd, 32'hc27b053d, 32'h428ea715, 32'hc2c38188, 32'hc1e4f696};
test_weights[1256:1263] = '{32'hc2c05ea8, 32'hc27e9e79, 32'hc25c944a, 32'h40d27498, 32'hc245424d, 32'hbe77feb9, 32'hc248076e, 32'hc2083755};
test_bias[157:157] = '{32'hc291c7b5};
test_output[157:157] = '{32'h44eaaf1b};
test_input[1264:1271] = '{32'h42ace70a, 32'hc1bb36dd, 32'h4218c882, 32'hc1af2572, 32'h42c48469, 32'hc2b1752d, 32'hc2b20b6a, 32'hc24637c7};
test_weights[1264:1271] = '{32'h427cce92, 32'h427c7844, 32'hc2a44c06, 32'h42a1e54e, 32'h4206ac10, 32'h41a2e50e, 32'hc13919b2, 32'h4296a172};
test_bias[158:158] = '{32'hbf9290d2};
test_output[158:158] = '{32'hc504d1f3};
test_input[1272:1279] = '{32'h423d7d79, 32'hc1a74df4, 32'hc2854886, 32'h42be5a0d, 32'h4164c1c4, 32'h427a4a45, 32'h428f83c3, 32'hc2bde814};
test_weights[1272:1279] = '{32'h42c47bda, 32'h422ade82, 32'h428a32eb, 32'hc0b3bc68, 32'hc21bc6a3, 32'h419a70fd, 32'h428e69b4, 32'hc291b596};
test_bias[159:159] = '{32'hc0a2b60e};
test_output[159:159] = '{32'h46307a6e};
test_input[1280:1287] = '{32'hc2764979, 32'h4280998a, 32'h4143b2bc, 32'hc196966b, 32'h40d965a6, 32'hc22ed2dd, 32'h4061f255, 32'h42a1f0b7};
test_weights[1280:1287] = '{32'h414b7887, 32'h425ff128, 32'hc295fe89, 32'hc267d90b, 32'hc16247e2, 32'hc2c49416, 32'hc2b71188, 32'hc12bace0};
test_bias[160:160] = '{32'hc180b2c6};
test_output[160:160] = '{32'h45baf288};
test_input[1288:1295] = '{32'hc2311963, 32'hc2b386f2, 32'h42b81b9f, 32'hc2b6082f, 32'h42a16f17, 32'hc2c350de, 32'hc2c0c86e, 32'hc1b2f2c5};
test_weights[1288:1295] = '{32'hc28919a2, 32'hc2aa231f, 32'hc2b9e88a, 32'h424af3c1, 32'hc2b87f09, 32'hc2976214, 32'h42b3ed2f, 32'hc20e2a97};
test_bias[161:161] = '{32'hc29ba5e8};
test_output[161:161] = '{32'hc624411c};
test_input[1296:1303] = '{32'hc295477b, 32'hc0dc6f53, 32'hc27d1466, 32'h41e49f4f, 32'h40cefea4, 32'h42273a5e, 32'h42b3d009, 32'h42a9eba6};
test_weights[1296:1303] = '{32'hc289e211, 32'h418c86c9, 32'h42b5717a, 32'hc299c38f, 32'h42611afb, 32'hc2b42d59, 32'hc1de644e, 32'h42478916};
test_bias[162:162] = '{32'hc2132846};
test_output[162:162] = '{32'hc590246a};
test_input[1304:1311] = '{32'h41d6ddb9, 32'hc2484841, 32'hc230019c, 32'h419a9461, 32'h41ce3f9f, 32'h42689554, 32'hc2bf5400, 32'hc231149e};
test_weights[1304:1311] = '{32'hc1c651f1, 32'hc2618b5e, 32'hc1e0a5e7, 32'hc1e78cc6, 32'hc273f1dd, 32'hc1e27cf8, 32'hc2484140, 32'h41e11de1};
test_bias[163:163] = '{32'hc037cfb2};
test_output[163:163] = '{32'h4545409d};
test_input[1312:1319] = '{32'h42bfc66d, 32'hc232200c, 32'hc2bd62bd, 32'h41bd7d5d, 32'h42875bbe, 32'h42b1d2c1, 32'h423d8112, 32'hc2c4a9c7};
test_weights[1312:1319] = '{32'hc265685b, 32'h4202838f, 32'hc28f3161, 32'h41c4cab4, 32'h423aa76b, 32'hc20a243c, 32'h4024962e, 32'h421a737d};
test_bias[164:164] = '{32'h4144270c};
test_output[164:164] = '{32'hc545d34d};
test_input[1320:1327] = '{32'h424bd46d, 32'h429cdbfa, 32'hc2498ac3, 32'hc25f5a63, 32'hc1334bd3, 32'hc207ce3b, 32'h40928f09, 32'hc0a23a35};
test_weights[1320:1327] = '{32'hc18c13c8, 32'hc194b396, 32'h41da48e3, 32'hc203cb74, 32'h4197c67b, 32'hc1ab2a75, 32'h41b0646c, 32'h42ae97b7};
test_bias[165:165] = '{32'hc2b41194};
test_output[165:165] = '{32'hc4e15bbe};
test_input[1328:1335] = '{32'h42249f49, 32'h421cd28f, 32'hc286942a, 32'h3f79cc96, 32'hc2a701f3, 32'h41658263, 32'h4189b827, 32'hc08f37af};
test_weights[1328:1335] = '{32'hc2144434, 32'hc2490721, 32'h4233acde, 32'hc288bb6a, 32'hc1cd4ff6, 32'h42a6263d, 32'h428ab977, 32'hc21fac39};
test_bias[166:166] = '{32'h42bd1829};
test_output[166:166] = '{32'hc4dee509};
test_input[1336:1343] = '{32'h421c055a, 32'hc2270eb1, 32'h4283ad84, 32'hc29a169e, 32'hc2782e69, 32'hc1da734b, 32'h429d0266, 32'h4298a0c6};
test_weights[1336:1343] = '{32'h429fec00, 32'hc27b69f7, 32'h429c269e, 32'h42021a23, 32'h42b51111, 32'h42642301, 32'h425c84b2, 32'hc2636b6a};
test_bias[167:167] = '{32'hc24bfc0f};
test_output[167:167] = '{32'h448ebf32};
test_input[1344:1351] = '{32'hc280ee75, 32'hc27ebc4a, 32'h428d88f7, 32'h42c249ce, 32'h4106218d, 32'hc0c367ca, 32'h3fd89789, 32'h410dbed0};
test_weights[1344:1351] = '{32'hc1ba4b69, 32'h42820bbb, 32'hc1984002, 32'h4297d743, 32'h429e23e6, 32'hc284ee4c, 32'h424ef8fb, 32'hc1cfa906};
test_bias[168:168] = '{32'h4108d14e};
test_output[168:168] = '{32'h45871cc3};
test_input[1352:1359] = '{32'h425ef99f, 32'hc0bdf73c, 32'hc0ba8a81, 32'hc2352bf9, 32'h4181d18d, 32'h4182dcf7, 32'h42049380, 32'h4191d656};
test_weights[1352:1359] = '{32'hc283dddb, 32'h41db7bb6, 32'h41e15d1b, 32'hc2abf2d2, 32'hc292484c, 32'hc2016546, 32'h42b5bbfe, 32'hc220dfa9};
test_bias[169:169] = '{32'hc06b280a};
test_output[169:169] = '{32'h43e131a1};
test_input[1360:1367] = '{32'h4278aded, 32'h41e431bd, 32'h429ee4f1, 32'hc0f590fa, 32'hc29b8f79, 32'hc19195ca, 32'hc24dd255, 32'hc28adbe9};
test_weights[1360:1367] = '{32'h42af38c2, 32'h4215e491, 32'hc2acfb6c, 32'hc254d94f, 32'hc2559aa2, 32'hc23b6f85, 32'h4232246e, 32'h4289cb09};
test_bias[170:170] = '{32'hc23dcc5a};
test_output[170:170] = '{32'hc500faec};
test_input[1368:1375] = '{32'hc2914a12, 32'hc2b2b98b, 32'h41d934a4, 32'hc2ad87f4, 32'h4289f03e, 32'hc28621c4, 32'hc2bd8fd0, 32'hc284c61b};
test_weights[1368:1375] = '{32'h41d0aae5, 32'h42a57c8a, 32'hc221f1e9, 32'hc27efa0b, 32'hc2a261b9, 32'h42bf50e1, 32'hc213122a, 32'hc2b3e966};
test_bias[171:171] = '{32'hc22913f8};
test_output[171:171] = '{32'hc5e90f9a};
test_input[1376:1383] = '{32'h42a89a66, 32'hc068e08b, 32'hc25bb43a, 32'hc2bc6cd5, 32'h4232e71b, 32'h41e3c740, 32'hc23eb19f, 32'h425147a9};
test_weights[1376:1383] = '{32'h42a4d1af, 32'hc2579581, 32'hc220c477, 32'h41116255, 32'h42a90176, 32'hc28f2c1e, 32'hbf1a2c73, 32'hc26ef5ba};
test_bias[172:172] = '{32'h4226358d};
test_output[172:172] = '{32'h45e06632};
test_input[1384:1391] = '{32'hc23a2567, 32'h42c19e01, 32'hc29596bb, 32'hc0a74f64, 32'hc2a47606, 32'h423ae5bf, 32'hc2aa9261, 32'hc288be4c};
test_weights[1384:1391] = '{32'h42886181, 32'h4251ec60, 32'h4269af5a, 32'hc28da3ca, 32'hbebe7803, 32'h4260be9d, 32'hc032f5a1, 32'h410acfdd};
test_bias[173:173] = '{32'h414cb247};
test_output[173:173] = '{32'h435de587};
test_input[1392:1399] = '{32'hc2b589ba, 32'h4254d243, 32'h42bdb16b, 32'hc1c25c80, 32'h425924da, 32'hc2af5f3f, 32'hc21a7b0e, 32'h42480e66};
test_weights[1392:1399] = '{32'hc175329a, 32'hc1321961, 32'hc236bd9f, 32'hc2a38b87, 32'h42adadcc, 32'h42b3f4f5, 32'h429e8e1d, 32'hc12e9fea};
test_bias[174:174] = '{32'hc2471a61};
test_output[174:174] = '{32'hc602f29b};
test_input[1400:1407] = '{32'hc23cdd2e, 32'hc2b67242, 32'h42c174b5, 32'h41e8260a, 32'hc2639afd, 32'h4295c4e6, 32'h428aad22, 32'h426b1b2a};
test_weights[1400:1407] = '{32'h4278b5ba, 32'hc232d528, 32'h42a52e7e, 32'h41203413, 32'h42ba29e4, 32'hc2317c65, 32'hc183ebd9, 32'hc207d348};
test_bias[175:175] = '{32'hc1a56b08};
test_output[175:175] = '{32'hc5135169};
test_input[1408:1415] = '{32'h4290d7ea, 32'hc1a81a9e, 32'h42477309, 32'hc0aabc7e, 32'hc2ba65f0, 32'h429ceeb0, 32'h422b3b30, 32'hc29ff46b};
test_weights[1408:1415] = '{32'h42270109, 32'h41428318, 32'h41c3302c, 32'hc287c601, 32'hc26b6652, 32'hc2bdbb0c, 32'hc268b908, 32'h415f97db};
test_bias[176:176] = '{32'hc179b795};
test_output[176:176] = '{32'hc49a79b7};
test_input[1416:1423] = '{32'h411d16d8, 32'h425c64ee, 32'hc285dbcc, 32'h41b41344, 32'h4273ac2e, 32'hc23683a6, 32'hc2156d6d, 32'h41d6b18a};
test_weights[1416:1423] = '{32'hc29adba0, 32'hc2a1bcb9, 32'h422b695b, 32'h40f997b0, 32'h4223c043, 32'hc1104d75, 32'h414de971, 32'hc2448eb8};
test_bias[177:177] = '{32'hc015641c};
test_output[177:177] = '{32'hc5d4a7a7};
test_input[1424:1431] = '{32'hc21434ef, 32'hc2c6554f, 32'h427909f8, 32'h42bcd3d3, 32'hc26a427f, 32'h4119e478, 32'hc2a88619, 32'hc1a564b7};
test_weights[1424:1431] = '{32'h42940268, 32'h3f72c8a6, 32'hc2613ce5, 32'hc237c613, 32'hc2597591, 32'hc208a85f, 32'hc2b177b8, 32'hc0c5a83b};
test_bias[178:178] = '{32'hc27bd2e0};
test_output[178:178] = '{32'hc38d53db};
test_input[1432:1439] = '{32'hc2631d50, 32'h4279b7ab, 32'h420a29fc, 32'h4187fa80, 32'hc20dfbfd, 32'h4248b436, 32'hc2863df2, 32'hc0de3e2a};
test_weights[1432:1439] = '{32'h4258b0c0, 32'h42b5ef57, 32'hc0ed611d, 32'hc2a3e71b, 32'hc2aa4409, 32'h41d08507, 32'hc1cc553a, 32'h42ac0a49};
test_bias[179:179] = '{32'h41ee2924};
test_output[179:179] = '{32'h45c8f3b3};
test_input[1440:1447] = '{32'h41cb6154, 32'h4293f91a, 32'h42a1dac4, 32'hc19ceb5e, 32'hc2c79ba2, 32'hc2c58257, 32'h42b5e1e8, 32'hc179c0de};
test_weights[1440:1447] = '{32'hc18fb9b2, 32'hc0de8ad7, 32'h423583fe, 32'hc2af9ac2, 32'hc2ba69d6, 32'h40990712, 32'hc2175269, 32'h425d230c};
test_bias[180:180] = '{32'h42a8221f};
test_output[180:180] = '{32'h460d2905};
test_input[1448:1455] = '{32'h42a8779c, 32'hc253a8b4, 32'h428e4886, 32'h4275255b, 32'hc26cb4d1, 32'h42944555, 32'hc2560cb8, 32'h41bf7a83};
test_weights[1448:1455] = '{32'hc016fb0d, 32'h42b3db7f, 32'h42ab960e, 32'hc1d6ae08, 32'h3eb235ad, 32'hc21fa57d, 32'hc2c7d16c, 32'h4199cd3f};
test_bias[181:181] = '{32'hc298cced};
test_output[181:181] = '{32'h450cc3c6};
test_input[1456:1463] = '{32'h419240bb, 32'hc1e9ed1e, 32'h415151c7, 32'h4200c454, 32'hc2307cf7, 32'h422a7535, 32'h402fc131, 32'h42a1a10c};
test_weights[1456:1463] = '{32'h422af9ae, 32'h42ab3fc3, 32'h41cfbdc3, 32'hc276e643, 32'hc0bce64d, 32'h4261f0b6, 32'hc2466520, 32'hc205383d};
test_bias[182:182] = '{32'hc276d41f};
test_output[182:182] = '{32'hc5607824};
test_input[1464:1471] = '{32'h42b2dd6d, 32'hc2c0aa37, 32'hc23be731, 32'hc210632c, 32'hc226fd5e, 32'h429526da, 32'h41707716, 32'hc1e3994f};
test_weights[1464:1471] = '{32'hc2c017cb, 32'hc107a126, 32'h4111bae2, 32'hc2b984bc, 32'h429ab240, 32'h4281a4b9, 32'hc17d6af9, 32'h42a7e273};
test_bias[183:183] = '{32'h41c5e71f};
test_output[183:183] = '{32'hc5b6c82a};
test_input[1472:1479] = '{32'hc214f1be, 32'h424fd37d, 32'h42a7fafc, 32'hc2b237db, 32'hc210a138, 32'h42ac9859, 32'hc1364cf2, 32'hc15596dc};
test_weights[1472:1479] = '{32'hc1809da5, 32'h41d10b74, 32'hc2a2c149, 32'h419ce8d9, 32'hc034e97f, 32'h409db022, 32'h4145f26f, 32'h427066b3};
test_bias[184:184] = '{32'hc1d015d0};
test_output[184:184] = '{32'hc5dce176};
test_input[1480:1487] = '{32'h42a1dcb2, 32'h425a07c5, 32'h4250e435, 32'hc2465a27, 32'hbfa72ec6, 32'h42bcc231, 32'h41bbaa08, 32'h42b05849};
test_weights[1480:1487] = '{32'h42b03075, 32'hc116e955, 32'hc281b8c4, 32'h4215b9f3, 32'hc20009b1, 32'h4081b2f3, 32'h42bd3b04, 32'h41cc0e97};
test_bias[185:185] = '{32'h418cfa57};
test_output[185:185] = '{32'h45c4548d};
test_input[1488:1495] = '{32'hc09c96ba, 32'hc285ded6, 32'hc147397e, 32'h42697ea3, 32'hc25fe732, 32'h4196ecd7, 32'h429db5eb, 32'hc243899d};
test_weights[1488:1495] = '{32'hc2b2a9f5, 32'hc1c609f9, 32'hc2c37ac1, 32'hc21fd799, 32'h422c6112, 32'h4295efec, 32'hbf2e6af8, 32'h429440b2};
test_bias[186:186] = '{32'h429e7124};
test_output[186:186] = '{32'hc5621957};
test_input[1496:1503] = '{32'h41cdb0ba, 32'hc1027008, 32'hc095b415, 32'h41efdc0c, 32'hc2a6be07, 32'h428a0db7, 32'h42884367, 32'hc2611885};
test_weights[1496:1503] = '{32'h4295e262, 32'hc2ab3625, 32'hc289104d, 32'h42593029, 32'hc04d54ff, 32'h42522c69, 32'hc2acacd7, 32'hc2552454};
test_bias[187:187] = '{32'h42a476d5};
test_output[187:187] = '{32'h45b11182};
test_input[1504:1511] = '{32'h40ed39bb, 32'hc2b29cbd, 32'h42b8ecd1, 32'h42698768, 32'h42b6ebfa, 32'h41b321cd, 32'h4220a699, 32'hc2859272};
test_weights[1504:1511] = '{32'h428ec4f2, 32'hc2babbf8, 32'hc2c32014, 32'hc23620e9, 32'h42a82b04, 32'hc1bb31f5, 32'h4253f19c, 32'h4208a16f};
test_bias[188:188] = '{32'hc279391d};
test_output[188:188] = '{32'h458159f4};
test_input[1512:1519] = '{32'h4237756d, 32'h4278fe44, 32'h40a7ced2, 32'hc2b46613, 32'hc2113935, 32'hc0643a0e, 32'hbf9cdec3, 32'h4255abf4};
test_weights[1512:1519] = '{32'h428cd855, 32'h418f4ade, 32'h42b4aa12, 32'hc2a6df4f, 32'hc1e84e80, 32'h42c72d7e, 32'h42610bca, 32'h40d8f1da};
test_bias[189:189] = '{32'hc29dba59};
test_output[189:189] = '{32'h464f27aa};
test_input[1520:1527] = '{32'h416f0b65, 32'hc2bbc334, 32'h41023056, 32'hc1877257, 32'hc2005e93, 32'h42403f3b, 32'hc2bf0318, 32'hc286a4db};
test_weights[1520:1527] = '{32'hc1ea5a86, 32'h42a27b38, 32'hc27e648f, 32'hc130de3f, 32'h429f5a5a, 32'h429c9086, 32'h42a33b88, 32'h4205b9a0};
test_bias[190:190] = '{32'h412efdfa};
test_output[190:190] = '{32'hc6869052};
test_input[1528:1535] = '{32'hc29ac1fb, 32'h420c8200, 32'h420988c5, 32'hc25e5159, 32'hc26e4164, 32'h4247cd72, 32'h42b271ee, 32'hc2541e2e};
test_weights[1528:1535] = '{32'h42a91dbc, 32'hc0bb6be7, 32'hc1fce750, 32'h42c1cfe4, 32'hc2a9dfe7, 32'hc205a920, 32'h420d35c8, 32'h42a01e42};
test_bias[191:191] = '{32'h427c1fcf};
test_output[191:191] = '{32'hc629c128};
test_input[1536:1543] = '{32'h4282d4df, 32'h424c97f7, 32'h4242759d, 32'hc292ce6b, 32'h4235fc93, 32'h4286476a, 32'hc00bdcbf, 32'h422d3281};
test_weights[1536:1543] = '{32'hc280e7d1, 32'h4202bdae, 32'hc1dc3a87, 32'hc2a74fca, 32'hc1295092, 32'hc224d975, 32'h429767ef, 32'h4275f5c1};
test_bias[192:192] = '{32'hc19dcadd};
test_output[192:192] = '{32'h44b9d849};
test_input[1544:1551] = '{32'h427912a2, 32'hc2599e5d, 32'h42c25d30, 32'hc23018d9, 32'h42437f99, 32'h424ac298, 32'h42b66a63, 32'hc1de998d};
test_weights[1544:1551] = '{32'hc2583461, 32'hbe2e6718, 32'h429fb31c, 32'h426aa627, 32'hc1ee0426, 32'h42c1422c, 32'hc1162c8a, 32'hc256ea18};
test_bias[193:193] = '{32'hc280f806};
test_output[193:193] = '{32'h45b67bc3};
test_input[1552:1559] = '{32'hc2a593ec, 32'hc2bad0b4, 32'h421afcc7, 32'hc237bbd4, 32'hc289c980, 32'hc0693d2c, 32'hc1b04ba6, 32'hc1b11f52};
test_weights[1552:1559] = '{32'h42b8fea2, 32'hc26a5b9c, 32'h427a3cc5, 32'hc265ee6d, 32'h41f700d0, 32'h42bbad9e, 32'h42a476d4, 32'h424809a2};
test_bias[194:194] = '{32'hc1b85e5a};
test_output[194:194] = '{32'hc51e4335};
test_input[1560:1567] = '{32'hc0cb2d90, 32'hc211d490, 32'h4293b22c, 32'hc1e0150a, 32'hc20f4a29, 32'h42ba1ae8, 32'h425400d4, 32'h409cd0ee};
test_weights[1560:1567] = '{32'h41a27a83, 32'h420eb2a7, 32'hc270b476, 32'h42c64b93, 32'h41f381c5, 32'h42441700, 32'hc213df8d, 32'hc13fbca0};
test_bias[195:195] = '{32'h429002c0};
test_output[195:195] = '{32'hc5deab14};
test_input[1568:1575] = '{32'h419b79b0, 32'hc0ac7a6b, 32'h3ffb279f, 32'h4279b951, 32'h423b2ce5, 32'h42043195, 32'hc22dc9dc, 32'hc0f3e6c6};
test_weights[1568:1575] = '{32'hc27a9cb1, 32'hc1951ac2, 32'hc2ae6a38, 32'h41e712fa, 32'hc298ba36, 32'h429674dc, 32'h42382ad2, 32'hc2a74fe8};
test_bias[196:196] = '{32'h41231d41};
test_output[196:196] = '{32'hc4f09820};
test_input[1576:1583] = '{32'hc2ac7a1e, 32'hc168ba15, 32'h413a51ce, 32'h42c056ac, 32'h42b5d3d5, 32'h427095e1, 32'hc1e38333, 32'hc259c1f5};
test_weights[1576:1583] = '{32'hc1994b55, 32'hc088233b, 32'hc297cee3, 32'h42a036c0, 32'hc084a711, 32'h42b76e59, 32'h4235c890, 32'hc2a6f090};
test_bias[197:197] = '{32'h429dba35};
test_output[197:197] = '{32'h4684d87f};
test_input[1584:1591] = '{32'h42339e1c, 32'h42ac2ef6, 32'hc0d2a67d, 32'h42be36b7, 32'hc2965409, 32'h428538c4, 32'h42b4ff5e, 32'h42c696cb};
test_weights[1584:1591] = '{32'h42299426, 32'hc11bd7e1, 32'hc23510ad, 32'h41ef57c4, 32'h4259416d, 32'hc2891f82, 32'hc281a27d, 32'hc280351f};
test_bias[198:198] = '{32'hc285b37a};
test_output[198:198] = '{32'hc682c587};
test_input[1592:1599] = '{32'h4239dc39, 32'h429d06a9, 32'h3e9de0db, 32'hc276df07, 32'h419ddcf5, 32'hc1d272c2, 32'h406942a4, 32'hc2ba2a7e};
test_weights[1592:1599] = '{32'h429a8df5, 32'h4293809e, 32'hc2b09471, 32'h429832f2, 32'hc2276cdf, 32'h42bb5844, 32'hc2c0975e, 32'hc251c515};
test_bias[199:199] = '{32'hc22b2f9f};
test_output[199:199] = '{32'h45b6f6c1};
test_input[1600:1607] = '{32'hc21a16cb, 32'h406fef99, 32'hc10b3f0a, 32'hc2969cb7, 32'hc2322227, 32'h42438b7f, 32'h40bdbf0c, 32'hc26c75a6};
test_weights[1600:1607] = '{32'hc25cdee8, 32'h428042eb, 32'h4281aa67, 32'hc2ad76e8, 32'hc217cde0, 32'h420a53ff, 32'h4286b596, 32'h4262ec49};
test_bias[200:200] = '{32'hc2307ba5};
test_output[200:200] = '{32'h46083449};
test_input[1608:1615] = '{32'h40c0e5dd, 32'h3fc7adf2, 32'hc24a52ea, 32'hc1e4f8e5, 32'hc1e90bdb, 32'hc2b0493a, 32'hc2b571c9, 32'h414a2cfe};
test_weights[1608:1615] = '{32'h414fb651, 32'hc2878392, 32'h402e3ff2, 32'hc20d08e4, 32'h41490fbf, 32'h4228cb3a, 32'hc2c2feb3, 32'h42996c59};
test_bias[201:201] = '{32'h42c3f263};
test_output[201:201] = '{32'h45d07759};
test_input[1616:1623] = '{32'h40f0f3de, 32'hc2c377ff, 32'h41e2410a, 32'hc29b540a, 32'h4229d457, 32'h4170247f, 32'h419b5f14, 32'hc216e5ec};
test_weights[1616:1623] = '{32'hc03a7a55, 32'hc1a6cf38, 32'hc2924435, 32'h3fa6de25, 32'hc214a9be, 32'hc2242088, 32'h418c73f9, 32'hc188cb02};
test_bias[202:202] = '{32'h427091f3};
test_output[202:202] = '{32'hc4a2a8c8};
test_input[1624:1631] = '{32'hc29517ec, 32'h41f36437, 32'h429bf07c, 32'hc24ac84d, 32'hc2b26054, 32'h423cf032, 32'hc28f635f, 32'h412ed30d};
test_weights[1624:1631] = '{32'h42ab860b, 32'h42998ea0, 32'h4197e339, 32'hc273f855, 32'h41172a02, 32'h41096a46, 32'h41a8c545, 32'h41e471fc};
test_bias[203:203] = '{32'hc21ab370};
test_output[203:203] = '{32'hc491225a};
test_input[1632:1639] = '{32'h4272cecb, 32'hc182861c, 32'h42c24199, 32'hc20d239f, 32'h41f3e985, 32'hc284221e, 32'hc298a48e, 32'hc0ff7372};
test_weights[1632:1639] = '{32'h42842930, 32'hc25e2e8e, 32'hc28497c0, 32'hc2c1dd91, 32'hc23a8e76, 32'h428a6cb8, 32'hc103b8af, 32'hc2117ace};
test_bias[204:204] = '{32'hc2809fa9};
test_output[204:204] = '{32'hc54a9cab};
test_input[1640:1647] = '{32'hc20158f5, 32'hc243f94d, 32'hc255bc1f, 32'hc2b11432, 32'h421441d7, 32'hc20026b7, 32'h40f2bbfe, 32'h414efd7c};
test_weights[1640:1647] = '{32'h42a168bc, 32'hc27a78bc, 32'hc27c72c6, 32'hc20a6cdc, 32'h407fbd79, 32'hc1825816, 32'hc2b26e69, 32'hc23a8886};
test_bias[205:205] = '{32'h42c29fe1};
test_output[205:205] = '{32'h45c76ed0};
test_input[1648:1655] = '{32'h4121a14c, 32'hc295a643, 32'hc25b076c, 32'hc215017b, 32'hc1bbdc05, 32'h41ac9baf, 32'h41098de2, 32'h411ecbf1};
test_weights[1648:1655] = '{32'h4201453b, 32'h4204c6fc, 32'h420f494e, 32'h3fd4bf58, 32'h42c7331e, 32'hc29525d7, 32'h418ac60c, 32'h427f49a8};
test_bias[206:206] = '{32'hc2a6918c};
test_output[206:206] = '{32'hc5e82a41};
test_input[1656:1663] = '{32'h428d171e, 32'hc22e57ed, 32'hc21e52ea, 32'h416c28d2, 32'h425b4882, 32'hc133e994, 32'h423be867, 32'h42b3c4d8};
test_weights[1656:1663] = '{32'hc172a3fc, 32'h4175454d, 32'h41f0774e, 32'h42098d52, 32'h429a7e58, 32'hc2129604, 32'h428dc8cd, 32'h428642f9};
test_bias[207:207] = '{32'h4216d57f};
test_output[207:207] = '{32'h4635b2c4};
test_input[1664:1671] = '{32'h428636f6, 32'hc27c3298, 32'h429d8a0f, 32'hc22dd4ea, 32'h41a2e404, 32'h423ead3e, 32'hc2a31681, 32'h4220afe3};
test_weights[1664:1671] = '{32'hc2af236b, 32'h41194773, 32'h4289276d, 32'h42c30e88, 32'hc29c8248, 32'hc24e7c9f, 32'hc0ac39dd, 32'h40967be4};
test_bias[208:208] = '{32'h42419e21};
test_output[208:208] = '{32'hc607dc50};
test_input[1672:1679] = '{32'hc2a044e6, 32'h3f0af3d2, 32'h427b044a, 32'h42b820ca, 32'h42b87681, 32'hc22d041e, 32'hc269d590, 32'h418613c3};
test_weights[1672:1679] = '{32'hc280d5a7, 32'h429ed1ce, 32'hc28a9f83, 32'hc2928619, 32'h42916cfc, 32'hc24ed15e, 32'hc1be8f96, 32'h42971e44};
test_bias[209:209] = '{32'h425d47d1};
test_output[209:209] = '{32'h45b43e26};
test_input[1680:1687] = '{32'hc29aa0b4, 32'h41d96320, 32'h429a5fbd, 32'hc1d6b754, 32'hbf7b791d, 32'h4283b71e, 32'h40838a0d, 32'hc24908b6};
test_weights[1680:1687] = '{32'h425de202, 32'hc1f6180a, 32'h42122b1d, 32'h41e92a31, 32'h42a72885, 32'hc2c611b1, 32'h4146256d, 32'hc2c3b7a2};
test_bias[210:210] = '{32'hc201f90e};
test_output[210:210] = '{32'hc5948f03};
test_input[1688:1695] = '{32'hc1c91ad6, 32'h42b13063, 32'hc272c235, 32'hc271c1f5, 32'hc1226abd, 32'hc24fca2c, 32'h3ff8c933, 32'hc1eee7aa};
test_weights[1688:1695] = '{32'h4242623f, 32'h4294e32e, 32'h42c3c7b0, 32'hc224136e, 32'h40c47e5e, 32'hbf14ef32, 32'hc2bf6a23, 32'hc2b36c74};
test_bias[211:211] = '{32'h423fcaa3};
test_output[211:211] = '{32'h458a26b2};
test_input[1696:1703] = '{32'hc297640d, 32'hc20c1d3d, 32'hc22425a1, 32'h41cd4068, 32'h4206ccc6, 32'h42bc820a, 32'h422b6487, 32'hc29b9a57};
test_weights[1696:1703] = '{32'h42265cf1, 32'hc20d381d, 32'h3fe1e1bc, 32'h41dbbe5b, 32'h4143665e, 32'h42b171f6, 32'h424055cb, 32'hc2a47a3e};
test_bias[212:212] = '{32'hc2874ab5};
test_output[212:212] = '{32'h467836e8};
test_input[1704:1711] = '{32'h429ded67, 32'h426df90d, 32'hc2bbed3f, 32'h425ee552, 32'hc10db8fb, 32'hc2a85c97, 32'h42b85a83, 32'hc22498df};
test_weights[1704:1711] = '{32'hc2976919, 32'hc2be896b, 32'hc2a56598, 32'hc29b15ac, 32'hc283630d, 32'h4187ff25, 32'hc2bebe25, 32'hc2938bc9};
test_bias[213:213] = '{32'h42668ff5};
test_output[213:213] = '{32'hc6665bd4};
test_input[1712:1719] = '{32'h428e779b, 32'hc2604b6f, 32'h42794955, 32'h42b05436, 32'h4184bf4f, 32'h42bab811, 32'hc2228443, 32'h408cd385};
test_weights[1712:1719] = '{32'hc24502aa, 32'hc2aaaa2c, 32'h4225e427, 32'h427d5c2a, 32'hc1d9b074, 32'h429b1ef5, 32'hc29563ad, 32'hc28a7628};
test_bias[214:214] = '{32'hc2acb23d};
test_output[214:214] = '{32'h46937d61};
test_input[1720:1727] = '{32'hc285b250, 32'hc1fff788, 32'h425d9c90, 32'hc28f0256, 32'hc252a950, 32'h429f8e7b, 32'h42bccb7a, 32'h4206bf86};
test_weights[1720:1727] = '{32'hc18d4227, 32'hc2a4a811, 32'hc24a5e8c, 32'hbfb15735, 32'hc26e19ad, 32'hc0bd82df, 32'hc1e95ae0, 32'hc1fdb3b6};
test_bias[215:215] = '{32'hc18b1594};
test_output[215:215] = '{32'hc2844488};
test_input[1728:1735] = '{32'h424c98bc, 32'h4216ff68, 32'hc1985552, 32'h41240581, 32'h429cd5b5, 32'hc2bb50db, 32'hc0a231de, 32'h41b02cfe};
test_weights[1728:1735] = '{32'hc2b76c8d, 32'h405942f8, 32'hc23cdaa0, 32'h429c2bb6, 32'h42ac1930, 32'hc1eae47f, 32'hc18f4b41, 32'h41533f14};
test_bias[216:216] = '{32'hc27a5796};
test_output[216:216] = '{32'h45d94a81};
test_input[1736:1743] = '{32'hc2003e1f, 32'h4159ff6f, 32'hc2858b8a, 32'h42b0c73d, 32'hc2200608, 32'h41930536, 32'h42b0f625, 32'hc25ed6ef};
test_weights[1736:1743] = '{32'h422a5da3, 32'hc1c4724a, 32'hc2c4b37c, 32'h425ccad3, 32'hc1660bd9, 32'h4096ba19, 32'hc2a11304, 32'h41aa157c};
test_bias[217:217] = '{32'hc1df1d1f};
test_output[217:217] = '{32'h450156a2};
test_input[1744:1751] = '{32'hc1bac784, 32'hc1abcc72, 32'h42078d0f, 32'h428ebdd9, 32'h42604873, 32'hc28efa12, 32'h424bbb5c, 32'hc29361c8};
test_weights[1744:1751] = '{32'hc29a27cb, 32'h42169c2c, 32'hc0446c59, 32'h4266f48c, 32'hc289df7d, 32'hc243fe75, 32'hc29b73ee, 32'h41b37bc9};
test_bias[218:218] = '{32'h428fc5bd};
test_output[218:218] = '{32'hc45fb92e};
test_input[1752:1759] = '{32'hc185621b, 32'hc17480ea, 32'h422df53a, 32'hc110daff, 32'hc29c082a, 32'hc27c19f5, 32'hc29db1a0, 32'hc133fe6c};
test_weights[1752:1759] = '{32'hc27efc03, 32'hc19c66a8, 32'hc20ef11a, 32'hc196d9a8, 32'h40397e95, 32'hc22b944a, 32'hc2c3a493, 32'h41be941d};
test_bias[219:219] = '{32'hc2b89d81};
test_output[219:219] = '{32'h46194098};
test_input[1760:1767] = '{32'h3fdaad90, 32'h41443c32, 32'h421febac, 32'hc26280df, 32'hc2b37765, 32'h42b7d2df, 32'hc2522fc4, 32'h42becea5};
test_weights[1760:1767] = '{32'h428fa5b6, 32'hc23d8964, 32'h428b3ad2, 32'hc29486ad, 32'h42b374d9, 32'h42881645, 32'h42389b2d, 32'hc29c94e3};
test_bias[220:220] = '{32'hc227967a};
test_output[220:220] = '{32'hc5a29ece};
test_input[1768:1775] = '{32'hc1b8f1f6, 32'h424bc0fc, 32'h42308e25, 32'h427cf325, 32'h42037ff9, 32'h42b64b3f, 32'h42117361, 32'hc2731d7a};
test_weights[1768:1775] = '{32'hc130c5ac, 32'h41a60672, 32'hc257bffd, 32'hc2895d10, 32'h42baa02e, 32'h41f0e63a, 32'h429fdd7c, 32'h42afd15d};
test_bias[221:221] = '{32'h42009874};
test_output[221:221] = '{32'hc4fa6d6c};
test_input[1776:1783] = '{32'h4184eede, 32'h4296e5ff, 32'h42815c1a, 32'h4064a05b, 32'hc06bbc66, 32'h41ea540e, 32'h421e0f1d, 32'hc1658bed};
test_weights[1776:1783] = '{32'hc1e6a67b, 32'hc23a2252, 32'hc2c0e25c, 32'hc0f33fd2, 32'h41703a0d, 32'hc2204729, 32'h4227d89c, 32'h42b8e91e};
test_bias[222:222] = '{32'h42587dc1};
test_output[222:222] = '{32'hc62d68ca};
test_input[1784:1791] = '{32'h42b99726, 32'h426801be, 32'h42927425, 32'h422ff571, 32'hc282cb4f, 32'hc2a09a07, 32'h42af7519, 32'h42bfbfe8};
test_weights[1784:1791] = '{32'h41f7703f, 32'hc2a6cdc6, 32'hc26b91dd, 32'hc2c4b877, 32'hc2968b7a, 32'hc19b3abf, 32'h42b52eeb, 32'hc24205f6};
test_bias[223:223] = '{32'h4225d675};
test_output[223:223] = '{32'hc444de24};
test_input[1792:1799] = '{32'h42326ddf, 32'h42093884, 32'h4284bec0, 32'hc2b90bc6, 32'hc14a36e7, 32'hc0cabbee, 32'h417e50f2, 32'hc275adb7};
test_weights[1792:1799] = '{32'hc29cff4a, 32'h41295d91, 32'h421504f8, 32'h42140f9e, 32'hc26cc11b, 32'hc20908a3, 32'hc285ad28, 32'h429106b6};
test_bias[224:224] = '{32'h425b1497};
test_output[224:224] = '{32'hc6062b24};
test_input[1800:1807] = '{32'h408e857f, 32'h42972dc8, 32'h3ee84fba, 32'hc2b1eb64, 32'h42bc7f4b, 32'h41eb7f9e, 32'h4174cba2, 32'h42839648};
test_weights[1800:1807] = '{32'h41991fb7, 32'hc215ffa3, 32'h429fa57c, 32'h409406a9, 32'hc1afd1eb, 32'h42a4505c, 32'hc24d65e8, 32'h42998516};
test_bias[225:225] = '{32'h4145837c};
test_output[225:225] = '{32'h44bb70e1};
test_input[1808:1815] = '{32'h42ae39e0, 32'h42b74dc4, 32'hc21e7696, 32'h428be4fa, 32'h40321d66, 32'h41b47d52, 32'h421b6da5, 32'hc24c0e2e};
test_weights[1808:1815] = '{32'h41f60596, 32'hc23d3579, 32'h40761d69, 32'hc2b39d4f, 32'hc1e3d8a3, 32'h42a39a30, 32'h427505e3, 32'hc25c7545};
test_bias[226:226] = '{32'h426cd035};
test_output[226:226] = '{32'hc4862618};
test_input[1816:1823] = '{32'hc04862fe, 32'h428b3f06, 32'hc2095928, 32'hc25e95fa, 32'hc29c55d7, 32'hbfffde31, 32'h42a4993e, 32'h412f2ca3};
test_weights[1816:1823] = '{32'h421123d9, 32'h42472ee7, 32'h42c7d43c, 32'hc2397d48, 32'h42b6575c, 32'hc184c00e, 32'hc0f6b15a, 32'h42c0724e};
test_bias[227:227] = '{32'h422fb1d0};
test_output[227:227] = '{32'hc580fba1};
test_input[1824:1831] = '{32'hc0f87ee0, 32'hc2112d35, 32'hc253299b, 32'h41df5489, 32'hc25eab75, 32'hbff2098e, 32'hc2455f3b, 32'hc16bf75b};
test_weights[1824:1831] = '{32'h4229d31b, 32'h42c401f9, 32'hc2834382, 32'h41509a8b, 32'h421cab87, 32'hc1f80dda, 32'h429c544a, 32'hc2659a35};
test_bias[228:228] = '{32'hc1e77d22};
test_output[228:228] = '{32'hc5a31793};
test_input[1832:1839] = '{32'hc2497a5a, 32'h427fdbf1, 32'h42119500, 32'hc217f47c, 32'hc19a7f8f, 32'hc21e3dc1, 32'h42af7090, 32'hc20938f0};
test_weights[1832:1839] = '{32'hc2c0946a, 32'hc26a99b4, 32'hc2b4dd8d, 32'hc1f6e399, 32'h42a432a5, 32'hc29ef2a7, 32'h429de0af, 32'hc2ab6bf8};
test_bias[229:229] = '{32'hc180b8a1};
test_output[229:229] = '{32'h46224b55};
test_input[1840:1847] = '{32'h4115fb77, 32'h4026b802, 32'hc2c68d5d, 32'h429e1bda, 32'hc1fd8338, 32'hc28d40b3, 32'h42a24388, 32'h425549ca};
test_weights[1840:1847] = '{32'hc29271eb, 32'h420a5eab, 32'hc247eb0f, 32'h4271b805, 32'hc29b1c4a, 32'hc2c1ccbd, 32'hc2bb5acb, 32'hc1b81a42};
test_bias[230:230] = '{32'hbf19491c};
test_output[230:230] = '{32'h461640b1};
test_input[1848:1855] = '{32'h42bc2b5d, 32'hc203cd93, 32'h42c5546c, 32'h42bdd076, 32'h4228ec55, 32'h3fd7b693, 32'h428c3275, 32'h41c1ddf3};
test_weights[1848:1855] = '{32'h42c3ce06, 32'h423db82a, 32'h4258bb9d, 32'hc275e604, 32'h42c3c093, 32'h41b51e95, 32'hc2b1fad3, 32'h419530c3};
test_bias[231:231] = '{32'h401a14bf};
test_output[231:231] = '{32'h45ad5d68};
test_input[1856:1863] = '{32'h42252bd9, 32'hc2bcfcc0, 32'hc265aab6, 32'h4228c980, 32'hc29e2883, 32'h4261a035, 32'h427e6ec7, 32'hc250833f};
test_weights[1856:1863] = '{32'hc28adb31, 32'h412f7265, 32'hc10e6a76, 32'h4298c034, 32'h429e311f, 32'hc14f099c, 32'h41c1e61f, 32'h42451655};
test_bias[232:232] = '{32'h42bc5a8c};
test_output[232:232] = '{32'hc5fcb3ed};
test_input[1864:1871] = '{32'h421b4ed1, 32'h40e73f64, 32'h413ef117, 32'hc2af4dbf, 32'h42c3d6a8, 32'hc0bdef19, 32'hc2beccba, 32'hc2a0db00};
test_weights[1864:1871] = '{32'h4249ec3c, 32'hc216f714, 32'h425d643a, 32'hc2b3c6fb, 32'hc2c48312, 32'h41f8cd18, 32'h41ef4d60, 32'h42a1f8c1};
test_bias[233:233] = '{32'h41b81a1d};
test_output[233:233] = '{32'hc60b6ce4};
test_input[1872:1879] = '{32'hc2956dae, 32'h42a75055, 32'h420bbea5, 32'h4034187f, 32'hc2bd42c4, 32'h4264f3db, 32'h41a08a53, 32'hc224a189};
test_weights[1872:1879] = '{32'hc29e83c6, 32'h429ef9c0, 32'h4220e3fb, 32'h421722f2, 32'h42a40d9c, 32'h42bd5ef7, 32'hc2821c89, 32'hc0908760};
test_bias[234:234] = '{32'hc1e86a18};
test_output[234:234] = '{32'h46257e95};
test_input[1880:1887] = '{32'hc246f37b, 32'h42c0c37c, 32'h424aa02e, 32'hc1eff110, 32'hc107d05a, 32'hc2c6638f, 32'h421e4e25, 32'h416c197b};
test_weights[1880:1887] = '{32'h4294a949, 32'hc2bccb4b, 32'hc0fcecfa, 32'hbf8f6f42, 32'h42114e65, 32'h4282975e, 32'h4206087f, 32'h41d89106};
test_bias[235:235] = '{32'h42418e7f};
test_output[235:235] = '{32'hc68dfa9d};
test_input[1888:1895] = '{32'h42c5c3e7, 32'h42a8f75a, 32'h42c4e63a, 32'hc1cc5db3, 32'hc1939a0c, 32'h429bc85d, 32'hc282de0b, 32'hc28a8561};
test_weights[1888:1895] = '{32'h413b032c, 32'hc199a8dc, 32'hc26741d4, 32'hc2b2f963, 32'hc22754a3, 32'hbf714b70, 32'hc23d24c2, 32'hc245cc94};
test_bias[236:236] = '{32'hc2ba063e};
test_output[236:236] = '{32'h454b3ae0};
test_input[1896:1903] = '{32'h42b4713d, 32'h410785cc, 32'hc2a9f7f2, 32'hc1eaeb4c, 32'hc2253f01, 32'hc229740b, 32'hc2174e06, 32'h428ec22e};
test_weights[1896:1903] = '{32'hc20690bc, 32'hbfa4c5e2, 32'hc228e38d, 32'h41b5aca3, 32'hc2aa8873, 32'hc27189dd, 32'h4272af4f, 32'h4295b4c8};
test_bias[237:237] = '{32'h4242b122};
test_output[237:237] = '{32'h460d723a};
test_input[1904:1911] = '{32'h41fe2d9f, 32'hc2743470, 32'h427a8f81, 32'h41d9bfd5, 32'hc2a52c84, 32'hc225da2e, 32'h429bfdad, 32'h42601ce0};
test_weights[1904:1911] = '{32'hc155ae83, 32'hc2c58f54, 32'hc0c9e96c, 32'h429da409, 32'hc21b4990, 32'h420d5a9b, 32'hc089e150, 32'hc20118ed};
test_bias[238:238] = '{32'hc1ec32e0};
test_output[238:238] = '{32'h45d85c3b};
test_input[1912:1919] = '{32'hc2719d2d, 32'hc22c3a0a, 32'h42b991db, 32'h42c60b92, 32'h41591b28, 32'hc296929e, 32'h42468392, 32'hc2b94ae5};
test_weights[1912:1919] = '{32'hc1f76daa, 32'hc0f6cc1f, 32'h41cda91a, 32'h42a7f132, 32'h42b9c4fd, 32'h41ff0eba, 32'h42a8e6cb, 32'h42a2c78b};
test_bias[239:239] = '{32'hc2c79cbd};
test_output[239:239] = '{32'h4601de2e};
test_input[1920:1927] = '{32'h429e7816, 32'hc1a1ddf3, 32'hc1ddafc8, 32'h4273f41e, 32'h41eb2a77, 32'h40512f59, 32'h42b0d223, 32'h41b0f792};
test_weights[1920:1927] = '{32'hc2211d4c, 32'hc283b24c, 32'h42779afd, 32'hc22f4533, 32'h42826196, 32'h428c9cd5, 32'hbe9b7774, 32'hc280832e};
test_bias[240:240] = '{32'h405d921a};
test_output[240:240] = '{32'hc5ad4bf0};
test_input[1928:1935] = '{32'h4207d4ee, 32'hc26fc165, 32'h420b237e, 32'hc1b1b44e, 32'hc21ab110, 32'h421007b5, 32'h416743ad, 32'hc201460b};
test_weights[1928:1935] = '{32'h429839e5, 32'hc22a82fd, 32'hc2a8a5f8, 32'hc084ce50, 32'h41aaa789, 32'h42c4513e, 32'h42188a23, 32'hc2aa273b};
test_bias[241:241] = '{32'hc18061e9};
test_output[241:241] = '{32'h46019396};
test_input[1936:1943] = '{32'h428810fc, 32'h42261f4c, 32'hc25a7379, 32'hc2311620, 32'h4267d3b7, 32'h428c394d, 32'hc226003b, 32'h42802a82};
test_weights[1936:1943] = '{32'hc1bbf4f0, 32'hc1fcf262, 32'hc25af373, 32'h411d9c66, 32'h4245591d, 32'h420e7730, 32'h42c13626, 32'hc1a8e19f};
test_bias[242:242] = '{32'hc295306e};
test_output[242:242] = '{32'hc3db2380};
test_input[1944:1951] = '{32'h42a5684b, 32'hc2a6678e, 32'h4228c60d, 32'h4047fdcc, 32'hc28d1587, 32'hc22b1060, 32'hc2a6ab44, 32'h429647cc};
test_weights[1944:1951] = '{32'hc264da08, 32'hc11c40c5, 32'hc2bfb242, 32'hc26ec3d1, 32'hc10b5d49, 32'hc2ac924c, 32'hc293ffcb, 32'h42909f65};
test_bias[243:243] = '{32'h42a120de};
test_output[243:243] = '{32'h45f4db81};
test_input[1952:1959] = '{32'h428e966d, 32'hc1c2bbcb, 32'h429f6b6f, 32'h41ac7700, 32'h42b31510, 32'h42a668bd, 32'h4226f443, 32'h41ec8bcf};
test_weights[1952:1959] = '{32'hc243bf7f, 32'hc19e611d, 32'hc002d801, 32'h42a6f378, 32'h42a358f2, 32'hc247e4fa, 32'h4242cffb, 32'h42913ab5};
test_bias[244:244] = '{32'hc288f693};
test_output[244:244] = '{32'h45b84120};
test_input[1960:1967] = '{32'h42c1bf34, 32'h417146c5, 32'hc2877225, 32'hc0ef4805, 32'h3f47ce32, 32'hc2275840, 32'hc26af5cb, 32'hc2874eaf};
test_weights[1960:1967] = '{32'h42877518, 32'h42703719, 32'h4144afeb, 32'h423d5243, 32'h421be711, 32'h428367ee, 32'h3fdafd4e, 32'hbeaa3d37};
test_bias[245:245] = '{32'hc07debae};
test_output[245:245] = '{32'h45597f89};
test_input[1968:1975] = '{32'hc106bd6c, 32'h408c70d6, 32'hc21b20b7, 32'h42c1b0a4, 32'h417175a1, 32'hc163381e, 32'hc1951cff, 32'h41dcd414};
test_weights[1968:1975] = '{32'h41614250, 32'hc19b2587, 32'h41b1f70c, 32'h42c00ffe, 32'hc1d9e100, 32'hc1b0877e, 32'hc22e1146, 32'h4224614d};
test_bias[246:246] = '{32'hc16b314b};
test_output[246:246] = '{32'h461d4b8e};
test_input[1976:1983] = '{32'h41a49b67, 32'hc2a4328e, 32'h41187280, 32'h4287fe64, 32'h41591efd, 32'h421da905, 32'h42b90120, 32'h42037a7f};
test_weights[1976:1983] = '{32'hc1e35a82, 32'hc28d46ac, 32'hc19c4ecb, 32'hc2463626, 32'h429e05ae, 32'h427251ed, 32'hc0a2b454, 32'hc26cf89e};
test_bias[247:247] = '{32'hc1b759d6};
test_output[247:247] = '{32'h452765b3};
test_input[1984:1991] = '{32'h4240a805, 32'h429abd18, 32'h4163cac2, 32'h411db181, 32'hc2994e26, 32'hc2adf4e2, 32'hc299396d, 32'h41acde9f};
test_weights[1984:1991] = '{32'h42af8bc3, 32'h42899ee6, 32'hc13ef591, 32'hc2b6d59b, 32'h424f2dff, 32'h419993d1, 32'hc1c41313, 32'hc22f9288};
test_bias[248:248] = '{32'h42b207fa};
test_output[248:248] = '{32'h45712b42};
test_input[1992:1999] = '{32'hc2c4f129, 32'hc2ac0b49, 32'h42b3306c, 32'h424f55e7, 32'hc1e69789, 32'hc2219906, 32'hc1d09960, 32'h419f2b42};
test_weights[1992:1999] = '{32'h4264759f, 32'h42514894, 32'hc19760ae, 32'h412b6cfe, 32'h4280f720, 32'h42bea1a9, 32'h42869b4a, 32'hc16bac62};
test_bias[249:249] = '{32'h42539df5};
test_output[249:249] = '{32'hc69432a1};
test_input[2000:2007] = '{32'hc20b764e, 32'h427dfc4e, 32'hc178276f, 32'hc0c71e7a, 32'hc18f6e29, 32'h42952f04, 32'h42224420, 32'h41b9e5b8};
test_weights[2000:2007] = '{32'h429e2c36, 32'hc24ad066, 32'h427c775f, 32'hc1f3a81f, 32'hc282368c, 32'h429c5753, 32'hc2bb9c05, 32'h418c1070};
test_bias[250:250] = '{32'hc210a17f};
test_output[250:250] = '{32'hc5482c2e};
test_input[2008:2015] = '{32'h42c085f2, 32'h420fcb58, 32'h42b411e8, 32'h419ed757, 32'hc1c26ebb, 32'hc20ac36b, 32'h429281ba, 32'h3e48d582};
test_weights[2008:2015] = '{32'h4207ba83, 32'hc1a3fadc, 32'hc1883fbc, 32'h42b5aad5, 32'hc2393dbc, 32'hc2c3300a, 32'h4212cdd6, 32'hc2b6568a};
test_bias[251:251] = '{32'hc277621d};
test_output[251:251] = '{32'h461afe0d};
test_input[2016:2023] = '{32'h42b50384, 32'h42262075, 32'hc2c132d9, 32'h428a0ebd, 32'hc215e64a, 32'h428dd6cd, 32'h42b3681c, 32'hc2bc6eae};
test_weights[2016:2023] = '{32'h42b60ec2, 32'h428b08e7, 32'h424df051, 32'h42af2d26, 32'h423a3ddc, 32'h42936a6c, 32'hc2a1464d, 32'h41a76b7c};
test_bias[252:252] = '{32'h41c0f3c6};
test_output[252:252] = '{32'h45cb20b1};
test_input[2024:2031] = '{32'h41bca04a, 32'h4285df16, 32'h42b3fe88, 32'hc2c24a0b, 32'hc1f1652f, 32'h42a88c4c, 32'hc2336416, 32'h42a9fbfa};
test_weights[2024:2031] = '{32'hc20e6752, 32'h4278c372, 32'hc28230f6, 32'h418c1a18, 32'hc157ca31, 32'hc269b4ab, 32'h42ae3e7d, 32'h4272e3e5};
test_bias[253:253] = '{32'hc20b48a5};
test_output[253:253] = '{32'hc5eb724a};
test_input[2032:2039] = '{32'hc2bbb63c, 32'h42a62f74, 32'h427d1fb4, 32'h4232963c, 32'h420b28e6, 32'hc29e9898, 32'h421159c6, 32'hc11aa39e};
test_weights[2032:2039] = '{32'hc16542af, 32'hc2a716f0, 32'hc2b4bba2, 32'hc24c31c4, 32'h429a47df, 32'hc2ac486e, 32'hc29edb42, 32'h429ec811};
test_bias[254:254] = '{32'hc2c3d248};
test_output[254:254] = '{32'hc5f4bd2e};
test_input[2040:2047] = '{32'hc18cca65, 32'hc18f5884, 32'hbee57e1a, 32'h42b352ed, 32'hc2378739, 32'hc1d70956, 32'h41cb54e6, 32'hc1fdad68};
test_weights[2040:2047] = '{32'hc1a6cd3b, 32'hc19ee4a0, 32'h41f5c359, 32'h41ad9509, 32'h42a72762, 32'hc0b7340d, 32'hc2429b55, 32'hc2b83792};
test_bias[255:255] = '{32'hc2c4d4af};
test_output[255:255] = '{32'h440bdf52};
test_input[2048:2055] = '{32'hc18d9ac7, 32'h42a1fcab, 32'h4280ae6f, 32'hc2bdbffd, 32'hc24f3d14, 32'h4191cc43, 32'hc1694c0d, 32'hbfa7bffb};
test_weights[2048:2055] = '{32'h42531db1, 32'h429a3976, 32'hc2c74817, 32'h42c4bfc9, 32'hc28a2539, 32'hc1fdf35a, 32'hc2814233, 32'h424759ea};
test_bias[256:256] = '{32'h42a1f78d};
test_output[256:256] = '{32'hc5ca55da};
test_input[2056:2063] = '{32'h42a4fbc3, 32'h42b0c596, 32'h42444bb0, 32'h42ac5d4f, 32'h415c20f1, 32'h4258fd75, 32'h42697527, 32'hc17c5e55};
test_weights[2056:2063] = '{32'h420801b1, 32'hc2be5c28, 32'hc2887947, 32'h42a403e7, 32'hc10dec58, 32'hc1dac8bc, 32'hc2ae81f0, 32'h41574e50};
test_bias[257:257] = '{32'h4231f1a0};
test_output[257:257] = '{32'hc608ca94};
test_input[2064:2071] = '{32'h422e1d08, 32'h4167d12f, 32'h429ebe96, 32'hc0ac0e29, 32'hc2a44891, 32'hc2954997, 32'hc2743d42, 32'h428715a8};
test_weights[2064:2071] = '{32'h42a9caab, 32'h42ab303e, 32'h41dd51ac, 32'hc1b5a5ad, 32'h429de370, 32'hc21b0ebe, 32'h42aea404, 32'h418dee49};
test_bias[258:258] = '{32'hc273f0de};
test_output[258:258] = '{32'hc405088a};
test_input[2072:2079] = '{32'hc15efc04, 32'hc28245f4, 32'hc00f495f, 32'hc19c4c72, 32'h42211fcb, 32'h41a3f2e8, 32'h41022b46, 32'h42bfa2b7};
test_weights[2072:2079] = '{32'hc2bcc2dd, 32'hc23d26c8, 32'h42681691, 32'hc1312b21, 32'hc21b47e6, 32'h42171f88, 32'hc295e6ee, 32'hc25546e3};
test_bias[259:259] = '{32'hc258d386};
test_output[259:259] = '{32'hc50206a8};
test_input[2080:2087] = '{32'h423f3b45, 32'h42999607, 32'hc23ad944, 32'h40f0fc0f, 32'h42a0f6b8, 32'hc2616853, 32'h428e20bf, 32'h42805171};
test_weights[2080:2087] = '{32'hc2804725, 32'hc2998b90, 32'hc2c5c931, 32'hc1a950f4, 32'h4176d152, 32'hc1f28955, 32'hc2b76a93, 32'h413c7b77};
test_bias[260:260] = '{32'h42019bb9};
test_output[260:260] = '{32'hc5e38692};
test_input[2088:2095] = '{32'hc2858146, 32'h420f6968, 32'h42a3b5ba, 32'h428c68bb, 32'h4242f024, 32'h429094f0, 32'hc1c32a6f, 32'h41d95afa};
test_weights[2088:2095] = '{32'h3f8c628f, 32'h41813625, 32'hc2a7d68d, 32'h4292c8f6, 32'h42c75b47, 32'hc2962155, 32'h41540d7f, 32'hbfc2eee3};
test_bias[261:261] = '{32'hc226fa50};
test_output[261:261] = '{32'hc508a07f};
test_input[2096:2103] = '{32'hc2949929, 32'h425a7347, 32'hc235de35, 32'hc193b44a, 32'h41a190ad, 32'h422f0f0c, 32'h42b3ef1d, 32'h4299e656};
test_weights[2096:2103] = '{32'hc25ddc0e, 32'h42aa7fb9, 32'hc0a0cc91, 32'h41461076, 32'h42b2cfb2, 32'h428954fb, 32'hc22234ce, 32'h428a5228};
test_bias[262:262] = '{32'hc2983ab7};
test_output[262:262] = '{32'h466d434b};
test_input[2104:2111] = '{32'h42951082, 32'hc2a27dd6, 32'hc036fb4c, 32'hc05b5f02, 32'h41a133c9, 32'h426fea24, 32'hc2877c9b, 32'hc104d96d};
test_weights[2104:2111] = '{32'h41eeb853, 32'hc284deaf, 32'h427c9b83, 32'hc1f04f44, 32'hc29abb20, 32'h4251ee8b, 32'hc17d5105, 32'hc263fe78};
test_bias[263:263] = '{32'hc24e2ebc};
test_output[263:263] = '{32'h46260cb4};
test_input[2112:2119] = '{32'h42960e7d, 32'h42bbe6ab, 32'h4234dcdf, 32'hc2775f3f, 32'h421cf111, 32'h422bb5ef, 32'hc2164aec, 32'hc2476d6c};
test_weights[2112:2119] = '{32'h4297305b, 32'hc2ab66c3, 32'hc2999d2b, 32'hc2adcb62, 32'h42514606, 32'hc2ad43bd, 32'h423c2e70, 32'hc1e3daa2};
test_bias[264:264] = '{32'h420d7fcb};
test_output[264:264] = '{32'hc51993e7};
test_input[2120:2127] = '{32'hc2280277, 32'h42998cd8, 32'h428383a3, 32'hc21d5a4a, 32'h42867425, 32'hc23035c7, 32'h3e9eaa22, 32'h406152f6};
test_weights[2120:2127] = '{32'hc29fd5c4, 32'hc0bdbdcf, 32'hc0d79ad3, 32'hc1f96c17, 32'h419c838d, 32'h42136c24, 32'h41e4f287, 32'h428e6abd};
test_bias[265:265] = '{32'hc18121c8};
test_output[265:265] = '{32'h4562403a};
test_input[2128:2135] = '{32'h42a0cd96, 32'hc2243be9, 32'h42758e3d, 32'h425b4c32, 32'h421c2d4b, 32'h41479000, 32'hc198de57, 32'h420e0dc3};
test_weights[2128:2135] = '{32'h42c699cb, 32'h4204ce08, 32'h427349a9, 32'h4256ec7b, 32'hc2a44229, 32'hc25aa095, 32'hc1439236, 32'h420a1740};
test_bias[266:266] = '{32'hc27420f9};
test_output[266:266] = '{32'h4628e9c0};
test_input[2136:2143] = '{32'hc297130a, 32'hc0e41592, 32'h406fdedf, 32'h42b74970, 32'h42ac7254, 32'hc28f2899, 32'hc1244ba6, 32'h429895eb};
test_weights[2136:2143] = '{32'hc2405b4b, 32'h414bb993, 32'h4165bdd7, 32'h41e95082, 32'hc2959e0d, 32'hc2b527b3, 32'h416fd5b2, 32'h428a04c4};
test_bias[267:267] = '{32'h41d4dcc3};
test_output[267:267] = '{32'h4632bc7f};
test_input[2144:2151] = '{32'hc215a54b, 32'hc2971d16, 32'h429be9ab, 32'h42c6167d, 32'hc2a0bb2d, 32'h41eb1aa9, 32'h417b5890, 32'h42c5faff};
test_weights[2144:2151] = '{32'hc1ba4326, 32'hc2c2ddb8, 32'hc214cf59, 32'h42be8256, 32'h42a0cf05, 32'hc202289a, 32'hc2845bfb, 32'hc0fddd54};
test_bias[268:268] = '{32'hc263877f};
test_output[268:268] = '{32'h45aad92f};
test_input[2152:2159] = '{32'h42b0b648, 32'h4282c44d, 32'hc251ce15, 32'h4287e118, 32'hc1bac391, 32'hc1cf7e45, 32'h428b164c, 32'hc2b94321};
test_weights[2152:2159] = '{32'hc2922d5b, 32'h407ebb4f, 32'hc205209b, 32'h40242d78, 32'h42492e9a, 32'h4298056e, 32'hc2389f91, 32'hc2976ff6};
test_bias[269:269] = '{32'hc1b2dd98};
test_output[269:269] = '{32'hc56398c5};
test_input[2160:2167] = '{32'hc1101a78, 32'hc2b31657, 32'hc25ee3d3, 32'hc2b0a9f0, 32'hc2b23faf, 32'h42c1ef22, 32'hc295283a, 32'h4290011d};
test_weights[2160:2167] = '{32'hc17ff09e, 32'h42bdbc21, 32'hc20f6d87, 32'h4293a8c4, 32'h4254c09b, 32'h4294020c, 32'hc28f3a60, 32'h41580330};
test_bias[270:270] = '{32'h4191f53a};
test_output[270:270] = '{32'hc5805b12};
test_input[2168:2175] = '{32'hc2554e20, 32'hc24fd501, 32'hc27b374e, 32'h4144b624, 32'hc2910d96, 32'h4249e813, 32'hc22ea357, 32'hc2b63916};
test_weights[2168:2175] = '{32'h42933ca5, 32'h42b9882c, 32'hc20bf0d2, 32'hc2bf7132, 32'hc224f2ab, 32'h42ae6c0f, 32'h4200f09f, 32'h427726b6};
test_bias[271:271] = '{32'hc2a3caf0};
test_output[271:271] = '{32'hc5e8da76};
test_input[2176:2183] = '{32'h42b21d64, 32'hc0df75ab, 32'hc2b3ac16, 32'h4277aa9b, 32'hc1d87c1f, 32'h425cd0ea, 32'hc1e4eaf3, 32'h42bfe217};
test_weights[2176:2183] = '{32'h4134f279, 32'hc289cee9, 32'hc08e8e5c, 32'hc2b1b7e8, 32'hc22b9dfb, 32'hc22c4f76, 32'h42a54ac1, 32'hc175c112};
test_bias[272:272] = '{32'h42910598};
test_output[272:272] = '{32'hc6065179};
test_input[2184:2191] = '{32'h4262d2ad, 32'h418360b8, 32'h4280a7b9, 32'h42b9d22c, 32'hc25b8b1f, 32'hc1b216d9, 32'hbf04fcc7, 32'h42283833};
test_weights[2184:2191] = '{32'h414e09b9, 32'hc295b4f7, 32'h41675286, 32'hbfefdcbd, 32'h416ca278, 32'h42aa22aa, 32'h4138d92b, 32'h41d8b51e};
test_bias[273:273] = '{32'hc28ebc37};
test_output[273:273] = '{32'hc4ad579e};
test_input[2192:2199] = '{32'h42acf528, 32'h417cc76f, 32'h41e20ef6, 32'hc1b8887a, 32'hc2adf44c, 32'hc247facf, 32'h42bc5243, 32'h42bdce03};
test_weights[2192:2199] = '{32'hc2354823, 32'h3f89d542, 32'hc2bdd439, 32'h428ebadc, 32'h42a92c5b, 32'hc28d9173, 32'h426bb8f3, 32'hc036286c};
test_bias[274:274] = '{32'h427fc002};
test_output[274:274] = '{32'hc5d18f4b};
test_input[2200:2207] = '{32'hc20bfc73, 32'h423e1862, 32'h41f27bed, 32'hc21a4b20, 32'hc1f97065, 32'h429090fa, 32'hc282ebe0, 32'hc29dc07e};
test_weights[2200:2207] = '{32'h4236ff76, 32'hc212d00c, 32'hc2aadbb5, 32'h42983c79, 32'h4290d4ca, 32'h42c08661, 32'h41c61bbd, 32'hc1617b40};
test_bias[275:275] = '{32'h412efaa3};
test_output[275:275] = '{32'hc591e95d};
test_input[2208:2215] = '{32'hc1b3cfb7, 32'hc25a3dd4, 32'hc29087db, 32'hc2948138, 32'h42658ce5, 32'hc1bbb195, 32'hc183687b, 32'h42ac37ee};
test_weights[2208:2215] = '{32'hc24d7593, 32'h4094905d, 32'hc292585f, 32'hc2a49910, 32'h423e1391, 32'h423303fa, 32'h42b85479, 32'h42787c3a};
test_bias[276:276] = '{32'hc2bb0fa8};
test_output[276:276] = '{32'h468a6d70};
test_input[2216:2223] = '{32'h42958c29, 32'h42abff1a, 32'h42847668, 32'hc20d2e55, 32'h4131cb14, 32'h4138e490, 32'h422c5369, 32'h42bb0312};
test_weights[2216:2223] = '{32'hc29bf1d0, 32'h429c125b, 32'hc1ae6e82, 32'h41c3c2c8, 32'h425485ef, 32'hc2a14c9c, 32'hc1912c75, 32'h42a7c0f6};
test_bias[277:277] = '{32'h42306e0c};
test_output[277:277] = '{32'h45a6c4f1};
test_input[2224:2231] = '{32'hc2a134f9, 32'hc2b9e6bf, 32'hc1e5c171, 32'hc1b74ccd, 32'hc1388297, 32'hbfcc69fe, 32'hc2a787ef, 32'h3f720a19};
test_weights[2224:2231] = '{32'hc26115ed, 32'h4295769d, 32'hc2af2122, 32'hc288e8b0, 32'hc2a489d8, 32'hc21538c4, 32'h42396b6d, 32'hc1861ddc};
test_bias[278:278] = '{32'hc2132a53};
test_output[278:278] = '{32'hc49cd67c};
test_input[2232:2239] = '{32'hc2aa458a, 32'hc2b4f5b5, 32'h42083c0a, 32'h4222b06e, 32'hc0d70217, 32'h42230e3d, 32'hc28bd82b, 32'h42a86c3a};
test_weights[2232:2239] = '{32'h41b64efc, 32'h420f6c19, 32'hc2af6e6a, 32'h41cc8180, 32'h421261d5, 32'hc2770e07, 32'hc2686236, 32'hc2172747};
test_bias[279:279] = '{32'hc1c7216b};
test_output[279:279] = '{32'hc60d4274};
test_input[2240:2247] = '{32'hc2c0530f, 32'hc22df892, 32'h42b4f1b3, 32'hbf9646f1, 32'hc268c345, 32'hc184b59b, 32'hc120b31e, 32'hc193e44e};
test_weights[2240:2247] = '{32'h42706106, 32'h4241bab6, 32'hc1623557, 32'hc1fde77e, 32'hc263a914, 32'h42918b45, 32'h40fe225f, 32'hc26378ce};
test_bias[280:280] = '{32'hc1d80fa6};
test_output[280:280] = '{32'hc5bdef08};
test_input[2248:2255] = '{32'hbf7dcf1d, 32'h42275489, 32'h4125bb21, 32'h42a484ba, 32'hc29e64c4, 32'hc03b5e8b, 32'hc28574e4, 32'h42a267ef};
test_weights[2248:2255] = '{32'hc18a45c8, 32'h42a2c96d, 32'hc2777b14, 32'h42b6b021, 32'hc1c5e871, 32'hc0c96ffc, 32'h41bdc60a, 32'hc0e977ed};
test_bias[281:281] = '{32'h42ab643c};
test_output[281:281] = '{32'h461f1c22};
test_input[2256:2263] = '{32'h42786165, 32'hc24b1365, 32'hc1d84df4, 32'h4265ba10, 32'hc22c85ad, 32'hbfbcbaf4, 32'h4299c375, 32'hc257df04};
test_weights[2256:2263] = '{32'hc26a4d43, 32'h41b8e945, 32'h42ab1473, 32'hc2007c90, 32'h41872245, 32'hc2bc8fc5, 32'h42c7fcb6, 32'hc11e8b09};
test_bias[282:282] = '{32'h41ba074a};
test_output[282:282] = '{32'hc4a40617};
test_input[2264:2271] = '{32'h429ba947, 32'hc0d7e7d9, 32'hc286fce4, 32'h4237b9d4, 32'h4253d485, 32'hc24b5e24, 32'hc28a877a, 32'hc1a4003f};
test_weights[2264:2271] = '{32'hc28b74c6, 32'hc2c5a0a4, 32'h42c12375, 32'h41a729af, 32'hc151d1c3, 32'h429d0271, 32'h4295a15c, 32'hc1a51063};
test_bias[283:283] = '{32'h41c9b9ac};
test_output[283:283] = '{32'hc69a3407};
test_input[2272:2279] = '{32'h424adcc5, 32'h427e0516, 32'hc2b9d410, 32'h42bba497, 32'h41c988c9, 32'h42b6f987, 32'hc1a7fdcd, 32'h42b7142c};
test_weights[2272:2279] = '{32'hc21a473d, 32'hc29dc8e1, 32'h420b9d95, 32'h42b330f7, 32'h42a3f4ce, 32'h41e40020, 32'hc29ecab6, 32'hc2a9cc61};
test_bias[284:284] = '{32'hc2448cc5};
test_output[284:284] = '{32'hc54d42a1};
test_input[2280:2287] = '{32'h419b98d1, 32'h42131659, 32'hc2ad094a, 32'hc28818d6, 32'hc231e49b, 32'h422b466a, 32'h4288e575, 32'hc1876a30};
test_weights[2280:2287] = '{32'h42828cd9, 32'hc28c1521, 32'h4143f06b, 32'hc2be5977, 32'h41cf29ca, 32'h422353b2, 32'h4285a7ea, 32'hc2746170};
test_bias[285:285] = '{32'hc1dbf671};
test_output[285:285] = '{32'h4620c282};
test_input[2288:2295] = '{32'hc2429ae3, 32'h42b937ef, 32'h409aa74d, 32'hc2acb7bb, 32'h41a5b9e5, 32'hbf0097ca, 32'hc2b0c94c, 32'hc2918775};
test_weights[2288:2295] = '{32'hc0cbb96a, 32'h42074fa5, 32'h415e6666, 32'h42bebf5e, 32'hc2b4f020, 32'hc2aee8f1, 32'h429568ae, 32'hc2477ee5};
test_bias[286:286] = '{32'h42709588};
test_output[286:286] = '{32'hc613fc3d};
test_input[2296:2303] = '{32'hc1c04ec3, 32'hc29d7ff4, 32'hc0c34fe5, 32'hc288243b, 32'hc283d9f3, 32'hc1f241e2, 32'hc272aeeb, 32'hc1b43cda};
test_weights[2296:2303] = '{32'h42b06afe, 32'h4204e76b, 32'h42a30934, 32'h4236e85e, 32'h42b0d36b, 32'h427facbe, 32'h4277cf6e, 32'hc2b20a34};
test_bias[287:287] = '{32'hc2b4e414};
test_output[287:287] = '{32'hc68c4604};
test_input[2304:2311] = '{32'hc2ac6e87, 32'h4089030c, 32'h42951d5f, 32'hbff1d8e1, 32'hc2a2c51a, 32'hc237d07d, 32'h420ff1a4, 32'h42210469};
test_weights[2304:2311] = '{32'h42240eed, 32'hc1c536a8, 32'h41ea5f2f, 32'hc2adca10, 32'hc082759c, 32'h429691e4, 32'hc2bc8a66, 32'hc29d3c97};
test_bias[288:288] = '{32'h424e404b};
test_output[288:288] = '{32'hc62aba66};
test_input[2312:2319] = '{32'h42b183c3, 32'h41c92a32, 32'h42aaf17b, 32'h429b5492, 32'hc1479850, 32'h4208e39c, 32'hc25f788b, 32'h41c42709};
test_weights[2312:2319] = '{32'hc2c5046d, 32'hc1d5fb97, 32'hc246c581, 32'hc1c8ad4d, 32'hc1ea78f5, 32'h419ecbbc, 32'hc291bac9, 32'h427f6ad9};
test_bias[289:289] = '{32'h420c1b79};
test_output[289:289] = '{32'hc60afc6f};
test_input[2320:2327] = '{32'h41e46d84, 32'hc2bb7916, 32'hc21ee61f, 32'h4259ea71, 32'hc2658110, 32'h42304d8f, 32'h424173f9, 32'h42c41e62};
test_weights[2320:2327] = '{32'hc281fb34, 32'h41b3d875, 32'h4193350d, 32'h4282d4a4, 32'hc1f1e73e, 32'h421174b6, 32'hc2483aa1, 32'h42c1a429};
test_bias[290:290] = '{32'hc28aae1b};
test_output[290:290] = '{32'h460feda7};
test_input[2328:2335] = '{32'h4269af87, 32'h4116afa6, 32'h41ea880f, 32'h42442b8f, 32'hc26be7fd, 32'hc2270f1b, 32'hc2762e45, 32'h42592df7};
test_weights[2328:2335] = '{32'hc23c7f49, 32'h42c2354c, 32'h421346d3, 32'h4197d0be, 32'hc156f620, 32'h42b34ce7, 32'hc2672f0b, 32'h42803ea1};
test_bias[291:291] = '{32'h42195f18};
test_output[291:291] = '{32'h458644b0};
test_input[2336:2343] = '{32'h4011bb94, 32'h42b0b12d, 32'hc2bdf374, 32'h41a6747d, 32'h423145e8, 32'hc1e21565, 32'h42980fdb, 32'hc09dccda};
test_weights[2336:2343] = '{32'hc02f2380, 32'hc286c4f6, 32'h42494a6c, 32'h417aeff9, 32'h41d97dde, 32'h42bc7e1e, 32'h427bd841, 32'h42582617};
test_bias[292:292] = '{32'hc13487fa};
test_output[292:292] = '{32'hc5e60eb4};
test_input[2344:2351] = '{32'h427a8cda, 32'h42be1776, 32'hc2c169b5, 32'hc272ba9e, 32'h4281074a, 32'hc2ac1c61, 32'hc2977a5a, 32'h41e820bc};
test_weights[2344:2351] = '{32'hc252e43f, 32'hc08e563b, 32'hc21d4789, 32'h428c3731, 32'h40859c2f, 32'hc10e4020, 32'hc0da58b1, 32'hc21a700e};
test_bias[293:293] = '{32'h4128d919};
test_output[293:293] = '{32'hc569780b};
test_input[2352:2359] = '{32'hc1c59d57, 32'hc29219ec, 32'h413c87d3, 32'hc25b1f87, 32'h42593623, 32'hc23d55a4, 32'hc1ab3887, 32'hc23c1c54};
test_weights[2352:2359] = '{32'h42852916, 32'hc239378e, 32'h41a7ba7a, 32'hc261aa5a, 32'h42b2beca, 32'h4139a159, 32'h408ab0a4, 32'hc2912f56};
test_bias[294:294] = '{32'h423a723f};
test_output[294:294] = '{32'h46472cdd};
test_input[2360:2367] = '{32'h42c74f04, 32'hc2c261d6, 32'hc2b0700c, 32'hc20155a1, 32'hc1c39adc, 32'hc1e97279, 32'hc2ad47f6, 32'hc04d9ecc};
test_weights[2360:2367] = '{32'h42a58a44, 32'h42c1f4af, 32'h42a401ab, 32'h42a5509f, 32'h4274300b, 32'hc244b1dd, 32'h4226438f, 32'h42a14883};
test_bias[295:295] = '{32'hc29732e6};
test_output[295:295] = '{32'hc66b961d};
test_input[2368:2375] = '{32'hc12b9b0e, 32'h41c22b29, 32'hc233d465, 32'hc1a9f77c, 32'h405f7fef, 32'hc0bf0508, 32'h4293b306, 32'h42505fda};
test_weights[2368:2375] = '{32'hc24d70dc, 32'hc2b644f6, 32'hc1a38d73, 32'hc27c079e, 32'h4200195d, 32'h4113fb81, 32'h40cc9e16, 32'hc1fbb15d};
test_bias[296:296] = '{32'h4289835a};
test_output[296:296] = '{32'hc3de55d6};
test_input[2376:2383] = '{32'h421ec785, 32'hbee0275f, 32'hc28322c9, 32'h41699aab, 32'hc2bfd66e, 32'h422dcd29, 32'h429e6e64, 32'hc29be667};
test_weights[2376:2383] = '{32'hc213a69e, 32'h41e12b2a, 32'h42a1024b, 32'h41043923, 32'hc292aa15, 32'h42adb5c6, 32'h4091b4b2, 32'h42840ab5};
test_bias[297:297] = '{32'hc28c483d};
test_output[297:297] = '{32'hc42ad89b};
test_input[2384:2391] = '{32'h41c2943e, 32'h42949d39, 32'h42c55649, 32'h4292088f, 32'h42b82638, 32'hc0ebc6a8, 32'h41bd7bbc, 32'hc2ba6557};
test_weights[2384:2391] = '{32'h42b32f11, 32'h4165ec40, 32'hc28304fe, 32'hc126412f, 32'hc25b7ec7, 32'h421211f4, 32'hc2ac20e5, 32'hc2399465};
test_bias[298:298] = '{32'h4251e7b3};
test_output[298:298] = '{32'hc5d9798f};
test_input[2392:2399] = '{32'hc2c6a3f7, 32'h4072a311, 32'hc2763037, 32'hc29f2722, 32'h4210b158, 32'h41795651, 32'h42391721, 32'h41cf42af};
test_weights[2392:2399] = '{32'hc2bf2a8c, 32'h426d3cf3, 32'hc2c2fcdd, 32'h4285418e, 32'hc07b37ae, 32'h42a08d29, 32'h42576a3f, 32'h4084e938};
test_bias[299:299] = '{32'h401ce90c};
test_output[299:299] = '{32'h465cbe8c};
test_input[2400:2407] = '{32'h4281a630, 32'hc0a59079, 32'h4244a193, 32'hc262acfc, 32'h4281c778, 32'hc1fbfaed, 32'hc2a9be19, 32'hc23d6ce1};
test_weights[2400:2407] = '{32'h428aead0, 32'hc1b58bb5, 32'h42829efa, 32'hc23bf937, 32'h41c7ff5d, 32'hc2c13317, 32'hc1e73401, 32'h420bccaa};
test_bias[300:300] = '{32'hc2a9f1db};
test_output[300:300] = '{32'h4677fcf5};
test_input[2408:2415] = '{32'h424b6e6a, 32'hc12a312e, 32'h419c1fb5, 32'h4290ccaa, 32'hc198655c, 32'h423403ed, 32'hc1e50a71, 32'h429ef87e};
test_weights[2408:2415] = '{32'h4211e94d, 32'h41a0e7d1, 32'h41a981e8, 32'hc2c17548, 32'hc12251cc, 32'h41483367, 32'hc24b6976, 32'h42092771};
test_bias[301:301] = '{32'h41e48d34};
test_output[301:301] = '{32'h418f0e15};
test_input[2416:2423] = '{32'h42281226, 32'h4196ef99, 32'h426c7ed2, 32'h427a1ca9, 32'hc25dbf28, 32'hc29a63b1, 32'h4283693f, 32'hc29a050c};
test_weights[2416:2423] = '{32'hc2568140, 32'h42ae2a37, 32'h4170018c, 32'hc286691e, 32'hc2758c7d, 32'h42c67719, 32'h42af7ae8, 32'h3f9bbaf8};
test_bias[302:302] = '{32'h3c34422b};
test_output[302:302] = '{32'hc51cf675};
test_input[2424:2431] = '{32'h427b42d3, 32'h424e212f, 32'h41361091, 32'h3fe69c78, 32'h4203b268, 32'h425d1c75, 32'hc2a7f6ff, 32'h4190b586};
test_weights[2424:2431] = '{32'hc2bb2a85, 32'hc1b5e993, 32'h4285be05, 32'h42154ad7, 32'hc2879d15, 32'hc1d108e4, 32'hc0b2ddc1, 32'hc1c617a3};
test_bias[303:303] = '{32'hc26a7cd5};
test_output[303:303] = '{32'hc61b401b};
test_input[2432:2439] = '{32'h4292ce6e, 32'hc272da22, 32'hc2ab83c2, 32'hc2bc4d8f, 32'hc20490a5, 32'h40b0557b, 32'h4157ac57, 32'h42423e2e};
test_weights[2432:2439] = '{32'h42acfcdd, 32'h41c2c43c, 32'h42a11281, 32'h426ba736, 32'h41f9e582, 32'hc2732daf, 32'hc1eba27f, 32'h4292840d};
test_bias[304:304] = '{32'h42018940};
test_output[304:304] = '{32'hc5b3ff9e};
test_input[2440:2447] = '{32'h41ffa9b6, 32'h41eb72d3, 32'h420fd827, 32'hc226ec18, 32'hc070e13f, 32'hc2158e80, 32'hc0aa8ef8, 32'hc1faea01};
test_weights[2440:2447] = '{32'h425a5b82, 32'hc1ded4e5, 32'h42b7bf9d, 32'h4289f13a, 32'h4267bf4b, 32'h415d7e7f, 32'h420272f5, 32'h41bfa829};
test_bias[305:305] = '{32'hc2b5549b};
test_output[305:305] = '{32'hc3c8870f};
test_input[2448:2455] = '{32'hc1aa6eac, 32'hc2b95f31, 32'hc0ad56b3, 32'hc29dc6c1, 32'h4296437c, 32'hc2ba3517, 32'h42821c30, 32'h41489a69};
test_weights[2448:2455] = '{32'h3e3cda0b, 32'h4218997a, 32'h41d0e87c, 32'hc2203f8d, 32'h41a0744e, 32'hc2577e6e, 32'hc28cd8ed, 32'hc2a83d0c};
test_bias[306:306] = '{32'hbc85116b};
test_output[306:306] = '{32'h43b6db22};
test_input[2456:2463] = '{32'hc2449021, 32'h4218abbe, 32'h42ad324d, 32'h429b981d, 32'h4184ee70, 32'h428c51f2, 32'h421e4781, 32'h428dd950};
test_weights[2456:2463] = '{32'h423f1b53, 32'h42848ad6, 32'h41881034, 32'hc2b4cc74, 32'hc27dec6d, 32'hc2369736, 32'hc2968016, 32'h42203637};
test_bias[307:307] = '{32'hc2837a21};
test_output[307:307] = '{32'hc619b9b1};
test_input[2464:2471] = '{32'h423b679e, 32'hc2a1f61e, 32'h4284498b, 32'h420e5130, 32'hc20fec17, 32'hc0c49255, 32'hc26edd00, 32'hc2c7edb2};
test_weights[2464:2471] = '{32'h429064b0, 32'h42520c65, 32'hc2a28577, 32'h4156a55f, 32'h425fec18, 32'h42889f3b, 32'h42b0f43d, 32'hc25f6621};
test_bias[308:308] = '{32'hc2b7a107};
test_output[308:308] = '{32'hc5f9cd81};
test_input[2472:2479] = '{32'hc2bd55f5, 32'hc188dc1f, 32'h429d3f86, 32'h426ea5ea, 32'hc2c72bbf, 32'h42b0c797, 32'hc1f7ee1c, 32'h41b2c03b};
test_weights[2472:2479] = '{32'h421590bd, 32'hc158b2ad, 32'h42b78886, 32'h42506565, 32'hc2a80c63, 32'hc1fb571e, 32'h42c72881, 32'h42b8e6c9};
test_bias[309:309] = '{32'h40d04d27};
test_output[309:309] = '{32'h46352045};
test_input[2480:2487] = '{32'hc2965f4f, 32'h427b7687, 32'hc2a847c9, 32'h4266d390, 32'hc1d220c7, 32'h4167c17d, 32'hc0ef3b4b, 32'h40bd6eec};
test_weights[2480:2487] = '{32'hc25e745f, 32'hc26beb0c, 32'h42a754fd, 32'h428290a1, 32'h42a1be24, 32'hc2098617, 32'h42c00b44, 32'h42b6d16e};
test_bias[310:310] = '{32'h426ea831};
test_output[310:310] = '{32'hc5ad10cd};
test_input[2488:2495] = '{32'hc1e1659a, 32'hc29dec4b, 32'h41bd3e5d, 32'hc29fe4c4, 32'hc2b041b7, 32'h42b7b658, 32'h42b0fe0c, 32'h423e3cb3};
test_weights[2488:2495] = '{32'hc281472b, 32'hc1afef7d, 32'hc274fede, 32'h420dd424, 32'hc205a325, 32'hc29ad331, 32'h42afcbcb, 32'h4261bd8d};
test_bias[311:311] = '{32'h428b82e6};
test_output[311:311] = '{32'h45b04058};
test_input[2496:2503] = '{32'h4144250d, 32'h421975a0, 32'hbe82364d, 32'hc21e8b8d, 32'hc263d86c, 32'h413f128d, 32'hc2534225, 32'hbfcd1b11};
test_weights[2496:2503] = '{32'hc235afef, 32'hc2031db1, 32'h4270b45b, 32'hbf67d7dd, 32'h42087090, 32'h42bb45c6, 32'hc13757e8, 32'hc1b2ff55};
test_bias[312:312] = '{32'h420901a7};
test_output[312:312] = '{32'hc4f2e775};
test_input[2504:2511] = '{32'hc2036689, 32'h4243b880, 32'hc1c206c5, 32'h41bcfbc6, 32'h425e491d, 32'hc2baf356, 32'h4212501d, 32'h42b2ca6b};
test_weights[2504:2511] = '{32'h423b5aec, 32'hc2388222, 32'h422b8602, 32'h422bf332, 32'h4243e84e, 32'hc2983bef, 32'h41c10b96, 32'h42824556};
test_bias[313:313] = '{32'hc0df4d55};
test_output[313:313] = '{32'h4646ac51};
test_input[2512:2519] = '{32'h429c2680, 32'hc2b56a8e, 32'hc20effeb, 32'h428e4ff8, 32'h4287edbd, 32'h422e1198, 32'h4183c48e, 32'hc2ad398a};
test_weights[2512:2519] = '{32'hc2616b98, 32'h42b13868, 32'h422286b6, 32'h41abd968, 32'hc20140d5, 32'h4243df12, 32'hc20872da, 32'h3fb99fe5};
test_bias[314:314] = '{32'h4222c2ef};
test_output[314:314] = '{32'hc64c468d};
test_input[2520:2527] = '{32'hc2b64381, 32'h42764b63, 32'h422209d6, 32'h42c6e3b1, 32'h4282faf8, 32'h42333c78, 32'hc18e5f89, 32'h422647f1};
test_weights[2520:2527] = '{32'hc2a2646a, 32'h4287a63b, 32'h4258511a, 32'h4238f871, 32'h42a7ab28, 32'hc299facd, 32'h42b2a4cc, 32'hc2abf119};
test_bias[315:315] = '{32'h41cf2047};
test_output[315:315] = '{32'h466e8fee};
test_input[2528:2535] = '{32'h42087316, 32'h41fa0019, 32'h42865794, 32'hc2474448, 32'hc28c9f33, 32'h41bbcaba, 32'h42b2aaf8, 32'h41f80ba6};
test_weights[2528:2535] = '{32'hc294434e, 32'hc2c7c926, 32'hc20902d0, 32'hc1bb5cb9, 32'h42a469fb, 32'h42330407, 32'hc2c74d48, 32'h40c3eb95};
test_bias[316:316] = '{32'hc226e44d};
test_output[316:316] = '{32'hc69e5842};
test_input[2536:2543] = '{32'hc29a1e34, 32'h4295413c, 32'hc259752d, 32'hc22520d7, 32'h41c1f27b, 32'h423c4876, 32'hc21c8fb3, 32'hc2445d8e};
test_weights[2536:2543] = '{32'hc2978253, 32'hc1646a7b, 32'hc2833f74, 32'h427b1b4e, 32'h428b1f4e, 32'hc28a8739, 32'hc254df1c, 32'hc2b30b9d};
test_bias[317:317] = '{32'h424c79d8};
test_output[317:317] = '{32'h46273cd1};
test_input[2544:2551] = '{32'hc29c887a, 32'h40b570e4, 32'h40157d4b, 32'h42841f5f, 32'h42ba9cdd, 32'h42b4c727, 32'h42124f13, 32'hc0347592};
test_weights[2544:2551] = '{32'h41bd5799, 32'h42c5245d, 32'h42480f6b, 32'hc2a8e434, 32'h41f7300f, 32'h42756fc9, 32'h42c45063, 32'h41a6513e};
test_bias[318:318] = '{32'hc28bc594};
test_output[318:318] = '{32'h45a07e12};
test_input[2552:2559] = '{32'h42c572a7, 32'hc25d8bc9, 32'hc27fed6c, 32'h41476490, 32'h4154d051, 32'hc2b101fe, 32'hc1fdf8ce, 32'h4216748d};
test_weights[2552:2559] = '{32'h41d35a4b, 32'hc0a2fe92, 32'hc19a7055, 32'hc1b7b331, 32'h42bde3af, 32'hc156e99a, 32'hc1a48d07, 32'hc2858026};
test_bias[319:319] = '{32'hc26ec110};
test_output[319:319] = '{32'h4588ac19};
test_input[2560:2567] = '{32'hc2b4ce04, 32'hc11a6f93, 32'hc289a754, 32'hc28f08cc, 32'hc1cb2d13, 32'h419cdbda, 32'hc185e4c8, 32'h4234cf99};
test_weights[2560:2567] = '{32'hc2c4410e, 32'hc2b93013, 32'hc2a96dc3, 32'hc29b9cda, 32'h425f2c7a, 32'h429857fd, 32'h418f0bb9, 32'hc0b345cd};
test_bias[320:320] = '{32'hc18c9a63};
test_output[320:320] = '{32'h46a17477};
test_input[2568:2575] = '{32'hc2c2b82c, 32'hc2a6dd49, 32'hc204223e, 32'hc2a3e078, 32'h42abe591, 32'h4059a2c5, 32'hc1bba8e3, 32'hc24a973a};
test_weights[2568:2575] = '{32'hc2a8b70f, 32'hc29622c9, 32'hc0e80ded, 32'hc1d8fc56, 32'h42a16c27, 32'hc2a05f70, 32'h42aeebb9, 32'hc2ae12bb};
test_bias[321:321] = '{32'hc10fb499};
test_output[321:321] = '{32'h46cabc10};
test_input[2576:2583] = '{32'h40e8f43e, 32'hc2b97ea1, 32'h424fbf3d, 32'hc2a8c792, 32'hc1934cce, 32'h4229948e, 32'h422bff55, 32'hc22907da};
test_weights[2576:2583] = '{32'hc129ddac, 32'hc163f1e6, 32'h42952a93, 32'h42095d97, 32'h40523bf9, 32'hc1b78eec, 32'hc2bdc3b8, 32'h42bbc9cb};
test_bias[322:322] = '{32'hc21be03f};
test_output[322:322] = '{32'hc5d7a1de};
test_input[2584:2591] = '{32'h40a6185b, 32'hc2bd3a76, 32'h41fbcbeb, 32'hc1f82c0c, 32'h429ec666, 32'h4271eb8d, 32'hc1e0e0b2, 32'hc1ec9994};
test_weights[2584:2591] = '{32'h4141aeba, 32'hc2a0a392, 32'hc20f215d, 32'hc208663e, 32'h4188f2ba, 32'hc222f007, 32'hc22389e5, 32'h41139d77};
test_bias[323:323] = '{32'h41850f8c};
test_output[323:323] = '{32'h45e6b186};
test_input[2592:2599] = '{32'hc150b148, 32'hbf87856a, 32'hc1898f1d, 32'hc2c127e7, 32'h42a282d9, 32'h42264bad, 32'h41ad5a52, 32'hc2723aa6};
test_weights[2592:2599] = '{32'hc22dc545, 32'h4297eea6, 32'hc2bd9419, 32'hc17cd5a6, 32'hc227592e, 32'hc08e6afe, 32'hc10f185b, 32'hc2104edc};
test_bias[324:324] = '{32'hc2951077};
test_output[324:324] = '{32'h44f6c376};
test_input[2600:2607] = '{32'hc211a9d5, 32'hc121f672, 32'hc1ecf7ab, 32'hc29a4224, 32'hc0bb0a19, 32'hc254ca60, 32'h41ed78ca, 32'hc2c2afba};
test_weights[2600:2607] = '{32'hc195e05d, 32'h42ac7eb1, 32'hc26a7a24, 32'hc0c29ab3, 32'hc1c65868, 32'h42a81055, 32'h428ccb64, 32'h4262932e};
test_bias[325:325] = '{32'h41a1635e};
test_output[325:325] = '{32'hc5b296a6};
test_input[2608:2615] = '{32'h41e969b2, 32'h428dd083, 32'h40266a45, 32'hc281343d, 32'hc2b88d76, 32'hc2c0b359, 32'h4299d298, 32'hc04b2828};
test_weights[2608:2615] = '{32'hc1ba9d4e, 32'hc2942f70, 32'h4291b65f, 32'h42191817, 32'hc254894e, 32'hc2a7e03a, 32'hc2a952ec, 32'hc27c1afb};
test_bias[326:326] = '{32'h421a4605};
test_output[326:326] = '{32'hc4bb78c5};
test_input[2616:2623] = '{32'h423d1eec, 32'h4038e748, 32'h41d3ae5e, 32'hc28f67b5, 32'hc2a58304, 32'hc289f302, 32'hc2825298, 32'h40f89c48};
test_weights[2616:2623] = '{32'hc1843600, 32'hc1963356, 32'hc1ef5bd9, 32'hc27dd64e, 32'hc2b4da5c, 32'h42b016d2, 32'h42312763, 32'h42208047};
test_bias[327:327] = '{32'hc1b4ed96};
test_output[327:327] = '{32'h44d91358};
test_input[2624:2631] = '{32'h41afe673, 32'hc2a430ac, 32'hc1b22084, 32'hc20ae161, 32'hc2806910, 32'h42bd4379, 32'h42855788, 32'h4267c1b8};
test_weights[2624:2631] = '{32'hc2007cc5, 32'h417cde06, 32'hc2699772, 32'hc24a7ce1, 32'h426ac8d6, 32'h42bf0b3b, 32'h42ae0529, 32'hc2a2e0e5};
test_bias[328:328] = '{32'h41685084};
test_output[328:328] = '{32'h45e7f013};
test_input[2632:2639] = '{32'h41c1375b, 32'h42c2493b, 32'hc1b71b96, 32'hc1b2d95a, 32'h42a0bbb2, 32'h4294611e, 32'h42a1bf50, 32'h411d4502};
test_weights[2632:2639] = '{32'hc234142e, 32'h41d5fda8, 32'hc0e8c9cd, 32'hc2ae4983, 32'h4240f12e, 32'h42a8bf93, 32'h428226e0, 32'hc2bc9d08};
test_bias[329:329] = '{32'hc20a222d};
test_output[329:329] = '{32'h468d1ef8};
test_input[2640:2647] = '{32'h42535a0e, 32'hc2855057, 32'hc2afce6a, 32'hc22a016b, 32'hc2a74346, 32'h41e528d8, 32'h4142fe25, 32'h42b872c9};
test_weights[2640:2647] = '{32'h4226fa8b, 32'h4263e68b, 32'h428b5608, 32'h4214c14f, 32'h42c27972, 32'hc21f674e, 32'h42a40fff, 32'hc29e09e5};
test_bias[330:330] = '{32'hc28d128c};
test_output[330:330] = '{32'hc6c2c13c};
test_input[2648:2655] = '{32'h428fed06, 32'hc155ffdd, 32'hc28ff3e2, 32'h4224aa92, 32'hc28b74db, 32'hc2460f9e, 32'h4169cb5d, 32'hc2907035};
test_weights[2648:2655] = '{32'h424a8d9c, 32'hbfc58fe9, 32'hc21c8a58, 32'hc1f89ae0, 32'hc1f7feb2, 32'h417b4a81, 32'hc2bea469, 32'hc1777767};
test_bias[331:331] = '{32'hc1d3d87a};
test_output[331:331] = '{32'h45c45e27};
test_input[2656:2663] = '{32'h42c53f5d, 32'hc1f83878, 32'h429d0a55, 32'hc2831356, 32'hc0cc68d1, 32'hc2aab457, 32'h420c95a1, 32'h41e755b4};
test_weights[2656:2663] = '{32'h428c4db9, 32'h41ab4e07, 32'h41cbecc9, 32'hc04d488e, 32'h42c6155b, 32'h42a338c6, 32'hc280fba5, 32'hc29499e4};
test_bias[332:332] = '{32'hc2817c60};
test_output[332:332] = '{32'hc561c411};
test_input[2664:2671] = '{32'hc1bb0846, 32'hc2861b80, 32'h42949ce9, 32'h42a8af8b, 32'h41f63600, 32'h422eb544, 32'hc1899c13, 32'hc2721b67};
test_weights[2664:2671] = '{32'h420d39c4, 32'hc2b43b52, 32'hc28c2777, 32'hc1fa53cd, 32'h4081db8a, 32'h42c36753, 32'h4269f2f5, 32'hc13664f7};
test_bias[333:333] = '{32'h425b8b5c};
test_output[333:333] = '{32'h44bbbb92};
test_input[2672:2679] = '{32'h428b9306, 32'h41b10669, 32'h428c4997, 32'h41cbab5d, 32'hc25462d1, 32'hc2968f50, 32'h421dc0d8, 32'hc1e541e2};
test_weights[2672:2679] = '{32'hc183f83e, 32'h41833464, 32'hc2112b77, 32'h41be2dcf, 32'hc21f3339, 32'h4092e73a, 32'hc19e8569, 32'hc23fb1a2};
test_bias[334:334] = '{32'h424c77c0};
test_output[334:334] = '{32'hc39f11e2};
test_input[2680:2687] = '{32'hc241d582, 32'h42840cc6, 32'h420abac8, 32'h4234d5a8, 32'h42917be5, 32'h425ab918, 32'h424c3960, 32'hc24388ed};
test_weights[2680:2687] = '{32'hc23890d8, 32'hbf0e6529, 32'h42bc835c, 32'hc230e522, 32'hc2a2d0e3, 32'hc2c33e45, 32'h42716113, 32'h428cfe25};
test_bias[335:335] = '{32'hc2c0f4c9};
test_output[335:335] = '{32'hc600f1e2};
test_input[2688:2695] = '{32'hc23301f6, 32'hc274d75c, 32'h4290b775, 32'h42398a37, 32'hc1b0a563, 32'hc1ade2e0, 32'h428ea5d6, 32'hc2bab507};
test_weights[2688:2695] = '{32'hc2871533, 32'h401fe811, 32'hc2ada426, 32'h424b1f01, 32'hc2064282, 32'hc27e57a2, 32'h41b300cb, 32'h421d8c0d};
test_bias[336:336] = '{32'h409263bc};
test_output[336:336] = '{32'hc47c91dc};
test_input[2696:2703] = '{32'h428e9e9b, 32'hc216693c, 32'h420765da, 32'h42c7646e, 32'h42a6adac, 32'h420afb57, 32'hc2925785, 32'hc20be5b6};
test_weights[2696:2703] = '{32'h4270345b, 32'hc2bdad3f, 32'hc299e695, 32'hc2c0a0b6, 32'hc0f3f353, 32'hc273ce1b, 32'hc2ab5be8, 32'h42a88792};
test_bias[337:337] = '{32'hc1e4dacf};
test_output[337:337] = '{32'hc56ea021};
test_input[2704:2711] = '{32'h42b5c728, 32'hc10e624b, 32'h425881e7, 32'hc0422c2e, 32'hc0a1e83d, 32'h429ca2f1, 32'hc206cdab, 32'hc1e8ffaa};
test_weights[2704:2711] = '{32'h42b0ba0a, 32'h42a0ceea, 32'hc234488a, 32'hc2a260d5, 32'h424c1a19, 32'h429772cd, 32'hc2c70db2, 32'h4219efce};
test_bias[338:338] = '{32'h41b3d259};
test_output[338:338] = '{32'h464bead4};
test_input[2712:2719] = '{32'hc04237eb, 32'h42afd21a, 32'hc2c535cb, 32'h42a6103f, 32'h42121e8c, 32'hc191f26d, 32'h424fd48a, 32'h3e97b9ed};
test_weights[2712:2719] = '{32'hc274df53, 32'hc2bcb92d, 32'h4219e285, 32'h4236a6bb, 32'hc1054d7a, 32'hc2b3d353, 32'h41949b1b, 32'hc200a73a};
test_bias[339:339] = '{32'hc2915f07};
test_output[339:339] = '{32'hc5b8257c};
test_input[2720:2727] = '{32'h429357f5, 32'h4217bde9, 32'hc151f838, 32'h42b1d791, 32'h4261577c, 32'hc2a62ec4, 32'h429eaae1, 32'hc21db4ae};
test_weights[2720:2727] = '{32'hc2ab4406, 32'hc2c7bd02, 32'h4234129b, 32'hc1d0fd65, 32'h423f983d, 32'h421de0a1, 32'h4167443c, 32'h42799dfa};
test_bias[340:340] = '{32'h42c21fd7};
test_output[340:340] = '{32'hc6676346};
test_input[2728:2735] = '{32'h424c44cf, 32'hc28de62c, 32'h429e124b, 32'hc1980e92, 32'hc28b9eef, 32'h421262d7, 32'h42b6b5bb, 32'h425f66e7};
test_weights[2728:2735] = '{32'hc28a8448, 32'hc29d3fef, 32'h428e9e1e, 32'h41a58940, 32'h41e9d8a0, 32'hc195520f, 32'hc2a25083, 32'hc27a8728};
test_bias[341:341] = '{32'hc252b5be};
test_output[341:341] = '{32'hc5c82256};
test_input[2736:2743] = '{32'hc20fe41e, 32'h42304b0a, 32'hc2bb6a46, 32'hc0977f31, 32'hc2a3e39a, 32'hc23ff9a5, 32'h42a32ddc, 32'hc1c70acd};
test_weights[2736:2743] = '{32'h4280ca03, 32'h42038857, 32'h42c1722d, 32'h422fd5fc, 32'hc2784829, 32'h42560ca5, 32'h4103e512, 32'h424c725b};
test_bias[342:342] = '{32'hc1bca590};
test_output[342:342] = '{32'hc600ce4c};
test_input[2744:2751] = '{32'h42bc8797, 32'h425eb0f2, 32'h4245db5e, 32'hc27111ea, 32'h428f0882, 32'h4211f486, 32'h41c23c9f, 32'hc199acea};
test_weights[2744:2751] = '{32'h42a38357, 32'hc23b73fc, 32'hc2713a64, 32'hc193d3f0, 32'h40f44b73, 32'h42099bdc, 32'hc25a9217, 32'hc20c5b0d};
test_bias[343:343] = '{32'hc23495bf};
test_output[343:343] = '{32'h45875e98};
test_input[2752:2759] = '{32'h425b21f6, 32'h429365b6, 32'h424857ba, 32'h425c1658, 32'hc2c4724a, 32'h41be133d, 32'h4232511a, 32'hc22f88af};
test_weights[2752:2759] = '{32'h421db6a3, 32'hc1258866, 32'h42b6d227, 32'h41802f8f, 32'hc1e1bc24, 32'hc2be6ada, 32'h4120e765, 32'h41cd42a9};
test_bias[344:344] = '{32'h424f1ed3};
test_output[344:344] = '{32'h45d2a8f1};
test_input[2760:2767] = '{32'hc2b3aaa2, 32'h4297d29c, 32'h41c44eae, 32'hc20d7a4e, 32'h426581e3, 32'hc2384b30, 32'h42b18d82, 32'hc03f2305};
test_weights[2760:2767] = '{32'hc1e57400, 32'h4296f8cb, 32'hc1d3afff, 32'hc27b8bc0, 32'h429b023f, 32'hc29cd4f3, 32'h420ba591, 32'h42994725};
test_bias[345:345] = '{32'hc20686d5};
test_output[345:345] = '{32'h46a254d6};
test_input[2768:2775] = '{32'hc2a9c3b8, 32'hc2961c26, 32'hc2a218fe, 32'h421e7b41, 32'h42c45df1, 32'hc2074915, 32'h422b0dc5, 32'hc0b0eb7f};
test_weights[2768:2775] = '{32'hc2552c63, 32'h42009026, 32'hc2ab6ff9, 32'h41f5a937, 32'hc2b99126, 32'h424c731c, 32'h40ec3e67, 32'hc2a3b74a};
test_bias[346:346] = '{32'hc1b6052d};
test_output[346:346] = '{32'h4336685f};
test_input[2776:2783] = '{32'hc2ba675e, 32'h424ee5ea, 32'hc21f84cb, 32'h427dd90d, 32'hc2a6429e, 32'hc2b196dd, 32'hc23de356, 32'hc2a84a03};
test_weights[2776:2783] = '{32'h41eda70c, 32'hc23dcce5, 32'hc23ec721, 32'h42b3af3b, 32'hc27e4b71, 32'hc1eff6b6, 32'h420c558e, 32'h42716d54};
test_bias[347:347] = '{32'h41ffb262};
test_output[347:347] = '{32'h45620ab6};
test_input[2784:2791] = '{32'h416f7ce7, 32'h41c58be0, 32'hc1892593, 32'h429a7a0e, 32'h417642ce, 32'h42ace553, 32'h42763c5e, 32'h42bf5180};
test_weights[2784:2791] = '{32'hbffb3b44, 32'hc28b9caf, 32'hc1c6f339, 32'hc2a11c97, 32'h42ae63d2, 32'hc29098cf, 32'h4289c2e0, 32'hc29e6718};
test_bias[348:348] = '{32'hc2b9a741};
test_output[348:348] = '{32'hc67836f4};
test_input[2792:2799] = '{32'h42b3e020, 32'h42af1ba7, 32'hc28c3934, 32'hc159ac38, 32'h42150671, 32'hc235d427, 32'h420eefa4, 32'h41c74fe1};
test_weights[2792:2799] = '{32'h428994e3, 32'h41e311a6, 32'h4261b0dc, 32'hc1e99bcd, 32'h4283a8ec, 32'h426a982c, 32'hc22fe53f, 32'h428082e2};
test_bias[349:349] = '{32'hc150ee6b};
test_output[349:349] = '{32'h4599a313};
test_input[2800:2807] = '{32'hc2679dca, 32'hc29fe424, 32'hc20a6240, 32'hc24afbfa, 32'h429aa849, 32'h42a13409, 32'hc25e4fb2, 32'hc11bf861};
test_weights[2800:2807] = '{32'h418b2ac5, 32'hc1755aeb, 32'hc2bd2bc1, 32'hc2867a95, 32'h42a080cb, 32'hc252c1db, 32'hc26a4b46, 32'hc2546f20};
test_bias[350:350] = '{32'hc280c133};
test_output[350:350] = '{32'h46446ab9};
test_input[2808:2815] = '{32'h40b52a43, 32'hc2028379, 32'hc1fe5afe, 32'hc136bb84, 32'hc2ace47d, 32'h42aa5467, 32'hc27c2802, 32'h4253dbce};
test_weights[2808:2815] = '{32'hbfcc4cca, 32'hc208adb0, 32'h42b4ee54, 32'hc24f0168, 32'hc1f93508, 32'h42c13d85, 32'h41fe759f, 32'h41820266};
test_bias[351:351] = '{32'hc1ebc4f7};
test_output[351:351] = '{32'h4605e120};
test_input[2816:2823] = '{32'hc214f06e, 32'hc22051de, 32'h42821e83, 32'h429ef55c, 32'hc1f0ee6b, 32'hc2a72321, 32'h417e4d16, 32'hc1eab94b};
test_weights[2816:2823] = '{32'hc262a23c, 32'h4292574e, 32'hc28829c5, 32'h41f952b5, 32'h427711dc, 32'h42160938, 32'h428fb61f, 32'h412bc75d};
test_bias[352:352] = '{32'hc16a510c};
test_output[352:352] = '{32'hc5d96def};
test_input[2824:2831] = '{32'h423c49f7, 32'h41de3ea0, 32'hc298288e, 32'hc2c728b5, 32'h41b401d7, 32'h426859e5, 32'h42aa0675, 32'hc2c48f9f};
test_weights[2824:2831] = '{32'h42121263, 32'hc26019f3, 32'hc1834763, 32'h4198c593, 32'hc1e10426, 32'h429ae6a9, 32'hc2ac3bfd, 32'hc1b80681};
test_bias[353:353] = '{32'hc2877626};
test_output[353:353] = '{32'hc4db1239};
test_input[2832:2839] = '{32'hc15f696e, 32'h428d4c61, 32'hc10fb955, 32'h41b95c43, 32'hc2882d97, 32'h422c4aa9, 32'h41e7fb88, 32'hc2a38122};
test_weights[2832:2839] = '{32'hc29adf73, 32'hc190c869, 32'hc1ffdf37, 32'h42b518f0, 32'hc0bce6fa, 32'h41dce35b, 32'h42a9640d, 32'hc29b3531};
test_bias[354:354] = '{32'h420a9e46};
test_output[354:354] = '{32'h46451892};
test_input[2840:2847] = '{32'hc295cf11, 32'h42bbc6c2, 32'hc2223a1a, 32'h424fb2fe, 32'h425f709d, 32'h410f2f46, 32'hc2698c0b, 32'hc29c5dec};
test_weights[2840:2847] = '{32'hc2c68b88, 32'h40b57222, 32'hc1d8ab07, 32'hc20853d4, 32'h4299edc9, 32'hc2c4c26d, 32'hc108d8e1, 32'hc251638d};
test_bias[355:355] = '{32'h428a239d};
test_output[355:355] = '{32'h46704401};
test_input[2848:2855] = '{32'hc2c386eb, 32'hc1e4b017, 32'h42ae20e7, 32'h418ff736, 32'hc1816a2b, 32'h4282b968, 32'hc0e2ce7f, 32'hc2b04bde};
test_weights[2848:2855] = '{32'hc1c53677, 32'hc2c0ee82, 32'h41a59a73, 32'h42b064b7, 32'hc2a6af62, 32'h426da144, 32'h42be97ca, 32'h42ad5f38};
test_bias[356:356] = '{32'hc1bd77b2};
test_output[356:356] = '{32'h45aa3f54};
test_input[2856:2863] = '{32'h4287df10, 32'h41b834fe, 32'hc1a73cf9, 32'hc26689e5, 32'h4183ce72, 32'hc25d6be8, 32'hc132a6f3, 32'hc2c135fb};
test_weights[2856:2863] = '{32'hc01489b8, 32'h42b9e5e8, 32'hbf591ae2, 32'h4250cd1b, 32'hc1e71983, 32'h42399bbd, 32'hc152eea8, 32'h41d74354};
test_bias[357:357] = '{32'hc2b522ff};
test_output[357:357] = '{32'hc5ce1cf7};
test_input[2864:2871] = '{32'h40a46d4c, 32'h422f9825, 32'h427f18d7, 32'h42b09a6a, 32'hc261a84f, 32'hc220aa13, 32'h42740b01, 32'hc2873506};
test_weights[2864:2871] = '{32'h4090811c, 32'hc21c2dbc, 32'hc1007b13, 32'h42a00950, 32'hc25d93c9, 32'h40ede32b, 32'hc2ad7e0e, 32'hc27291e5};
test_bias[358:358] = '{32'h409fa802};
test_output[358:358] = '{32'h45cb2b97};
test_input[2872:2879] = '{32'hc221c367, 32'h42a797d2, 32'h420aaa71, 32'h4275309d, 32'hc2a1e891, 32'hc2647182, 32'hc236e12a, 32'h424eb168};
test_weights[2872:2879] = '{32'h42bb18b7, 32'h41ff3383, 32'hc1ace008, 32'h42b8ecef, 32'hc21b1046, 32'h427f4405, 32'h42c015d8, 32'hc259505a};
test_bias[359:359] = '{32'h42ae2626};
test_output[359:359] = '{32'hc56e1184};
test_input[2880:2887] = '{32'h41ccfb16, 32'hc2926aad, 32'hc294573f, 32'h41cb7fb6, 32'hc1aa7118, 32'h410007df, 32'h41481ec7, 32'h42b692b1};
test_weights[2880:2887] = '{32'h42aebf7b, 32'h4252dea0, 32'h4297b461, 32'hc17c815b, 32'hc23d6a67, 32'h41006867, 32'hc1b531e2, 32'h4122b691};
test_bias[360:360] = '{32'h42b1ef05};
test_output[360:360] = '{32'hc5b68750};
test_input[2888:2895] = '{32'h42379ef3, 32'h4162b46b, 32'h424de989, 32'h41958823, 32'hc225fa90, 32'h42bfb359, 32'h41a30721, 32'hc2ba1dcd};
test_weights[2888:2895] = '{32'h42c314c6, 32'h3ee1add3, 32'h42bc0184, 32'h4294a647, 32'hc1859ad3, 32'hc1fe8d9d, 32'h42aa4f95, 32'hc2b47270};
test_bias[361:361] = '{32'hc2aea3c5};
test_output[361:361] = '{32'h468fbebb};
test_input[2896:2903] = '{32'hc29b2246, 32'h41519b4d, 32'h4295b7ca, 32'hc1b8d680, 32'h42c5aa73, 32'h40a3c97c, 32'hc282491a, 32'hc2684090};
test_weights[2896:2903] = '{32'h41e90397, 32'h4297c451, 32'hc2a1243a, 32'h4229452a, 32'h414e612e, 32'h42c77054, 32'hc2a12d01, 32'h41e730a9};
test_bias[362:362] = '{32'hc1e22898};
test_output[362:362] = '{32'hc5381a1a};
test_input[2904:2911] = '{32'h419205f1, 32'hc269a285, 32'hc29a716a, 32'hc1227af1, 32'h42954b02, 32'hc009b892, 32'h42270e81, 32'h42839022};
test_weights[2904:2911] = '{32'h42953d42, 32'hc1e201d4, 32'hc25cc4a7, 32'hc1f152fb, 32'hc1ca8136, 32'h41832441, 32'h4254d06e, 32'h414e5b79};
test_bias[363:363] = '{32'hc2a5a966};
test_output[363:363] = '{32'h46070cf1};
test_input[2912:2919] = '{32'hc1b5bc46, 32'h429754f8, 32'hc24e6a5f, 32'h42afc1ff, 32'h42bbc947, 32'hc218b04b, 32'hc2acebcb, 32'h429214de};
test_weights[2912:2919] = '{32'hc124c1e8, 32'hc25f6952, 32'h4096c0ca, 32'hc24b544d, 32'h41a41142, 32'h42c77f9b, 32'hc2b811d1, 32'hc22d6f27};
test_bias[364:364] = '{32'h42b2d82b};
test_output[364:364] = '{32'hc5b244ef};
test_input[2920:2927] = '{32'hc21dbb0c, 32'hbfb7191e, 32'hc2aeaa72, 32'h3fef356c, 32'hc25b825d, 32'h41a16408, 32'hc295d094, 32'h42af5dcb};
test_weights[2920:2927] = '{32'h40cfc7b2, 32'h424d4a8b, 32'h4250a825, 32'h425c75b5, 32'hc29898b2, 32'h42889fc6, 32'hc2a7af1f, 32'hc2aa735c};
test_bias[365:365] = '{32'hc2a97e18};
test_output[365:365] = '{32'hc3f71153};
test_input[2928:2935] = '{32'hc2c2c40b, 32'h426b9960, 32'hc20c0d49, 32'hc15bdc50, 32'h42769451, 32'hc295e1e5, 32'hc2773a25, 32'hc088b8ec};
test_weights[2928:2935] = '{32'hc2908710, 32'hc1272396, 32'h423cc3ad, 32'hc17d8e7b, 32'hc296babc, 32'h42a6ffdc, 32'h41e15ee1, 32'hc1f9a48c};
test_bias[366:366] = '{32'hc2910162};
test_output[366:366] = '{32'hc5ed62a3};
test_input[2936:2943] = '{32'hc0f6453a, 32'h428c46e1, 32'hc14aa73e, 32'hc2c65ff6, 32'h4250b5db, 32'h42bfc95b, 32'h4260457a, 32'h41988210};
test_weights[2936:2943] = '{32'hc29284a3, 32'hc2a89a7d, 32'h42b9a517, 32'hc2be9dbb, 32'h41bf040f, 32'hc1c71828, 32'h41255340, 32'hc21d075f};
test_bias[367:367] = '{32'h429b2777};
test_output[367:367] = '{32'h44d41328};
test_input[2944:2951] = '{32'h41352116, 32'hc2896aaf, 32'h42865459, 32'h41725483, 32'hc1c89149, 32'hc1c244e1, 32'hc224cda5, 32'hc1986312};
test_weights[2944:2951] = '{32'hc1aec146, 32'h42139ec4, 32'hc1f62afd, 32'h42102c61, 32'h4272e0e8, 32'h42be2a6b, 32'h42af60d6, 32'h3e2c60b9};
test_bias[368:368] = '{32'hc28f4819};
test_output[368:368] = '{32'hc638bb14};
test_input[2952:2959] = '{32'hc28d3813, 32'h420ab300, 32'h41d793bb, 32'hc18457ca, 32'hc285ec0a, 32'hc2071f7a, 32'h41c49be0, 32'h421ec33c};
test_weights[2952:2959] = '{32'h42a1a853, 32'hc277b6e4, 32'h415e321d, 32'h41d52f02, 32'hc1fa1e08, 32'h418deb6d, 32'h42a74b6c, 32'hc2c4e5fe};
test_bias[369:369] = '{32'h427b8156};
test_output[369:369] = '{32'hc6005fb0};
test_input[2960:2967] = '{32'hc257f370, 32'hc238978d, 32'hc17dc540, 32'hc0812247, 32'h42c0cde4, 32'h42c65d96, 32'hc282c699, 32'hc29cf011};
test_weights[2960:2967] = '{32'h41313fe8, 32'h422c7487, 32'hc242482c, 32'hc28d36c4, 32'h3fdcae35, 32'h41cf94e4, 32'h41a279f9, 32'hc1e542cf};
test_bias[370:370] = '{32'hc2b2d51c};
test_output[370:370] = '{32'h44fed5ac};
test_input[2968:2975] = '{32'hc2659abe, 32'h3f2405f0, 32'h42be374d, 32'hc29316f7, 32'hc2bb8202, 32'h42a1bf82, 32'hc249d6e1, 32'h42144193};
test_weights[2968:2975] = '{32'h429df899, 32'h42a063f9, 32'h42accfa0, 32'h409a2db2, 32'hc063060b, 32'hc2a0885d, 32'hc2379e97, 32'h42a2b63d};
test_bias[371:371] = '{32'hc24b689e};
test_output[371:371] = '{32'h451c705a};
test_input[2976:2983] = '{32'h40237ab2, 32'h402497a4, 32'h428d4daf, 32'hc21d3707, 32'h42b662f3, 32'h417a36a9, 32'h429ac173, 32'h42782726};
test_weights[2976:2983] = '{32'h427c6bf4, 32'hc27288c7, 32'hc2801404, 32'hc21ff13b, 32'h41c244f9, 32'hc24f8510, 32'h42a02cf5, 32'hc2bd5714};
test_bias[372:372] = '{32'hc147f45e};
test_output[372:372] = '{32'hc49a228a};
test_input[2984:2991] = '{32'hc293df68, 32'hc2c22d3e, 32'h42743532, 32'h42821264, 32'hc209e30c, 32'h41b5e547, 32'h403017c4, 32'hc2a70731};
test_weights[2984:2991] = '{32'hc2b5458b, 32'h42af8733, 32'hc0dbff73, 32'hc2a6f22a, 32'h427655b3, 32'hc1e9e6ff, 32'h427d8148, 32'hc1b15676};
test_bias[373:373] = '{32'h42a5313b};
test_output[373:373] = '{32'hc6026df1};
test_input[2992:2999] = '{32'hc2895268, 32'hc1e82cb6, 32'h40890d75, 32'h429af64a, 32'hc2c03bab, 32'h419547e1, 32'hc0cce4ad, 32'h40f54796};
test_weights[2992:2999] = '{32'h420bcf59, 32'h42520892, 32'hc231812e, 32'h41904701, 32'h42b88497, 32'h429971d0, 32'hc2369c63, 32'h427c66b8};
test_bias[374:374] = '{32'hc0d534c3};
test_output[374:374] = '{32'hc6129c84};
test_input[3000:3007] = '{32'hc27c3c12, 32'h429d1cf4, 32'hc1e6e722, 32'hc1130f09, 32'hc2ac87c7, 32'hc209a446, 32'h428aabf1, 32'hc27a56ab};
test_weights[3000:3007] = '{32'h425f32a9, 32'h42878028, 32'h41da9917, 32'h42bf4b8b, 32'h41560680, 32'hc211abc4, 32'h42a83aa9, 32'hc21a3b40};
test_bias[375:375] = '{32'hc2a207ad};
test_output[375:375] = '{32'h46033d29};
test_input[3008:3015] = '{32'hc2bc3122, 32'hc226db68, 32'hc15364b6, 32'hc1b38ea3, 32'h42c0e9f4, 32'hc2a35f9f, 32'h42942b75, 32'hc24b5af7};
test_weights[3008:3015] = '{32'hc274322c, 32'h42847d07, 32'hc28ba023, 32'hc28f25e3, 32'h426c41c4, 32'h42a29c05, 32'hc0ea56c3, 32'h42006e15};
test_bias[376:376] = '{32'hc2101ca2};
test_output[376:376] = '{32'h45132baf};
test_input[3016:3023] = '{32'hc271c3e4, 32'hc28cfd4e, 32'hc1494407, 32'h4286c170, 32'hc1c795c9, 32'h4287ae5d, 32'hc2b30341, 32'h415b3ca7};
test_weights[3016:3023] = '{32'h42b9ffb1, 32'h42b7523a, 32'hc21b36ca, 32'hc13a5399, 32'h421e4a66, 32'h41fe377b, 32'h4269cacb, 32'h42844228};
test_bias[377:377] = '{32'hc2809dca};
test_output[377:377] = '{32'hc673c112};
test_input[3024:3031] = '{32'h42b0cee3, 32'h417b2ed5, 32'h42a8ada5, 32'h42a3a1c2, 32'hc29fbaf0, 32'hc18d3fbd, 32'h42727287, 32'h41d28938};
test_weights[3024:3031] = '{32'hc2b0ecdb, 32'hc1de5cb6, 32'h41a89c1e, 32'hc1b5cea8, 32'h42c0590c, 32'hc2961e6c, 32'hc29077c7, 32'hc29349b4};
test_bias[378:378] = '{32'h4294fc14};
test_output[378:378] = '{32'hc6a39039};
test_input[3032:3039] = '{32'hc2c6b9d5, 32'hc2bb174e, 32'h41aa581a, 32'hc2035553, 32'hc282fc4f, 32'hc22ce95b, 32'h42a29a49, 32'hc29bd298};
test_weights[3032:3039] = '{32'hc29d1f89, 32'hc2b07cd2, 32'hc277f0f8, 32'h42661374, 32'h4193f2d7, 32'h42517f88, 32'h4222018b, 32'hc293a66f};
test_bias[379:379] = '{32'h420533a8};
test_output[379:379] = '{32'h46902e74};
test_input[3040:3047] = '{32'h42a85a0b, 32'hc287f85a, 32'h42ad0006, 32'hc268a6ad, 32'h4212c085, 32'h429961c9, 32'h4293fcbb, 32'h426f49fe};
test_weights[3040:3047] = '{32'h41093769, 32'h405ae1e1, 32'h4252f197, 32'hc2333404, 32'h42bbd626, 32'hc03fd26a, 32'hc1c06314, 32'h405e7183};
test_bias[380:380] = '{32'hc24228d2};
test_output[380:380] = '{32'h46109236};
test_input[3048:3055] = '{32'hc2602212, 32'h41ce7bff, 32'hbf838f14, 32'hbeee28eb, 32'hc20e11a2, 32'hc2816365, 32'h424bac78, 32'hc2b33896};
test_weights[3048:3055] = '{32'hc07f626f, 32'hc1578f62, 32'h420bfbb2, 32'hc29af21e, 32'h41fc0e97, 32'hc098b593, 32'h4223d5d9, 32'hc11d1f1c};
test_bias[381:381] = '{32'hc29805c6};
test_output[381:381] = '{32'h44f464b6};
test_input[3056:3063] = '{32'hc139e585, 32'h4229d101, 32'hc0049489, 32'h428e8ed6, 32'hc2668a9f, 32'hc25c82d7, 32'hc22df867, 32'h4291b491};
test_weights[3056:3063] = '{32'h40b6958e, 32'h42a42218, 32'h4163a872, 32'hc1a3ed32, 32'h42721911, 32'h42910cbf, 32'h42b77b28, 32'h422413c4};
test_bias[382:382] = '{32'hc28d2873};
test_output[382:382] = '{32'hc5cf3804};
test_input[3064:3071] = '{32'h42223287, 32'h41c0c39e, 32'hc2bc466d, 32'hc1e59547, 32'h40a891fa, 32'h420fb2f6, 32'hc206f48b, 32'h4159873a};
test_weights[3064:3071] = '{32'hc2b76c11, 32'hc2b0a178, 32'hc1113b8f, 32'hc2b35e64, 32'h421309b4, 32'h4241c78d, 32'h4209ae22, 32'h421ccf94};
test_bias[383:383] = '{32'hc237fc6a};
test_output[383:383] = '{32'hc490dc2a};
test_input[3072:3079] = '{32'h4273d0fe, 32'hbe30c573, 32'h428f8dcb, 32'h42c0e576, 32'hc20696c0, 32'hc27c76a6, 32'h42b45ffd, 32'h4246fe08};
test_weights[3072:3079] = '{32'h402c81b3, 32'h42c517a4, 32'h4296d30d, 32'hc24b39b5, 32'hc2148b3c, 32'hc296c2e0, 32'h423a2b0d, 32'h41418adb};
test_bias[384:384] = '{32'hc202ecbb};
test_output[384:384] = '{32'h4632a6fe};
test_input[3080:3087] = '{32'hc2b6d80d, 32'hc1879fcd, 32'h41bf2056, 32'h40bbd0fb, 32'hc294bdf6, 32'hc1d11e1d, 32'hc13423ca, 32'h426fee82};
test_weights[3080:3087] = '{32'h4264e834, 32'h4137c0ef, 32'h42749161, 32'h42c39508, 32'hc1e4a841, 32'hc031d9f3, 32'h428c747a, 32'h41facf2a};
test_bias[385:385] = '{32'h4206d6c0};
test_output[385:385] = '{32'hc28bcada};
test_input[3088:3095] = '{32'hc213b602, 32'hc221bc84, 32'h428793f7, 32'hc1cd3b53, 32'hc19a3991, 32'hc0b66e36, 32'h42586314, 32'hc22b6bf7};
test_weights[3088:3095] = '{32'hc2bf7e14, 32'hc28ab9f8, 32'hc1efcb2f, 32'h42bfce7f, 32'hc26d11f9, 32'h41fef25f, 32'hc233d231, 32'h4295fca9};
test_bias[386:386] = '{32'h40d9b0bb};
test_output[386:386] = '{32'hc530e036};
test_input[3096:3103] = '{32'hc231e387, 32'hc2b8edf1, 32'hc26b8a4b, 32'hc2ad3309, 32'h420569f1, 32'h4184b3a0, 32'hc2acee39, 32'h42423b1c};
test_weights[3096:3103] = '{32'h421737e2, 32'h4231ec52, 32'h418ca697, 32'hc1f01e71, 32'h40b8f8ff, 32'h428e47f0, 32'hc27a357c, 32'h4291e703};
test_bias[387:387] = '{32'h42a58b4d};
test_output[387:387] = '{32'h45c10347};
test_input[3104:3111] = '{32'hc2afcbed, 32'hc0a264af, 32'h41e9e143, 32'h42bf8015, 32'h405eb958, 32'hc27917df, 32'hbf22c1d6, 32'hc2a0aac0};
test_weights[3104:3111] = '{32'h42bf84c6, 32'hc219b8a4, 32'h429825ad, 32'hc2190d03, 32'h41b08088, 32'hc22791b2, 32'h418a0731, 32'h4136d931};
test_bias[388:388] = '{32'h40b755c3};
test_output[388:388] = '{32'hc5f6db95};
test_input[3112:3119] = '{32'hc295a390, 32'hc1a142d2, 32'h414da803, 32'h426d418a, 32'hc20bacff, 32'h42aad46b, 32'hc29fd965, 32'h428aedc1};
test_weights[3112:3119] = '{32'hc23dbc4e, 32'hc0d398b3, 32'h41b9fb37, 32'hc1aa1928, 32'h42a8d422, 32'hc1862881, 32'h3ebd51ea, 32'h425742f0};
test_bias[389:389] = '{32'hc1a2f827};
test_output[389:389] = '{32'h44fd86b7};
test_input[3120:3127] = '{32'hbf26bac0, 32'h42779148, 32'hc191dc2c, 32'h429fe1cd, 32'hc28f0236, 32'hc1ffff0a, 32'h41615a54, 32'hc2adb7fc};
test_weights[3120:3127] = '{32'hc2392fbc, 32'h414ec44f, 32'h4209d6b1, 32'h42b8f92b, 32'h42a53e2b, 32'hc0fa7092, 32'h42be04a9, 32'hc0767a56};
test_bias[390:390] = '{32'hc29c32ef};
test_output[390:390] = '{32'h455cc644};
test_input[3128:3135] = '{32'hc298f350, 32'hc29b1aa2, 32'hc2b2477d, 32'h41b8b8af, 32'hc0c51ca6, 32'hc29f12ca, 32'hc2a6ff50, 32'hc0ca8489};
test_weights[3128:3135] = '{32'h42982514, 32'hc2a23065, 32'hc1c56fc5, 32'hc1663769, 32'h423e4ed9, 32'h3eda7d0c, 32'h413246fd, 32'hc25a3e3e};
test_bias[391:391] = '{32'hc23008df};
test_output[391:391] = '{32'h44acdff6};
test_input[3136:3143] = '{32'hc29cfe34, 32'hc29ea85f, 32'h420eacb4, 32'hc2995e95, 32'h4245aa01, 32'h41fb7cb6, 32'hc2742186, 32'h42c2d062};
test_weights[3136:3143] = '{32'hc29e0bcd, 32'hc10778b1, 32'hc234de84, 32'h42a7702f, 32'h417dc428, 32'h4271c25e, 32'hc25eb44c, 32'h42753d04};
test_bias[392:392] = '{32'h416b14e0};
test_output[392:392] = '{32'h462a7975};
test_input[3144:3151] = '{32'h41abe121, 32'h42b54093, 32'h4210b409, 32'h42996d1c, 32'hc2aa1b85, 32'h42681f6d, 32'hc2b6dbeb, 32'hc185a445};
test_weights[3144:3151] = '{32'h428e9c2e, 32'h428f689d, 32'h415d32fb, 32'hc24fe929, 32'hc2a0307e, 32'hc08bcb0f, 32'h429f8d99, 32'hc2837c2e};
test_bias[393:393] = '{32'h420c3e8f};
test_output[393:393] = '{32'h459a69f2};
test_input[3152:3159] = '{32'h42028945, 32'h410d7ffc, 32'hc2ab45e9, 32'hc2ab65c4, 32'h4102f44a, 32'hc2643ef3, 32'hc2c4c3d9, 32'hc294a7a0};
test_weights[3152:3159] = '{32'hc2c4fbdc, 32'hc26a46fc, 32'h4172b1cb, 32'h42bc6574, 32'h4298ec99, 32'hc2be7161, 32'h416fab98, 32'hc1991909};
test_bias[394:394] = '{32'h419afe1f};
test_output[394:394] = '{32'hc5dd2361};
test_input[3160:3167] = '{32'h421be4b7, 32'h42bc8102, 32'hc27d138a, 32'hc27d347b, 32'h42b762d1, 32'h4283712f, 32'h428748bc, 32'hc29d31ad};
test_weights[3160:3167] = '{32'h4298d142, 32'h42aff3ed, 32'h41b8b066, 32'h42c3f862, 32'h427c50e4, 32'hc0973e2c, 32'h4293f965, 32'h41ae584e};
test_bias[395:395] = '{32'h423cf73d};
test_output[395:395] = '{32'h46420bb2};
test_input[3168:3175] = '{32'hc2c31382, 32'h4275ef00, 32'hc2416675, 32'hc2b344bd, 32'hc29d2b23, 32'hc1da78b8, 32'hc29e3cd2, 32'hc2c37cb5};
test_weights[3168:3175] = '{32'hc2b8bc62, 32'hc2439b50, 32'hc27dfaff, 32'hc238efd7, 32'h4042b114, 32'h4156deea, 32'h41fc92c9, 32'h4202969a};
test_bias[396:396] = '{32'hc295bfb8};
test_output[396:396] = '{32'h45d5fa48};
test_input[3176:3183] = '{32'hc2013333, 32'hc1f98158, 32'hc291cf13, 32'hc2bf9ae4, 32'hc2c030a2, 32'hc2b8081f, 32'hbeea2e1e, 32'hc24511b4};
test_weights[3176:3183] = '{32'h416096dd, 32'hc107eb79, 32'h42a4dcfd, 32'hc297269a, 32'hc12022cf, 32'hc294ad8c, 32'hc2705148, 32'h4266ec99};
test_bias[397:397] = '{32'h422bb544};
test_output[397:397] = '{32'h45bdb429};
test_input[3184:3191] = '{32'hc20449a1, 32'hc002aa25, 32'h426c4c1a, 32'h428acd79, 32'h4214d7e8, 32'hc1e564cc, 32'hc24751d6, 32'hc29376d6};
test_weights[3184:3191] = '{32'h425333f7, 32'hc0f2439b, 32'h42b4f28a, 32'hc1c74941, 32'hc29fe214, 32'h42c09797, 32'hc2a75d1c, 32'h4234a9ea};
test_bias[398:398] = '{32'hc2462ced};
test_output[398:398] = '{32'hc53f4b3d};
test_input[3192:3199] = '{32'h42b930f5, 32'hc1d4dc03, 32'hbfd0b1db, 32'hc208a066, 32'h4287ee8e, 32'hc2339e51, 32'hc265d9b2, 32'hc2978f85};
test_weights[3192:3199] = '{32'h417bf6bf, 32'h410e2249, 32'h4275063b, 32'h4285d12f, 32'hc22668d3, 32'h42590c40, 32'h40f653af, 32'hc29185e1};
test_bias[399:399] = '{32'h42c65d03};
test_output[399:399] = '{32'hc49d1b57};
test_input[3200:3207] = '{32'hc27719f9, 32'hc22f3f7f, 32'hc2bd579b, 32'hc0144342, 32'h41749ca3, 32'h41a2fb12, 32'h425d6056, 32'h41831d43};
test_weights[3200:3207] = '{32'hc1489f74, 32'h41238864, 32'h42a3a093, 32'hc1ce4a8a, 32'hc26de31f, 32'h42b4e0fd, 32'hc251ad5e, 32'hc20448fc};
test_bias[400:400] = '{32'hc2966e7f};
test_output[400:400] = '{32'hc61b5fa1};
test_input[3208:3215] = '{32'hc2b64419, 32'hc2720d51, 32'hc1a554cc, 32'h429d1930, 32'hc14f6917, 32'hc2a99c6b, 32'h42bd3650, 32'h425c5e17};
test_weights[3208:3215] = '{32'hc2752956, 32'hc2aa63da, 32'hc267f67e, 32'h41ff6d78, 32'h422495c9, 32'hc18c8dca, 32'hc29215e2, 32'h42b6a116};
test_bias[401:401] = '{32'h42c7df20};
test_output[401:401] = '{32'h4654e149};
test_input[3216:3223] = '{32'hc291e207, 32'h42767c5c, 32'hc289975f, 32'hc211d3fd, 32'h40c08d5a, 32'h4135addd, 32'hc1d20cb4, 32'h422ef7a9};
test_weights[3216:3223] = '{32'hc2a2e7d6, 32'h42a38370, 32'hc2becae2, 32'h42831b04, 32'hc2a5240f, 32'h40147945, 32'hc1f1566d, 32'h4271b4c5};
test_bias[402:402] = '{32'hc2574417};
test_output[402:402] = '{32'h468d1e54};
test_input[3224:3231] = '{32'h423ace85, 32'hc262d675, 32'hc2889603, 32'hc2ae6377, 32'hc1c44903, 32'hc2270971, 32'h42a9fea1, 32'hc270679b};
test_weights[3224:3231] = '{32'hc26bdb4e, 32'h42c4afec, 32'h424eccf0, 32'h4247a4e2, 32'h42876889, 32'hc2b608fd, 32'h423ecd11, 32'hc2bda5f0};
test_bias[403:403] = '{32'h42437d07};
test_output[403:403] = '{32'hc5857bdf};
test_input[3232:3239] = '{32'hc1b783e1, 32'h423934b8, 32'hc28bf507, 32'hc2722176, 32'h41736ae3, 32'h428e9c09, 32'h4273971a, 32'h42c588af};
test_weights[3232:3239] = '{32'h40cbf82e, 32'hc2826af4, 32'hc271ecba, 32'hc1922d7b, 32'h421578b6, 32'hc2aeca7b, 32'hc2a938ca, 32'hc2b5bcd7};
test_bias[404:404] = '{32'h41ab4098};
test_output[404:404] = '{32'hc689788d};
test_input[3240:3247] = '{32'hc294cf76, 32'h42400175, 32'h42c1f34d, 32'hc27676c4, 32'hc225e72e, 32'h42449bd1, 32'h4247c5c0, 32'h411e12aa};
test_weights[3240:3247] = '{32'hc23b6374, 32'h42adc804, 32'h4190055a, 32'h4206c834, 32'h4265b254, 32'hc1dbde90, 32'hc21bb21e, 32'h4286e8a9};
test_bias[405:405] = '{32'hc21c206f};
test_output[405:405] = '{32'h450e4fb8};
test_input[3248:3255] = '{32'hc29a18ee, 32'h42981046, 32'h427cf6b9, 32'hc240babc, 32'hc236c611, 32'hc13d95ca, 32'hc2688bd6, 32'hc2aec020};
test_weights[3248:3255] = '{32'h41b527d6, 32'h42607903, 32'h4055513f, 32'hc2346cbf, 32'hc2535496, 32'hc2c23212, 32'hc2aa120d, 32'hc22b4629};
test_bias[406:406] = '{32'hc19db0b3};
test_output[406:406] = '{32'h4685dffe};
test_input[3256:3263] = '{32'hc2974929, 32'hc24c5919, 32'h420cad3c, 32'h411745cc, 32'h420e7e75, 32'hc1cc2ad4, 32'hc23de39f, 32'h41a10f66};
test_weights[3256:3263] = '{32'h42c1b8e7, 32'hc2be3499, 32'h429ed665, 32'h42a440e7, 32'h41f8e8e2, 32'h4251d902, 32'hc26acfa3, 32'hc212c053};
test_bias[407:407] = '{32'hc2b142f4};
test_output[407:407] = '{32'h4530e3a6};
test_input[3264:3271] = '{32'hc24c8f82, 32'h410dcd0b, 32'hc2a93e9f, 32'h428e9d50, 32'hc2ab5d88, 32'hc2bb356d, 32'hc28ce305, 32'h421ee370};
test_weights[3264:3271] = '{32'hc232862a, 32'h42c005b7, 32'hc29e781f, 32'hc220833e, 32'hc28ac44f, 32'h4236ecaf, 32'hc2a78c26, 32'h428dfa95};
test_bias[408:408] = '{32'h42a23c1a};
test_output[408:408] = '{32'h4688470c};
test_input[3272:3279] = '{32'h4250bccf, 32'h4256b756, 32'h4198545e, 32'h42b4a3f3, 32'h4286a873, 32'h3fff3f03, 32'hc2b2c312, 32'hc2475516};
test_weights[3272:3279] = '{32'hc21142e0, 32'h426e032d, 32'h421f2a5f, 32'h42be3b0a, 32'hc1d49ef1, 32'h40c25314, 32'hc25af23e, 32'hc25a63e5};
test_bias[409:409] = '{32'h42408639};
test_output[409:409] = '{32'h468126eb};
test_input[3280:3287] = '{32'h42700530, 32'hc0d9af5b, 32'h41f9bd03, 32'hc2c2a837, 32'hc2a0901a, 32'h42b6d438, 32'h42a3c80d, 32'h421ad920};
test_weights[3280:3287] = '{32'hc239c6e0, 32'h42a8e5ef, 32'h42b6492b, 32'h40a82b7b, 32'hc2c5a8c6, 32'hc1575b18, 32'h426f4815, 32'hc2bd5fb8};
test_bias[410:410] = '{32'h429185fb};
test_output[410:410] = '{32'h45da30f6};
test_input[3288:3295] = '{32'h3f34a506, 32'h4249724e, 32'hc2529b4c, 32'hc1682cba, 32'h41e8b682, 32'h42965e73, 32'hc07115fc, 32'h4278ac64};
test_weights[3288:3295] = '{32'h42727393, 32'hc1bb76d3, 32'h425ec986, 32'h426d7777, 32'hc2ae696a, 32'hc1a5b9c7, 32'h428db6bf, 32'h42b3b5b5};
test_bias[411:411] = '{32'hc133ac08};
test_output[411:411] = '{32'hc56859aa};
test_input[3296:3303] = '{32'hc211be1d, 32'hc16965f0, 32'h4155c326, 32'h41ae274d, 32'hc2aa3cff, 32'hc2949d1e, 32'hc1a88bcc, 32'hc130499c};
test_weights[3296:3303] = '{32'hc2ba631e, 32'h41536669, 32'h42bf0cb9, 32'hc28cca10, 32'h4238ed81, 32'hc167b142, 32'h420c0436, 32'h42669976};
test_bias[412:412] = '{32'h42b11c4d};
test_output[412:412] = '{32'hc49595cc};
test_input[3304:3311] = '{32'h41dfb3bc, 32'hc09ee9d0, 32'hc2301d6d, 32'h41b834ac, 32'h429ca40d, 32'h41df597b, 32'hc1a22284, 32'h42a24acc};
test_weights[3304:3311] = '{32'h41aeed53, 32'h4239746f, 32'h425b1bd6, 32'h42c0340b, 32'h4128b5f4, 32'hc161224a, 32'hc1f984e8, 32'h42852723};
test_bias[413:413] = '{32'h42ad0886};
test_output[413:413] = '{32'h45d28246};
test_input[3312:3319] = '{32'h41b50539, 32'hc28de9e2, 32'h4259019b, 32'h411dc9fc, 32'h425e4956, 32'h41e888fa, 32'hc2030446, 32'hc1ca3493};
test_weights[3312:3319] = '{32'hc2005428, 32'h415e0f43, 32'h418ff0cb, 32'hc1e91b9a, 32'h42b03c7b, 32'h401b88df, 32'hc2c6217b, 32'h42a0e58e};
test_bias[414:414] = '{32'hc18e1e26};
test_output[414:414] = '{32'h45a09993};
test_input[3320:3327] = '{32'h42c6f86b, 32'h409ac2ba, 32'h4248c62c, 32'h42aeef07, 32'h42bfc0f7, 32'h41c72b50, 32'h429e4ed4, 32'hc21e1c82};
test_weights[3320:3327] = '{32'h426dbb57, 32'h41e84907, 32'h429663b9, 32'h427899d8, 32'h41bee727, 32'h4271f40d, 32'h42311a11, 32'hc1cc47dd};
test_bias[415:415] = '{32'h42c20d94};
test_output[415:415] = '{32'h46b8e88c};
test_input[3328:3335] = '{32'hc2b5399c, 32'h401086b6, 32'hc27188d1, 32'h4291b88c, 32'hc29907c7, 32'hc0506103, 32'hc2b8b598, 32'hc25ec852};
test_weights[3328:3335] = '{32'hc150bdc8, 32'hc20ea306, 32'h42bd6b01, 32'hc23bdc65, 32'h410abf39, 32'hc292fd48, 32'hc28077c4, 32'h4211f5c2};
test_bias[416:416] = '{32'h428ed3cc};
test_output[416:416] = '{32'hc58c5fde};
test_input[3336:3343] = '{32'h42bd4c46, 32'h42575bd6, 32'h42ae3578, 32'hc2931412, 32'h3f1f0a6b, 32'hc2572e3f, 32'hc18abdaf, 32'h42a88499};
test_weights[3336:3343] = '{32'hc1801ccc, 32'h42890209, 32'h4281d6fd, 32'h4289aedc, 32'hc235bc3e, 32'h42b00f15, 32'hc207c234, 32'hc2218f90};
test_bias[417:417] = '{32'hc2949ebc};
test_output[417:417] = '{32'hc598bf9b};
test_input[3344:3351] = '{32'h41967229, 32'h428a0259, 32'hc28caac1, 32'hc262ee0d, 32'h42b533db, 32'h42bb7e84, 32'hc187cfe3, 32'h40c6e0d7};
test_weights[3344:3351] = '{32'hc20f543f, 32'hc1e967fb, 32'h415a3e86, 32'hc2365a2d, 32'h42594e85, 32'h420ae86c, 32'h42abfacb, 32'h429fe857};
test_bias[418:418] = '{32'hc2b6c9b5};
test_output[418:418] = '{32'h45bd7959};
test_input[3352:3359] = '{32'hc2a67bac, 32'h42066780, 32'h41a3afff, 32'hc25895bd, 32'h42218a71, 32'h42635528, 32'hc15d9a08, 32'h42399854};
test_weights[3352:3359] = '{32'hc2372134, 32'hc15b6492, 32'h419fb726, 32'hc2352dde, 32'hc2bf1b8b, 32'hc1f24021, 32'h429f6ba1, 32'h41c5c001};
test_bias[419:419] = '{32'hc200ec28};
test_output[419:419] = '{32'h442082ea};
test_input[3360:3367] = '{32'h426608ff, 32'hc242878f, 32'hc1f81f88, 32'h41c7ab15, 32'h427d7287, 32'h4297cce5, 32'hc1fa9284, 32'hc24d4cd6};
test_weights[3360:3367] = '{32'h41206af3, 32'hc06ae6d6, 32'hc04a24ba, 32'h414d231b, 32'hc27f1e9e, 32'h421ca39e, 32'hc2674537, 32'hc2878dc0};
test_bias[420:420] = '{32'h42584624};
test_output[420:420] = '{32'h45aa3dc4};
test_input[3368:3375] = '{32'hc24e2dfd, 32'hc27971dc, 32'h40acf891, 32'hc1984dcb, 32'hc0bdf19a, 32'h426a42b7, 32'hc2b0e9f9, 32'hc25add13};
test_weights[3368:3375] = '{32'h42a1e139, 32'hc2c2c42a, 32'h423d9141, 32'h41cf7868, 32'hc2339b11, 32'hc09eabb4, 32'hc1eb164b, 32'h41ef4788};
test_bias[421:421] = '{32'hc2bd98a9};
test_output[421:421] = '{32'h451cb806};
test_input[3376:3383] = '{32'h42bfca8b, 32'hc2c00bdb, 32'hc190750c, 32'h42a26242, 32'h403e4884, 32'hc2b420f4, 32'h42a19229, 32'h422d248f};
test_weights[3376:3383] = '{32'h424519c8, 32'h42885462, 32'h41b60e16, 32'h4144c435, 32'hc290a5ed, 32'hc1965f59, 32'hc25548c1, 32'h42bc0535};
test_bias[422:422] = '{32'hc28f9e3c};
test_output[422:422] = '{32'hc2818bf0};
test_input[3384:3391] = '{32'hc118f975, 32'h4280256e, 32'h42366b6a, 32'hc2c65968, 32'hc14cbabe, 32'hc269b3e9, 32'hc28d2a45, 32'hc18196fd};
test_weights[3384:3391] = '{32'hc2694897, 32'h42afa2c3, 32'hc261bd61, 32'hc2c3a19c, 32'hc0f57553, 32'h427c55dc, 32'hc04e82ef, 32'h4211cb71};
test_bias[423:423] = '{32'h425999df};
test_output[423:423] = '{32'h46131e96};
test_input[3392:3399] = '{32'hc2a47b97, 32'h42901ec7, 32'h4218e4a4, 32'h424558bc, 32'hc26f0e7a, 32'hc245b74d, 32'hc2998cec, 32'h41ef0509};
test_weights[3392:3399] = '{32'h42bd27dd, 32'hc204f738, 32'hc1f8c4b8, 32'hc2c42864, 32'hc1fe88f8, 32'h40be3358, 32'h412aa83f, 32'h42a7f3e5};
test_bias[424:424] = '{32'hc2a0e566};
test_output[424:424] = '{32'hc64adeca};
test_input[3400:3407] = '{32'hc29eb727, 32'h4213992e, 32'hc243fcb1, 32'hc209053c, 32'hc1d91f64, 32'hc26b19c9, 32'hc27f09ed, 32'h409cde1c};
test_weights[3400:3407] = '{32'h42af59c8, 32'h42963c7b, 32'h423ca2af, 32'h409f3431, 32'hc13a0d97, 32'h41cc19fc, 32'h4298fb97, 32'hc2a1353e};
test_bias[425:425] = '{32'hc23ab005};
test_output[425:425] = '{32'hc64dc6eb};
test_input[3408:3415] = '{32'hc1ed944c, 32'h3f9ea0cb, 32'hc25a29fa, 32'hc17a78c8, 32'hc28a2bed, 32'hc15e207b, 32'h3fea2370, 32'h42c0f6a9};
test_weights[3408:3415] = '{32'h421cc9cd, 32'h424a747a, 32'h42a3aebb, 32'h427b4f31, 32'h4281f51d, 32'hc285af2a, 32'h41bb1797, 32'h423c5e7f};
test_bias[426:426] = '{32'hc0096154};
test_output[426:426] = '{32'hc5acac34};
test_input[3416:3423] = '{32'hc13d84ee, 32'hc1f0bfca, 32'hc2182183, 32'h4246a8e0, 32'hc1a59008, 32'hc2a28db9, 32'hc2124256, 32'h401bde1c};
test_weights[3416:3423] = '{32'hc2b74868, 32'h4219161e, 32'h424cbba2, 32'h42836afb, 32'h42aa30d4, 32'h4244a51f, 32'hc0fc7d42, 32'hc2a5e4f8};
test_bias[427:427] = '{32'h41e8359d};
test_output[427:427] = '{32'hc589356c};
test_input[3424:3431] = '{32'hc295f5fd, 32'h42b0e533, 32'h41c32476, 32'h42329d3e, 32'h42a9a613, 32'hc299f8bf, 32'h429650e1, 32'h42009d15};
test_weights[3424:3431] = '{32'h42a2f565, 32'hc1aa9bbd, 32'h429e48fd, 32'hc2b5ed49, 32'hc1936cf3, 32'h4226d111, 32'h4289df5b, 32'h4205c0b4};
test_bias[428:428] = '{32'h42942df0};
test_output[428:428] = '{32'hc605e976};
test_input[3432:3439] = '{32'h41d898b6, 32'hc269e906, 32'hc2b4f7a7, 32'hc21b8627, 32'h41956570, 32'h416a30bc, 32'h42877a5f, 32'h420f92ce};
test_weights[3432:3439] = '{32'h42c408cc, 32'hc28e94d3, 32'h410a0539, 32'hc236b92f, 32'hc298f71f, 32'h4179ce9e, 32'hc2001a9d, 32'hc187bacd};
test_bias[429:429] = '{32'h42bef959};
test_output[429:429] = '{32'h4575f9bd};
test_input[3440:3447] = '{32'h3fff025b, 32'hc04be015, 32'hc2156aa3, 32'h4225f5d2, 32'hc134d2cf, 32'hc22b8df8, 32'hc1fb0c52, 32'h429b34d7};
test_weights[3440:3447] = '{32'h424b67c0, 32'h4234b46e, 32'hc28489a5, 32'hc284b056, 32'h420cb407, 32'h4236bf0a, 32'hc1b3e93e, 32'hc2001c54};
test_bias[430:430] = '{32'h422f5fd5};
test_output[430:430] = '{32'hc589e565};
test_input[3448:3455] = '{32'hc26f5468, 32'hc1bcf181, 32'hc22fa942, 32'h41efc0ee, 32'h42b40974, 32'h41185520, 32'hc2c0321b, 32'hc2721b37};
test_weights[3448:3455] = '{32'h424972e9, 32'h42295de7, 32'h42ad42ac, 32'hc2b09d39, 32'h41e548e9, 32'hc2828460, 32'hc294ddd3, 32'hc266b4bd};
test_bias[431:431] = '{32'hc2b270ad};
test_output[431:431] = '{32'h45001169};
test_input[3456:3463] = '{32'hc24d8f67, 32'h41b81576, 32'hc2264586, 32'h42832f24, 32'h41e94b2f, 32'h428f1489, 32'hc2b36c6b, 32'hc2708ea0};
test_weights[3456:3463] = '{32'h42948d46, 32'h41efef2a, 32'hc1c260d6, 32'hc2c44268, 32'hc1627d99, 32'h42bfd2cd, 32'hc0e2e3a1, 32'hc265318e};
test_bias[432:432] = '{32'hc260371b};
test_output[432:432] = '{32'h44f025dd};
test_input[3464:3471] = '{32'h42b0009c, 32'h4246279b, 32'h42052a8e, 32'h4219210f, 32'hc2b3ea28, 32'h42073dd1, 32'h411eed60, 32'h42ac678b};
test_weights[3464:3471] = '{32'h42c21421, 32'h42b7f8f2, 32'hc29cbba7, 32'h42b66f4a, 32'h41c8da2d, 32'hc1e5e5d3, 32'hc265e60b, 32'h420acf86};
test_bias[433:433] = '{32'hc1047b44};
test_output[433:433] = '{32'h464da6a1};
test_input[3472:3479] = '{32'hc29156dc, 32'hc25a8214, 32'hc2283fe1, 32'hc225b279, 32'h40eaab9d, 32'h42a38275, 32'hc1772a1a, 32'hc2861fc1};
test_weights[3472:3479] = '{32'h42b3d9c7, 32'h42a6e69d, 32'hc00aee7d, 32'h426ea77a, 32'h416c72f6, 32'hc29ce02d, 32'hc2b15784, 32'h424b3c4e};
test_bias[434:434] = '{32'hc2a79a07};
test_output[434:434] = '{32'hc6ab16c1};
test_input[3480:3487] = '{32'h3f422baa, 32'h42833d12, 32'h41ec7f8e, 32'h41978f43, 32'h40a0fc75, 32'h41686495, 32'h40a3e88a, 32'hc295ffcd};
test_weights[3480:3487] = '{32'h42ae7863, 32'hc2008aa2, 32'h42882840, 32'h421837e0, 32'hc27e0b5b, 32'hc0d5b02d, 32'h4244d884, 32'hc26b5a7e};
test_bias[435:435] = '{32'h429a7bd5};
test_output[435:435] = '{32'h459cc504};
test_input[3488:3495] = '{32'h41a7412e, 32'hc2a658bc, 32'hc2b8e99e, 32'hc1ecdaee, 32'hc2293deb, 32'h42b56d80, 32'h4107444e, 32'hc19dbdba};
test_weights[3488:3495] = '{32'hc22d95b6, 32'hc234993a, 32'h42b11844, 32'hc20f3d83, 32'h3f8e6d48, 32'h418adf64, 32'h428cf1f8, 32'h42876684};
test_bias[436:436] = '{32'h424223a8};
test_output[436:436] = '{32'hc5571818};
test_input[3496:3503] = '{32'h40ed2e4f, 32'h4273ab55, 32'hc1955f51, 32'hc2c2a9b6, 32'hc181f750, 32'h420640bf, 32'hc20c2d7a, 32'h424dce80};
test_weights[3496:3503] = '{32'h4209963c, 32'h421b77b2, 32'h41c3f986, 32'h41e6eec3, 32'hc19790d0, 32'h42c60a56, 32'h4242cd0a, 32'h42904cc2};
test_bias[437:437] = '{32'h42c6903d};
test_output[437:437] = '{32'h459f1d47};
test_input[3504:3511] = '{32'h3cca62a3, 32'hc297c96b, 32'h42045933, 32'hc24e8724, 32'h41ea15f0, 32'hc2c6bf3b, 32'h428db55c, 32'hc266e51f};
test_weights[3504:3511] = '{32'h409194db, 32'hc16238ec, 32'h42065e23, 32'h41a9cb64, 32'h42b9e7de, 32'h409b749a, 32'hc2342c52, 32'hc0bca890};
test_bias[438:438] = '{32'hc22f5668};
test_output[438:438] = '{32'h43d76d59};
test_input[3512:3519] = '{32'hc238725d, 32'h421cb0ad, 32'h42340f95, 32'hc28394b0, 32'hc2942a4e, 32'h428fbac1, 32'h42a94f91, 32'h42c29576};
test_weights[3512:3519] = '{32'h42882cf5, 32'h4232c853, 32'hc18a9842, 32'h4299da92, 32'h429c52ae, 32'hbe8e3e11, 32'hc24b20fa, 32'hc1824c6a};
test_bias[439:439] = '{32'h414f9dd9};
test_output[439:439] = '{32'hc693bd72};
test_input[3520:3527] = '{32'hc26ec279, 32'hc2b36f06, 32'hc1547563, 32'h42bdcf32, 32'hc2a1dd71, 32'h41c40098, 32'h40fd7882, 32'h429dab02};
test_weights[3520:3527] = '{32'hc1fd8117, 32'h4287a2eb, 32'hc14691a6, 32'hc2880157, 32'h42a03c0b, 32'hc24e0636, 32'hbf915c9e, 32'hc298e97f};
test_bias[440:440] = '{32'h41a4b865};
test_output[440:440] = '{32'hc6bd6764};
test_input[3528:3535] = '{32'h41d464ee, 32'hbfe5a6e5, 32'hc141f056, 32'h425bccb0, 32'hc2a06120, 32'hc24f6b05, 32'h42296c9f, 32'h41ef83f5};
test_weights[3528:3535] = '{32'hc2aeb72c, 32'h429f5bdf, 32'hc1af701a, 32'h429d9654, 32'hc2936943, 32'hc2c7b538, 32'h4231fc69, 32'h42700338};
test_bias[441:441] = '{32'h42acc0e1};
test_output[441:441] = '{32'h4684ba39};
test_input[3536:3543] = '{32'h429f4c0f, 32'hc293e827, 32'hc27af1c5, 32'h42ad1c73, 32'h429ec9b5, 32'hc28a2260, 32'h3fe6f0de, 32'h41ff51c1};
test_weights[3536:3543] = '{32'hc2630a45, 32'hc22e471b, 32'h40b935c5, 32'h41934c3b, 32'h41c4a930, 32'hc2ba8849, 32'hc2a33ed6, 32'hc26f3056};
test_bias[442:442] = '{32'h427a7bf1};
test_output[442:442] = '{32'h45c5e0d1};
test_input[3544:3551] = '{32'h423f7332, 32'hc0870717, 32'h42460c13, 32'hc22c00cb, 32'h41d862f6, 32'hc20c70a4, 32'h42c066ac, 32'h40b833e3};
test_weights[3544:3551] = '{32'h4225055a, 32'h406d7d77, 32'h42b9bdc1, 32'hc11bc4e8, 32'h42253e7f, 32'hc29a8a46, 32'hc1373028, 32'h4297e807};
test_bias[443:443] = '{32'hc1eeba01};
test_output[443:443] = '{32'h461e0029};
test_input[3552:3559] = '{32'h413e7d39, 32'hc2b27306, 32'hc1b48aff, 32'hc2a73b79, 32'h42736130, 32'h42411334, 32'hc2ab1dac, 32'hc1b8596d};
test_weights[3552:3559] = '{32'h421fa0a0, 32'h42c656b0, 32'hc1ee22e5, 32'hc2a9b199, 32'h41887396, 32'hc2b5147e, 32'h4072f11d, 32'h41a9c120};
test_bias[444:444] = '{32'h428ffd5f};
test_output[444:444] = '{32'hc59248be};
test_input[3560:3567] = '{32'hc2329433, 32'h428c70cd, 32'hc2a368ae, 32'h41e22851, 32'h41bf4265, 32'hc1e88a55, 32'hc1f3a646, 32'h4166882a};
test_weights[3560:3567] = '{32'h3ff43aa8, 32'h4070bad1, 32'h4073e683, 32'hc1ea801e, 32'h42ac208a, 32'h42138865, 32'h42b1dcb5, 32'h41fab301};
test_bias[445:445] = '{32'hc2c276cd};
test_output[445:445] = '{32'hc5119d90};
test_input[3568:3575] = '{32'h42c564de, 32'h42c0148d, 32'h421c3156, 32'h42bba638, 32'h4262a19d, 32'hc09d82f3, 32'h41e53f2e, 32'h413d7cc2};
test_weights[3568:3575] = '{32'h42aafd1b, 32'hc1d13cad, 32'hbfaddf79, 32'hc174a2c9, 32'hc2ab8ef8, 32'hc1bd36f1, 32'h405c14c1, 32'hc276e7e8};
test_bias[446:446] = '{32'hc1906765};
test_output[446:446] = '{32'hc46ee88d};
test_input[3576:3583] = '{32'h428e62a9, 32'h4263de1f, 32'h40848d57, 32'h42116309, 32'h421b8298, 32'h42ac31f4, 32'h42003844, 32'hc2972195};
test_weights[3576:3583] = '{32'hc2b62416, 32'hc200604e, 32'hc1a818ab, 32'h420b8a5a, 32'hc26a9a43, 32'h42132ed6, 32'h422d22a4, 32'h429ff013};
test_bias[447:447] = '{32'hc2c2edb8};
test_output[447:447] = '{32'hc62bd000};
test_input[3584:3591] = '{32'hc11ddbc5, 32'hc2378b2d, 32'h423e734e, 32'hc253185c, 32'h4184e530, 32'hc2c28e61, 32'hc21e6615, 32'hbfaf70a8};
test_weights[3584:3591] = '{32'hc2afb897, 32'hc14e058f, 32'h423792f5, 32'hc2629698, 32'h420a4e10, 32'hc22e3aea, 32'h424b6c59, 32'h425fc953};
test_bias[448:448] = '{32'h3e3e3ad1};
test_output[448:448] = '{32'h461225ea};
test_input[3592:3599] = '{32'hc0b93e9a, 32'h40ab92e7, 32'h420d1280, 32'h4281b1b2, 32'hc2787cca, 32'h4260bb7a, 32'h42c36f14, 32'h41ae960a};
test_weights[3592:3599] = '{32'hc0d00a51, 32'h417ee3b5, 32'h425dd1a7, 32'hc25d7d74, 32'hc222d9b0, 32'hc288f8a8, 32'h41bf4f0c, 32'hc26a5b02};
test_bias[449:449] = '{32'hc244679c};
test_output[449:449] = '{32'hc4e3ae3b};
test_input[3600:3607] = '{32'hc0f72d32, 32'hc05225d5, 32'hc22c2ba4, 32'h42bde031, 32'h40e5d1a6, 32'h4228512d, 32'h4278a8a5, 32'h42c4edfe};
test_weights[3600:3607] = '{32'h42ac6c7d, 32'h425f792b, 32'hc2265b1c, 32'h42b23351, 32'hc24af362, 32'h429f1803, 32'h427b096f, 32'h42bbb3a5};
test_bias[450:450] = '{32'hc19f641e};
test_output[450:450] = '{32'h46c7422f};
test_input[3608:3615] = '{32'h42305415, 32'h3ebe5815, 32'h41e10d48, 32'hc13feac6, 32'hc23d57d2, 32'h42a49c5c, 32'hc2ac777f, 32'h4269e0a1};
test_weights[3608:3615] = '{32'hc237d0e3, 32'h424078dd, 32'hc2a3d469, 32'h41c14acd, 32'hc2aa7c23, 32'hc2376077, 32'hc2a7189b, 32'h429e0234};
test_bias[451:451] = '{32'h424830c9};
test_output[451:451] = '{32'h45eb6df1};
test_input[3616:3623] = '{32'h428e8226, 32'hc2b4dbef, 32'hc1db31b0, 32'hc2ae3697, 32'hc28841e1, 32'hc2c6f632, 32'hc2060e5f, 32'hc2c30935};
test_weights[3616:3623] = '{32'hc2a21448, 32'h42a6e3f0, 32'hc1dc33ff, 32'hc260a87c, 32'hc23d014e, 32'h420f522d, 32'h41c48022, 32'h41e5423b};
test_bias[452:452] = '{32'h419a2d4a};
test_output[452:452] = '{32'hc6358683};
test_input[3624:3631] = '{32'hc23d9951, 32'h426f8b9f, 32'hc2c7026d, 32'h425df213, 32'h4287a190, 32'h42491c44, 32'hc282a186, 32'h4134ee0c};
test_weights[3624:3631] = '{32'h4215304f, 32'hc1325618, 32'hc2c60c95, 32'hc24c7f68, 32'h4176d107, 32'h429c2f4f, 32'hc2bc0bce, 32'hc08ca1ee};
test_bias[453:453] = '{32'hc29db304};
test_output[453:453] = '{32'h4673397d};
test_input[3632:3639] = '{32'h420e59c0, 32'hc2036dcd, 32'h41f9f32b, 32'hc246e683, 32'hc2b1e1e3, 32'h42a7b7bb, 32'h41c215af, 32'h4224bc8d};
test_weights[3632:3639] = '{32'hc271f7a3, 32'h4273cf05, 32'h42c5452f, 32'hc299af5b, 32'hc171e7a8, 32'hc2c0b3d0, 32'h4286dd64, 32'hc14e769b};
test_bias[454:454] = '{32'h427eef22};
test_output[454:454] = '{32'hc5303b2d};
test_input[3640:3647] = '{32'hc274df14, 32'h42c2e2f4, 32'hc118991a, 32'hc2b7cf08, 32'h4220d527, 32'hc267cefe, 32'h424d5c1b, 32'hc21d130b};
test_weights[3640:3647] = '{32'h40e79a16, 32'h42c01910, 32'h423eb540, 32'hc2a5e96e, 32'hc2c70bd1, 32'hc2a980c5, 32'h422e0048, 32'hc23c4f65};
test_bias[455:455] = '{32'hc2715967};
test_output[455:455] = '{32'h46a43227};
test_input[3648:3655] = '{32'h429f3113, 32'h429f8eab, 32'h425bf2d7, 32'hc18c66d0, 32'h411c87c8, 32'h427a1574, 32'h423e03b3, 32'h423714bb};
test_weights[3648:3655] = '{32'h4203a375, 32'h419b3e5d, 32'h429167fa, 32'hc22ada4d, 32'h42b344d3, 32'hc2810241, 32'h41270add, 32'hc16ff00a};
test_bias[456:456] = '{32'h42b295d2};
test_output[456:456] = '{32'h45b0cee7};
test_input[3656:3663] = '{32'hc254e4fd, 32'hc1ea3208, 32'hc1c620fd, 32'h42b86d3c, 32'h407a4e5f, 32'h423805fa, 32'h42c327c8, 32'h42ab11c4};
test_weights[3656:3663] = '{32'hc2aab1c9, 32'hc1b9a77b, 32'hc10d5763, 32'h425f216d, 32'hc2582961, 32'h41019f54, 32'hc20121e4, 32'hc2c5049d};
test_bias[457:457] = '{32'h41f06ed8};
test_output[457:457] = '{32'hc4480652};
test_input[3664:3671] = '{32'hc1dd586f, 32'h4186bf33, 32'hc19b7df5, 32'h41f37b83, 32'hc21078fa, 32'h4231b8db, 32'hc24b7af3, 32'hc20f403f};
test_weights[3664:3671] = '{32'h41ab0428, 32'hc084f1ff, 32'hc24da0c6, 32'h4187f527, 32'h4143a73a, 32'h417a13eb, 32'h428a003c, 32'hc1427956};
test_bias[458:458] = '{32'hc2b396e4};
test_output[458:458] = '{32'hc5008d00};
test_input[3672:3679] = '{32'h41889c9f, 32'hc248f1d2, 32'h4292b30f, 32'h429576c0, 32'h41c3cc10, 32'h4272f601, 32'h420dcfe5, 32'hc1146e1b};
test_weights[3672:3679] = '{32'h427c1ac1, 32'h41e2548e, 32'h42946d47, 32'hc1e3433b, 32'hc289566d, 32'hc2af67a5, 32'h4283f3b2, 32'h4154f7e5};
test_bias[459:459] = '{32'h4209538a};
test_output[459:459] = '{32'hc4dec760};
test_input[3680:3687] = '{32'h421cadad, 32'h42aa4f6e, 32'h428c8f2e, 32'hbd52afda, 32'hc28bf37d, 32'h419d2b30, 32'hc273bb96, 32'h40a263ef};
test_weights[3680:3687] = '{32'hc2b9541f, 32'h40a0c791, 32'h42916986, 32'h3ecedad6, 32'h42a23686, 32'h4293379f, 32'hc1fd9545, 32'h42143d7c};
test_bias[460:460] = '{32'hc283c841};
test_output[460:460] = '{32'hc385e099};
test_input[3688:3695] = '{32'hc1832cdc, 32'hc2764388, 32'h42a53cb6, 32'h4220a8a2, 32'h4214e6b9, 32'hc2693a1f, 32'h4248a599, 32'h42ae8c70};
test_weights[3688:3695] = '{32'h410c5ddf, 32'hc09b329e, 32'h42182262, 32'h423545aa, 32'hc1a93a6d, 32'h429c1b57, 32'hc25a5350, 32'hc15d3039};
test_bias[461:461] = '{32'hc24f6064};
test_output[461:461] = '{32'hc583cc31};
test_input[3696:3703] = '{32'h41e07065, 32'hc286b95f, 32'hc2888063, 32'hc29740c2, 32'hc28cf98b, 32'hc230491a, 32'hc213518e, 32'hc0627023};
test_weights[3696:3703] = '{32'h41f952ee, 32'hc0b5dc0a, 32'hc2b04d78, 32'h42805258, 32'h4290ad02, 32'h428acdb0, 32'hc292f549, 32'h423a06d8};
test_bias[462:462] = '{32'hc2be98ac};
test_output[462:462] = '{32'hc54d9dec};
test_input[3704:3711] = '{32'h42b4289f, 32'hc20310f0, 32'hc2c0d6a6, 32'hc2c66edd, 32'hc0ee5cd5, 32'h42a74c5a, 32'h428e050a, 32'hc2c6c82a};
test_weights[3704:3711] = '{32'hc1fa50ad, 32'hc1f41b6b, 32'hc106b6a7, 32'h40e3bbbe, 32'hc1c3dee9, 32'hc289967a, 32'hc238da84, 32'hc2a6060a};
test_bias[463:463] = '{32'h427834a1};
test_output[463:463] = '{32'hc50ce18d};
test_input[3712:3719] = '{32'h42c21e93, 32'hbfd47df6, 32'h42462e9c, 32'h428d342e, 32'h429c6cd5, 32'h40e79168, 32'h424a6bd2, 32'h41efe175};
test_weights[3712:3719] = '{32'h41c53e72, 32'hc2126f8f, 32'h41c36d58, 32'hc254babc, 32'hc287f3ad, 32'h429367d9, 32'h42b40b50, 32'h42769e64};
test_bias[464:464] = '{32'hc15693bb};
test_output[464:464] = '{32'h44bda1b5};
test_input[3720:3727] = '{32'hc24df7aa, 32'hc138f853, 32'h427853ca, 32'h42526a39, 32'hc0cbd87b, 32'h417d6578, 32'hc29cbf68, 32'hc1f26d40};
test_weights[3720:3727] = '{32'hc2c45e2a, 32'hc2b71f0a, 32'hc271726a, 32'h420fde03, 32'h41ad6b43, 32'hc1d0f727, 32'hc0262e01, 32'hc2968486};
test_bias[465:465] = '{32'h4294adc0};
test_output[465:465] = '{32'h45c3cbad};
test_input[3728:3735] = '{32'hc2162c94, 32'hc2417d46, 32'h423b8bba, 32'h3ff694dc, 32'h41a9f564, 32'hc24618a1, 32'h41f9e348, 32'h40eba7bc};
test_weights[3728:3735] = '{32'h42b269ef, 32'hc2404fbb, 32'h42184d1d, 32'hc2449aa7, 32'hc2166d6f, 32'h40ed177d, 32'hc27b03a7, 32'hc18ccca9};
test_bias[466:466] = '{32'h426bf279};
test_output[466:466] = '{32'hc51e1a56};
test_input[3736:3743] = '{32'hc275b7bc, 32'h4090e029, 32'h429a1220, 32'h41fe0b48, 32'h40ceac18, 32'hc095826d, 32'hc24a0301, 32'h42a299ce};
test_weights[3736:3743] = '{32'hc2acc4f8, 32'hc256d6f1, 32'hc1e83f2a, 32'h41de6ce9, 32'h4257553d, 32'h41d82a01, 32'hc1dbdc2c, 32'h428c2e77};
test_bias[467:467] = '{32'h428783a3};
test_output[467:467] = '{32'h462d35cb};
test_input[3744:3751] = '{32'hc1732ea3, 32'h42c79313, 32'hc1f5a77b, 32'hbedfc0df, 32'hc208714d, 32'h428a8b42, 32'h419ba30b, 32'h4127550f};
test_weights[3744:3751] = '{32'h3ff63a56, 32'hc1067a11, 32'hc2c482fc, 32'h42a16634, 32'hc274fc03, 32'h420515c3, 32'hc266781d, 32'hc1bd5ac1};
test_bias[468:468] = '{32'h41e6f9fc};
test_output[468:468] = '{32'h45a181f2};
test_input[3752:3759] = '{32'hc29b759c, 32'hc1aeb696, 32'h416e3d22, 32'h41656025, 32'hc25242e4, 32'h419be3af, 32'h41e4d650, 32'h42658786};
test_weights[3752:3759] = '{32'hc21e864e, 32'hc29597d5, 32'hc1e22424, 32'h417e8b7c, 32'hc23fad24, 32'hbf234d75, 32'hc2289912, 32'h42b83b8f};
test_bias[469:469] = '{32'h4289293a};
test_output[469:469] = '{32'h462ea192};
test_input[3760:3767] = '{32'h42b15a3d, 32'hc24da311, 32'hc2a36155, 32'hc19d48a1, 32'hc2200c00, 32'h42ad7298, 32'hc216a341, 32'h42ab584a};
test_weights[3760:3767] = '{32'hc1e55cfb, 32'h4245470e, 32'hc293ab63, 32'hc26ddab5, 32'hc2c11b6e, 32'hc1a5995d, 32'h424383dc, 32'h41fdc896};
test_bias[470:470] = '{32'h41bb364d};
test_output[470:470] = '{32'h459f1aa6};
test_input[3768:3775] = '{32'hc210f668, 32'h423b893c, 32'h429d9afb, 32'hc2957e16, 32'hc2c7ac07, 32'hc2adb220, 32'h4201a494, 32'hc2bc6f52};
test_weights[3768:3775] = '{32'hc03ecd22, 32'hc1a85037, 32'hc297a694, 32'h42b61d9a, 32'h408c3234, 32'hc290345e, 32'h42a33a3e, 32'hc2801783};
test_bias[471:471] = '{32'hc1d0d3a3};
test_output[471:471] = '{32'h444c8061};
test_input[3776:3783] = '{32'hc2942af7, 32'hc274c97c, 32'hc205c4b7, 32'hc2a94d3a, 32'h428b2460, 32'h41d52b11, 32'h429a2c5b, 32'h41083bae};
test_weights[3776:3783] = '{32'hc2aa6c3b, 32'h42554b64, 32'hc22cfea1, 32'hc0f38004, 32'h42128249, 32'h41bab60c, 32'hc1dbe836, 32'h414c29a5};
test_bias[472:472] = '{32'hc1c38212};
test_output[472:472] = '{32'h45c41aa8};
test_input[3784:3791] = '{32'h422ee3b0, 32'h42737c1c, 32'h414ec1f6, 32'h4197c5aa, 32'hc2c644ce, 32'h4194b425, 32'hc25f1da8, 32'h4242db70};
test_weights[3784:3791] = '{32'h41a23c23, 32'h429fe814, 32'hc2947e52, 32'h414e255e, 32'h41b91136, 32'hc121f121, 32'h4241d698, 32'hc17036b4};
test_bias[473:473] = '{32'hc19389fe};
test_output[473:473] = '{32'hc45ff1ed};
test_input[3792:3799] = '{32'h421a68ec, 32'h41f09830, 32'h4214ef86, 32'hc21ced51, 32'h41f15451, 32'h42a3a222, 32'hc1c61d4a, 32'hc26e17bf};
test_weights[3792:3799] = '{32'hc281e6a0, 32'hc0b9e6b0, 32'h41b041f2, 32'h420fdcc3, 32'hc2c7d1b7, 32'hc2865040, 32'hc2657305, 32'hc2a72817};
test_bias[474:474] = '{32'h41d1bb46};
test_output[474:474] = '{32'hc5a77b82};
test_input[3800:3807] = '{32'h41df56fc, 32'h423a72c7, 32'h422ea459, 32'hc22c5e23, 32'h42505646, 32'hc0a46cc8, 32'h41b01101, 32'h42891767};
test_weights[3800:3807] = '{32'h417383da, 32'h41c2e43b, 32'hc1fabda2, 32'hc2c13303, 32'h4224f6c7, 32'h42a4d9ef, 32'hc2977be7, 32'hc2a3911f};
test_bias[475:475] = '{32'hc2388d8a};
test_output[475:475] = '{32'hc49afb39};
test_input[3808:3815] = '{32'hc2984abb, 32'h40b70936, 32'h42427bab, 32'h42873aa4, 32'hc0e9a045, 32'hc236d1c9, 32'h42ae3de4, 32'hc29f79c9};
test_weights[3808:3815] = '{32'h424ed56c, 32'hc2889f59, 32'h40ae0504, 32'h42bed3ff, 32'h429881aa, 32'hc1e015c0, 32'hc246ada9, 32'hc25df113};
test_bias[476:476] = '{32'h42ad3f23};
test_output[476:476] = '{32'h454ded42};
test_input[3816:3823] = '{32'h416af9a1, 32'hc29d97e2, 32'h42ad3f63, 32'h422e98f2, 32'h42bd90fa, 32'hc298597b, 32'h41bc8f59, 32'h427db2b0};
test_weights[3816:3823] = '{32'h4089dcc9, 32'h4200c0a5, 32'h4259021a, 32'h41ec4a02, 32'hc20117f8, 32'h421538c9, 32'h42c3c31f, 32'hc1b98f38};
test_bias[477:477] = '{32'hc216d99e};
test_output[477:477] = '{32'hc4c6592a};
test_input[3824:3831] = '{32'hc240eeb1, 32'h4296c390, 32'h4188fd06, 32'hc1890929, 32'hc1b37398, 32'hc22aa30d, 32'hc27e3a49, 32'h40462803};
test_weights[3824:3831] = '{32'hc1f2a097, 32'h42803c86, 32'hc2038842, 32'hc0fe3375, 32'h429d1bd3, 32'hc2832f07, 32'hc1b064f6, 32'hc0b95915};
test_bias[478:478] = '{32'h427edbeb};
test_output[478:478] = '{32'h46028175};
test_input[3832:3839] = '{32'hc24e0eda, 32'hc13c4205, 32'h4119a379, 32'hc2475f3e, 32'hc2a31fbb, 32'hc095bb9e, 32'hc2a9a1e3, 32'hc29d6322};
test_weights[3832:3839] = '{32'h420fce85, 32'hc282c1fc, 32'hc2b71ad9, 32'h42006ac5, 32'h422926e1, 32'hc2affd42, 32'h4172870e, 32'hc18cdb05};
test_bias[479:479] = '{32'h4222c8db};
test_output[479:479] = '{32'hc5c9d687};
test_input[3840:3847] = '{32'hc297ff34, 32'hc2bca45f, 32'h42b8f19e, 32'hc2a3b4f5, 32'h428fa19f, 32'h42892818, 32'h4294f04b, 32'h41bcadab};
test_weights[3840:3847] = '{32'h42c25250, 32'hc2963dab, 32'hc272379c, 32'h42bfdf1c, 32'h42609faa, 32'hc26d910a, 32'h426c97b6, 32'h428ff403};
test_bias[480:480] = '{32'h42c4f56a};
test_output[480:480] = '{32'hc5ed31c3};
test_input[3848:3855] = '{32'hc2a54ad8, 32'hc1886bcf, 32'hc27d88a9, 32'h42b49490, 32'h41c8f06e, 32'h4294e07a, 32'hc24c2ea7, 32'h42c5d5ef};
test_weights[3848:3855] = '{32'h42841a6d, 32'h416c42d3, 32'hc2417e03, 32'hc2a8fd38, 32'hc20fec9b, 32'h4084ee0e, 32'hc21814f3, 32'hc10a2a70};
test_bias[481:481] = '{32'hc0274667};
test_output[481:481] = '{32'hc618e103};
test_input[3856:3863] = '{32'hc26f61f5, 32'h42908b45, 32'hc27d9c99, 32'h4253f65d, 32'h420c6360, 32'h4222614a, 32'h424770e2, 32'h42b4973b};
test_weights[3856:3863] = '{32'h42a57324, 32'hc22b9bf0, 32'hc0bf11a1, 32'hc2373a40, 32'hc1f49a70, 32'h4265c563, 32'hc11eab10, 32'hc2bf5d5a};
test_bias[482:482] = '{32'h42354a10};
test_output[482:482] = '{32'hc68c1447};
test_input[3864:3871] = '{32'hc1eb5c60, 32'hc29ab81a, 32'hc2b5db56, 32'h40f4e439, 32'h40a4d98c, 32'hc1897109, 32'h420e1192, 32'hc2730ccc};
test_weights[3864:3871] = '{32'hc0d9e6d0, 32'hc2b04274, 32'h41612661, 32'h4212a2ad, 32'hc25853b2, 32'h41e3095b, 32'hc19572e7, 32'h4116dd42};
test_bias[483:483] = '{32'hc1206b50};
test_output[483:483] = '{32'h457a666e};
test_input[3872:3879] = '{32'hc2af863a, 32'h414bb695, 32'h429bb033, 32'hc26bdcbc, 32'h4279497b, 32'h41f607a7, 32'hbea053ce, 32'hc2813086};
test_weights[3872:3879] = '{32'h4186acc6, 32'h41e125e7, 32'hc19411ca, 32'hc00446cf, 32'hc1bf18a0, 32'h42b9a5e0, 32'hc2199f47, 32'hc2450fb6};
test_bias[484:484] = '{32'h4254ec1e};
test_output[484:484] = '{32'h4507f870};
test_input[3880:3887] = '{32'h4294c4f9, 32'h41fe6fbf, 32'h426a876c, 32'hc2a2739b, 32'hc202db93, 32'h42a2bc5c, 32'hc160d67b, 32'hc2a74b58};
test_weights[3880:3887] = '{32'hc196fbe2, 32'hc21d29ab, 32'hc19386ce, 32'h41af754c, 32'hc2a0fc34, 32'hc2996a19, 32'h42815896, 32'h42017762};
test_bias[485:485] = '{32'h42b76019};
test_output[485:485] = '{32'hc645a3a2};
test_input[3888:3895] = '{32'hc2b04887, 32'hc24b0a2d, 32'hc2ae7642, 32'h422bab89, 32'hc155bfbe, 32'h426eefdc, 32'h429288ba, 32'hc2b64268};
test_weights[3888:3895] = '{32'hc2c56651, 32'hc2c0b060, 32'hc23540ac, 32'hc289c16c, 32'hc25dc2f6, 32'h422fbc57, 32'hc2a7caf9, 32'h427bcd0c};
test_bias[486:486] = '{32'h41f28e83};
test_output[486:486] = '{32'h45be93ff};
test_input[3896:3903] = '{32'hc2706c76, 32'hc227cdc2, 32'hc2bb15af, 32'hc1f475f4, 32'h413261b5, 32'hc18352b5, 32'hc2b21320, 32'hc10c152b};
test_weights[3896:3903] = '{32'hc1d10ce3, 32'h4216cc75, 32'h4231b2e8, 32'h413763ad, 32'hc25b419c, 32'h42ad4769, 32'h4271844b, 32'hc2b2629d};
test_bias[487:487] = '{32'hc17faf47};
test_output[487:487] = '{32'hc62e649b};
test_input[3904:3911] = '{32'hc1557015, 32'hc00e6e58, 32'hc25e24ef, 32'h42abf942, 32'h429b29cc, 32'h42c129aa, 32'hc223eea4, 32'h427aaf90};
test_weights[3904:3911] = '{32'hc2bf2285, 32'h415f2914, 32'hc2bba4c7, 32'hc0772093, 32'h42aee5af, 32'hc12db035, 32'h42c6d933, 32'hc14a0f0f};
test_bias[488:488] = '{32'hc2b39454};
test_output[488:488] = '{32'h45d7b25d};
test_input[3912:3919] = '{32'hc13d87c9, 32'h42261614, 32'hc1c44593, 32'h42ac10b5, 32'hc233007d, 32'h3ffe5070, 32'h41c5c536, 32'h42a1c7f6};
test_weights[3912:3919] = '{32'h427eccd0, 32'h425cf58d, 32'hc1aeaede, 32'h423743ea, 32'h41b94b7b, 32'hc10ffbe9, 32'h42ab0910, 32'hc2934f5d};
test_bias[489:489] = '{32'h41b6d4bc};
test_output[489:489] = '{32'h448ea221};
test_input[3920:3927] = '{32'hc12b6087, 32'hc2826263, 32'h4283461f, 32'hc2479f73, 32'h42bbce4e, 32'h41565305, 32'h416806b5, 32'hc1c26f3f};
test_weights[3920:3927] = '{32'hc1e8a7a5, 32'hc255cc00, 32'hc22759f7, 32'h4283951e, 32'hc0857754, 32'h4146dac0, 32'hc14885c7, 32'hc2a6ba12};
test_bias[490:490] = '{32'h42752e56};
test_output[490:490] = '{32'hc40a41cf};
test_input[3928:3935] = '{32'hc261b86c, 32'hc2550107, 32'h42722448, 32'hc25071f5, 32'h41c39a75, 32'hc2587dd2, 32'h4284277f, 32'hc22b514d};
test_weights[3928:3935] = '{32'h42b44b34, 32'hc223a9fc, 32'hc25ba85a, 32'h42c49f9d, 32'h42b06588, 32'h41177c72, 32'hc2afbb6c, 32'hc2ac0fd5};
test_bias[491:491] = '{32'hc2a9f882};
test_output[491:491] = '{32'hc63a3741};
test_input[3936:3943] = '{32'h42c3f990, 32'h424de178, 32'hc1763811, 32'hc2b787c9, 32'hc04cd855, 32'h428a712e, 32'hc1ac1082, 32'hc1b0bcb2};
test_weights[3936:3943] = '{32'hc1990c04, 32'h41e25a88, 32'h40a36e9f, 32'hc1f73d8a, 32'hc1f4603f, 32'h41bb8e95, 32'h41e21c03, 32'h41e5eaef};
test_bias[492:492] = '{32'hc2932cb8};
test_output[492:492] = '{32'h452b75d6};
test_input[3944:3951] = '{32'hc250d5e2, 32'hc22ae956, 32'h428a5153, 32'h4153a35b, 32'h4136cc50, 32'h42b79264, 32'h40b7127c, 32'h41965c64};
test_weights[3944:3951] = '{32'hc292f3c6, 32'hc23ce4f9, 32'h41a56cb1, 32'hc28553c7, 32'h423c965c, 32'hc241ceb4, 32'h42b65547, 32'hc10f5658};
test_bias[493:493] = '{32'hc1d64c5e};
test_output[493:493] = '{32'h4530400d};
test_input[3952:3959] = '{32'hbe79e518, 32'hc2a70951, 32'h4225f772, 32'h3ff695d0, 32'hc1a0173d, 32'hc28f3c12, 32'h419575a0, 32'hc21cdc00};
test_weights[3952:3959] = '{32'h42071032, 32'h3fe0f5a4, 32'hc26316ca, 32'h418d0c93, 32'hc14adc1c, 32'hc299d2be, 32'hc2a31686, 32'hc29c159e};
test_bias[494:494] = '{32'hc29bafef};
test_output[494:494] = '{32'h4594435b};
test_input[3960:3967] = '{32'h4251e295, 32'hc21d656a, 32'h41a7573b, 32'hc1ac03a6, 32'h42a39d96, 32'h422451a3, 32'h40d79a37, 32'hc28e7a08};
test_weights[3960:3967] = '{32'hc0f8765f, 32'h426b60ea, 32'h4014fe8e, 32'h409597c5, 32'h42a7dd34, 32'hc071e2c6, 32'hc1eed66b, 32'h42b0fd10};
test_bias[495:495] = '{32'hc273b472};
test_output[495:495] = '{32'hc5245ef3};
test_input[3968:3975] = '{32'hc04ebb15, 32'hc2bd2512, 32'hc238057b, 32'hc290ecd6, 32'h42a434ff, 32'h42541b9f, 32'hc0f752d0, 32'h42ae8b52};
test_weights[3968:3975] = '{32'hc2063b02, 32'hc2b3dd14, 32'h4281b5d4, 32'h4240ed30, 32'hc295ad62, 32'hc2436a5c, 32'h41d5d9ea, 32'h42c01473};
test_bias[496:496] = '{32'hc27bad7b};
test_output[496:496] = '{32'h44bcf944};
test_input[3976:3983] = '{32'hc2a45f33, 32'h421a9ab0, 32'hc17ead77, 32'hc242bb5c, 32'hc2891d2c, 32'hc12e6f2a, 32'h421985e8, 32'hbf993c28};
test_weights[3976:3983] = '{32'h4148180d, 32'h429069e2, 32'h40d620ee, 32'h42243d50, 32'h4285c17f, 32'hc2a86211, 32'hc2c6b606, 32'hc1138a57};
test_bias[497:497] = '{32'h4265aa53};
test_output[497:497] = '{32'hc5f252a4};
test_input[3984:3991] = '{32'h42537158, 32'hc1b00872, 32'h4288e094, 32'hc28ffabf, 32'h427e0731, 32'h42a7d771, 32'hc2b52798, 32'hc1aa7f80};
test_weights[3984:3991] = '{32'hc1bcc8fd, 32'h4215e764, 32'hc2546226, 32'hc2b3580d, 32'h41a19b07, 32'h4180074a, 32'h41a5a57b, 32'h4194eb39};
test_bias[498:498] = '{32'hc0b4d16b};
test_output[498:498] = '{32'h448935ca};
test_input[3992:3999] = '{32'h4294f567, 32'h42356b68, 32'hc28e710f, 32'hc2257257, 32'h4204dbc7, 32'hc1a8248d, 32'hc28cd3c8, 32'hc1c08565};
test_weights[3992:3999] = '{32'h427a11fb, 32'h4218a2ca, 32'hc29a4990, 32'hc0fd304e, 32'hc236227b, 32'h4258e1cc, 32'h421665ab, 32'h4253b0b4};
test_bias[499:499] = '{32'h429331e2};
test_output[499:499] = '{32'h45b267d7};
test_input[4000:4007] = '{32'hc28cdae7, 32'h42bcc1aa, 32'h4248d972, 32'h42a47d9c, 32'h4159d33a, 32'hc230d568, 32'h41a7a441, 32'h4238586b};
test_weights[4000:4007] = '{32'h3f2e1376, 32'h418dfd5e, 32'h421e7504, 32'hc28ce4e5, 32'hc175a4bf, 32'hc29e832b, 32'h4007cb05, 32'h428f34a0};
test_bias[500:500] = '{32'h4284a2d8};
test_output[500:500] = '{32'h458d7ed4};
test_input[4008:4015] = '{32'h428eda82, 32'h41cf8d04, 32'hc2369371, 32'h4252d170, 32'h420f9ec9, 32'hc25d9d79, 32'h41220733, 32'h424060c3};
test_weights[4008:4015] = '{32'hc299b755, 32'hc12d4080, 32'h42c621d1, 32'hc2b2d1d4, 32'h41c58e64, 32'h41fa0afc, 32'hc24ec109, 32'h42646dfa};
test_bias[501:501] = '{32'h428b9c77};
test_output[501:501] = '{32'hc653d33c};
test_input[4016:4023] = '{32'h42515cfa, 32'h41451b0e, 32'h418170c9, 32'h42022543, 32'hc2c006fd, 32'hc10d57df, 32'h42b56f64, 32'hc1580f09};
test_weights[4016:4023] = '{32'hc16167ee, 32'hc29f9b34, 32'h41376ab6, 32'hc29958f6, 32'h4246a017, 32'hc28f031a, 32'h427f3639, 32'hc22cdaca};
test_bias[502:502] = '{32'h429050bd};
test_output[502:502] = '{32'hc4d73def};
test_input[4024:4031] = '{32'hc16e03e5, 32'hc1514062, 32'hc29996cf, 32'hc2325d18, 32'hc21182c5, 32'hc2c7d8bc, 32'h42bd0a1e, 32'hc2b46317};
test_weights[4024:4031] = '{32'hc2a4565a, 32'h42a2fe8f, 32'h42904e30, 32'hc1af0443, 32'h424f6de7, 32'hc21f4a92, 32'hc257581a, 32'h425ec71d};
test_bias[503:503] = '{32'h424a5331};
test_output[503:503] = '{32'hc64165a0};
test_input[4032:4039] = '{32'hc259b71d, 32'h42266bf5, 32'hc2c19061, 32'h426ffd36, 32'h42166bde, 32'hc2845a32, 32'hc288345e, 32'h42c782ca};
test_weights[4032:4039] = '{32'h42c5d71e, 32'hc2b11223, 32'h429cff85, 32'hc1e321ed, 32'h42091ae8, 32'hc082fc69, 32'hc2a7795b, 32'h422d68c5};
test_bias[504:504] = '{32'h42a0f284};
test_output[504:504] = '{32'hc5d165e8};
test_input[4040:4047] = '{32'hc24539ce, 32'h428887e4, 32'h420e1216, 32'h42843fa7, 32'h4172bb3c, 32'hc2b1c33b, 32'h42020847, 32'h41b31025};
test_weights[4040:4047] = '{32'hc29f9ebe, 32'h41ae3543, 32'h42ab0d59, 32'h424785c7, 32'hc20bc9c7, 32'h42935c7e, 32'h41b42051, 32'h40a290f1};
test_bias[505:505] = '{32'hc17910c3};
test_output[505:505] = '{32'h45ac2654};
test_input[4048:4055] = '{32'h423c5d14, 32'hc2bfa228, 32'h4130e027, 32'hc2c4bda4, 32'hc28c2dcf, 32'hc1c70c79, 32'hc08e473f, 32'hc2053210};
test_weights[4048:4055] = '{32'hc20b79f8, 32'h42bfa1ab, 32'hc2ac087d, 32'hc0050d3d, 32'h42026142, 32'hc28cea22, 32'hc0a3690e, 32'h4278b1d8};
test_bias[506:506] = '{32'h429fb527};
test_output[506:506] = '{32'hc65bd1ad};
test_input[4056:4063] = '{32'h42a45381, 32'h42ae9e7e, 32'hc2a510f5, 32'hc203348b, 32'h426307ff, 32'hc235b872, 32'h4223bc5b, 32'h413f6a96};
test_weights[4056:4063] = '{32'h425a7e97, 32'h41c261f8, 32'h429e4ccc, 32'hc146fc91, 32'h427c4675, 32'h411142f6, 32'h40a4bd5f, 32'h40dbbb99};
test_bias[507:507] = '{32'hc25bc202};
test_output[507:507] = '{32'h457320f1};
test_input[4064:4071] = '{32'hc1740ed2, 32'h4259d7f6, 32'hc2425fd6, 32'hc298bf5b, 32'hc237ccdc, 32'hc298892d, 32'h428100e6, 32'hc20844a8};
test_weights[4064:4071] = '{32'h42812da1, 32'hc1a48696, 32'hc28de896, 32'hc2b7e057, 32'hc20ec53a, 32'hc1f2b1bd, 32'hbff3217f, 32'h41b2d694};
test_bias[508:508] = '{32'h426e356c};
test_output[508:508] = '{32'h46339674};
test_input[4072:4079] = '{32'hc1c9a3ef, 32'hc28d4b23, 32'h42a92eb6, 32'hc20befb4, 32'h428aff62, 32'h42579fa9, 32'hc0c37926, 32'h41c157fe};
test_weights[4072:4079] = '{32'h42c25e2b, 32'h422cf362, 32'hc1979e4c, 32'h4206a8fa, 32'hc246fbe8, 32'h425d48ab, 32'hc27f1ce7, 32'h427b840d};
test_bias[509:509] = '{32'h42b4bb94};
test_output[509:509] = '{32'hc5d344e1};
test_input[4080:4087] = '{32'hc0404036, 32'h41f0d8ce, 32'hc2349ca1, 32'h41d95be1, 32'h3f65a950, 32'h42c21782, 32'hc23ab0bb, 32'h4196b15f};
test_weights[4080:4087] = '{32'h41faa8e6, 32'h420f1024, 32'hc1a52358, 32'h419a3dd3, 32'h42c03313, 32'h41a4f4ee, 32'hc1d7dbd6, 32'hc281b77b};
test_bias[510:510] = '{32'h4094a2e7};
test_output[510:510] = '{32'h458ec089};
test_input[4088:4095] = '{32'hc2bddafc, 32'h3fb1f045, 32'hc185a0d3, 32'h419dba35, 32'h4252e479, 32'hbf2cd4fd, 32'hc1e91059, 32'h41cb346b};
test_weights[4088:4095] = '{32'h4180f36b, 32'hc26f2cf2, 32'hc267b22e, 32'h425eaf0f, 32'h428eec6a, 32'hc2bf8416, 32'h42a393e2, 32'h4140f9dc};
test_bias[511:511] = '{32'hc2b35a70};
test_output[511:511] = '{32'h45046272};
test_input[4096:4103] = '{32'h42b60f93, 32'hc2046381, 32'hc2ab8c75, 32'hc2b97943, 32'hc24c2068, 32'h3fb83173, 32'h42381621, 32'h4022bd6c};
test_weights[4096:4103] = '{32'h4094f4ae, 32'hc28caecb, 32'hc24b154f, 32'h420808d1, 32'h4276f1f5, 32'h420e7952, 32'h4292673b, 32'hc1e2cec5};
test_bias[512:512] = '{32'h427e32c4};
test_output[512:512] = '{32'h4583af10};
test_input[4104:4111] = '{32'h42be2baa, 32'h428588ac, 32'h406e3f39, 32'hc1439334, 32'h42897331, 32'hc24be49c, 32'hc29554e8, 32'h42a98a79};
test_weights[4104:4111] = '{32'h4134dd8d, 32'h40a29a18, 32'hc2947041, 32'h416abfa2, 32'h4162d431, 32'h429ad70f, 32'hc16604e7, 32'h42512d50};
test_bias[513:513] = '{32'hc1fe0a9e};
test_output[513:513] = '{32'h45585199};
test_input[4112:4119] = '{32'h4294d538, 32'h4295ba64, 32'hc1409b88, 32'h428614b8, 32'h42baa8e8, 32'h426024ca, 32'hc14c6df9, 32'hc1308441};
test_weights[4112:4119] = '{32'h42b07378, 32'hc1c4b37a, 32'hc25e69b0, 32'hc2255c19, 32'hc2807dd9, 32'h4070cb9d, 32'h41135171, 32'hc29d2965};
test_bias[514:514] = '{32'h418d0d58};
test_output[514:514] = '{32'hc515bb46};
test_input[4120:4127] = '{32'h42834c14, 32'h4177774d, 32'hc2165523, 32'h41fd99f8, 32'h42bac11f, 32'h4180bc56, 32'hc2b47e8a, 32'hc286c67f};
test_weights[4120:4127] = '{32'hc1c91e17, 32'h4151c510, 32'hc28a5c62, 32'h42217132, 32'hc2b3bab5, 32'h4261451b, 32'h42b61dab, 32'h41e1038a};
test_bias[515:515] = '{32'h42000571};
test_output[515:515] = '{32'hc66c7941};
test_input[4128:4135] = '{32'h41f4140b, 32'h41c94231, 32'hc20190c0, 32'hc268e13d, 32'h42b4963c, 32'h42159d97, 32'h4212aa8a, 32'h414e2175};
test_weights[4128:4135] = '{32'h4255af03, 32'h420813d4, 32'hc286168e, 32'h4290f7eb, 32'h3ddb57da, 32'hc2c6fb1f, 32'hc296e2f5, 32'hc2b2c1de};
test_bias[516:516] = '{32'hc1949798};
test_output[516:516] = '{32'hc5e15525};
test_input[4136:4143] = '{32'hbeef426c, 32'hc2c1180e, 32'hc1f9706c, 32'hc1f71ebc, 32'hc218b9fd, 32'hc1a7e1ec, 32'h42ae53fb, 32'hc1c1f812};
test_weights[4136:4143] = '{32'hc281184f, 32'hc2a4b832, 32'hc1853cef, 32'h41904b27, 32'hc2a4daeb, 32'h41d7bedf, 32'hc1c07dfe, 32'hc290153d};
test_bias[517:517] = '{32'hc2003f14};
test_output[517:517] = '{32'h461e7a27};
test_input[4144:4151] = '{32'hc19cdc41, 32'h429913d4, 32'h4174b297, 32'h42694496, 32'hc1314505, 32'hc19f305e, 32'h402b6371, 32'h42a7e461};
test_weights[4144:4151] = '{32'hc24b9fc5, 32'h42b27eb6, 32'hc2a419d8, 32'h42a73a3f, 32'hc2307cf5, 32'h42511bb8, 32'h41d7a4cc, 32'h42a85fd0};
test_bias[518:518] = '{32'h42baae88};
test_output[518:518] = '{32'h468da72f};
test_input[4152:4159] = '{32'h427facf2, 32'hc2b9ddc5, 32'hc28c694b, 32'h42488f01, 32'hc2a3f309, 32'hc1b41c7e, 32'hc28bb336, 32'hc11ca269};
test_weights[4152:4159] = '{32'hc113bdbb, 32'h3fb9bc96, 32'hc292e10e, 32'h428734c6, 32'h42ae9c01, 32'h41f64ef9, 32'h423f0438, 32'h42b98608};
test_bias[519:519] = '{32'h4150b412};
test_output[519:519] = '{32'hc58521e0};
test_input[4160:4167] = '{32'hc23c7684, 32'hc189488e, 32'h41e51781, 32'h41ac9e22, 32'h428d673b, 32'h422cb2cf, 32'h42bdf581, 32'h42b6a39d};
test_weights[4160:4167] = '{32'hc2b5ee4b, 32'hc19846b7, 32'hc09d41bb, 32'h4208705d, 32'h41e5b2dc, 32'hc29aa52a, 32'h41292b1d, 32'hbbb36340};
test_bias[520:520] = '{32'hc295d401};
test_output[520:520] = '{32'h4596e202};
test_input[4168:4175] = '{32'h42c43fd4, 32'hc2aa4c49, 32'hc1b50732, 32'h41cc299a, 32'hc286a084, 32'h4202ccc9, 32'hc2bc2edd, 32'h4297620b};
test_weights[4168:4175] = '{32'h42876b09, 32'h415cae8d, 32'h42960978, 32'hc281d30d, 32'hc1c68c9e, 32'h42995e71, 32'h42892c9f, 32'h42c543ce};
test_bias[521:521] = '{32'hc08878df};
test_output[521:521] = '{32'h45e42bd1};
test_input[4176:4183] = '{32'hc1212628, 32'h4224b300, 32'hc1a662c3, 32'hc10f7cf3, 32'h4189ec9c, 32'h41cb4065, 32'hc1e0552a, 32'hc237497f};
test_weights[4176:4183] = '{32'h4287e58b, 32'h41daff81, 32'h42afba56, 32'hc27b6de6, 32'hc23c2440, 32'h4247b3b1, 32'hc2ae22df, 32'hc2ac3be3};
test_bias[522:522] = '{32'hc2225661};
test_output[522:522] = '{32'h45bafc8a};
test_input[4184:4191] = '{32'hc1ab123a, 32'h41d77544, 32'h428af7f1, 32'hc113d661, 32'h4206018d, 32'hc163b9b9, 32'hc1c61d9c, 32'hc0c78af4};
test_weights[4184:4191] = '{32'hc280a614, 32'hc25c7dd2, 32'hc1f2afbd, 32'hc29c7161, 32'h4240f609, 32'h425cc510, 32'h40b63273, 32'hc1de80b6};
test_bias[523:523] = '{32'hc2b80054};
test_output[523:523] = '{32'hc434cb54};
test_input[4192:4199] = '{32'hc293dc34, 32'hc2472068, 32'hc1e28dff, 32'h422b618c, 32'h42b43a6e, 32'hc295822a, 32'hc2afd62e, 32'h401a1d5d};
test_weights[4192:4199] = '{32'h403e1327, 32'hc1fb56ba, 32'h426158d2, 32'hbf82aa24, 32'hc176751c, 32'hc0ebedb0, 32'hc22ece0d, 32'h421467e5};
test_bias[524:524] = '{32'hc26a45fe};
test_output[524:524] = '{32'h452b542c};
test_input[4200:4207] = '{32'hc14f03f3, 32'h416c3c14, 32'hc240ce39, 32'h4253c0f0, 32'hc1841ba5, 32'h4256d393, 32'hc2239e19, 32'hc196da80};
test_weights[4200:4207] = '{32'h42945e85, 32'h41f8ae32, 32'hc29a6d6e, 32'h4216eaa9, 32'h428eb763, 32'hc26433b1, 32'hc248066a, 32'hc29fc04d};
test_bias[525:525] = '{32'h420ab59a};
test_output[525:525] = '{32'h458e91e7};
test_input[4208:4215] = '{32'h4276eb4c, 32'h414b795c, 32'h42ba9202, 32'h4278d273, 32'hc2a28f0f, 32'h4254a21a, 32'h41e1cc31, 32'hbfd8e22c};
test_weights[4208:4215] = '{32'h41a45e58, 32'h4297f4ef, 32'hbf288672, 32'hc20646c5, 32'h4206290a, 32'h42849809, 32'h3fe1ab09, 32'h4250060b};
test_bias[526:526] = '{32'h420ac5a0};
test_output[526:526] = '{32'h445bd8d1};
test_input[4216:4223] = '{32'h42adbe96, 32'h424bde18, 32'hc2008bc0, 32'hc2c57b4c, 32'h42c36f1a, 32'hc20e9d92, 32'hc219eb39, 32'h422945c8};
test_weights[4216:4223] = '{32'h4266d8f5, 32'h429b5ebc, 32'h4265d04b, 32'hc2c0ec1f, 32'hc25fed51, 32'h42c1e65e, 32'h4253ad76, 32'hc29c798e};
test_bias[527:527] = '{32'h42b883ae};
test_output[527:527] = '{32'h451a54a8};
test_input[4224:4231] = '{32'hc1361284, 32'hc227d277, 32'h42a2525d, 32'hc1c43bc2, 32'hc2b192e7, 32'h41bb5fb3, 32'hc2be1a34, 32'h412a2252};
test_weights[4224:4231] = '{32'h4282363f, 32'hc2414c9d, 32'hc297393e, 32'hc2ac73e6, 32'hc2a3cda1, 32'h423673e3, 32'h420dc055, 32'h42b1e31e};
test_bias[528:528] = '{32'h4223fa2d};
test_output[528:528] = '{32'h4549773a};
test_input[4232:4239] = '{32'hc2990bbb, 32'h427a9c1e, 32'h423eb551, 32'h411fd802, 32'hc2a531d6, 32'h4031125b, 32'hc0ecd4b3, 32'hc152520e};
test_weights[4232:4239] = '{32'hbf2acf21, 32'h412d3618, 32'h42bb242c, 32'h429fff1b, 32'h421e79a3, 32'h42596834, 32'hc2bafb8f, 32'h4192816c};
test_bias[529:529] = '{32'hc299690a};
test_output[529:529] = '{32'h454aa27a};
test_input[4240:4247] = '{32'hc21f3931, 32'hc21d8f92, 32'hc1703653, 32'h4209325a, 32'h41edd119, 32'hc255de89, 32'hc29c44f6, 32'hc2b41ad0};
test_weights[4240:4247] = '{32'hc2296035, 32'hc098ee41, 32'hc2a73bd3, 32'h41bac426, 32'hc267d639, 32'h420c39f2, 32'hc27fcffe, 32'h42a1ef24};
test_bias[530:530] = '{32'hc2952f63};
test_output[530:530] = '{32'hc4fe8ba6};
test_input[4248:4255] = '{32'hc1eec815, 32'hbf60db89, 32'h42483e65, 32'h427eeec3, 32'h421db7aa, 32'h42a28f12, 32'h419e9e5e, 32'hc2592886};
test_weights[4248:4255] = '{32'h4220e315, 32'hc060b792, 32'hc11478e3, 32'hc2c0828a, 32'h41a72b92, 32'hc205d16f, 32'hc2972ab4, 32'hc1432fff};
test_bias[531:531] = '{32'h410c8e36};
test_output[531:531] = '{32'hc6245d97};
test_input[4256:4263] = '{32'hc2997302, 32'hc09acf4a, 32'h42448fc2, 32'h4282ab96, 32'h42a5b157, 32'h429d97cd, 32'h42a71a27, 32'h42973408};
test_weights[4256:4263] = '{32'hc1ae0872, 32'hc2b4d4e2, 32'hc2b7d29f, 32'hc2c35ce0, 32'hc2625111, 32'hc2848f00, 32'h42924d54, 32'hc26c9f19};
test_bias[532:532] = '{32'hc2928502};
test_output[532:532] = '{32'hc685df69};
test_input[4264:4271] = '{32'h428438c1, 32'h41318b5c, 32'h421cc592, 32'h420ad27e, 32'h42a3e576, 32'h42ab9a2f, 32'hc1a642a6, 32'hc29f4a9f};
test_weights[4264:4271] = '{32'h41897e9c, 32'hc21eccbe, 32'hc1ec9993, 32'hc18528d5, 32'hc03ad8e4, 32'h421a8622, 32'h42b4b98d, 32'h4217ef27};
test_bias[533:533] = '{32'hc1e0285b};
test_output[533:533] = '{32'hc5350f88};
test_input[4272:4279] = '{32'h421d15b8, 32'hc2578659, 32'h42bfe34e, 32'h4109ca3f, 32'hc20845cf, 32'hc1461668, 32'h42634bbc, 32'hc2377072};
test_weights[4272:4279] = '{32'hc29f3940, 32'hc29eb802, 32'hc1cda150, 32'hc29ab4ea, 32'h4231fdbe, 32'hc2799177, 32'h409f1ed3, 32'h426fa774};
test_bias[534:534] = '{32'h4250f692};
test_output[534:534] = '{32'hc5a098bc};
test_input[4280:4287] = '{32'hc2a1a872, 32'hbf380d04, 32'h42abf1f4, 32'h423d84cd, 32'h42871de0, 32'h42729954, 32'h41a2d998, 32'h42b91e25};
test_weights[4280:4287] = '{32'hc28a99b3, 32'h4173e271, 32'hc228861b, 32'h41759485, 32'hc0d59a38, 32'h4267df2f, 32'hc2349235, 32'h40e7b2f6};
test_bias[535:535] = '{32'h42574f46};
test_output[535:535] = '{32'h45adebca};
test_input[4288:4295] = '{32'hc2a26042, 32'hc29a6fab, 32'hc1fc9604, 32'h42424803, 32'hc2089572, 32'hc136ad7f, 32'h427bb48f, 32'h421afd96};
test_weights[4288:4295] = '{32'hc22a8fcf, 32'h42ac9a65, 32'hc243bf41, 32'h42c6000f, 32'hc25d68fa, 32'hc015af4f, 32'h42c7936e, 32'hc2bdf8a3};
test_bias[536:536] = '{32'hc2a2983d};
test_output[536:536] = '{32'h45ed0d9a};
test_input[4296:4303] = '{32'hc2909f00, 32'h419e0c2f, 32'hc25b4da1, 32'h419f071c, 32'h4234db50, 32'h419c64de, 32'h4293c6cb, 32'hc13fdebd};
test_weights[4296:4303] = '{32'h40d1b4ec, 32'hc2bceb96, 32'h41a5a1c8, 32'h4146c09c, 32'h41c77bdf, 32'hc2c26504, 32'hc2b0a5de, 32'h41ad7561};
test_bias[537:537] = '{32'h4292c416};
test_output[537:537] = '{32'hc627668d};
test_input[4304:4311] = '{32'h42b83a95, 32'hc29e7d97, 32'hc2b623fa, 32'h428faa1c, 32'h42a290dd, 32'h41ccd9c3, 32'hc25f71ec, 32'h4132a52c};
test_weights[4304:4311] = '{32'h42606c76, 32'hc293c481, 32'h41aa1b18, 32'h424e7462, 32'hc2205b69, 32'hc2a023b5, 32'h41fcac57, 32'hc1e46dcb};
test_bias[538:538] = '{32'hc2920c45};
test_output[538:538] = '{32'h45a6893b};
test_input[4312:4319] = '{32'hc2ab4b2e, 32'h42852893, 32'h42168de9, 32'h428df1a4, 32'hc20044a6, 32'h40d5069c, 32'hc180f1c3, 32'hc1caca4b};
test_weights[4312:4319] = '{32'h42735872, 32'hc20e0d95, 32'h42a3918d, 32'h42913628, 32'hc2857fd9, 32'hc20b488c, 32'h40796a53, 32'h41c1790a};
test_bias[539:539] = '{32'h42810390};
test_output[539:539] = '{32'h44f434ad};
test_input[4320:4327] = '{32'hc2142b21, 32'hc26bfb75, 32'hc16ebcc3, 32'h42207274, 32'h42bbec03, 32'hc2581a99, 32'hc21fd97d, 32'hc28be6a7};
test_weights[4320:4327] = '{32'h42ad2861, 32'hc1b19737, 32'h42c60290, 32'h42b48210, 32'h3f2b2fa9, 32'hc2570232, 32'h4253d7c1, 32'h42462d51};
test_bias[540:540] = '{32'h42b31e11};
test_output[540:540] = '{32'hc50e81fc};
test_input[4328:4335] = '{32'hc2bd504b, 32'h4140897a, 32'h42769793, 32'hc2607770, 32'hc273267d, 32'h4053f115, 32'h40a59926, 32'hc27d2cd4};
test_weights[4328:4335] = '{32'hc23083b4, 32'h4287925a, 32'hc2c12b42, 32'hc239dbd0, 32'hc2399a16, 32'hc2c13c19, 32'h4229c29a, 32'hc2c5fa7f};
test_bias[541:541] = '{32'h4124e769};
test_output[541:541] = '{32'h462647b7};
test_input[4336:4343] = '{32'hc2250bf7, 32'h41412e55, 32'h42987655, 32'hc2b7cb81, 32'hc2542d31, 32'hc2bc6b67, 32'h4100b170, 32'h427c8fd1};
test_weights[4336:4343] = '{32'h41bd26ac, 32'hc1bf00d4, 32'h40a50ed0, 32'h4193729e, 32'hc06f85e7, 32'h42624936, 32'h41dd0131, 32'hc1e23acb};
test_bias[542:542] = '{32'hc202fea4};
test_output[542:542] = '{32'hc6112e36};
test_input[4344:4351] = '{32'h424c8624, 32'h40ab669e, 32'h41f5f721, 32'h41d2c7a4, 32'h4284662c, 32'h42201dfd, 32'h42892e33, 32'hc2c2887e};
test_weights[4344:4351] = '{32'h4203d84c, 32'hc27cb599, 32'hc2acadae, 32'h42bf8eeb, 32'h400f512f, 32'hc26159a1, 32'h41f3906d, 32'hc24a461e};
test_bias[543:543] = '{32'h423fe91e};
test_output[543:543] = '{32'h45c09f14};
test_input[4352:4359] = '{32'h42043dac, 32'hc282479f, 32'hc20e7a6e, 32'h42c3f15c, 32'hbfc1ecc8, 32'h42bf7da6, 32'hc2b9565b, 32'h4249755a};
test_weights[4352:4359] = '{32'h4207355d, 32'hc2092fa5, 32'h42851695, 32'h4235dd2f, 32'hc2864810, 32'hc2925ddf, 32'h41c67c5d, 32'hc2a18219};
test_bias[544:544] = '{32'hc2be79c7};
test_output[544:544] = '{32'hc5f7d919};
test_input[4360:4367] = '{32'hc2b29c0e, 32'h418811a6, 32'h427b4539, 32'h42aef875, 32'h42c1d6cf, 32'hc1dbcfbd, 32'hc1a837e6, 32'hc17546b2};
test_weights[4360:4367] = '{32'hc1877a09, 32'hc222296a, 32'hc136030e, 32'hc24f4343, 32'hc11690d2, 32'h42560203, 32'hc2c4fc0e, 32'hc205a3ad};
test_bias[545:545] = '{32'h4293600e};
test_output[545:545] = '{32'hc581b0ec};
test_input[4368:4375] = '{32'hc2241212, 32'hc2b88f66, 32'hc2298efd, 32'h421d8672, 32'hc2894ded, 32'hc240e48e, 32'h429ada79, 32'h425e63f4};
test_weights[4368:4375] = '{32'hc2925aba, 32'h42905d76, 32'h42295332, 32'hc2c74218, 32'h42002333, 32'hc29f4e8b, 32'h41dd2c9e, 32'h41179a98};
test_bias[546:546] = '{32'h4235104c};
test_output[546:546] = '{32'hc59cf671};
test_input[4376:4383] = '{32'hc18b3b6c, 32'h41705723, 32'hc00c6251, 32'h428b8347, 32'hc1dd66c4, 32'hc21b1280, 32'h417948b9, 32'h407e63ea};
test_weights[4376:4383] = '{32'hc196e085, 32'hc14fe475, 32'hc2b06ac1, 32'h420ee7bf, 32'h42c4a9a3, 32'hc230b840, 32'h408ce6d6, 32'h42858917};
test_bias[547:547] = '{32'h42a5717b};
test_output[547:547] = '{32'h450b2d4f};
test_input[4384:4391] = '{32'hc1c54479, 32'hc2c13a91, 32'h42510963, 32'h421a7cd3, 32'hc26cc9ab, 32'h42a14808, 32'h429e944c, 32'hc2bdc6ed};
test_weights[4384:4391] = '{32'h41c9dcc9, 32'h42a53cb8, 32'h40ed9e77, 32'h42acd75f, 32'hc1df5ebc, 32'hc2c51a22, 32'h41c4116f, 32'h4109d060};
test_bias[548:548] = '{32'h422ae59a};
test_output[548:548] = '{32'hc61c50fc};
test_input[4392:4399] = '{32'hc2810e2d, 32'h4282404a, 32'hc27279e6, 32'h42ad307c, 32'hc24ff659, 32'h42b5703b, 32'hc2084880, 32'h42a6f5eb};
test_weights[4392:4399] = '{32'h42be7263, 32'hc22e2113, 32'hc282dc15, 32'h41f1fe81, 32'hc2c796de, 32'h41d78664, 32'hc18f1fa4, 32'h423fb60a};
test_bias[549:549] = '{32'h41789616};
test_output[549:549] = '{32'h461a2281};
test_input[4400:4407] = '{32'hc0aad4ce, 32'hc2be65e2, 32'h427c41be, 32'hc2bd06be, 32'h420234dc, 32'hc29d2edf, 32'h429f8eb1, 32'h4225026f};
test_weights[4400:4407] = '{32'hc21094cc, 32'h413fc4c4, 32'hc297da53, 32'h40d2c617, 32'h42413717, 32'hc2411e28, 32'hc23d8650, 32'h41b52e3d};
test_bias[550:550] = '{32'hc12f7965};
test_output[550:550] = '{32'hc5708cd3};
test_input[4408:4415] = '{32'hc25b5455, 32'hc2523d17, 32'hc2a1bb04, 32'hc1d456d7, 32'h42bb63b0, 32'hc1ba28d5, 32'h429dc3b9, 32'h42798f1d};
test_weights[4408:4415] = '{32'h42bb6a5c, 32'hc2966d14, 32'hc2b6c89a, 32'h423e18f2, 32'h41c4afd3, 32'hc2b11175, 32'hc2292c6f, 32'hc244e7e0};
test_bias[551:551] = '{32'hc28f1822};
test_output[551:551] = '{32'h4530cbe1};
test_input[4416:4423] = '{32'h41ede839, 32'h3f4d12a6, 32'h421775cf, 32'hc126190a, 32'h42196a5b, 32'h42b605a6, 32'hc245098d, 32'hc2b635b1};
test_weights[4416:4423] = '{32'hc2c3f626, 32'hbf712ca9, 32'h42671d38, 32'hc2413982, 32'hc2328aad, 32'h4260db7a, 32'h3fe0d1fe, 32'hc2a28b28};
test_bias[552:552] = '{32'hc11b96ea};
test_output[552:552] = '{32'h4623dba3};
test_input[4424:4431] = '{32'hc2af78cd, 32'h42843288, 32'hc29ac5d2, 32'h41d01cf6, 32'h40d8206d, 32'hc268fe2d, 32'h411039cf, 32'hc1efaccb};
test_weights[4424:4431] = '{32'hc298a8d9, 32'hc216b3e2, 32'hc21b337c, 32'hc1961328, 32'hc21a6afa, 32'hc2769e96, 32'hc2c2b63b, 32'h42ac48e5};
test_bias[553:553] = '{32'h4041ab8b};
test_output[553:553] = '{32'h45ce231a};
test_input[4432:4439] = '{32'h42a8c336, 32'h4190d6e4, 32'hc2be7534, 32'h41bf32cc, 32'hc26149c4, 32'h41820c32, 32'h42086fe7, 32'hc1f3f43e};
test_weights[4432:4439] = '{32'h418805b3, 32'h426fbffc, 32'hc1a3571b, 32'h42051d58, 32'hc25f1776, 32'h42747593, 32'h429534a7, 32'h4165839b};
test_bias[554:554] = '{32'hc2863878};
test_output[554:554] = '{32'h4632a9a1};
test_input[4440:4447] = '{32'h427c7167, 32'h4295f8ff, 32'hc2998dda, 32'h424d8383, 32'h41a19e91, 32'hc0bab470, 32'hc2675038, 32'hc2b74b96};
test_weights[4440:4447] = '{32'h3d16d921, 32'h4288e4bf, 32'h42b0f194, 32'h4220f8b0, 32'h4205bcde, 32'h42a7e5ab, 32'h42a4e434, 32'h41d2ab5e};
test_bias[555:555] = '{32'h423c291b};
test_output[555:555] = '{32'hc5cc5422};
test_input[4448:4455] = '{32'h428aa1a3, 32'hc2a447dc, 32'hc1fdaa26, 32'hc29b0fe2, 32'hc28bd2b4, 32'h41e86c25, 32'h4247d77e, 32'hc22d7f37};
test_weights[4448:4455] = '{32'h3f3a3d64, 32'hc20da066, 32'hc1554886, 32'hc2a4809c, 32'h4249c865, 32'hc291110d, 32'hc2b670aa, 32'hc1554c33};
test_bias[556:556] = '{32'hc1b80b88};
test_output[556:556] = '{32'h42f475de};
test_input[4456:4463] = '{32'hc247486f, 32'h4118702c, 32'h42afab03, 32'hc0840284, 32'h42063b0c, 32'hc2c56218, 32'h3ec009b7, 32'hc1bcdc27};
test_weights[4456:4463] = '{32'hc23edb45, 32'hc202cd5a, 32'h42b7349f, 32'h42bb6012, 32'h420f1fce, 32'hc2c2a288, 32'h41c2efde, 32'hc11f050e};
test_bias[557:557] = '{32'h423ec7b5};
test_output[557:557] = '{32'h46a2ab1d};
test_input[4464:4471] = '{32'hc29a4f50, 32'hbf08bf01, 32'hc19acf82, 32'hc1c0404c, 32'hc1332402, 32'hc236066c, 32'hc101f6e3, 32'h427d00cb};
test_weights[4464:4471] = '{32'h425ad1ed, 32'h4296c42b, 32'hc188da49, 32'hc288af72, 32'h42952583, 32'h42afa1a1, 32'hc2310e82, 32'hc2433980};
test_bias[558:558] = '{32'h42966f1b};
test_output[558:558] = '{32'hc618abf8};
test_input[4472:4479] = '{32'h42a3ed8f, 32'h421d6070, 32'hc293b5c7, 32'h4210aef3, 32'hc2b2edac, 32'hc230b263, 32'hc29fc7d1, 32'hc1d02421};
test_weights[4472:4479] = '{32'hc1873626, 32'h41cf1f0e, 32'h41d22142, 32'hc1895583, 32'h428640b7, 32'h41953bde, 32'hc14b548a, 32'h3f4a425f};
test_bias[559:559] = '{32'hc2b53d72};
test_output[559:559] = '{32'hc60a5382};
test_input[4480:4487] = '{32'h41d8bece, 32'hc2b74ae6, 32'h427e78a6, 32'h41dfdf9b, 32'h426e6b95, 32'h426d70c5, 32'hc2871d6f, 32'h4192bf03};
test_weights[4480:4487] = '{32'hc223d37d, 32'h42994d80, 32'hc017c7c0, 32'hc1715ada, 32'hc2a4acec, 32'h4231e9ee, 32'hc2ba316d, 32'hc20e4538};
test_bias[560:560] = '{32'hc2775609};
test_output[560:560] = '{32'hc5a8bed2};
test_input[4488:4495] = '{32'hc1d1b5c5, 32'hc1f33345, 32'h4236ed9c, 32'h42b517de, 32'hc1d294fd, 32'h4259a5b3, 32'h423c777b, 32'hc2b7ac13};
test_weights[4488:4495] = '{32'h425041c1, 32'h42bada7b, 32'hc2832112, 32'hc1de0c5d, 32'hc10b862c, 32'hc20c9799, 32'hc2a62182, 32'hc1eb3612};
test_bias[561:561] = '{32'hbf55908a};
test_output[561:561] = '{32'hc645180d};
test_input[4496:4503] = '{32'hc1584d28, 32'h419d6ce0, 32'hc255212f, 32'hc1c04627, 32'h424419ab, 32'h415454d8, 32'hc2b1b005, 32'h41a33c84};
test_weights[4496:4503] = '{32'h419fb05e, 32'hc2792caa, 32'hc2921d27, 32'hc2987fbf, 32'h41f5759a, 32'hc28a8b02, 32'h41f2d66e, 32'h401a5611};
test_bias[562:562] = '{32'hc22b9f1b};
test_output[562:562] = '{32'h4504bf93};
test_input[4504:4511] = '{32'hc2a9a1a2, 32'hc2836809, 32'hc28fcd50, 32'hbf5f6751, 32'hc2bdd966, 32'hc254864c, 32'h42c6f9a8, 32'h4215d52d};
test_weights[4504:4511] = '{32'hc233ba4d, 32'hc1a251cc, 32'h42b10b3a, 32'h423d47f2, 32'hc2a45922, 32'hc1b81b17, 32'h42868295, 32'h42b62a14};
test_bias[563:563] = '{32'hc1afc327};
test_output[563:563] = '{32'h468b63b1};
test_input[4512:4519] = '{32'h4298e4e4, 32'h4192a4f6, 32'h423f262b, 32'hc2175d31, 32'hc22484d1, 32'hc29cf828, 32'h4212e580, 32'hbfad45d7};
test_weights[4512:4519] = '{32'h42b1d399, 32'hc13ab1a2, 32'hc25b724a, 32'hc23b5a96, 32'h41cd5722, 32'h42aedafa, 32'hc0e2c77f, 32'h4296dec1};
test_bias[564:564] = '{32'hc29a98e3};
test_output[564:564] = '{32'hc523f1b9};
test_input[4520:4527] = '{32'hc27ad3a6, 32'h42c4ffc6, 32'h42c031e9, 32'hc29edd3c, 32'hc2c0405a, 32'hc214be73, 32'hc1d36b18, 32'hc241dad5};
test_weights[4520:4527] = '{32'h42c7cc11, 32'hc28b3a66, 32'hc2321dad, 32'hc1897529, 32'h41ffb788, 32'hc2946ee3, 32'h41bfb414, 32'hc292b2b0};
test_bias[565:565] = '{32'hc2a75899};
test_output[565:565] = '{32'hc6531a38};
test_input[4528:4535] = '{32'hc1b328a0, 32'h41ee7475, 32'hc27ad19f, 32'h426b3626, 32'h41974e13, 32'h422e7d0a, 32'h42b694c0, 32'hc1686fe4};
test_weights[4528:4535] = '{32'h42082b69, 32'h41b41ce5, 32'h42687b7f, 32'h425b78b7, 32'hc21105d1, 32'hc1029ad1, 32'hc2a88c0a, 32'hc2020a92};
test_bias[566:566] = '{32'hc200b137};
test_output[566:566] = '{32'hc609918f};
test_input[4536:4543] = '{32'hc2ab5a9f, 32'hc247e72a, 32'hc2897554, 32'h424b0d31, 32'h4202f27e, 32'hc2441bcd, 32'h41d33be2, 32'hc2b81d5b};
test_weights[4536:4543] = '{32'hc25c513e, 32'h41354950, 32'h42878a06, 32'h4262067a, 32'hc1eddd04, 32'hc2751f8f, 32'h4218595e, 32'h40987a1d};
test_bias[567:567] = '{32'h4233a15d};
test_output[567:567] = '{32'h459c73a9};
test_input[4544:4551] = '{32'h4164c61e, 32'hc26adcff, 32'hc1fdeac3, 32'h413eb712, 32'h42c5caaf, 32'h4136ad0d, 32'h42c5f873, 32'hc250b65a};
test_weights[4544:4551] = '{32'hc2a59504, 32'h4227910e, 32'hc29b58c9, 32'hc29848ab, 32'h42bfb57c, 32'hc1294d5c, 32'h4218bc34, 32'hc22ca898};
test_bias[568:568] = '{32'h40035345};
test_output[568:568] = '{32'h464febf5};
test_input[4552:4559] = '{32'h407d6016, 32'hc1957209, 32'h4213b20f, 32'hc2c4e35c, 32'h4218b48d, 32'h42c732e9, 32'h41d5f449, 32'hc14e6e5c};
test_weights[4552:4559] = '{32'h427ba518, 32'hc25a7c79, 32'h3f9f6180, 32'hc2042b5d, 32'h3f7fe202, 32'hc28c454e, 32'h42c4252e, 32'h420c4ced};
test_bias[569:569] = '{32'hc21584ab};
test_output[569:569] = '{32'hc376162f};
test_input[4560:4567] = '{32'hc2447019, 32'h4177c037, 32'hc1677ce8, 32'hc25422e6, 32'hc257817f, 32'hc1962f22, 32'hc1a4d6f7, 32'h42932033};
test_weights[4560:4567] = '{32'hc2c3fdf7, 32'h42868218, 32'hc138376d, 32'hc2a6ffb0, 32'h426f5f7b, 32'h424d5f0c, 32'h42b7fed9, 32'h40967a0d};
test_bias[570:570] = '{32'h42c14042};
test_output[570:570] = '{32'h45963e01};
test_input[4568:4575] = '{32'hc2bbcc94, 32'h422516a9, 32'hc0d05542, 32'h414a3bde, 32'h425dade4, 32'h426d400d, 32'hc109eb61, 32'h42c5df15};
test_weights[4568:4575] = '{32'hc0463f28, 32'h429adea5, 32'hc25314fa, 32'hc18801a9, 32'h41534088, 32'hc2796fcb, 32'hc22b4b69, 32'hc1dcf59d};
test_bias[571:571] = '{32'hc29f3906};
test_output[571:571] = '{32'hc4e052eb};
test_input[4576:4583] = '{32'hbf254686, 32'hc2a778b0, 32'h426b9bb2, 32'hc1cd7404, 32'hc238fa71, 32'h42aa7605, 32'hc280c4de, 32'h4258a59b};
test_weights[4576:4583] = '{32'hc27e3445, 32'hc24a3116, 32'hc19f2764, 32'h4227082f, 32'hc2236c7d, 32'hc2c33adb, 32'hc2206672, 32'h41e519c8};
test_bias[572:572] = '{32'h42b8741c};
test_output[572:572] = '{32'hc32fd31e};
test_input[4584:4591] = '{32'h42a2ee4f, 32'h428b8cac, 32'hc2800565, 32'hc22a2731, 32'hc19f384d, 32'h428921dc, 32'h412d84ec, 32'h4294ae82};
test_weights[4584:4591] = '{32'hc20d7c2b, 32'h41ae8017, 32'h41f2a48d, 32'hc23ddbd6, 32'h428c3f31, 32'h42a753b0, 32'h42bff6b1, 32'hc25a63ab};
test_bias[573:573] = '{32'h4222eaca};
test_output[573:573] = '{32'h42a36fad};
test_input[4592:4599] = '{32'hc217b0fe, 32'h4215f6ef, 32'hc217d52c, 32'hc218cd3e, 32'h42932333, 32'hc2c60f3b, 32'h41fa7144, 32'hc28eb071};
test_weights[4592:4599] = '{32'hc1023c4f, 32'hc210e499, 32'hc2c5ee22, 32'h42c7d2ed, 32'h3f0c5451, 32'hc1d3e580, 32'hc24f8ffa, 32'h4283e8bf};
test_bias[574:574] = '{32'hc293dc6d};
test_output[574:574] = '{32'hc5979087};
test_input[4600:4607] = '{32'h3fe813b9, 32'hc290beb1, 32'h42bef575, 32'h42c2bf9d, 32'h42b9d2f1, 32'hc1d03674, 32'h428df87e, 32'hc199a076};
test_weights[4600:4607] = '{32'hc2b79cd9, 32'hc290d222, 32'h42313e32, 32'hc245c81a, 32'h428a2b12, 32'hc28ac35d, 32'hc22073d4, 32'h4242d8a3};
test_bias[575:575] = '{32'h42b0baa8};
test_output[575:575] = '{32'h460cf07f};
test_input[4608:4615] = '{32'hc29083b1, 32'hc0e2a18e, 32'hc1d774a6, 32'h4239b43d, 32'hc2c0e6a5, 32'h41fea4e7, 32'h420a75ef, 32'hc2887bc5};
test_weights[4608:4615] = '{32'hc224ad59, 32'hc06b4524, 32'h429971c1, 32'hc255b25c, 32'h4156f807, 32'hc1a9e574, 32'h41fd8824, 32'h41d9d340};
test_bias[576:576] = '{32'hc2afbbb5};
test_output[576:576] = '{32'hc588745f};
test_input[4616:4623] = '{32'h425bb2c0, 32'hc2000d0d, 32'h42c3c2b3, 32'h422e4712, 32'h412b5fa9, 32'h421542a4, 32'h42456c60, 32'hc0053457};
test_weights[4616:4623] = '{32'hc289799c, 32'hc17b465b, 32'h42890ffd, 32'h422004a8, 32'hc24e84c3, 32'h4269a690, 32'hbf22d8e4, 32'h420836e6};
test_bias[577:577] = '{32'h4214ea0a};
test_output[577:577] = '{32'h45d29ea9};
test_input[4624:4631] = '{32'hc19befbf, 32'hc2b8cfca, 32'h411cf717, 32'h42690ce0, 32'hc2604939, 32'hc153f674, 32'h419a86d9, 32'hc1fdcdcd};
test_weights[4624:4631] = '{32'h429af0f6, 32'h421a5d7f, 32'h42807ce8, 32'hc28b06c5, 32'hc25348fb, 32'hc26e3028, 32'hc10acf44, 32'hc24ee260};
test_bias[578:578] = '{32'hc28bc1de};
test_output[578:578] = '{32'hc550dd73};
test_input[4632:4639] = '{32'h42a6765d, 32'h4124a9d1, 32'hc2b54c12, 32'hc246b9c4, 32'h428b855f, 32'h42be6862, 32'hc22f4d28, 32'hc2b6b577};
test_weights[4632:4639] = '{32'hc1f36139, 32'h42bde458, 32'h425e0c13, 32'hc27bd9ee, 32'hc2c2c961, 32'h428fb56c, 32'h4261db5b, 32'h42c1e4b7};
test_bias[579:579] = '{32'hc28f8969};
test_output[579:579] = '{32'hc6677cbe};
test_input[4640:4647] = '{32'hc2571423, 32'h3fc76326, 32'h429755bb, 32'hc2278d96, 32'hc28823e0, 32'hc2536ed3, 32'h425b7029, 32'h42afe752};
test_weights[4640:4647] = '{32'h42ab3f6c, 32'h429bc2cd, 32'h42b5812c, 32'hc2973350, 32'h4156ee8b, 32'hc2649212, 32'hc13d1f73, 32'hc170dffa};
test_bias[580:580] = '{32'h42b92ea6};
test_output[580:580] = '{32'h45b489bd};
test_input[4648:4655] = '{32'h4261a667, 32'h42ab42da, 32'h421e163a, 32'h41810d8a, 32'h4197cd34, 32'h42b176e1, 32'h410e36e5, 32'hc245253c};
test_weights[4648:4655] = '{32'h4295dee2, 32'h42ba0cfb, 32'hc23a9c54, 32'h426b773f, 32'h420af0a5, 32'hc2c50f2e, 32'h42838b9f, 32'hc2c1e767};
test_bias[581:581] = '{32'hc18cfc29};
test_output[581:581] = '{32'h4605c2b1};
test_input[4656:4663] = '{32'h4128959e, 32'hbf93ef8b, 32'hc1dca430, 32'hc267a3fb, 32'h422581f8, 32'h425b057d, 32'h410a5b7b, 32'hc2090eb0};
test_weights[4656:4663] = '{32'h42a0b925, 32'h42b3184d, 32'h422ee124, 32'h414e9c52, 32'h42b6e9ac, 32'hc2c498eb, 32'hc23179a2, 32'h42a7cbad};
test_bias[582:582] = '{32'h42572ebf};
test_output[582:582] = '{32'hc5bbe920};
test_input[4664:4671] = '{32'h423be02d, 32'h413b3bd5, 32'hc284d7bd, 32'h41327581, 32'hc1f4beac, 32'hc27ae3eb, 32'hc1100aa9, 32'h41b58c8b};
test_weights[4664:4671] = '{32'hc2978b69, 32'hc209d305, 32'hc2c0519a, 32'hc23af69d, 32'hc21d1325, 32'h4269941b, 32'hc1f3b9ba, 32'h4085bedc};
test_bias[583:583] = '{32'h41a494fa};
test_output[583:583] = '{32'hc32810b4};
test_input[4672:4679] = '{32'hc1f78629, 32'hc1cc00e6, 32'h429b2417, 32'h4176419e, 32'h4185cc44, 32'h41a17085, 32'hc2a0ee26, 32'h41c2cd7b};
test_weights[4672:4679] = '{32'hc22a5e8f, 32'hc2043aa3, 32'hc297dba8, 32'hc290dd10, 32'h428f6269, 32'h428142b5, 32'hc110ee7b, 32'h42b7a2a5};
test_bias[584:584] = '{32'h42ba12c9};
test_output[584:584] = '{32'h443347c6};
test_input[4680:4687] = '{32'h421e1c51, 32'hbff36228, 32'h41c5abb9, 32'hc1a88a3f, 32'h421eef7b, 32'h42485ba4, 32'h42ae1914, 32'hc1963972};
test_weights[4680:4687] = '{32'hc29db861, 32'h42b17de8, 32'h42c7e135, 32'hc1684955, 32'hc2811c06, 32'hc0e97276, 32'h4219407c, 32'h429e72be};
test_bias[585:585] = '{32'hc2951502};
test_output[585:585] = '{32'hc4d085b1};
test_input[4688:4695] = '{32'hc26ec10c, 32'hc211db69, 32'hc2c1c60b, 32'hc2b4a66c, 32'hc246df30, 32'h42c3c09d, 32'h41387c80, 32'h42b87821};
test_weights[4688:4695] = '{32'hc2600725, 32'hc2bd0f38, 32'h42805b36, 32'hc25f672e, 32'hc2a617e3, 32'hc2c749d2, 32'hc22cdd80, 32'h4286d33b};
test_bias[586:586] = '{32'h415c00f8};
test_output[586:586] = '{32'h45b2efd0};
test_input[4696:4703] = '{32'hc221817f, 32'h421e5acd, 32'h41a62953, 32'h41fc076c, 32'hc067c94f, 32'hc2665fab, 32'hc26b4a69, 32'h42c0236d};
test_weights[4696:4703] = '{32'h41a827f0, 32'h4099ef52, 32'h3eff7b34, 32'h42a4cb63, 32'hc1e6ea1d, 32'h4267159e, 32'hc2b4454a, 32'hc2aa8275};
test_bias[587:587] = '{32'h42bcdbb7};
test_output[587:587] = '{32'hc57e4b4f};
test_input[4704:4711] = '{32'h4271c411, 32'h42382911, 32'h4095c97c, 32'h419a7c74, 32'h422758b6, 32'hc1397908, 32'hc0523a2a, 32'hc277b010};
test_weights[4704:4711] = '{32'hc1d71909, 32'h423b3f86, 32'h42023ddd, 32'hc2b806bd, 32'hc092f1fb, 32'hc208730d, 32'hc2903295, 32'hc288941f};
test_bias[588:588] = '{32'h4177c5e2};
test_output[588:588] = '{32'h45605ee5};
test_input[4712:4719] = '{32'hc258ba91, 32'h4179992a, 32'hc2a92d61, 32'h426a9dee, 32'h41337656, 32'hc2770900, 32'hc0ecccc1, 32'hc2bc438a};
test_weights[4712:4719] = '{32'h4232f773, 32'hc229c6c9, 32'hc1db5fb0, 32'hc2243276, 32'h428da72e, 32'h4210247b, 32'h413b4ef5, 32'hc28bef90};
test_bias[589:589] = '{32'hc293955c};
test_output[589:589] = '{32'h44e38703};
test_input[4720:4727] = '{32'hc1b78057, 32'hc2984d02, 32'h42687910, 32'h428bc8c2, 32'hc2c13b64, 32'hc268c5fd, 32'h41a54631, 32'h41d15a0e};
test_weights[4720:4727] = '{32'h4295d169, 32'hc0534be1, 32'h41a4921f, 32'h428cfdf6, 32'hc198a205, 32'hc2c1588f, 32'h4164f627, 32'hc2a8812c};
test_bias[590:590] = '{32'h421242c2};
test_output[590:590] = '{32'h46203157};
test_input[4728:4735] = '{32'h422a6ac1, 32'hc239bdbb, 32'h42b1de5b, 32'hc2a1d139, 32'h40b3d7b8, 32'hc216d758, 32'hc2b1ecd3, 32'hc2969acf};
test_weights[4728:4735] = '{32'hc1eb0d81, 32'h42c01f7c, 32'h426a029d, 32'h414c2c3e, 32'hc2169331, 32'h4257a23e, 32'h42ab78b2, 32'hc199999c};
test_bias[591:591] = '{32'h41f4045e};
test_output[591:591] = '{32'hc61b45b3};
test_input[4736:4743] = '{32'hc294a776, 32'h427366f6, 32'hc1df8b4c, 32'hc2acf5b4, 32'h4264141f, 32'hbf3d3ede, 32'h4242c445, 32'hc2ae9387};
test_weights[4736:4743] = '{32'h4246e00e, 32'hc2a92b76, 32'h413957bf, 32'hc2c3403d, 32'hc19a65cb, 32'hc2069da8, 32'h419abf00, 32'h40b67cfc};
test_bias[592:592] = '{32'h429e333d};
test_output[592:592] = '{32'hc49f7e6e};
test_input[4744:4751] = '{32'h429f411c, 32'hc0a45bca, 32'h4286aade, 32'hc0f70785, 32'h41d796dc, 32'hc23aa67d, 32'hc2957dcf, 32'hc1a19a1c};
test_weights[4744:4751] = '{32'h422c7a94, 32'h41ae367b, 32'h41aa5e48, 32'h41a23500, 32'hc11dec0e, 32'h41a95fae, 32'h420f0153, 32'h42205aea};
test_bias[593:593] = '{32'h420aab7f};
test_output[593:593] = '{32'hc2cc7946};
test_input[4752:4759] = '{32'hc112985e, 32'h42011fa6, 32'hc23997e8, 32'h426f36a9, 32'hc21a8537, 32'h4287ed79, 32'h42023db1, 32'h429d7423};
test_weights[4752:4759] = '{32'h4246dc11, 32'h41aa9e30, 32'hc25822e1, 32'h42b43586, 32'h419db977, 32'hc2bbc2ee, 32'h41c618df, 32'h42b767ae};
test_bias[594:594] = '{32'h42c2e25b};
test_output[594:594] = '{32'h460e56a1};
test_input[4760:4767] = '{32'hc28648b9, 32'h42bf277d, 32'hc2a65b31, 32'hc2ab34b4, 32'h41c1fa0d, 32'h421487fd, 32'hc28c35c8, 32'hc2873abf};
test_weights[4760:4767] = '{32'hc23ce9bf, 32'h4056f86c, 32'hc14a2b5e, 32'hc1a79955, 32'hc26eb0ec, 32'hc2c133b2, 32'h42b6815f, 32'h4283942f};
test_bias[595:595] = '{32'hc222ccb6};
test_output[595:595] = '{32'hc615bf68};
test_input[4768:4775] = '{32'h428fe9e9, 32'hc034b996, 32'hc1831254, 32'h4239d244, 32'hc2bd0fc2, 32'hc24f9829, 32'h4277f051, 32'h41c247c1};
test_weights[4768:4775] = '{32'hc2a808d6, 32'h428e3d95, 32'hc1e99887, 32'hc20d98bc, 32'h41937ec5, 32'hc24053ea, 32'h41c99ac9, 32'h4120ce43};
test_bias[596:596] = '{32'hc296999a};
test_output[596:596] = '{32'hc59a0960};
test_input[4776:4783] = '{32'hc28f6f7a, 32'h4240036b, 32'hc2892ee8, 32'h426a502c, 32'hc209e31a, 32'hc174d3b9, 32'hc29c2d31, 32'h41962a69};
test_weights[4776:4783] = '{32'h428db3de, 32'hc1d77796, 32'hc27623d7, 32'h42a62a05, 32'hc28be085, 32'hc13dd8b2, 32'h42b3da23, 32'h41ab11e4};
test_bias[597:597] = '{32'h404d1923};
test_output[597:597] = '{32'hc4a3f69d};
test_input[4784:4791] = '{32'h420f196c, 32'hc226c081, 32'h426e5ecb, 32'hc2644eb6, 32'hc20b94b9, 32'h42410e4c, 32'h42a4f8d2, 32'h421888f1};
test_weights[4784:4791] = '{32'hc2ae45d1, 32'hc23db2b4, 32'hc2a49b8f, 32'h428808be, 32'h426eb9ea, 32'h429ed1c3, 32'h4267284a, 32'hc1b7381c};
test_bias[598:598] = '{32'h4214edb3};
test_output[598:598] = '{32'hc584b386};
test_input[4792:4799] = '{32'hc1a133aa, 32'h409a7290, 32'h42ba8991, 32'hc262919d, 32'h423e514d, 32'h41a754fb, 32'hc10dfd65, 32'hc2a59141};
test_weights[4792:4799] = '{32'h42b16c27, 32'h41ab5c69, 32'hc298158f, 32'h426e78e0, 32'h401c5a94, 32'hc1cd6ff6, 32'hc20bb6bb, 32'h402a92f8};
test_bias[599:599] = '{32'hc2436b97};
test_output[599:599] = '{32'hc643d74f};
test_input[4800:4807] = '{32'hc2866cd9, 32'h42c63c5a, 32'h42816da4, 32'hc2452d5b, 32'h4196342e, 32'h42be23f8, 32'hc0d795a2, 32'h41c10a29};
test_weights[4800:4807] = '{32'h420646b0, 32'h41cafeaa, 32'h4217238b, 32'hc21fb693, 32'h421b0770, 32'hc23b930c, 32'hc1e0ed39, 32'h42b6d3e1};
test_bias[600:600] = '{32'hc23e88f3};
test_output[600:600] = '{32'h454d953c};
test_input[4808:4815] = '{32'h40343de4, 32'hc2b9f5f8, 32'h4282d5a0, 32'h425ed543, 32'hc183738e, 32'h4295ba5d, 32'hc263656d, 32'hbb0763bb};
test_weights[4808:4815] = '{32'hc213ff43, 32'h42951d60, 32'hc259acd0, 32'h4261cb09, 32'h4231341d, 32'hc2a94ec3, 32'h42c0e809, 32'hc22198be};
test_bias[601:601] = '{32'hc2b783d6};
test_output[601:601] = '{32'hc69cf886};
test_input[4816:4823] = '{32'hc2c68fbe, 32'h42706f6e, 32'hc0e8f0a5, 32'hc27a1f2c, 32'h42a105b4, 32'h4210dbc2, 32'hc2812ca3, 32'h4211f48a};
test_weights[4816:4823] = '{32'hc03431f6, 32'hc28f0bcd, 32'hc09ce6fc, 32'h421d2bb7, 32'h42aea81e, 32'h42af50ee, 32'h4207b1cf, 32'h42b7e706};
test_bias[602:602] = '{32'hc2107d4f};
test_output[602:602] = '{32'h4598e415};
test_input[4824:4831] = '{32'hc14c758b, 32'hc18e5616, 32'h42895f7d, 32'hc2347768, 32'hc2a8033e, 32'h41908b65, 32'hc1d33713, 32'hc11597b5};
test_weights[4824:4831] = '{32'h42865373, 32'h42992ecd, 32'hc2909feb, 32'h4256128c, 32'h42b294d2, 32'hc191b344, 32'h4141ffe4, 32'h4286d86f};
test_bias[603:603] = '{32'h415ce5fb};
test_output[603:603] = '{32'hc68f8249};
test_input[4832:4839] = '{32'h4285318b, 32'h411c9923, 32'hc2af1c19, 32'hc1a9931b, 32'h41e8fd1a, 32'h42415cf8, 32'hc2c1b522, 32'hc2a440f3};
test_weights[4832:4839] = '{32'h41a1a9b2, 32'h426f184a, 32'h42a8b2c9, 32'hc224a05d, 32'h42a3f75a, 32'h41a86fb7, 32'h42a08298, 32'hc216577d};
test_bias[604:604] = '{32'hc2a1a803};
test_output[604:604] = '{32'hc5b9bce5};
test_input[4840:4847] = '{32'hc264d6c5, 32'h42134c13, 32'h41c9b865, 32'h42060b44, 32'hc2841e0b, 32'h422f5643, 32'h423d5b29, 32'hc149e952};
test_weights[4840:4847] = '{32'h41c97be3, 32'hc2adcbf0, 32'hc1d629d6, 32'hc21d6287, 32'hbf5a85c4, 32'h42ba2080, 32'h3f9cca8d, 32'hc2633af9};
test_bias[605:605] = '{32'hc2887af8};
test_output[605:605] = '{32'hc4dfffad};
test_input[4848:4855] = '{32'h3ff48dfc, 32'h423ff13c, 32'h41cd8087, 32'h42a71e26, 32'hc18fc497, 32'h42a41c75, 32'hc29ed96a, 32'hc0d02ea6};
test_weights[4848:4855] = '{32'h41b6dc06, 32'h428c6bb5, 32'hc250e361, 32'hc17bc2ba, 32'h41aa8d72, 32'h422843c5, 32'hc286cd6f, 32'hc1e63763};
test_bias[606:606] = '{32'hc181dd7a};
test_output[606:606] = '{32'h461215b5};
test_input[4856:4863] = '{32'h42beacbd, 32'hc013fd99, 32'h425a1263, 32'h418335b2, 32'hc21b83bb, 32'h42c04f35, 32'hc2b9f659, 32'h420bb8eb};
test_weights[4856:4863] = '{32'h427090e7, 32'h428b769a, 32'hc08cf904, 32'h4265c85e, 32'hc23649df, 32'h41896bd3, 32'h42a47d3f, 32'h4288b323};
test_bias[607:607] = '{32'hc253b9bf};
test_output[607:607] = '{32'h45890ae2};
test_input[4864:4871] = '{32'hc171227c, 32'h4230bb73, 32'h425e63e4, 32'hc1f914e5, 32'hc21cd873, 32'h406d07ca, 32'hc299d17a, 32'h42abe6d6};
test_weights[4864:4871] = '{32'hc1d33e01, 32'hc2a256f3, 32'hc257fe26, 32'hc25742af, 32'h42c69cb8, 32'h419914d2, 32'h42819370, 32'h42715f90};
test_bias[608:608] = '{32'hc0f0b78d};
test_output[608:608] = '{32'hc5fe6e79};
test_input[4872:4879] = '{32'hc2ae0fed, 32'h41bca85b, 32'h418841f2, 32'hc273894a, 32'h4194adbe, 32'hc1ba92b7, 32'hc1f000d2, 32'hc171f6f9};
test_weights[4872:4879] = '{32'hc29c0a64, 32'h421c1f48, 32'hc05ed492, 32'hc20949ac, 32'hc07c5189, 32'hc1de5370, 32'hc1e9635c, 32'hc27e01b8};
test_bias[609:609] = '{32'h429c588e};
test_output[609:609] = '{32'h463f162e};
test_input[4880:4887] = '{32'h421e7642, 32'hc2ab89a2, 32'hc1abff76, 32'hc2846c86, 32'hc1524f82, 32'hc1ff2849, 32'hc23ea7bb, 32'h42b078ab};
test_weights[4880:4887] = '{32'h42b534da, 32'h42506d33, 32'hc26897ad, 32'hc292505d, 32'h41cd9a08, 32'hc2984fcb, 32'hc2c2d68b, 32'h413f0b4d};
test_bias[610:610] = '{32'hc22b0994};
test_output[610:610] = '{32'h464a7e0c};
test_input[4888:4895] = '{32'h416d0fdc, 32'hc1e747d4, 32'h41c077d8, 32'hc21e113f, 32'hc2c125b6, 32'hc2ae5621, 32'hc2c6a5f0, 32'h4287b665};
test_weights[4888:4895] = '{32'hc2a4fcd3, 32'hc296bd84, 32'hc223018e, 32'h41beea63, 32'h41e0d6f7, 32'h429d242b, 32'hc26bc047, 32'h4286e72e};
test_bias[611:611] = '{32'h42b2bd3f};
test_output[611:611] = '{32'hc118404e};
test_input[4896:4903] = '{32'hc2926ba4, 32'h4293a21c, 32'hc2a55950, 32'hc0c8fc82, 32'h41858545, 32'h41d5e921, 32'hc2527e20, 32'h4213c832};
test_weights[4896:4903] = '{32'h4210d5c2, 32'hc0af6767, 32'hc2b57b29, 32'h429b494d, 32'hc20d91cf, 32'hc16460eb, 32'hc223893c, 32'hc2b59324};
test_bias[612:612] = '{32'h416b1e6c};
test_output[612:612] = '{32'h44e0cc61};
test_input[4904:4911] = '{32'hc2c2e95e, 32'h4215be41, 32'h41f5bf4f, 32'h423990f8, 32'h42918996, 32'hc0f327c8, 32'hc0bf9bb4, 32'hc2637edd};
test_weights[4904:4911] = '{32'hc25d2f34, 32'h42bb676d, 32'hc28ec8fb, 32'hc2b06d83, 32'hc1e9dbf8, 32'hc291d00e, 32'hc04cfebf, 32'hc2897584};
test_bias[613:613] = '{32'h425b3a42};
test_output[613:613] = '{32'h459ce7c4};
test_input[4912:4919] = '{32'h4062b6bd, 32'h429da8a2, 32'hc28a9c1a, 32'h41b137de, 32'h4269109d, 32'hc23f7dc5, 32'hc244661f, 32'h40f8d170};
test_weights[4912:4919] = '{32'hc28e2c3b, 32'hc2c3cc53, 32'hc1f222cb, 32'h429ca047, 32'hc273d186, 32'hc2b7d0ac, 32'h4164c45b, 32'h429932f9};
test_bias[614:614] = '{32'h421431e5};
test_output[614:614] = '{32'hc551dc48};
test_input[4920:4927] = '{32'hc2602046, 32'h4165c07e, 32'hc25dbb21, 32'hc1a5a8d1, 32'h4203bc0b, 32'hc240e05f, 32'hc2117170, 32'h41039f0c};
test_weights[4920:4927] = '{32'h41acfe1b, 32'hc2813b6a, 32'h4286293a, 32'h4275c604, 32'hc2979cde, 32'h4121c6f4, 32'hc278102d, 32'h42bc835b};
test_bias[615:615] = '{32'hbfad209c};
test_output[615:615] = '{32'hc5dd6b69};
test_input[4928:4935] = '{32'hc22be875, 32'hc23cd2e8, 32'h40b85c71, 32'hc23f9ac1, 32'h41106992, 32'h42099ada, 32'hc209f265, 32'hc084bddf};
test_weights[4928:4935] = '{32'h428577d5, 32'hc04d0afe, 32'h41c2343c, 32'h41f77b7c, 32'hc2973a2e, 32'hc220ed13, 32'h41ce2faf, 32'h426c7729};
test_bias[616:616] = '{32'h41c9c860};
test_output[616:616] = '{32'hc5e210bc};
test_input[4936:4943] = '{32'h42c6f21d, 32'hc24a3451, 32'hc233136e, 32'h42a5c6e9, 32'h4206d8fe, 32'h40cd955a, 32'hc1c0671c, 32'hc2b8a12d};
test_weights[4936:4943] = '{32'h3fb49488, 32'hc130515c, 32'h421e69d5, 32'hc2763138, 32'h41495f87, 32'h42b3405c, 32'h4295e759, 32'h4293e643};
test_bias[617:617] = '{32'h422e13dd};
test_output[617:617] = '{32'hc6570b8e};
test_input[4944:4951] = '{32'hc2b99f31, 32'hc2764dec, 32'hc28d8f8d, 32'h414cc6b3, 32'h41e25e24, 32'h4217c9f2, 32'h41efb5e2, 32'hc1da8efa};
test_weights[4944:4951] = '{32'hc25567ae, 32'hc233660b, 32'hc2060d92, 32'h42ab37d7, 32'h41dc3e02, 32'h4280c1d2, 32'h41bb38d4, 32'hc184a12c};
test_bias[618:618] = '{32'h42976c0c};
test_output[618:618] = '{32'h46744366};
test_input[4952:4959] = '{32'h419d2613, 32'hc16d7f46, 32'hc29a254c, 32'h4102e2f9, 32'hc2bc5d6f, 32'h42b68fd7, 32'hc134c947, 32'hc2838fa9};
test_weights[4952:4959] = '{32'h41e049c4, 32'hc01b749a, 32'hc197564e, 32'h428891e2, 32'h416dbddb, 32'h42258b1d, 32'hc2271c07, 32'hc0c31327};
test_bias[619:619] = '{32'h42a8837d};
test_output[619:619] = '{32'h45b997e2};
test_input[4960:4967] = '{32'h41cb120a, 32'h425dbc2d, 32'h41bbc074, 32'h41d3c976, 32'h42bfda07, 32'hc2aa09e7, 32'hc245d6db, 32'hc18c7fbb};
test_weights[4960:4967] = '{32'h4297014b, 32'h401b1e8d, 32'h41ef5250, 32'h41c9eecb, 32'h42614664, 32'h42aa2c9c, 32'hc18a8488, 32'hc0ee0860};
test_bias[620:620] = '{32'hc2672910};
test_output[620:620] = '{32'h451d6cf1};
test_input[4968:4975] = '{32'h3e34cbb9, 32'hc1ba7e73, 32'h3fe8aa50, 32'h41389909, 32'hc2b8e16b, 32'h42839bad, 32'hc2b106b8, 32'hc2a1a64d};
test_weights[4968:4975] = '{32'h402c2d15, 32'h41481060, 32'hc2350fb6, 32'h42b1c011, 32'h4217a8ef, 32'h429fe496, 32'h3f3ed533, 32'hc2ab2e64};
test_bias[621:621] = '{32'h422f306f};
test_output[621:621] = '{32'h46115eb9};
test_input[4976:4983] = '{32'h4271fac8, 32'hc0955695, 32'hc1209495, 32'hc2c399c8, 32'h4297e02a, 32'hc2537ce6, 32'h428b8e5f, 32'hc239da5b};
test_weights[4976:4983] = '{32'h42a549ba, 32'hc2b543cd, 32'h423d2106, 32'h412a535d, 32'hc2c1193a, 32'h41b70987, 32'hc298dc3b, 32'hc29db9d1};
test_bias[622:622] = '{32'hc2332c9c};
test_output[622:622] = '{32'hc5c66264};
test_input[4984:4991] = '{32'hc2a89fbe, 32'h42849a93, 32'hc268c187, 32'h3f895182, 32'hc2229541, 32'hc26d2d44, 32'h42867ff6, 32'hc20b3da0};
test_weights[4984:4991] = '{32'h3fdd8f8b, 32'h42043e6b, 32'hc2a0117d, 32'hc21459f7, 32'hc2a56a50, 32'h426c54c7, 32'hc284e799, 32'h41664729};
test_bias[623:623] = '{32'h42211d9c};
test_output[623:623] = '{32'h44c7063d};
test_input[4992:4999] = '{32'hc2b96f14, 32'hc1b9429a, 32'hc2617c85, 32'hc129a131, 32'h41374591, 32'h425169c0, 32'h4236f797, 32'hc2217a4b};
test_weights[4992:4999] = '{32'hc1b49d46, 32'h41e89969, 32'h4235b5b0, 32'h40a087d7, 32'h41b137cc, 32'h41522eea, 32'hc2554b86, 32'h41b85a2b};
test_bias[624:624] = '{32'hc19ba556};
test_output[624:624] = '{32'hc56396d9};
test_input[5000:5007] = '{32'h41923f29, 32'hc28f7eae, 32'h42990a5b, 32'hc27be452, 32'hc28c0295, 32'h4189c794, 32'h42838fe1, 32'h42747f36};
test_weights[5000:5007] = '{32'h4260dca0, 32'hc236becb, 32'hc09bbf44, 32'hbf614e4f, 32'hc1b5a3d0, 32'h42304d76, 32'h416e29ca, 32'hc1b9d005};
test_bias[625:625] = '{32'hc19d559a};
test_output[625:625] = '{32'h45b7a705};
test_input[5008:5015] = '{32'hc1ddb302, 32'h41b0bc48, 32'h4007f504, 32'h427836b6, 32'h41bc4bfd, 32'h42a0c855, 32'hc029d875, 32'hc1775036};
test_weights[5008:5015] = '{32'h3f861698, 32'h41272006, 32'h4268c4e1, 32'hc2b880f0, 32'hc29b1727, 32'h42bc4af8, 32'h426227fb, 32'h4183aff6};
test_bias[626:626] = '{32'hc265fec8};
test_output[626:626] = '{32'hc2eba245};
test_input[5016:5023] = '{32'hc13805b3, 32'hc273e4e4, 32'h41deb76f, 32'hc26dbd40, 32'h42474fdd, 32'h41259e6f, 32'h422ae720, 32'h4253d868};
test_weights[5016:5023] = '{32'hc0b91604, 32'hc27981be, 32'hc23cb10c, 32'hc26cea2c, 32'hc2626a6b, 32'h42b3db7b, 32'hc218e0aa, 32'h41c87661};
test_bias[627:627] = '{32'h42276ef3};
test_output[627:627] = '{32'h457533bc};
test_input[5024:5031] = '{32'hc17ae95e, 32'h42b8c269, 32'hc20c7230, 32'hc29f1553, 32'hc234ae90, 32'h42bb95d7, 32'hc1d85a71, 32'h4293d15e};
test_weights[5024:5031] = '{32'hc27e74c7, 32'h4105c0d6, 32'h413d0444, 32'hc1315011, 32'h42908f21, 32'h40a0f564, 32'hc1f115b6, 32'h42b4350e};
test_bias[628:628] = '{32'hc232e473};
test_output[628:628] = '{32'h45d6c927};
test_input[5032:5039] = '{32'hc010a6ac, 32'h41209de9, 32'h42af63a6, 32'hc22b577e, 32'h42184706, 32'h42b53438, 32'hc2a9cad8, 32'hc20a14d8};
test_weights[5032:5039] = '{32'hc252ef39, 32'hc24ccf4b, 32'h41d54c83, 32'h41418583, 32'h42a39542, 32'hc28bfa35, 32'hc008c146, 32'h41f3c8b8};
test_bias[629:629] = '{32'hc25c7f50};
test_output[629:629] = '{32'hc52a7c92};
test_input[5040:5047] = '{32'hbf9a74f7, 32'h42276591, 32'hc2b69edf, 32'h41b3bb70, 32'hc1f44ed4, 32'h4144df36, 32'hc1cca31f, 32'hc2bdb260};
test_weights[5040:5047] = '{32'hc18c05f4, 32'hc28714c9, 32'hc1a024fa, 32'h418bbf83, 32'h4260b7f6, 32'hc0d0cfae, 32'hc28b674b, 32'h420bd5e0};
test_bias[630:630] = '{32'hc28c50aa};
test_output[630:630] = '{32'hc579005f};
test_input[5048:5055] = '{32'h41be91f9, 32'hc2ad595e, 32'h4201ef0b, 32'hc29cb540, 32'hc1968246, 32'hc18c0b4a, 32'hc28ceb76, 32'hc26f0e8d};
test_weights[5048:5055] = '{32'hc2a106bc, 32'h423552d8, 32'h41600ebd, 32'hc2c53ae5, 32'hc2998c89, 32'h42a735ad, 32'h42bdc99a, 32'hbfaa3d07};
test_bias[631:631] = '{32'h420bbd47};
test_output[631:631] = '{32'hc58500ee};
test_input[5056:5063] = '{32'h416d7760, 32'hc27785b9, 32'hc19f2e68, 32'h42ac3ecf, 32'h41b356b5, 32'hc1435b75, 32'hc1d7e9f8, 32'hc26ebd5f};
test_weights[5056:5063] = '{32'h420b7440, 32'hc23388dd, 32'hc22fd51d, 32'h4288b3d5, 32'hc25e825c, 32'hc219eea6, 32'hc206e759, 32'h425d6092};
test_bias[632:632] = '{32'hc17630f3};
test_output[632:632] = '{32'h45d6b4c8};
test_input[5064:5071] = '{32'h42a9b450, 32'h4280c826, 32'hc128d350, 32'h417c95d3, 32'h423b7b32, 32'h41b138eb, 32'h41cd5c8a, 32'hc2c28c91};
test_weights[5064:5071] = '{32'h4118613f, 32'hc2914a26, 32'hc29b38c1, 32'hc27c42f3, 32'h422ffb18, 32'h42b12910, 32'h418d9a81, 32'hbf42a18a};
test_bias[633:633] = '{32'h41c4fe93};
test_output[633:633] = '{32'h4404c623};
test_input[5072:5079] = '{32'hc2b6b4a2, 32'h42107103, 32'h4135b67b, 32'hc2071778, 32'h423a89cf, 32'h405e1c5e, 32'h42aa9e72, 32'h42ade066};
test_weights[5072:5079] = '{32'h429fdcf5, 32'hc281a1b4, 32'hc24738d5, 32'h4236b661, 32'hc2895216, 32'hc23dfc5b, 32'hc25c1310, 32'h42525865};
test_bias[634:634] = '{32'h422ef560};
test_output[634:634] = '{32'hc66d6ed4};
test_input[5080:5087] = '{32'h416381fc, 32'hc2c01143, 32'hc11fb8f0, 32'hc2836bb6, 32'hc2991959, 32'h41b950fc, 32'hc2954c44, 32'hc2248401};
test_weights[5080:5087] = '{32'hc2b16a95, 32'hc1c1aebb, 32'hc1931a69, 32'h41aa91ed, 32'h41f6e4c6, 32'h42642662, 32'h426c87f1, 32'hc2acf184};
test_bias[635:635] = '{32'h4200b493};
test_output[635:635] = '{32'hc4fc91e7};
test_input[5088:5095] = '{32'h42a62362, 32'h429ee17b, 32'hc2992e7c, 32'hc2a55181, 32'hc29a7616, 32'hc2396e72, 32'h420cb3f3, 32'hc17e4c6a};
test_weights[5088:5095] = '{32'h42568a7e, 32'hc286b5b3, 32'h42653ba5, 32'hc243ec1a, 32'hc23a430b, 32'hc2c2f3b4, 32'hc28ed4d0, 32'h41a15c99};
test_bias[636:636] = '{32'hc1956b67};
test_output[636:636] = '{32'h457bbd94};
test_input[5096:5103] = '{32'hc1f45400, 32'h4232d336, 32'hc0a06224, 32'h427f5fb5, 32'h41c52ca7, 32'hc26c94f4, 32'h420fc8f0, 32'hc20d3081};
test_weights[5096:5103] = '{32'hc1e348c7, 32'hc2c491f4, 32'hc1682fff, 32'hc2b95cad, 32'hc1e63c92, 32'hc2bdd413, 32'hc24862f0, 32'hc290155c};
test_bias[637:637] = '{32'h4252e9a7};
test_output[637:637] = '{32'hc56575e5};
test_input[5104:5111] = '{32'h424d6e5e, 32'h4280b23b, 32'h42495f92, 32'hc2b1629a, 32'h42450be7, 32'h42c5e0df, 32'h41a9a568, 32'hc187763b};
test_weights[5104:5111] = '{32'hc2a40076, 32'hc2a41254, 32'hc26bcd4a, 32'hc25bf950, 32'hc29afcf4, 32'hc2a9253c, 32'hc151ba5d, 32'hc22d5035};
test_bias[638:638] = '{32'h4255bce9};
test_output[638:638] = '{32'hc69670c7};
test_input[5112:5119] = '{32'h40ae8c87, 32'h42325e93, 32'hc2b962eb, 32'hc247048d, 32'hc2ad10e6, 32'h4266cabc, 32'h429fa4b5, 32'hc2c41401};
test_weights[5112:5119] = '{32'h419a9bf5, 32'hc2abaa47, 32'hc186df87, 32'hc204fe06, 32'h4206f45e, 32'h418e7931, 32'h429918b7, 32'h41d9403d};
test_bias[639:639] = '{32'h41644069};
test_output[639:639] = '{32'h44852193};
test_input[5120:5127] = '{32'h41ddce1f, 32'h417635a0, 32'h412f7409, 32'h4215bbc0, 32'h42487c4a, 32'hc1aca6ce, 32'hc29f516f, 32'hc241516c};
test_weights[5120:5127] = '{32'hc2b32f4c, 32'h415fabdb, 32'h425cf4f2, 32'h422bfc79, 32'h428f363b, 32'h428067a0, 32'hc1bb99bb, 32'hc2258cbd};
test_bias[640:640] = '{32'hc2856f19};
test_output[640:640] = '{32'h45b9fa59};
test_input[5128:5135] = '{32'h427e6595, 32'h423dcd18, 32'hc28d4964, 32'h42be9654, 32'h42038d7b, 32'hc2aaf879, 32'hc20a440d, 32'h42a51a55};
test_weights[5128:5135] = '{32'h4251bb40, 32'h425eeaf7, 32'h420c2a82, 32'h42ae8e70, 32'hc15090d6, 32'hc0f72441, 32'h4282d791, 32'hc191142f};
test_bias[641:641] = '{32'h3f94e8db};
test_output[641:641] = '{32'h46019ba7};
test_input[5136:5143] = '{32'hc21d8376, 32'h429956b0, 32'hc29f65fc, 32'hc194366e, 32'hc11350d0, 32'hc2b69e06, 32'h4267a408, 32'h42a5d5b8};
test_weights[5136:5143] = '{32'h417e8dbd, 32'hc26fab96, 32'hc1c2fa73, 32'h41e17ae8, 32'hc223b60f, 32'h42892c60, 32'hc2adf783, 32'h428f9523};
test_bias[642:642] = '{32'hc1d8e70d};
test_output[642:642] = '{32'hc6097579};
test_input[5144:5151] = '{32'hc2137a41, 32'hc283cc72, 32'h424c188e, 32'h4094d406, 32'hc28da492, 32'hc14f5f80, 32'hc23b0f87, 32'hc294bbac};
test_weights[5144:5151] = '{32'h420821b3, 32'hc1878f47, 32'h42808c91, 32'hc16551c4, 32'hc2b34e9b, 32'hc25edfe3, 32'hc254ab36, 32'h42130de8};
test_bias[643:643] = '{32'hc206e306};
test_output[643:643] = '{32'h461a23f9};
test_input[5152:5159] = '{32'hc2c1a036, 32'hc2aa33cc, 32'hc1aafe88, 32'h40f05a31, 32'hc21b66d2, 32'h42addd66, 32'h423f9cc6, 32'h42707007};
test_weights[5152:5159] = '{32'hc24af1f2, 32'h4291b005, 32'hc13f2660, 32'h42c47f92, 32'hc25843bc, 32'hc2447501, 32'hc29ff760, 32'h410505b7};
test_bias[644:644] = '{32'h4185f7c8};
test_output[644:644] = '{32'hc5b48f85};
test_input[5160:5167] = '{32'h429014b0, 32'hbfa984e1, 32'h42583d09, 32'h423640a1, 32'h42563239, 32'hc138ea88, 32'h40ff7dc2, 32'h429c18fd};
test_weights[5160:5167] = '{32'hc20a9051, 32'h425f9f46, 32'h428d07dc, 32'hc2079e0f, 32'h40ffa51d, 32'h3e7f115d, 32'hc2a00133, 32'hbfe11d2b};
test_bias[645:645] = '{32'hc282ecd4};
test_output[645:645] = '{32'hc433b96e};
test_input[5168:5175] = '{32'h421ff70e, 32'hc15c7d42, 32'h422c4860, 32'h42a62838, 32'hc28a0b51, 32'h423d2067, 32'h415dd7b8, 32'hc15b1fa7};
test_weights[5168:5175] = '{32'hc2a1ab98, 32'h428481f0, 32'hc2b365d8, 32'h422c9174, 32'hc1133888, 32'hc23b77cb, 32'h423ea75a, 32'h4291ed55};
test_bias[646:646] = '{32'hc27d1674};
test_output[646:646] = '{32'hc5c83b95};
test_input[5176:5183] = '{32'h42272654, 32'hc0399bf1, 32'h418a007c, 32'hc2363ebc, 32'h42179d14, 32'h4215df8d, 32'h42919382, 32'h42b2c0d2};
test_weights[5176:5183] = '{32'h423b9d0e, 32'hc2193075, 32'hc22d329c, 32'hc2508d01, 32'h42aa7a3b, 32'hc2beab51, 32'h42c1a9a4, 32'h40c80bd3};
test_bias[647:647] = '{32'hc28d07c8};
test_output[647:647] = '{32'h462a3b14};
test_input[5184:5191] = '{32'hc2891d3a, 32'h41a88cae, 32'hc292ed93, 32'hc2391c46, 32'hc1be9515, 32'h429515fe, 32'hc2bc017d, 32'h426bcb81};
test_weights[5184:5191] = '{32'hc234b366, 32'hc28a24da, 32'h423d06f7, 32'hc180f087, 32'h42b472e6, 32'hc2a0c772, 32'hc28ecf18, 32'hc2a46054};
test_bias[648:648] = '{32'h41e0b2f6};
test_output[648:648] = '{32'hc5e51355};
test_input[5192:5199] = '{32'hc232e445, 32'h42a3824f, 32'hc29be85e, 32'hc283fd52, 32'hc212898c, 32'h3f9a4f26, 32'hc29e0553, 32'h4117e342};
test_weights[5192:5199] = '{32'h418bfe0d, 32'hc2b82ad9, 32'hc2130c25, 32'hc2abdcd5, 32'h420a7c58, 32'h42a6b71f, 32'hc0fb3499, 32'hc261658b};
test_bias[649:649] = '{32'h421d69e8};
test_output[649:649] = '{32'hc44c523c};
test_input[5200:5207] = '{32'hc0db32af, 32'h423f2e98, 32'h40fd02ce, 32'hc1b2c55d, 32'h42795ae3, 32'h42a66727, 32'hc12f46d7, 32'hc2608adf};
test_weights[5200:5207] = '{32'h41a9bbc7, 32'hc255dd75, 32'hc2a0a690, 32'h42481e4c, 32'h4215dbfb, 32'hc0b01d4d, 32'hc20821ed, 32'hc2a806d1};
test_bias[650:650] = '{32'h42102bbb};
test_output[650:650] = '{32'h451f4c0e};
test_input[5208:5215] = '{32'h425e4936, 32'h42756f84, 32'hc2acde9e, 32'h42bf6842, 32'hc27ff677, 32'hc23e976d, 32'h41cc3ee5, 32'h416b303d};
test_weights[5208:5215] = '{32'hc2918f58, 32'h429df2cd, 32'hc28dca22, 32'hc2070c11, 32'hc1af24ef, 32'hc15ec2a5, 32'h420a5365, 32'hc28a9ede};
test_bias[651:651] = '{32'hc16740b0};
test_output[651:651] = '{32'h45af5f14};
test_input[5216:5223] = '{32'hc218e668, 32'hc2c6b2c6, 32'hc109d33d, 32'h423bfd3f, 32'hc235d113, 32'hc2a970fe, 32'hc1fe0018, 32'hc2ae2684};
test_weights[5216:5223] = '{32'hc25841f5, 32'h422dfc40, 32'hc1bd85e6, 32'h42b7abe1, 32'h4153448d, 32'hc19c09fa, 32'hc2395e92, 32'hc28573fc};
test_bias[652:652] = '{32'h41ed917a};
test_output[652:652] = '{32'h462613da};
test_input[5224:5231] = '{32'hc24852c6, 32'hc2603b82, 32'h428bd451, 32'h42247ef5, 32'h42a1faa4, 32'hc20173cf, 32'h42bcc39c, 32'h42b2404e};
test_weights[5224:5231] = '{32'hc2371c0b, 32'hc29e4db0, 32'hc222d856, 32'hc27db7d3, 32'h42153647, 32'h42995489, 32'hc289b53c, 32'hc2450608};
test_bias[653:653] = '{32'hc2a771c1};
test_output[653:653] = '{32'hc60f1568};
test_input[5232:5239] = '{32'hc29ebc73, 32'h42978538, 32'h408cade3, 32'h420da775, 32'h42958d57, 32'h42b6968d, 32'h41a0b94d, 32'h42c3015d};
test_weights[5232:5239] = '{32'h40c18679, 32'h40867c8e, 32'hc27eed29, 32'h42583aa2, 32'hc240fa85, 32'hc1883845, 32'h41feef23, 32'h42377007};
test_bias[654:654] = '{32'hc1088fd9};
test_output[654:654] = '{32'h44b0b439};
test_input[5240:5247] = '{32'hc21ce6f6, 32'h42c5660e, 32'hc2960c35, 32'hc13dcf7d, 32'hc03384ce, 32'hc2796c27, 32'h41bd5670, 32'h414b2ae4};
test_weights[5240:5247] = '{32'h4287613e, 32'h41ede32a, 32'h42778318, 32'h3e98f018, 32'h422eb3af, 32'h42ae0672, 32'h4190ffb4, 32'h42c5352b};
test_bias[655:655] = '{32'h42905cda};
test_output[655:655] = '{32'hc5ff092d};
test_input[5248:5255] = '{32'h42542a04, 32'hc141ea41, 32'hc28fd480, 32'hc2b8bf2b, 32'h40c9f409, 32'h4293bfc0, 32'h42c75142, 32'hc28f258d};
test_weights[5248:5255] = '{32'hc2b58651, 32'hc2ba6b9a, 32'h42168673, 32'h428afa0d, 32'h4177845d, 32'h42c55fef, 32'h42378f69, 32'hc2876fb4};
test_bias[656:656] = '{32'hc1b5e2b0};
test_output[656:656] = '{32'h45787f3e};
test_input[5256:5263] = '{32'hc167003d, 32'h41e8bec4, 32'h4210c073, 32'h42b060e2, 32'hc292caac, 32'h42c26fbd, 32'h42bad57b, 32'hc1dac261};
test_weights[5256:5263] = '{32'hc2867ecd, 32'hc2b217e3, 32'hc2b195e5, 32'hc2a5e10f, 32'hc2bd7a96, 32'h425104bb, 32'h42a2f3d9, 32'h42ba343a};
test_bias[657:657] = '{32'h42969524};
test_output[657:657] = '{32'h459d174f};
test_input[5264:5271] = '{32'h425f490e, 32'h420bf701, 32'h42bf8739, 32'h421fc91d, 32'hc2bf3dff, 32'h42b9abf7, 32'h42a01440, 32'hc281c6cb};
test_weights[5264:5271] = '{32'hc1e9589e, 32'h4260cce6, 32'h421d667a, 32'hc2a76690, 32'h42c13a73, 32'hc2aaf566, 32'hc2a58ced, 32'hc2c069b7};
test_bias[658:658] = '{32'h4233ff0e};
test_output[658:658] = '{32'hc682d8d8};
test_input[5272:5279] = '{32'h42a6d03e, 32'h423b6138, 32'h41cd973a, 32'h426ab6ec, 32'hc1e61c2c, 32'hc25e7329, 32'hc28e1433, 32'hc285ad83};
test_weights[5272:5279] = '{32'hc1f17769, 32'h42a52cbe, 32'h419c1ee1, 32'hc140d323, 32'h420f8b5e, 32'h42034d4c, 32'hc2864fe5, 32'h40bba5ac};
test_bias[659:659] = '{32'h42139ea5};
test_output[659:659] = '{32'h4528f9fb};
test_input[5280:5287] = '{32'h41d4fd37, 32'hc233d6a5, 32'h42ac38c4, 32'h42870440, 32'hc2041dd2, 32'h42498d57, 32'h42b0b322, 32'h42a7d74c};
test_weights[5280:5287] = '{32'hc24e415e, 32'hc231974f, 32'hc2b21b1d, 32'h42735aef, 32'h41777071, 32'hc2ba51e2, 32'hc2179f3c, 32'hc037d6ee};
test_bias[660:660] = '{32'hc22f3aaa};
test_output[660:660] = '{32'hc6380312};
test_input[5288:5295] = '{32'h42785c7e, 32'hc24ac068, 32'hc230ce59, 32'hc298b784, 32'h4170f49a, 32'h42ace065, 32'hc2bb511b, 32'hc22ccd38};
test_weights[5288:5295] = '{32'hc17d6c63, 32'h4288ede4, 32'hc1b9f44c, 32'h4217d3b8, 32'hc2009e7f, 32'hc2aca82c, 32'hc2ad77f3, 32'hc2b4826c};
test_bias[661:661] = '{32'h41dc7955};
test_output[661:661] = '{32'hc50acfda};
test_input[5296:5303] = '{32'hc28b3b78, 32'h41e3d808, 32'hc2c690a9, 32'h42c2d2d4, 32'hc13a5706, 32'hc1187266, 32'h4217012d, 32'h4224ec2d};
test_weights[5296:5303] = '{32'hc284aa24, 32'hc276bcc7, 32'h427f1ab9, 32'h41a644cd, 32'h42c30cba, 32'hc28648d1, 32'h40dccb1d, 32'hc1098ce2};
test_bias[662:662] = '{32'hc21fd7b1};
test_output[662:662] = '{32'hc501c4ca};
test_input[5304:5311] = '{32'h426d1e3d, 32'h41b199dd, 32'h429e3b65, 32'hc183fcc9, 32'hc279bf13, 32'hc20034c2, 32'hc294e251, 32'hc23daade};
test_weights[5304:5311] = '{32'h4112b9a5, 32'hc1d6440a, 32'hc292d89d, 32'h427c37ac, 32'h41e124c2, 32'h422ad0ec, 32'h42be362f, 32'h4169bfe2};
test_bias[663:663] = '{32'h42462641};
test_output[663:663] = '{32'hc68aaa51};
test_input[5312:5319] = '{32'h425c3deb, 32'h42c1db8b, 32'h41cba9b8, 32'h4123f2bb, 32'h4288e65b, 32'h425c1438, 32'hc27eebed, 32'hc2114e4e};
test_weights[5312:5319] = '{32'h42b62481, 32'h41fc1cd9, 32'h42887247, 32'h3f77ac4e, 32'hc2b7e89e, 32'hc21159c1, 32'h42b50283, 32'hc0b1af1a};
test_bias[664:664] = '{32'hc14f1d05};
test_output[664:664] = '{32'hc57d8ec5};
test_input[5320:5327] = '{32'h4154b675, 32'h4012f38e, 32'hc284dc3d, 32'h4101cef5, 32'hc2a0074e, 32'h41e3c18f, 32'hc184401c, 32'hc2bbfc08};
test_weights[5320:5327] = '{32'h42a042ef, 32'hc0caeaa9, 32'hc28a8e42, 32'h4288a362, 32'h4117b9a4, 32'hc23b4b5d, 32'h42ae12b4, 32'h428134f6};
test_bias[665:665] = '{32'hc2289e7f};
test_output[665:665] = '{32'hc556ddb0};
test_input[5328:5335] = '{32'hc2a4c32d, 32'h41c246ca, 32'h413edcce, 32'hc2a5105c, 32'hc2a42196, 32'h41ffde3d, 32'hc2b8cc26, 32'h4206f322};
test_weights[5328:5335] = '{32'h41b3df21, 32'h4188851e, 32'h42bae75d, 32'h41bcbefa, 32'h421f699d, 32'h420493d4, 32'hc1c1b663, 32'hc2a2930b};
test_bias[666:666] = '{32'hc2288e90};
test_output[666:666] = '{32'hc59d1fbf};
test_input[5336:5343] = '{32'hc187d5ee, 32'hc23a2366, 32'hc09ed01d, 32'hc0c29047, 32'h4274d047, 32'hc2b782f1, 32'hc1167caf, 32'h4290168a};
test_weights[5336:5343] = '{32'hc1fbcd8b, 32'h425f58a2, 32'hc2bd2490, 32'h42bed545, 32'h4197f571, 32'hc293a40d, 32'h4280dcd4, 32'h41f3afec};
test_bias[667:667] = '{32'h4240cf3a};
test_output[667:667] = '{32'h45e7303d};
test_input[5344:5351] = '{32'h41f24cbe, 32'h4293c815, 32'h41f0a644, 32'hc264109e, 32'hc24b955c, 32'h4255eb0d, 32'hc25842e0, 32'h41d2e903};
test_weights[5344:5351] = '{32'h4262fa08, 32'hc20d62a1, 32'h42a19956, 32'hc1ff2ae6, 32'h41f59deb, 32'h41e6f4b8, 32'h42b36bc5, 32'h3f9ac7aa};
test_bias[668:668] = '{32'h421ef3d8};
test_output[668:668] = '{32'hc4b42942};
test_input[5352:5359] = '{32'h42b38246, 32'h42244d26, 32'h42567681, 32'hc247c7ce, 32'h42613eeb, 32'hc21d59e7, 32'hc2c00c54, 32'h42b3a6cb};
test_weights[5352:5359] = '{32'h41fc6a40, 32'hc2a9cabe, 32'hc293760a, 32'hc2bc15f8, 32'h422fb40f, 32'h41fa6388, 32'hc2889a25, 32'h41de8c40};
test_bias[669:669] = '{32'h41c90d08};
test_output[669:669] = '{32'h4622b5d9};
test_input[5360:5367] = '{32'hc10fd63d, 32'hc201a439, 32'hc2b1c52e, 32'hc23d317f, 32'hc28345ac, 32'hc287159a, 32'hc2864289, 32'h41f3e589};
test_weights[5360:5367] = '{32'h42850a4a, 32'h426da5ff, 32'h425fe27b, 32'h42a10853, 32'h429d0e94, 32'hc2299c4c, 32'h42683910, 32'h42557654};
test_bias[670:670] = '{32'h41c7d981};
test_output[670:670] = '{32'hc6778a20};
test_input[5368:5375] = '{32'hc29b1e5e, 32'hc26e874f, 32'hc1fc62c6, 32'hc2b22f77, 32'hc21dd28d, 32'hc2b2e8e8, 32'hc2a24e15, 32'h42780f8c};
test_weights[5368:5375] = '{32'h41c3ab84, 32'h425c1ac1, 32'h41ef1ae4, 32'h42c7a6f0, 32'h42bee5c4, 32'hc2be7a14, 32'hc08cb976, 32'hc298613d};
test_bias[671:671] = '{32'h42883c35};
test_output[671:671] = '{32'hc663859a};
test_input[5376:5383] = '{32'hc1a18716, 32'hc2a3ea59, 32'hc1ae57cf, 32'hc224cdaa, 32'h41dd4ddc, 32'h428643c9, 32'h425df191, 32'hc1d233ba};
test_weights[5376:5383] = '{32'hc26bc78c, 32'hc2985c36, 32'h415e81e2, 32'h4299a686, 32'hc1915c23, 32'hc2c72eeb, 32'hc1175699, 32'hc0f25ba6};
test_bias[672:672] = '{32'hc25a252a};
test_output[672:672] = '{32'hc5613734};
test_input[5384:5391] = '{32'h42a7eac4, 32'hc2c3e246, 32'hc261872d, 32'hc225a47a, 32'hc14e9922, 32'hc2a39da3, 32'h41e18250, 32'hc2b49cd6};
test_weights[5384:5391] = '{32'hc2938c78, 32'hc2069788, 32'hc204ad00, 32'hc169e54e, 32'hc27a6aac, 32'h41bcb954, 32'hc1a235cc, 32'hc2a87970};
test_bias[673:673] = '{32'h427d85ba};
test_output[673:673] = '{32'h45ad940d};
test_input[5392:5399] = '{32'hc217244d, 32'hc2943c59, 32'hc25a3581, 32'h426f663b, 32'h42602814, 32'h4298ffa8, 32'h41ea9ce5, 32'h42c0554a};
test_weights[5392:5399] = '{32'hc2c1c766, 32'hc17d7d14, 32'h42ad0688, 32'hc10b707d, 32'h42312bb1, 32'h427e74c0, 32'hc265fca4, 32'hc2667b1e};
test_bias[674:674] = '{32'h406f0a51};
test_output[674:674] = '{32'hc38c6a0a};
test_input[5400:5407] = '{32'h4215c029, 32'h4194a644, 32'hc1ab5988, 32'hc2aea8b5, 32'hc290ca43, 32'h3da56a88, 32'h41e67973, 32'hc23dfd43};
test_weights[5400:5407] = '{32'h41c69bd9, 32'hc200a97c, 32'hc1264bcb, 32'hc118883d, 32'hc1edcbbf, 32'h427db0fc, 32'hc29a8393, 32'h428ec48a};
test_bias[675:675] = '{32'h41a66451};
test_output[675:675] = '{32'hc5003870};
test_input[5408:5415] = '{32'hc29e60d7, 32'h423f3f61, 32'hc258b3f5, 32'h41bf41dd, 32'h428f5151, 32'h41d401ad, 32'h42a2e0c8, 32'hc2a61963};
test_weights[5408:5415] = '{32'h4289b427, 32'h4228d5ff, 32'h423cd4ba, 32'hc2426653, 32'hc280da27, 32'h41b2cc90, 32'h41071e64, 32'hbf4ab006};
test_bias[676:676] = '{32'h42b68f9f};
test_output[676:676] = '{32'hc6217505};
test_input[5416:5423] = '{32'h411b73b6, 32'hc2ac98b2, 32'h42b541ac, 32'hc22adc85, 32'hc0a1df63, 32'h4233a75c, 32'h42c15db3, 32'h419fe254};
test_weights[5416:5423] = '{32'h42883958, 32'hc2baffc6, 32'hc2b44bd8, 32'hc22f37d3, 32'hc29f36b3, 32'h41a2a640, 32'h42aeeb05, 32'h422bd4b4};
test_bias[677:677] = '{32'h421c2aa5};
test_output[677:677] = '{32'h464cb3e4};
test_input[5424:5431] = '{32'hc1d9a852, 32'hc2504091, 32'h42beb3a4, 32'h4281cff7, 32'hc2a436a7, 32'hc2bdc1af, 32'hc1e70160, 32'h4206fdb0};
test_weights[5424:5431] = '{32'hc1411786, 32'h424e6976, 32'hc29fa26c, 32'hc2af30c8, 32'h418c5b86, 32'hc040a72a, 32'h42857530, 32'h42b5d317};
test_bias[678:678] = '{32'h422f27ec};
test_output[678:678] = '{32'hc6742124};
test_input[5432:5439] = '{32'hc2962222, 32'hc2a884c4, 32'h41e40548, 32'h41d86987, 32'h41f310c2, 32'hc24d8396, 32'h42b7d375, 32'hc1e2cbc2};
test_weights[5432:5439] = '{32'hc24c349e, 32'hc299b184, 32'hc2bb0be7, 32'h41bc0ada, 32'hc2b56760, 32'hc29d00df, 32'h42a9c9bb, 32'hc29bb8a4};
test_bias[679:679] = '{32'h4285dfb5};
test_output[679:679] = '{32'h46996036};
test_input[5440:5447] = '{32'hc280edbe, 32'hc158b2ec, 32'h42c3a720, 32'hc25c4fc4, 32'h41bbd3bc, 32'h4018d8ce, 32'hc183063b, 32'h4039d613};
test_weights[5440:5447] = '{32'h423a37a2, 32'h4261f534, 32'h42901ee9, 32'hc136dd8f, 32'hc2731df3, 32'hc10814fe, 32'hc195d913, 32'h4275e186};
test_bias[680:680] = '{32'hc26e7c0a};
test_output[680:680] = '{32'h4534b10a};
test_input[5448:5455] = '{32'hc2843b1e, 32'hc2791816, 32'hc2163612, 32'hc226476a, 32'h415511dd, 32'h4295740b, 32'h42c7063b, 32'hc2bfbebf};
test_weights[5448:5455] = '{32'h41187426, 32'h4162eb1d, 32'hc0f319ec, 32'hc2a777db, 32'h42b29279, 32'h422f76a4, 32'hc2a4ce79, 32'hc2a82359};
test_bias[681:681] = '{32'hc2961eea};
test_output[681:681] = '{32'h45cb44ec};
test_input[5456:5463] = '{32'h4263f891, 32'h42c38681, 32'hc297ac8a, 32'hc2a7d756, 32'h4271b05e, 32'hc1705394, 32'hc287fbe4, 32'h42c18e55};
test_weights[5456:5463] = '{32'hc20bbaf5, 32'h428c68dd, 32'hc23055e3, 32'hc26a4ad0, 32'hc1f4c436, 32'hc1983de1, 32'h411f0d8b, 32'hc2b83064};
test_bias[682:682] = '{32'hc2873177};
test_output[682:682] = '{32'h44ef0490};
test_input[5464:5471] = '{32'hc2860813, 32'h4236ffae, 32'hc28bed9c, 32'h414802cf, 32'hc27c27e0, 32'h42232a3b, 32'h425eaf8a, 32'h41e04cd9};
test_weights[5464:5471] = '{32'hc18486e0, 32'h426234bc, 32'h401f7ffc, 32'h41fa672b, 32'hc09b8757, 32'h4293a0c7, 32'hc2939749, 32'hc2bf6134};
test_bias[683:683] = '{32'h42922f18};
test_output[683:683] = '{32'h44006269};
test_input[5472:5479] = '{32'hc2970df6, 32'hc29ef06a, 32'hc26ded06, 32'h4287db78, 32'h4086d4de, 32'h415db6cf, 32'hc299e3a2, 32'h42854afe};
test_weights[5472:5479] = '{32'h42b1385e, 32'h425690ba, 32'h4293e3b4, 32'hc2183f13, 32'hc1bf65ed, 32'hc28c020a, 32'hc2455318, 32'h4279a63f};
test_bias[684:684] = '{32'hc28cd170};
test_output[684:684] = '{32'hc62dd459};
test_input[5480:5487] = '{32'hc2981bc1, 32'h42a74613, 32'h4289f2a4, 32'h41f37f1d, 32'h4229d148, 32'h420f2ab2, 32'hc2b34957, 32'hc1357f93};
test_weights[5480:5487] = '{32'hc1fb62fa, 32'h42648e36, 32'h42461dbe, 32'hc1ed9543, 32'h42a0e473, 32'h42673fd5, 32'hc200f036, 32'hc2bc1048};
test_bias[685:685] = '{32'h3faf7bf2};
test_output[685:685] = '{32'h46956675};
test_input[5488:5495] = '{32'h422e1b02, 32'h425a0ba9, 32'hc099302a, 32'h4181e1bc, 32'hc213427e, 32'h423328ca, 32'hc278a122, 32'hc28cde56};
test_weights[5488:5495] = '{32'h42b8cbc0, 32'h42a3e01c, 32'h4179ec93, 32'h42612c92, 32'h428f546a, 32'h41bee724, 32'h424a10ec, 32'hc2c6572b};
test_bias[686:686] = '{32'hc29291f4};
test_output[686:686] = '{32'h46342697};
test_input[5496:5503] = '{32'h428cec7e, 32'h4203b04d, 32'h429c2688, 32'h424d70ae, 32'hc237ccf6, 32'h418d94d1, 32'hc2875a1d, 32'hc0c4bd7b};
test_weights[5496:5503] = '{32'h4225df2b, 32'hc2b1283a, 32'hbfb21c54, 32'hc2ae65f5, 32'hc1f7db70, 32'hc2477210, 32'hc2abce4e, 32'h42277c07};
test_bias[687:687] = '{32'hc0b04de7};
test_output[687:687] = '{32'h44bccb46};
test_input[5504:5511] = '{32'hc0e5fbae, 32'h418cb8e5, 32'h42bb4c9d, 32'hc07ea935, 32'hc2a1cfb5, 32'h42873764, 32'h42a6bb59, 32'hbf3b89bd};
test_weights[5504:5511] = '{32'hc209b7b1, 32'hc277ebc7, 32'h427c1fce, 32'h420c085a, 32'h424f21a0, 32'hc255c33a, 32'h42982817, 32'h42819dbc};
test_bias[688:688] = '{32'h42adb5fe};
test_output[688:688] = '{32'h455abe4d};
test_input[5512:5519] = '{32'h429f0063, 32'hc1a47962, 32'h426c7187, 32'h42508d0b, 32'h4254d0a9, 32'hc2c2ff3e, 32'h4156eacd, 32'hc2584c55};
test_weights[5512:5519] = '{32'hc29b9c9e, 32'hc060a6ff, 32'h41f39310, 32'hc26b9876, 32'hc2a86571, 32'h41b958d7, 32'hc253e261, 32'hc1cd3c51};
test_bias[689:689] = '{32'h42849714};
test_output[689:689] = '{32'hc6511462};
test_input[5520:5527] = '{32'h4235c3dd, 32'hc25c0ac0, 32'h3f305012, 32'h40c4bc82, 32'hc23e75dc, 32'h418c2e2a, 32'hc08451c9, 32'hc238e8dd};
test_weights[5520:5527] = '{32'h41342320, 32'h42670fd2, 32'hc2a47d3f, 32'hc2a7ee52, 32'hc2c17723, 32'hc2ba6b5d, 32'hc2350ab6, 32'hc28e6092};
test_bias[690:690] = '{32'hc2403170};
test_output[690:690] = '{32'h4545baab};
test_input[5528:5535] = '{32'hc2125dc1, 32'h41caec69, 32'hc2817351, 32'h426f494e, 32'h42078b0c, 32'hc284ce42, 32'hc1c69f44, 32'hc2111042};
test_weights[5528:5535] = '{32'h420fb6c3, 32'hc1fc12c9, 32'h40a8a695, 32'hc2c14dac, 32'h42012ce0, 32'h42af3a2d, 32'h41dcf704, 32'hc23adfaa};
test_bias[691:691] = '{32'hc26eb7de};
test_output[691:691] = '{32'hc63bae34};
test_input[5536:5543] = '{32'h420c484d, 32'h429779f6, 32'hc19606c6, 32'h42823233, 32'h42bdb9bc, 32'hc283f983, 32'hc09d437e, 32'hc1098685};
test_weights[5536:5543] = '{32'h42abedeb, 32'hc122800b, 32'h428ceda7, 32'h4087ef62, 32'hc1a35aa7, 32'h41ca2277, 32'h424fad03, 32'h423e59a5};
test_bias[692:692] = '{32'hc253a9ab};
test_output[692:692] = '{32'hc5430b48};
test_input[5544:5551] = '{32'h41067b99, 32'hc29d0b85, 32'hc28615ef, 32'h4249d5f5, 32'h42a56f3f, 32'h42230c21, 32'h429b4cf7, 32'hc20db24a};
test_weights[5544:5551] = '{32'h420c5e8f, 32'h41ab17af, 32'h429a8212, 32'h4297ef6a, 32'h42288bef, 32'hc2c1802b, 32'h415d18e4, 32'h41d64d37};
test_bias[693:693] = '{32'h42a41a85};
test_output[693:693] = '{32'hc53a69be};
test_input[5552:5559] = '{32'h4265f546, 32'h428944a2, 32'hc127fd0f, 32'hc28b1fc6, 32'h4153e43a, 32'h4149b444, 32'hc298fe95, 32'h427b5906};
test_weights[5552:5559] = '{32'h42ac9294, 32'hc2b2242a, 32'h41468c18, 32'h42b6f4ca, 32'h42b0a402, 32'h42938b5d, 32'hc2b568ef, 32'hc1a7c8cf};
test_bias[694:694] = '{32'hc1f48355};
test_output[694:694] = '{32'h422de3ea};
test_input[5560:5567] = '{32'h407b9846, 32'h4205b836, 32'hc2ab87a9, 32'hc2b742a3, 32'h42135fef, 32'hc186313b, 32'h421d684d, 32'h4210f8fc};
test_weights[5560:5567] = '{32'h415dac67, 32'h40b132af, 32'hc15a06e0, 32'hc1e69e16, 32'h413dac46, 32'hc221ca5b, 32'hc26efefb, 32'h4096f5ac};
test_bias[695:695] = '{32'h420522d5};
test_output[695:695] = '{32'h453c9f95};
test_input[5568:5575] = '{32'hc287ee99, 32'hc28f641d, 32'h41bb2d06, 32'hc23bafa0, 32'hc2a4d005, 32'h406c4433, 32'h422085a5, 32'hc2aa9d5c};
test_weights[5568:5575] = '{32'h41faad77, 32'hc2aebe80, 32'hc1d98feb, 32'h429ed2e8, 32'h420381c4, 32'h4299d14d, 32'hc2a239d1, 32'hc246e476};
test_bias[696:696] = '{32'hc28e4249};
test_output[696:696] = '{32'hc4d93795};
test_input[5576:5583] = '{32'hc187b1aa, 32'hc2531a63, 32'h421bd5df, 32'hc2575bd4, 32'h42c79808, 32'hc2c1fe59, 32'h41cd9241, 32'hc26f13fc};
test_weights[5576:5583] = '{32'hc17cc14d, 32'hc2934394, 32'hc17aa4bb, 32'h424f9e37, 32'hc2add0ef, 32'hc28c2684, 32'h41cd0a6a, 32'hc28c9642};
test_bias[697:697] = '{32'h4180fda7};
test_output[697:697] = '{32'h456a5279};
test_input[5584:5591] = '{32'hc2c1f8c3, 32'h42ada0cd, 32'h427cee45, 32'h42991c32, 32'h4294f752, 32'h426fe968, 32'h41e728bf, 32'h4280de63};
test_weights[5584:5591] = '{32'hc10e9f25, 32'h42637ac3, 32'h4232da2c, 32'hc1e357f3, 32'hc069d021, 32'h429d65cf, 32'h4253eff6, 32'hc1b75648};
test_bias[698:698] = '{32'h42b8cdca};
test_output[698:698] = '{32'h462ca0e6};
test_input[5592:5599] = '{32'hc2500b1d, 32'hc28571e1, 32'h41ec8911, 32'h41f23d7f, 32'h42b5ba4e, 32'hc19aaabe, 32'h4275a3d9, 32'hc2816acc};
test_weights[5592:5599] = '{32'hc1da4b02, 32'hc2a93cae, 32'hc268bac8, 32'hc1ab9e7e, 32'hc2a14c53, 32'hc2447b4c, 32'h429ae1ac, 32'h41e22099};
test_bias[699:699] = '{32'hc27a3c9f};
test_output[699:699] = '{32'h44939d01};
test_input[5600:5607] = '{32'hc28bc9cb, 32'hc1e602ae, 32'h4256bffe, 32'h4167e4b9, 32'hc23cbdd0, 32'h4271ecb1, 32'h417c8b4e, 32'hc1e4fa59};
test_weights[5600:5607] = '{32'h429f1b10, 32'h42a47a1f, 32'hc124d715, 32'h40af6372, 32'hc2b0b9b4, 32'h4266b44d, 32'hc260ddbc, 32'h40ea1004};
test_bias[700:700] = '{32'hc2a1b955};
test_output[700:700] = '{32'hc4efc711};
test_input[5608:5615] = '{32'hc13f1481, 32'h41e2a91b, 32'hc28f0bb2, 32'hc286ac33, 32'hc1fd76ab, 32'hc02b3709, 32'hc2828ace, 32'h421fe906};
test_weights[5608:5615] = '{32'hc27cbf9a, 32'h428929a1, 32'h42b081d3, 32'hc250c1aa, 32'h42bca2ca, 32'hc28518b9, 32'h42a590d9, 32'hc23c9e40};
test_bias[701:701] = '{32'h4205b0d9};
test_output[701:701] = '{32'hc61ed5fb};
test_input[5616:5623] = '{32'hc2605df7, 32'h422c4c29, 32'hc295d040, 32'hc1b3e3ff, 32'h3f7f47cf, 32'hc1c88dcd, 32'hc237dce0, 32'h427ae7e0};
test_weights[5616:5623] = '{32'h4206b278, 32'hc1d4e664, 32'hc1f9d3ad, 32'hc207f124, 32'hc21afd2b, 32'hc125a9af, 32'h424c407f, 32'hc28e0ae9};
test_bias[702:702] = '{32'hc112b546};
test_output[702:702] = '{32'hc5cbd05d};
test_input[5624:5631] = '{32'hc24e8d84, 32'hc1bb657a, 32'hc2a21abb, 32'h42c5c393, 32'h414b6674, 32'h42928179, 32'h423dcfe5, 32'h42a714e0};
test_weights[5624:5631] = '{32'h426bba49, 32'hc2a35b73, 32'h42aef746, 32'hc2a612da, 32'h4263310a, 32'h42af3b59, 32'hc228d905, 32'h42c691b7};
test_bias[703:703] = '{32'h42669d2f};
test_output[703:703] = '{32'hc537e579};
test_input[5632:5639] = '{32'hc2009e9a, 32'hc287075a, 32'hc1dba27e, 32'h42729906, 32'h425e5e8c, 32'h416e1498, 32'hc0e9ac86, 32'hbfc0c688};
test_weights[5632:5639] = '{32'hc236ecf6, 32'h4266977d, 32'hc18309c6, 32'h41ee67b7, 32'h42b30b6b, 32'h40036846, 32'h4117f8d4, 32'hc1a1d0fa};
test_bias[704:704] = '{32'hc0954efd};
test_output[704:704] = '{32'h4595fa0d};
test_input[5640:5647] = '{32'hbfc1d014, 32'hc1e7bdd2, 32'h42c252e3, 32'h4184cd17, 32'hc28249e6, 32'hc2c552e3, 32'h4201a1db, 32'h41223878};
test_weights[5640:5647] = '{32'h4295b9c2, 32'hc206844c, 32'h424bb5d1, 32'h42813007, 32'h42a9f073, 32'h41ec9542, 32'h4267baf0, 32'h428a1ab8};
test_bias[705:705] = '{32'hc17c09fe};
test_output[705:705] = '{32'h44778782};
test_input[5648:5655] = '{32'h429b83db, 32'hc29c7b42, 32'hc2af7b7d, 32'hc26ff395, 32'hc225a9b7, 32'h424676f6, 32'h422dd5d0, 32'h426e514d};
test_weights[5648:5655] = '{32'hc2119d84, 32'h418ca98f, 32'hc28a4039, 32'h428f0eb0, 32'hc25ae278, 32'h415b0900, 32'hbdb5781f, 32'hc285971d};
test_bias[706:706] = '{32'hc28268c0};
test_output[706:706] = '{32'hc55cf30a};
test_input[5656:5663] = '{32'h423831e0, 32'h40fd4c71, 32'hc1eac3d5, 32'h4244976d, 32'h41122450, 32'hc2b4e96c, 32'h41904792, 32'hc177a9be};
test_weights[5656:5663] = '{32'h428cbfae, 32'h412f8eed, 32'h42788a5a, 32'hbfa76068, 32'hc02754c1, 32'hc2a25634, 32'h42c20f7c, 32'hc2aba0ab};
test_bias[707:707] = '{32'h42164b00};
test_output[707:707] = '{32'h463987bb};
test_input[5664:5671] = '{32'h42551e82, 32'h426dc9ad, 32'hc2adadc0, 32'hc2c195f1, 32'h4280a799, 32'h42b6e49b, 32'h41b9f0bc, 32'hc1cc608a};
test_weights[5664:5671] = '{32'h42ac2f0d, 32'hc2c5c955, 32'h42218ef3, 32'hc25ce1e5, 32'hc1d2d300, 32'hc1c0f3e3, 32'hc27b2113, 32'h42970483};
test_bias[708:708] = '{32'h4229d4b3};
test_output[708:708] = '{32'hc5d1681a};
test_input[5672:5679] = '{32'hc2b7ad00, 32'hc28942ae, 32'hc2644168, 32'h423c1add, 32'hc29741b4, 32'h42049c7d, 32'hc22c49d7, 32'h407f0957};
test_weights[5672:5679] = '{32'hc2c3cb2d, 32'hc244d0d5, 32'h42bbe60a, 32'hc29a856f, 32'h42b59c0d, 32'h426f1cf6, 32'h422d23ef, 32'hc238d75c};
test_bias[709:709] = '{32'hc1f898ed};
test_output[709:709] = '{32'hc5608112};
test_input[5680:5687] = '{32'hc195a174, 32'h428a982c, 32'h3fb0e725, 32'h42a3e91f, 32'hc29c6f69, 32'hc1c4c7c8, 32'h42bb9af3, 32'hc1f61eb8};
test_weights[5680:5687] = '{32'hc2b6dd42, 32'hc09a6ec0, 32'h426987c1, 32'hc2a8a373, 32'h3f74d35f, 32'hc11d8be3, 32'h4211ba5c, 32'hc2bb657f};
test_bias[710:710] = '{32'hc2bb8300};
test_output[710:710] = '{32'h4465eab1};
test_input[5688:5695] = '{32'h42937139, 32'h40eda9cb, 32'hc1891b6e, 32'h422bb87e, 32'hc278df40, 32'h4235a882, 32'hc2084367, 32'h4271be8a};
test_weights[5688:5695] = '{32'hc153131f, 32'h428e9305, 32'hc2ad9bab, 32'hc1691058, 32'hc0b0df86, 32'hc2384951, 32'hc25b77c4, 32'hc1f264a3};
test_bias[711:711] = '{32'h42a726ae};
test_output[711:711] = '{32'hc496f59e};
test_input[5696:5703] = '{32'h42b745ef, 32'hc21670e1, 32'h41f13996, 32'h3f47fd75, 32'h42a14947, 32'hc2571817, 32'hc2afba6b, 32'hc28600c8};
test_weights[5696:5703] = '{32'hc28ff510, 32'h41eaa457, 32'h41b73c55, 32'hc265f3e3, 32'hc169ac30, 32'h42bb4ed8, 32'h42907d5b, 32'hc09afb5c};
test_bias[712:712] = '{32'hc16f04c0};
test_output[712:712] = '{32'hc696d295};
test_input[5704:5711] = '{32'h42bae842, 32'hc19f6b87, 32'hc2b49050, 32'hc10a5523, 32'hc282678b, 32'h429cf815, 32'hc2177f0d, 32'h4159c3fa};
test_weights[5704:5711] = '{32'hc231cd50, 32'h426c1fc0, 32'h42c30e08, 32'hc19d56be, 32'h412abce2, 32'h4206e544, 32'hc2147879, 32'h42ac7389};
test_bias[713:713] = '{32'hc2895045};
test_output[713:713] = '{32'hc6147e5e};
test_input[5712:5719] = '{32'hc2bfa72c, 32'h427bcd2e, 32'hc289a6ed, 32'hc2bc81f2, 32'hc1e2d6ef, 32'h4297d992, 32'hc27571e8, 32'h425ac4ee};
test_weights[5712:5719] = '{32'hc2471a26, 32'hc2677bbe, 32'h42c569ee, 32'h42b3ba69, 32'h42662ffa, 32'h42833358, 32'hc2932ecb, 32'hc1dfca71};
test_bias[714:714] = '{32'h427e232a};
test_output[714:714] = '{32'hc5f1d4e5};
test_input[5720:5727] = '{32'hc287f926, 32'hc1ad975d, 32'hc1dc4bf7, 32'h42a78041, 32'hc02468e9, 32'h42b982a5, 32'h41cb2714, 32'h421b7493};
test_weights[5720:5727] = '{32'h409f48ed, 32'h4181d5d1, 32'h41c2d57e, 32'h41cf032c, 32'h426dbe5e, 32'hc2aed07c, 32'h4287545a, 32'hc1e9ef91};
test_bias[715:715] = '{32'hc236403c};
test_output[715:715] = '{32'hc5d82f78};
test_input[5728:5735] = '{32'hbff30289, 32'h41b16beb, 32'hc1c4b140, 32'hc2bf7264, 32'hc295783f, 32'h42414fdc, 32'hc2a9984f, 32'h421bfca8};
test_weights[5728:5735] = '{32'h405afc29, 32'h4110f318, 32'hc2346fa5, 32'hc2992130, 32'h4271e5c6, 32'hc242bf0e, 32'hc2bebbc5, 32'h426c7c4d};
test_bias[716:716] = '{32'hc1d4a48f};
test_output[716:716] = '{32'h463d7791};
test_input[5736:5743] = '{32'hc005675b, 32'hc2929c0b, 32'hc15bdacd, 32'hbf1679fc, 32'h42249af1, 32'h4157b717, 32'hc2b5b642, 32'hc2409730};
test_weights[5736:5743] = '{32'h41f9badc, 32'h42a9fb20, 32'hc2c48d93, 32'h421157cc, 32'h40edf25b, 32'h420378e4, 32'h41276552, 32'hc191397d};
test_bias[717:717] = '{32'h42c7e452};
test_output[717:717] = '{32'hc5830d70};
test_input[5744:5751] = '{32'h42795360, 32'hc1d2c518, 32'h423969f0, 32'hc2a04af6, 32'h422102cc, 32'hc2c6109d, 32'hc2b234ef, 32'hc268613c};
test_weights[5744:5751] = '{32'hc297c6c6, 32'h427fb399, 32'hc260bf8c, 32'h42b58d07, 32'hc2085fc4, 32'h4090e5a4, 32'h427a8ecb, 32'h41f613d2};
test_bias[718:718] = '{32'h42c269d9};
test_output[718:718] = '{32'hc6c6544b};
test_input[5752:5759] = '{32'h41df5d5f, 32'h42151b34, 32'h423736ec, 32'h42aa2d8d, 32'hc1c86d32, 32'h42c6aa80, 32'h421c674e, 32'hc201c99f};
test_weights[5752:5759] = '{32'h424a208c, 32'h424a3e85, 32'h42109602, 32'h42503bb1, 32'h40c1aeba, 32'h428ac535, 32'hc1ad6e94, 32'h421f4d95};
test_bias[719:719] = '{32'hc2893ce2};
test_output[719:719] = '{32'h465963c1};
test_input[5760:5767] = '{32'hc1afce41, 32'h429bd332, 32'hc2597abc, 32'hc244e6ac, 32'h42bb7b6b, 32'hc2aae22c, 32'h42b7f7a0, 32'hc260094f};
test_weights[5760:5767] = '{32'hc1d45fbd, 32'hc2b5a080, 32'h4224399a, 32'hc2c15a32, 32'hc2ada374, 32'hc2971014, 32'hc1d8ba1b, 32'h42159cd8};
test_bias[720:720] = '{32'hc22c2cd6};
test_output[720:720] = '{32'hc620a137};
test_input[5768:5775] = '{32'hc2a8af43, 32'h420688f1, 32'hc21e15b4, 32'h425249f2, 32'h413031e7, 32'hc2485257, 32'hc1b4e9bb, 32'h42a8a1a7};
test_weights[5768:5775] = '{32'hc0c08419, 32'h4260982d, 32'hc1925bda, 32'h42bbac8f, 32'h42bc9570, 32'hc22cfefc, 32'hc2a61a16, 32'hc1608d91};
test_bias[721:721] = '{32'h423aff18};
test_output[721:721] = '{32'h463b77ee};
test_input[5776:5783] = '{32'hc27793da, 32'hc2c5a589, 32'hc13cc51d, 32'h429b95b9, 32'hc1d28dc7, 32'hbf85010f, 32'h42239edb, 32'hc2a7d321};
test_weights[5776:5783] = '{32'hc0a17103, 32'h4205d0d1, 32'hc2a5339f, 32'hc2a5562b, 32'h42bc37a7, 32'h42488a83, 32'h42add6b7, 32'h4231b744};
test_bias[722:722] = '{32'h428c9f70};
test_output[722:722] = '{32'hc62d262d};
test_input[5784:5791] = '{32'hc271835d, 32'h41c66ca4, 32'h40f92e76, 32'h42663a2c, 32'h42aaeda5, 32'hc2c56092, 32'hc22ce6a0, 32'h42255b7b};
test_weights[5784:5791] = '{32'hc27da2c6, 32'h42ac275a, 32'hc1cce98e, 32'hc1a88423, 32'h42227207, 32'hc143db2e, 32'h4234711b, 32'h42b2f1b2};
test_bias[723:723] = '{32'hc25a0898};
test_output[723:723] = '{32'h462ab32b};
test_input[5792:5799] = '{32'h423521b3, 32'hc283b4ac, 32'h42c16242, 32'hc2bc2530, 32'hc1f6dbf8, 32'h42bed4d0, 32'h41deff81, 32'h42b9e356};
test_weights[5792:5799] = '{32'h42ba2d52, 32'hc1f322cc, 32'hc22e6509, 32'h42be6518, 32'h42b6e206, 32'hc2971dcc, 32'hc265b25c, 32'hc2488df7};
test_bias[724:724] = '{32'hc287fedf};
test_output[724:724] = '{32'hc6b6247d};
test_input[5800:5807] = '{32'h4217cf0e, 32'hc20da118, 32'h425d875e, 32'hc1a272ae, 32'hc29a8f7d, 32'h4247ba87, 32'h42090816, 32'hc235a55c};
test_weights[5800:5807] = '{32'hc2a3cdc1, 32'hc12c7ddf, 32'h421c5cfc, 32'hc2828b6c, 32'hc2c21912, 32'hc2b44bf4, 32'hc2657469, 32'hc21758b4};
test_bias[725:725] = '{32'hc22c62e4};
test_output[725:725] = '{32'h4559057c};
test_input[5808:5815] = '{32'h42a848f5, 32'h427ad462, 32'h42267476, 32'hc286c035, 32'h411750f7, 32'h420ae176, 32'hc1b00242, 32'h403956e0};
test_weights[5808:5815] = '{32'hc2b8165c, 32'h409a7bed, 32'hc293dd92, 32'hc1b68ba7, 32'hc1e9c3dd, 32'h42a1865f, 32'h40ae9320, 32'h42a4eb4b};
test_bias[726:726] = '{32'h418ff17d};
test_output[726:726] = '{32'hc5c5664a};
test_input[5816:5823] = '{32'h41f31782, 32'hc287e996, 32'hc2bf6974, 32'h41ba18dc, 32'h4226fba7, 32'h42883381, 32'hc24af139, 32'hc1c11f15};
test_weights[5816:5823] = '{32'h41881ed9, 32'hc2658c75, 32'h428b3d1f, 32'hc292a0ec, 32'hc27fa744, 32'hc242ad72, 32'hc0040f21, 32'hc1051a46};
test_bias[727:727] = '{32'h41fde863};
test_output[727:727] = '{32'hc615f37c};
test_input[5824:5831] = '{32'h42a6db37, 32'h4163d7db, 32'hc1e095b4, 32'hc20593d4, 32'hc1c313a4, 32'hbfdffd6d, 32'hc18bc224, 32'h408ad968};
test_weights[5824:5831] = '{32'h427b3aa6, 32'h4255565e, 32'h4271f979, 32'h423e8386, 32'h41ac20b4, 32'h4174729b, 32'hc21f98a0, 32'hc15aa664};
test_bias[728:728] = '{32'h4285ad56};
test_output[728:728] = '{32'h4532fccb};
test_input[5832:5839] = '{32'h421685aa, 32'hc2c7d427, 32'h42058c19, 32'h428a4184, 32'h41c7dd30, 32'hc269f075, 32'hc104e6b6, 32'hc17b9b46};
test_weights[5832:5839] = '{32'hc24b87c6, 32'hc29bf366, 32'hc2c33999, 32'hc1c54c96, 32'h41a6b22d, 32'hc23f06f3, 32'hc22d9951, 32'h419f94c7};
test_bias[729:729] = '{32'hc28f9c47};
test_output[729:729] = '{32'h45834749};
test_input[5840:5847] = '{32'h4222b533, 32'hc293dfc5, 32'h42a3de85, 32'h42c6ca77, 32'h419fe556, 32'h42aff184, 32'hc27de1c1, 32'hc2c1297d};
test_weights[5840:5847] = '{32'h422f22ac, 32'h420b9ee4, 32'h4217eaaa, 32'h428b91d1, 32'hc200dbe5, 32'h41fc4cc6, 32'h41643d21, 32'h429d03d0};
test_bias[730:730] = '{32'h4294e111};
test_output[730:730] = '{32'h453958bf};
test_input[5848:5855] = '{32'hc23ded86, 32'hc1822403, 32'hc2900056, 32'h42bb81ad, 32'h41ae710d, 32'h3fda3f57, 32'hc1a7def5, 32'h42b7e37e};
test_weights[5848:5855] = '{32'hc22d8664, 32'h42b39019, 32'h42926e99, 32'h4114d2b0, 32'h42bfa26d, 32'hc281e646, 32'hc2791bd0, 32'h422246f6};
test_bias[731:731] = '{32'hc2a14b01};
test_output[731:731] = '{32'h4543e986};
test_input[5856:5863] = '{32'h41e2cfd1, 32'hc1691c5a, 32'h42645c8a, 32'h425c1759, 32'h426b7854, 32'hc2a66ada, 32'hc1654edc, 32'h41413abc};
test_weights[5856:5863] = '{32'h41873408, 32'h409ee359, 32'h42923eaf, 32'h3f6173ed, 32'hc2ad1de7, 32'hc249772c, 32'hc1e15bf5, 32'h425b1560};
test_bias[732:732] = '{32'h42ab2556};
test_output[732:732] = '{32'h4598606e};
test_input[5864:5871] = '{32'hc0e106b2, 32'hc2b077e9, 32'h42b68713, 32'hc2bac8c7, 32'h4288212a, 32'hc150945e, 32'hc19546c4, 32'h426c46f0};
test_weights[5864:5871] = '{32'h41ebe232, 32'h41c2e7f7, 32'h410d949c, 32'hc2b43db7, 32'h4299b9e2, 32'hc1900580, 32'hc1da5a09, 32'h423ed499};
test_bias[733:733] = '{32'hc2645ac4};
test_output[733:733] = '{32'h4673cee0};
test_input[5872:5879] = '{32'h4296855a, 32'h428802e3, 32'h42aee6bc, 32'hc06d32ab, 32'hc167f7e1, 32'h42bbc331, 32'hc2400038, 32'h429a5b33};
test_weights[5872:5879] = '{32'hc21cb9e4, 32'hc20f15d3, 32'h429c1111, 32'hc2bf6db2, 32'h42980f2c, 32'h4293e130, 32'hc0a36cd0, 32'hc2c32ca8};
test_bias[734:734] = '{32'h428d2f94};
test_output[734:734] = '{32'h43d25fe2};
test_input[5880:5887] = '{32'h42252df8, 32'h42a2cee5, 32'hc27a8fff, 32'hc1f518d3, 32'h40b2948d, 32'h42ac675a, 32'h4284fae9, 32'h4260e852};
test_weights[5880:5887] = '{32'h423d5883, 32'h42118c01, 32'hc13333d6, 32'h429245f9, 32'h428b40e2, 32'h41000c1d, 32'hc2a1f605, 32'h413c2a5d};
test_bias[735:735] = '{32'h42467c90};
test_output[735:735] = '{32'hc3596e07};
test_input[5888:5895] = '{32'hc2a375c0, 32'h40419bb2, 32'hc2aeb540, 32'h42688d62, 32'hc2c67c8c, 32'h426c1ab2, 32'hc2c6eafe, 32'h4281e513};
test_weights[5888:5895] = '{32'h4284c954, 32'h4241f4d3, 32'hc2a85194, 32'hc2348f92, 32'h42b1b678, 32'h4176e026, 32'h42352bfb, 32'h4281db96};
test_bias[736:736] = '{32'h417c4163};
test_output[736:736] = '{32'hc608702c};
test_input[5896:5903] = '{32'hc243a1fe, 32'hc28aad99, 32'hc1f56649, 32'h421db90a, 32'hc2ad1357, 32'hc2a4d2c9, 32'h415fb80d, 32'h4245eaf9};
test_weights[5896:5903] = '{32'h4188f2b4, 32'h42aa2836, 32'h418d48ff, 32'hc25959d3, 32'h42b9bc3b, 32'h420c839d, 32'hc1ef091f, 32'h4239050c};
test_bias[737:737] = '{32'hc2c6842a};
test_output[737:737] = '{32'hc6912981};
test_input[5904:5911] = '{32'h427c44de, 32'hc2a2eae1, 32'h42700b1b, 32'hc1e09d2a, 32'h423d132f, 32'h4284534a, 32'hc2274b28, 32'h3fac5035};
test_weights[5904:5911] = '{32'hc2a9891e, 32'h418839d0, 32'hc284255e, 32'h42907902, 32'h3fddc9a1, 32'hc26a4d9f, 32'h42b60585, 32'h420fc8b3};
test_bias[738:738] = '{32'hc28a6ace};
test_output[738:738] = '{32'hc69ef682};
test_input[5912:5919] = '{32'h41ecba03, 32'h42b6155d, 32'hc279bb65, 32'h42bb93b2, 32'h4286fc04, 32'h41fd8c8d, 32'hc287294e, 32'hc2aea8bb};
test_weights[5912:5919] = '{32'h411a2215, 32'h42765be5, 32'h42c26c99, 32'hc0d48929, 32'h42abdd56, 32'hc2bf48c6, 32'h4281ea1c, 32'h40ef2c17};
test_bias[739:739] = '{32'hc1b2328d};
test_output[739:739] = '{32'hc5418321};
test_input[5920:5927] = '{32'hc217e483, 32'h42903143, 32'hc1efee5c, 32'h42a112d6, 32'h4185e4c5, 32'hc2ad3294, 32'h42a2d36a, 32'hc1d88133};
test_weights[5920:5927] = '{32'hc2c48564, 32'hc22886a4, 32'h421c0820, 32'h40f2b6f5, 32'hc23a9ec5, 32'h4245ae15, 32'hc2a811d4, 32'hc264d751};
test_bias[740:740] = '{32'h421bde92};
test_output[740:740] = '{32'hc61f1087};
test_input[5928:5935] = '{32'hc225f8ee, 32'hc19ca3a7, 32'hc21b5430, 32'h42784e18, 32'h41b08d39, 32'hc21e3739, 32'h4190996d, 32'h429f2ce4};
test_weights[5928:5935] = '{32'h423cee68, 32'hc1b1736e, 32'h428e3546, 32'h422fc46e, 32'h4254b4da, 32'hc2373999, 32'h408d87b2, 32'hc14f36a7};
test_bias[741:741] = '{32'h426eba6a};
test_output[741:741] = '{32'h4405d6c5};
test_input[5936:5943] = '{32'h42b914c3, 32'hc22f875a, 32'hc2c17967, 32'hc2b5272e, 32'h41d75559, 32'hc2ae2aac, 32'h428c18b8, 32'hc2815024};
test_weights[5936:5943] = '{32'h425ecad4, 32'hc2274f8a, 32'h4219c19f, 32'hc1cfc7d0, 32'h427a5b6e, 32'hc186862d, 32'hc1f8e165, 32'hc2646a42};
test_bias[742:742] = '{32'h3eebdc02};
test_output[742:742] = '{32'h4620b916};
test_input[5944:5951] = '{32'hc2066254, 32'h41970616, 32'h4243e13a, 32'hc190dae3, 32'h4297f8cb, 32'h4192a6f6, 32'hc2a5f5e2, 32'h42851d0c};
test_weights[5944:5951] = '{32'h42a29f35, 32'hc2c62247, 32'hc291035f, 32'hc2b5ea16, 32'hc29ebf06, 32'h42a0cba7, 32'hc15960ef, 32'h3f158165};
test_bias[743:743] = '{32'h4142863c};
test_output[743:743] = '{32'hc61a7275};
test_input[5952:5959] = '{32'h4244c3af, 32'hc2a9893f, 32'h4210183e, 32'h41dc86df, 32'h42b2dabe, 32'h425f763c, 32'hc063222a, 32'hc29d959e};
test_weights[5952:5959] = '{32'hc2821c39, 32'hc2c6e319, 32'h419a68af, 32'hc2406f89, 32'hc288f9a9, 32'h41bb17e9, 32'h424cd716, 32'hc2af37b0};
test_bias[744:744] = '{32'hc205ae8a};
test_output[744:744] = '{32'h45ca21b5};
test_input[5960:5967] = '{32'h4296b3fc, 32'h41c8743a, 32'h42a37c5d, 32'hbf4a0014, 32'hc1ce1de1, 32'hc2be8b1c, 32'h4188dafd, 32'hc2c007a7};
test_weights[5960:5967] = '{32'h404b2d67, 32'hc1a5cfd5, 32'h42b7b2a9, 32'hc1870991, 32'hc1881827, 32'hc2036419, 32'hc2a1e640, 32'h41f9d334};
test_bias[745:745] = '{32'h425f0667};
test_output[745:745] = '{32'h45ca8c5e};
test_input[5968:5975] = '{32'h42ad6468, 32'hc25bdd4c, 32'hc2af4b6b, 32'hc2299aff, 32'h420a9e39, 32'hc1ec7fc5, 32'hc2516067, 32'hc2c5b94b};
test_weights[5968:5975] = '{32'h42b5ae74, 32'h4258d4d4, 32'hc08e9991, 32'hc28b2641, 32'hc25fa0b7, 32'hc2b86ad6, 32'hc2a18ba4, 32'hc184b238};
test_bias[746:746] = '{32'h42a31979};
test_output[746:746] = '{32'h4669f9ac};
test_input[5976:5983] = '{32'hc2384626, 32'h42567721, 32'hc2150698, 32'h4201b5bc, 32'h4185a779, 32'hc2a1c0bb, 32'h40b0e243, 32'hc25ca198};
test_weights[5976:5983] = '{32'h428ebba3, 32'h3fec8a27, 32'h42b70b5d, 32'h4233c371, 32'h42c39dc3, 32'h41ef92e7, 32'h41a841ca, 32'hc2194e24};
test_bias[747:747] = '{32'h4267cc99};
test_output[747:747] = '{32'hc5638dc9};
test_input[5984:5991] = '{32'h42b75a35, 32'h42abc511, 32'hc209d236, 32'h426c873d, 32'h42103fe2, 32'h4283d2ad, 32'hc29559d6, 32'hc273a2e6};
test_weights[5984:5991] = '{32'h423acf97, 32'h41cef413, 32'h42bbefff, 32'hc2035a05, 32'hc24e93c1, 32'hc28bf75b, 32'h429cd68c, 32'hc2a80458};
test_bias[748:748] = '{32'hc13d5808};
test_output[748:748] = '{32'hc5b871de};
test_input[5992:5999] = '{32'h4266b833, 32'h41e9462c, 32'hc20c09e1, 32'h42053efe, 32'h42bdb7e9, 32'hc26c87a7, 32'hc00e0f5e, 32'hc2be2353};
test_weights[5992:5999] = '{32'hc29a8e53, 32'h42be3048, 32'h41b8100e, 32'h42471b43, 32'h421ea130, 32'hc2be271d, 32'h42c27938, 32'h41a81a61};
test_bias[749:749] = '{32'hc24f47c7};
test_output[749:749] = '{32'h45c47638};
test_input[6000:6007] = '{32'hc1d6b8ff, 32'h41ac1eb1, 32'hc292fc3f, 32'h42a5f275, 32'h423d624b, 32'h41962a14, 32'hc2037b9a, 32'h41ac7548};
test_weights[6000:6007] = '{32'h4087d95f, 32'hc1ad230c, 32'hc2a4fcc0, 32'h3f9b00c1, 32'h41d3fdd2, 32'hc2b535c9, 32'h42baeedc, 32'h41baeae0};
test_bias[750:750] = '{32'hc14e52e9};
test_output[750:750] = '{32'h451fbf77};
test_input[6008:6015] = '{32'h428a25f5, 32'h42aa9304, 32'h4268b18c, 32'h421a08d7, 32'hc2814116, 32'hc1deeed8, 32'hc1a78e49, 32'h422af833};
test_weights[6008:6015] = '{32'h3fabf493, 32'hc26cb905, 32'h4244ff13, 32'h42a74d23, 32'hc2878b3c, 32'hc2965e65, 32'h41174dff, 32'h3f5d188c};
test_bias[751:751] = '{32'hc21ad59a};
test_output[751:751] = '{32'h45e77716};
test_input[6016:6023] = '{32'hc1f69cac, 32'hc1d61c7c, 32'h42c75eb3, 32'h42b0df82, 32'hc21b5767, 32'h42aac098, 32'h424ae8f7, 32'h428d24fd};
test_weights[6016:6023] = '{32'h42c4bbdd, 32'h42046df9, 32'h422eb87d, 32'h4130d06f, 32'hc1028288, 32'h42ac6af8, 32'hc1b1f6fa, 32'h41c41804};
test_bias[752:752] = '{32'hc2b3bb8b};
test_output[752:752] = '{32'h46160696};
test_input[6024:6031] = '{32'h42962551, 32'h41297cef, 32'h429fe109, 32'h4222abe4, 32'hc204022d, 32'h428d9aa5, 32'h42742d6c, 32'h3ff76b0e};
test_weights[6024:6031] = '{32'h42b197ca, 32'h428f4232, 32'hc2969cc9, 32'hc2b05aa2, 32'hc2b0b9af, 32'hc1902deb, 32'h41bcecd7, 32'h425402cc};
test_bias[753:753] = '{32'hc1c23e37};
test_output[753:753] = '{32'h4474bdda};
test_input[6032:6039] = '{32'h42a006a2, 32'hc2766ade, 32'hc23e1e8f, 32'hc16bc6a9, 32'h412d1c2d, 32'hc254ded8, 32'hc2a0e084, 32'hc27799bb};
test_weights[6032:6039] = '{32'h426ecddf, 32'hc241137f, 32'h42141d8e, 32'hc15058ba, 32'hc0a3f6a1, 32'h42850e9d, 32'h429331a6, 32'h415659c4};
test_bias[754:754] = '{32'h424b1384};
test_output[754:754] = '{32'hc58080de};
test_input[6040:6047] = '{32'hbe0fbf25, 32'hc2b1d296, 32'h4276247c, 32'h427ae917, 32'hc2b0a5aa, 32'h4295ca1f, 32'h42409497, 32'hc2b8eafa};
test_weights[6040:6047] = '{32'hc2c3ff60, 32'h41c2311c, 32'hc26e7cc7, 32'h4204ff4f, 32'h429cd690, 32'hc20e5fc8, 32'hc23f8368, 32'h419a518c};
test_bias[755:755] = '{32'h409399ff};
test_output[755:755] = '{32'hc687f772};
test_input[6048:6055] = '{32'hc2876d38, 32'hc2aab844, 32'h42960ab0, 32'h41801e97, 32'h419f7cce, 32'hc12f5742, 32'hc2ae6b25, 32'hc26ba2a8};
test_weights[6048:6055] = '{32'hbfbf02bc, 32'h429f7fc1, 32'hc1217c1e, 32'hc2229378, 32'h401a9506, 32'h42331d37, 32'h42a21c1e, 32'hc203de0d};
test_bias[756:756] = '{32'h40fb0425};
test_output[756:756] = '{32'hc655af7b};
test_input[6056:6063] = '{32'h4296868e, 32'hc25994d4, 32'hc2a12f2f, 32'h41be9171, 32'hc277eb70, 32'hc2178a9c, 32'h41d975b1, 32'hc22bbaeb};
test_weights[6056:6063] = '{32'hc1c85640, 32'h428a923b, 32'hc2aa58bb, 32'hc25044c5, 32'hc2bddc99, 32'hc289c3b1, 32'hc28f8307, 32'hc2858706};
test_bias[757:757] = '{32'hc2852186};
test_output[757:757] = '{32'h461184a0};
test_input[6064:6071] = '{32'hc28f66d3, 32'hc2a716f2, 32'hc2645a35, 32'hc2b64a54, 32'h421c23c2, 32'h429b5698, 32'hc27345aa, 32'hc2a207c1};
test_weights[6064:6071] = '{32'hc1f2a1c3, 32'hc24b65e8, 32'hc0e4001f, 32'h42c6ecd5, 32'hc286617e, 32'hc20dbb19, 32'h423b0044, 32'h423f109a};
test_bias[758:758] = '{32'h41777250};
test_output[758:758] = '{32'hc65f9155};
test_input[6072:6079] = '{32'hc2a234cd, 32'h42825b2e, 32'hc25cccd2, 32'hc2949e30, 32'hc29d262f, 32'hc261024c, 32'hc21e785d, 32'h429e950a};
test_weights[6072:6079] = '{32'h425bfe6d, 32'h41960b23, 32'hc21f05f1, 32'hc2b3545e, 32'hc209646e, 32'hc2711844, 32'h42419725, 32'hc2b27845};
test_bias[759:759] = '{32'h42b597ad};
test_output[759:759] = '{32'h452f6997};
test_input[6080:6087] = '{32'hc26f9e74, 32'hc1833831, 32'h42836b3e, 32'hc2865501, 32'h424c4216, 32'hc2876ce2, 32'h42394e62, 32'h41e242c4};
test_weights[6080:6087] = '{32'h4202819a, 32'h4170b6e4, 32'hc11e28e6, 32'hc107fa19, 32'hc262cdff, 32'h401756a6, 32'hc21f89ac, 32'h41ae4733};
test_bias[760:760] = '{32'h42597834};
test_output[760:760] = '{32'hc5cb85cd};
test_input[6088:6095] = '{32'hc20147ba, 32'h419ba9fd, 32'hc2a5000d, 32'hc2a1b297, 32'h41da254f, 32'h41b766d8, 32'h41a3e2e5, 32'hc2845eca};
test_weights[6088:6095] = '{32'h42c0c923, 32'hc288208a, 32'hc2afc903, 32'hc201415c, 32'hc1829614, 32'h41ef4725, 32'h4253e35b, 32'hc2894aae};
test_bias[761:761] = '{32'hc2b03c24};
test_output[761:761] = '{32'h462f136a};
test_input[6096:6103] = '{32'hc2b15a42, 32'hc2947f16, 32'h4255c691, 32'h3f0e7925, 32'h42250769, 32'h421cbe89, 32'hc23b6ac2, 32'hc20dd6ca};
test_weights[6096:6103] = '{32'hc22ab875, 32'hc1cb06c4, 32'hc2a96bdb, 32'h428a1a4c, 32'hc276e83a, 32'h41055399, 32'h429cf3eb, 32'hc200c62a};
test_bias[762:762] = '{32'h42c4b49d};
test_output[762:762] = '{32'hc5594ff9};
test_input[6104:6111] = '{32'h4234814d, 32'h429d4633, 32'h41d7149f, 32'hc25c6a6d, 32'hc22f4622, 32'hc15344fa, 32'h42a705bd, 32'hc29eada3};
test_weights[6104:6111] = '{32'hbfccaad7, 32'h4117e8ee, 32'hc2c6c56d, 32'hc1d4aa1e, 32'h426cc7ce, 32'hc1db05be, 32'hc1dbd296, 32'h40f435e0};
test_bias[763:763] = '{32'h41db9caf};
test_output[763:763] = '{32'hc5b02e34};
test_input[6112:6119] = '{32'hc1b09c48, 32'hc295410d, 32'hc11ab5a5, 32'hc2a710c0, 32'h41455208, 32'h42534967, 32'h3f63fdd0, 32'hc140edca};
test_weights[6112:6119] = '{32'hc2a69fbd, 32'h42c03464, 32'hc0fc0213, 32'h42a80b5c, 32'h42b6c98d, 32'hc283feb9, 32'hc2b68cc2, 32'h42548525};
test_bias[764:764] = '{32'h42c1136c};
test_output[764:764] = '{32'hc66e6dc8};
test_input[6120:6127] = '{32'h42ad4036, 32'hc21af178, 32'h417cf79f, 32'h42926ba3, 32'hc213737c, 32'hc12f7c9f, 32'hc23185b7, 32'hc25292b9};
test_weights[6120:6127] = '{32'h42499624, 32'h428a7137, 32'hc2444479, 32'hc1fdac41, 32'h41972e71, 32'hc0a81163, 32'h42297739, 32'hc284f6f4};
test_bias[765:765] = '{32'h41d6b245};
test_output[765:765] = '{32'hc3cabe31};
test_input[6128:6135] = '{32'hc298920d, 32'hc2624dbb, 32'hc29cbe56, 32'h428155be, 32'h429e634f, 32'hc18c9d41, 32'h4180cf8d, 32'h42af2e37};
test_weights[6128:6135] = '{32'hc2b3a8d8, 32'h41e86006, 32'hc229dd3d, 32'hc238f666, 32'hbbe9e291, 32'h4284d43d, 32'h41f794a6, 32'h428de27a};
test_bias[766:766] = '{32'h429a1402};
test_output[766:766] = '{32'h462e81ef};
test_input[6136:6143] = '{32'h420afc50, 32'hc2099c02, 32'hc29bb05f, 32'h41b2f774, 32'hc12b468f, 32'h42b9d04f, 32'hc238320e, 32'h4228582a};
test_weights[6136:6143] = '{32'h42b83c27, 32'hc2b1c998, 32'hc1474904, 32'hc1721b2d, 32'hc2aec657, 32'h42a79de1, 32'h3e653bd9, 32'h42c3f8ef};
test_bias[767:767] = '{32'hc2467210};
test_output[767:767] = '{32'h4699b77c};
test_input[6144:6151] = '{32'hc1aab0b0, 32'h409b17d9, 32'h4093a660, 32'hc2b8e389, 32'h4199ac1e, 32'h42a51e3e, 32'h428fc7ca, 32'hc2651767};
test_weights[6144:6151] = '{32'hc1e528f9, 32'h421fa532, 32'hc254f751, 32'h42abb7c5, 32'hc16109ab, 32'hc07ee8fd, 32'hc2be6ae9, 32'hc248951d};
test_bias[768:768] = '{32'hc07477b7};
test_output[768:768] = '{32'hc63ac693};
test_input[6152:6159] = '{32'h413c6490, 32'hc1f561aa, 32'h42b56128, 32'h41fd6050, 32'hc29c7aba, 32'hc107d247, 32'h42a5398c, 32'hc28a3480};
test_weights[6152:6159] = '{32'h40124c5b, 32'hc2bbf7b5, 32'h41f649e6, 32'h42114adb, 32'h42bd1d95, 32'h3f36988e, 32'h423cde91, 32'hc249eb7f};
test_bias[769:769] = '{32'h42bf5b7c};
test_output[769:769] = '{32'h45d8a45b};
test_input[6160:6167] = '{32'h42297010, 32'h3f0efa08, 32'h42a0b744, 32'hc214cb80, 32'hc24f2670, 32'hc0985ca5, 32'hc2471418, 32'hc2972615};
test_weights[6160:6167] = '{32'hc104b6ca, 32'hc2956ece, 32'h42956ccd, 32'hc2c43449, 32'hc03c2c01, 32'h4198d6bf, 32'h42a35004, 32'h41f631b4};
test_bias[770:770] = '{32'h42c12560};
test_output[770:770] = '{32'h453d40eb};
test_input[6168:6175] = '{32'hc1872ced, 32'h42593a5f, 32'hc2bc5159, 32'hc2b9f8f8, 32'hc1760963, 32'hc1e17191, 32'h42779216, 32'hc25afcf6};
test_weights[6168:6175] = '{32'hc25c2abd, 32'hc1a1b677, 32'h418bcd32, 32'hc2b6006e, 32'hc2a389a1, 32'hc0b9e13c, 32'h42981c08, 32'hc28ff4f3};
test_bias[771:771] = '{32'hc2648c23};
test_output[771:771] = '{32'h468228db};
test_input[6176:6183] = '{32'h40a85fc4, 32'hc241f4ea, 32'hbf29edb9, 32'h42231d52, 32'h40d9c57c, 32'h429b7af6, 32'h423b7f88, 32'h428802c8};
test_weights[6176:6183] = '{32'hc1d93eef, 32'h42983777, 32'h42ba045d, 32'h42027b79, 32'h428cb677, 32'h42bdae1c, 32'hc2b934f9, 32'h4272fafb};
test_bias[772:772] = '{32'h428472d4};
test_output[772:772] = '{32'h45a0ba9e};
test_input[6184:6191] = '{32'h410dd99a, 32'h4298eee9, 32'h42b39796, 32'hc2aa592b, 32'h41d5b103, 32'h42a769d5, 32'hc1ece599, 32'hc279ad4a};
test_weights[6184:6191] = '{32'h426e822b, 32'hc2794f01, 32'h42912202, 32'hc27ebabc, 32'h40420747, 32'hc2053d04, 32'hc1d66b9a, 32'hc235eb44};
test_bias[773:773] = '{32'hc195b50d};
test_output[773:773] = '{32'h460685ea};
test_input[6192:6199] = '{32'hc1e66af0, 32'hc20fe0ed, 32'h4250a3c0, 32'h42c5188c, 32'hc139150e, 32'hc2982e8e, 32'h3fcf5e13, 32'h4293a3c2};
test_weights[6192:6199] = '{32'h42c0ed50, 32'hc075e480, 32'h40b304e6, 32'hc206be00, 32'hc2a6c7f8, 32'hc297b523, 32'hc229c48d, 32'hc2af6b18};
test_bias[774:774] = '{32'hc16120df};
test_output[774:774] = '{32'hc5ab88c1};
test_input[6200:6207] = '{32'hc189a2f4, 32'h426e8141, 32'h426e414a, 32'h42231383, 32'hc2bba1fb, 32'h4297fe3a, 32'h4251deb0, 32'hc1077a19};
test_weights[6200:6207] = '{32'hc255ab77, 32'hc26bd1ef, 32'hc1eba9fc, 32'hc0d24c73, 32'h425b1eb7, 32'h4129a8b8, 32'h417e75ee, 32'h3f138285};
test_bias[775:775] = '{32'hc2082b5a};
test_output[775:775] = '{32'hc5fee5a1};
test_input[6208:6215] = '{32'hc0bcc465, 32'hc2be1c86, 32'h4270cd43, 32'h41dda647, 32'h429fb0d4, 32'hc1f17342, 32'h42bd2d96, 32'hc2bb2621};
test_weights[6208:6215] = '{32'h412a0754, 32'hc1562bce, 32'hc2c4bd8a, 32'h426be8d3, 32'hc0e1499b, 32'hc04abd01, 32'hc20561d9, 32'hc2b781d3};
test_bias[776:776] = '{32'hc1f61db0};
test_output[776:776] = '{32'h44e80604};
test_input[6216:6223] = '{32'h42a29448, 32'h421a40c1, 32'h418bee87, 32'hc1288981, 32'hc2b68486, 32'hc2254cbd, 32'hc29bf859, 32'hc28514fa};
test_weights[6216:6223] = '{32'h42aedf7b, 32'h4226e508, 32'hc2a2015e, 32'h425c3098, 32'h41c3504f, 32'hc18170ec, 32'h426bfc64, 32'h429d02d2};
test_bias[777:777] = '{32'hc0efa387};
test_output[777:777] = '{32'hc591fc79};
test_input[6224:6231] = '{32'hc2c6489f, 32'hc290a248, 32'h429922ec, 32'hc1bb7cf0, 32'hc2bd0ad9, 32'h42b34739, 32'h41bbb898, 32'hc1863c02};
test_weights[6224:6231] = '{32'h428a5367, 32'hc235d597, 32'hc0ae08cf, 32'h410da9b4, 32'h4299e5c9, 32'hc2bef5c3, 32'h4290b3ef, 32'hc1939ff9};
test_bias[778:778] = '{32'h42a2132a};
test_output[778:778] = '{32'hc68c2221};
test_input[6232:6239] = '{32'hc2b417c8, 32'h410e61b3, 32'hc2b59603, 32'h40c8e7c1, 32'hc269cef5, 32'hc2c64b9d, 32'h413fc547, 32'h4292ffe7};
test_weights[6232:6239] = '{32'hc2880fe2, 32'hc288b648, 32'h42a45390, 32'hc197adc2, 32'hc2870f99, 32'h429eae68, 32'h42b1f639, 32'hc238918e};
test_bias[779:779] = '{32'h4266ed01};
test_output[779:779] = '{32'hc600de4a};
test_input[6240:6247] = '{32'hc2bcc9b0, 32'h422d3d5b, 32'h420dd30c, 32'hc2a9911f, 32'h42065e2f, 32'hc21b4c09, 32'hc2685cd4, 32'hc2ba667c};
test_weights[6240:6247] = '{32'hc2047b2f, 32'h40e48218, 32'hc284a7cb, 32'h410b6c2e, 32'hc24606b7, 32'hc2a3a3f3, 32'h42c25a91, 32'h4197acdc};
test_bias[780:780] = '{32'h421939af};
test_output[780:780] = '{32'hc5ac58b5};
test_input[6248:6255] = '{32'hc273ae31, 32'h42926a8c, 32'hc1ce6b7d, 32'hc26fd110, 32'hc2b07ea6, 32'hc0fea51f, 32'h424ecaa8, 32'h42ba0cd0};
test_weights[6248:6255] = '{32'h42876043, 32'hc2ae3ee2, 32'hc263310c, 32'hc20c2def, 32'h427679ec, 32'h42919f76, 32'hc2af2c65, 32'hc070fefc};
test_bias[781:781] = '{32'hc2ac0e78};
test_output[781:781] = '{32'hc68bf916};
test_input[6256:6263] = '{32'hc29359b0, 32'hc2b684db, 32'h41c530ad, 32'h42868209, 32'h41aa5ef4, 32'hc253efbf, 32'h40825612, 32'h4269d6a2};
test_weights[6256:6263] = '{32'h4200afa9, 32'hc24ea78d, 32'hc281f356, 32'hc1db7d09, 32'hc25d4b9d, 32'hc20dc8d1, 32'h4276b109, 32'hc1e47904};
test_bias[782:782] = '{32'hc19b5422};
test_output[782:782] = '{32'hc4e602a3};
test_input[6264:6271] = '{32'hc2b88442, 32'hc210a845, 32'h42328b31, 32'h4188dca8, 32'hc2a1f8d1, 32'h42924a6e, 32'h41dc936c, 32'h421369d3};
test_weights[6264:6271] = '{32'h42178736, 32'hc265bdc9, 32'h42c47f83, 32'h423b4128, 32'h4204aa16, 32'h419baa67, 32'hc1df4348, 32'h4243702c};
test_bias[783:783] = '{32'h424fae8f};
test_output[783:783] = '{32'h45604dca};
test_input[6272:6279] = '{32'h425d7ddc, 32'h420158c8, 32'hc1932678, 32'h41fe128e, 32'h42389041, 32'h42a50e5d, 32'hc29c6635, 32'h42881168};
test_weights[6272:6279] = '{32'hc246d8d0, 32'hc03de166, 32'h42970bdf, 32'h41c492b3, 32'h42547d10, 32'hc234927a, 32'h42a4db98, 32'h42bfd945};
test_bias[784:784] = '{32'h42af7d60};
test_output[784:784] = '{32'hc58e9f5c};
test_input[6280:6287] = '{32'hc2b5af32, 32'h426e89d2, 32'hc1c4efea, 32'hc1d71b12, 32'hc285385c, 32'hc1d857fb, 32'hc189a536, 32'h4297bea6};
test_weights[6280:6287] = '{32'h42bd6544, 32'h41e32ce9, 32'hc1b98a36, 32'h41146db6, 32'h429fbe0f, 32'h4223c550, 32'h40dc2bc5, 32'hc2291348};
test_bias[785:785] = '{32'h4213d61e};
test_output[785:785] = '{32'hc67ebe0e};
test_input[6288:6295] = '{32'h41b152c9, 32'hc0eee701, 32'hc24b56e4, 32'h42b563bf, 32'h41caf6dc, 32'hc2500fb7, 32'h42aceac4, 32'hc213955a};
test_weights[6288:6295] = '{32'hc28f165e, 32'h42a836b4, 32'hc20e6b5c, 32'hc184a0c5, 32'h42400951, 32'h427aeb0b, 32'hc2093d40, 32'hc1c55587};
test_bias[786:786] = '{32'h42c67e6e};
test_output[786:786] = '{32'hc5b8a9ea};
test_input[6296:6303] = '{32'hc266c647, 32'h3ff26e53, 32'h412970dd, 32'hc2bde467, 32'h3f379b38, 32'h424d4d9c, 32'h4288f021, 32'hc15a1405};
test_weights[6296:6303] = '{32'h42aaf87d, 32'h411fb9bf, 32'hc2b79c98, 32'hc23644cc, 32'h41f1ac80, 32'h42c6d3a8, 32'hc17e0b91, 32'hc0b7346c};
test_bias[787:787] = '{32'h42986f16};
test_output[787:787] = '{32'h4524864e};
test_input[6304:6311] = '{32'h421766fc, 32'h421559f6, 32'h424b8101, 32'h41f4ca00, 32'hc2800fcd, 32'h422847dc, 32'h4236d64b, 32'h42986f58};
test_weights[6304:6311] = '{32'hc2a467b6, 32'h41a4ba1d, 32'hc1851b20, 32'hc2a6ed1c, 32'h42487bc5, 32'hc228901c, 32'hc1df8426, 32'h42b930da};
test_bias[788:788] = '{32'h429de14b};
test_output[788:788] = '{32'hc5980edb};
test_input[6312:6319] = '{32'hc27f5195, 32'hc2c64128, 32'hc293462d, 32'h42210b14, 32'h4216ca7d, 32'hc12e88be, 32'h428ce5cd, 32'h4266b63a};
test_weights[6312:6319] = '{32'hc1f351be, 32'h42311c1b, 32'hc265bbf9, 32'hc2b84f17, 32'hc20834ac, 32'h424b7abc, 32'hc29ebd04, 32'hc0d782e3};
test_bias[789:789] = '{32'h42af1cc2};
test_output[789:789] = '{32'hc616ee84};
test_input[6320:6327] = '{32'h42be0609, 32'h42b4c340, 32'hc2723865, 32'h425ab1bb, 32'hc2218cf8, 32'h404a3ee5, 32'hc2b148b0, 32'h4203f4f3};
test_weights[6320:6327] = '{32'hc117389a, 32'hc22484ac, 32'h429c6fc1, 32'h4231837f, 32'hc22bf34e, 32'h42ac7012, 32'hc2a398cc, 32'h421e4878};
test_bias[790:790] = '{32'hc12a8569};
test_output[790:790] = '{32'h4562ca28};
test_input[6328:6335] = '{32'hc2a01546, 32'hc1921c14, 32'h423f05df, 32'hc2c71972, 32'hc17f4978, 32'h423fd8eb, 32'hc220b8dd, 32'hc1980bea};
test_weights[6328:6335] = '{32'hc23a8d0e, 32'hc1a6ff79, 32'h42c46b0c, 32'h42064386, 32'h42ae08a5, 32'h42435a49, 32'h42c237ce, 32'h42584b50};
test_bias[791:791] = '{32'hc20629ba};
test_output[791:791] = '{32'h44b5b36f};
test_input[6336:6343] = '{32'h41cacc26, 32'h42617223, 32'hc2487de2, 32'hc18f51b7, 32'h428c915e, 32'hc2488b24, 32'h42a90637, 32'h42b1baf8};
test_weights[6336:6343] = '{32'hc205c266, 32'hc2bbef2d, 32'hc2b193eb, 32'h419a876e, 32'h429f02de, 32'hc2c201a5, 32'h423b9795, 32'h40eb681a};
test_bias[792:792] = '{32'hc1b822fb};
test_output[792:792] = '{32'h464b37e6};
test_input[6344:6351] = '{32'hc26f30f4, 32'h41931533, 32'hc284ffb6, 32'h41bf7847, 32'hc1b85ffd, 32'hc229c5bf, 32'h4212bd5a, 32'hc10b7408};
test_weights[6344:6351] = '{32'h42c5007c, 32'h42689424, 32'hc299c774, 32'h42808d4b, 32'hc20df007, 32'h41df7150, 32'hc0d8e4fe, 32'hc243fab9};
test_bias[793:793] = '{32'h41dee029};
test_output[793:793] = '{32'h44d09e21};
test_input[6352:6359] = '{32'hc123ec0e, 32'hc25899a3, 32'h42b25be7, 32'h426ada0e, 32'h42b8e7be, 32'h42ad54c4, 32'hc1aae609, 32'h420d784e};
test_weights[6352:6359] = '{32'hc2991eaa, 32'h4082d50d, 32'h42ad5d44, 32'hc24158ea, 32'h4234aacf, 32'hc29be0f7, 32'h4186b22c, 32'hc21c433a};
test_bias[794:794] = '{32'hc0dad6b4};
test_output[794:794] = '{32'h448d069a};
test_input[6360:6367] = '{32'hc14fc02c, 32'hc24e0387, 32'h424dece5, 32'hc1c669c1, 32'h3fcb32d4, 32'hc1b15b71, 32'h429ce017, 32'hc1430e52};
test_weights[6360:6367] = '{32'h429ece97, 32'h4286f689, 32'h42c7d24d, 32'hc1dc2b48, 32'h41c75d87, 32'hc23f0768, 32'h4251d75b, 32'hc2069325};
test_bias[795:795] = '{32'hc255eb78};
test_output[795:795] = '{32'h45d74b6b};
test_input[6368:6375] = '{32'hc2244a82, 32'hc280296b, 32'h42963669, 32'hc2917fb8, 32'hc1ec36ad, 32'h418bfb60, 32'h4133bda1, 32'hc29baf67};
test_weights[6368:6375] = '{32'h428fe682, 32'h428925b5, 32'hc242a8a1, 32'hc22e55ee, 32'h418df18e, 32'h4206dcc1, 32'h41d9889d, 32'h42c74622};
test_bias[796:796] = '{32'h40f5f2db};
test_output[796:796] = '{32'hc66daa41};
test_input[6376:6383] = '{32'h42ad9f16, 32'h418e1664, 32'hc1b46aa1, 32'hc1ce08c8, 32'h428dfbdc, 32'hc29fa9ed, 32'h4210aa95, 32'h42ad5428};
test_weights[6376:6383] = '{32'hc1bdbe80, 32'hc1940f4e, 32'h42bf459d, 32'h426b468e, 32'hc22dd104, 32'h41a11053, 32'hc2398d97, 32'hc2be20a5};
test_bias[797:797] = '{32'hc2a6f043};
test_output[797:797] = '{32'hc6a21e8d};
test_input[6384:6391] = '{32'h42a622a6, 32'hc1c27d2e, 32'h41aee82d, 32'h42c53c73, 32'hc2ac1960, 32'h4213d8df, 32'hc1ddb10a, 32'h426f2bfe};
test_weights[6384:6391] = '{32'hc2ba7afd, 32'hc2856121, 32'h40efaf93, 32'h428a7a76, 32'h41acc0df, 32'hc25220aa, 32'h41924a8e, 32'h42353070};
test_bias[798:798] = '{32'hc259bc62};
test_output[798:798] = '{32'hc44420a6};
test_input[6392:6399] = '{32'h41e7908d, 32'h41f46167, 32'h426cadaa, 32'h412f9d12, 32'h42a7a69c, 32'hc22f95be, 32'h41312dfc, 32'hc2028e5d};
test_weights[6392:6399] = '{32'hbf18f6e1, 32'hc270a33c, 32'hc2adcbb2, 32'h428bc47f, 32'hc2999797, 32'h42c42349, 32'h41e32c73, 32'hc2bbb7de};
test_bias[799:799] = '{32'h42845aa6};
test_output[799:799] = '{32'hc6535fa3};
test_input[6400:6407] = '{32'hc205f207, 32'h4285db45, 32'hc2116736, 32'hc11ac5c1, 32'hc295b89e, 32'hc27bd077, 32'h4251ee76, 32'h4297ff8b};
test_weights[6400:6407] = '{32'h41df3d51, 32'h4291cc5e, 32'h42b68652, 32'h4278b79a, 32'h41e25d5a, 32'h428ba41b, 32'hc2abc2f9, 32'h3f5ffe4a};
test_bias[800:800] = '{32'hc2a90c4a};
test_output[800:800] = '{32'hc62c1553};
test_input[6408:6415] = '{32'h427e519c, 32'h422eff79, 32'h42c214e0, 32'h41551194, 32'h42282962, 32'h42bbe426, 32'hc2083349, 32'h411a3512};
test_weights[6408:6415] = '{32'hc2a0e1a1, 32'h42ac7018, 32'h416f263a, 32'hc1df7048, 32'hc2761a59, 32'hc11a8187, 32'h42308f77, 32'hc297d7fe};
test_bias[801:801] = '{32'h42ac7f6d};
test_output[801:801] = '{32'hc5b89085};
test_input[6416:6423] = '{32'h421262d6, 32'h42b52ccf, 32'hc2adb147, 32'h41075967, 32'hc2bd08b0, 32'hc29f2f24, 32'h42a83604, 32'hc2400d69};
test_weights[6416:6423] = '{32'h4288879c, 32'hc130fd23, 32'h40c1ac0b, 32'h42a1f7ae, 32'hc2138c9f, 32'hc19dbcd9, 32'h42bc0a04, 32'hc222a8bf};
test_bias[802:802] = '{32'hc299faf1};
test_output[802:802] = '{32'h4680dcf3};
test_input[6424:6431] = '{32'h41ea1c57, 32'h409bbf35, 32'hc1544330, 32'hc2a4cfa4, 32'hc2144402, 32'h4287d912, 32'h42448e0c, 32'h4231bdd8};
test_weights[6424:6431] = '{32'hc225cd7b, 32'hc10e8771, 32'h4267e090, 32'hc21697de, 32'h41023c8e, 32'hc240cb83, 32'hc25b3e22, 32'h40d2ab89};
test_bias[803:803] = '{32'hc2926801};
test_output[803:803] = '{32'hc59b643e};
test_input[6432:6439] = '{32'hc2b71c9b, 32'h424ef7cd, 32'hc1d4588d, 32'h41dbd101, 32'h415dafc7, 32'hc290aeed, 32'hc25010b0, 32'h41a42446};
test_weights[6432:6439] = '{32'hc25c4df3, 32'h40129c38, 32'h41c9d55c, 32'hc267ff97, 32'h41b11e5c, 32'hc1353eee, 32'h42a4cb6e, 32'hc2964431};
test_bias[804:804] = '{32'h42927e67};
test_output[804:804] = '{32'hc4d84ab6};
test_input[6440:6447] = '{32'hc2a22072, 32'hc2a8242f, 32'hc0cb4ba5, 32'h41bf2f84, 32'hc277f54d, 32'h41883f18, 32'hc2a565f5, 32'hc2802ffe};
test_weights[6440:6447] = '{32'hc200dcd7, 32'h422dc0bb, 32'h41f5f70c, 32'hc142ce12, 32'h42669bc7, 32'h4294a0df, 32'hc219210a, 32'h42aa8b4f};
test_bias[805:805] = '{32'hc1328e03};
test_output[805:805] = '{32'hc5c00c27};
test_input[6448:6455] = '{32'h41249d7b, 32'h42afe4bd, 32'h42b890e2, 32'hc260378c, 32'hc289e11d, 32'h4280dc31, 32'hc2651b43, 32'hc2038583};
test_weights[6448:6455] = '{32'hc24a0b9a, 32'h425c5b99, 32'hc2369bdd, 32'hc1395d5d, 32'hc150197b, 32'hc29ecc2a, 32'h4282e2e5, 32'h42402b59};
test_bias[806:806] = '{32'h427bd016};
test_output[806:806] = '{32'hc6084960};
test_input[6456:6463] = '{32'hc28edf62, 32'h426195ce, 32'hc2c426ae, 32'hc129e305, 32'hc1efe062, 32'hc1829deb, 32'hc1bd1d8f, 32'hc2992126};
test_weights[6456:6463] = '{32'hc20dcd01, 32'h41c9f2bc, 32'hc2033135, 32'h422d14e1, 32'h42025c24, 32'hc2ab5871, 32'h42b17f74, 32'hc21068b7};
test_bias[807:807] = '{32'h42503d22};
test_output[807:807] = '{32'h45f5693d};
test_input[6464:6471] = '{32'hc19010ff, 32'hc2191906, 32'h41637494, 32'h409e509f, 32'hc1334308, 32'hc25e3a20, 32'hc2508963, 32'h421e7be1};
test_weights[6464:6471] = '{32'h42846243, 32'h4165347f, 32'hc2762d82, 32'hc2c190dd, 32'h423d09b0, 32'hc203a9e4, 32'hc1e0d876, 32'hc29e15dc};
test_bias[808:808] = '{32'hbea4b457};
test_output[808:808] = '{32'hc55859eb};
test_input[6472:6479] = '{32'h42b29b69, 32'h4291f743, 32'hc287b8c0, 32'h42bcaeaa, 32'h42922a1a, 32'hc20edda2, 32'h42a0d810, 32'h428759a8};
test_weights[6472:6479] = '{32'hc2bdcd58, 32'hc170c46e, 32'hc031f04c, 32'hc08e2ce3, 32'hc2870c40, 32'h42b1d883, 32'hc2886c6f, 32'h4216be19};
test_bias[809:809] = '{32'h3fe3fe8a};
test_output[809:809] = '{32'hc6a2e034};
test_input[6480:6487] = '{32'hc2593f76, 32'hc297f478, 32'hc25e9c92, 32'hc2ab1d15, 32'hbfeaa0ef, 32'hc2a57040, 32'hc26fab60, 32'h42a356ce};
test_weights[6480:6487] = '{32'h4193238a, 32'hc28b587d, 32'hc2a5526b, 32'hc17449bd, 32'hc11fd460, 32'hc2ba83ab, 32'h42282e8e, 32'hc2a166ff};
test_bias[810:810] = '{32'hc1ef8f47};
test_output[810:810] = '{32'h460966c5};
test_input[6488:6495] = '{32'h42b797e6, 32'hc28b1bb8, 32'hc2b79923, 32'h421f7613, 32'hc2c29a5c, 32'hc2819474, 32'h41129ff7, 32'h426dccad};
test_weights[6488:6495] = '{32'h421ac388, 32'hc2a7561d, 32'h42659068, 32'h42253e21, 32'hc215bfea, 32'hc1d82e7c, 32'h410e02fc, 32'h42266029};
test_bias[811:811] = '{32'h41efd078};
test_output[811:811] = '{32'h46567caf};
test_input[6496:6503] = '{32'hc273eb68, 32'hc2980845, 32'h42a50349, 32'h42971e4c, 32'hc2b44eb1, 32'hc149269b, 32'hc28db672, 32'h428940ef};
test_weights[6496:6503] = '{32'h42c4cf04, 32'h42b47133, 32'h425aab81, 32'hc190e20e, 32'hc1943142, 32'h42ab91cd, 32'h429fb690, 32'hc0f0340f};
test_bias[812:812] = '{32'hc28e8314};
test_output[812:812] = '{32'hc670288d};
test_input[6504:6511] = '{32'hc2560fa4, 32'hc1c923b8, 32'hc1c03263, 32'hc1bc3358, 32'hc12fb6c1, 32'h4184a62f, 32'h42b6cd60, 32'hc28f6938};
test_weights[6504:6511] = '{32'hc2c54eee, 32'h429c9ff6, 32'hc28508b0, 32'hc2a940f9, 32'h412959e3, 32'h420e0e78, 32'h423f56bd, 32'h410ff5a4};
test_bias[813:813] = '{32'h4284c8ce};
test_output[813:813] = '{32'h462e75b9};
test_input[6512:6519] = '{32'hc1dbeb22, 32'hc25c67ad, 32'hc298155e, 32'h41eda1d0, 32'hc1391470, 32'hc2126cfa, 32'h42b0d01c, 32'hc1351252};
test_weights[6512:6519] = '{32'hc192547e, 32'hc25abd24, 32'h4288a6fb, 32'hc0989712, 32'hc2a11916, 32'hc2932105, 32'h41dfc307, 32'h42a9d8b1};
test_bias[814:814] = '{32'hc0a2583c};
test_output[814:814] = '{32'h454ee060};
test_input[6520:6527] = '{32'hc25b9958, 32'hc0bcd682, 32'hc27b46b6, 32'hc29ee121, 32'h41eb91a1, 32'hc2a2eeaa, 32'h420737ea, 32'hc2202583};
test_weights[6520:6527] = '{32'hc1e3d3ba, 32'h42aedf6f, 32'h419bc669, 32'h41041610, 32'hc2c1389c, 32'h4198dce0, 32'hc239c24c, 32'h421873e6};
test_bias[815:815] = '{32'h42a7da37};
test_output[815:815] = '{32'hc600d36c};
test_input[6528:6535] = '{32'h42b47877, 32'hc2850323, 32'h42b9dd0a, 32'hc295e6bc, 32'h40820805, 32'h428f70ba, 32'h4262c6c1, 32'h426b22a1};
test_weights[6528:6535] = '{32'hc29de2f7, 32'h420f3be6, 32'h4194c270, 32'hc14208d2, 32'hc2c2e862, 32'h423b64d2, 32'h426afe18, 32'hbff27729};
test_bias[816:816] = '{32'hc25ccdb7};
test_output[816:816] = '{32'hc438f6ff};
test_input[6536:6543] = '{32'hc2958464, 32'hc27f614b, 32'hc2ac2b6a, 32'h42282613, 32'hc2a40f2c, 32'h4216f779, 32'h427257bb, 32'hc291ed9a};
test_weights[6536:6543] = '{32'h420b4bbc, 32'hc29ffabf, 32'hc252ff84, 32'h428b2656, 32'h4217213e, 32'hc25bd226, 32'hc13fecb2, 32'hc2a68ea0};
test_bias[817:817] = '{32'hc2bb97f2};
test_output[817:817] = '{32'h461d0e90};
test_input[6544:6551] = '{32'h4297d850, 32'hc2630008, 32'h427a9378, 32'h42bf85d0, 32'h420fd41f, 32'h42a730b7, 32'h42693029, 32'h418ca787};
test_weights[6544:6551] = '{32'hbeb56400, 32'hc18246dd, 32'hc124f62c, 32'h41e0d0ba, 32'h41ba8506, 32'hc2b8ff09, 32'hc229f7f7, 32'hc2800d50};
test_bias[818:818] = '{32'h42659d19};
test_output[818:818] = '{32'hc5ea485a};
test_input[6552:6559] = '{32'h3f211488, 32'hc1acba73, 32'h42b30607, 32'hc1637f4a, 32'hc09064ff, 32'hc26c21f5, 32'hc1e1f2ee, 32'h4223a8b2};
test_weights[6552:6559] = '{32'h41a9cfba, 32'hbf5c13f7, 32'hc251fc51, 32'h41adc846, 32'h41cf46e6, 32'h42bb092a, 32'hc28e2228, 32'hc2372157};
test_bias[819:819] = '{32'hc1c445b6};
test_output[819:819] = '{32'hc6242067};
test_input[6560:6567] = '{32'hc2053e04, 32'h42b6065e, 32'h424fab2f, 32'hc2b157b9, 32'h424c1c7d, 32'h42c4d10b, 32'h42c73bb2, 32'hc22019ab};
test_weights[6560:6567] = '{32'hc21853e1, 32'hbeb3b9c4, 32'hc29a2255, 32'h4278b7ad, 32'h42b25f1f, 32'h42559cbe, 32'hc2ad60f8, 32'h41006b7b};
test_bias[820:820] = '{32'hc29ba924};
test_output[820:820] = '{32'hc5ea9492};
test_input[6568:6575] = '{32'hc2ad60bd, 32'h421dedc6, 32'h420548c0, 32'h4203eb32, 32'hc1c52f17, 32'hc2bf2998, 32'hc2bf006d, 32'hc295e091};
test_weights[6568:6575] = '{32'h415b50e2, 32'hc2215f56, 32'hc29cce42, 32'hc0d1b11a, 32'h42855c07, 32'hc248ed9a, 32'hc2b9db74, 32'hc29ce7b8};
test_bias[821:821] = '{32'hc224bb72};
test_output[821:821] = '{32'h463f92fb};
test_input[6576:6583] = '{32'h40a0d11b, 32'hc29a383d, 32'h41db9f9e, 32'hc28eebcc, 32'hc205499a, 32'h4105b200, 32'hc27c54d7, 32'h427a2a89};
test_weights[6576:6583] = '{32'hc270b6d3, 32'h42ae9de8, 32'h42af97d1, 32'hc285a74b, 32'hc242d8a8, 32'h422d334e, 32'hc2a5d4c8, 32'hc29b9cfa};
test_bias[822:822] = '{32'hc282376d};
test_output[822:822] = '{32'h45183416};
test_input[6584:6591] = '{32'h42b15039, 32'h4272e162, 32'hc2a21c2e, 32'h424556b9, 32'h4218ac7a, 32'h4184bda7, 32'h426cbab0, 32'h420583c6};
test_weights[6584:6591] = '{32'h4292e001, 32'h41d7ffea, 32'h4294d069, 32'hc28bd096, 32'hc1add934, 32'hc180ae2f, 32'hc1c825e8, 32'h4239497b};
test_bias[823:823] = '{32'hc2393664};
test_output[823:823] = '{32'hc5166e3f};
test_input[6592:6599] = '{32'h4256e1d5, 32'h415e2df3, 32'h42acd22d, 32'h41e34537, 32'h42c5400e, 32'h421fb41a, 32'h428c38ee, 32'h424ec9ee};
test_weights[6592:6599] = '{32'h4101ce03, 32'hc1522a9e, 32'hc29ed55a, 32'hc1ebb12c, 32'hc26c575f, 32'hc20ba9f5, 32'h428ed40b, 32'hc2928345};
test_bias[824:824] = '{32'h41e2348b};
test_output[824:824] = '{32'hc651ad16};
test_input[6600:6607] = '{32'h4270be53, 32'hc2964285, 32'hc2bc49ee, 32'h42b4e302, 32'h42ab3f20, 32'h42022e72, 32'hbf2ac056, 32'h42b73b5d};
test_weights[6600:6607] = '{32'h41554506, 32'h41c7fb9e, 32'h426a668e, 32'hc2434092, 32'h4246415d, 32'h421cd313, 32'h422fd32d, 32'h429e10f8};
test_bias[825:825] = '{32'h42561e55};
test_output[825:825] = '{32'h44de2521};
test_input[6608:6615] = '{32'hc28c8e9a, 32'h4271e3b0, 32'hc27176dc, 32'hc2c4d0e2, 32'h4097fe66, 32'h41c90b7b, 32'h422b0c36, 32'h42451412};
test_weights[6608:6615] = '{32'h418f6988, 32'hc20a71e4, 32'h4190ac7e, 32'hc149eb72, 32'hc28dfc8b, 32'h4228809b, 32'h42ac5584, 32'h42ae49c5};
test_bias[826:826] = '{32'hc0fbbda1};
test_output[826:826] = '{32'h45ab893b};
test_input[6616:6623] = '{32'h42977092, 32'h42b31e2f, 32'hc2a324a8, 32'h423c2b58, 32'hc20b04f9, 32'hc2bd3e22, 32'hc2883445, 32'hc0ae065e};
test_weights[6616:6623] = '{32'hc2196bdb, 32'h421913b5, 32'h42c72be8, 32'hc2b3f15e, 32'hc133ec2c, 32'h4223a652, 32'hc15b1bc0, 32'hc0b05ae6};
test_bias[827:827] = '{32'h428d8243};
test_output[827:827] = '{32'hc65f1f16};
test_input[6624:6631] = '{32'h427a538d, 32'hc1fe84d8, 32'hc1e8033e, 32'h427fbaf6, 32'hc2074f8d, 32'hc23aa7e3, 32'h416b2dfb, 32'hc18a0420};
test_weights[6624:6631] = '{32'h42183319, 32'h42a36659, 32'h4098c5cd, 32'h42b58365, 32'hc2aedc5d, 32'hc2613921, 32'hc2c44977, 32'h4241e9ba};
test_bias[828:828] = '{32'h42b87007};
test_output[828:828] = '{32'h460a306c};
test_input[6632:6639] = '{32'h4280d463, 32'hc0b5e41b, 32'hc2208cce, 32'hc2b7d075, 32'hc29da5fc, 32'h42b626f5, 32'hc1fba482, 32'hc1a2f89c};
test_weights[6632:6639] = '{32'h41cd0090, 32'hc294d839, 32'h42979f1c, 32'h42a18dda, 32'h41e6d57a, 32'hc2a01931, 32'h40f6a948, 32'h424928d6};
test_bias[829:829] = '{32'hc1236cd4};
test_output[829:829] = '{32'hc696469b};
test_input[6640:6647] = '{32'h425e5140, 32'h415edac2, 32'hc216aaec, 32'hc2b9a215, 32'hc255b188, 32'hc27f2212, 32'h402b84b4, 32'hc217b642};
test_weights[6640:6647] = '{32'hc1c67b76, 32'hc1957e4e, 32'hc2b49e75, 32'h42aafdfd, 32'hc08fea2d, 32'hc2b3c838, 32'hc28d5aba, 32'h42c00b2d};
test_bias[830:830] = '{32'hc28008bc};
test_output[830:830] = '{32'hc57fe861};
test_input[6648:6655] = '{32'hc099db6f, 32'hc24cd503, 32'h429e86e0, 32'h428fb42d, 32'h406ab3db, 32'h41b010d5, 32'hc26ae832, 32'h42b4c780};
test_weights[6648:6655] = '{32'hc28772dc, 32'h426c2b48, 32'h4283e13a, 32'h41e8df4b, 32'hc260d3d0, 32'h42c46ca7, 32'h428c2e9a, 32'hc1df6c32};
test_bias[831:831] = '{32'h42540c46};
test_output[831:831] = '{32'hc13e51b2};
test_input[6656:6663] = '{32'hc12eec76, 32'h42bb934e, 32'h41b8969a, 32'hc2b132f1, 32'h428251ae, 32'h40b587dd, 32'hc1fcc6af, 32'hc06534da};
test_weights[6656:6663] = '{32'h42635e20, 32'h42557c65, 32'h42288eb0, 32'hc27432d3, 32'hc1e0a4fb, 32'h413010b7, 32'hc06da43c, 32'hc1ba4929};
test_bias[832:832] = '{32'hc210b36d};
test_output[832:832] = '{32'h460f2ab2};
test_input[6664:6671] = '{32'h41b1730a, 32'h41e47282, 32'h42a28cb0, 32'hc1561b39, 32'h41dbabed, 32'h421841b5, 32'h424847b6, 32'h424ac815};
test_weights[6664:6671] = '{32'hc240e53b, 32'hc286ffe9, 32'h42282b8f, 32'h426a132d, 32'hc2b87f86, 32'hc24c5865, 32'hc192cc41, 32'hc1c3b1ea};
test_bias[833:833] = '{32'hc181c89f};
test_output[833:833] = '{32'hc5db3fd6};
test_input[6672:6679] = '{32'hc2c1c4e7, 32'h42648ad4, 32'hc258843a, 32'h42b6c35b, 32'hc237d1b3, 32'h42b55e1f, 32'hc2bf292e, 32'hc1835e51};
test_weights[6672:6679] = '{32'hc2460f98, 32'h415673ed, 32'h42b21013, 32'h42b077a1, 32'h425589c5, 32'hc2b1b143, 32'hc23ff656, 32'h4137d989};
test_bias[834:834] = '{32'hc20dae36};
test_output[834:834] = '{32'h4526376c};
test_input[6680:6687] = '{32'h426e4824, 32'hc234281a, 32'hc1fb5eb2, 32'h4294ce3b, 32'hc27aca78, 32'h41107cbd, 32'hc2952f60, 32'hc1fde1ea};
test_weights[6680:6687] = '{32'hc24c037a, 32'h41ea514f, 32'h428eb95a, 32'h42887b51, 32'hc19b6bab, 32'h3ffd828e, 32'hc186ee03, 32'hc151ac83};
test_bias[835:835] = '{32'hc2a40046};
test_output[835:835] = '{32'h44a32f0d};
test_input[6688:6695] = '{32'h41f0db3c, 32'h42a20217, 32'hc293b81a, 32'h4200c340, 32'hc1640390, 32'h40856832, 32'hc2adb361, 32'h42922d8b};
test_weights[6688:6695] = '{32'h42675209, 32'hc2835a2a, 32'h423c664c, 32'hc0282fcb, 32'hc2b6590c, 32'hbf31a501, 32'hc2a81897, 32'hc0fd49eb};
test_bias[836:836] = '{32'h414e1999};
test_output[836:836] = '{32'h445e043d};
test_input[6696:6703] = '{32'h42132872, 32'h424b57a6, 32'hc13b7d64, 32'hc1c580b0, 32'hc29f6003, 32'hc2a641ad, 32'hc1e415a4, 32'hc08a2a7e};
test_weights[6696:6703] = '{32'h415205dd, 32'hc1fae019, 32'h42bc6f73, 32'hc1f3752e, 32'h4273e238, 32'hc2682e2c, 32'hc2b6efca, 32'h41b8f2e3};
test_bias[837:837] = '{32'h428106fd};
test_output[837:837] = '{32'h44866229};
test_input[6704:6711] = '{32'h4132b7ab, 32'hc2b242eb, 32'h41ee93bb, 32'h421fea3d, 32'h4180afc2, 32'hc2b11cdd, 32'h41ccd08b, 32'hc170764d};
test_weights[6704:6711] = '{32'hc21d7310, 32'h421595e3, 32'hc29aabc5, 32'h42089e64, 32'hc2ae2723, 32'hbffac21f, 32'hc287940e, 32'hc27d4a10};
test_bias[838:838] = '{32'h41388f02};
test_output[838:838] = '{32'hc5d1c9c6};
test_input[6712:6719] = '{32'h426dffc1, 32'hc20959bd, 32'h422292df, 32'h4222355d, 32'hc16795a5, 32'hc2af511d, 32'hc2aa0925, 32'h427da045};
test_weights[6712:6719] = '{32'h413abece, 32'h40e2a223, 32'hc2c48a97, 32'hc28f724d, 32'hc2206504, 32'h423f6aae, 32'hc19d3313, 32'hc2171a6f};
test_bias[839:839] = '{32'h421b7c44};
test_output[839:839] = '{32'hc627fe13};
test_input[6720:6727] = '{32'h42a76cc1, 32'hc2ba0ac6, 32'h42847cad, 32'hc1eab269, 32'h423288ed, 32'h420a4776, 32'hc207ddab, 32'h42c37627};
test_weights[6720:6727] = '{32'hc2bbb0eb, 32'h41d234a1, 32'hc0e4c538, 32'h41445c19, 32'hc144570c, 32'h4213c863, 32'h424a806a, 32'hc0c4cef9};
test_bias[840:840] = '{32'hc20cb089};
test_output[840:840] = '{32'hc64760a9};
test_input[6728:6735] = '{32'hc2bb47cf, 32'hc2b3d9fb, 32'hc24f884d, 32'hbfc9d9f0, 32'h42a69de0, 32'hc2bc7c33, 32'hc28840e6, 32'hc260064a};
test_weights[6728:6735] = '{32'h424516d3, 32'h41ac0b1f, 32'h425daf29, 32'hc1f33ef9, 32'hc1210096, 32'hc24e6c54, 32'h4202fcdc, 32'hbe89d082};
test_bias[841:841] = '{32'h41b97391};
test_output[841:841] = '{32'hc5ebb609};
test_input[6736:6743] = '{32'hc2b2fb01, 32'h419c3215, 32'hc22b3efd, 32'hbf87fc6e, 32'hc26a93f9, 32'h42b04e6e, 32'hc1823bfb, 32'hc2bb9c8e};
test_weights[6736:6743] = '{32'hc2977562, 32'hc297ba31, 32'h425c2474, 32'hc241e114, 32'hc2511832, 32'h414e1e00, 32'hc1213aa6, 32'h4129d9dc};
test_bias[842:842] = '{32'h42401941};
test_output[842:842] = '{32'h45c844d6};
test_input[6744:6751] = '{32'h429c6da5, 32'hc27c0d33, 32'hc21e6577, 32'hc1ce7013, 32'hc2781708, 32'hc2a86db9, 32'hc2564a97, 32'h415dc5d8};
test_weights[6744:6751] = '{32'h42394622, 32'h3fc5f89b, 32'hc0f5739b, 32'h4289f314, 32'h428b29e8, 32'hc15694c9, 32'h4157a954, 32'hc17bb0bc};
test_bias[843:843] = '{32'h3f48309e};
test_output[843:843] = '{32'hc501c67a};
test_input[6752:6759] = '{32'h41c823af, 32'h4224a0ff, 32'hc20902e0, 32'h415dbfb5, 32'hc1c2c885, 32'hc2719c44, 32'hc027d024, 32'h427a79cd};
test_weights[6752:6759] = '{32'hc2ab72b1, 32'hc1a4d316, 32'h402e54ec, 32'hc25c523e, 32'hc1134729, 32'h42b23e59, 32'h42b73577, 32'h41857477};
test_bias[844:844] = '{32'h42704522};
test_output[844:844] = '{32'hc5fe7ea2};
test_input[6760:6767] = '{32'hc20f0c54, 32'hc1443b2d, 32'hc18cb150, 32'h420cde57, 32'h40e97c6c, 32'hc1dc01cb, 32'hc2bee7fc, 32'hc16ec60b};
test_weights[6760:6767] = '{32'hc260f989, 32'hc2556128, 32'h41ea2e6d, 32'h42a522d1, 32'hc2c753a0, 32'h42119a3c, 32'h40ec4232, 32'hc1bc8938};
test_bias[845:845] = '{32'hc08bf6cc};
test_output[845:845] = '{32'h4539cfca};
test_input[6768:6775] = '{32'h41e835a9, 32'hc21a212e, 32'hc2876cfc, 32'hc235c971, 32'hc26fabfd, 32'h42254163, 32'hc1b21c7b, 32'hc2650ee2};
test_weights[6768:6775] = '{32'h424e6e40, 32'hc1ba515f, 32'hc118df75, 32'hc0e296d8, 32'hc264fc8a, 32'h428b871f, 32'hc28e5b06, 32'h42b7c832};
test_bias[846:846] = '{32'h4160fe2d};
test_output[846:846] = '{32'h45bbe910};
test_input[6776:6783] = '{32'h42c757fa, 32'h4273be6e, 32'h41977f4d, 32'h42228c45, 32'hc2984c78, 32'h421636d6, 32'hc20cd92b, 32'h428f955c};
test_weights[6776:6783] = '{32'hc0ceacb7, 32'h42b9504a, 32'h41d0a00b, 32'h42831c6d, 32'hc22dadd2, 32'h41e9c113, 32'h41c85a69, 32'h42aadbd5};
test_bias[847:847] = '{32'hc18fefc4};
test_output[847:847] = '{32'h468b0a53};
test_input[6784:6791] = '{32'h42b5c42b, 32'hc2941d8b, 32'hc1fea342, 32'h419d4480, 32'h429ea191, 32'hc10ca9ca, 32'hc20fc3d2, 32'h4285b521};
test_weights[6784:6791] = '{32'hc2811b9c, 32'h42bd7f0c, 32'hc2c3c706, 32'hc2bbd153, 32'hbfd5efb7, 32'h416edcef, 32'h429a0ec3, 32'h4098d207};
test_bias[848:848] = '{32'h42bb0b95};
test_output[848:848] = '{32'hc65e663b};
test_input[6792:6799] = '{32'hc2138433, 32'h4206bd60, 32'h3fdff9fc, 32'h42c36de0, 32'h424fd1c0, 32'h42803dd8, 32'h4271909d, 32'h42502bc0};
test_weights[6792:6799] = '{32'h427a0812, 32'hc2b21a76, 32'hc15c76d7, 32'hc27976ad, 32'h426a73c4, 32'h41714d9f, 32'h421995fd, 32'h428b0181};
test_bias[849:849] = '{32'h4243cbf0};
test_output[849:849] = '{32'hc4b23e9b};
test_input[6800:6807] = '{32'h4288fdfc, 32'hc1a6e917, 32'hc25b2551, 32'h4021dff8, 32'hc21384fd, 32'h401b8b34, 32'h421a5c36, 32'h424cbd79};
test_weights[6800:6807] = '{32'h42ac486a, 32'hc27209a9, 32'hc190106c, 32'h4205ba1a, 32'h40f2ba77, 32'h42a490e0, 32'h427dd166, 32'h42aebd09};
test_bias[850:850] = '{32'h42ac6d8f};
test_output[850:850] = '{32'h466ce478};
test_input[6808:6815] = '{32'hc231ad33, 32'hc29a5c05, 32'h403c99d5, 32'hc28afd7b, 32'h42529d8f, 32'hc1017af8, 32'h4280d177, 32'hc2ae2cbd};
test_weights[6808:6815] = '{32'hc2a328d5, 32'hc2c10bf4, 32'h429f3867, 32'hc299323b, 32'hc250139b, 32'hc185c62a, 32'h42976786, 32'h40be011d};
test_bias[851:851] = '{32'hc237c0a6};
test_output[851:851] = '{32'h468f48ab};
test_input[6816:6823] = '{32'hc2997c43, 32'hc1dc7a60, 32'h42b41b42, 32'hc12ddcd3, 32'h401ee8c2, 32'h427bf37f, 32'hc27e43ac, 32'h4184e7c1};
test_weights[6816:6823] = '{32'hc205d348, 32'hc2762755, 32'h3f6eca88, 32'hc20e2bb5, 32'hc2abb753, 32'hc2b664c7, 32'h4231ca5b, 32'hc08aff29};
test_bias[852:852] = '{32'h40a757e6};
test_output[852:852] = '{32'hc580a039};
test_input[6824:6831] = '{32'h41ac2db7, 32'h420685b6, 32'hc21230d1, 32'h42640e0e, 32'h409ee0d9, 32'hc210a925, 32'hc29ae16e, 32'hc239cee7};
test_weights[6824:6831] = '{32'h415e06a3, 32'h4292e18f, 32'h42b7d091, 32'h4173635d, 32'hc2136164, 32'hc217b8f2, 32'hc18ad304, 32'hc204b7c1};
test_bias[853:853] = '{32'h425c6160};
test_output[853:853] = '{32'h4589ae52};
test_input[6832:6839] = '{32'hc1d30c72, 32'hc2922946, 32'hc1919e9d, 32'hc1ec3a30, 32'h428c5ffa, 32'h4260eed2, 32'h42a4a44d, 32'h41394ade};
test_weights[6832:6839] = '{32'h421896b0, 32'h42151490, 32'h4136edab, 32'h41f28f2e, 32'hc282afdf, 32'hc23b4ca3, 32'hc280a29c, 32'h42a55a6a};
test_bias[854:854] = '{32'h429e980b};
test_output[854:854] = '{32'hc67edb4b};
test_input[6840:6847] = '{32'hc1014ea1, 32'hc08becc4, 32'h422c8e77, 32'h41d7a5f3, 32'h42a00420, 32'h424d7dd3, 32'h40ed4ee3, 32'hc268a458};
test_weights[6840:6847] = '{32'hc18523cb, 32'hc2c0e2e5, 32'hc2c18789, 32'hc1ab3904, 32'h42b32535, 32'hc1f68d98, 32'hc26299b3, 32'h4226e1ef};
test_bias[855:855] = '{32'h423581ab};
test_output[855:855] = '{32'hc4b0a0e4};
test_input[6848:6855] = '{32'h42607145, 32'h415c4906, 32'hc1f5f8fd, 32'hc1c9928d, 32'hbf129bb2, 32'h4123a547, 32'hc20d440e, 32'h414b02e2};
test_weights[6848:6855] = '{32'h4259c9e7, 32'hc27dedbb, 32'h40ecdc6f, 32'hc1c9479b, 32'hc2c08a41, 32'h41f2d58f, 32'h42b50553, 32'hc26e0540};
test_bias[856:856] = '{32'hc2028121};
test_output[856:856] = '{32'hc480e47f};
test_input[6856:6863] = '{32'hc1cb5c30, 32'h421d18fb, 32'h41121fa0, 32'hc284cbc9, 32'hc271398e, 32'hc21466f5, 32'hc11fb45d, 32'h429d4fc1};
test_weights[6856:6863] = '{32'h42621c84, 32'hc2b08180, 32'h41a13189, 32'h42254743, 32'h42ba39e6, 32'hc26b3f92, 32'h41f2cb7d, 32'h418f9116};
test_bias[857:857] = '{32'h424ce99d};
test_output[857:857] = '{32'hc6182027};
test_input[6864:6871] = '{32'h42627f97, 32'h3fcc1cef, 32'hc232eb5c, 32'hc2627133, 32'h416586fb, 32'hc20f4735, 32'hc2849751, 32'hc2324abb};
test_weights[6864:6871] = '{32'h427b51b9, 32'h40daaf07, 32'hc2b7ce3c, 32'hc2bf6b32, 32'h42b910c4, 32'h42aba035, 32'hc1ee8e7a, 32'hc157a0a4};
test_bias[858:858] = '{32'hc19725f2};
test_output[858:858] = '{32'h465957b0};
test_input[6872:6879] = '{32'h41a96366, 32'hc24c54f8, 32'hc2c77c93, 32'h42212c3b, 32'h4202b635, 32'h429cdb6e, 32'h4209c72c, 32'hc257b6a1};
test_weights[6872:6879] = '{32'hc29bba50, 32'hc23bfbfa, 32'hc235bbda, 32'h40648ea9, 32'h40e9e558, 32'hc25fb4d6, 32'h41ee1a4c, 32'hc10418ee};
test_bias[859:859] = '{32'h42c63202};
test_output[859:859] = '{32'h45321bb7};
test_input[6880:6887] = '{32'h42575352, 32'h41d4a660, 32'h424738a0, 32'h40a7387f, 32'h4219c6ed, 32'h40e61f41, 32'h41bc707e, 32'h4264e986};
test_weights[6880:6887] = '{32'h42888c22, 32'h41dff071, 32'h3fdca37f, 32'h42c2013f, 32'hc2b6ac36, 32'h4235e91a, 32'h401f40dd, 32'h425ba835};
test_bias[860:860] = '{32'h42a5df2f};
test_output[860:860] = '{32'h459fbfaf};
test_input[6888:6895] = '{32'h425554f8, 32'hc08b2a43, 32'hc2afce64, 32'h426e5640, 32'h424b2bbc, 32'hc1d8c278, 32'h427ba4ea, 32'h42a23e73};
test_weights[6888:6895] = '{32'hc2917d0f, 32'hc280361a, 32'h42521303, 32'h41b615e8, 32'hc29e2842, 32'h40dc25b5, 32'hc2368c48, 32'h408fd521};
test_bias[861:861] = '{32'hc1de215a};
test_output[861:861] = '{32'hc65479ea};
test_input[6896:6903] = '{32'hc254e1ee, 32'h42b9267c, 32'h421dcc19, 32'h41d8ecfa, 32'hc284f9b7, 32'hc2c10c72, 32'h427c2fad, 32'h4215cb73};
test_weights[6896:6903] = '{32'hc2812b32, 32'hc295a409, 32'hc0a36d04, 32'hc1e05fa9, 32'hc2a9d0d6, 32'h4260afea, 32'h4257b4b9, 32'h42861d88};
test_bias[862:862] = '{32'h42a8f378};
test_output[862:862] = '{32'h44dcf66f};
test_input[6904:6911] = '{32'hc20aaf41, 32'hc2ab67a7, 32'h4181db02, 32'h4188de6f, 32'hc1b154ea, 32'hc29be8ad, 32'hc21a2574, 32'hc1db3d59};
test_weights[6904:6911] = '{32'hc2257fc4, 32'hc27016b5, 32'hc21f9bb6, 32'h4297420b, 32'h428ba99c, 32'hc28facd6, 32'h4208ef21, 32'h41e68fd9};
test_bias[863:863] = '{32'h428c2c0e};
test_output[863:863] = '{32'h461057cb};
test_input[6912:6919] = '{32'h41173542, 32'h423ea210, 32'h421e9e54, 32'h421523d9, 32'hc1b96fd5, 32'hc2c0500a, 32'h42a7fdf3, 32'hc09ab79e};
test_weights[6912:6919] = '{32'hc2a96e50, 32'h41cc8bcc, 32'hc2619a54, 32'h428f1c39, 32'hc29c9a9b, 32'h42ad3be4, 32'h42b34b49, 32'h42171255};
test_bias[864:864] = '{32'h420dbe82};
test_output[864:864] = '{32'h44d6cc3b};
test_input[6920:6927] = '{32'hc26be95d, 32'h4137a5ca, 32'hc2c33559, 32'h420f1d90, 32'hc25d0b7a, 32'h426c9387, 32'h4298b413, 32'hc24189b7};
test_weights[6920:6927] = '{32'hc1b2aa87, 32'hc256836b, 32'hc1b9443a, 32'hc24ed949, 32'hc1cb3c7f, 32'h421744ca, 32'h41e3a06b, 32'hc2a86a24};
test_bias[865:865] = '{32'h42a594d0};
test_output[865:865] = '{32'h462d2794};
test_input[6928:6935] = '{32'hc24877ea, 32'h41114e3f, 32'h42a46b8e, 32'h4255cb81, 32'hc140552e, 32'h40449983, 32'h428bd09e, 32'h3ff4738b};
test_weights[6928:6935] = '{32'hc247cbce, 32'hc2a786a6, 32'h428861e3, 32'hc2ab8975, 32'h3f862d79, 32'h42a2ab31, 32'h425f9840, 32'hc230e5a7};
test_bias[866:866] = '{32'h402dec57};
test_output[866:866] = '{32'h45d55d01};
test_input[6936:6943] = '{32'h424b1c61, 32'hc1b0ec72, 32'h42bbf309, 32'h41e8f8c1, 32'hc1cc37a2, 32'hc1bc68d7, 32'h42a7f9b5, 32'hc20a0691};
test_weights[6936:6943] = '{32'h4166828e, 32'hc2a024a2, 32'h4249d636, 32'h3f31e88d, 32'h42ada31e, 32'hc1fec5f8, 32'hc1966289, 32'hc2a56773};
test_bias[867:867] = '{32'h409f5170};
test_output[867:867] = '{32'h45dd31a4};
test_input[6944:6951] = '{32'hc0cf9b64, 32'h41345240, 32'hc2838014, 32'h42a8a549, 32'h42b1934e, 32'hc10a38f2, 32'h40adf0bf, 32'hc271b4dd};
test_weights[6944:6951] = '{32'h41bf82da, 32'hc2982a6f, 32'h42866766, 32'hc29e3266, 32'h42964cbc, 32'hc0fc25df, 32'hc2b19ad8, 32'hc200e0c4};
test_bias[868:868] = '{32'hc199bd65};
test_output[868:868] = '{32'hc574ba79};
test_input[6952:6959] = '{32'h41ba1fa3, 32'hc2bf772d, 32'hc28f6733, 32'hc2a9c994, 32'h42b2abe7, 32'hc2c32cef, 32'h42b639da, 32'h42b90f64};
test_weights[6952:6959] = '{32'hc2215774, 32'h41c29cfe, 32'hc285c7e7, 32'h423ee6ea, 32'h4284fcd7, 32'h42261529, 32'hc29a31c1, 32'h4276f1bc};
test_bias[869:869] = '{32'hc1c73cc6};
test_output[869:869] = '{32'hc4f66c00};
test_input[6960:6967] = '{32'h426ae8de, 32'h424218be, 32'hc2695ad7, 32'hc25a2642, 32'h418ce8f6, 32'hc26aeb05, 32'h41a31976, 32'hc29f4d98};
test_weights[6960:6967] = '{32'hc2a994ac, 32'h42a721bd, 32'hc2027f06, 32'hc07a07c8, 32'hc2a66dd0, 32'h42c2c129, 32'hc2acb647, 32'hc27d70c1};
test_bias[870:870] = '{32'h423ef27d};
test_output[870:870] = '{32'hc5262fe9};
test_input[6968:6975] = '{32'hc2609f56, 32'h42379a7e, 32'h42469d4b, 32'hc1910bd3, 32'h4262e487, 32'hc11db01c, 32'hc1cf300a, 32'hc2b0c70b};
test_weights[6968:6975] = '{32'hc2842f1b, 32'hc2bf51f1, 32'h42b59e91, 32'hc1175533, 32'hc281d135, 32'h428dd967, 32'h41dd6b80, 32'hc27bc264};
test_bias[871:871] = '{32'h42486aed};
test_output[871:871] = '{32'h458d25cf};
test_input[6976:6983] = '{32'hc28cc489, 32'h420dd5b1, 32'h429b12b1, 32'h3f857d6b, 32'h42b393af, 32'hc2129b87, 32'h42429e0a, 32'hc2825638};
test_weights[6976:6983] = '{32'hc217c1f8, 32'hc287c103, 32'hc27e520e, 32'hbe1d6eec, 32'h428368c3, 32'h41913289, 32'h4194204c, 32'hc277138b};
test_bias[872:872] = '{32'hc08511a6};
test_output[872:872] = '{32'h45ab8fa3};
test_input[6984:6991] = '{32'hc289f4f6, 32'hc29da5ce, 32'hc1ddc373, 32'hc1ffdebc, 32'hc2ad5493, 32'h427ab790, 32'hc175e5f7, 32'h40352931};
test_weights[6984:6991] = '{32'hc22341b3, 32'h40a2811a, 32'h426188d5, 32'hc2af90e3, 32'h415a05ed, 32'hc1c7f993, 32'hc1ef7533, 32'h420c5e14};
test_bias[873:873] = '{32'hc1f4339c};
test_output[873:873] = '{32'h44b4185f};
test_input[6992:6999] = '{32'hc28c724c, 32'h42b507d3, 32'h422677bb, 32'h4292c7be, 32'hc241d918, 32'hc1c4e37f, 32'hc21ad1d0, 32'h42b1d10c};
test_weights[6992:6999] = '{32'hc2181fb1, 32'hc2a1a789, 32'hc2b7b0f2, 32'h426ab513, 32'hc0c57c94, 32'h4217fb6b, 32'h4225d9e9, 32'hc2a84de2};
test_bias[874:874] = '{32'hc2085e9d};
test_output[874:874] = '{32'hc65978ed};
test_input[7000:7007] = '{32'hc29c7ff1, 32'hc224ec35, 32'hc22f2b6b, 32'hc2929cec, 32'h418fd8b1, 32'hc29167de, 32'hc2a5a123, 32'h42c3cd14};
test_weights[7000:7007] = '{32'h42286e63, 32'hc24b4fa0, 32'h42a86322, 32'h42b1ecba, 32'h4283d3c2, 32'hc282c026, 32'hc2b2d3b9, 32'h423e7653};
test_bias[875:875] = '{32'h41a79b0c};
test_output[875:875] = '{32'h45ceccf2};
test_input[7008:7015] = '{32'hc19f3c5d, 32'hc2bedc2c, 32'h41f62c16, 32'h416607be, 32'hc28d6813, 32'hc25ff777, 32'h423c5186, 32'h42a48345};
test_weights[7008:7015] = '{32'hc2ba839a, 32'hc26dd15f, 32'hc0bd185d, 32'hc239b218, 32'h42a707f5, 32'h421109a5, 32'h4150d491, 32'h429066c0};
test_bias[876:876] = '{32'h42927341};
test_output[876:876] = '{32'h45a7e2a4};
test_input[7016:7023] = '{32'h423004e5, 32'h40307c74, 32'hc24c6ad8, 32'h428b1e4d, 32'h41c05273, 32'hc292a64f, 32'h42572981, 32'h4205df98};
test_weights[7016:7023] = '{32'h423f4d1e, 32'hc257ec52, 32'h42c5e74d, 32'h41a562f7, 32'h41f8fe44, 32'hc1dbbf7f, 32'h4280031a, 32'h415064b6};
test_bias[877:877] = '{32'hc2a3d2ad};
test_output[877:877] = '{32'h459900ec};
test_input[7024:7031] = '{32'hc2b691bb, 32'h4221e353, 32'hc04e0574, 32'h42a1a5f2, 32'hc1026f06, 32'hc23faf4d, 32'hc22c993b, 32'hc2868e08};
test_weights[7024:7031] = '{32'hc2be34a7, 32'hc2b682e3, 32'hc1002f26, 32'h41b78b5d, 32'hc2ae7f9e, 32'hc25dcfdb, 32'hc2c5567f, 32'h41c67792};
test_bias[878:878] = '{32'hc20d62a6};
test_output[878:878] = '{32'h4647d831};
test_input[7032:7039] = '{32'hc06dca57, 32'h41d32af6, 32'hc2a1eb89, 32'hc144c362, 32'h41c94bdd, 32'h423c97ed, 32'hc2b442d8, 32'hc25f3b24};
test_weights[7032:7039] = '{32'hc2852e43, 32'h42b5a507, 32'hc2be5a9b, 32'hc2aa5f02, 32'h42badb5f, 32'hc20d6e6a, 32'hc00e00b1, 32'h42124362};
test_bias[879:879] = '{32'h4251c6ad};
test_output[879:879] = '{32'h4620d5ba};
test_input[7040:7047] = '{32'h429bee22, 32'h4292b4c7, 32'hc21fafbe, 32'h4264068d, 32'h42bbe8d5, 32'hbf882acc, 32'h42b27690, 32'hc2895a9e};
test_weights[7040:7047] = '{32'h414f68a8, 32'h427cf517, 32'h428e2c79, 32'hc2570545, 32'hc23653e0, 32'h42abb00b, 32'hc18bcbbc, 32'h41d3c100};
test_bias[880:880] = '{32'h413f6998};
test_output[880:880] = '{32'hc5f9bf5f};
test_input[7048:7055] = '{32'h42b05533, 32'hc21235b4, 32'hc18defdb, 32'h41cc2ae3, 32'h41a7c41c, 32'h428b9a1b, 32'h42a0fa2a, 32'hc2402d8a};
test_weights[7048:7055] = '{32'hc29092d4, 32'h4143b631, 32'h4296ceb4, 32'hc23ccba4, 32'h42851050, 32'hc2859694, 32'hc2bef180, 32'hc08af6fe};
test_bias[881:881] = '{32'h42879066};
test_output[881:881] = '{32'hc69c8b92};
test_input[7056:7063] = '{32'h4197cc22, 32'h427ff886, 32'hc2c3b7e7, 32'h424d0069, 32'hc2b6fa27, 32'h41ea3adb, 32'h4162580d, 32'h42c08c5b};
test_weights[7056:7063] = '{32'hc2111162, 32'h422d0c06, 32'h427a8a14, 32'h42c6a1be, 32'hc01ab59f, 32'hc2b25645, 32'hc2bec776, 32'h40bcda73};
test_bias[882:882] = '{32'h4210dd42};
test_output[882:882] = '{32'hc502dc00};
test_input[7064:7071] = '{32'hc19437d6, 32'h427c0d17, 32'hc21c0591, 32'h4116aee7, 32'h42979bf4, 32'hc2b7d4ca, 32'hc2748446, 32'h41ff4d1e};
test_weights[7064:7071] = '{32'hc29a5ca0, 32'h429103af, 32'h42a64f64, 32'hc2b9d158, 32'hc265290c, 32'hbe86c22d, 32'hc2a78134, 32'hc283dab9};
test_bias[883:883] = '{32'h412eb53a};
test_output[883:883] = '{32'h441319ce};
test_input[7072:7079] = '{32'h41dba2ac, 32'h4259de51, 32'hc16fbe94, 32'hc1e6d304, 32'h429d50cb, 32'h422c4ba2, 32'hc247e8b5, 32'h41cdc8ea};
test_weights[7072:7079] = '{32'h41edd28d, 32'hc2b55461, 32'h427c3032, 32'h4280b30b, 32'hc23da31a, 32'hc21d7de1, 32'hc29b6776, 32'hc2a54557};
test_bias[884:884] = '{32'hc29708f7};
test_output[884:884] = '{32'hc626a963};
test_input[7080:7087] = '{32'h429f69a4, 32'h427cf734, 32'h42479335, 32'h421ffb90, 32'hc224d0ab, 32'hc2b9f57f, 32'hc28a809f, 32'h42874e39};
test_weights[7080:7087] = '{32'hc2c5a61c, 32'h40d2a582, 32'hc1d4412e, 32'h428596e3, 32'hc296ad4e, 32'h420cd2af, 32'hc1b867c6, 32'hc2389849};
test_bias[885:885] = '{32'h41176ca7};
test_output[885:885] = '{32'hc5f3b36a};
test_input[7088:7095] = '{32'hc271db02, 32'h3e7e10b3, 32'h42911ec3, 32'h41cd5ddf, 32'hc064a305, 32'hc2872f35, 32'h420e5450, 32'h4266d20b};
test_weights[7088:7095] = '{32'hc1f6556d, 32'h42555350, 32'hc2a66765, 32'hc25ef88a, 32'h42b29d34, 32'h429bdf10, 32'hc2c3b490, 32'hc10c07dd};
test_bias[886:886] = '{32'h423e5c3c};
test_output[886:886] = '{32'hc66c3cf5};
test_input[7096:7103] = '{32'hc17ecac4, 32'h40f49d82, 32'h42a64544, 32'hc2953091, 32'hc226da01, 32'hc227a6fb, 32'hbf573dc0, 32'h422308c2};
test_weights[7096:7103] = '{32'h429cde7e, 32'hc241cd3e, 32'hc26fd40c, 32'hc234e6df, 32'h42c1760e, 32'hc29a64a5, 32'h420879bb, 32'hc2c230f8};
test_bias[887:887] = '{32'hc220c187};
test_output[887:887] = '{32'hc5fbc0a3};
test_input[7104:7111] = '{32'h40dce251, 32'h41aecc9b, 32'h42ac6cf7, 32'h42441f44, 32'hc2ada59f, 32'hc2a48391, 32'hc2111456, 32'hc2ac2539};
test_weights[7104:7111] = '{32'h41ef380c, 32'h4207d449, 32'hc1ad4643, 32'hc251f808, 32'h429579f0, 32'h429f5812, 32'h42aaba85, 32'hc11d65e9};
test_bias[888:888] = '{32'hc2848a57};
test_output[888:888] = '{32'hc69345eb};
test_input[7112:7119] = '{32'h429144ad, 32'hc2136edf, 32'h42acd5f6, 32'hc2927960, 32'hc1a6381f, 32'hc2ad3495, 32'h42bb5081, 32'h42b81542};
test_weights[7112:7119] = '{32'h4199ed2d, 32'hc2c19a7e, 32'h428104c2, 32'h41779382, 32'hc14cd343, 32'h4272b030, 32'hc1ac035d, 32'hc18b4642};
test_bias[889:889] = '{32'hc280dc65};
test_output[889:889] = '{32'h44388210};
test_input[7120:7127] = '{32'h426621da, 32'hc28714b3, 32'hc1f5d656, 32'h4241c566, 32'h42a00084, 32'hc2c1e071, 32'hc25f29d6, 32'hc1302b02};
test_weights[7120:7127] = '{32'hc2aea726, 32'hc1971fd6, 32'hc2bcad72, 32'hc2a194ea, 32'h428f7d7d, 32'h41d82c6a, 32'hc269d25e, 32'hbf246948};
test_bias[890:890] = '{32'hc1005ddf};
test_output[890:890] = '{32'h44ca31a3};
test_input[7128:7135] = '{32'h41f39e62, 32'hc18ba134, 32'h41ebe47a, 32'h42ad408e, 32'h428bf354, 32'h420e571a, 32'hc28a0a17, 32'hc201363e};
test_weights[7128:7135] = '{32'h4230c891, 32'hc2077120, 32'h40914a5c, 32'h4186f8ff, 32'hc29a1ad5, 32'hc1804f87, 32'hc25588a0, 32'h4205aa73};
test_bias[891:891] = '{32'hc23c0511};
test_output[891:891] = '{32'h42ff9b9c};
test_input[7136:7143] = '{32'hc1a47b6e, 32'hc17701dd, 32'h427aec88, 32'h42196539, 32'hc2552175, 32'h41eba759, 32'hc29cf8ba, 32'hc2aaa247};
test_weights[7136:7143] = '{32'hc1a1c3a5, 32'h41ffb607, 32'hc0a39bab, 32'hc236acef, 32'hc27b6af4, 32'h4208b7dd, 32'h42ba8080, 32'h42b78211};
test_bias[892:892] = '{32'hc172dd01};
test_output[892:892] = '{32'hc64a709e};
test_input[7144:7151] = '{32'hc277cf80, 32'h41afebf7, 32'hc29a3ccd, 32'h42a6956c, 32'h42aa3038, 32'hc14743be, 32'h401072f0, 32'h4291e42d};
test_weights[7144:7151] = '{32'hc0c519ab, 32'h42b94d42, 32'h42bab364, 32'h418f5e3f, 32'h4283875a, 32'h42562965, 32'h427cc647, 32'hc2685774};
test_bias[893:893] = '{32'hc1991899};
test_output[893:893] = '{32'hc51a79a5};
test_input[7152:7159] = '{32'hc166dbf3, 32'hc166a05c, 32'hc2887ea8, 32'hc2189f3a, 32'hc1a31559, 32'hc1e26fe8, 32'h4209cf17, 32'h421b857a};
test_weights[7152:7159] = '{32'hc24d3201, 32'hc2346782, 32'h4239128f, 32'hc1933ca0, 32'h40b37656, 32'h42973142, 32'hc2c1e8bc, 32'hc29cce5f};
test_bias[894:894] = '{32'hc0059f6c};
test_output[894:894] = '{32'hc617b7cc};
test_input[7160:7167] = '{32'hc2854533, 32'h423aa39d, 32'hc26ebfdd, 32'h4205f66d, 32'h42973e2c, 32'h40114e59, 32'hc03b81a2, 32'hc1f29a1d};
test_weights[7160:7167] = '{32'hc2744b5a, 32'hc12a3a6e, 32'h423aeb28, 32'h3f5ef2d2, 32'hc25d4977, 32'hc19d8222, 32'hc08d7a78, 32'hc212453b};
test_bias[895:895] = '{32'hc2c0d0e1};
test_output[895:895] = '{32'hc5155860};
test_input[7168:7175] = '{32'h42a9fd09, 32'h42acd6b1, 32'hc2058a34, 32'hc29d111e, 32'hc29eff28, 32'hc1c666b6, 32'hc1ce3892, 32'hc0fe196f};
test_weights[7168:7175] = '{32'h4275e146, 32'h416f4021, 32'hc1e317cf, 32'hc120b697, 32'hc280a800, 32'hc12de964, 32'hc2c4cd35, 32'h3fc04636};
test_bias[896:896] = '{32'h405027ea};
test_output[896:896] = '{32'h467c930f};
test_input[7176:7183] = '{32'hc29d1dc9, 32'h4295837e, 32'h4250d4f3, 32'h421cf239, 32'h42bb29a7, 32'h427d05da, 32'h4290b8c2, 32'hc1fcf1d2};
test_weights[7176:7183] = '{32'h4167c562, 32'h422b7dd1, 32'hc220d5cd, 32'hc1a95420, 32'hc28d0dc4, 32'hc2626a17, 32'hc2b32cd8, 32'hc28f798e};
test_bias[897:897] = '{32'hc2ba0d92};
test_output[897:897] = '{32'hc66fda63};
test_input[7184:7191] = '{32'h42ab801d, 32'hc246a7dc, 32'h426ed9de, 32'hc2939485, 32'hbfa16740, 32'h4104289e, 32'hc1de0c64, 32'hc2545bf9};
test_weights[7184:7191] = '{32'hc23b1abe, 32'hc284bff5, 32'h40a85719, 32'h424c3a9d, 32'h42ac388b, 32'h40f3ad4e, 32'h41d468d3, 32'h4206419a};
test_bias[898:898] = '{32'hc27e42ab};
test_output[898:898] = '{32'hc5d46108};
test_input[7192:7199] = '{32'hc1a9a1c6, 32'h42355983, 32'h40cec565, 32'hc1c57e4d, 32'h422da668, 32'hc24da498, 32'h41f150a1, 32'hc296bea5};
test_weights[7192:7199] = '{32'hc274fa1e, 32'hc0861600, 32'h42a32fad, 32'h42a72b2d, 32'h4204e5fa, 32'h42b3f901, 32'h414b2147, 32'hc1c676a9};
test_bias[899:899] = '{32'hc2c43d63};
test_output[899:899] = '{32'hc4b618f1};
test_input[7200:7207] = '{32'hc295aeee, 32'h4244a708, 32'hc1337682, 32'hc2955b5c, 32'h41fde4a8, 32'h42660718, 32'h423730db, 32'hc2a7f42e};
test_weights[7200:7207] = '{32'hc2bd0a7d, 32'hc0327b73, 32'hc2b77cbe, 32'h42715811, 32'h408ca361, 32'hbe451afd, 32'hc25c8567, 32'hc2b25e49};
test_bias[900:900] = '{32'h41a3014a};
test_output[900:900] = '{32'h4605f63c};
test_input[7208:7215] = '{32'h42528f6a, 32'h4141c442, 32'h42269984, 32'hc2364848, 32'h42850f8f, 32'h41accb37, 32'h4219fc5a, 32'hbee7de3b};
test_weights[7208:7215] = '{32'h41914587, 32'h42be9ea2, 32'h4196b344, 32'hc1d72a86, 32'hc292847d, 32'hc2bb7008, 32'hc130f986, 32'h4227697b};
test_bias[901:901] = '{32'hc2a8e8a1};
test_output[901:901] = '{32'hc54eb090};
test_input[7216:7223] = '{32'h42556117, 32'h420f2098, 32'h4284dc2c, 32'h42151263, 32'h42b17b56, 32'h410d84b7, 32'hc1316269, 32'h420ef10b};
test_weights[7216:7223] = '{32'hc17ea9d1, 32'hc20fb127, 32'hc2bc1d3a, 32'h41a84c6f, 32'h429ca9c1, 32'h42c3d91f, 32'hc2a11ea3, 32'h428c8c75};
test_bias[902:902] = '{32'hc28b7f09};
test_output[902:902] = '{32'h455e15a7};
test_input[7224:7231] = '{32'hc2ae23ca, 32'hc2949939, 32'h41fc65ec, 32'h4254b7d9, 32'hc271592d, 32'hc2002739, 32'hc217116c, 32'hc28dc19c};
test_weights[7224:7231] = '{32'hc08f0686, 32'hc1e264f6, 32'h42a2fdb9, 32'hc1fcdf3e, 32'h42250bd8, 32'h429a7185, 32'hc2c66fbb, 32'hc2bce765};
test_bias[903:903] = '{32'hc28c8857};
test_output[903:903] = '{32'h4609574e};
test_input[7232:7239] = '{32'h42900999, 32'hc2ba31aa, 32'hc2af53aa, 32'h40553a2c, 32'h428eab65, 32'hc2baab29, 32'hc1b844cc, 32'h422f289a};
test_weights[7232:7239] = '{32'hc2c2b392, 32'hc2a04d12, 32'h425ba6f7, 32'hc2baec58, 32'hc26f4eda, 32'h42bc2aa2, 32'h41721bf7, 32'h418f68e1};
test_bias[904:904] = '{32'h42874102};
test_output[904:904] = '{32'hc68686d8};
test_input[7240:7247] = '{32'hc195f4d4, 32'h42a2111c, 32'hc1f409f2, 32'hc1809353, 32'h42b1dbaf, 32'h427d76e9, 32'hc298444f, 32'hc18e2334};
test_weights[7240:7247] = '{32'h3f89ded4, 32'h422b14d2, 32'h42a90bfa, 32'h413eadfa, 32'hc2918955, 32'hc203bc80, 32'h421433ee, 32'hc2959a27};
test_bias[905:905] = '{32'hc1f7ed6c};
test_output[905:905] = '{32'hc612f4b2};
test_input[7248:7255] = '{32'h42ba6dfd, 32'h42c56aa6, 32'hc1d4de78, 32'hc2aed758, 32'hc1dbc661, 32'hc20feaa7, 32'h427c8c95, 32'h4251ccc8};
test_weights[7248:7255] = '{32'h42bae2ce, 32'hc1a2223c, 32'h42bff8c3, 32'hc2466f65, 32'hc283f7ab, 32'hc28e9720, 32'h424f04f1, 32'h42b5c45b};
test_bias[906:906] = '{32'hc218d4d2};
test_output[906:906] = '{32'h46a3055c};
test_input[7256:7263] = '{32'hc21db6cc, 32'h426e958d, 32'h42b84217, 32'hc24fabda, 32'h423d0f6b, 32'hc2bfd102, 32'hc23ba89a, 32'hc0f68495};
test_weights[7256:7263] = '{32'hc2394b08, 32'hc26f50f8, 32'hc21c9208, 32'h42a62588, 32'hc233ba02, 32'hc1fb0101, 32'hc28785b5, 32'hc13c66c8};
test_bias[907:907] = '{32'h424fc38b};
test_output[907:907] = '{32'hc5aa713c};
test_input[7264:7271] = '{32'hc2161413, 32'h42b0a781, 32'h4203b1e7, 32'hc24e6bf1, 32'hc1d72c3b, 32'h42c679f0, 32'hc2003cdc, 32'h42a71aa3};
test_weights[7264:7271] = '{32'h424ad219, 32'hbd6af278, 32'h429d4bc6, 32'hc11e3152, 32'hc1fedac5, 32'h42478a71, 32'h42875607, 32'hc2a10db0};
test_bias[908:908] = '{32'h42715fdb};
test_output[908:908] = '{32'hc4e5b878};
test_input[7272:7279] = '{32'hc2a81892, 32'hc2557de6, 32'h42b1f637, 32'h4265cc1e, 32'hc20d9f56, 32'hc1ecd8e3, 32'hc203d50d, 32'hc1a713d4};
test_weights[7272:7279] = '{32'h415ded11, 32'hc233153a, 32'h4237ac97, 32'h422d6562, 32'hc1eec73c, 32'hc208d5c5, 32'h427875cd, 32'hc25f153b};
test_bias[909:909] = '{32'h41c14b72};
test_output[909:909] = '{32'h460ccd1e};
test_input[7280:7287] = '{32'hc1e72e34, 32'h4129386b, 32'h426cd3e7, 32'hc24c5511, 32'h40cd4e1d, 32'hc1fc4f3a, 32'hc2bf8e3d, 32'h42b44414};
test_weights[7280:7287] = '{32'hc1f85503, 32'hc29ab37b, 32'hc242117b, 32'hc1b38d77, 32'hc0d54669, 32'hc26d2b24, 32'hc1c008bc, 32'h411a2946};
test_bias[910:910] = '{32'h418aa7b2};
test_output[910:910] = '{32'h45524fd6};
test_input[7288:7295] = '{32'h42c18d78, 32'h41c9cdfc, 32'h429338db, 32'hc1ce4269, 32'hc18b33c9, 32'hc08326d5, 32'h4287ce20, 32'hc1e886c8};
test_weights[7288:7295] = '{32'hc2457fa3, 32'hc2b13c00, 32'h42aa6333, 32'hc23bb61b, 32'h42340128, 32'h405a314d, 32'hc2ae7086, 32'h41fd5444};
test_bias[911:911] = '{32'h42144a78};
test_output[911:911] = '{32'hc5defb13};
test_input[7296:7303] = '{32'h42a3afb7, 32'hc03ab3f9, 32'h423fdf33, 32'h42088752, 32'hc234207f, 32'h429a2947, 32'h41e7c940, 32'hc20450d5};
test_weights[7296:7303] = '{32'h428ce9a9, 32'h42b408e6, 32'hc2a742a8, 32'hc253af09, 32'h42b1bb54, 32'hc274ccc6, 32'h4234181c, 32'h425b9f2f};
test_bias[912:912] = '{32'h42acacc0};
test_output[912:912] = '{32'hc613ca77};
test_input[7304:7311] = '{32'h4252705c, 32'hc2828bc7, 32'h423f036a, 32'hc2303612, 32'hc28c90a5, 32'hc2b1f58e, 32'h41c34d75, 32'h42967945};
test_weights[7304:7311] = '{32'hc191a657, 32'hc1a7c52f, 32'hc26eff7e, 32'h4174f956, 32'h426b62e0, 32'h4293508b, 32'h425b9926, 32'h4295b0a1};
test_bias[913:913] = '{32'h42bea0ba};
test_output[913:913] = '{32'hc5d29f3f};
test_input[7312:7319] = '{32'h42979683, 32'h41e24cda, 32'h4247143b, 32'hc21a065e, 32'hc04b804c, 32'hc1c160ac, 32'hc202df8d, 32'h41be3944};
test_weights[7312:7319] = '{32'h423ee169, 32'hc29170c3, 32'h41af90f0, 32'hc2c17011, 32'hc2b3ff3a, 32'hc2619cd1, 32'h3fa5d4a3, 32'h4141dd27};
test_bias[914:914] = '{32'hc1bb58ad};
test_output[914:914] = '{32'h4600e0c5};
test_input[7320:7327] = '{32'hc293fce4, 32'h41b9df87, 32'h420618c1, 32'h42a0e99e, 32'h429b8d49, 32'h42befed9, 32'hc2b65111, 32'hc2b1c147};
test_weights[7320:7327] = '{32'h40f23f35, 32'hc1956e9b, 32'hc28f5dca, 32'h41d474cf, 32'hc16895f6, 32'h41ce7b8e, 32'hc28db75e, 32'hc11c428d};
test_bias[915:915] = '{32'h42986873};
test_output[915:915] = '{32'h45e9a94e};
test_input[7328:7335] = '{32'h42b4d25b, 32'hc11b52a7, 32'hc21d53a9, 32'h41e8d75d, 32'h429bb745, 32'h4291eacd, 32'hc2934e1b, 32'h4271bfbd};
test_weights[7328:7335] = '{32'h421df590, 32'hc0bfb746, 32'h414b9865, 32'h41d71dad, 32'h41849429, 32'hc196af65, 32'hc21c9c0c, 32'h40fc9de1};
test_bias[916:916] = '{32'hc2a66bc1};
test_output[916:916] = '{32'h45de01f2};
test_input[7336:7343] = '{32'h42573b15, 32'h4291de23, 32'h4279a485, 32'hc09706d2, 32'hc22dac21, 32'hc203ce06, 32'hc19ed644, 32'hc1ea53fd};
test_weights[7336:7343] = '{32'h42ad90a1, 32'hc19f9abc, 32'h423d94b0, 32'hc27867a4, 32'hc2bdf783, 32'h4063860e, 32'hc1683a96, 32'hc21bdacf};
test_bias[917:917] = '{32'hc2a654d0};
test_output[917:917] = '{32'h4638aad1};
test_input[7344:7351] = '{32'h40db6dcd, 32'hc22b967a, 32'hc285d9d5, 32'h42a70fe8, 32'h41a79c34, 32'h420de8d0, 32'hc25e38c0, 32'h41874feb};
test_weights[7344:7351] = '{32'h4172a219, 32'h41ffe9c9, 32'h42153e3c, 32'hc29a67b1, 32'hc2474c42, 32'hc2b7535a, 32'h425dfe7d, 32'hc2c0d77d};
test_bias[918:918] = '{32'hc116011d};
test_output[918:918] = '{32'hc69642d9};
test_input[7352:7359] = '{32'h42a893d5, 32'h427c7ed8, 32'h42147035, 32'hc2a71fb7, 32'h429ed772, 32'hc2237f4b, 32'hc2bfeae6, 32'hc24cc4b5};
test_weights[7352:7359] = '{32'hc1955384, 32'h4206e139, 32'h42c4e9fb, 32'h42c6289e, 32'hc1cd39d7, 32'hc189d2c3, 32'h42827239, 32'hc22f17ae};
test_bias[919:919] = '{32'h429d1c2b};
test_output[919:919] = '{32'hc611fb9c};
test_input[7360:7367] = '{32'h41cbb532, 32'h428b8d6e, 32'hc2b05942, 32'hc1a1f822, 32'h4280bced, 32'h41d4145c, 32'h4290117b, 32'h3f958018};
test_weights[7360:7367] = '{32'hc26e9352, 32'h42bca4c5, 32'hc1b290a4, 32'h40819bd9, 32'hc1a13d56, 32'hc227c871, 32'hc1dea493, 32'hc297f386};
test_bias[920:920] = '{32'hc2831c51};
test_output[920:920] = '{32'h4514c6c3};
test_input[7368:7375] = '{32'hc1e3656b, 32'hc2998d8d, 32'h42885eba, 32'hc25b84e5, 32'hc0118e6c, 32'hc0f78a38, 32'hc28c5ae7, 32'hc227b34a};
test_weights[7368:7375] = '{32'h42456c3a, 32'hc290aae2, 32'h42a2a5c4, 32'h4210c83b, 32'h40d5ac90, 32'h3f58cfe5, 32'hc20865f8, 32'hc2558d1c};
test_bias[921:921] = '{32'hc259351f};
test_output[921:921] = '{32'h463fa234};
test_input[7376:7383] = '{32'h42b31fc4, 32'hc1ec8e3b, 32'h426e4173, 32'h41230ea3, 32'hc231c095, 32'h42c6f8a7, 32'hc28f288e, 32'h429fc6a6};
test_weights[7376:7383] = '{32'hc2349f0a, 32'hc267719a, 32'h41dfa7c7, 32'hc23a20ae, 32'h410b4b13, 32'hc1872ae5, 32'hc26c5b97, 32'hc2b969e9};
test_bias[922:922] = '{32'hc27dee71};
test_output[922:922] = '{32'hc5c990f2};
test_input[7384:7391] = '{32'h424a7571, 32'hc2368369, 32'h42729d9d, 32'hc29d383f, 32'hc2b61c97, 32'h3cf58927, 32'h4278c5d4, 32'h40c9c968};
test_weights[7384:7391] = '{32'hc1b4aab6, 32'hc0c8bad8, 32'h425e21b5, 32'h428f3c3e, 32'hc211fbf4, 32'h42b48146, 32'h42005a2c, 32'hc2bb5ed1};
test_bias[923:923] = '{32'hc1850330};
test_output[923:923] = '{32'h44c7782a};
test_input[7392:7399] = '{32'hbe81fbec, 32'h42077d89, 32'hc24d87ef, 32'h42ac99ba, 32'h419c605b, 32'h425b9837, 32'hc0155730, 32'hc211a72f};
test_weights[7392:7399] = '{32'hbf41cd2f, 32'h42c7e97c, 32'h41d3d2c8, 32'h4281488f, 32'hc2396ad9, 32'hc2b67184, 32'h4254dd4f, 32'h4221be28};
test_bias[924:924] = '{32'hc089426a};
test_output[924:924] = '{32'h42b24c22};
test_input[7400:7407] = '{32'h41dee8b6, 32'hc26f4b93, 32'h425c5d04, 32'h42c75cb2, 32'hc2bf5066, 32'h423c1115, 32'hc2c48e98, 32'h40dabb8b};
test_weights[7400:7407] = '{32'h42426010, 32'hc29df042, 32'h41dec61a, 32'hc23d0a67, 32'h42a639d4, 32'hc2403d6c, 32'h41ddffaa, 32'h422a630d};
test_bias[925:925] = '{32'hc0b3bb35};
test_output[925:925] = '{32'hc61858e5};
test_input[7408:7415] = '{32'h420975eb, 32'h42906f10, 32'h42a8dfda, 32'hc296ec5d, 32'h414e9fd1, 32'hc2c4f7db, 32'hc15863ad, 32'hc205cb5c};
test_weights[7408:7415] = '{32'h41872282, 32'hc2b447e6, 32'hc27b71f5, 32'h408ff8ed, 32'h40893189, 32'hc210dcd2, 32'hc2b5be0e, 32'h415d8d8e};
test_bias[926:926] = '{32'hc281bd23};
test_output[926:926] = '{32'hc5e2ac61};
test_input[7416:7423] = '{32'h4126e984, 32'hc28590a1, 32'h42540b82, 32'h420b8e28, 32'h4274454b, 32'hc223ab29, 32'h40e0a1eb, 32'h42907f32};
test_weights[7416:7423] = '{32'hc203b62c, 32'hc24bccf4, 32'h426e1a57, 32'h42b72879, 32'h416bf3db, 32'hc195530c, 32'h4297bbdb, 32'h41c9e267};
test_bias[927:927] = '{32'hc2ba3d0b};
test_output[927:927] = '{32'h465062b4};
test_input[7424:7431] = '{32'h42b4f36c, 32'h41e3d513, 32'hc13bd30c, 32'h41537c3c, 32'h42a2969e, 32'h41648391, 32'hc1d0c2de, 32'h42b6c577};
test_weights[7424:7431] = '{32'h41aeafb2, 32'hc1a00777, 32'hc27e11bb, 32'h42835b83, 32'h3feb4557, 32'hc2a5b90e, 32'h42afb74d, 32'h427488bf};
test_bias[928:928] = '{32'h42b7d97b};
test_output[928:928] = '{32'h45a7dd38};
test_input[7432:7439] = '{32'h42bd5594, 32'hc2c7b2be, 32'hc206806a, 32'hc274b912, 32'hc22fa83e, 32'h41f3d1ab, 32'hc2a2a1d7, 32'h424bf5e9};
test_weights[7432:7439] = '{32'h422b3d7b, 32'h4266e00a, 32'h420f702d, 32'h3fcd4a32, 32'h4263d76c, 32'hc28a9a01, 32'hc12166e9, 32'h418574d5};
test_bias[929:929] = '{32'hc2aff347};
test_output[929:929] = '{32'hc5bce770};
test_input[7440:7447] = '{32'h428a0112, 32'hc25eea6e, 32'h42971f6d, 32'hc2850d76, 32'h42b4d89b, 32'h42ad782c, 32'hc13c1746, 32'hc1925bfa};
test_weights[7440:7447] = '{32'hc24a9038, 32'h415597cb, 32'h42a9b808, 32'hc080623a, 32'h41f4c27a, 32'h429826b2, 32'hc15dfaa2, 32'hc25a2137};
test_bias[930:930] = '{32'h4271143f};
test_output[930:930] = '{32'h464b8a86};
test_input[7448:7455] = '{32'h4292b777, 32'hc18961f2, 32'h41cde4a8, 32'hc1d8cc6c, 32'hc2812246, 32'h42c5de88, 32'hc1eeb70e, 32'h423f6bd7};
test_weights[7448:7455] = '{32'hc26d07e6, 32'h42bbb84e, 32'h420fc79c, 32'hc2a31240, 32'h42105fd1, 32'h423a7bdf, 32'hc28f5e8e, 32'h4284ce85};
test_bias[931:931] = '{32'hc1783581};
test_output[931:931] = '{32'h4594b87a};
test_input[7456:7463] = '{32'hc19ff4d7, 32'h42af235c, 32'hc19cb559, 32'h4195bc28, 32'h426b6e1a, 32'h422e7b50, 32'hc29ed607, 32'hc25267e7};
test_weights[7456:7463] = '{32'h4238fc4a, 32'hc29edca6, 32'hc263310d, 32'hc1c0c4d0, 32'hc19663f4, 32'hc2b865da, 32'h4132f65d, 32'h41c4675f};
test_bias[932:932] = '{32'hc2b61cad};
test_output[932:932] = '{32'hc66466f7};
test_input[7464:7471] = '{32'hc18082cc, 32'hc1812a08, 32'hc2937324, 32'hc21e9171, 32'h41d77ca4, 32'hc1e0b382, 32'hc2a25184, 32'h42b3d64a};
test_weights[7464:7471] = '{32'hc286ba1b, 32'hc121a9ab, 32'h42b252f4, 32'h42802b13, 32'h4282b728, 32'h4238c83d, 32'h42a3c0b9, 32'h42c2fefa};
test_bias[933:933] = '{32'hc09429c3};
test_output[933:933] = '{32'hc5a543c0};
test_input[7472:7479] = '{32'h42523c33, 32'hc2a704c1, 32'hc24dbdf2, 32'h4118c028, 32'hc2200e22, 32'hc2257413, 32'hc2c101c6, 32'h4294a79c};
test_weights[7472:7479] = '{32'h422d9ae5, 32'hc29bef9e, 32'h42ab3466, 32'hc15cc669, 32'hc050036e, 32'hc1c9be6a, 32'h42b2ff7e, 32'hc227804b};
test_bias[934:934] = '{32'hc23bb4ba};
test_output[934:934] = '{32'hc5c6ee39};
test_input[7480:7487] = '{32'h4156aec0, 32'hc20aff7c, 32'h42b0e3c8, 32'h42b9fd3c, 32'h429974bd, 32'h42c2dc95, 32'hc10b3a0c, 32'hc0baa692};
test_weights[7480:7487] = '{32'h411f8b7c, 32'h42b29a9f, 32'hc29a556b, 32'hbfe7620f, 32'hbee4502a, 32'hc28470f6, 32'hc1f8c5f5, 32'hc0812315};
test_bias[935:935] = '{32'hc1557b0e};
test_output[935:935] = '{32'hc67c9f82};
test_input[7488:7495] = '{32'h4285d04b, 32'h4289bd01, 32'hc28244ce, 32'h3f00bc99, 32'hc2195725, 32'hc10985e8, 32'h42806f49, 32'h42658301};
test_weights[7488:7495] = '{32'hc1ebc2e5, 32'h41c6df7d, 32'h42904e77, 32'h425a4f64, 32'hc1d11060, 32'h4256d480, 32'hc2bc40a3, 32'h4236a428};
test_bias[936:936] = '{32'hc25a4da0};
test_output[936:936] = '{32'hc5f5f7cd};
test_input[7496:7503] = '{32'hc1aef2b0, 32'h40e3eeea, 32'hc227bfd5, 32'hc264af15, 32'hc2b588b7, 32'hc2b9a38c, 32'h422960e6, 32'h410b355b};
test_weights[7496:7503] = '{32'h42a11bbf, 32'hc2872d38, 32'h429bcc05, 32'hc277a4ae, 32'h423c5d1d, 32'h420757ec, 32'h4273d2d1, 32'h4295b536};
test_bias[937:937] = '{32'hc27787ee};
test_output[937:937] = '{32'hc5c23622};
test_input[7504:7511] = '{32'h42809828, 32'h42b29e40, 32'hbf67487a, 32'h3eceb776, 32'hc27c1cac, 32'hc253fca9, 32'hc258aaf1, 32'hc108d85b};
test_weights[7504:7511] = '{32'h4290cc78, 32'hc1afcf0e, 32'h40ad20b4, 32'hc2bfaef4, 32'hc23a24a7, 32'h42a0a3ca, 32'hc23c0f29, 32'hc26c4793};
test_bias[938:938] = '{32'hc29fd227};
test_output[938:938] = '{32'h45864924};
test_input[7512:7519] = '{32'hc21355b4, 32'hc2243389, 32'hc20a3c4a, 32'hc2b10aea, 32'h424ae19a, 32'hbf91a593, 32'h42b40cea, 32'h42b120ea};
test_weights[7512:7519] = '{32'hc2c08ec0, 32'h428821a2, 32'h4294e8dc, 32'hc2270256, 32'hc2ad1764, 32'hc221f992, 32'hc1425e8c, 32'h424362cd};
test_bias[939:939] = '{32'hc1688319};
test_output[939:939] = '{32'h443b5ac5};
test_input[7520:7527] = '{32'h41e42a52, 32'hc258e7f4, 32'hc28fa1cc, 32'h426bf984, 32'hc2ba59c3, 32'hc2a84be3, 32'hc27d6aa9, 32'h415389dd};
test_weights[7520:7527] = '{32'h4254c008, 32'hc2a5810f, 32'h422a52db, 32'hc2883ffd, 32'h42999cb1, 32'hc2447071, 32'hc26383ab, 32'hc130cb23};
test_bias[940:940] = '{32'hbffd62e5};
test_output[940:940] = '{32'hc4204860};
test_input[7528:7535] = '{32'h40fcbcb8, 32'hc2abc6dd, 32'hc23d46cc, 32'h42b6029a, 32'hc28bcad3, 32'hc19eeb00, 32'hc29ebed2, 32'h420122db};
test_weights[7528:7535] = '{32'h42a60bb4, 32'hc216083c, 32'hc2415f11, 32'h41e8bf58, 32'hc2ac5a75, 32'h4287ba89, 32'h42b218fa, 32'h4109c960};
test_bias[941:941] = '{32'h426a448b};
test_output[941:941] = '{32'h45d32227};
test_input[7536:7543] = '{32'hc13877c3, 32'h42684764, 32'h423b59b1, 32'hc1bd8cb3, 32'h42237672, 32'hc24e4251, 32'h427b9d85, 32'h42a2bf01};
test_weights[7536:7543] = '{32'hc2b548e7, 32'hc26d7bff, 32'h4152246a, 32'h424d50d3, 32'hc1577886, 32'h41e4285d, 32'h41e100d7, 32'hc1b7e1fd};
test_bias[942:942] = '{32'hc1e18a6d};
test_output[942:942] = '{32'hc5a10fc0};
test_input[7544:7551] = '{32'hc294609c, 32'h417e28c6, 32'hc1b26da0, 32'hc29dde1a, 32'h4225b8cf, 32'h422c3436, 32'h4273c2a3, 32'h421c513d};
test_weights[7544:7551] = '{32'hc2a24160, 32'h42712d20, 32'h4266e025, 32'hc144fbec, 32'hc095c09f, 32'h42be7e08, 32'h42a5f33b, 32'hc214b8cc};
test_bias[943:943] = '{32'hc16dad50};
test_output[943:943] = '{32'h465d30d1};
test_input[7552:7559] = '{32'h40816e69, 32'hc22d00bf, 32'h40ac2e17, 32'h4243c734, 32'hc2b61870, 32'hc26ea027, 32'h42674954, 32'h41f5c0d7};
test_weights[7552:7559] = '{32'hc281bdf8, 32'h420853f0, 32'h42754c23, 32'h41f15584, 32'h4286d0ac, 32'hc211fd1a, 32'h41a38e0b, 32'h41ca2760};
test_bias[944:944] = '{32'h422ba06d};
test_output[944:944] = '{32'hc4ec174e};
test_input[7560:7567] = '{32'hc18fd3ce, 32'hc2c64ab9, 32'h422dba6b, 32'h41e90c39, 32'h4164824d, 32'hc0936a11, 32'h420c85a3, 32'h3f381ecc};
test_weights[7560:7567] = '{32'hc2613952, 32'hc288dbe3, 32'hc25ffb9a, 32'hc248a357, 32'h4101c061, 32'h42c51063, 32'h42993815, 32'h42465aae};
test_bias[945:945] = '{32'hc281f254};
test_output[945:945] = '{32'h45c29c38};
test_input[7568:7575] = '{32'hc290b7c4, 32'hc225a99d, 32'hc0dd02bb, 32'h4185cc4a, 32'hc2913a47, 32'h3e37d49b, 32'hc2b205c3, 32'h40b66833};
test_weights[7568:7575] = '{32'h42563b4d, 32'hc178a490, 32'hc25d0df7, 32'h42bda778, 32'h4284b44b, 32'h40c4cd3c, 32'h41d5754f, 32'h41b3dc0f};
test_bias[946:946] = '{32'hc24a19c1};
test_output[946:946] = '{32'hc602ea0f};
test_input[7576:7583] = '{32'hc2a5ee73, 32'hc2b175c1, 32'hc2240a19, 32'hc174f817, 32'h4214851a, 32'h4236d70c, 32'h42833bf2, 32'h42a2ddd3};
test_weights[7576:7583] = '{32'h410465bf, 32'hc2340c4c, 32'hc2b37cbe, 32'hc29de417, 32'h425df7f0, 32'hc2a1ab0e, 32'h42926698, 32'h4224048a};
test_bias[947:947] = '{32'hbf9de3b1};
test_output[947:947] = '{32'h4665bc2b};
test_input[7584:7591] = '{32'hc254af6a, 32'hc1bceb80, 32'h40442503, 32'h42b93d01, 32'h41d55477, 32'hc276d4b1, 32'hc1b61976, 32'h42907e7f};
test_weights[7584:7591] = '{32'hc2457452, 32'h42c100da, 32'h42a9b44f, 32'hc2a5185d, 32'hc2961778, 32'h41f169b0, 32'hc250fdfe, 32'hc26c5311};
test_bias[948:948] = '{32'hbf87ecc8};
test_output[948:948] = '{32'hc65a7c7c};
test_input[7592:7599] = '{32'hc21b1df0, 32'hc211da04, 32'hc241bee5, 32'h4282c91d, 32'hc2c1b2e2, 32'hc2b2f645, 32'h420ea20a, 32'hc1580340};
test_weights[7592:7599] = '{32'hc29426dc, 32'hc2a5f530, 32'hc1c54fbb, 32'hc28ce562, 32'h42576a83, 32'h42961bac, 32'hc1e6f634, 32'hc00d3f9c};
test_bias[949:949] = '{32'hc2bbd628};
test_output[949:949] = '{32'hc624ac80};
test_input[7600:7607] = '{32'hc2048c5a, 32'h4172c7c4, 32'h42a6c035, 32'hbda29029, 32'h4205b7e4, 32'hc21b0386, 32'hc27f3a35, 32'hc2953677};
test_weights[7600:7607] = '{32'h42a0fce5, 32'hc25dc8b4, 32'hc20d298a, 32'hc1bd7303, 32'h421467f5, 32'h41e08e0c, 32'hc1d46ea7, 32'hc2afc37c};
test_bias[950:950] = '{32'hc202b546};
test_output[950:950] = '{32'h44f031d0};
test_input[7608:7615] = '{32'hc2c63918, 32'hc2bfac37, 32'h414d4c38, 32'hc2293c61, 32'h42bdcffe, 32'h41f251f5, 32'hbe488b66, 32'hc2001b13};
test_weights[7608:7615] = '{32'h42223fb7, 32'h4293c709, 32'h420f78f9, 32'h40bc9acf, 32'hc22537cd, 32'h412c4887, 32'h4288251d, 32'h427c7f50};
test_bias[951:951] = '{32'h41e2306f};
test_output[951:951] = '{32'hc680d64e};
test_input[7616:7623] = '{32'h427ca139, 32'h42b0a6fa, 32'hc29c54c8, 32'h4285072b, 32'hc21772f4, 32'hc2ba539f, 32'hc2ad6a4c, 32'h429aa73a};
test_weights[7616:7623] = '{32'h41f8e71f, 32'hc29b3cc9, 32'h4104067f, 32'h42660046, 32'hc26e94b8, 32'hc1450d08, 32'hc18c656a, 32'h410f95ae};
test_bias[952:952] = '{32'h425b0fb8};
test_output[952:952] = '{32'h4577ce0d};
test_input[7624:7631] = '{32'hc297daa0, 32'h42bb03e6, 32'h4273fb53, 32'hc275f455, 32'hc08f026b, 32'h42914842, 32'hc1cf6232, 32'hc2ad3ee3};
test_weights[7624:7631] = '{32'h4195ee07, 32'h41824d3c, 32'h427583eb, 32'h4175701b, 32'hc2263fa8, 32'h41552b90, 32'h422d7dd9, 32'hc23fe12d};
test_bias[953:953] = '{32'h42b48d9a};
test_output[953:953] = '{32'h45e03b62};
test_input[7632:7639] = '{32'hc232e583, 32'h424c199f, 32'h41897f79, 32'h420ef5fd, 32'hc25cda1a, 32'h42506d65, 32'h41ecb91f, 32'hc1e5aa28};
test_weights[7632:7639] = '{32'h410361c8, 32'h42c28c12, 32'hc2c0e2f3, 32'hc2102714, 32'h42b11d5b, 32'hc2ae4d04, 32'h422fc310, 32'hc2c1b802};
test_bias[954:954] = '{32'h417dc538};
test_output[954:954] = '{32'hc5663639};
test_input[7640:7647] = '{32'h41a61e7c, 32'h4299ae32, 32'hc1a2c6a1, 32'h411a790e, 32'h4044c6ef, 32'h41048cda, 32'hc1faef56, 32'h4186aafe};
test_weights[7640:7647] = '{32'h4294f81a, 32'hc2c50b0e, 32'hc1e3e496, 32'hc29ee6a6, 32'hc29bb6ff, 32'h4236a540, 32'h4242bd12, 32'hc2b7c43e};
test_bias[955:955] = '{32'h42561df7};
test_output[955:955] = '{32'hc60e1251};
test_input[7648:7655] = '{32'hc2b4fd88, 32'h4283839b, 32'h4249df93, 32'h428cb8ce, 32'h427271c9, 32'h423260bb, 32'hc24de741, 32'hc1bdc2bd};
test_weights[7648:7655] = '{32'h42c6eb00, 32'hc18e87a0, 32'h423bec33, 32'hc265e2dd, 32'hc26515ab, 32'h42bd6f71, 32'h41d0f044, 32'h42189cb1};
test_bias[956:956] = '{32'hc29043fe};
test_output[956:956] = '{32'hc65196f5};
test_input[7656:7663] = '{32'h42a3bd8e, 32'h42b29d26, 32'hc29c417d, 32'hc20c507f, 32'hc1b64922, 32'h41e69c46, 32'h42b36f9c, 32'hc29d8bdc};
test_weights[7656:7663] = '{32'hc25fd614, 32'hc2c651c4, 32'hc203c0be, 32'h42a6f5ed, 32'h42b87c3b, 32'h42147176, 32'h4290692a, 32'hc202ed73};
test_bias[957:957] = '{32'h42c70cc0};
test_output[957:957] = '{32'hc5b1201d};
test_input[7664:7671] = '{32'h425cd0f5, 32'hc1e4f88f, 32'hc28b7d8d, 32'h42052622, 32'h3e6ed757, 32'h428b432f, 32'hc2a1ed0b, 32'hc28efd95};
test_weights[7664:7671] = '{32'hc28b2015, 32'h41356339, 32'h420a4b5c, 32'h410ba91b, 32'hc12ff884, 32'hc06df46e, 32'hc26d544f, 32'hc1cd5173};
test_bias[958:958] = '{32'h429885fd};
test_output[958:958] = '{32'h43280981};
test_input[7672:7679] = '{32'h42886b42, 32'hc270fcf3, 32'h42be99dd, 32'hc281ca7e, 32'hc294a988, 32'hc28b9f3e, 32'hc1ab102a, 32'h42b3ade6};
test_weights[7672:7679] = '{32'hc277522b, 32'hc1ac5e35, 32'h42a4489f, 32'hc22658bd, 32'h4272dbf8, 32'h406f7750, 32'hc123f829, 32'hc28c8900};
test_bias[959:959] = '{32'hc2b4d3a0};
test_output[959:959] = '{32'hc5516af2};
test_input[7680:7687] = '{32'hc22bcdda, 32'hc20ee8a2, 32'h42aa6a93, 32'hc255e9e1, 32'h423a581b, 32'h4265a0df, 32'h42c628ef, 32'hc2076243};
test_weights[7680:7687] = '{32'hc1d7b841, 32'h429c6b97, 32'h410f0777, 32'hc16432ac, 32'hc2b98f82, 32'hc295822d, 32'hc03aa295, 32'hc17d2435};
test_bias[960:960] = '{32'h42abb68b};
test_output[960:960] = '{32'hc603239d};
test_input[7688:7695] = '{32'hc2b783c9, 32'hc1dc653c, 32'hc1c4d294, 32'h41d36f6d, 32'h422e391b, 32'hc1c679a3, 32'h4012644a, 32'h418b3335};
test_weights[7688:7695] = '{32'hc228f1ca, 32'h41e72acf, 32'hc12a87f6, 32'hc2a9f467, 32'h3fef5655, 32'hc249583b, 32'h415b2ce3, 32'hc2227805};
test_bias[961:961] = '{32'hc1cb98ed};
test_output[961:961] = '{32'h44d7a40e};
test_input[7696:7703] = '{32'h42a9c9f7, 32'h41d09977, 32'h4286796f, 32'h4294a0b4, 32'h42991771, 32'hc2801718, 32'hc1e3fbcd, 32'hc2874a09};
test_weights[7696:7703] = '{32'h41e0f4a3, 32'hc23788fa, 32'h429228c1, 32'h42463000, 32'h42394eb7, 32'hc22782ae, 32'h41d96071, 32'hc2a65bbd};
test_bias[962:962] = '{32'hc1a4a1e9};
test_output[962:962] = '{32'h46a2dcaa};
test_input[7704:7711] = '{32'h428c916f, 32'h42860dc4, 32'hc2af2452, 32'h4197a80b, 32'hc2c5f6f0, 32'hc24076f2, 32'hc271e18d, 32'h429702c4};
test_weights[7704:7711] = '{32'h4248d2b5, 32'h428a5d86, 32'hc29befa0, 32'hc1e41774, 32'h420618fb, 32'hc1a64672, 32'hc1cbcd85, 32'hc2b26fa0};
test_bias[963:963] = '{32'h4224ba88};
test_output[963:963] = '{32'h45da1fe5};
test_input[7712:7719] = '{32'hc223a928, 32'h40d9e973, 32'h41fe8e10, 32'hc28a9817, 32'h42643c3b, 32'h42bc5738, 32'h41b0fe16, 32'hc21fcbfb};
test_weights[7712:7719] = '{32'hc0892d55, 32'h41d8ecf7, 32'h41eddf55, 32'h4252cc68, 32'hc1c069b2, 32'h42485db5, 32'h42ac0559, 32'hc1b95bf5};
test_bias[964:964] = '{32'h41733574};
test_output[964:964] = '{32'h45702bc6};
test_input[7720:7727] = '{32'h42c149d5, 32'h40bca3d4, 32'h42b56f45, 32'h42b8e69b, 32'h42b1840a, 32'h42b01949, 32'hc25fcbdc, 32'hc0618a45};
test_weights[7720:7727] = '{32'h40eb4f79, 32'h42a0f21e, 32'hc29a3200, 32'hc1c33556, 32'h42afd7c2, 32'h4257f9f1, 32'h4234052c, 32'hc27e9e3a};
test_bias[965:965] = '{32'h42a40ee3};
test_output[965:965] = '{32'h450e94d3};
test_input[7728:7735] = '{32'hc2686aeb, 32'hc21dfcb8, 32'h42a49331, 32'hc210a671, 32'hc1a80b44, 32'h420a0485, 32'hc29558ba, 32'hc20f3ec9};
test_weights[7728:7735] = '{32'h4187b8e3, 32'h4286639b, 32'hc1b4b5f8, 32'hc28fe4a9, 32'hc14adb55, 32'hc20bc68d, 32'hc1ecc5e7, 32'h41f7b49c};
test_bias[966:966] = '{32'hc1a5ecff};
test_output[966:966] = '{32'hc52c3a0f};
test_input[7736:7743] = '{32'h41db3366, 32'h424a6177, 32'hc2c4ba11, 32'hc14efe5d, 32'hc0906cdf, 32'h42545151, 32'hc250d623, 32'hc0d88bb1};
test_weights[7736:7743] = '{32'hc2a52c0b, 32'hc296318a, 32'hc28055bb, 32'hc12f2eeb, 32'h4191e03e, 32'hc28e60df, 32'hc19d50a3, 32'h426a4b7a};
test_bias[967:967] = '{32'h423e46be};
test_output[967:967] = '{32'hc52e824d};
test_input[7744:7751] = '{32'h421a2dfe, 32'hc2af324e, 32'h41d41501, 32'hc184b3a0, 32'h41a1e4b2, 32'hc2bd9721, 32'h4103c2de, 32'hc2c6c81d};
test_weights[7744:7751] = '{32'h421208a2, 32'hc10d75dd, 32'h424ab6dd, 32'h41a78249, 32'hc16c8298, 32'hc292853b, 32'h4270122f, 32'hc1af6932};
test_bias[968:968] = '{32'hc07cd70f};
test_output[968:968] = '{32'h46433421};
test_input[7752:7759] = '{32'h4038661c, 32'h42719131, 32'hc2b5f03a, 32'hc2ab45a0, 32'hc295f33b, 32'hc2b78faa, 32'hc2152450, 32'hc2a12c28};
test_weights[7752:7759] = '{32'h415abc96, 32'hc22bb0ba, 32'hc2747b78, 32'h411216ae, 32'hc2b370c3, 32'hc23b4308, 32'h41e734c6, 32'h429548da};
test_bias[969:969] = '{32'hc21973db};
test_output[969:969] = '{32'h45bf2ed1};
test_input[7760:7767] = '{32'h42c4d562, 32'hc1c9aea1, 32'h42c6ae21, 32'h410a1629, 32'hc2b5584c, 32'h407038f4, 32'hc23d41d2, 32'hc1a71944};
test_weights[7760:7767] = '{32'h412ca15c, 32'hc165df23, 32'h42a5244e, 32'h425c078c, 32'h42893ab2, 32'h41b04a4c, 32'hc289a4b3, 32'h42ad8496};
test_bias[970:970] = '{32'hc1424c02};
test_output[970:970] = '{32'h45a894b2};
test_input[7768:7775] = '{32'hc18f1057, 32'hc1c07182, 32'hc237284b, 32'hc0fad65e, 32'hc253dcc9, 32'h4211e849, 32'hc266e6eb, 32'h41cc18ba};
test_weights[7768:7775] = '{32'h42634fb6, 32'hc24e44c9, 32'h41940b80, 32'hc24fafa0, 32'hc23c909c, 32'h41b39ca7, 32'h4291a615, 32'hc1e67ba1};
test_bias[971:971] = '{32'h4208f812};
test_output[971:971] = '{32'hc4e19d55};
test_input[7776:7783] = '{32'hc07c724b, 32'h420814c4, 32'h423c189c, 32'h42a3b8ae, 32'h42190f40, 32'h41dae29b, 32'h42bbf8ca, 32'hc20eaadb};
test_weights[7776:7783] = '{32'h41f00238, 32'hbf8f9874, 32'h4226eade, 32'hc2963c7f, 32'hc25065ba, 32'hc2734006, 32'hc27ef90c, 32'h42986467};
test_bias[972:972] = '{32'hc1bf26cc};
test_output[972:972] = '{32'hc682bad9};
test_input[7784:7791] = '{32'hc29d5dec, 32'h41b1d02d, 32'hc21518d3, 32'h42b0d9ca, 32'hc2a3a9c8, 32'h41fbafb5, 32'h42b30d3a, 32'hc1bf132d};
test_weights[7784:7791] = '{32'h425fd486, 32'hc28b0f74, 32'h4291494e, 32'h42855cfb, 32'h4227a16a, 32'h408a307e, 32'h423b25e9, 32'h427cbb18};
test_bias[973:973] = '{32'hc248dd57};
test_output[973:973] = '{32'hc555fe26};
test_input[7792:7799] = '{32'h420e9886, 32'h41b35c52, 32'h41f2895f, 32'hc1b4600e, 32'hc28d194d, 32'h41dbda94, 32'hc274c497, 32'hc2af5835};
test_weights[7792:7799] = '{32'h41a64f87, 32'hc001ec61, 32'h4220d0f4, 32'hc2810c38, 32'h41bf9e20, 32'hc211df04, 32'h424fd0c4, 32'h4281874c};
test_bias[974:974] = '{32'hc1f5609c};
test_output[974:974] = '{32'hc6004a6c};
test_input[7800:7807] = '{32'hc0fccf58, 32'h428e9c33, 32'h41bff7df, 32'hc2957a6b, 32'h42557ae6, 32'hc03edaf8, 32'h422a8e26, 32'h41bc61f1};
test_weights[7800:7807] = '{32'h42b10f20, 32'h41f04727, 32'h42043689, 32'h425e1b8f, 32'hc22a1ee2, 32'h42ba4f28, 32'h4177b9df, 32'hc273ab75};
test_bias[975:975] = '{32'hc23d70a2};
test_output[975:975] = '{32'hc5a51fae};
test_input[7808:7815] = '{32'hc1bf394d, 32'hc2b7d497, 32'hc0b13be7, 32'hbead65f8, 32'hc276d503, 32'hc27224d7, 32'h42aa4e12, 32'h426f0548};
test_weights[7808:7815] = '{32'h4107e555, 32'h42481b93, 32'h41606a57, 32'hc22c3198, 32'hc2c4fd49, 32'h42c0646c, 32'hc2396aeb, 32'h42aafe01};
test_bias[976:976] = '{32'hc2427247};
test_output[976:976] = '{32'hc55a8bf2};
test_input[7816:7823] = '{32'h42b90e0e, 32'h423f10aa, 32'h420b6e61, 32'hbf876e91, 32'hc2c6c6e9, 32'hbed79215, 32'hbf1c5eae, 32'h4247e576};
test_weights[7816:7823] = '{32'hc286f150, 32'h42a8c8be, 32'h429cd79e, 32'hc1cb0cc5, 32'hc280c8ec, 32'h41032829, 32'h427f3a7b, 32'h42097632};
test_bias[977:977] = '{32'hc2987d0f};
test_output[977:977] = '{32'h46058caa};
test_input[7824:7831] = '{32'hc22fc929, 32'hc2372887, 32'hc1926e60, 32'hc031a979, 32'hc27c4174, 32'hc2b133a0, 32'hc27a09df, 32'hc23a9a62};
test_weights[7824:7831] = '{32'h42b2fc42, 32'h429377fd, 32'hc23cc25f, 32'h41bce2df, 32'h42c77b04, 32'hc2245242, 32'hc2c56fe0, 32'h42164715};
test_bias[978:978] = '{32'hc23ec028};
test_output[978:978] = '{32'hc595b558};
test_input[7832:7839] = '{32'hc29b83f3, 32'hc2608d56, 32'h42557ca1, 32'h41e01fa8, 32'h4140d77d, 32'hc2901e3b, 32'h4111933d, 32'h4192958c};
test_weights[7832:7839] = '{32'hc26a7447, 32'h42bcc543, 32'hc2ab8e90, 32'hc22034c3, 32'hc2a3628e, 32'h4206e042, 32'hc2584115, 32'hc23add45};
test_bias[979:979] = '{32'h420a188d};
test_output[979:979] = '{32'hc62e8378};
test_input[7840:7847] = '{32'hc1edba03, 32'hc256828b, 32'hc28bcd48, 32'hc11ed2fd, 32'hc25cb5a1, 32'hc218de25, 32'h4193f82a, 32'h42bd445a};
test_weights[7840:7847] = '{32'hc05c4a5f, 32'h41f71a00, 32'hc274abc9, 32'h42b282f2, 32'h42807941, 32'h42b6f6ef, 32'hc28ff6cd, 32'h42b8b517};
test_bias[980:980] = '{32'hc2c58436};
test_output[980:980] = '{32'h450388cc};
test_input[7848:7855] = '{32'h429911ec, 32'h4275fe4e, 32'h41467ffd, 32'h415495d8, 32'h4251df8d, 32'h41250be5, 32'h42a35154, 32'h411c3b0a};
test_weights[7848:7855] = '{32'h41be401c, 32'h421f8ac4, 32'hc023b935, 32'h428f0a60, 32'h41291503, 32'hc2015be1, 32'hc1af3e63, 32'hc204b234};
test_bias[981:981] = '{32'hc157f290};
test_output[981:981] = '{32'h454d6309};
test_input[7856:7863] = '{32'h4285db99, 32'hc2b31d86, 32'h4296d69a, 32'hc27d0322, 32'h41aa7df6, 32'h4267c21b, 32'hc217e329, 32'h42376f86};
test_weights[7856:7863] = '{32'h4232b798, 32'hc29538af, 32'h41f9f4e7, 32'hc24706a8, 32'hc1925efb, 32'hc2054e33, 32'hc2a76682, 32'hc2aa6ce4};
test_bias[982:982] = '{32'h420f9081};
test_output[982:982] = '{32'h463e061f};
test_input[7864:7871] = '{32'hc171a3a7, 32'h41dff7d0, 32'hc2842a7b, 32'h4238bada, 32'hc1f34c61, 32'h428cf6f9, 32'hc29587a5, 32'hc2967634};
test_weights[7864:7871] = '{32'hc23200f2, 32'hc0ea608c, 32'hc2b25068, 32'hc2a5fe8b, 32'hc1fd716e, 32'hc230ce39, 32'hc18746f5, 32'hc22c95af};
test_bias[983:983] = '{32'h4180abd7};
test_output[983:983] = '{32'h459920a9};
test_input[7872:7879] = '{32'hc1a0d0eb, 32'hc2afde9c, 32'hc2bccc2e, 32'h40ea021e, 32'h42af2fce, 32'h4245c4d3, 32'h42923889, 32'h42c36384};
test_weights[7872:7879] = '{32'h419d6fa3, 32'h40f96035, 32'h428f6fde, 32'h429d919d, 32'h4267317c, 32'hc260b9d1, 32'h4263be75, 32'h4294b839};
test_bias[984:984] = '{32'hc2b7bc05};
test_output[984:984] = '{32'h45c64b53};
test_input[7880:7887] = '{32'h42c6929e, 32'hc2853a4d, 32'h42396781, 32'hc2135409, 32'h41cbc0f7, 32'h429b1af9, 32'h4299ffcc, 32'h42570261};
test_weights[7880:7887] = '{32'h416d6b92, 32'h4267e5d9, 32'hc23d48b4, 32'h411bbeae, 32'h42788a60, 32'hc0400b96, 32'h42358532, 32'h4240ce1e};
test_bias[985:985] = '{32'hc23d01f9};
test_output[985:985] = '{32'h4518f39f};
test_input[7888:7895] = '{32'h4218b7fb, 32'hc2bd53de, 32'hc22ed4ec, 32'hc1801c7a, 32'hc0d4ea22, 32'h42abc28e, 32'hc1fd4267, 32'hc2750762};
test_weights[7888:7895] = '{32'h421fdcdb, 32'h42997b81, 32'hc1a0e697, 32'hc2a448eb, 32'h4177f049, 32'hc29bccbb, 32'hc252639a, 32'hc10542ba};
test_bias[986:986] = '{32'hc2bc0afc};
test_output[986:986] = '{32'hc6010073};
test_input[7896:7903] = '{32'h425318f4, 32'hc11c4b94, 32'h42572d78, 32'h4188f5e4, 32'hc26acc29, 32'h42a83ee5, 32'hc1e7411d, 32'h420fe149};
test_weights[7896:7903] = '{32'hc2112572, 32'h42c11ce5, 32'hc2ab5466, 32'h42372a43, 32'h41bbfffb, 32'hc22bde70, 32'hc2960c1e, 32'h429fd2f7};
test_bias[987:987] = '{32'hc1618073};
test_output[987:987] = '{32'hc5cfbbc4};
test_input[7904:7911] = '{32'h42a06047, 32'h42c7d0cb, 32'h41113e63, 32'hc2543b65, 32'hc1733b53, 32'hc2b34dcc, 32'h42b2bb8a, 32'hc0c086b0};
test_weights[7904:7911] = '{32'h4260b248, 32'hc2110594, 32'hc2a55561, 32'hc282fdf5, 32'h42960d4b, 32'hc21c210e, 32'h42c715c4, 32'hc2ba4417};
test_bias[988:988] = '{32'hc2717224};
test_output[988:988] = '{32'h467005c1};
test_input[7912:7919] = '{32'h404e1918, 32'h428a7242, 32'h42aa6e01, 32'h42bc5560, 32'h411bdc9d, 32'h42bb621c, 32'h4249de49, 32'h41657860};
test_weights[7912:7919] = '{32'hc21ad912, 32'h42c68bd5, 32'h4232000e, 32'hc222a894, 32'h4245aca6, 32'hc2bafbeb, 32'hc2b33610, 32'h4245cbb5};
test_bias[989:989] = '{32'hc13a19a5};
test_output[989:989] = '{32'hc5a8838c};
test_input[7920:7927] = '{32'h4114a3f2, 32'h4208afe6, 32'hc255941f, 32'h426c53e3, 32'hc130f31e, 32'h427f3923, 32'hc21bed45, 32'h42233115};
test_weights[7920:7927] = '{32'h41ffb7e2, 32'h42934460, 32'h41a5c525, 32'hc1d4a5aa, 32'h41bbfd8f, 32'h428e1fd5, 32'h42072457, 32'hc2ac6c1b};
test_bias[990:990] = '{32'hc0e09dcb};
test_output[990:990] = '{32'hc3d757f6};
test_input[7928:7935] = '{32'h4291d467, 32'hc256ddf4, 32'hc2bcfea1, 32'h42629eae, 32'h428ee187, 32'hc28212d4, 32'h422b3219, 32'h42b6527c};
test_weights[7928:7935] = '{32'h41f29a49, 32'h4289e1eb, 32'h4277c83b, 32'h428d552d, 32'hc2c6a76b, 32'hc27fb8a1, 32'hc0dcd643, 32'hc2b27be4};
test_bias[991:991] = '{32'hc0c79068};
test_output[991:991] = '{32'hc665f573};
test_input[7936:7943] = '{32'hc2a75111, 32'hc2b405b8, 32'hc28a2e2c, 32'h41a32027, 32'h422cf238, 32'hc0cfc318, 32'h425f8600, 32'h420838b8};
test_weights[7936:7943] = '{32'hc2517118, 32'hc24a397f, 32'h41c395d0, 32'hc282584d, 32'hc2c47e8d, 32'h425b6f13, 32'h41ae7388, 32'h42542380};
test_bias[992:992] = '{32'hc25d36ce};
test_output[992:992] = '{32'h4585b265};
test_input[7944:7951] = '{32'h42bbef22, 32'hc2aac7bf, 32'hc23c2651, 32'h42c05ad0, 32'hc0dc76dc, 32'h4183e86c, 32'hc2225b51, 32'h4282fc49};
test_weights[7944:7951] = '{32'hc20dd45d, 32'h429873d3, 32'hc290ecaa, 32'h42a54fe6, 32'h4298a8e6, 32'h422db38d, 32'hc26f000b, 32'h4260d59f};
test_bias[993:993] = '{32'hc2be9909};
test_output[993:993] = '{32'h45f134b9};
test_input[7952:7959] = '{32'hc191751a, 32'hc2b2ae72, 32'hc0efc35f, 32'h41bae5a5, 32'h4121aef4, 32'hc21cc952, 32'hc243f56a, 32'hc26d40f2};
test_weights[7952:7959] = '{32'h41df58bc, 32'h4288f798, 32'hc12f8de6, 32'h42843d72, 32'h424bd39e, 32'hc0fe4a22, 32'hc2355ba8, 32'h42c37745};
test_bias[994:994] = '{32'h41ee4abb};
test_output[994:994] = '{32'hc5f134b9};
test_input[7960:7967] = '{32'h418619da, 32'h42746468, 32'h425d94ca, 32'h42029a7e, 32'hc191fe46, 32'h428b73bc, 32'h426d496e, 32'h427a5d74};
test_weights[7960:7967] = '{32'hc28bae08, 32'h42789384, 32'hc23edab1, 32'hc11b270f, 32'hc2151fdc, 32'h41e1af89, 32'hc03f21d0, 32'h4216894c};
test_bias[995:995] = '{32'h42baf650};
test_output[995:995] = '{32'h458f4db2};
test_input[7968:7975] = '{32'hc1228b05, 32'h42918873, 32'hc2b940ff, 32'hc22de53b, 32'h426e095f, 32'h41e42591, 32'hc2bed46a, 32'h4196f1ea};
test_weights[7968:7975] = '{32'hc1289909, 32'hc060fbda, 32'h42bc6ff9, 32'hc159a1c2, 32'hc22184cb, 32'h418a3fbc, 32'h41b266c1, 32'hc297f478};
test_bias[996:996] = '{32'hc233cbbd};
test_output[996:996] = '{32'hc657a40e};
test_input[7976:7983] = '{32'hc15259ea, 32'h42830a32, 32'h423f3e46, 32'h411ab05c, 32'hc095c51e, 32'hc25559e2, 32'hc205f1b7, 32'h40d92050};
test_weights[7976:7983] = '{32'h41f12725, 32'hc2442990, 32'hc1e213c6, 32'h4106b4ba, 32'hbfd9255d, 32'h42733360, 32'hc298492d, 32'h42868de0};
test_bias[997:997] = '{32'hc283874d};
test_output[997:997] = '{32'hc5a1adb9};
test_input[7984:7991] = '{32'hc2bb7d43, 32'hc2b287da, 32'h42971263, 32'hc2c6c244, 32'h41fd1831, 32'h41d3a6bb, 32'h4215ebe0, 32'hc2abbbf9};
test_weights[7984:7991] = '{32'hc22f5e51, 32'hc28e6ca1, 32'hc23a7ea1, 32'h428e08d4, 32'h42c3568a, 32'h424b3e8b, 32'hc1baf40c, 32'h424a3e34};
test_bias[998:998] = '{32'h4267d26a};
test_output[998:998] = '{32'hc4517922};
test_input[7992:7999] = '{32'hc28dc186, 32'h4104af3f, 32'hc210d303, 32'h41157b22, 32'hc26f5f59, 32'hc251b763, 32'h41f4e375, 32'hc22aa4ae};
test_weights[7992:7999] = '{32'h41c6df5c, 32'hc2afc41e, 32'hc1564953, 32'h42bf804b, 32'h428abbbd, 32'hc2431760, 32'h41c48102, 32'h42a2765d};
test_bias[999:999] = '{32'h4289297d};
test_output[999:999] = '{32'hc5a731a7};
test_input[8000:8007] = '{32'h40ed1a06, 32'hc2131e21, 32'h42839b5d, 32'h4181617b, 32'h42a416e7, 32'h4228c0be, 32'hc243b800, 32'h42aad3e7};
test_weights[8000:8007] = '{32'hc21a4b61, 32'hc29c5103, 32'h420fb9bc, 32'hc03ab6bf, 32'h4254f8d7, 32'h41e8e694, 32'hc250dc3f, 32'h41e4e9c1};
test_bias[1000:1000] = '{32'h42a65df5};
test_output[1000:1000] = '{32'h46738294};
test_input[8008:8015] = '{32'hc099ef9f, 32'hc29ffe80, 32'h4232cc52, 32'h40f4139d, 32'h4296b862, 32'h413185bc, 32'hc23a5716, 32'h423f111e};
test_weights[8008:8015] = '{32'hc227dee1, 32'hc21703c8, 32'h428688a0, 32'h42925543, 32'h42a78131, 32'h41a3f81e, 32'hc208cc45, 32'h4240ee45};
test_bias[1001:1001] = '{32'h4249dcfd};
test_output[1001:1001] = '{32'h4686f2ff};
test_input[8016:8023] = '{32'hc2ba5a44, 32'hc1f229ce, 32'h42af8917, 32'hc2b875a7, 32'hc066fe68, 32'h420b08f0, 32'hc27f94a4, 32'hc21cc19a};
test_weights[8016:8023] = '{32'h424d0133, 32'h420577db, 32'h42074c22, 32'h42730c73, 32'h42b0b6ec, 32'h420f493c, 32'h42a3a0ab, 32'hc20d137c};
test_bias[1002:1002] = '{32'h41e2677b};
test_output[1002:1002] = '{32'hc630bea7};
test_input[8024:8031] = '{32'h415d724f, 32'hc12d7192, 32'hbfd88f61, 32'h40d86701, 32'h42679391, 32'hc22c6e1a, 32'h42b6765b, 32'hc2985ae3};
test_weights[8024:8031] = '{32'h41ab71e4, 32'hc27fd564, 32'h40b5c9a0, 32'h42585e4b, 32'hc22ecbbf, 32'hc26550a9, 32'h41c16a99, 32'hc190e0e8};
test_bias[1003:1003] = '{32'hbf8671a6};
test_output[1003:1003] = '{32'h45983dc5};
test_input[8032:8039] = '{32'hc2461194, 32'h416b9512, 32'hc10173f8, 32'hbfe6b2d8, 32'hc127815d, 32'h42436131, 32'h426d7d72, 32'h41affeec};
test_weights[8032:8039] = '{32'hc26a86ce, 32'h41a73594, 32'h4065b08b, 32'h42b511c2, 32'hc1f6254b, 32'h4296ef7d, 32'h42a071a2, 32'h4227c1cb};
test_bias[1004:1004] = '{32'hc22a3c17};
test_output[1004:1004] = '{32'h4645f8cc};
test_input[8040:8047] = '{32'h3f96153a, 32'h423bf9e3, 32'hc23b038a, 32'h428d112c, 32'h421d9f2a, 32'hc10061f3, 32'hc1c76b65, 32'h42a91798};
test_weights[8040:8047] = '{32'hc2a5e4cf, 32'h425e8bf7, 32'hc1876845, 32'h419f948d, 32'hc28195e5, 32'h428d4fcc, 32'h429bc0bc, 32'h42b990a7};
test_bias[1005:1005] = '{32'hc2a17e66};
test_output[1005:1005] = '{32'h45e7cf5a};
test_input[8048:8055] = '{32'hc2a1632a, 32'h4290cde5, 32'h42c2cfcd, 32'h41a466aa, 32'h4257fd92, 32'hc1ce7658, 32'h4292f655, 32'h42479f36};
test_weights[8048:8055] = '{32'hc248c0db, 32'h42bc0eba, 32'h4209e104, 32'hc121bdf1, 32'h429df732, 32'h4107707f, 32'hc2a5546a, 32'h41eb1b8d};
test_bias[1006:1006] = '{32'h4259f5db};
test_output[1006:1006] = '{32'h4652f353};
test_input[8056:8063] = '{32'hc21e9285, 32'hc1a40c97, 32'hc29716f8, 32'hc04639c6, 32'h41f70d8f, 32'h3cc53833, 32'h41b8f071, 32'h41e8b617};
test_weights[8056:8063] = '{32'h3e1c48e3, 32'hc22b47e9, 32'h4023828a, 32'hc1aaad96, 32'hc23420bd, 32'hbf9c4e2d, 32'hc2919e9e, 32'hc2a66d13};
test_bias[1007:1007] = '{32'h41339c31};
test_output[1007:1007] = '{32'hc59410e6};
test_input[8064:8071] = '{32'hc1897113, 32'h427fa310, 32'h428f6033, 32'hc28f144e, 32'hc292cfac, 32'h41fba9dd, 32'hc2b21e47, 32'h421b7a09};
test_weights[8064:8071] = '{32'h42b415d3, 32'hc246da76, 32'hc288f2be, 32'hc29eeb56, 32'h421937fd, 32'hc28faf5c, 32'hc2c4a2eb, 32'hc187f0ef};
test_bias[1008:1008] = '{32'h423e408f};
test_output[1008:1008] = '{32'hc45b3b8a};
test_input[8072:8079] = '{32'hc29803c5, 32'h427e7b46, 32'h42414512, 32'h423fcb53, 32'hc2c303ff, 32'hc21d3515, 32'h427b49aa, 32'hc2853a5e};
test_weights[8072:8079] = '{32'hc058fecf, 32'hc2ad7063, 32'h4110f4f8, 32'hc22887a9, 32'h41a1115d, 32'h420de822, 32'hbf5769ae, 32'hc08bef8d};
test_bias[1009:1009] = '{32'h42832eef};
test_output[1009:1009] = '{32'hc61a9d38};
test_input[8080:8087] = '{32'hc20eb086, 32'h41198f67, 32'h42a1d2e7, 32'hc151e6cb, 32'hc28e58e8, 32'h427009f9, 32'h414cc545, 32'h428b84e3};
test_weights[8080:8087] = '{32'h424ce425, 32'h427957e5, 32'hc24e447f, 32'h41b89e61, 32'h42825c63, 32'hc168f9dc, 32'hc2230a1f, 32'hc16b227c};
test_bias[1010:1010] = '{32'h42559e21};
test_output[1010:1010] = '{32'hc64699d1};
test_input[8088:8095] = '{32'hc27cccfc, 32'h422183db, 32'h40f9e680, 32'h4062b350, 32'h421ba0bc, 32'h42b1eaae, 32'h42c552a2, 32'h420ae1dc};
test_weights[8088:8095] = '{32'h41c6460c, 32'h41d54854, 32'hc2b77491, 32'h42a91845, 32'hc28130ba, 32'h4280b2c2, 32'hc1c52d5d, 32'hc1952ef9};
test_bias[1011:1011] = '{32'hc258d981};
test_output[1011:1011] = '{32'hc44f3ad7};
test_input[8096:8103] = '{32'h425d3780, 32'h42ae0dac, 32'h42a56e66, 32'hc24a227f, 32'h4244138e, 32'h426c7904, 32'h42741134, 32'h423c5ead};
test_weights[8096:8103] = '{32'hc1ec20b9, 32'h421fc3c9, 32'hc28f466b, 32'hbfbd84fc, 32'h4161bb45, 32'h42aaff06, 32'h4206d25b, 32'h420e6c19};
test_bias[1012:1012] = '{32'hc284c226};
test_output[1012:1012] = '{32'h45a8ef40};
test_input[8104:8111] = '{32'h41f89ec4, 32'h42902e1c, 32'hc2a8fe75, 32'h4144a383, 32'h427b8d01, 32'hc2afda5e, 32'h42872d70, 32'h41a753f8};
test_weights[8104:8111] = '{32'h41886bd6, 32'hc1e9b9a2, 32'hc0d4e4c1, 32'hc2b17dd8, 32'hc25cb417, 32'h42902afd, 32'h41772c61, 32'hc227acc7};
test_bias[1013:1013] = '{32'hc1fbebea};
test_output[1013:1013] = '{32'hc6380354};
test_input[8112:8119] = '{32'hc1ad52a4, 32'h41d03d68, 32'h41640377, 32'hc1075cda, 32'h41212b8e, 32'h42a48d12, 32'hc0982470, 32'h425872b3};
test_weights[8112:8119] = '{32'hc232bcc6, 32'h4123e420, 32'h42225e03, 32'h42043d2a, 32'h4257921e, 32'hc2a6b536, 32'hc1dbae9c, 32'hc24866cd};
test_bias[1014:1014] = '{32'h41b172e2};
test_output[1014:1014] = '{32'hc5e55f3d};
test_input[8120:8127] = '{32'hc20696c7, 32'hc23db15b, 32'hc0a1a6a6, 32'hc27bf3b2, 32'h42a8da3a, 32'hc10b61cc, 32'hc20980ba, 32'hc29d23b9};
test_weights[8120:8127] = '{32'hc2a51eca, 32'h42c1a5ce, 32'hc2b7b496, 32'h42b67e5b, 32'h42962337, 32'hc23bcf36, 32'h417282fe, 32'hc25b37fa};
test_bias[1015:1015] = '{32'h4287d183};
test_output[1015:1015] = '{32'h455ae6fc};
test_input[8128:8135] = '{32'h419c84d4, 32'hc28bdd5e, 32'h41943e70, 32'h405aa0d5, 32'hc269be16, 32'hc288833e, 32'hc211d31f, 32'hc1db0d6e};
test_weights[8128:8135] = '{32'h41a1b906, 32'hc1b2ec53, 32'h421838e2, 32'hc2bac0be, 32'hc1855f94, 32'hc2b4dad3, 32'h42421efb, 32'h42313a09};
test_bias[1016:1016] = '{32'hc2bc469d};
test_output[1016:1016] = '{32'h45c87d8b};
test_input[8136:8143] = '{32'h41d06935, 32'h418f620f, 32'h42c65d2a, 32'hc1af5fb4, 32'h4215582f, 32'hc2bebf2b, 32'h42116f57, 32'hc2465b42};
test_weights[8136:8143] = '{32'hc2c2f9cf, 32'hc266fddd, 32'hc24757d6, 32'hc15e94c7, 32'hc11257a9, 32'hc276f7a9, 32'h41405c43, 32'hc29ef242};
test_bias[1017:1017] = '{32'hc253b04b};
test_output[1017:1017] = '{32'h44cf761d};
test_input[8144:8151] = '{32'hc28039f9, 32'hc276b163, 32'h42475be8, 32'h41d53253, 32'hc2be7517, 32'hc0828646, 32'hc02a372b, 32'hc28c7be6};
test_weights[8144:8151] = '{32'hc1dc3b86, 32'hc2886ec0, 32'hc172e8bb, 32'h4268de24, 32'h424d0e8b, 32'hc0796a6c, 32'h42684386, 32'h420e3581};
test_bias[1018:1018] = '{32'hc25a7fcb};
test_output[1018:1018] = '{32'hc449566a};
test_input[8152:8159] = '{32'h4284fdf3, 32'hc2908b98, 32'hc29c2b8f, 32'h42b24942, 32'hc26449df, 32'hc27efb44, 32'h422c30c5, 32'h41e660fb};
test_weights[8152:8159] = '{32'hc2b626c5, 32'h4296ba9d, 32'hc2439c08, 32'h42957854, 32'h42bb9d25, 32'h41fdb8f4, 32'hc21f62f6, 32'h4226043e};
test_bias[1019:1019] = '{32'h42850ec0};
test_output[1019:1019] = '{32'hc60a4d58};
test_input[8160:8167] = '{32'hc23e5032, 32'hc1591dcb, 32'hc0ce06b3, 32'hc2ae5618, 32'h41d2a6e3, 32'h42893658, 32'hc2b2477a, 32'h42b38f28};
test_weights[8160:8167] = '{32'h408fe5cc, 32'h42a2164d, 32'h42a0cc8e, 32'h42a928b6, 32'h42c75464, 32'h4246816e, 32'hc29def4f, 32'hc285c209};
test_bias[1020:1020] = '{32'hc2a2e756};
test_output[1020:1020] = '{32'hc50adab2};
test_input[8168:8175] = '{32'h41e56a07, 32'h426c328a, 32'hc2c6e9a7, 32'h4229366c, 32'hc12462b6, 32'hc2bcb034, 32'hc2afb761, 32'h42a48161};
test_weights[8168:8175] = '{32'h42b0e1a9, 32'hc2a15e58, 32'h425d44f4, 32'hc15ca433, 32'h41c8e01c, 32'hc251a7e0, 32'h404882e8, 32'hc05ce5d2};
test_bias[1021:1021] = '{32'h410b23a9};
test_output[1021:1021] = '{32'hc582855f};
test_input[8176:8183] = '{32'hc22cce6e, 32'hc05667b8, 32'hc185ab3f, 32'h42979f23, 32'hc28c249b, 32'h420c5c2c, 32'hc2892635, 32'hc2794c5c};
test_weights[8176:8183] = '{32'h4198a918, 32'hc280e3b0, 32'h41ceaf9f, 32'hc23418d0, 32'hc2174876, 32'h41a3bb81, 32'hc18fed21, 32'h428d99a6};
test_bias[1022:1022] = '{32'hc282f94a};
test_output[1022:1022] = '{32'hc5874c4d};
test_input[8184:8191] = '{32'hc2c123ac, 32'hc2b18d8a, 32'h428ac7fd, 32'h41b13aac, 32'h41fe8afd, 32'hc2977b2e, 32'h42a67513, 32'hc1e31222};
test_weights[8184:8191] = '{32'h42c75237, 32'hbff503c9, 32'hc19dc002, 32'h42206cbc, 32'hc2bd7e15, 32'h41cb1b7f, 32'h422c7b9e, 32'hc2050a5c};
test_bias[1023:1023] = '{32'hc15277e5};
test_output[1023:1023] = '{32'hc621bf56};
test_input[8192:8199] = '{32'h4270c1f6, 32'h425e31ac, 32'hc1c17da4, 32'h4288b50b, 32'h422618ac, 32'hc1ae1cea, 32'hc2661016, 32'h42b5d95c};
test_weights[8192:8199] = '{32'h4242c595, 32'hc1ddda46, 32'h3f938b4c, 32'hc1ce4993, 32'hc2aba992, 32'h4208a6e5, 32'hc2a47b4b, 32'h423cd3a8};
test_bias[1024:1024] = '{32'hc1a6e929};
test_output[1024:1024] = '{32'h45862ebf};
test_input[8200:8207] = '{32'h41574943, 32'h41592276, 32'hc1fd30c5, 32'hc2367b1d, 32'hc2c32810, 32'h40cb7939, 32'h4282753e, 32'h42c67263};
test_weights[8200:8207] = '{32'h421d2bfe, 32'h4282bbf1, 32'hc2a35ceb, 32'h427f0c3b, 32'h418e90d1, 32'hc2b9f081, 32'h42a0bd31, 32'hc0bb325a};
test_bias[1025:1025] = '{32'h4291b5a6};
test_output[1025:1025] = '{32'h455a8d84};
test_input[8208:8215] = '{32'h42b2575a, 32'h40e722c2, 32'hc296a72c, 32'h3f8cd14b, 32'hc23e3f3f, 32'h4229791f, 32'hc2a69de6, 32'hc1e3ffac};
test_weights[8208:8215] = '{32'hc2abc435, 32'hc1bd3035, 32'h42aebddc, 32'h41c2f10d, 32'hc29b3aee, 32'h424f19b3, 32'h41a827f4, 32'h40b13605};
test_bias[1026:1026] = '{32'h42bc5e13};
test_output[1026:1026] = '{32'hc62124dc};
test_input[8216:8223] = '{32'h418af221, 32'hc1cb065d, 32'hc29f63bf, 32'hc1ccce6b, 32'h42a825b5, 32'hc269b8d3, 32'hc1460618, 32'hc29b0327};
test_weights[8216:8223] = '{32'hc2352cca, 32'hc22c70f3, 32'hc2972e98, 32'h42600518, 32'h42bcd5b2, 32'h428a0fa3, 32'hc199c7b9, 32'h4181ddcc};
test_bias[1027:1027] = '{32'hc2446a95};
test_output[1027:1027] = '{32'h45f1a7c8};
test_input[8224:8231] = '{32'hbfaa2390, 32'h425f7208, 32'hc27cae93, 32'hc116cf67, 32'h429b4ae7, 32'h41a13008, 32'h41aac959, 32'h428812f7};
test_weights[8224:8231] = '{32'h423e8f7c, 32'h42bb0a4f, 32'h3e2355c9, 32'h40895191, 32'hc0396500, 32'hc2af0a49, 32'h42a8ff91, 32'h4211afb1};
test_bias[1028:1028] = '{32'hc2652bd4};
test_output[1028:1028] = '{32'h45e59510};
test_input[8232:8239] = '{32'hc21df1fd, 32'hc2c75a81, 32'hc1800cef, 32'hc2169712, 32'hc2a9b983, 32'h42ad23a2, 32'hc2811629, 32'h4223401f};
test_weights[8232:8239] = '{32'hc2768c4a, 32'h3f2ef155, 32'hc2c4d11d, 32'h425ccfef, 32'hc28ba97e, 32'hc2319825, 32'hc1d164a5, 32'hc2414e60};
test_bias[1029:1029] = '{32'hc2c58ef4};
test_output[1029:1029] = '{32'h455eb4f8};
test_input[8240:8247] = '{32'hc2105ff9, 32'hc21cdad8, 32'hc2081ad4, 32'hc072f036, 32'h41d43430, 32'hc2a2bcd2, 32'hc2bfef66, 32'h42a19824};
test_weights[8240:8247] = '{32'h41e48b9d, 32'h427abdff, 32'hc1c8ac50, 32'hc2ab8b35, 32'h41a9971b, 32'h412e0c04, 32'hc26baeb1, 32'hc10ee580};
test_bias[1030:1030] = '{32'hc1590d0e};
test_output[1030:1030] = '{32'h450ee51a};
test_input[8248:8255] = '{32'h42c24b43, 32'hc29815ca, 32'h41661ede, 32'h418f6517, 32'hc2691faa, 32'h4209e5ac, 32'h406ce221, 32'h417627c0};
test_weights[8248:8255] = '{32'hc1ebb60e, 32'hc2aeb8a3, 32'h4186b683, 32'h42403187, 32'h40633be1, 32'h42af29ef, 32'hc19540fd, 32'hc294f416};
test_bias[1031:1031] = '{32'h422a56f9};
test_output[1031:1031] = '{32'h45cbe2c2};
test_input[8256:8263] = '{32'hc1e95b0b, 32'h4257e075, 32'hc13b6c6b, 32'hc20d53fb, 32'h42b1550c, 32'h41e4d68c, 32'hc1fcb78a, 32'hc2936ef8};
test_weights[8256:8263] = '{32'hc28b0804, 32'h4293fb3b, 32'hc231a712, 32'hc29edaed, 32'hc28c53f1, 32'h427300b7, 32'h42bb108c, 32'hc1d9a3b2};
test_bias[1032:1032] = '{32'hc0401ee1};
test_output[1032:1032] = '{32'h45747f1a};
test_input[8264:8271] = '{32'h3fd04599, 32'hc25c03c3, 32'h42b31099, 32'hc29d5e52, 32'h41d9ba93, 32'hc2a7d53f, 32'h42a08a08, 32'h411393d7};
test_weights[8264:8271] = '{32'h42adfc9f, 32'h41e072cf, 32'hc257867d, 32'hc22c01e9, 32'hc0eec409, 32'hc1da7e66, 32'h427a6cd6, 32'hc290e505};
test_bias[1033:1033] = '{32'h423aca3f};
test_output[1033:1033] = '{32'h456427dd};
test_input[8272:8279] = '{32'hc293dc1b, 32'hc25b2857, 32'h42ad9002, 32'h425d7a8d, 32'hc25792c5, 32'hc2394e6e, 32'h429d84cc, 32'hc1cfe39d};
test_weights[8272:8279] = '{32'hc02e6c8c, 32'hc00593d0, 32'hc1206455, 32'hc0014d74, 32'h41800e52, 32'h424880b3, 32'hc146f3ab, 32'hc2817a5b};
test_bias[1034:1034] = '{32'h42bc2073};
test_output[1034:1034] = '{32'hc53edbd6};
test_input[8280:8287] = '{32'h402d26c6, 32'hc290152f, 32'hc238ecc3, 32'h419a2813, 32'hc0cae4bb, 32'h41a1cdb9, 32'hc20dd7fa, 32'hc249552e};
test_weights[8280:8287] = '{32'hc2b0217b, 32'h42427413, 32'h421d8ee5, 32'hc2a52462, 32'h42466087, 32'hc2776967, 32'h423620a4, 32'h4271a504};
test_bias[1035:1035] = '{32'hc2b961d0};
test_output[1035:1035] = '{32'hc65267fe};
test_input[8288:8295] = '{32'h4250ba27, 32'h4210d45e, 32'hc1ce5621, 32'h419ff88c, 32'hc1e4d464, 32'hc241aeee, 32'hc2a22b89, 32'h42bef807};
test_weights[8288:8295] = '{32'h4273914d, 32'hc25d4b5e, 32'hc2aca51c, 32'h41bd2aa5, 32'hc2c4aeca, 32'hc0e7c62f, 32'h41cdbd64, 32'h421bffaa};
test_bias[1036:1036] = '{32'h4244ad33};
test_output[1036:1036] = '{32'h460853d2};
test_input[8296:8303] = '{32'h423054cb, 32'h4282e6de, 32'hc26e5587, 32'hc26d8734, 32'hc11e6330, 32'h4129a91e, 32'h42b46341, 32'hc2b0d911};
test_weights[8296:8303] = '{32'hc2b5ffb6, 32'hc23f66c6, 32'hc14c22c7, 32'h4286edd6, 32'h41b4416f, 32'h41377e89, 32'h42972def, 32'hc2c175ee};
test_bias[1037:1037] = '{32'hc2c19524};
test_output[1037:1037] = '{32'h45957b70};
test_input[8304:8311] = '{32'hc29e0213, 32'h42c5ae3e, 32'hc2425b86, 32'hc208e4aa, 32'h42710f7d, 32'hc299c5d8, 32'h41b6cdd6, 32'hc1aa98df};
test_weights[8304:8311] = '{32'hc045b4d1, 32'hc208f4dd, 32'h41b7c40d, 32'h4268f2e8, 32'hc2931a3b, 32'hc2a61d9a, 32'hc2b13419, 32'hc2b7c0eb};
test_bias[1038:1038] = '{32'hbff37964};
test_output[1038:1038] = '{32'hc5885956};
test_input[8312:8319] = '{32'hc1919642, 32'hc2844d3e, 32'h40abe39d, 32'hc15b5d73, 32'h429db1b0, 32'hc2bd79b7, 32'h427a56d4, 32'h42b81df8};
test_weights[8312:8319] = '{32'h412a9545, 32'hc18ca900, 32'h41956fa3, 32'hc223ea47, 32'hc2114084, 32'hc2ac0a7b, 32'hc2a283a6, 32'h413782d4};
test_bias[1039:1039] = '{32'h4292deed};
test_output[1039:1039] = '{32'h453914b0};
test_input[8320:8327] = '{32'h42c009a2, 32'h42bc7c32, 32'h425df04f, 32'hc1b841b2, 32'h4177bbab, 32'h42324ca4, 32'hc1e55264, 32'h411f0cb0};
test_weights[8320:8327] = '{32'h429daf00, 32'h42b1e99e, 32'h3f9f7407, 32'hc2c3c794, 32'h4213fc36, 32'h41c0b6da, 32'hc2af7d79, 32'h420a5902};
test_bias[1040:1040] = '{32'h42b40d6a};
test_output[1040:1040] = '{32'h46b2b254};
test_input[8328:8335] = '{32'h42aeeb42, 32'h41bb4953, 32'hc2c0cf80, 32'h41cf0df4, 32'hbde66c95, 32'hc2b11ef5, 32'h41fa2885, 32'h4284ced4};
test_weights[8328:8335] = '{32'h4295c8d9, 32'hc1cd51d6, 32'hc26845a9, 32'hc0f42e2b, 32'h418a3695, 32'h3f5d83d6, 32'hc26e2025, 32'h411bfab2};
test_bias[1041:1041] = '{32'hc29ea0e3};
test_output[1041:1041] = '{32'h461be6cf};
test_input[8336:8343] = '{32'h409da601, 32'h427156ce, 32'hc2b06f93, 32'h42878b29, 32'hc2a45306, 32'hc16318e9, 32'hc263747f, 32'h41d0c34b};
test_weights[8336:8343] = '{32'hc18c02a1, 32'h41393040, 32'hc2b4b5c0, 32'hc23359c1, 32'h424cf95e, 32'h42980be3, 32'h42441846, 32'hc1f1441c};
test_bias[1042:1042] = '{32'h42ab0fcc};
test_output[1042:1042] = '{32'hc54a2243};
test_input[8344:8351] = '{32'h429584cb, 32'hc292a369, 32'h42c4209f, 32'hc23f8bd7, 32'h41b1b6d5, 32'hc245203a, 32'h42a116fc, 32'h4292f05f};
test_weights[8344:8351] = '{32'hc177c0c7, 32'hc2844ba3, 32'h40dc012f, 32'h42c3c154, 32'h40c71457, 32'hc2b2ec7d, 32'h41269324, 32'hc0feb685};
test_bias[1043:1043] = '{32'hc1214d1c};
test_output[1043:1043] = '{32'h458bb11b};
test_input[8352:8359] = '{32'h42ab7ef0, 32'hc2bd6e27, 32'hc29c3808, 32'h41ab194a, 32'hc2a57839, 32'h42bc3914, 32'hc2187208, 32'h423e9647};
test_weights[8352:8359] = '{32'hc160828a, 32'h41b6e60b, 32'hc295f1d1, 32'h42b044be, 32'hc1a4ddd5, 32'h41f08d40, 32'h42a9818a, 32'hc2c1625a};
test_bias[1044:1044] = '{32'h42c25d92};
test_output[1044:1044] = '{32'h4491ea23};
test_input[8360:8367] = '{32'h401491a6, 32'h422e31d9, 32'hbf9a3d69, 32'h426d64fe, 32'hc18561a4, 32'hc1c0b1bc, 32'hc28732ad, 32'hc266c4ea};
test_weights[8360:8367] = '{32'h41e4f90d, 32'hc18477e9, 32'h4291e22e, 32'hc2aca82c, 32'hc289be8f, 32'hc2bb70a3, 32'hc28619b1, 32'hc1662248};
test_bias[1045:1045] = '{32'hc275f231};
test_output[1045:1045] = '{32'h45318831};
test_input[8368:8375] = '{32'hc292ac7d, 32'h41917d36, 32'h419cf037, 32'hc27d1f9a, 32'h42a28ad7, 32'h414f550b, 32'h42ad11db, 32'hc2902734};
test_weights[8368:8375] = '{32'h4217b853, 32'hc286cbc1, 32'h428c4984, 32'h40c799f7, 32'hc2a82c7b, 32'h4237753d, 32'hc2428a3a, 32'h42b3fc46};
test_bias[1046:1046] = '{32'hc0f3de88};
test_output[1046:1046] = '{32'hc69c0063};
test_input[8376:8383] = '{32'hc19572f6, 32'hc2ae109b, 32'hc2884637, 32'hc222a8c3, 32'hc21833c7, 32'h42539957, 32'h42ba44f3, 32'hc293b557};
test_weights[8376:8383] = '{32'hc17ee5c2, 32'h4042887f, 32'hc2a07679, 32'h42a43965, 32'h42b08d70, 32'hc2561cc7, 32'h429e1d98, 32'hc2489b28};
test_bias[1047:1047] = '{32'hc23ec6ca};
test_output[1047:1047] = '{32'h45da6b03};
test_input[8384:8391] = '{32'h42afe0c0, 32'h41cb7c09, 32'h417de185, 32'hc2c5a2f6, 32'hc23be9c1, 32'h4285d53f, 32'hc2714214, 32'hc26e8c67};
test_weights[8384:8391] = '{32'hc0f2d019, 32'h41e45d8c, 32'hc155b34b, 32'h411f7e55, 32'h41e608e6, 32'h40ebd665, 32'hc295eb7c, 32'h42b27ee2};
test_bias[1048:1048] = '{32'h42827c58};
test_output[1048:1048] = '{32'hc52abe8c};
test_input[8392:8399] = '{32'h42840b2d, 32'h42252407, 32'h42b8f0ca, 32'hc2c75b2c, 32'h42aaeed0, 32'hc267a53f, 32'hc1882d51, 32'hc2221640};
test_weights[8392:8399] = '{32'hc266fca2, 32'h42c71599, 32'h42a25942, 32'hc1ada5c3, 32'hc194c403, 32'h4289d74e, 32'h427e4dac, 32'hc2849ba4};
test_bias[1049:1049] = '{32'hc2a93ef2};
test_output[1049:1049] = '{32'h45b891e3};
test_input[8400:8407] = '{32'hc283365d, 32'h42a891c8, 32'hc2650b1e, 32'hc1a27137, 32'h42a79a0a, 32'h3f7883c5, 32'h41cc3a63, 32'hc10c9580};
test_weights[8400:8407] = '{32'h42315833, 32'hc2915b65, 32'hc24034e5, 32'hc2b5fae6, 32'h42b200de, 32'hc2aaae14, 32'hc207ef95, 32'hc1a3be71};
test_bias[1050:1050] = '{32'h41de1ca0};
test_output[1050:1050] = '{32'h450e843d};
test_input[8408:8415] = '{32'h41596f9d, 32'hc2511ce0, 32'h425a9f30, 32'h41c240f4, 32'hc045633c, 32'h4230e79b, 32'hc2a22026, 32'hc27dba24};
test_weights[8408:8415] = '{32'h41bf1e30, 32'h4110f323, 32'h419d4e0a, 32'hc2b2bd06, 32'hc2b0cfa2, 32'hc1de0c58, 32'hc2aa6fac, 32'h41ebbb9f};
test_bias[1051:1051] = '{32'h403729ba};
test_output[1051:1051] = '{32'h4531a955};
test_input[8416:8423] = '{32'h427f703b, 32'h428a4e45, 32'hc2831b69, 32'hc2c5ae6e, 32'hc2899540, 32'h42ab922f, 32'hc1ca4bb1, 32'hc21c6a00};
test_weights[8416:8423] = '{32'hc2108148, 32'h42b4c3c8, 32'hc2903d7e, 32'hc17af2cc, 32'hc20dc022, 32'hc19b792e, 32'hc272a951, 32'hc0647120};
test_bias[1052:1052] = '{32'hc2937d13};
test_output[1052:1052] = '{32'h4644beb6};
test_input[8424:8431] = '{32'h42b821db, 32'h428c92a9, 32'h42ab0342, 32'hc24da242, 32'hc1b20914, 32'h420e2482, 32'h4194c75f, 32'hc201c6f9};
test_weights[8424:8431] = '{32'h41d38f0f, 32'hc2049463, 32'hc298eb36, 32'h41aa1d7f, 32'h4264b128, 32'h42c3667c, 32'hc2990a30, 32'hc2499e05};
test_bias[1053:1053] = '{32'hc25ea0e0};
test_output[1053:1053] = '{32'hc5a18e6c};
test_input[8432:8439] = '{32'h4269143e, 32'h42adefd2, 32'h4286a01a, 32'hc28faee7, 32'hc1526716, 32'hc1e2d0e6, 32'h41bc7553, 32'hc2a4e3c2};
test_weights[8432:8439] = '{32'h41f85382, 32'hc2914a80, 32'hc2c453d4, 32'h41abaa8d, 32'hbffb1a8f, 32'h42b68228, 32'hc26ffdbb, 32'hc293b83f};
test_bias[1054:1054] = '{32'h423f0f9e};
test_output[1054:1054] = '{32'hc6240058};
test_input[8440:8447] = '{32'h429e9be5, 32'h4289516b, 32'hc2a8cee2, 32'h42b3652f, 32'hc233c064, 32'h428761d5, 32'hc21ec621, 32'hc21e8632};
test_weights[8440:8447] = '{32'h4246003b, 32'hc295ed55, 32'hc2c1877d, 32'hc2166558, 32'hc23e29ef, 32'h42bd9831, 32'hc2a012a4, 32'hc2883e86};
test_bias[1055:1055] = '{32'hc299b13e};
test_output[1055:1055] = '{32'h468c0d35};
test_input[8448:8455] = '{32'hc220f0d1, 32'hc20d3cb9, 32'h410d874d, 32'h40e33ab5, 32'hc2704480, 32'h421537bc, 32'h428e3b19, 32'h4169c8ce};
test_weights[8448:8455] = '{32'h4252eb58, 32'hc25308fe, 32'h4273c2db, 32'hc2a40f72, 32'h4260b4e3, 32'hc22488f3, 32'hc2c7da32, 32'hc2c09bd2};
test_bias[1056:1056] = '{32'h4156e9a5};
test_output[1056:1056] = '{32'hc6563bfe};
test_input[8456:8463] = '{32'hc034515f, 32'hc1fb7993, 32'h41e5c110, 32'h4259f3fc, 32'hc1a73bb0, 32'h42825b78, 32'hc1285b48, 32'h416b4bf8};
test_weights[8456:8463] = '{32'h41cafc3c, 32'hc29b52c5, 32'hc28b84ca, 32'h42c5842a, 32'hc107b25b, 32'hc20400e4, 32'hc2948b5a, 32'hc281ede5};
test_bias[1057:1057] = '{32'h4153b7e4};
test_output[1057:1057] = '{32'h4561d300};
test_input[8464:8471] = '{32'hc1eb8572, 32'hc1cd0e0c, 32'h418dc68c, 32'h42586d9e, 32'hc2afc749, 32'h418db21a, 32'h425b39e2, 32'hc27bb449};
test_weights[8464:8471] = '{32'h42933bc2, 32'hc23305bb, 32'h4231da4f, 32'h4272cd7e, 32'hc2c12a84, 32'h41e3d174, 32'h420f6d36, 32'hc2869a64};
test_bias[1058:1058] = '{32'h423115ea};
test_output[1058:1058] = '{32'h468ee351};
test_input[8472:8479] = '{32'h41e3811b, 32'h419565c1, 32'hc2852731, 32'hc2acf33b, 32'h4206ce54, 32'h42a7b718, 32'hc218da59, 32'h414b37a0};
test_weights[8472:8479] = '{32'hc2a1821e, 32'h42aa2cac, 32'hc27929e1, 32'h41de49ea, 32'hc2148548, 32'h428b5a2a, 32'h41d1c3d7, 32'hc191e3e7};
test_bias[1059:1059] = '{32'h4195cede};
test_output[1059:1059] = '{32'h4589eba8};
test_input[8480:8487] = '{32'hc1bd9777, 32'h41da9930, 32'hc2b2e6d5, 32'h42575471, 32'hc10aef85, 32'h41be9532, 32'h42aadd97, 32'h42505ca0};
test_weights[8480:8487] = '{32'h4187f9c7, 32'h42a4d5ad, 32'h41c7e5f5, 32'h421bcd6b, 32'hc2800e11, 32'hc2ba694c, 32'h409c9391, 32'h429d6b6f};
test_bias[1060:1060] = '{32'h42bb4e98};
test_output[1060:1060] = '{32'h45919152};
test_input[8488:8495] = '{32'hc234ec2b, 32'h42064004, 32'h42c0a056, 32'hc2b6870d, 32'h420d0e78, 32'h427b073d, 32'h4285a2d8, 32'hc21dce97};
test_weights[8488:8495] = '{32'h4131f9de, 32'hc2a7a450, 32'h4293640e, 32'h42260e07, 32'h41eb693c, 32'hc28d9211, 32'hc1df09b3, 32'h422866c4};
test_bias[1061:1061] = '{32'h41c8bfba};
test_output[1061:1061] = '{32'hc5d7f419};
test_input[8496:8503] = '{32'h3d6d1f76, 32'hc2598181, 32'hc1396d48, 32'h42267e09, 32'hc2925f82, 32'hc2af48f2, 32'hc21c4daa, 32'h408f0f98};
test_weights[8496:8503] = '{32'h414ceb0e, 32'h41cbc41a, 32'hc260ec35, 32'hc21e34a8, 32'h417270ed, 32'h4283085c, 32'h429328a0, 32'hc2b56d70};
test_bias[1062:1062] = '{32'hc1adbde5};
test_output[1062:1062] = '{32'hc643d117};
test_input[8504:8511] = '{32'h42c5e931, 32'h40b6cd02, 32'h4244c22e, 32'hc24fa0d7, 32'hc2c0bb1a, 32'h4265fdab, 32'hc22b13ac, 32'hc2a50f9b};
test_weights[8504:8511] = '{32'hc10eae15, 32'h426eeac3, 32'h42b31e5d, 32'h42579d35, 32'hc1bccdf5, 32'hc1b53757, 32'hc113893d, 32'hc24f9a74};
test_bias[1063:1063] = '{32'hc2815384};
test_output[1063:1063] = '{32'h45cfd918};
test_input[8512:8519] = '{32'hc258e9d0, 32'h426c9882, 32'hc2bc6f49, 32'hc27f1f7a, 32'h427c050d, 32'h416c1f33, 32'h42b08425, 32'hc24b3b50};
test_weights[8512:8519] = '{32'h4221c41b, 32'h42857b4c, 32'hc2a8a2af, 32'h4269c257, 32'hc2abfa2c, 32'hc1e3aca6, 32'hc2221197, 32'h41b31166};
test_bias[1064:1064] = '{32'h42a6d79b};
test_output[1064:1064] = '{32'hc58c8093};
test_input[8520:8527] = '{32'hc1271bf2, 32'hc2ba61f5, 32'h42309e02, 32'h408b6d35, 32'h42514e62, 32'hc2b13dd9, 32'hc28dc67e, 32'h42220b17};
test_weights[8520:8527] = '{32'h42b49773, 32'h419d74dc, 32'h427092bc, 32'h423120f9, 32'hc2b8bfee, 32'h409e0bc0, 32'hc20d4954, 32'h42b49d6b};
test_bias[1065:1065] = '{32'h41d5c06a};
test_output[1065:1065] = '{32'h44773aaf};
test_input[8528:8535] = '{32'hc2a94aa5, 32'h40d527a3, 32'h41ece100, 32'h428101a6, 32'h421e3097, 32'h4194d6d2, 32'hc090a88b, 32'h3ed3b082};
test_weights[8528:8535] = '{32'h4206a15e, 32'hc2344633, 32'h41a973b2, 32'h424600d7, 32'h40361e3b, 32'h42a903c2, 32'hc2ad2c00, 32'h423a3ff2};
test_bias[1066:1066] = '{32'hc26d95a3};
test_output[1066:1066] = '{32'h45293064};
test_input[8536:8543] = '{32'h41442a82, 32'h42b00768, 32'h4110c001, 32'hc27b6a4c, 32'h4190c8dc, 32'hc2c10b66, 32'hc2a312e5, 32'hc17a585f};
test_weights[8536:8543] = '{32'hc1fef16c, 32'h422ab2b6, 32'h417d325e, 32'hc27048f4, 32'h4180e1c5, 32'hc2ac8cfe, 32'hc246f9ef, 32'hc23d3012};
test_bias[1067:1067] = '{32'hc243829c};
test_output[1067:1067] = '{32'h46a154a8};
test_input[8544:8551] = '{32'hc13cb32d, 32'h4278b8a9, 32'h42a589a4, 32'hc0a80451, 32'h42c5df1b, 32'h4251db23, 32'h42479020, 32'hc03b6c40};
test_weights[8544:8551] = '{32'h423ee52c, 32'h41d637a2, 32'hc2ba6c11, 32'h4259fa0d, 32'hc29832d0, 32'h42b842f1, 32'hc25d8842, 32'hc2bb0bc3};
test_bias[1068:1068] = '{32'hc28d3944};
test_output[1068:1068] = '{32'hc63de895};
test_input[8552:8559] = '{32'h421ff3c6, 32'hc299e222, 32'hc2832806, 32'hc20295df, 32'h423eb59e, 32'hc266ef77, 32'hc1d0513b, 32'h428ec226};
test_weights[8552:8559] = '{32'hc1f9f66a, 32'h429cb74a, 32'h3eaa1f7d, 32'h415dfc0d, 32'h4288c6dc, 32'h42605398, 32'hbf946bfb, 32'h41a5aa8d};
test_bias[1069:1069] = '{32'h428917fc};
test_output[1069:1069] = '{32'hc5c04c14};
test_input[8560:8567] = '{32'h41248e7a, 32'h4248e7fd, 32'h424f0210, 32'hc184f42a, 32'h42a10664, 32'h429cd0e6, 32'hc224178b, 32'hc28e618d};
test_weights[8560:8567] = '{32'h42a06114, 32'hc2097fd0, 32'h425d9670, 32'h42743a3f, 32'h422977ea, 32'h422e5de7, 32'h4288e852, 32'hc1e0a54b};
test_bias[1070:1070] = '{32'h423c5653};
test_output[1070:1070] = '{32'h45db4b28};
test_input[8568:8575] = '{32'h426dd8e9, 32'h42aca781, 32'hc2a993c7, 32'h4218f6ea, 32'hc0aa7646, 32'h415dd44b, 32'hc2c21696, 32'hc2426cab};
test_weights[8568:8575] = '{32'hc2be50a3, 32'h427d1ea9, 32'hc2011dba, 32'h413641eb, 32'h429f8d0d, 32'hc19572ef, 32'h424c023c, 32'hc2a2a652};
test_bias[1071:1071] = '{32'h41d42038};
test_output[1071:1071] = '{32'h44a560b3};
test_input[8576:8583] = '{32'h415c652c, 32'h40fed40b, 32'hc29e929a, 32'hc211ff93, 32'hc2804f12, 32'h41f7571b, 32'h42a175a3, 32'h42c268ce};
test_weights[8576:8583] = '{32'h429994c9, 32'h42664e27, 32'h42a7a3d4, 32'h42340aa7, 32'hc2117868, 32'h41b9a7ee, 32'hc2b24fbf, 32'h42239d07};
test_bias[1072:1072] = '{32'hc1793718};
test_output[1072:1072] = '{32'hc5d9769b};
test_input[8584:8591] = '{32'hc2b666c1, 32'h42b4ec7e, 32'h4289794b, 32'hc28e30eb, 32'h42750068, 32'hc27be83f, 32'h42ae91cb, 32'hc23e7f13};
test_weights[8584:8591] = '{32'hc28a963f, 32'h420b1c06, 32'h42afb6ef, 32'h3dba6c15, 32'h427bc128, 32'hc1ddaa80, 32'h424575c3, 32'h42a772e9};
test_bias[1073:1073] = '{32'h4206329b};
test_output[1073:1073] = '{32'h46a79a84};
test_input[8592:8599] = '{32'hc2ab6975, 32'hc29b00ed, 32'h42870c3b, 32'hc2125b7b, 32'hc20d9f73, 32'h4287a439, 32'hc1b8a32d, 32'hc2c4786b};
test_weights[8592:8599] = '{32'hc1fbffeb, 32'h40c03e06, 32'hc2a0a6c2, 32'h421281b0, 32'h41ca4f07, 32'hc1b936b8, 32'h426af727, 32'h42aa5902};
test_bias[1074:1074] = '{32'hc2791652};
test_output[1074:1074] = '{32'hc6831906};
test_input[8600:8607] = '{32'h41e1f0d7, 32'hc2ae8169, 32'h428d4a57, 32'h422ba420, 32'h421522e7, 32'hc20ea690, 32'h42ba28c1, 32'h3f427f11};
test_weights[8600:8607] = '{32'hc1ff6c88, 32'h41e38379, 32'hc2c3479c, 32'hc202888e, 32'h42456790, 32'hc2036db9, 32'hc0ebc991, 32'h41d95cb1};
test_bias[1075:1075] = '{32'h418315c1};
test_output[1075:1075] = '{32'hc6119901};
test_input[8608:8615] = '{32'hbfd7d609, 32'hc0d83231, 32'h422001bb, 32'hc2161e10, 32'h418d41d7, 32'h42ae9d09, 32'h42c485e7, 32'h42056bd0};
test_weights[8608:8615] = '{32'h40f900eb, 32'h42b29fbc, 32'h41a32c3a, 32'hc297ebf4, 32'h424597b5, 32'hc1ef75f7, 32'h4285062a, 32'h429a5fca};
test_bias[1076:1076] = '{32'hc2b49624};
test_output[1076:1076] = '{32'h462163b7};
test_input[8616:8623] = '{32'hc289b3f1, 32'h41edc8da, 32'hc2ab2026, 32'hc273b066, 32'h4259bce4, 32'h42628ce1, 32'hc2447e23, 32'h427bac44};
test_weights[8616:8623] = '{32'hc1146738, 32'h422bbfd4, 32'h3f9eb531, 32'hc2a248db, 32'h42bc533b, 32'hc29c1141, 32'h4194e1ea, 32'hc2b1b988};
test_bias[1077:1077] = '{32'h42b493c2};
test_output[1077:1077] = '{32'h44826667};
test_input[8624:8631] = '{32'hc1afae1a, 32'h42866aac, 32'h42a158e4, 32'hc20e9956, 32'h403c497c, 32'h42c7b762, 32'hc29d7b23, 32'h4293c1df};
test_weights[8624:8631] = '{32'hc28d904e, 32'hc14aefd5, 32'h4253b690, 32'hc2c416a0, 32'hc2b546ef, 32'h41fa08ea, 32'hc28ca24e, 32'h4220a818};
test_bias[1078:1078] = '{32'hc2a24524};
test_output[1078:1078] = '{32'h469a40c0};
test_input[8632:8639] = '{32'hc1890b31, 32'hc28793fe, 32'hc28033cd, 32'hc2a5c086, 32'h423097a8, 32'hc1b88a27, 32'h420461b9, 32'hc2365c5f};
test_weights[8632:8639] = '{32'h40c6e189, 32'h429b359c, 32'hc2c75bac, 32'h411fee69, 32'h423b3585, 32'h427d7169, 32'h42a9a385, 32'hc29044db};
test_bias[1079:1079] = '{32'h41e2139b};
test_output[1079:1079] = '{32'h45d854d3};
test_input[8640:8647] = '{32'h41a11471, 32'hc266ab89, 32'h42ad947d, 32'hc29e5086, 32'h41f495e9, 32'h4290a195, 32'hc27de9d2, 32'hc24d8ec0};
test_weights[8640:8647] = '{32'h410775b3, 32'h42561fe5, 32'hc2490c52, 32'hc2286c93, 32'hc1eb7d52, 32'h42a52382, 32'h42be4e5a, 32'h3e87f871};
test_bias[1080:1080] = '{32'hc276e635};
test_output[1080:1080] = '{32'hc59bf1c2};
test_input[8648:8655] = '{32'hc2a35612, 32'hc279f2b7, 32'hc2a225c0, 32'h4198a034, 32'h42a71c8a, 32'h412d77a3, 32'h41d148e8, 32'h419f739d};
test_weights[8648:8655] = '{32'hc29df014, 32'h42048146, 32'hc0ddb89e, 32'hc29767ed, 32'hc1d60055, 32'hc2593d82, 32'hc293c581, 32'h403a996a};
test_bias[1081:1081] = '{32'hc160e8af};
test_output[1081:1081] = '{32'hc498013d};
test_input[8656:8663] = '{32'hc2ace4d0, 32'hc2981579, 32'hc2b94cb8, 32'h42b46fff, 32'h42801932, 32'hc29ff4b5, 32'h42830df4, 32'h42937694};
test_weights[8656:8663] = '{32'h427c7dc9, 32'h4251eeed, 32'h42aae24e, 32'hc28e5dd6, 32'h4266de4d, 32'hc0bbcc55, 32'hc2413987, 32'hc2877d0c};
test_bias[1082:1082] = '{32'h4283793e};
test_output[1082:1082] = '{32'hc6d884c5};
test_input[8664:8671] = '{32'h42674ef6, 32'hc2bc8780, 32'h429748de, 32'hbdd4153e, 32'h4292f3fb, 32'hc210f35f, 32'h419ed89a, 32'h41ad8e3b};
test_weights[8664:8671] = '{32'h419d30b2, 32'hc28e67d1, 32'hc091874c, 32'h429e4172, 32'hc1593e22, 32'h42a6e3e8, 32'hc2bf8412, 32'h426e9e06};
test_bias[1083:1083] = '{32'hc20b6fb6};
test_output[1083:1083] = '{32'h45310672};
test_input[8672:8679] = '{32'hc20e09d2, 32'hc2760978, 32'hc20169fa, 32'hc277bf4e, 32'h420c6893, 32'h41c5896a, 32'h42b143ff, 32'h4233ba4f};
test_weights[8672:8679] = '{32'h42c43f53, 32'hc196b918, 32'h427f1012, 32'h429fa326, 32'hc1621a71, 32'hc2628139, 32'hc28462f1, 32'h41abfe06};
test_bias[1084:1084] = '{32'hc2b6b035};
test_output[1084:1084] = '{32'hc67d6af3};
test_input[8680:8687] = '{32'hc22d08b6, 32'h42c69726, 32'hc29032f7, 32'hc2b7b8d0, 32'h428e36a5, 32'hc2c5164a, 32'h41bd34cb, 32'h42abca28};
test_weights[8680:8687] = '{32'hbffa9eb0, 32'h41d9b0ad, 32'h42735c76, 32'hc2891056, 32'hc05c60f6, 32'hc21ba115, 32'hc16f40d9, 32'h422f18dd};
test_bias[1085:1085] = '{32'hc1ccf0ad};
test_output[1085:1085] = '{32'h463645ad};
test_input[8688:8695] = '{32'h41650e7c, 32'hc2b020ca, 32'h426f1ed8, 32'h4252bcee, 32'hc0e657dd, 32'h41bf94f9, 32'h42861019, 32'hc1518516};
test_weights[8688:8695] = '{32'h42abe59c, 32'h429f0d76, 32'h4271ee01, 32'h42bf908c, 32'hc233bce4, 32'hc2943e6f, 32'h429eb384, 32'hc2c0f0c6};
test_bias[1086:1086] = '{32'h40072d14};
test_output[1086:1086] = '{32'h45faad90};
test_input[8696:8703] = '{32'h42841d86, 32'h428dd950, 32'hc27a0f42, 32'hc2989d4d, 32'hc211bbde, 32'hc291aa19, 32'h422f29ef, 32'h42a27b42};
test_weights[8696:8703] = '{32'h429142ee, 32'hc2b9da2a, 32'hc25334ee, 32'hc282aa02, 32'hc2809a19, 32'h422057bf, 32'hc0977f55, 32'h421ea0cc};
test_bias[1087:1087] = '{32'h421f6431};
test_output[1087:1087] = '{32'h460c2b05};
test_input[8704:8711] = '{32'h4141ff48, 32'hc26452af, 32'hc29c39e5, 32'hc0a99f36, 32'hc1dd8f64, 32'h4212d928, 32'h42805851, 32'h42afeeb1};
test_weights[8704:8711] = '{32'hc20eb62b, 32'hc2aab564, 32'hc21e6326, 32'hc1f917f5, 32'hc1ae224b, 32'h42837edc, 32'hc23b68cf, 32'hc013fb4d};
test_bias[1088:1088] = '{32'h42043364};
test_output[1088:1088] = '{32'h45eb894b};
test_input[8712:8719] = '{32'hc29b3b0e, 32'h419d0991, 32'hc0a49321, 32'hc273a770, 32'h40f7fb17, 32'h42b32ccc, 32'h429d435e, 32'hc2c4972e};
test_weights[8712:8719] = '{32'hc1c9c5c2, 32'hc25395b4, 32'hc299c6c9, 32'hc1dad6b8, 32'h426c07d3, 32'h42348911, 32'hc008c8e2, 32'hc2ae360d};
test_bias[1089:1089] = '{32'hc2763e7e};
test_output[1089:1089] = '{32'h46771870};
test_input[8720:8727] = '{32'h42c44eaa, 32'hc2818b45, 32'h3f9894ec, 32'hc287942f, 32'h42a19487, 32'h42479e4d, 32'hc292ea6d, 32'hc138b36f};
test_weights[8720:8727] = '{32'h42941a2b, 32'h42513a25, 32'hc2110e95, 32'hc203eeed, 32'h42bdf9ff, 32'h42adeebc, 32'h42896877, 32'hc2603b53};
test_bias[1090:1090] = '{32'h42c518d9};
test_output[1090:1090] = '{32'h46576809};
test_input[8728:8735] = '{32'hc0be201b, 32'h4287198b, 32'h418002b4, 32'h4263341c, 32'hc1c78ea2, 32'h408b6844, 32'h415ed1f4, 32'hc25802ba};
test_weights[8728:8735] = '{32'h41ac3662, 32'hc29c48b8, 32'h427c3007, 32'h4290ce6d, 32'hc2b90085, 32'h418787ed, 32'hc0d2acae, 32'h42aaf55e};
test_bias[1091:1091] = '{32'h429ff305};
test_output[1091:1091] = '{32'hc51e3977};
test_input[8736:8743] = '{32'hc0d2fe41, 32'hc2c4311a, 32'hc262c2be, 32'h41d635db, 32'hc2b22a74, 32'h424a26c8, 32'hc1e433d8, 32'hc2c7a962};
test_weights[8736:8743] = '{32'h421ec353, 32'hc298538a, 32'h4219cfc4, 32'h42103536, 32'hc27534e6, 32'h42477f22, 32'hc2a51671, 32'hc2a093df};
test_bias[1092:1092] = '{32'h42abe312};
test_output[1092:1092] = '{32'h46bee0a5};
test_input[8744:8751] = '{32'hc20c05c6, 32'hc1ca1215, 32'hc2968a35, 32'h410e91d4, 32'hc1e84d9d, 32'hc20520b7, 32'hc2b6c689, 32'h41e3782c};
test_weights[8744:8751] = '{32'hc17ed5b3, 32'h4249e422, 32'h421a7c3c, 32'h418ab4a0, 32'hc185abba, 32'h40c1b891, 32'h429dd013, 32'h41a6caf0};
test_bias[1093:1093] = '{32'h4130fc92};
test_output[1093:1093] = '{32'hc6190578};
test_input[8752:8759] = '{32'h42a150ac, 32'h41447c8c, 32'h42c29102, 32'hc2b21d71, 32'hc22b497e, 32'h429cdc21, 32'h427c0dc6, 32'h41faa6d1};
test_weights[8752:8759] = '{32'h428e305a, 32'hc1185e99, 32'h4061b8f0, 32'hc2789bf7, 32'h42586635, 32'hc0c79567, 32'hc0adaca5, 32'hc288d1e0};
test_bias[1094:1094] = '{32'h4293ce79};
test_output[1094:1094] = '{32'h45c43273};
test_input[8760:8767] = '{32'h42c6d3a9, 32'hc26b79b9, 32'hc20e6986, 32'h4235f0fc, 32'hc2658877, 32'h42a0b294, 32'h427fc559, 32'hc24bf42a};
test_weights[8760:8767] = '{32'h40995d94, 32'hc2ae279e, 32'hc29e7a10, 32'hc1ce916e, 32'hc119a287, 32'hc2b99a10, 32'h41954707, 32'hc24900be};
test_bias[1095:1095] = '{32'hc0d23e65};
test_output[1095:1095] = '{32'h457fc9ae};
test_input[8768:8775] = '{32'h42767b54, 32'h426320b9, 32'h426bc307, 32'hc2a48129, 32'h410b0a7e, 32'h420eb1c1, 32'hc22f13ab, 32'hc2959ef1};
test_weights[8768:8775] = '{32'h42c285ba, 32'hc26f2c8c, 32'hc2392ced, 32'hc27336e2, 32'h420afc55, 32'h41b8833c, 32'h426a8312, 32'hc26a4197};
test_bias[1096:1096] = '{32'h428e38cc};
test_output[1096:1096] = '{32'h45f64d67};
test_input[8776:8783] = '{32'h42104a26, 32'h425da1e5, 32'h423955dd, 32'hc12f6570, 32'hc2b22d8d, 32'hc2c38969, 32'hc28a5a26, 32'hc2024e1e};
test_weights[8776:8783] = '{32'h41d12eb0, 32'hc27978e7, 32'h41ecfb89, 32'hc2a1081b, 32'hc2466ad8, 32'h41b47113, 32'h42956508, 32'h42c7e469};
test_bias[1097:1097] = '{32'hc24f0634};
test_output[1097:1097] = '{32'hc5cbb187};
test_input[8784:8791] = '{32'h42841bfd, 32'h41370fff, 32'hc1048743, 32'h421fc399, 32'h415c0737, 32'hc290fc44, 32'h41b10e0c, 32'h420b3684};
test_weights[8784:8791] = '{32'hc2687341, 32'h422c5c50, 32'hc2194b82, 32'h426614e3, 32'h426bda25, 32'h42490218, 32'hc2bdef21, 32'hc1fce1d9};
test_bias[1098:1098] = '{32'hc249da31};
test_output[1098:1098] = '{32'hc5d4f990};
test_input[8792:8799] = '{32'hc2a8cc80, 32'hc28572dc, 32'h41d667ab, 32'h42842fcb, 32'h4251f5fd, 32'h41dc8e37, 32'hc10bd1ea, 32'hc1733cf5};
test_weights[8792:8799] = '{32'hc210af70, 32'h41b1e7eb, 32'h41f155cd, 32'h4154f14b, 32'h4247e380, 32'hc201b496, 32'hc27a3172, 32'hc24cd355};
test_bias[1099:1099] = '{32'h427f609f};
test_output[1099:1099] = '{32'h45c738cb};
test_input[8800:8807] = '{32'h41257391, 32'hc1c7745d, 32'hc26671c0, 32'hc1df6842, 32'h423b3a82, 32'h418d0952, 32'h414ddb1c, 32'hc2a188e2};
test_weights[8800:8807] = '{32'h3fddabad, 32'h3fc341fd, 32'hc18cb515, 32'h42ac8c16, 32'hc1e3e4f6, 32'h424e1a18, 32'hc1bb1091, 32'hc29e314c};
test_bias[1100:1100] = '{32'hc212f415};
test_output[1100:1100] = '{32'h45838d8b};
test_input[8808:8815] = '{32'h422c3491, 32'hc295d7b2, 32'hc19b071f, 32'h4285190a, 32'hc1d09f82, 32'h42879deb, 32'h426a0ca2, 32'h412b3736};
test_weights[8808:8815] = '{32'h42030a63, 32'hc22d293b, 32'h402ff338, 32'hc2003670, 32'h42aa4cf5, 32'h418c2522, 32'hc1d20017, 32'hc24fc5a7};
test_bias[1101:1101] = '{32'hc295fff7};
test_output[1101:1101] = '{32'hc43706a5};
test_input[8816:8823] = '{32'h42c2b6c8, 32'hc230ac0e, 32'h4238f52e, 32'hc2aadab8, 32'h4298ae75, 32'hc1595b16, 32'hc04be0b9, 32'h421f9b63};
test_weights[8816:8823] = '{32'hc2475298, 32'hc248aa61, 32'h415b1bee, 32'h427a10a1, 32'h42166e32, 32'hc1b61066, 32'hc10a7e9b, 32'hc1691a1b};
test_bias[1102:1102] = '{32'h42a00453};
test_output[1102:1102] = '{32'hc590e48c};
test_input[8824:8831] = '{32'h4283bd79, 32'hc2183120, 32'h41c0b57c, 32'hc14e12d4, 32'h4273aaa8, 32'hc2b5b237, 32'h429bd748, 32'h4163ed6e};
test_weights[8824:8831] = '{32'hc1aad8e3, 32'hc1d92a24, 32'hc1cbbb3e, 32'h42bc585a, 32'h423f610b, 32'hc2bee5c6, 32'h417de21b, 32'h421e757c};
test_bias[1103:1103] = '{32'hc2acbe2f};
test_output[1103:1103] = '{32'h462d7017};
test_input[8832:8839] = '{32'hc1bccbbb, 32'h3fc2e0e1, 32'hc268689b, 32'hc1949483, 32'hc24346a6, 32'h3c3da099, 32'h420bde23, 32'hc27cab3a};
test_weights[8832:8839] = '{32'hc20cc87f, 32'h423edb08, 32'hc211c66d, 32'h417c3a29, 32'hc127b0ba, 32'h42a1b9cc, 32'hc2459d0c, 32'h42208b57};
test_bias[1104:1104] = '{32'h409f4646};
test_output[1104:1104] = '{32'hc47e5173};
test_input[8840:8847] = '{32'hc23b6d6c, 32'hc243e27d, 32'h4209f238, 32'hc27405cc, 32'hbf9cfe88, 32'hc2ae9cc3, 32'hc22f4eaa, 32'h4231c498};
test_weights[8840:8847] = '{32'hc03fec87, 32'hc281f5fc, 32'h4257f0b0, 32'hc2306fd9, 32'h425cb81c, 32'hc2708be5, 32'hc1828ac2, 32'hc28c66a8};
test_bias[1105:1105] = '{32'h424079c1};
test_output[1105:1105] = '{32'h46273597};
test_input[8848:8855] = '{32'hc28c125c, 32'hc28f8792, 32'hc2adce67, 32'hc2a561c5, 32'hc2b3bc80, 32'hc179c658, 32'h4280d238, 32'hc2224ff5};
test_weights[8848:8855] = '{32'h42baf58c, 32'hc1e27b4e, 32'h42a03084, 32'hc2c2102a, 32'h42c4f1e2, 32'hc29f6fec, 32'h42a07d42, 32'h42000601};
test_bias[1106:1106] = '{32'h42c06fdd};
test_output[1106:1106] = '{32'hc5dd988c};
test_input[8856:8863] = '{32'h417e497e, 32'hc2429439, 32'hc296fb38, 32'hc2773aed, 32'hc2a4189d, 32'h424c88d3, 32'h429407e7, 32'h42b0a98a};
test_weights[8856:8863] = '{32'hc25795cb, 32'hc2297e59, 32'h42644217, 32'h422797b1, 32'hc22f1dd8, 32'hc217a420, 32'h40105720, 32'hc270b83c};
test_bias[1107:1107] = '{32'hc1fcd337};
test_output[1107:1107] = '{32'hc6100ee0};
test_input[8864:8871] = '{32'hc18a1b7b, 32'hc26ecce9, 32'h402877ea, 32'hc0c69da4, 32'h41fafe08, 32'hc2bd3241, 32'hc23f8405, 32'h41f22b99};
test_weights[8864:8871] = '{32'h4255cafe, 32'hc2a1ee85, 32'hc28bdc28, 32'hc23a7a75, 32'hc128d358, 32'hc0f0679d, 32'hc23c965e, 32'hc260ed39};
test_bias[1108:1108] = '{32'hc1134772};
test_output[1108:1108] = '{32'h459a6e87};
test_input[8872:8879] = '{32'h426a7fb7, 32'h425a05ee, 32'h4247a514, 32'h3f0325e1, 32'h42237074, 32'hc17d3b60, 32'hc2a56d4c, 32'h422b0578};
test_weights[8872:8879] = '{32'h413b096a, 32'h4149f32b, 32'h414f14da, 32'h41acd614, 32'hc232024c, 32'h42aa67d7, 32'h40a1def9, 32'hc1b55002};
test_bias[1109:1109] = '{32'h429af44e};
test_output[1109:1109] = '{32'hc518e786};
test_input[8880:8887] = '{32'h41d386a9, 32'h42138d01, 32'h414cb64c, 32'hc2c7fa96, 32'hc29783ed, 32'h42ae4fdc, 32'h4288dc0f, 32'hc2186fb9};
test_weights[8880:8887] = '{32'hc28ac76a, 32'hc2703417, 32'h42c0d8b2, 32'h422bd0ad, 32'h41964976, 32'h416915eb, 32'hc1004c2f, 32'h41d0e019};
test_bias[1110:1110] = '{32'h411c0a23};
test_output[1110:1110] = '{32'hc6097a32};
test_input[8888:8895] = '{32'hc01f9043, 32'h411f4564, 32'h42bcc8c1, 32'h428fea67, 32'h42212e50, 32'h42a15fb9, 32'h423d36cd, 32'h4217f58e};
test_weights[8888:8895] = '{32'hc2a91fe8, 32'hc2aec5bf, 32'hc194b7fd, 32'hc1bab388, 32'hc2a3ca68, 32'hc237495c, 32'h42920713, 32'h413a6760};
test_bias[1111:1111] = '{32'hc2a9751e};
test_output[1111:1111] = '{32'hc5e3751f};
test_input[8896:8903] = '{32'hc28f5261, 32'hc18db890, 32'h41ac2191, 32'h4268a1ad, 32'h42a4fe50, 32'hc02da7bd, 32'h421a1922, 32'h4275ef4b};
test_weights[8896:8903] = '{32'h42919496, 32'h41e3a118, 32'h42760ffa, 32'hc277d3ab, 32'h4203f8bf, 32'hc26a3056, 32'h42858eab, 32'h421524e7};
test_bias[1112:1112] = '{32'hc27bb703};
test_output[1112:1112] = '{32'hc39e8e2a};
test_input[8904:8911] = '{32'hc28b8531, 32'h42c54b2d, 32'hc28b7ab2, 32'hc1b79c48, 32'h424017a6, 32'hc12788d0, 32'h41b7c5b0, 32'h42c1fef5};
test_weights[8904:8911] = '{32'hc233a251, 32'hc2b42903, 32'h40e56e7e, 32'hc2204fc1, 32'h427f23fd, 32'h41b9067a, 32'h42808fc8, 32'h42705c1c};
test_bias[1113:1113] = '{32'h42134357};
test_output[1113:1113] = '{32'h4596ec8b};
test_input[8912:8919] = '{32'h4278dc74, 32'hc140b9d9, 32'h4086ed51, 32'hc19f3f45, 32'hc1d1cc7e, 32'h42a0afe0, 32'h429a4f9a, 32'h42b5319a};
test_weights[8912:8919] = '{32'h4291996b, 32'hc29daa95, 32'hc2836526, 32'h422e2038, 32'h40d92258, 32'h4275cd75, 32'h42023f4c, 32'hbed242c8};
test_bias[1114:1114] = '{32'h42a66e8d};
test_output[1114:1114] = '{32'h4636134f};
test_input[8920:8927] = '{32'h42577d7f, 32'h41c9a562, 32'h424fb297, 32'h41d4a3ce, 32'h428a4e58, 32'hc24f2610, 32'h41d6eb1c, 32'hc2bc31ae};
test_weights[8920:8927] = '{32'hc296aa5b, 32'hc2c07687, 32'hc2a116eb, 32'hc27e3652, 32'h42052b39, 32'h426b170b, 32'h42908d88, 32'hc2a7c1b9};
test_bias[1115:1115] = '{32'hc1e24504};
test_output[1115:1115] = '{32'hc54dab95};
test_input[8928:8935] = '{32'hc2b2d02c, 32'hc23a4c8f, 32'h41f6bf25, 32'hc12c2cfd, 32'h41effb4c, 32'hc25610c2, 32'hc199d143, 32'hc286f2a4};
test_weights[8928:8935] = '{32'h428ca4a6, 32'h419fc785, 32'hc29afe01, 32'h41fce767, 32'hc2536a3a, 32'h422ebe0d, 32'hc29fd725, 32'h4106159b};
test_bias[1116:1116] = '{32'h4271899d};
test_output[1116:1116] = '{32'hc6489ea2};
test_input[8936:8943] = '{32'hc21b8c0f, 32'h41afce23, 32'hc241ce98, 32'hc2973440, 32'h428d8218, 32'hc29adc4f, 32'h42486da4, 32'h42c63167};
test_weights[8936:8943] = '{32'h410e6334, 32'h4121d1a9, 32'hc1a1ddb8, 32'hc2afacf6, 32'h408d8c59, 32'hc2941911, 32'hc2bb8860, 32'hc1026ff8};
test_bias[1117:1117] = '{32'hc2172b80};
test_output[1117:1117] = '{32'h45f9feb0};
test_input[8944:8951] = '{32'hc2b8abe6, 32'h42ac8605, 32'h4206b394, 32'h4191391c, 32'hc2a8df40, 32'hc26a16d7, 32'h4229b910, 32'hc18fc54f};
test_weights[8944:8951] = '{32'hc28894fb, 32'hc236c2e1, 32'hc215fa20, 32'h4077bda0, 32'hc2a18d14, 32'h42a66dee, 32'h42389d01, 32'hc2c119d8};
test_bias[1118:1118] = '{32'hc1bf931d};
test_output[1118:1118] = '{32'h45d43fc5};
test_input[8952:8959] = '{32'hc2b6b31c, 32'hc1fcfc2a, 32'h4217b80f, 32'hc2911bf4, 32'h422ed40e, 32'h40d8fb6f, 32'h419b0a4f, 32'h41cac0de};
test_weights[8952:8959] = '{32'hc21456ff, 32'hc2a00fe7, 32'hc212cb0f, 32'h41ce1f51, 32'h42394b55, 32'hc189b03c, 32'hc1e28e3c, 32'hc2336ad6};
test_bias[1119:1119] = '{32'h4130845b};
test_output[1119:1119] = '{32'h4534a8f2};
test_input[8960:8967] = '{32'h4229f0db, 32'h42bd12dd, 32'h4290e626, 32'hc2a97dec, 32'hc2ba6d8b, 32'h3ea343d8, 32'hc2bc6bce, 32'hc2bdf4c1};
test_weights[8960:8967] = '{32'h40f5891a, 32'h4238a9e2, 32'hc2aa2edd, 32'h426b4646, 32'hc105447f, 32'h414dec99, 32'hc2916eee, 32'h40ddde8c};
test_bias[1120:1120] = '{32'hc2b78eff};
test_output[1120:1120] = '{32'h43d2e21e};
test_input[8968:8975] = '{32'hc0195b34, 32'h4217bcb2, 32'h41c1f1e8, 32'h42abb5f2, 32'h41a83985, 32'h4249653e, 32'hc19bee24, 32'h42aef8eb};
test_weights[8968:8975] = '{32'h419ce7ff, 32'h42ae6b6b, 32'h4269428a, 32'hc26984e9, 32'h4298350c, 32'hc285086a, 32'hc2af04b5, 32'h42237218};
test_bias[1121:1121] = '{32'h42a445cd};
test_output[1121:1121] = '{32'h454cca8d};
test_input[8976:8983] = '{32'h426d97fa, 32'h42052175, 32'h42282a66, 32'hc2951002, 32'h42bf80e4, 32'hc2be908d, 32'h42b1f9d3, 32'h4142be76};
test_weights[8976:8983] = '{32'hc20d4c44, 32'h42b4a34e, 32'h42421222, 32'hc288bf5f, 32'h4220b0c8, 32'hc2190445, 32'h4205e136, 32'h42500587};
test_bias[1122:1122] = '{32'h41e16725};
test_output[1122:1122] = '{32'h4695cd66};
test_input[8984:8991] = '{32'h4295165a, 32'hc039ab8f, 32'h4183a3dc, 32'hc1ad65ba, 32'hc18c7378, 32'h401a4541, 32'h417c9bfb, 32'hc2be51bf};
test_weights[8984:8991] = '{32'h4232eaed, 32'h42aa7e05, 32'h42a11f75, 32'h42a863a3, 32'h426cbf96, 32'h40b3dc42, 32'hc24931f3, 32'h42105e3d};
test_bias[1123:1123] = '{32'hc1f1bec8};
test_output[1123:1123] = '{32'hc5288abd};
test_input[8992:8999] = '{32'h42b323d8, 32'h3fb2a9de, 32'hc2948ad9, 32'h40e182b5, 32'h41ff03a2, 32'hc2b50a32, 32'hc1b91a30, 32'hc137357d};
test_weights[8992:8999] = '{32'hc2c0ac49, 32'h42c1ce24, 32'h4231b35b, 32'h42b15ad0, 32'hc1b37c8b, 32'h4200d7e2, 32'h42a66984, 32'h4182807a};
test_bias[1124:1124] = '{32'hc297c061};
test_output[1124:1124] = '{32'hc684b5ea};
test_input[9000:9007] = '{32'h4273a967, 32'hc2a089c2, 32'h4290ccc5, 32'hc29299f8, 32'h4285f60c, 32'hc2989c3b, 32'hc0c6f38c, 32'hc2c0adbf};
test_weights[9000:9007] = '{32'h428b1f37, 32'hc1986707, 32'h41bc4db0, 32'h4224ceff, 32'h418e6f89, 32'h41d5bc3d, 32'hc1fb5861, 32'h42817eb1};
test_bias[1125:1125] = '{32'hc08ed078};
test_output[1125:1125] = '{32'hc518a74d};
test_input[9008:9015] = '{32'hc21f2020, 32'hc29e79d8, 32'h421ca866, 32'h42863424, 32'hc2a9d3bc, 32'h41b6a8af, 32'h42c7a103, 32'h42784627};
test_weights[9008:9015] = '{32'h422d2029, 32'h427a9b2c, 32'hc275d832, 32'h41e06024, 32'hc2b5554a, 32'hc24bc93c, 32'h420d0543, 32'h4297eae4};
test_bias[1126:1126] = '{32'h42a9af8f};
test_output[1126:1126] = '{32'h45eed652};
test_input[9016:9023] = '{32'h4292b5c7, 32'hc1c74817, 32'h41a888fb, 32'h415b683d, 32'hc2ae11b5, 32'hc139befa, 32'h4152f0ef, 32'hc28a2f16};
test_weights[9016:9023] = '{32'h4250c73f, 32'hc29adb46, 32'h4057293c, 32'h42a5993f, 32'h41aaea13, 32'hc2b91ad0, 32'hc2b656a9, 32'hc188aa2d};
test_bias[1127:1127] = '{32'h41a52bd2};
test_output[1127:1127] = '{32'h45c10dfa};
test_input[9024:9031] = '{32'h425b5d9a, 32'hc0d35250, 32'h42395959, 32'hc2b46042, 32'h40f243ea, 32'h41817a39, 32'h427ea70c, 32'h42ac3d9c};
test_weights[9024:9031] = '{32'h42784cad, 32'hc2612d7e, 32'hc29fd730, 32'h416381fd, 32'hc2c3e05a, 32'hc2bf14ea, 32'hc29ccb98, 32'hc29b3387};
test_bias[1128:1128] = '{32'h429a153c};
test_output[1128:1128] = '{32'hc66bd9ad};
test_input[9032:9039] = '{32'hc296c1a4, 32'h4252fb6a, 32'hc0d60755, 32'h420b273d, 32'h422077d4, 32'h4291093c, 32'h429ed8f4, 32'h42a991af};
test_weights[9032:9039] = '{32'hc2b43a87, 32'hc1af46cc, 32'h428e9f1d, 32'h42c575ee, 32'hc29504d9, 32'hc21c12a0, 32'hc1035034, 32'h4239cd9b};
test_bias[1129:1129] = '{32'h422b0dc2};
test_output[1129:1129] = '{32'h45becac3};
test_input[9040:9047] = '{32'h429a4c5a, 32'hc2a6b183, 32'hc2367d6b, 32'hc2ad5e9f, 32'hc1a75f43, 32'h429fc2ff, 32'hc28f04fa, 32'h4292f2e2};
test_weights[9040:9047] = '{32'hc2aa3f6f, 32'h41158281, 32'h42c14c81, 32'hc2504a5d, 32'h41b2c775, 32'h418ae35d, 32'h427576f0, 32'h429dd3ad};
test_bias[1130:1130] = '{32'hc207d6fb};
test_output[1130:1130] = '{32'hc59a9317};
test_input[9048:9055] = '{32'hc24d407d, 32'hc2b0520e, 32'hc14c5fc0, 32'hc09c9907, 32'h42ba1add, 32'hc1f72140, 32'h4257e72b, 32'h40cac9e8};
test_weights[9048:9055] = '{32'h420367fd, 32'hc28aa894, 32'hc2a654e1, 32'h416fd124, 32'hc235c5cb, 32'h42846e42, 32'h42addc7c, 32'hc2c26958};
test_bias[1131:1131] = '{32'h4281cf12};
test_output[1131:1131] = '{32'h454d24e0};
test_input[9056:9063] = '{32'hc0951455, 32'h42966146, 32'hc2463003, 32'hc14ce595, 32'h418f0f30, 32'h421e2dc4, 32'h42b63011, 32'h41c7a846};
test_weights[9056:9063] = '{32'h41c1adfa, 32'hc26643d8, 32'h41630f98, 32'hc246292c, 32'h41f294d5, 32'hc240fd75, 32'hc22d91d6, 32'h40fb8286};
test_bias[1132:1132] = '{32'hc2008863};
test_output[1132:1132] = '{32'hc6170178};
test_input[9064:9071] = '{32'hc17f95b1, 32'h4186c0ea, 32'hc25772b2, 32'h4224f2eb, 32'h42c22cb2, 32'h419346e8, 32'h424639ce, 32'h4241c13e};
test_weights[9064:9071] = '{32'hc2a7ee67, 32'hc10b8320, 32'h423a5eb4, 32'h3f8721a2, 32'hc0f9426b, 32'h42884c34, 32'h420a6ae0, 32'h4107d3bc};
test_bias[1133:1133] = '{32'h41d29f2c};
test_output[1133:1133] = '{32'h44ac63c0};
test_input[9072:9079] = '{32'h410a66ae, 32'h41d1313d, 32'h4262d0e6, 32'hc1d290b8, 32'h423d7f4e, 32'h4208c8ac, 32'hc1657b1d, 32'hc26f4e4b};
test_weights[9072:9079] = '{32'h42b210d1, 32'hc10336af, 32'h42300858, 32'hc2aa2097, 32'hc29ea3ef, 32'h4291ecaf, 32'h419ab6b4, 32'hc2bb7cd2};
test_bias[1134:1134] = '{32'h420c1bf9};
test_output[1134:1134] = '{32'h4612c56a};
test_input[9080:9087] = '{32'hc2c79869, 32'hc2387eed, 32'hc1232494, 32'hc261e7ce, 32'hc197f9a5, 32'hc2be7494, 32'hc2c57d50, 32'hc280b8f6};
test_weights[9080:9087] = '{32'hc1892fa3, 32'h42ad4e30, 32'h429f07ec, 32'h4204bd98, 32'hc2a0eaea, 32'hc2af1f65, 32'hc28c6b7b, 32'hc2a9f9b0};
test_bias[1135:1135] = '{32'h429bf745};
test_output[1135:1135] = '{32'h4687c242};
test_input[9088:9095] = '{32'hc21ce016, 32'hc284b782, 32'h42bb9376, 32'hc2973f0a, 32'h421e498a, 32'hc28f0c6c, 32'hc2b9f2c1, 32'hc27f510b};
test_weights[9088:9095] = '{32'hc1c14f02, 32'h409ac27b, 32'hc2b24262, 32'hc2a6fffd, 32'h42828e91, 32'hbfbe82ac, 32'h41f79e70, 32'h421dba78};
test_bias[1136:1136] = '{32'h41ac3721};
test_output[1136:1136] = '{32'hc5802c52};
test_input[9096:9103] = '{32'hc2657b11, 32'h41a088c8, 32'h42a34a68, 32'hc2158736, 32'h41f131de, 32'h412e0f01, 32'h41968d2f, 32'hc20e1671};
test_weights[9096:9103] = '{32'h4253ab82, 32'h4250de61, 32'h3fa92657, 32'hc24eb3a3, 32'hc296ef61, 32'h426b2384, 32'hc0fe44a0, 32'h42149570};
test_bias[1137:1137] = '{32'hc2ac718c};
test_output[1137:1137] = '{32'hc54437a3};
test_input[9104:9111] = '{32'h422b3b3b, 32'h412b6945, 32'h4188a035, 32'h427b0f44, 32'h412223fa, 32'hc29c6dc5, 32'hc2a452ec, 32'h425ef8b6};
test_weights[9104:9111] = '{32'h418c53ff, 32'h427d00bb, 32'hc297a3d5, 32'h42894323, 32'hc19df8b7, 32'hc28ed5a6, 32'h42422475, 32'hc1d01c80};
test_bias[1138:1138] = '{32'h429933a3};
test_output[1138:1138] = '{32'h458b8dff};
test_input[9112:9119] = '{32'h42b58093, 32'h428b1875, 32'hc247c4fa, 32'h4133d07e, 32'h426c2369, 32'hc2078ca7, 32'h414072b8, 32'hc29ef836};
test_weights[9112:9119] = '{32'h42b7f4fe, 32'h420854c7, 32'hc20026e4, 32'hc181eae3, 32'h427bd264, 32'hc1c838f8, 32'hc245ba2a, 32'h42851e53};
test_bias[1139:1139] = '{32'hc1511173};
test_output[1139:1139] = '{32'h4628c6b3};
test_input[9120:9127] = '{32'hc2994ab4, 32'hc136b4d3, 32'hc280243e, 32'h40d52f3f, 32'h42823258, 32'hc22194de, 32'hc27866fc, 32'hc2764881};
test_weights[9120:9127] = '{32'h424eaffd, 32'hc298e8b6, 32'h4294a5ac, 32'h42938aa3, 32'hc1b68e37, 32'hc27878e4, 32'h42aa3339, 32'h42712395};
test_bias[1140:1140] = '{32'hc233ee7b};
test_output[1140:1140] = '{32'hc6703e98};
test_input[9128:9135] = '{32'hc22974cf, 32'h42253308, 32'h4274f10b, 32'hc2976927, 32'h41440059, 32'hc261de1b, 32'h42883475, 32'h41d9bc82};
test_weights[9128:9135] = '{32'h41248c92, 32'hc142997c, 32'h42326c45, 32'h41d5e81e, 32'hc1639346, 32'h42a4e09b, 32'h4217e482, 32'hc253e71f};
test_bias[1141:1141] = '{32'h41eb28da};
test_output[1141:1141] = '{32'hc572e753};
test_input[9136:9143] = '{32'hc1035aa9, 32'hc1eb0f18, 32'h429d5246, 32'h41a24cde, 32'hc2034f14, 32'h4252eefe, 32'hc214a10c, 32'h410b128f};
test_weights[9136:9143] = '{32'hc2b7a63b, 32'h40b62414, 32'hc2a2d8fc, 32'h4192d0b1, 32'hc2a932dd, 32'h42ba6e9b, 32'hc290310e, 32'h427b6de3};
test_bias[1142:1142] = '{32'hc26eed82};
test_output[1142:1142] = '{32'h45a922b0};
test_input[9144:9151] = '{32'hc2917878, 32'h429d11d2, 32'hc2914822, 32'hc1512906, 32'hc1df443f, 32'hc22d6062, 32'h4249e3ff, 32'h41952b0e};
test_weights[9144:9151] = '{32'h427dab9f, 32'h40fe8cc3, 32'h426f0984, 32'hc2571809, 32'h4135bb0d, 32'h42b84b7a, 32'hc28a7ae4, 32'h42979cc3};
test_bias[1143:1143] = '{32'h421e470f};
test_output[1143:1143] = '{32'hc65a6acf};
test_input[9152:9159] = '{32'h42abdcda, 32'hc2c48fa6, 32'h42b7673d, 32'h420a15dd, 32'hc2add00e, 32'h410a2877, 32'hc1f1850c, 32'hc2b0e651};
test_weights[9152:9159] = '{32'hc2c1c98f, 32'hc27e935c, 32'h429efb18, 32'h42676795, 32'h4284aa91, 32'h42808ce7, 32'hc1b6ca87, 32'hc1fef286};
test_bias[1144:1144] = '{32'hc26724b0};
test_output[1144:1144] = '{32'h45aa822e};
test_input[9160:9167] = '{32'hc27a8618, 32'hc1d0cbee, 32'hc24add18, 32'h4259da13, 32'h41551215, 32'hc20935f2, 32'h419e3933, 32'hc0960184};
test_weights[9160:9167] = '{32'hc2c35063, 32'hc28e0c38, 32'h41d602b4, 32'hc11b4da5, 32'h42bdd84a, 32'hc0a4a235, 32'h422c6557, 32'hc27784a1};
test_bias[1145:1145] = '{32'hc2bb0507};
test_output[1145:1145] = '{32'h4605f8d5};
test_input[9168:9175] = '{32'h426e54c7, 32'h41baa072, 32'h429a7da0, 32'h42ad5ec9, 32'h40e50d7f, 32'h424fa03f, 32'hc0be1ec5, 32'hc28b84df};
test_weights[9168:9175] = '{32'hc0e49c02, 32'hc09596db, 32'h41270cac, 32'hc220ff73, 32'hc1980e86, 32'hc2b1de07, 32'h40184f14, 32'hc1eaf323};
test_bias[1146:1146] = '{32'h42a101d9};
test_output[1146:1146] = '{32'hc5b6f36e};
test_input[9176:9183] = '{32'h40adda10, 32'h41fd94e2, 32'hc2be257c, 32'hc2c499cb, 32'h42078e73, 32'h41a0b554, 32'h420c9250, 32'hc13a9a71};
test_weights[9176:9183] = '{32'h40219512, 32'hc2c02a01, 32'h425dc095, 32'hc205e33c, 32'h4193887d, 32'hc23da2d8, 32'h4241dd0d, 32'h42c1634c};
test_bias[1147:1147] = '{32'hc1d29b0d};
test_output[1147:1147] = '{32'hc595b39f};
test_input[9184:9191] = '{32'hc147d5e3, 32'h412656f5, 32'h42232f67, 32'hc2905a7e, 32'h408e02ca, 32'hc28f9d2d, 32'hc0e69db6, 32'h4274b5da};
test_weights[9184:9191] = '{32'h42b59010, 32'h42881be4, 32'h42a62a1d, 32'hc2b3e56f, 32'hc2192085, 32'hc2b108e8, 32'h4222b904, 32'hc0a063f6};
test_bias[1148:1148] = '{32'h41b98941};
test_output[1148:1148] = '{32'h466b63c9};
test_input[9192:9199] = '{32'hc285f047, 32'h424e3529, 32'h42ae6f63, 32'h3fb8f884, 32'h429c3fb2, 32'h4142d4f3, 32'h40f2b28c, 32'hc2c09048};
test_weights[9192:9199] = '{32'h428fc3c2, 32'hc0e7fc35, 32'h42c60d42, 32'h42300dec, 32'hc19c77e6, 32'hc210e031, 32'h42af0f8f, 32'h41a17c41};
test_bias[1149:1149] = '{32'hc204be7e};
test_output[1149:1149] = '{32'h4366e228};
test_input[9200:9207] = '{32'hc2361be2, 32'hc2842544, 32'hc2a30db7, 32'h4218f849, 32'h41c73eaa, 32'hc295a810, 32'hc2799c1b, 32'h42c16ae8};
test_weights[9200:9207] = '{32'hc200b45a, 32'hc13ddb44, 32'hc1aa20bb, 32'hc1497eb7, 32'hc108912e, 32'h42b13d5a, 32'hc1d000ac, 32'h42164eb0};
test_bias[1150:1150] = '{32'hc286cf37};
test_output[1150:1150] = '{32'h44e6c992};
test_input[9208:9215] = '{32'hc285f83c, 32'h422c570a, 32'h42ad3d36, 32'h428f8e71, 32'hc168eeee, 32'h41515244, 32'h429c45e6, 32'hc19a6381};
test_weights[9208:9215] = '{32'hc1fc1ede, 32'h42b0daa0, 32'hc2616b8c, 32'h421f37d0, 32'h4206b319, 32'hc264a94d, 32'h4228118c, 32'h4001967c};
test_bias[1151:1151] = '{32'hc233b398};
test_output[1151:1151] = '{32'h45b70c12};
test_input[9216:9223] = '{32'hc1178aa2, 32'hc1d91904, 32'hc218a12f, 32'hc2655ba5, 32'h409aa325, 32'h42a58293, 32'h42008b1d, 32'hc1ceef3b};
test_weights[9216:9223] = '{32'hc29a72f8, 32'h40d91411, 32'h41948e24, 32'hc18f75f2, 32'h41a76426, 32'hc274d22d, 32'h42353f1d, 32'h4235fb83};
test_bias[1152:1152] = '{32'hc2ab7704};
test_output[1152:1152] = '{32'hc573f585};
test_input[9224:9231] = '{32'h41b6245c, 32'hc206b5ee, 32'h42569ad6, 32'hc249c8cc, 32'h42c4b474, 32'h42bd6e3d, 32'h42726c25, 32'hc28b4f7b};
test_weights[9224:9231] = '{32'hbfda7a44, 32'h4214d9c2, 32'h4226a518, 32'h42350c61, 32'hbfd7b1b7, 32'hc2a54aa5, 32'hc17b9eac, 32'hc2234311};
test_bias[1153:1153] = '{32'h41c74d77};
test_output[1153:1153] = '{32'hc5e7d792};
test_input[9232:9239] = '{32'hc27068f6, 32'h41816435, 32'hc242a221, 32'hc29127ce, 32'h42698399, 32'h414a186c, 32'hc2b534b7, 32'hc0124bc2};
test_weights[9232:9239] = '{32'h408e93e0, 32'h4228a899, 32'h4240bb64, 32'hc293e380, 32'hc2a7c7c0, 32'hc1c2345a, 32'hc281059b, 32'hc23b133f};
test_bias[1154:1154] = '{32'hc2625550};
test_output[1154:1154] = '{32'h4580fcb5};
test_input[9240:9247] = '{32'hc0910f6e, 32'h429c8320, 32'h41bdc8db, 32'hc22dc3e7, 32'hc20c2e63, 32'h42bdfeed, 32'hc1ec6930, 32'h42107dac};
test_weights[9240:9247] = '{32'h4246e668, 32'h42b0d4ed, 32'hc1e095ea, 32'h4195dc05, 32'hc1ac0790, 32'h42599fe4, 32'hc2207269, 32'h425e1822};
test_bias[1155:1155] = '{32'hc28025ef};
test_output[1155:1155] = '{32'h465edbc8};
test_input[9248:9255] = '{32'h424a55f0, 32'h414cb93c, 32'hc209a4fc, 32'hc2ad7c97, 32'h420b9e21, 32'hbe2110a9, 32'h3d4a03af, 32'hc1be2b6e};
test_weights[9248:9255] = '{32'hc243e8be, 32'hc26742ae, 32'h429b3c87, 32'h419e8071, 32'hc24cd973, 32'h4280b5f7, 32'hc14b57ad, 32'h428e380b};
test_bias[1156:1156] = '{32'hc2771978};
test_output[1156:1156] = '{32'hc62e54c3};
test_input[9256:9263] = '{32'h42016655, 32'hc29a698c, 32'hc24b131b, 32'hc1237bf2, 32'h4252b2dc, 32'h42b6b300, 32'h40782528, 32'h417dfe84};
test_weights[9256:9263] = '{32'h4299178f, 32'h4283fb8c, 32'h41382ecb, 32'hc28d6448, 32'h42a11c1a, 32'h42978e92, 32'h40e083d6, 32'h41acfeb0};
test_bias[1157:1157] = '{32'hc20500fb};
test_output[1157:1157] = '{32'h460cf818};
test_input[9264:9271] = '{32'hc2939f39, 32'hc2b5d477, 32'h426398f6, 32'h41a76061, 32'h42429ee4, 32'hc235af1d, 32'hc29ef305, 32'hc25531ea};
test_weights[9264:9271] = '{32'h40a5fab2, 32'h4205f3fd, 32'hc25cf591, 32'h41f9c445, 32'h429eead8, 32'h40d8cea7, 32'hc2211346, 32'h421619b3};
test_bias[1158:1158] = '{32'hc238f06f};
test_output[1158:1158] = '{32'hc4969d9c};
test_input[9272:9279] = '{32'h418e504b, 32'h4081f917, 32'hc21b68df, 32'h42aae75b, 32'h4297c1d7, 32'hc2628ae5, 32'h423e34b1, 32'h429cde60};
test_weights[9272:9279] = '{32'h42072292, 32'hc2217d39, 32'h41383b1f, 32'hc158fcb5, 32'h41bc150f, 32'hc01bf40c, 32'hc28637db, 32'h422a0472};
test_bias[1159:1159] = '{32'hc1dd3f6c};
test_output[1159:1159] = '{32'h4458edcd};
test_input[9280:9287] = '{32'hbf8993be, 32'hc2223bbf, 32'hc2431e78, 32'hc263e3f5, 32'h4282f055, 32'h41fec49d, 32'hc2a7a6ad, 32'h42a91282};
test_weights[9280:9287] = '{32'h415d7923, 32'hc214865f, 32'h429a0ed7, 32'h417e0d95, 32'hc017528d, 32'h42666fc5, 32'h42c64e92, 32'h4222e223};
test_bias[1160:1160] = '{32'hc2b24acc};
test_output[1160:1160] = '{32'hc5c98c18};
test_input[9288:9295] = '{32'hc20684c4, 32'hc29cdab4, 32'hc2a7080c, 32'hc2c43572, 32'hc1fabcf0, 32'h426b5d48, 32'h42a5a703, 32'h42815f90};
test_weights[9288:9295] = '{32'hc291afc4, 32'hc1ca22fd, 32'h42c01b91, 32'hc245bba2, 32'hc2c59998, 32'h42b5f20d, 32'h42a0f473, 32'h4261d7d7};
test_bias[1161:1161] = '{32'h422611d1};
test_output[1161:1161] = '{32'h469cc7cc};
test_input[9296:9303] = '{32'hc21a9338, 32'hc1f651d9, 32'h4260a035, 32'hc0d44ece, 32'hc243f6a8, 32'hc1a943a2, 32'hc2b5fb0b, 32'hc2a1c71f};
test_weights[9296:9303] = '{32'hc2123372, 32'hc2856484, 32'h429d84e3, 32'hc25fddc9, 32'hc24782f5, 32'hc2bfdd46, 32'hc2a44726, 32'hc28f3426};
test_bias[1162:1162] = '{32'hc1db50d3};
test_output[1162:1162] = '{32'h46cae770};
test_input[9304:9311] = '{32'h42a28481, 32'h42aea52c, 32'hc132cda3, 32'hc1582d79, 32'h428231a8, 32'hc2816e3f, 32'h41163693, 32'hc276cb0a};
test_weights[9304:9311] = '{32'h4290cdce, 32'h42a55a2b, 32'hc2639d19, 32'h4188b6f3, 32'hc1b52de8, 32'hc26a0cb1, 32'hc296807f, 32'hc18b1141};
test_bias[1163:1163] = '{32'hc22b0480};
test_output[1163:1163] = '{32'h467c3dda};
test_input[9312:9319] = '{32'h42317c34, 32'hc2929d9e, 32'h42b0cdb1, 32'h42857548, 32'h425a4add, 32'h42b34a23, 32'hc18c9005, 32'h4262d9ba};
test_weights[9312:9319] = '{32'h42a5c542, 32'hc288cf10, 32'h3f04b846, 32'h411ac595, 32'h42c5dffe, 32'hc26a66ce, 32'hc2b0fc47, 32'hc21ff127};
test_bias[1164:1164] = '{32'hc244a9c3};
test_output[1164:1164] = '{32'h4608fee8};
test_input[9320:9327] = '{32'hc1683fb3, 32'h420f5e1f, 32'h42bd252f, 32'h4212f115, 32'hc1f6b953, 32'hc27e84d0, 32'hc14b9295, 32'hc192b7f7};
test_weights[9320:9327] = '{32'h412436a2, 32'h41ecae67, 32'h4258b49f, 32'h4235b0eb, 32'h41a78d99, 32'hc2a1eb3e, 32'h42a75f9c, 32'hc1976ca0};
test_bias[1165:1165] = '{32'h41b9b723};
test_output[1165:1165] = '{32'h4633eae0};
test_input[9328:9335] = '{32'h42c7c9da, 32'h41fc2ce3, 32'h42ac3817, 32'h41d77aad, 32'h429d6fb0, 32'hc21aab07, 32'h42bd9a44, 32'hc299020b};
test_weights[9328:9335] = '{32'h40f72109, 32'h4196c353, 32'hc237cbe2, 32'hc2bb0324, 32'hc29337fd, 32'hc1e4af81, 32'hc162e523, 32'h3f832920};
test_bias[1166:1166] = '{32'h41f18de9};
test_output[1166:1166] = '{32'hc62edd7a};
test_input[9336:9343] = '{32'h40940700, 32'h420461a5, 32'h41809c7c, 32'h421f027c, 32'h41eaadbc, 32'h4242e856, 32'hc2b8238d, 32'hc0a106a9};
test_weights[9336:9343] = '{32'hc23cd1ae, 32'hc15991ec, 32'h429a8101, 32'h4248403c, 32'h40f7860b, 32'hc1d3b596, 32'h416f7f88, 32'hc1d3fe93};
test_bias[1167:1167] = '{32'h41c05a17};
test_output[1167:1167] = '{32'h438c26f0};
test_input[9344:9351] = '{32'hc21cfd05, 32'hc1ebcbc3, 32'h418485fe, 32'h423cea7f, 32'hc20fb812, 32'hc29f91de, 32'h42907335, 32'h41ea9184};
test_weights[9344:9351] = '{32'hc2a3f210, 32'h4275169a, 32'hc27b31ca, 32'hc28f64e7, 32'hc14d064f, 32'hc22be238, 32'hc0c9cb60, 32'h3fcafe30};
test_bias[1168:1168] = '{32'h4245b886};
test_output[1168:1168] = '{32'h4400849c};
test_input[9352:9359] = '{32'h42a6b7c1, 32'h423f31eb, 32'hc2406e9d, 32'hc0afbef5, 32'h4248a9fa, 32'h41c31be2, 32'hc2689f19, 32'hc2522882};
test_weights[9352:9359] = '{32'hc2689d82, 32'h428a8bfe, 32'hc2899777, 32'hc15e78ca, 32'hc2b9871b, 32'h42866e88, 32'hc1bea4db, 32'hc17c1630};
test_bias[1169:1169] = '{32'h4252e581};
test_output[1169:1169] = '{32'h4489b41d};
test_input[9360:9367] = '{32'hc26d8667, 32'h4187d0de, 32'h41cf717e, 32'hc2826d1e, 32'hc2bff02b, 32'h421f917c, 32'h4266b14a, 32'hbfb9bcc7};
test_weights[9360:9367] = '{32'hc2be921d, 32'hc1ee85a9, 32'h42b98a42, 32'h41f96001, 32'hc2458f7f, 32'h4297a955, 32'h4148d189, 32'h4225b97c};
test_bias[1170:1170] = '{32'h42649ea2};
test_output[1170:1170] = '{32'h465aea73};
test_input[9368:9375] = '{32'hc10fd0c6, 32'hc28e60ae, 32'hc24f2451, 32'hc20282ee, 32'h428f8663, 32'h4230585e, 32'hc29c4a19, 32'hc2b503db};
test_weights[9368:9375] = '{32'hc2aadc5b, 32'h42b8e1f0, 32'h42b673c0, 32'h426485e0, 32'hc20bf15d, 32'hc2248ae9, 32'hc29aadbe, 32'hc287159e};
test_bias[1171:1171] = '{32'h4106e052};
test_output[1171:1171] = '{32'hc58e8129};
test_input[9376:9383] = '{32'h42bb421e, 32'h428cba94, 32'h40d65ad2, 32'hc1939ef8, 32'hc1627e01, 32'hc2a52ac8, 32'h40841a6a, 32'hc0e4f05d};
test_weights[9376:9383] = '{32'hc1d59097, 32'hc1910058, 32'hc0d414a5, 32'h41cc27b9, 32'h41f37b6d, 32'hc2649584, 32'hc27c1bae, 32'hc26e77c9};
test_bias[1172:1172] = '{32'h413222e4};
test_output[1172:1172] = '{32'h432fcd89};
test_input[9384:9391] = '{32'hc29df17c, 32'h415711b0, 32'h41f305b4, 32'hc2ad6d80, 32'h429ed651, 32'hc28e2ec1, 32'hc23028c5, 32'hc2a218c0};
test_weights[9384:9391] = '{32'hc0b16f86, 32'hc299bd8e, 32'h427714ce, 32'h424b4d47, 32'h419ec805, 32'h422e30d3, 32'hc28b4446, 32'hc1c0a1dc};
test_bias[1173:1173] = '{32'hc23bfc32};
test_output[1173:1173] = '{32'h43a2b3d4};
test_input[9392:9399] = '{32'hc122e5ed, 32'h420323e8, 32'h42b15d25, 32'hc106e85b, 32'hc1a2b97d, 32'h42032e4a, 32'h411e7b67, 32'h429665ef};
test_weights[9392:9399] = '{32'hc2594677, 32'hc23f1fdd, 32'h413c9145, 32'hc299828f, 32'h41aa7102, 32'hc129b0b0, 32'h42aba8e4, 32'h4272bc6f};
test_bias[1174:1174] = '{32'hc18b361a};
test_output[1174:1174] = '{32'h45a56e8d};
test_input[9400:9407] = '{32'hc1c969a3, 32'hc210609d, 32'hc059b118, 32'hc2312fe2, 32'h4295123a, 32'hc231ade4, 32'hc19ff980, 32'h42c1d67d};
test_weights[9400:9407] = '{32'hc2934751, 32'h42a46320, 32'h4214d620, 32'hc281a66d, 32'h4272579e, 32'hc2b6a339, 32'hc28a83f9, 32'hc261dd65};
test_bias[1175:1175] = '{32'h40377332};
test_output[1175:1175] = '{32'h45bf3c50};
test_input[9408:9415] = '{32'h41016a4f, 32'h4225c796, 32'hc2ba8e17, 32'hc24f98a1, 32'h41bfb959, 32'h425aece1, 32'h429b4318, 32'h424f47c8};
test_weights[9408:9415] = '{32'h42165fd6, 32'h428f7e7e, 32'h4157bde7, 32'h42839b19, 32'h41060d07, 32'h42bd59f6, 32'hc28ac410, 32'h42a02cd8};
test_bias[1176:1176] = '{32'h425e5d08};
test_output[1176:1176] = '{32'h452f6c17};
test_input[9416:9423] = '{32'hc27a1f00, 32'hc2c7d3a6, 32'h42c207ae, 32'h42456096, 32'h428901cd, 32'h41caf321, 32'hc22ea836, 32'h41b4ccf7};
test_weights[9416:9423] = '{32'hc2961dc7, 32'hc28c9214, 32'hc299b5ba, 32'hc252c087, 32'h41be514c, 32'h426840ba, 32'h42a81dd6, 32'h429433eb};
test_bias[1177:1177] = '{32'h41d67f67};
test_output[1177:1177] = '{32'h452e9bf6};
test_input[9424:9431] = '{32'h411e6da7, 32'hc2b0c8bb, 32'h42bd1067, 32'h42a554fc, 32'h41a10a38, 32'h42b93c51, 32'h425997d5, 32'h4219a67c};
test_weights[9424:9431] = '{32'h4205efb2, 32'hc294954c, 32'hc234af85, 32'h4299ff13, 32'h4167c082, 32'h422184f1, 32'hc2bc5fcb, 32'hc1636441};
test_bias[1178:1178] = '{32'h426e00b4};
test_output[1178:1178] = '{32'h45e7b60a};
test_input[9432:9439] = '{32'h41e1b64c, 32'h42ac1886, 32'hc2803551, 32'hc1db0148, 32'h42a74bdb, 32'h421c5320, 32'hc20cfd09, 32'h42bb0625};
test_weights[9432:9439] = '{32'hc23d8164, 32'hc18c8ddc, 32'h42610671, 32'h42267792, 32'hc20c4b45, 32'h4286ad89, 32'hbe11b04f, 32'h40ed2375};
test_bias[1179:1179] = '{32'hc1976574};
test_output[1179:1179] = '{32'hc5e188d2};
test_input[9440:9447] = '{32'hc219d9c5, 32'h42b6b1c0, 32'hc28a8cd4, 32'hc2914b90, 32'h41869fc9, 32'hc0fb86d4, 32'h41e14450, 32'hc1b23f98};
test_weights[9440:9447] = '{32'hc2866ae0, 32'hc2be0a2e, 32'h41e234c4, 32'h40474234, 32'hc1fb1517, 32'h42c3abe8, 32'h428dbe37, 32'hc212c86d};
test_bias[1180:1180] = '{32'h41fce8f4};
test_output[1180:1180] = '{32'hc5d2607d};
test_input[9448:9455] = '{32'hbfdfdc16, 32'h42c7b19a, 32'h3e3458a1, 32'hc21551a1, 32'hc213d887, 32'h41dbf166, 32'h423f27ad, 32'h42422da5};
test_weights[9448:9455] = '{32'hc1933321, 32'h41dbd75f, 32'h425f5a6e, 32'hc1ccf759, 32'hc25c607d, 32'hc0b0fdea, 32'h42a9caf4, 32'hc19d62f8};
test_bias[1181:1181] = '{32'hc2a62188};
test_output[1181:1181] = '{32'h46071621};
test_input[9456:9463] = '{32'h4284331a, 32'h4248a8d5, 32'hc29a2b61, 32'h42317ba6, 32'h424d5b7b, 32'h42a945be, 32'hc180175f, 32'h41dbce24};
test_weights[9456:9463] = '{32'h42b87d1b, 32'h42795007, 32'hc2a02693, 32'hc1b5ca94, 32'hc1271b53, 32'h421b4722, 32'h41abc1ab, 32'h42c1f7ea};
test_bias[1182:1182] = '{32'hc23d792f};
test_output[1182:1182] = '{32'h4697a67b};
test_input[9464:9471] = '{32'h426f921b, 32'h421c48a3, 32'hc200989e, 32'h42549940, 32'hc280c65c, 32'h421233bf, 32'hc2adf4aa, 32'h429e1c2c};
test_weights[9464:9471] = '{32'h41997974, 32'hc27e90da, 32'h41f6a8be, 32'h4224fb66, 32'hc28be6cf, 32'hc28b7c78, 32'h418501ac, 32'hc2b01b80};
test_bias[1183:1183] = '{32'h41c29020};
test_output[1183:1183] = '{32'hc5cd24f8};
test_input[9472:9479] = '{32'h4258bdfd, 32'hc2ac8a23, 32'hc24e1e18, 32'hc206732c, 32'h4209d96d, 32'hc15a5da0, 32'hc1d21fe4, 32'hc2bf508a};
test_weights[9472:9479] = '{32'hc21f9854, 32'h423ce62f, 32'hc20839ca, 32'hc29d7878, 32'hc1dd75ec, 32'hc295cae9, 32'hc2454692, 32'hc2c2fe41};
test_bias[1184:1184] = '{32'hc2637d54};
test_output[1184:1184] = '{32'h46097954};
test_input[9480:9487] = '{32'h420d5097, 32'h42422565, 32'hc2852eec, 32'h4199ea19, 32'hc2b5b837, 32'h421a8a54, 32'hc0fd6dd0, 32'hc2413f8f};
test_weights[9480:9487] = '{32'hc29c6231, 32'h422d257f, 32'hc27f562e, 32'h4292e347, 32'hc1f18157, 32'hc20b52bc, 32'hc2a58b22, 32'h427e5deb};
test_bias[1185:1185] = '{32'h41d97d89};
test_output[1185:1185] = '{32'h457aa0f5};
test_input[9488:9495] = '{32'h4251f399, 32'hc2c4e647, 32'h42988814, 32'h427fae6a, 32'h424f8d38, 32'h42a8172b, 32'h42c11f05, 32'h42b1db28};
test_weights[9488:9495] = '{32'h42424b1d, 32'h3e110c5d, 32'hc2939cc3, 32'h420bc3dd, 32'h424e8f90, 32'hc249299f, 32'h42adc254, 32'hc2b47813};
test_bias[1186:1186] = '{32'hc09bdbae};
test_output[1186:1186] = '{32'hc4ffe50d};
test_input[9496:9503] = '{32'h42a73c8f, 32'hc2a1585c, 32'h41f5fc8b, 32'hc28b5e29, 32'h4243d43e, 32'h429f7255, 32'hc2709ee0, 32'h417cbdc6};
test_weights[9496:9503] = '{32'hc200bab5, 32'hc2392198, 32'h421cd089, 32'h4104fc10, 32'h429c7d87, 32'hc1f487fe, 32'h41968189, 32'h4236a09d};
test_bias[1187:1187] = '{32'h429c474e};
test_output[1187:1187] = '{32'h452aa707};
test_input[9504:9511] = '{32'hc293cf6a, 32'hc0178596, 32'hc22504de, 32'h42650529, 32'hc2754a0b, 32'h42755b1d, 32'hc23aae8f, 32'hc085af85};
test_weights[9504:9511] = '{32'h42633ce6, 32'h428957ad, 32'hc218519b, 32'hc1752745, 32'h42867105, 32'hc2b65719, 32'hc23b62fd, 32'h4205e15c};
test_bias[1188:1188] = '{32'hc23b02c2};
test_output[1188:1188] = '{32'hc631d81b};
test_input[9512:9519] = '{32'hc2843ad1, 32'h42bdb03f, 32'h42b350d6, 32'h40019a42, 32'hc26c7d1e, 32'hc25b5e8b, 32'h42c66b1f, 32'hc2b7277e};
test_weights[9512:9519] = '{32'hc1988616, 32'hc2bb19d2, 32'h422ca60a, 32'h4233ab22, 32'hc2416ef7, 32'h41b7141c, 32'hc113da36, 32'hc24ee5bb};
test_bias[1189:1189] = '{32'hc2a67b61};
test_output[1189:1189] = '{32'h44d32a97};
test_input[9520:9527] = '{32'h42b0abeb, 32'hc208e942, 32'h42267b6a, 32'hc287f029, 32'h420e35e5, 32'h40596325, 32'hc0b14b8f, 32'hc2a5b427};
test_weights[9520:9527] = '{32'hc2c37011, 32'h42b53fa1, 32'h41cb4ff7, 32'h41c0037a, 32'hc01e8184, 32'hc1bf81db, 32'hc26b24b5, 32'hc2bd0847};
test_bias[1190:1190] = '{32'h42034204};
test_output[1190:1190] = '{32'hc585fc9b};
test_input[9528:9535] = '{32'hc28b584c, 32'hc21e7db1, 32'hc2ad915e, 32'hc2060659, 32'h42022fcd, 32'h42895ec0, 32'h42928857, 32'h42b84bdf};
test_weights[9528:9535] = '{32'h41c3dfcf, 32'h42725c8c, 32'hc0da0110, 32'hc1de8e4c, 32'h42931ddf, 32'hc209d745, 32'hc00c7e73, 32'h418dbe6d};
test_bias[1191:1191] = '{32'h4290c8d5};
test_output[1191:1191] = '{32'hc47cf7c5};
test_input[9536:9543] = '{32'hc16cb168, 32'hc130b4de, 32'hc2303cae, 32'hc2a6f5c5, 32'h427197eb, 32'hc11381af, 32'h42b64174, 32'hc21db58a};
test_weights[9536:9543] = '{32'h4295ed86, 32'hc2a00bab, 32'hc22143fc, 32'hc196ad83, 32'hc2563aa0, 32'h42b76037, 32'h42601e32, 32'h41930f3b};
test_bias[1192:1192] = '{32'h42285dee};
test_output[1192:1192] = '{32'h4558a90c};
test_input[9544:9551] = '{32'hc1dd468e, 32'hc1e68df2, 32'hc1e6dfcf, 32'hc2997165, 32'hc1c2156a, 32'hc1db20ab, 32'h4108cbb0, 32'hc2b807dc};
test_weights[9544:9551] = '{32'h41a5575d, 32'hc295bacd, 32'hc2862006, 32'h429a4d71, 32'hc1f87f8c, 32'h4283e107, 32'h42af91d6, 32'h42a0a9d0};
test_bias[1193:1193] = '{32'h429f6f8c};
test_output[1193:1193] = '{32'hc61c6fbf};
test_input[9552:9559] = '{32'h427e3339, 32'h4122ab90, 32'h42bcf2a5, 32'hc2a49401, 32'hc24fdec4, 32'h42ac8913, 32'hc1a26772, 32'hc1e516ef};
test_weights[9552:9559] = '{32'hc276f5a7, 32'hc20b26d5, 32'h41dfeedb, 32'h416ab3f0, 32'h41a1ed5c, 32'hc295d7c2, 32'hc2026bf3, 32'hc22e1acd};
test_bias[1194:1194] = '{32'h416cfadb};
test_output[1194:1194] = '{32'hc603bf96};
test_input[9560:9567] = '{32'h42a1c82a, 32'h42644f2b, 32'h42aa933a, 32'h4271678d, 32'hc2653648, 32'h414f2706, 32'h429809e4, 32'h425cb1df};
test_weights[9560:9567] = '{32'hc28fbddd, 32'hc2363b5d, 32'hc210ee02, 32'hc1a88d30, 32'hc2871450, 32'hbfbdf66e, 32'h41e99b73, 32'hc29145fb};
test_bias[1195:1195] = '{32'h41663c11};
test_output[1195:1195] = '{32'hc627288b};
test_input[9568:9575] = '{32'hc1b4c6a5, 32'h42845648, 32'h4238b7b4, 32'hc27c8737, 32'hc1dc3c3f, 32'hc2407211, 32'hc20fe44e, 32'hc2bbf372};
test_weights[9568:9575] = '{32'h42815ab3, 32'hc2971a5f, 32'hc1f56984, 32'hc1a3ceac, 32'hc1f49c7b, 32'h42872591, 32'h41a158fb, 32'h428d04f8};
test_bias[1196:1196] = '{32'h42b6b481};
test_output[1196:1196] = '{32'hc67df8e6};
test_input[9576:9583] = '{32'h40d43052, 32'hc29be26d, 32'h42164be2, 32'h413199f3, 32'h420bad16, 32'hc24f6b52, 32'h419b6eb2, 32'hc288ac2b};
test_weights[9576:9583] = '{32'hbfcc996d, 32'hc2bfb8c5, 32'hc2b00863, 32'h41107e55, 32'hc29126a6, 32'h42470ad1, 32'hc2a76586, 32'h41fb6a06};
test_bias[1197:1197] = '{32'hc2ab7b5d};
test_output[1197:1197] = '{32'hc5937fd4};
test_input[9584:9591] = '{32'h42978937, 32'hc1c3035d, 32'hc1451811, 32'h421049af, 32'h41a56d11, 32'hc1b27475, 32'hc2313a5f, 32'h41677888};
test_weights[9584:9591] = '{32'hc20c1ec7, 32'hc242b491, 32'h42852048, 32'h42b97b12, 32'h40e7a255, 32'h42bece61, 32'hc2929fad, 32'h4199aed3};
test_bias[1198:1198] = '{32'hc269efd9};
test_output[1198:1198] = '{32'h451f2fbc};
test_input[9592:9599] = '{32'hc2842f7f, 32'h4214d2a2, 32'h423c4137, 32'hc28e6d79, 32'h40e1964d, 32'h4229d412, 32'h42ae31a2, 32'hc1b3ca6b};
test_weights[9592:9599] = '{32'h408f686a, 32'h3ffc8c9c, 32'h4129e3f1, 32'hc299a1ba, 32'h41a1d4ce, 32'hc00bc578, 32'hc2a2a067, 32'h4224ddc7};
test_bias[1199:1199] = '{32'hc285e43c};
test_output[1199:1199] = '{32'hc50e633c};
test_input[9600:9607] = '{32'hc1b8cfb0, 32'hc2a5ba9b, 32'hc2afe165, 32'hc2bc4a33, 32'hc2a07abe, 32'h40f4d510, 32'h429708aa, 32'h41c1ea1a};
test_weights[9600:9607] = '{32'hc27a54c9, 32'hc174bc45, 32'hc24f5cbf, 32'h428fd06c, 32'h40f7b193, 32'hc2998f97, 32'hc2b2f28a, 32'hc2ae5235};
test_bias[1200:1200] = '{32'h422e6e71};
test_output[1200:1200] = '{32'hc614eff8};
test_input[9608:9615] = '{32'h4219fda9, 32'hc2a8dd54, 32'hc1b13d9e, 32'h429414e4, 32'h42bc69d0, 32'hc2bb588d, 32'h41eb0de2, 32'h41de567d};
test_weights[9608:9615] = '{32'hc214a6a9, 32'h42a864de, 32'hc2659015, 32'h42892725, 32'hc27a996f, 32'hc26b0120, 32'hc27dc1bd, 32'h427a8b80};
test_bias[1201:1201] = '{32'hbdcedbf1};
test_output[1201:1201] = '{32'hc5298932};
test_input[9616:9623] = '{32'h423e2e08, 32'h428ca3c9, 32'hc18b7d9e, 32'hc2195e6a, 32'h42c497e2, 32'h42994488, 32'h42b61d70, 32'h421826e9};
test_weights[9616:9623] = '{32'hc232270f, 32'hbf8dcbc2, 32'h4282fc1a, 32'hc2b489de, 32'h41c35ab9, 32'h41804707, 32'h429083c0, 32'h41f013f7};
test_bias[1202:1202] = '{32'hc283331b};
test_output[1202:1202] = '{32'h46324150};
test_input[9624:9631] = '{32'hc11190d2, 32'hc24dcfdf, 32'h415c066b, 32'hc2853857, 32'h41c35feb, 32'h41d06de6, 32'h421ea822, 32'hc1a1f20d};
test_weights[9624:9631] = '{32'hc2450325, 32'h41c63275, 32'hc1cfdbc9, 32'hc26c0034, 32'h42bd06dd, 32'hc2b701a9, 32'hc1858d86, 32'h41c99ff2};
test_bias[1203:1203] = '{32'h42258e2e};
test_output[1203:1203] = '{32'h44c069fb};
test_input[9632:9639] = '{32'h42c532d1, 32'h42b78a5b, 32'h4213c83a, 32'hc2219b83, 32'h408e3403, 32'h4214f141, 32'hc2657dc6, 32'h427dccbb};
test_weights[9632:9639] = '{32'hc175f1a3, 32'hc2bd4ebe, 32'hc29a746c, 32'h428df5ea, 32'hc24b61e8, 32'hc13a6182, 32'h423d2a64, 32'hc2108e40};
test_bias[1204:1204] = '{32'h42c241bb};
test_output[1204:1204] = '{32'hc6a7e793};
test_input[9640:9647] = '{32'h427899ab, 32'h42bbd5d4, 32'h41c24748, 32'h41fe859c, 32'h42103ad3, 32'h4247e6db, 32'hc021f156, 32'hc2a17d3d};
test_weights[9640:9647] = '{32'h42045502, 32'hc29997b2, 32'hc2275684, 32'hc233e82f, 32'hc2b5c632, 32'h41c28dd3, 32'h4263cb87, 32'h419d96dc};
test_bias[1205:1205] = '{32'h42171b97};
test_output[1205:1205] = '{32'hc63187e9};
test_input[9648:9655] = '{32'h419a072f, 32'hc2c48a14, 32'hc1e45882, 32'hc2b9b95c, 32'hc26a2a14, 32'h418f6b5a, 32'hc1647c3b, 32'h42c59945};
test_weights[9648:9655] = '{32'hc0ac97e3, 32'h428069ff, 32'h42c488a8, 32'hc2134529, 32'hc2c05d19, 32'h42a017ec, 32'hc27c3c2e, 32'h41e5363c};
test_bias[1206:1206] = '{32'hc28a0fa9};
test_output[1206:1206] = '{32'h459a03e5};
test_input[9656:9663] = '{32'hc1a4973e, 32'h42bf4c5d, 32'hc2b902bd, 32'h41dcdb23, 32'hc18d93bd, 32'h42903a3a, 32'h41b6e3c1, 32'hc2033745};
test_weights[9656:9663] = '{32'hc29424aa, 32'h41902d58, 32'hc2c24efd, 32'h41d95950, 32'hc20d35b5, 32'h42533923, 32'h42322004, 32'h41cf036b};
test_bias[1207:1207] = '{32'hc2ab0b33};
test_output[1207:1207] = '{32'h4688bb04};
test_input[9664:9671] = '{32'hc1d599cd, 32'hc17af152, 32'hc28d70e1, 32'hc27abe61, 32'h42a602fe, 32'hc2ab1f3b, 32'hc22b89c6, 32'h41f1f2c6};
test_weights[9664:9671] = '{32'hc230a494, 32'h424a50a3, 32'hc2c240ff, 32'hc2939e8b, 32'h4299b87e, 32'hc2903371, 32'hc2ac50d9, 32'h40880e1d};
test_bias[1208:1208] = '{32'hc21176c0};
test_output[1208:1208] = '{32'h46dc72d7};
test_input[9672:9679] = '{32'hc1bdc6b5, 32'h41f24af2, 32'h413cc90f, 32'hc1ced14f, 32'h42bd7e2f, 32'hc2b20bf3, 32'h429b5bf9, 32'h4223c860};
test_weights[9672:9679] = '{32'h4288aa7c, 32'hc291236f, 32'h4258b5b3, 32'h4252f1c8, 32'hc22e967a, 32'h41d03034, 32'h42c5d3c7, 32'h42a6c90b};
test_bias[1209:1209] = '{32'hc2a7436a};
test_output[1209:1209] = '{32'h419b8eae};
test_input[9680:9687] = '{32'h426ceafc, 32'h4246c85c, 32'h428eee96, 32'h41cb4f38, 32'hc1d29e87, 32'h42841b20, 32'hc24d9bdc, 32'hc2a873c5};
test_weights[9680:9687] = '{32'h4282eb7e, 32'h423e540e, 32'h411c14dc, 32'hc2849f02, 32'hc2c51dd6, 32'hc20c8494, 32'h419b92f2, 32'h42b3dde2};
test_bias[1210:1210] = '{32'hc10d00a1};
test_output[1210:1210] = '{32'hc53ef091};
test_input[9688:9695] = '{32'h428fd46b, 32'hc1a26616, 32'h408656b6, 32'h415da83a, 32'h42aa792d, 32'h418be148, 32'hc290be4a, 32'hc07d646b};
test_weights[9688:9695] = '{32'hc2a18d99, 32'hc2b9abe5, 32'hc21c97eb, 32'h429ccde7, 32'h424a09a9, 32'h428f2b5a, 32'hc25c110d, 32'hc2350d25};
test_bias[1211:1211] = '{32'h42a5b19e};
test_output[1211:1211] = '{32'h45d46f72};
test_input[9696:9703] = '{32'h426efaa0, 32'h42bcfa6d, 32'hc1ef8a7e, 32'h427c4c4d, 32'h422780ed, 32'hc0b7542b, 32'h42342598, 32'hc16ddf8e};
test_weights[9696:9703] = '{32'hc280470d, 32'h42b8fac6, 32'hc0deef04, 32'hc2c13878, 32'h42862a39, 32'h3ff81332, 32'hc2bbdcc0, 32'h42b7cad9};
test_bias[1212:1212] = '{32'hc20e7135};
test_output[1212:1212] = '{32'hc56e3e03};
test_input[9704:9711] = '{32'hc296d05d, 32'h42899728, 32'h426ac823, 32'hc1ce4f90, 32'h428a3871, 32'hc2743ecc, 32'h422041fb, 32'hc2bae437};
test_weights[9704:9711] = '{32'hc250bbaf, 32'h42b67f08, 32'hc0fded7b, 32'h41ec33d8, 32'h42a10808, 32'hc1c9adf3, 32'hc1e46dc6, 32'h41233ada};
test_bias[1213:1213] = '{32'hc2ad6fda};
test_output[1213:1213] = '{32'h46594412};
test_input[9712:9719] = '{32'h4285333e, 32'h42baad1e, 32'hc11723cb, 32'h428efa1e, 32'h41ad1447, 32'hc2b80b71, 32'h429e0ecf, 32'h42a4f4a4};
test_weights[9712:9719] = '{32'hc20284a4, 32'h41c1e615, 32'h42ab29ac, 32'h4280f83e, 32'h412789d1, 32'hc24da1dd, 32'hc229d7bf, 32'h42a3bf04};
test_bias[1214:1214] = '{32'hc15d7011};
test_output[1214:1214] = '{32'h463f1c81};
test_input[9720:9727] = '{32'hbf16b8f3, 32'hc284dc3a, 32'hc272b754, 32'h41840a0f, 32'hbfbca725, 32'h4204ff8e, 32'h429b25c4, 32'h4269142d};
test_weights[9720:9727] = '{32'hc271825b, 32'hc2bb32f0, 32'hc2b7d689, 32'h42b0c57e, 32'h41cc604e, 32'h4239c922, 32'h42a706dc, 32'h428ff872};
test_bias[1215:1215] = '{32'h4243490e};
test_output[1215:1215] = '{32'h46c75c75};
test_input[9728:9735] = '{32'h3c5fa470, 32'hc0a044a0, 32'h428aaa7d, 32'h41184b20, 32'hc1222912, 32'hc26b89ef, 32'h4246ec2b, 32'h4141c280};
test_weights[9728:9735] = '{32'hc2a1280b, 32'hc233a3e3, 32'h423850e1, 32'hc256483b, 32'hc2a38002, 32'h42c1ef97, 32'hc2357d2c, 32'h40ddc4fc};
test_bias[1216:1216] = '{32'hc2b6bb9b};
test_output[1216:1216] = '{32'hc5846407};
test_input[9736:9743] = '{32'h41bb70dc, 32'h42a7db82, 32'hc1f73b09, 32'hc0ea6ffd, 32'h41230fd9, 32'h42539f2d, 32'h42907a50, 32'hc279884a};
test_weights[9736:9743] = '{32'h42b23b5f, 32'h429b9b33, 32'h42ac652d, 32'hc29fd124, 32'h42867010, 32'h408c1c3f, 32'hc13e6598, 32'hc281d124};
test_bias[1217:1217] = '{32'h4293914b};
test_output[1217:1217] = '{32'h46277e2d};
test_input[9744:9751] = '{32'h4195304d, 32'h42a653dd, 32'hc29efd17, 32'hc2604e00, 32'hc2bf0cef, 32'h41b8eca0, 32'h42af09ba, 32'h42a8612f};
test_weights[9744:9751] = '{32'hc11cf2dc, 32'hc2b209ee, 32'hc1ed370b, 32'h4254f6cc, 32'h40a16559, 32'h425bbd28, 32'hc290f472, 32'h42012fdc};
test_bias[1218:1218] = '{32'hc1c4580f};
test_output[1218:1218] = '{32'hc62d0c6b};
test_input[9752:9759] = '{32'hc1827423, 32'h42c2764b, 32'h428f8d4f, 32'hc2153a5c, 32'h42503baf, 32'h4142b785, 32'hc0a5e6ea, 32'hc2236811};
test_weights[9752:9759] = '{32'h425e682d, 32'hbf8cb8b5, 32'hc22985a2, 32'hc2af2a9b, 32'h420d8b69, 32'hc292fac2, 32'h42bc35ba, 32'h420f25d8};
test_bias[1219:1219] = '{32'hc22817a5};
test_output[1219:1219] = '{32'hc4e502bd};
test_input[9760:9767] = '{32'h424a4bd7, 32'hc24b6f97, 32'h420415dc, 32'h42c59bb4, 32'h412e0a7e, 32'h429620b1, 32'h4217c713, 32'hc1c6616e};
test_weights[9760:9767] = '{32'hc2892052, 32'h410a3b5f, 32'h42c7fde2, 32'h428c0c80, 32'hc23ba70f, 32'h411e6d36, 32'h408b5829, 32'hc2c34fae};
test_bias[1220:1220] = '{32'h422149bc};
test_output[1220:1220] = '{32'h460f57ab};
test_input[9768:9775] = '{32'h4256999e, 32'hc27fb646, 32'h415d5768, 32'h42bd9ae8, 32'hc28b1ee9, 32'h42167171, 32'hc269ef46, 32'hc0fedaf9};
test_weights[9768:9775] = '{32'hc2bb14f3, 32'h41da9587, 32'h4297e9ff, 32'hc29341c6, 32'hc1d467d5, 32'h4298fa07, 32'h418e1787, 32'hc2bdef67};
test_bias[1221:1221] = '{32'h4285ed6b};
test_output[1221:1221] = '{32'hc5ffd2d4};
test_input[9776:9783] = '{32'hc18b969c, 32'h4004d067, 32'h427c8b39, 32'h421ff4d8, 32'hc29044e8, 32'hc2ad0ca6, 32'hc190ccd2, 32'h428058a2};
test_weights[9776:9783] = '{32'h424649f0, 32'hc216a0fb, 32'h423267f3, 32'hc25bd6a4, 32'h41a0d85b, 32'hc0135a03, 32'h429dcf5f, 32'h42875493};
test_bias[1222:1222] = '{32'h42325b32};
test_output[1222:1222] = '{32'h44acd504};
test_input[9784:9791] = '{32'hc2be80a2, 32'hc270deca, 32'h42a1b50c, 32'h42c1ba9b, 32'h42507423, 32'h42b48121, 32'h42b3963a, 32'hc1e965fb};
test_weights[9784:9791] = '{32'hc2b5a1c5, 32'hc20af06a, 32'hc2a91db0, 32'h420f1d21, 32'h417716d4, 32'hc2ae86fc, 32'h41848a26, 32'hc227b7b6};
test_bias[1223:1223] = '{32'hc22256ff};
test_output[1223:1223] = '{32'h4539a381};
test_input[9792:9799] = '{32'h42743fe6, 32'h412632f2, 32'h42319977, 32'hc18c9584, 32'h42a4402d, 32'hc2974da9, 32'hc1dfb1b8, 32'hc26403ef};
test_weights[9792:9799] = '{32'h426fd9c1, 32'h41287a83, 32'h428f691f, 32'h42a17c49, 32'hc28a0394, 32'hc2b4ceaf, 32'hc2b0976d, 32'hc29a6195};
test_bias[1224:1224] = '{32'hc19ad311};
test_output[1224:1224] = '{32'h4653d559};
test_input[9800:9807] = '{32'h40979cd7, 32'hc2a93912, 32'hc19e9893, 32'hc2bdfde7, 32'hc28b750c, 32'hc28319e5, 32'hc1016604, 32'h42217ab1};
test_weights[9800:9807] = '{32'h427c4eda, 32'hc232697b, 32'hc2ba13d2, 32'h42077d41, 32'hc2967687, 32'hc18c94d4, 32'h41423831, 32'hc2205a81};
test_bias[1225:1225] = '{32'hc2481d3d};
test_output[1225:1225] = '{32'h45e514f3};
test_input[9808:9815] = '{32'hc2b8623e, 32'hc298159b, 32'hbfa6adba, 32'hbfc92e0d, 32'hc18f759a, 32'h40c3f91a, 32'hc1ef2ed1, 32'h4160e094};
test_weights[9808:9815] = '{32'h42797f99, 32'hc28a868d, 32'hc1f0b12d, 32'hc2576dd3, 32'hc24f75b9, 32'hc1de3c4b, 32'h424dd916, 32'h3fa18e39};
test_bias[1226:1226] = '{32'hc18ad799};
test_output[1226:1226] = '{32'hc48e3fb6};
test_input[9816:9823] = '{32'h42a47ef8, 32'hc20b520c, 32'h422a78d9, 32'hc219c91c, 32'hc1fb7da2, 32'h422dd688, 32'h4145af7b, 32'hc09a9a99};
test_weights[9816:9823] = '{32'h4101e003, 32'hc1b9f763, 32'hc25202f6, 32'hc1b3f0be, 32'hc25551dc, 32'h421a6a4f, 32'hc298ea17, 32'h428d2f2f};
test_bias[1227:1227] = '{32'hc2894a11};
test_output[1227:1227] = '{32'h450384f4};
test_input[9824:9831] = '{32'h42c7230a, 32'hc29666f7, 32'h42b0fa86, 32'hc2adb22d, 32'h3f8cdddd, 32'h41927e43, 32'h427e73f6, 32'h41b075c2};
test_weights[9824:9831] = '{32'h42728c10, 32'hc2b7d35c, 32'hc27e6bab, 32'h41a16562, 32'hc2813af3, 32'hc2bc0701, 32'h414b1ff7, 32'h42c500be};
test_bias[1228:1228] = '{32'h420f864a};
test_output[1228:1228] = '{32'h45d443cc};
test_input[9832:9839] = '{32'h41939a3f, 32'h4156dcff, 32'h41eb3d0f, 32'h425a9327, 32'h422c793f, 32'hc141da0a, 32'h42884006, 32'h424e3764};
test_weights[9832:9839] = '{32'hc2632e66, 32'hc02c2ecd, 32'hc1f848c9, 32'h41aa3990, 32'h41fe11a9, 32'h413a8f05, 32'h42c3aedd, 32'h425faf58};
test_bias[1229:1229] = '{32'hc2452f38};
test_output[1229:1229] = '{32'h461a9560};
test_input[9840:9847] = '{32'h4146a344, 32'hc20bf443, 32'h414b4578, 32'h41591a8e, 32'hc2bd566b, 32'hc21a66d3, 32'h40d02b81, 32'h40f21364};
test_weights[9840:9847] = '{32'h42bf0c3a, 32'hc161696d, 32'hc2b8aaf1, 32'hc29b9e5c, 32'h41820f14, 32'hc0d828d8, 32'hc2406113, 32'hc21df4e5};
test_bias[1230:1230] = '{32'hc14b0ca9};
test_output[1230:1230] = '{32'hc51949d5};
test_input[9848:9855] = '{32'h427d7001, 32'hc248d4d3, 32'h42a310d5, 32'hc2a65073, 32'hc282789a, 32'hc2adef6a, 32'hbf9e423b, 32'h41a918ff};
test_weights[9848:9855] = '{32'hc247da81, 32'hc1e74333, 32'hc039e9dd, 32'h4220d8ff, 32'h42bfc3ab, 32'h420e1cba, 32'hc22c288d, 32'h4205eb0a};
test_bias[1231:1231] = '{32'h42bcb770};
test_output[1231:1231] = '{32'hc65761ed};
test_input[9856:9863] = '{32'h428c444e, 32'h41adb59e, 32'hbf088abd, 32'h425f6f8b, 32'hc282de93, 32'h424ebbed, 32'hc2119b25, 32'hc1217d74};
test_weights[9856:9863] = '{32'h4204ee6b, 32'h406310e1, 32'hc2751f3e, 32'hc15d9fa1, 32'h40da7c66, 32'h41034451, 32'hc0a77960, 32'hc27a03a2};
test_bias[1232:1232] = '{32'hc2a5e075};
test_output[1232:1232] = '{32'h4514e684};
test_input[9864:9871] = '{32'hc0920c91, 32'h429f5855, 32'hc1e8390a, 32'hc2b5a87a, 32'h42238e88, 32'h4251b7fb, 32'hc170647b, 32'hc12172de};
test_weights[9864:9871] = '{32'hc1aa88c3, 32'hc1509019, 32'h42b67891, 32'hc25d6f89, 32'hc238255e, 32'hc2a83bf1, 32'h425355b4, 32'h42af3da8};
test_bias[1233:1233] = '{32'h42b29e27};
test_output[1233:1233] = '{32'hc5c95575};
test_input[9872:9879] = '{32'hc1b0b374, 32'h40848038, 32'hc297c350, 32'hc2849232, 32'hc269e4fe, 32'h42ad4c5b, 32'h40cbd61c, 32'h429551d4};
test_weights[9872:9879] = '{32'h4250dc77, 32'hc24b73c5, 32'hc2c3f0f3, 32'hc2a01eee, 32'h3fbb7a66, 32'hc29290ce, 32'hc26cb0bf, 32'h42861653};
test_bias[1234:1234] = '{32'h42b8fd77};
test_output[1234:1234] = '{32'h4616fa53};
test_input[9880:9887] = '{32'h4108fa19, 32'h41801d29, 32'hc2986986, 32'hc2b1eac0, 32'hc21bb7e7, 32'hc2be6500, 32'h4259f550, 32'h427d82e3};
test_weights[9880:9887] = '{32'hc2a13966, 32'h41fd90e3, 32'hc2667dfa, 32'h4290b814, 32'hc1a52a43, 32'h4242370e, 32'hc21c75d6, 32'h419b1183};
test_bias[1235:1235] = '{32'hc1bc6a8c};
test_output[1235:1235] = '{32'hc5d9e996};
test_input[9888:9895] = '{32'hc1330b82, 32'hc254755e, 32'h42a5b80e, 32'hc1ae8d86, 32'h428d133d, 32'hc11a394a, 32'h42a7a1c7, 32'hc2669221};
test_weights[9888:9895] = '{32'hc1959cb6, 32'hc1ad7df8, 32'hc25b8e65, 32'h42991db5, 32'hc2bf30d5, 32'h422e2973, 32'h4241687f, 32'h428dc1c8};
test_bias[1236:1236] = '{32'h425f3c25};
test_output[1236:1236] = '{32'hc63b7507};
test_input[9896:9903] = '{32'hc2aa1b89, 32'hc22f9e99, 32'hc28657ba, 32'hbc47fdc7, 32'hc2ab5bac, 32'h42a32ac8, 32'hc213b092, 32'h42ae4206};
test_weights[9896:9903] = '{32'hc274d0a8, 32'hc2566afb, 32'hc1a6ab90, 32'h4099aca0, 32'hc259a3ef, 32'h42c589f0, 32'hc2c2362f, 32'h416d1743};
test_bias[1237:1237] = '{32'h42b027ff};
test_output[1237:1237] = '{32'h46d0259a};
test_input[9904:9911] = '{32'h40421611, 32'hc2191d27, 32'hc23a6172, 32'h42c26707, 32'hc2743180, 32'hc285855f, 32'h42b68348, 32'hc296383a};
test_weights[9904:9911] = '{32'h40ecbf04, 32'hc2580484, 32'h41c4cf8b, 32'h4246d6c0, 32'hc1820de4, 32'hc23364c9, 32'hc2a901c8, 32'h42bd82d8};
test_bias[1238:1238] = '{32'hc1b43a55};
test_output[1238:1238] = '{32'hc59f0aca};
test_input[9912:9919] = '{32'h40c78643, 32'h41a44a16, 32'h421e7500, 32'hc2295333, 32'hc2159c26, 32'h42370588, 32'hc28d5cd1, 32'h423760bb};
test_weights[9912:9919] = '{32'hc1b7738a, 32'h4217cc20, 32'hc26e1eab, 32'hc25fa012, 32'hc1993f4c, 32'h42624280, 32'hc207a345, 32'h3fb88b67};
test_bias[1239:1239] = '{32'hc2b17983};
test_output[1239:1239] = '{32'h45c59ba5};
test_input[9920:9927] = '{32'h423ae3a3, 32'hc2af3065, 32'hc185d7fd, 32'hc2928a78, 32'hc2a9950e, 32'hc1ba7b62, 32'hc256772d, 32'hc25fe1db};
test_weights[9920:9927] = '{32'hc279c3c0, 32'hc27a8a2d, 32'hc2b05198, 32'h428ca70b, 32'hc19205d9, 32'hc081f461, 32'h419b9aa3, 32'hc21bd706};
test_bias[1240:1240] = '{32'hc237e5f5};
test_output[1240:1240] = '{32'h44cb29eb};
test_input[9928:9935] = '{32'hc2614202, 32'h4129fda3, 32'h412414e8, 32'hc2aa90a1, 32'hbfa6e022, 32'hc2a668ed, 32'h42b9dade, 32'h4294abea};
test_weights[9928:9935] = '{32'hc255225f, 32'h42b8ee97, 32'hc2b7335e, 32'hc2c3b796, 32'hc22f7cc0, 32'h3e6d3a0a, 32'hc118220d, 32'h41e70a8c};
test_bias[1241:1241] = '{32'h42220599};
test_output[1241:1241] = '{32'h4646ebd1};
test_input[9936:9943] = '{32'hc2486185, 32'h42c7dd35, 32'h425a4187, 32'h4289b6f8, 32'hc20c7de4, 32'hc1a1033e, 32'hc1f12591, 32'hc1656fb6};
test_weights[9936:9943] = '{32'h423f47ed, 32'hc21f3132, 32'h409f83d2, 32'hc2bbf978, 32'hc20365af, 32'h421a925c, 32'h41ed0e65, 32'hc2aba017};
test_bias[1242:1242] = '{32'hc2a57180};
test_output[1242:1242] = '{32'hc63a9713};
test_input[9944:9951] = '{32'hc23c6794, 32'hc25eaf08, 32'hc134b181, 32'hc2bc647b, 32'hc1e6c6c8, 32'h42b54438, 32'hc2884f61, 32'hc20850b1};
test_weights[9944:9951] = '{32'h42b24652, 32'h428d508b, 32'hc2b12e50, 32'hc1fad93e, 32'h42794096, 32'hc2c2cdc3, 32'hc28ccc45, 32'h42909280};
test_bias[1243:1243] = '{32'hc271b115};
test_output[1243:1243] = '{32'hc643c47f};
test_input[9952:9959] = '{32'h41fb2311, 32'h40293ee4, 32'hc22a1c12, 32'h41822cb0, 32'h4233a214, 32'hc29ff67d, 32'h421b04a7, 32'hc2c735ae};
test_weights[9952:9959] = '{32'h422a96f8, 32'hc236da0c, 32'h41e60702, 32'h41addee2, 32'h423061ee, 32'h428a9783, 32'hc22442d5, 32'hc29ee8fa};
test_bias[1244:1244] = '{32'h42b7ee29};
test_output[1244:1244] = '{32'h4548139c};
test_input[9960:9967] = '{32'h413a0058, 32'hc25b1a47, 32'h42af7c51, 32'hc2b90f15, 32'hc24f13c3, 32'hc28adb66, 32'hc2b57457, 32'hc2b769c7};
test_weights[9960:9967] = '{32'h422ad87a, 32'hc097b6be, 32'hbf024dac, 32'hc248b599, 32'hc1c93590, 32'hc1c8c3ff, 32'hc2877da7, 32'hc2a83dd9};
test_bias[1245:1245] = '{32'hc2af3fd9};
test_output[1245:1245] = '{32'h46ad3808};
test_input[9968:9975] = '{32'hc27606f9, 32'hc0a4d8b0, 32'h421a97f2, 32'hc22ccdc5, 32'h42466639, 32'hc10cd40f, 32'h42859338, 32'h3f4cc65d};
test_weights[9968:9975] = '{32'hc21c2b1f, 32'h40db6f78, 32'h4298740e, 32'hc2054d80, 32'hc1fc1d89, 32'hc2b7f327, 32'h4164a8e7, 32'h41dafd9e};
test_bias[1246:1246] = '{32'hc2c4d76f};
test_output[1246:1246] = '{32'h45d6e13a};
test_input[9976:9983] = '{32'h42300d82, 32'h3f24b5b6, 32'hc289c85c, 32'h41df3f73, 32'hc211a23b, 32'h42427dc8, 32'hc2a636a7, 32'hc1bfdd1a};
test_weights[9976:9983] = '{32'h41f8b9b2, 32'h42480acf, 32'h42975097, 32'h42ac7bce, 32'h426060f0, 32'hc0a953fa, 32'h42c31e13, 32'h41269deb};
test_bias[1247:1247] = '{32'h4200ffb7};
test_output[1247:1247] = '{32'hc63bf72d};
test_input[9984:9991] = '{32'hc254430e, 32'h42a25e99, 32'h42c1fb8c, 32'hc290b8ec, 32'h40baeda2, 32'h42068b75, 32'h41aeee12, 32'h421dbad5};
test_weights[9984:9991] = '{32'hc15c369f, 32'hc1f8ff2a, 32'hc1334253, 32'hc29b250f, 32'hc181bd4f, 32'hc24d5c5b, 32'hc21ad152, 32'h401bff8e};
test_bias[1248:1248] = '{32'hbecf9b7b};
test_output[1248:1248] = '{32'h431dd9bb};
test_input[9992:9999] = '{32'hc1b59296, 32'h428f8be4, 32'hc2440ac0, 32'hc2c218fb, 32'hc0dd6a4a, 32'h418e0265, 32'h4182ae3f, 32'hc2c7e2d7};
test_weights[9992:9999] = '{32'h41caf95e, 32'hc1ad16f7, 32'hc277bbe0, 32'hc2a5247a, 32'hc22aedce, 32'hbf9ce088, 32'h425964fe, 32'h418560cf};
test_bias[1249:1249] = '{32'h42c330d1};
test_output[1249:1249] = '{32'h46050468};
test_input[10000:10007] = '{32'h420b5777, 32'hc2605b3a, 32'hc0cd2bbc, 32'h40f56732, 32'h42934e3c, 32'hc1a685c9, 32'h42c227ca, 32'h427f8b9a};
test_weights[10000:10007] = '{32'h42b1542b, 32'hc2274858, 32'hc254be05, 32'hc1b1b5ab, 32'h42b96e27, 32'hc22b1cc1, 32'h418a6a01, 32'hc2a428b7};
test_bias[1250:1250] = '{32'h412303df};
test_output[1250:1250] = '{32'h4618a8d5};
test_input[10008:10015] = '{32'hc2bd13c2, 32'hc1707efb, 32'hc2833dec, 32'h41c1eeaf, 32'hc230d2c0, 32'h426686a3, 32'h42aa703f, 32'hc1f02f58};
test_weights[10008:10015] = '{32'hc20a6b43, 32'hc233ef20, 32'hc284ad2f, 32'h41e92f59, 32'h3d8a91eb, 32'hc2c7ad49, 32'hc2bcab54, 32'hc241cece};
test_bias[1251:1251] = '{32'h426b55a4};
test_output[1251:1251] = '{32'hc54cb08e};
test_input[10016:10023] = '{32'h427c25c7, 32'h41a97f90, 32'h42b32f3c, 32'h42a4e0fe, 32'h426295be, 32'hc1c064e7, 32'h41bdc36f, 32'hc00b7e82};
test_weights[10016:10023] = '{32'hc25d7d76, 32'h41fb5b8d, 32'h42828969, 32'hc218d404, 32'h427ef7d7, 32'h4256bb57, 32'hc2492ebb, 32'hc2b640a4};
test_bias[1252:1252] = '{32'h428f365c};
test_output[1252:1252] = '{32'h449ebb92};
test_input[10024:10031] = '{32'hc2a31944, 32'h40b761d5, 32'h4201c2a8, 32'h41af2ac9, 32'h416104f5, 32'h415c8dd8, 32'h42129b26, 32'h4222f836};
test_weights[10024:10031] = '{32'h42396959, 32'hc29cd340, 32'h41fdf1a1, 32'h4230e02d, 32'hc18b8819, 32'h42097e1b, 32'hc2c1e16e, 32'hc1600311};
test_bias[1253:1253] = '{32'hc2bf1367};
test_output[1253:1253] = '{32'hc5c26f1a};
test_input[10032:10039] = '{32'h41b4a897, 32'hc26ef286, 32'h4210d4d3, 32'hc09d380f, 32'h429d4a53, 32'h426cf61a, 32'h41b0f63b, 32'hc287c51e};
test_weights[10032:10039] = '{32'h425bb7ce, 32'h425ecae4, 32'hc25171a5, 32'h42b1b74e, 32'h42bd031b, 32'h42ad4252, 32'h4239cb8c, 32'h42123a9b};
test_bias[1254:1254] = '{32'h42813f89};
test_output[1254:1254] = '{32'h45d31c7e};
test_input[10040:10047] = '{32'hc0b8bdc7, 32'hc232bc3e, 32'hc1ee1207, 32'hc1003ea1, 32'h42b6ff0f, 32'hc2117427, 32'hc1caf5f8, 32'hc0417ce2};
test_weights[10040:10047] = '{32'h41280db9, 32'hc258ce8c, 32'hc20bf709, 32'hc25514ff, 32'hc1dedadd, 32'hc26d3cba, 32'hc0310b0e, 32'h42a085d7};
test_bias[1255:1255] = '{32'h417eeed3};
test_output[1255:1255] = '{32'h454d0e18};
test_input[10048:10055] = '{32'hc224151c, 32'hc2909537, 32'h427bc4f8, 32'h41246a13, 32'h42aa3fea, 32'h420491c0, 32'hc2bc0538, 32'hc231d27f};
test_weights[10048:10055] = '{32'h40159f28, 32'h42662c68, 32'hc14ee891, 32'hc185a54e, 32'hc28067df, 32'h4130be2f, 32'h42b0f86c, 32'hc261bc20};
test_bias[1256:1256] = '{32'hc1cbbdc4};
test_output[1256:1256] = '{32'hc67cbf04};
test_input[10056:10063] = '{32'h429d80f0, 32'h42a398ba, 32'hc28610e6, 32'hc1487be4, 32'h428a10b7, 32'h424e6133, 32'h41e568f1, 32'h420062f5};
test_weights[10056:10063] = '{32'hc280f8d6, 32'h41dc33c9, 32'hc261c946, 32'h41075803, 32'h4223af32, 32'h41cd89b0, 32'hc2958ecc, 32'h40acea5a};
test_bias[1257:1257] = '{32'h42c44a3e};
test_output[1257:1257] = '{32'h454389a8};
test_input[10064:10071] = '{32'h42b5be0f, 32'hc2b5684a, 32'hc11bf5fc, 32'hc27ed1c1, 32'hc23c947e, 32'h4272ea91, 32'h4220e5d4, 32'h420f423f};
test_weights[10064:10071] = '{32'hc19b304d, 32'hc2be0e6f, 32'hc1272639, 32'hc263687f, 32'hc22dfeb0, 32'hc298ce41, 32'hc0e46d60, 32'hc2be2489};
test_bias[1258:1258] = '{32'h423519a9};
test_output[1258:1258] = '{32'h4587c23a};
test_input[10072:10079] = '{32'hc1ec40a2, 32'hc28629ba, 32'h418e88d3, 32'hc2c5aad2, 32'h42904964, 32'h4197221c, 32'hc2837932, 32'h426f6bdb};
test_weights[10072:10079] = '{32'hc1cdb8ee, 32'h4286d437, 32'h40c881ef, 32'hc1bf94b0, 32'hc2c21d0f, 32'hc10d0a68, 32'h4281b3e8, 32'h411fa9ac};
test_bias[1259:1259] = '{32'h4262700d};
test_output[1259:1259] = '{32'hc63c7884};
test_input[10080:10087] = '{32'hc1d88983, 32'hc277a597, 32'h42030294, 32'hc2b6e6f4, 32'h42a30fc6, 32'h428877cb, 32'h4245a402, 32'h429b0b99};
test_weights[10080:10087] = '{32'hc270a38f, 32'hc186c483, 32'h40b9b1c7, 32'hc26b7fb9, 32'hc1822bcc, 32'hc282f8ad, 32'h42ba4adc, 32'hc0aa8b28};
test_bias[1260:1260] = '{32'hc16e76c5};
test_output[1260:1260] = '{32'h45cf06fd};
test_input[10088:10095] = '{32'hc27cf753, 32'h420bdf90, 32'hc2afc867, 32'hc272f91a, 32'h42877053, 32'h41931164, 32'hc10202ab, 32'hc147f031};
test_weights[10088:10095] = '{32'h421f3de7, 32'hc22950b8, 32'hc1b2b578, 32'h421160ba, 32'hc219384a, 32'hc2339cad, 32'h42055525, 32'h42bf82d2};
test_bias[1261:1261] = '{32'hc251a170};
test_output[1261:1261] = '{32'hc60f75cc};
test_input[10096:10103] = '{32'h42990a45, 32'hc2922007, 32'h427eaf0a, 32'hc19400d1, 32'h42b3acd6, 32'h419412e7, 32'h41d6b9c9, 32'hc196085b};
test_weights[10096:10103] = '{32'h40185e93, 32'h42b253b1, 32'h423eb267, 32'hc2a92548, 32'hc29957d5, 32'hc27cce0a, 32'h42a3ff2a, 32'hc239f88b};
test_bias[1262:1262] = '{32'h429e1c64};
test_output[1262:1262] = '{32'hc5cf7139};
test_input[10104:10111] = '{32'h414649e2, 32'h40e47578, 32'h427b2a3c, 32'hc2a97cd5, 32'h42aa56fd, 32'h4198f321, 32'h41a2a351, 32'hc288879f};
test_weights[10104:10111] = '{32'h42646f8a, 32'h428f29b1, 32'h40c2ffd1, 32'h41aafdf9, 32'hc2c4e02c, 32'h42169e09, 32'h408e8ae9, 32'h4219f864};
test_bias[1263:1263] = '{32'hc2befbc0};
test_output[1263:1263] = '{32'hc6242a31};
test_input[10112:10119] = '{32'hc2a1e2bb, 32'h42bb0c84, 32'hc2aecb9d, 32'h41d12527, 32'h42c7b9a0, 32'h42ae37f7, 32'h4299b679, 32'hc219276e};
test_weights[10112:10119] = '{32'hc1a1f4fe, 32'h427e46de, 32'hc216a892, 32'hc27c60da, 32'hc253806e, 32'h42c7aba0, 32'hc1c156d9, 32'h41c660ea};
test_bias[1264:1264] = '{32'hc2a66220};
test_output[1264:1264] = '{32'h461861ea};
test_input[10120:10127] = '{32'hc2145070, 32'hc2ac7bf8, 32'hc26d8bd0, 32'hc222efc1, 32'h40e403cf, 32'hc1f916b4, 32'hc1d527e9, 32'hc203fd1c};
test_weights[10120:10127] = '{32'hc27a7801, 32'h429238a5, 32'hc1d24414, 32'hc0ead7ad, 32'hc23c2978, 32'hc2c3f4aa, 32'hc21ccefd, 32'hc28ac45b};
test_bias[1265:1265] = '{32'hc0c49043};
test_output[1265:1265] = '{32'h4574fa64};
test_input[10128:10135] = '{32'h40ca54ee, 32'hc1914355, 32'h40b542fa, 32'hc2a9be7d, 32'h427df0f4, 32'h423ac152, 32'hc29a5c57, 32'hc19af630};
test_weights[10128:10135] = '{32'hc1367952, 32'h4287b3eb, 32'h42a81434, 32'h42b7d660, 32'h42871c51, 32'hc235348e, 32'hc1ee7e68, 32'h3f88d297};
test_bias[1266:1266] = '{32'hc25faad7};
test_output[1266:1266] = '{32'hc5843bd3};
test_input[10136:10143] = '{32'h42082eca, 32'h41e27454, 32'hc2b630d2, 32'hc2a6b001, 32'hc275a190, 32'hc27e807e, 32'h413724d9, 32'h41c76826};
test_weights[10136:10143] = '{32'hc28cc8cd, 32'h40e93a03, 32'h41547d1b, 32'h4264bc1f, 32'h42405f62, 32'hc23bb1a7, 32'hc2b612f8, 32'hc2a9bcec};
test_bias[1267:1267] = '{32'h41e68db7};
test_output[1267:1267] = '{32'hc62ff97f};
test_input[10144:10151] = '{32'hc28709fa, 32'hc2bdfede, 32'h42aa5179, 32'h426796eb, 32'h4289a6bf, 32'hc2156a66, 32'h429c9524, 32'hc21e8a1d};
test_weights[10144:10151] = '{32'h426b8e0e, 32'hc2b1c7cb, 32'hc2805fd4, 32'h42bb7799, 32'h41b0d3ac, 32'h42b9071a, 32'h420af9ad, 32'h41d810ab};
test_bias[1268:1268] = '{32'hc1ec7d09};
test_output[1268:1268] = '{32'h45809574};
test_input[10152:10159] = '{32'hc193f1d1, 32'hc222c34a, 32'h42a5c65b, 32'hc1380063, 32'hc283d65f, 32'h41bc7d55, 32'h4251f20e, 32'h42be81e4};
test_weights[10152:10159] = '{32'h42b77a99, 32'h41efe84f, 32'hc2a0ccec, 32'hc2a8d91a, 32'h42b3d651, 32'h418ee05a, 32'hc22bc753, 32'hc200bf01};
test_bias[1269:1269] = '{32'hc296d394};
test_output[1269:1269] = '{32'hc6986fd2};
test_input[10160:10167] = '{32'h423813ab, 32'hc2894078, 32'h4219b26d, 32'hc180c9db, 32'hc2b17f4f, 32'h42adc4cc, 32'h4230e62e, 32'h415c5140};
test_weights[10160:10167] = '{32'h42b70668, 32'h4180130c, 32'hc2356b7e, 32'h41ba2bfa, 32'h42c3f871, 32'h41ed1b68, 32'h42be2103, 32'hc2b8d7ca};
test_bias[1270:1270] = '{32'h428703df};
test_output[1270:1270] = '{32'hc504e8c6};
test_input[10168:10175] = '{32'hc28e8140, 32'h4295c98e, 32'hc2958927, 32'h428101cb, 32'h4281b608, 32'hc197a4d7, 32'h42a04234, 32'h426de0a5};
test_weights[10168:10175] = '{32'hc25be50e, 32'hc12278ce, 32'h42b17aeb, 32'hc256884f, 32'hc2984ba0, 32'h4296db1b, 32'h42c4331c, 32'hc2a968b6};
test_bias[1271:1271] = '{32'hc2460552};
test_output[1271:1271] = '{32'hc62491d8};
test_input[10176:10183] = '{32'hc2a1aad2, 32'h42bcfa94, 32'h41b429d0, 32'hc22aceae, 32'hc21b7610, 32'h421f151c, 32'h42b72bce, 32'h41204dae};
test_weights[10176:10183] = '{32'h42939b8b, 32'h426a8178, 32'h42aa222e, 32'hc1dbb818, 32'hc29b76e8, 32'h4161f39b, 32'h41a3704c, 32'h42351b56};
test_bias[1272:1272] = '{32'hc299c647};
test_output[1272:1272] = '{32'h4604b352};
test_input[10184:10191] = '{32'h42495369, 32'hc25471ca, 32'h418a93d8, 32'h414ca060, 32'hc1eccf92, 32'hc1a460e2, 32'h42400dc1, 32'hc18e2ccc};
test_weights[10184:10191] = '{32'hbffbd571, 32'hc1cff05b, 32'h413178c9, 32'h426764ef, 32'hc2025f96, 32'h42a266c6, 32'hc2adcad6, 32'hc284ca61};
test_bias[1273:1273] = '{32'hc2c74679};
test_output[1273:1273] = '{32'hc4c5c243};
test_input[10192:10199] = '{32'h42b894cb, 32'h428fda45, 32'h42986390, 32'h40bc694e, 32'h42b99966, 32'h429d88ae, 32'h3e64f0e5, 32'h411bc9c5};
test_weights[10192:10199] = '{32'h4252f413, 32'h40b6e080, 32'h4065f069, 32'hc24cbfd0, 32'hc2c06883, 32'h427786c3, 32'hc1a5515c, 32'hc1831562};
test_bias[1274:1274] = '{32'h429d91a3};
test_output[1274:1274] = '{32'h448afa31};
test_input[10200:10207] = '{32'hc0af7acb, 32'h42b8feaf, 32'hc22d895f, 32'hc2444f2b, 32'hc16a8540, 32'hc2487151, 32'hc29f0109, 32'hc296b728};
test_weights[10200:10207] = '{32'hc2656e9f, 32'hc2a17faf, 32'hc2ae8624, 32'h429c716a, 32'h42b184c6, 32'hc20e1b8b, 32'hc2afd124, 32'h42b2fa8e};
test_bias[1275:1275] = '{32'hc1af913a};
test_output[1275:1275] = '{32'hc5cb494e};
test_input[10208:10215] = '{32'hc2828b4b, 32'h42ac1c62, 32'h42bd4df9, 32'h4040cd48, 32'h42c0f713, 32'hc154cbae, 32'hc14e146f, 32'h42c1ce06};
test_weights[10208:10215] = '{32'h413146a9, 32'h429fc9a4, 32'hc2489706, 32'h408baa62, 32'h42a4e98d, 32'hc2aacae1, 32'h42515637, 32'h41d7ea89};
test_bias[1276:1276] = '{32'h421a3d8d};
test_output[1276:1276] = '{32'h46432763};
test_input[10216:10223] = '{32'hbf2dc703, 32'hc28aa085, 32'hc1978d47, 32'h429a4c30, 32'h4125390f, 32'h426bd700, 32'h40ce0bb4, 32'h4297c22f};
test_weights[10216:10223] = '{32'hc26e7d71, 32'h4232fe57, 32'h429fa190, 32'hc1ad8c59, 32'h426e83b7, 32'h4212cc63, 32'hc21474ac, 32'hc20f362c};
test_bias[1277:1277] = '{32'hc2aed8eb};
test_output[1277:1277] = '{32'hc5cb7318};
test_input[10224:10231] = '{32'h42b8802e, 32'hc249402e, 32'hc2549fb4, 32'hc20fb19f, 32'hc2106e8f, 32'h4296a0ba, 32'hc2b5d64c, 32'h427d18d3};
test_weights[10224:10231] = '{32'hc212cc9f, 32'hc24242a1, 32'hc182ffea, 32'h42aba0e3, 32'h4115d6e1, 32'h414338d0, 32'hc0a9fd9c, 32'hc2051c2c};
test_bias[1278:1278] = '{32'hc222c991};
test_output[1278:1278] = '{32'hc58467f6};
test_input[10232:10239] = '{32'h40d25db1, 32'hc267cbb1, 32'h40357202, 32'hc2972d0d, 32'h428d69bd, 32'hbfc626eb, 32'h42ad25f2, 32'hc2be9aa4};
test_weights[10232:10239] = '{32'h41c11068, 32'hc29d68dc, 32'h42a2cf31, 32'hc21b5f25, 32'hc2a8c087, 32'hc2834249, 32'hc2b1bf00, 32'h429758f9};
test_bias[1279:1279] = '{32'hc1b6223c};
test_output[1279:1279] = '{32'hc649aae0};
test_input[10240:10247] = '{32'h41e0a88b, 32'h42b950bc, 32'hc04dc177, 32'h422311a0, 32'h40c698c1, 32'h421e1e6d, 32'hc1d57983, 32'h41d5035d};
test_weights[10240:10247] = '{32'hc212b08f, 32'h42717e5f, 32'h425535fd, 32'h42745f19, 32'hc2410dc4, 32'hc2ae7710, 32'hc26a50cf, 32'hc26ed1b5};
test_bias[1280:1280] = '{32'hc130f37a};
test_output[1280:1280] = '{32'h45419f85};
test_input[10248:10255] = '{32'hc1d383c1, 32'h4280d708, 32'h42886ab7, 32'hc25d98e0, 32'hc28dec4d, 32'hc2c4cf62, 32'h42835aab, 32'hc22f5c43};
test_weights[10248:10255] = '{32'hc282c431, 32'hc2c69082, 32'h428b4cbb, 32'h423781cd, 32'h42727fa9, 32'hc22e4f21, 32'h426f2548, 32'h42c459c3};
test_bias[1281:1281] = '{32'hc2814610};
test_output[1281:1281] = '{32'hc5361c16};
test_input[10256:10263] = '{32'h429857f3, 32'hc2392b20, 32'h41b79fe9, 32'hc2c5eb5b, 32'hc26d7512, 32'hc21384ae, 32'hc2550662, 32'hc2b21be7};
test_weights[10256:10263] = '{32'hc29692fa, 32'hc181d47e, 32'h3ed78e9b, 32'h42a563a2, 32'h4270c8b6, 32'h429fd8f0, 32'h428acd5a, 32'h4291ea9a};
test_bias[1282:1282] = '{32'hc1322ea0};
test_output[1282:1282] = '{32'hc6e97577};
test_input[10264:10271] = '{32'hc293c21f, 32'hc1e975c5, 32'hc1c05174, 32'hbfba55fc, 32'hc282c9b9, 32'hc2a43407, 32'hc2b7c9aa, 32'h4152b003};
test_weights[10264:10271] = '{32'h423003f6, 32'hc289b1a0, 32'h41e48841, 32'h42a6a045, 32'h421eaf50, 32'hc23befb7, 32'h422c2e7b, 32'h41e4a0b2};
test_bias[1283:1283] = '{32'hc2b22ee3};
test_output[1283:1283] = '{32'hc58b3833};
test_input[10272:10279] = '{32'h4292e5bf, 32'hc15e4e76, 32'hc153f074, 32'h42277783, 32'hbff8ff1d, 32'h41b95586, 32'hc1ffebb2, 32'h41816982};
test_weights[10272:10279] = '{32'h42b309ea, 32'h421356c2, 32'h4122927e, 32'hc29268dc, 32'hc04f1d4a, 32'h40ae0b1e, 32'hc2802c63, 32'h426d4f6a};
test_bias[1284:1284] = '{32'hc1bf32c8};
test_output[1284:1284] = '{32'h45baf0dc};
test_input[10280:10287] = '{32'h42bb1c44, 32'hc2828bf3, 32'h42b3ffe3, 32'hc121e71a, 32'h4223ba3c, 32'h427e54a0, 32'h426b1f5d, 32'hc254ba4e};
test_weights[10280:10287] = '{32'hc19e8300, 32'hc2b92c98, 32'hc2471d18, 32'h402761dd, 32'hc1e5a142, 32'hc0d3bedf, 32'hc28ccb09, 32'hc284ae93};
test_bias[1285:1285] = '{32'h420550ef};
test_output[1285:1285] = '{32'hc51b8da1};
test_input[10288:10295] = '{32'h42c3ab71, 32'hc2baa013, 32'hc1b10ee9, 32'h4265f708, 32'hc279041e, 32'hc20bacca, 32'h42c3df2d, 32'hc28febac};
test_weights[10288:10295] = '{32'hc24d3693, 32'hc1c36cb0, 32'hc233d1e6, 32'h42106775, 32'h42c16e54, 32'hc0448341, 32'hc2648030, 32'hc1ab9558};
test_bias[1286:1286] = '{32'hc22d0165};
test_output[1286:1286] = '{32'hc6173614};
test_input[10296:10303] = '{32'hc1d326ee, 32'h423ca17c, 32'h429786e6, 32'hc0425191, 32'h42953517, 32'h41741f2a, 32'h4205c766, 32'h41e2b91f};
test_weights[10296:10303] = '{32'hc10901fa, 32'h42a3a7e1, 32'h4099f34f, 32'hc2725b9d, 32'h429f8cdd, 32'h42b43c67, 32'hc1ef3172, 32'hc27a5d18};
test_bias[1287:1287] = '{32'h42770e16};
test_output[1287:1287] = '{32'h46107eee};
test_input[10304:10311] = '{32'hc2aa95e0, 32'h428e988b, 32'hc1a9f6d3, 32'h40a9960b, 32'hc0a340d9, 32'hc28fb470, 32'hc1b99804, 32'hc2c6f456};
test_weights[10304:10311] = '{32'h41d874e2, 32'h429d133f, 32'h4240253d, 32'hc2a3078a, 32'hc2bc9ad8, 32'h407c65b6, 32'h42331f3b, 32'hc132dea2};
test_bias[1288:1288] = '{32'h42156147};
test_output[1288:1288] = '{32'h450638b4};
test_input[10312:10319] = '{32'hc241848e, 32'hc2816119, 32'h427c3858, 32'h42ae177f, 32'h42660a99, 32'hc230e77b, 32'hc2a69730, 32'hc175276f};
test_weights[10312:10319] = '{32'hc25167ae, 32'h414c6634, 32'hc26e9953, 32'h42c75455, 32'h4299adb3, 32'hc20b030a, 32'h42617359, 32'hc221e7cf};
test_bias[1289:1289] = '{32'h42a3ef27};
test_output[1289:1289] = '{32'h46061fd1};
test_input[10320:10327] = '{32'h403b9df9, 32'hc21d880a, 32'hc1e51895, 32'hc29d064b, 32'h41fbdcbe, 32'h423a454e, 32'h42abd91e, 32'h42a38c4e};
test_weights[10320:10327] = '{32'hc17923c9, 32'hc09f2428, 32'h42860a2c, 32'h415acb9c, 32'hc2b1107c, 32'hc24e8c79, 32'h423cd5a0, 32'hc1699800};
test_bias[1290:1290] = '{32'hc292990f};
test_output[1290:1290] = '{32'hc5a3eac6};
test_input[10328:10335] = '{32'h4288d6eb, 32'hc1998335, 32'hc2800542, 32'hc10bae56, 32'h41c86a2a, 32'hc2bef4f4, 32'hc2215471, 32'hc183bd77};
test_weights[10328:10335] = '{32'h42a615e3, 32'hc204224a, 32'hc23bd935, 32'hc2ae1e4e, 32'hc2a2d894, 32'h41b24e0e, 32'hc22b4c40, 32'hc2b7e1ed};
test_bias[1291:1291] = '{32'h41104bfd};
test_output[1291:1291] = '{32'h460f30be};
test_input[10336:10343] = '{32'h3efde597, 32'h42908cfe, 32'hc15ff9b6, 32'hc1a07737, 32'h420eec83, 32'h426dbd32, 32'h419950ae, 32'hc285e2b3};
test_weights[10336:10343] = '{32'h4286153c, 32'h418b7d00, 32'hc17fc03e, 32'h41a7fb90, 32'hc297ec76, 32'hc249aaf9, 32'h41e7e236, 32'h42c6f08a};
test_bias[1292:1292] = '{32'h421428c0};
test_output[1292:1292] = '{32'hc626e3c9};
test_input[10344:10351] = '{32'hc17e44db, 32'hc2c263f0, 32'hc2bba519, 32'hc2653b16, 32'h429704df, 32'h429b5377, 32'hc2751f13, 32'h41be25f5};
test_weights[10344:10351] = '{32'hc1e9d87e, 32'hc1e710f2, 32'hc11e41c1, 32'hc2c3114b, 32'h3e8e3597, 32'h41563218, 32'hc04b24a5, 32'h42532ea9};
test_bias[1293:1293] = '{32'hc2b07ee4};
test_output[1293:1293] = '{32'h463ecc57};
test_input[10352:10359] = '{32'hc2399f03, 32'hc28d82d0, 32'hc21689a4, 32'h422e8b66, 32'hc2c30b94, 32'hbeef41b5, 32'hc2b228e5, 32'h41931bbc};
test_weights[10352:10359] = '{32'hc1d6a082, 32'h4299c21c, 32'h41af02bb, 32'hc2984c89, 32'hc128fc4c, 32'h42163d85, 32'h42505035, 32'h4257c5fd};
test_bias[1294:1294] = '{32'hc21d55d5};
test_output[1294:1294] = '{32'hc62c1b96};
test_input[10360:10367] = '{32'h411981ed, 32'h419fc2aa, 32'hbe2efc9e, 32'h42b0ee53, 32'h412559ff, 32'h42910e15, 32'h422d6764, 32'hc195ffdf};
test_weights[10360:10367] = '{32'h42282372, 32'h41a1c1f6, 32'h4064b2ae, 32'hc29b55d7, 32'h418b81ac, 32'h413289e1, 32'h42baad32, 32'h4268a0e8};
test_bias[1295:1295] = '{32'h427d2dbb};
test_output[1295:1295] = '{32'hc5007c1d};
test_input[10368:10375] = '{32'hc28e300e, 32'hc15f324c, 32'hc1c4c8df, 32'h41382ec5, 32'h421dc361, 32'h42a62c3f, 32'hc272d540, 32'hc2a9b1d1};
test_weights[10368:10375] = '{32'hc2c5ebb0, 32'h42a327e7, 32'h42a3506f, 32'h42bebc1d, 32'h42882b4a, 32'hc29f6d3a, 32'hc2758a3b, 32'hc1fd4907};
test_bias[1296:1296] = '{32'hc2711e18};
test_output[1296:1296] = '{32'h45e74c1e};
test_input[10376:10383] = '{32'hc1c8f7f9, 32'hc2a3eda8, 32'hc1916f4f, 32'h42a4c1a0, 32'hc2bb06c5, 32'hc26fe68c, 32'hc28bf40c, 32'h425f099d};
test_weights[10376:10383] = '{32'h419221e0, 32'h4298cbc2, 32'h427e192a, 32'hc2846c8e, 32'h4195a8c0, 32'hc20f21af, 32'h429a2383, 32'h42264842};
test_bias[1297:1297] = '{32'hbd9dfba4};
test_output[1297:1297] = '{32'hc67a2215};
test_input[10384:10391] = '{32'hc204912c, 32'h41bc8136, 32'h41396f4f, 32'h41daef65, 32'hc15dcbe3, 32'h41af127f, 32'hc0a38535, 32'h425d8e44};
test_weights[10384:10391] = '{32'h42c78bc3, 32'h40f17c11, 32'h400ef077, 32'h42b1ebbe, 32'h40a4a1d6, 32'h4237fccb, 32'h41b3f4d3, 32'hc1b2f845};
test_bias[1298:1298] = '{32'hc19fe752};
test_output[1298:1298] = '{32'hc48a64fd};
test_input[10392:10399] = '{32'hc20c9431, 32'hc2667094, 32'hc2327225, 32'h4298dbc9, 32'h429c2ebb, 32'h42a5148f, 32'hc274c60a, 32'hc234d890};
test_weights[10392:10399] = '{32'h425909f8, 32'hc28a106f, 32'h42727b15, 32'h42895447, 32'h41477939, 32'hc2a39339, 32'h3fb1291b, 32'h4247778e};
test_bias[1299:1299] = '{32'h3f2ad261};
test_output[1299:1299] = '{32'hc55ae246};
test_input[10400:10407] = '{32'h41968957, 32'hc266bc17, 32'hc182090b, 32'hc2a9a465, 32'hc251e152, 32'hc08ed004, 32'h421c4db1, 32'h425c8943};
test_weights[10400:10407] = '{32'hc242f659, 32'hc27bc5b4, 32'hc2bd636c, 32'hc23011f4, 32'h42180845, 32'hc2544ddc, 32'h40886272, 32'hc289fb55};
test_bias[1300:1300] = '{32'hc241ecd9};
test_output[1300:1300] = '{32'h451ef594};
test_input[10408:10415] = '{32'hc23664eb, 32'hc2098510, 32'h4280f87e, 32'h41a40a56, 32'hc2ace068, 32'hc22de075, 32'hc28864d9, 32'h41fe9c67};
test_weights[10408:10415] = '{32'h42bcbd38, 32'h428d94d0, 32'h423593f1, 32'hc29138a5, 32'hc16f75cd, 32'hc257fa5d, 32'h41699235, 32'h41c4a4bd};
test_bias[1301:1301] = '{32'h42827891};
test_output[1301:1301] = '{32'hc4e1b837};
test_input[10416:10423] = '{32'h42bb00a1, 32'hc1e9087b, 32'hc2b8eb4b, 32'hc28fef5c, 32'hc25db808, 32'h4275f0c6, 32'hc1b65871, 32'h416c6003};
test_weights[10416:10423] = '{32'hc0e1bda6, 32'hc1e68da6, 32'h406b7079, 32'hc1be77d2, 32'h4259eb58, 32'hc2921f8b, 32'hc2a5573e, 32'h40d5b1df};
test_bias[1302:1302] = '{32'hc2c70c16};
test_output[1302:1302] = '{32'hc57eb5d0};
test_input[10424:10431] = '{32'hc2209d43, 32'hc1e9aea4, 32'h42bcaeb6, 32'hc2087103, 32'hc1cb1bc9, 32'h41dde6a9, 32'h4129e541, 32'hc2b968a3};
test_weights[10424:10431] = '{32'hc2174080, 32'h426b9ea1, 32'hc18b32bf, 32'h421c7cfa, 32'hc2a5e131, 32'h42a1de0b, 32'hc270d2f1, 32'hc1c63586};
test_bias[1303:1303] = '{32'hc2af2e30};
test_output[1303:1303] = '{32'h452b650e};
test_input[10432:10439] = '{32'h42b25344, 32'h42994fbc, 32'hc23c3bb9, 32'h42611603, 32'h41867979, 32'h428057bb, 32'h41cc0dcc, 32'hc287b3fd};
test_weights[10432:10439] = '{32'h42828c1c, 32'hc28a5ca3, 32'h427e1466, 32'h42b21cf0, 32'h41e74e09, 32'hc20c2b87, 32'h42a0bced, 32'h42b59402};
test_bias[1304:1304] = '{32'h42223298};
test_output[1304:1304] = '{32'hc54dd55d};
test_input[10440:10447] = '{32'hc1ee7f4d, 32'h41953af1, 32'h424434ba, 32'hc1feb919, 32'hc1885c8f, 32'hc2a720ec, 32'h421c442a, 32'hc2464c1c};
test_weights[10440:10447] = '{32'hc058dfe2, 32'h41f3221c, 32'h4240891d, 32'hc09f1d97, 32'h41db2c81, 32'h4103f7d3, 32'h42236058, 32'hc0046156};
test_bias[1305:1305] = '{32'hc2c0cf46};
test_output[1305:1305] = '{32'h45630db9};
test_input[10448:10455] = '{32'h3f724af1, 32'h42967425, 32'hc11c6b2f, 32'hc20e78d4, 32'h421df5ae, 32'hc2009de9, 32'h4133758f, 32'h42264a4e};
test_weights[10448:10455] = '{32'h42a7ad71, 32'h4253c658, 32'h41190aec, 32'h40894596, 32'hc28b8438, 32'h4202ab27, 32'h422f29db, 32'hc2442580};
test_bias[1306:1306] = '{32'h42c43113};
test_output[1306:1306] = '{32'hc4b3d3a7};
test_input[10456:10463] = '{32'h40d4984e, 32'hc22b022a, 32'h417c9682, 32'h4255f3a5, 32'hc166e8b0, 32'hc2336fe4, 32'h4107bdeb, 32'h4202a0fb};
test_weights[10456:10463] = '{32'hc2a2e6a6, 32'h4298a338, 32'h42942ffd, 32'hc209df0c, 32'h42b967e1, 32'h4224b8f8, 32'hc2a0133e, 32'hc26e4181};
test_bias[1307:1307] = '{32'hc23a2c36};
test_output[1307:1307] = '{32'hc621772e};
test_input[10464:10471] = '{32'h420c3b9a, 32'hc2829139, 32'hc28a47d3, 32'hc261d53f, 32'h41bbd569, 32'h410c8a80, 32'hc22ff607, 32'h42acd3eb};
test_weights[10464:10471] = '{32'hc1a7ee38, 32'hc0fde9fd, 32'hc2339780, 32'h3e981015, 32'h42ab4457, 32'hc2afebe4, 32'hc22c55a2, 32'h3ff67137};
test_bias[1308:1308] = '{32'h42ae2390};
test_output[1308:1308] = '{32'h45c3821d};
test_input[10472:10479] = '{32'h422bdc53, 32'h42500814, 32'hc234a540, 32'hc1c5fa5a, 32'hc257977a, 32'hc271c992, 32'hc1e1a3f5, 32'h4135823b};
test_weights[10472:10479] = '{32'hc1dfac0a, 32'hc16cbe85, 32'h4160fadb, 32'hc0c5abb3, 32'h42a045b9, 32'h3ffb03d8, 32'hc29571c2, 32'hc1a1dd13};
test_bias[1309:1309] = '{32'hc1b03eb7};
test_output[1309:1309] = '{32'hc59d5579};
test_input[10480:10487] = '{32'h42a109b5, 32'h41a4f2d6, 32'hc1b18373, 32'h4283766d, 32'h427d1cbe, 32'hc29f2b81, 32'hc2afd5c9, 32'h418d8fe7};
test_weights[10480:10487] = '{32'h42bbff3d, 32'h4287b63c, 32'hc2bed7f9, 32'h41e3665c, 32'h42b89fd6, 32'h42600060, 32'hc1869d27, 32'hc0404413};
test_bias[1310:1310] = '{32'hc2788599};
test_output[1310:1310] = '{32'h4675587e};
test_input[10488:10495] = '{32'hc216183f, 32'h421d5767, 32'h419ba58b, 32'hc1fd1334, 32'h4285e4f8, 32'hc1c6d541, 32'h428ed4fb, 32'h429bcbf3};
test_weights[10488:10495] = '{32'h42706667, 32'hc28c85c7, 32'hc0bfb6f0, 32'hc2b0c70a, 32'h421e1138, 32'h42358e8e, 32'h41f80684, 32'h4109387e};
test_bias[1311:1311] = '{32'hc2ad3c43};
test_output[1311:1311] = '{32'h44f6b4d4};
test_input[10496:10503] = '{32'h41a1fa91, 32'h42c07121, 32'h420ff5a3, 32'hc2c2c8dd, 32'hc2aeafde, 32'h3f781917, 32'h427631ff, 32'hc201e50a};
test_weights[10496:10503] = '{32'h42942b6a, 32'hc2199b16, 32'hc1b4163d, 32'hc256e45f, 32'hc2baa927, 32'h42a6cee8, 32'h41de8dbf, 32'hc2c67d7f};
test_bias[1312:1312] = '{32'h41eb03f9};
test_output[1312:1312] = '{32'h46710092};
test_input[10504:10511] = '{32'h425727fd, 32'hc0d568e3, 32'hc2a71973, 32'h40324433, 32'hc2bf4b6b, 32'h427c9314, 32'hc2c393ec, 32'hc1866989};
test_weights[10504:10511] = '{32'h42a05bb5, 32'h3f283549, 32'hc1c1e846, 32'hc1d0a203, 32'h42a2756a, 32'h423e1551, 32'hc29615e7, 32'h40d5adf8};
test_bias[1313:1313] = '{32'h42640c44};
test_output[1313:1313] = '{32'h46091d2b};
test_input[10512:10519] = '{32'h420fad73, 32'hc17c82b1, 32'h40c6e7ad, 32'h4257ad70, 32'hc27f7d8c, 32'h42920a05, 32'h41532093, 32'h42980508};
test_weights[10512:10519] = '{32'hc18cc555, 32'h4267918d, 32'h40002020, 32'hc2643b73, 32'h42a6d675, 32'h42638057, 32'hc0e50c9b, 32'hc2a532f5};
test_bias[1314:1314] = '{32'hc212a46d};
test_output[1314:1314] = '{32'hc63e89c6};
test_input[10520:10527] = '{32'h4241fce5, 32'hc2666c85, 32'hc2aa354e, 32'h4215da84, 32'hc1d84114, 32'hc2b563c8, 32'h42a603c6, 32'h425f8f76};
test_weights[10520:10527] = '{32'hc0ea1a98, 32'hc243a8d8, 32'hbff5dd19, 32'hc099f1bc, 32'hc2ab0f32, 32'h41141a22, 32'hc18ba009, 32'hc1b45ef7};
test_bias[1315:1315] = '{32'h42bd6543};
test_output[1315:1315] = '{32'h44a312f1};
test_input[10528:10535] = '{32'hc1c5bdbc, 32'h4252040e, 32'hc21d6670, 32'hc19688d4, 32'hc28f4cd8, 32'h419457bd, 32'hc265a400, 32'h42ad8242};
test_weights[10528:10535] = '{32'h4235a656, 32'h428c67fc, 32'hc2afd070, 32'h3ee9b31f, 32'h41d773fb, 32'hc1324136, 32'hc1bed616, 32'h42b302b2};
test_bias[1316:1316] = '{32'h421f5911};
test_output[1316:1316] = '{32'h464bf050};
test_input[10536:10543] = '{32'hc2b91d41, 32'hc1a95764, 32'h42b3d1a8, 32'h42a7b41f, 32'h426a31bc, 32'h428b86bb, 32'hc2a030b1, 32'h42962eb7};
test_weights[10536:10543] = '{32'h40fb2480, 32'h4254eb7d, 32'hbf0eceeb, 32'h425c5087, 32'h4267d95d, 32'hc235bc20, 32'hc14f3bd9, 32'h4260bc03};
test_bias[1317:1317] = '{32'hc286783f};
test_output[1317:1317] = '{32'h45fe0194};
test_input[10544:10551] = '{32'h419d3455, 32'h420bab29, 32'hc273215a, 32'h419d5512, 32'h41654bb5, 32'h429b62b0, 32'h414469ff, 32'hc1b8ff71};
test_weights[10544:10551] = '{32'hc1fa27d6, 32'h41eb3607, 32'h41e2ad83, 32'hc2b02606, 32'hc04a72e3, 32'h428f8057, 32'h41ffa128, 32'h42b1414e};
test_bias[1318:1318] = '{32'h405ad299};
test_output[1318:1318] = '{32'h44504913};
test_input[10552:10559] = '{32'hc297d19b, 32'h42183a00, 32'h406cc928, 32'hc204861c, 32'hc2ac0a2f, 32'hc185f9ac, 32'hc2b685af, 32'hc1233c98};
test_weights[10552:10559] = '{32'h41a5d970, 32'hc2b32fbb, 32'hc2a37a39, 32'h41c90ea4, 32'hc1d0a9c4, 32'hc25291cc, 32'hc136f1b9, 32'hc119d0d0};
test_bias[1319:1319] = '{32'h421d826b};
test_output[1319:1319] = '{32'hc4e2862a};
test_input[10560:10567] = '{32'h420fe626, 32'h417e5079, 32'h427b2373, 32'h41c0de9c, 32'h41ae2dee, 32'h4114e71a, 32'hc2baefb7, 32'h4214f8ee};
test_weights[10560:10567] = '{32'h421e5f57, 32'h413517f5, 32'hc1ff9d9f, 32'h42a4dc0b, 32'hc1290405, 32'h42889ba2, 32'h42a941dc, 32'hc0e723a4};
test_bias[1320:1320] = '{32'h4208a404};
test_output[1320:1320] = '{32'hc5c04e9e};
test_input[10568:10575] = '{32'h413e507a, 32'hc18f3838, 32'h4223b384, 32'h428b933a, 32'h4272e297, 32'hc282f8fd, 32'h41ea1679, 32'h4182608d};
test_weights[10568:10575] = '{32'h4134322d, 32'hc27ac649, 32'hc19f3e27, 32'h409ee306, 32'hc0b9c8b9, 32'h41993042, 32'h425915f2, 32'h4107d966};
test_bias[1321:1321] = '{32'h42bd402b};
test_output[1321:1321] = '{32'h447aaf4a};
test_input[10576:10583] = '{32'h4182a8cc, 32'h427e99e6, 32'h42983060, 32'h4277ddb2, 32'hc1800477, 32'h4121c60a, 32'h428abf4e, 32'h42c0ae4f};
test_weights[10576:10583] = '{32'h42287caa, 32'h41957c0a, 32'hc270d301, 32'hc088957a, 32'h41fad0f7, 32'hc1d7c243, 32'hc1a64076, 32'h4255d620};
test_bias[1322:1322] = '{32'h4166e4ae};
test_output[1322:1322] = '{32'hc19f53a8};
test_input[10584:10591] = '{32'hc216ab22, 32'hc20c9dd3, 32'hc0eab477, 32'h419fd194, 32'hc1193e40, 32'h42959faf, 32'h42838144, 32'hc28470f1};
test_weights[10584:10591] = '{32'hc2abfecb, 32'hc1c9805b, 32'h429cce70, 32'hc122c76b, 32'hc2bcb604, 32'h41d78343, 32'h425c48bb, 32'hc009039a};
test_bias[1323:1323] = '{32'h42941725};
test_output[1323:1323] = '{32'h461dd988};
test_input[10592:10599] = '{32'hc26eb26c, 32'h426e6f9e, 32'hc1d692a8, 32'h42041ebf, 32'hc0a885c8, 32'hc2853e1b, 32'h42b0b059, 32'h42654136};
test_weights[10592:10599] = '{32'h416fe041, 32'hc29716b9, 32'h428e4252, 32'h41dba704, 32'hc044e8f4, 32'h41ae024f, 32'hc29dcb89, 32'h429af56d};
test_bias[1324:1324] = '{32'hc0f0fb42};
test_output[1324:1324] = '{32'hc6220290};
test_input[10600:10607] = '{32'h415dad6d, 32'hc289c8ca, 32'hc286bf2a, 32'hc242f332, 32'h42851f9e, 32'hc2827dd6, 32'hc2abf5ad, 32'hc219bcb1};
test_weights[10600:10607] = '{32'hc236e951, 32'h4298339c, 32'hc19a7dc0, 32'h4233c625, 32'hc09fde0f, 32'hc2640294, 32'h41b0cd30, 32'h40a0ddd2};
test_bias[1325:1325] = '{32'h4242eb69};
test_output[1325:1325] = '{32'hc5a97d62};
test_input[10608:10615] = '{32'hc29e6ad5, 32'h42c34cd8, 32'hc201e349, 32'h424c3739, 32'hc2bba023, 32'hc22d16a3, 32'h42a3a6bf, 32'h423cd326};
test_weights[10608:10615] = '{32'hc231562c, 32'h42b5fb1c, 32'h420a21d0, 32'hc06d1e1c, 32'hc24a2bfc, 32'hc28d4f1b, 32'h428ec229, 32'h42a5897f};
test_bias[1326:1326] = '{32'h4159a27b};
test_output[1326:1326] = '{32'h46dfcd82};
test_input[10616:10623] = '{32'h41ec58a5, 32'h416a6a35, 32'hc25dc6e9, 32'h42a017b9, 32'h42a671d5, 32'h4154c8b9, 32'hbfee2447, 32'h41677694};
test_weights[10616:10623] = '{32'hc2ab9565, 32'hbe26ab96, 32'h3dc5020c, 32'h42a88be2, 32'h4257799c, 32'hc22db56e, 32'hc285c229, 32'hc28ae313};
test_bias[1327:1327] = '{32'h422f679f};
test_output[1327:1327] = '{32'h45e34590};
test_input[10624:10631] = '{32'h411b6714, 32'h425bece7, 32'h40cd13e0, 32'hc2ae72b9, 32'h420e25a9, 32'h41cb1058, 32'h426a94f5, 32'h4214092f};
test_weights[10624:10631] = '{32'h42bd2447, 32'h42c59f62, 32'hc27ab2f7, 32'h4296f716, 32'h419988d4, 32'h4268f607, 32'hc22db19f, 32'h429d69e0};
test_bias[1328:1328] = '{32'hc25af7b6};
test_output[1328:1328] = '{32'h44e5b35c};
test_input[10632:10639] = '{32'h40306aae, 32'h4277b54a, 32'hc26cfc86, 32'h4265036c, 32'hc28ddf87, 32'hc1dbb63c, 32'hc2540718, 32'h41ccfaf5};
test_weights[10632:10639] = '{32'h42c283c3, 32'h42a3f492, 32'hc273e2b7, 32'hc1bcddfa, 32'hc0dfbf48, 32'hc2b65b2b, 32'h42bd8e23, 32'hc2ab8321};
test_bias[1329:1329] = '{32'h41f9cea3};
test_output[1329:1329] = '{32'h45557973};
test_input[10640:10647] = '{32'h4261a63e, 32'h41ec731f, 32'h422c3602, 32'h42c6aa5d, 32'h42a0f508, 32'hc24b0d58, 32'hc247bd09, 32'hc215707d};
test_weights[10640:10647] = '{32'h422a0966, 32'h42747eb4, 32'hc22c5ae0, 32'hc289088b, 32'h4288d738, 32'hc28ec73a, 32'h4215705d, 32'h424ec45a};
test_bias[1330:1330] = '{32'h42934261};
test_output[1330:1330] = '{32'h446db1ea};
test_input[10648:10655] = '{32'hc15b2394, 32'hc2c7e864, 32'hc20928c1, 32'hc25bec52, 32'hc2a2cba4, 32'hc2504793, 32'hc1fcfdf9, 32'h42b58b08};
test_weights[10648:10655] = '{32'h41654573, 32'hc1ecb070, 32'h41c6b47b, 32'hc2755229, 32'hc23be318, 32'h42a48814, 32'h42627a78, 32'h41477577};
test_bias[1331:1331] = '{32'h411bd633};
test_output[1331:1331] = '{32'h45825f10};
test_input[10656:10663] = '{32'hc2c31be3, 32'h4204e93e, 32'h42916450, 32'h40adc61d, 32'hc2b82ce6, 32'hc2a1fc48, 32'hc14edb75, 32'hc25bbe51};
test_weights[10656:10663] = '{32'hc2a536f3, 32'hc21c38f0, 32'h40d1257d, 32'hc181751b, 32'hc2c68b70, 32'hc24c79e5, 32'h42b17210, 32'hc20f6bdc};
test_bias[1332:1332] = '{32'hc1f97740};
test_output[1332:1332] = '{32'h46a5cb89};
test_input[10664:10671] = '{32'hc2c51eac, 32'h42b4b75e, 32'hc1b0fbbf, 32'h421fd8ff, 32'hc29a82fd, 32'hc267b7b1, 32'hc2088300, 32'hc222596e};
test_weights[10664:10671] = '{32'hc28700ae, 32'hc24dedb1, 32'hc2775339, 32'h4279c81d, 32'hc21336e6, 32'h41881372, 32'h41653bb5, 32'hc240c83a};
test_bias[1333:1333] = '{32'hc2ae2c73};
test_output[1333:1333] = '{32'h460e39d2};
test_input[10672:10679] = '{32'hc1b85d0a, 32'h42ac5cd5, 32'h426272c8, 32'h413d32c3, 32'h41b67e80, 32'h4288d14a, 32'hc2632907, 32'hc280b8ac};
test_weights[10672:10679] = '{32'hc219cd5b, 32'hc13a7474, 32'h41934f93, 32'hc18ecaf8, 32'h42b174e7, 32'h41cb8775, 32'hc15e6346, 32'h42b51903};
test_bias[1334:1334] = '{32'hc28b99e2};
test_output[1334:1334] = '{32'hc41da779};
test_input[10680:10687] = '{32'h40da85c1, 32'h42901a41, 32'hc22d24e7, 32'h42a4e376, 32'h42bd8f01, 32'h42880b45, 32'h41c34644, 32'h40c5d97b};
test_weights[10680:10687] = '{32'h41d482fd, 32'hc28781c9, 32'hc2831905, 32'h42b54e56, 32'h428dec1e, 32'hc2831cce, 32'h4196f9b6, 32'hc1e40a5d};
test_bias[1335:1335] = '{32'h4288ac80};
test_output[1335:1335] = '{32'h460097e5};
test_input[10688:10695] = '{32'hc2365598, 32'h41f9206f, 32'h4234d519, 32'hc272fe6a, 32'h41eeaa47, 32'h41886ca7, 32'hc2736740, 32'hc2add056};
test_weights[10688:10695] = '{32'h42bcb0d7, 32'hc138d5cc, 32'h42117369, 32'h42bf37f3, 32'h42c28957, 32'h428a8c17, 32'h429ce1de, 32'h42b7a122};
test_bias[1336:1336] = '{32'h42569112};
test_output[1336:1336] = '{32'hc68840a8};
test_input[10696:10703] = '{32'hc269fbf3, 32'hc2a67d6f, 32'hc2283375, 32'h41c0e904, 32'hc2a99d01, 32'h4295802f, 32'h4159441d, 32'h4083e892};
test_weights[10696:10703] = '{32'h4132dcb6, 32'hc289d72b, 32'h41de58a9, 32'hc2973865, 32'h425b5dbc, 32'h4205149f, 32'hc29287a8, 32'h42b4091f};
test_bias[1337:1337] = '{32'h429d02c1};
test_output[1337:1337] = '{32'hc41a790e};
test_input[10704:10711] = '{32'h42c481d5, 32'hc2c696d1, 32'hc26d901c, 32'hbfdcd5b2, 32'h419119a9, 32'hbfd51ade, 32'hc04af285, 32'h42aa0a1b};
test_weights[10704:10711] = '{32'h4277d247, 32'h4221b0ca, 32'hc0ae058b, 32'hc1ce2331, 32'h41a73439, 32'hc2820f0a, 32'h4255b070, 32'h41c8c26d};
test_bias[1338:1338] = '{32'h41e47a04};
test_output[1338:1338] = '{32'h4599c8b4};
test_input[10712:10719] = '{32'h41f0b472, 32'hc2499a94, 32'hc229ce76, 32'hc244f4c4, 32'h4184dccd, 32'hc108033d, 32'hc280bedb, 32'hc2abbc01};
test_weights[10712:10719] = '{32'h42659b35, 32'hc2803dc3, 32'hc2a25f4d, 32'hc25301e6, 32'hc0d966c2, 32'hc15b35d5, 32'hc1949a98, 32'hc11c61b0};
test_bias[1339:1339] = '{32'h41138fc2};
test_output[1339:1339] = '{32'h464bea95};
test_input[10720:10727] = '{32'h428c181a, 32'hc1b94321, 32'hc2685ee6, 32'hc19dcc37, 32'hc2b4989e, 32'h40eaeb15, 32'hbf2396a7, 32'hc26ce0fb};
test_weights[10720:10727] = '{32'hc2a00b49, 32'hc2c1daf4, 32'hc169ab27, 32'hc2804ce8, 32'h40ea7feb, 32'hc1e1d43f, 32'hc13b1ca9, 32'h42afbcc7};
test_bias[1340:1340] = '{32'hc29e29c9};
test_output[1340:1340] = '{32'hc5e6f865};
test_input[10728:10735] = '{32'h422c1973, 32'h427b96ba, 32'hc25b6a8c, 32'hc28924b3, 32'h421dcffa, 32'hbf9a91d3, 32'hc2600507, 32'hc2a7b342};
test_weights[10728:10735] = '{32'h41786529, 32'h42647e53, 32'hc1afcad9, 32'hc255f775, 32'h41154d0b, 32'hc2b1127f, 32'h42731d96, 32'hc2bb4af9};
test_bias[1341:1341] = '{32'h4214722b};
test_output[1341:1341] = '{32'h465c3afd};
test_input[10736:10743] = '{32'hc27ad863, 32'hc2524200, 32'h42c3105e, 32'hc2c33e73, 32'h42bc6180, 32'h428a40ea, 32'hc2483bac, 32'h426e5b86};
test_weights[10736:10743] = '{32'hc28424f3, 32'h41d02192, 32'h4136dbad, 32'hc239c67c, 32'h4030f7c8, 32'h422da787, 32'hc28d332f, 32'hc222b016};
test_bias[1342:1342] = '{32'hc2a61897};
test_output[1342:1342] = '{32'h4646a5e1};
test_input[10744:10751] = '{32'hc24c73c0, 32'h42341b8b, 32'h4280ec2e, 32'h42c436fa, 32'h42501f3f, 32'hc216a7b8, 32'hc20c44c8, 32'hc2077057};
test_weights[10744:10751] = '{32'hc142da95, 32'h4233d52d, 32'h42382879, 32'hc2122f2e, 32'h41b26dd7, 32'hc1b20758, 32'h4003a4fc, 32'h42931ec8};
test_bias[1343:1343] = '{32'h42c5cb25};
test_output[1343:1343] = '{32'h44c37965};
test_input[10752:10759] = '{32'hc12e0286, 32'hc2260915, 32'hc27433c5, 32'h42c642c3, 32'hc21dd7e0, 32'hc2702bb2, 32'h42a8f59f, 32'hc28111b9};
test_weights[10752:10759] = '{32'h4201b1ad, 32'hc25a9ddd, 32'h40dd6462, 32'hc28ae99d, 32'hc2c5595f, 32'h428cf33c, 32'hc2822042, 32'h4226a980};
test_bias[1344:1344] = '{32'h42156473};
test_output[1344:1344] = '{32'hc658d56f};
test_input[10760:10767] = '{32'h42bb114f, 32'hc146dc15, 32'h429fff4f, 32'h416ba41f, 32'h42a7c538, 32'hc28bc428, 32'hc2974555, 32'hc1e31cbc};
test_weights[10760:10767] = '{32'hbf87eb60, 32'h42196697, 32'hc0305bee, 32'h42aea5db, 32'hc26ddf61, 32'h426f261d, 32'h42c1f30b, 32'hc1f2f88e};
test_bias[1345:1345] = '{32'h4239f1de};
test_output[1345:1345] = '{32'hc66bfbe7};
test_input[10768:10775] = '{32'h429bf8cd, 32'h4182a871, 32'hc19538fd, 32'h42721de3, 32'hc1066b9b, 32'hc2793bc8, 32'hc2ae036f, 32'h4187f46e};
test_weights[10768:10775] = '{32'h4187923c, 32'hc2360ee8, 32'h3f734e8c, 32'h42af4871, 32'h4292ae29, 32'hc20528be, 32'h42740153, 32'hc2b5d795};
test_bias[1346:1346] = '{32'hc08b3a8d};
test_output[1346:1346] = '{32'h43e9372e};
test_input[10776:10783] = '{32'h42336b4e, 32'h42c4a202, 32'h42bb4097, 32'h427aa70d, 32'h42b6e4a5, 32'h41e59db2, 32'h4255f7c6, 32'h429b3bd7};
test_weights[10776:10783] = '{32'h4295a2a2, 32'h42c60935, 32'h42724fdd, 32'hc2399859, 32'h42bb8df7, 32'h41f0a28d, 32'hc22bdc9e, 32'hc2b783b5};
test_bias[1347:1347] = '{32'hc18f0880};
test_output[1347:1347] = '{32'h4677c046};
test_input[10784:10791] = '{32'hc2bd5903, 32'hc2339b15, 32'hc2a3b73b, 32'hc189e4fa, 32'h42148279, 32'hc2714442, 32'hc2330e54, 32'h4209fbcb};
test_weights[10784:10791] = '{32'hbfe01c94, 32'hc2c03532, 32'h426b86b8, 32'h42adb987, 32'h425c22da, 32'hc11ca9f7, 32'h4286a3e7, 32'hc0b477f0};
test_bias[1348:1348] = '{32'h42a46a32};
test_output[1348:1348] = '{32'hc51182cd};
test_input[10792:10799] = '{32'h429dafd0, 32'h42247cab, 32'hc2acfd87, 32'h41800f65, 32'hc2477efa, 32'hc298c798, 32'hc2b0d8a5, 32'hc256a329};
test_weights[10792:10799] = '{32'h4287ea73, 32'h4196eaec, 32'hc122e286, 32'hc22a2dfa, 32'hc29011df, 32'hc1c3322d, 32'hc1b1b515, 32'h42991a72};
test_bias[1349:1349] = '{32'hc1785698};
test_output[1349:1349] = '{32'h46167b1f};
test_input[10800:10807] = '{32'h42b97374, 32'hc2c38094, 32'hc2b6b6cc, 32'h41ecdd9e, 32'h42545eeb, 32'hbea9459d, 32'h42bf41a9, 32'hc2172e64};
test_weights[10800:10807] = '{32'hc2b763ec, 32'h42889a6d, 32'h4165ad71, 32'hc297c94b, 32'h41fd67b9, 32'hc292cd51, 32'h4299de6c, 32'h42b0294a};
test_bias[1350:1350] = '{32'hc1fa4fb2};
test_output[1350:1350] = '{32'hc64baae3};
test_input[10808:10815] = '{32'h42389873, 32'h426980b6, 32'hc2b2d784, 32'hc22e7588, 32'hc1bee65e, 32'h41ae0a38, 32'hc2628233, 32'hc20db9ca};
test_weights[10808:10815] = '{32'hc2294149, 32'h424498e6, 32'h404cfcdf, 32'hc2941454, 32'hc2c54775, 32'hc1e924a1, 32'h42a372a3, 32'hc0bad024};
test_bias[1351:1351] = '{32'h42b528c3};
test_output[1351:1351] = '{32'h449c13f9};
test_input[10816:10823] = '{32'hc21824bf, 32'h42a9fb2d, 32'hc075ae8e, 32'hc2a4709e, 32'hc2a09217, 32'h42aee342, 32'h41b0895a, 32'h41d32642};
test_weights[10816:10823] = '{32'h42722ee6, 32'h41cfffd4, 32'hc286bb4e, 32'hc283ea21, 32'hc2c496dc, 32'h4264b576, 32'h422c13c5, 32'hc0b55103};
test_bias[1352:1352] = '{32'hc2a59dd5};
test_output[1352:1352] = '{32'h4695f99e};
test_input[10824:10831] = '{32'h423d14cb, 32'h4284f66e, 32'h42b2d6fe, 32'hc26fb5df, 32'hc27b04f7, 32'h42bda9e6, 32'h42209aae, 32'h4285047a};
test_weights[10824:10831] = '{32'hc207b40d, 32'hc2c36292, 32'h41f32053, 32'hc285b3f5, 32'hc2242890, 32'h421cbe72, 32'h41f6ba19, 32'hc1cb2698};
test_bias[1353:1353] = '{32'h4207ab1d};
test_output[1353:1353] = '{32'h458ca186};
test_input[10832:10839] = '{32'hc2564746, 32'hc297f8f0, 32'hc2b099d4, 32'h42ab9ec9, 32'hc121fb03, 32'h419084a1, 32'hc1e23fe4, 32'hc20bc83f};
test_weights[10832:10839] = '{32'h424f7233, 32'h41807691, 32'h42c56893, 32'hc237deed, 32'h419377d9, 32'h42b21f6e, 32'hc22ff795, 32'hc2c3df10};
test_bias[1354:1354] = '{32'hc231f730};
test_output[1354:1354] = '{32'hc625d8bb};
test_input[10840:10847] = '{32'hc21dcd3b, 32'h423cb3b1, 32'hc2630a82, 32'hc21d25c6, 32'hc1c27fae, 32'hc240bf1f, 32'hc291e8b9, 32'h429fa5a4};
test_weights[10840:10847] = '{32'hc09b818a, 32'hc29dc774, 32'h42a62fef, 32'h42708848, 32'hc1e67829, 32'hc27305ae, 32'hc1f50626, 32'h425d4170};
test_bias[1355:1355] = '{32'hc1be97eb};
test_output[1355:1355] = '{32'hc3b16776};
test_input[10848:10855] = '{32'h40962827, 32'hc28e39fa, 32'h429474c8, 32'h422b3ac8, 32'h41dbafd1, 32'hc2abd7c5, 32'h42bd356d, 32'h4294be0e};
test_weights[10848:10855] = '{32'hc2036d45, 32'hc2a27d31, 32'h41483b85, 32'hc206a7a0, 32'hc2272454, 32'h41ce9a6d, 32'h423f66e3, 32'h41388ae6};
test_bias[1356:1356] = '{32'hc1950476};
test_output[1356:1356] = '{32'h45de36ea};
test_input[10856:10863] = '{32'hc20f8390, 32'hc2c754b2, 32'hc0ae66ea, 32'hc1c47ee7, 32'hc2ae49f9, 32'hc2570fa7, 32'h4212ae4f, 32'h42b3b651};
test_weights[10856:10863] = '{32'hc1900546, 32'h429ffff3, 32'h4239ac03, 32'hc212deec, 32'hc252f22f, 32'h3f80fa08, 32'hc293772b, 32'h413bfe6f};
test_bias[1357:1357] = '{32'h428f73db};
test_output[1357:1357] = '{32'hc5681379};
test_input[10864:10871] = '{32'hc157cad1, 32'hc1685c50, 32'hc226faec, 32'h41fb15c2, 32'hbedaac22, 32'h423bf29a, 32'h4107af27, 32'hc20361c2};
test_weights[10864:10871] = '{32'h4294c66e, 32'hc11941cf, 32'hc28f8f21, 32'h4172d458, 32'hc244a742, 32'hc1f3c11f, 32'h40ce71e0, 32'hc27a8da0};
test_bias[1358:1358] = '{32'hc165fce5};
test_output[1358:1358] = '{32'h454dfac3};
test_input[10872:10879] = '{32'h427d82c5, 32'hc20b33a3, 32'hc2b0ca3a, 32'hc2bfacc3, 32'hc272954d, 32'h424defd7, 32'h429b1a1f, 32'h423a9094};
test_weights[10872:10879] = '{32'h423f870f, 32'hc11a5707, 32'h4297bcf8, 32'h42129a70, 32'h42530b3e, 32'hc291613b, 32'hc29d29df, 32'hc0dcc326};
test_bias[1359:1359] = '{32'h42a020e6};
test_output[1359:1359] = '{32'hc69d3d16};
test_input[10880:10887] = '{32'hc20a7a6c, 32'hc0dd355c, 32'h41aec5f7, 32'h42c02704, 32'hc0b46bb8, 32'hc29ed733, 32'h3fd10e07, 32'hc245ccce};
test_weights[10880:10887] = '{32'h4229669b, 32'h428d257a, 32'h428a6b7b, 32'h41b1c84b, 32'h422771b9, 32'h42b62969, 32'h42933506, 32'h41920352};
test_bias[1360:1360] = '{32'h42673854};
test_output[1360:1360] = '{32'hc5cb2908};
test_input[10888:10895] = '{32'hc164655e, 32'hc215c011, 32'h42b3ea42, 32'hc2b58bf7, 32'h42527de2, 32'hc1989b46, 32'hc2900b84, 32'hc2c6621a};
test_weights[10888:10895] = '{32'h42ade417, 32'h426791b4, 32'hc292d368, 32'hc2af96c3, 32'hc2700a25, 32'h42c02b01, 32'hc28368cd, 32'hc24677c7};
test_bias[1361:1361] = '{32'hc2bbb605};
test_output[1361:1361] = '{32'h451de0d8};
test_input[10896:10903] = '{32'h42be17d5, 32'hc1ba4f45, 32'h420bfb70, 32'hc2915781, 32'hc2a8872e, 32'hc21da7ed, 32'hc26e5eab, 32'h3e41f479};
test_weights[10896:10903] = '{32'h41c9a133, 32'hc1f61262, 32'hc2b669b7, 32'hc2b45e9e, 32'h41d43715, 32'h41f98f37, 32'hc280b45a, 32'h421fb615};
test_bias[1362:1362] = '{32'hc2905b35};
test_output[1362:1362] = '{32'h45d3daee};
test_input[10904:10911] = '{32'h4296cfb3, 32'h4122e40f, 32'hc2a30a58, 32'hc2268ea0, 32'hc268b7ce, 32'hc20c19a5, 32'h42758b92, 32'h42b31021};
test_weights[10904:10911] = '{32'hc241b433, 32'h429545e9, 32'hc232f385, 32'hc12e2d5f, 32'hc2b82382, 32'h427e49ac, 32'h429607dc, 32'h41d5b2f7};
test_bias[1363:1363] = '{32'hc209f2c6};
test_output[1363:1363] = '{32'h46309231};
test_input[10912:10919] = '{32'hc2ab7d89, 32'h4261f2f7, 32'h4215ea8f, 32'hc2b92aaf, 32'hc2807f34, 32'h424149ef, 32'hc07c876f, 32'hc2357b58};
test_weights[10912:10919] = '{32'hc2600381, 32'h41d89f62, 32'h42c27881, 32'hc2959b02, 32'h418e3fbe, 32'hc2234bfc, 32'h4275a575, 32'hc2a30ace};
test_bias[1364:1364] = '{32'hc27cd85b};
test_output[1364:1364] = '{32'h468636b5};
test_input[10920:10927] = '{32'hc18b7eb4, 32'hc17269d6, 32'hc2055923, 32'h41df0f4b, 32'hc2bafe5e, 32'hc10105c7, 32'hc21f6dde, 32'hc192aac6};
test_weights[10920:10927] = '{32'hc1cc0052, 32'h4233be88, 32'h417b0871, 32'hc1c13568, 32'h42b98e9c, 32'hc2b6c55f, 32'h410df251, 32'hc23eb56d};
test_bias[1365:1365] = '{32'hc2362cde};
test_output[1365:1365] = '{32'hc60afcfa};
test_input[10928:10935] = '{32'h41273ab7, 32'hc2c2f11f, 32'h42857301, 32'hc27f9ce1, 32'h429e2143, 32'h42bfda1b, 32'hc2a8dbb5, 32'h428e34ff};
test_weights[10928:10935] = '{32'hc18cd7f0, 32'hc28fdf04, 32'hc2c6d1d6, 32'hc082c84b, 32'hc1945aae, 32'hc217e1fd, 32'h426e7ba3, 32'hc2be286c};
test_bias[1366:1366] = '{32'h429cf185};
test_output[1366:1366] = '{32'hc67fc24e};
test_input[10936:10943] = '{32'hc1a4feb9, 32'hc1981ab8, 32'hc27ea8a1, 32'hc1896086, 32'hc28c3940, 32'h42a7bb59, 32'hc25b1895, 32'hc29fe853};
test_weights[10936:10943] = '{32'h422b577b, 32'hc2a761a0, 32'hc2aecab1, 32'h42abd56a, 32'h429d6737, 32'h42051e39, 32'h411c8e83, 32'h42786a38};
test_bias[1367:1367] = '{32'h417048d7};
test_output[1367:1367] = '{32'hc5558d70};
test_input[10944:10951] = '{32'h41ccbf57, 32'hc2a338d7, 32'hc216a020, 32'h42c00d92, 32'hc024241e, 32'h4288450f, 32'hc200a283, 32'hc186ad50};
test_weights[10944:10951] = '{32'hc21b4789, 32'h42077615, 32'h40a5f20f, 32'h427ef35d, 32'hc2bacaf4, 32'h42aa9b98, 32'h42329ce0, 32'h429cce0c};
test_bias[1368:1368] = '{32'h41384485};
test_output[1368:1368] = '{32'h45ab1a22};
test_input[10952:10959] = '{32'hc2ad4213, 32'hc27430e7, 32'h420c0680, 32'hc29f160a, 32'h42bb5cbc, 32'h4243bc3c, 32'h41a972cc, 32'hc23ab63b};
test_weights[10952:10959] = '{32'h425b2e94, 32'h42281b82, 32'h42a40740, 32'hc25759c5, 32'hc2015eca, 32'hc24f53e2, 32'h41b2a0a2, 32'h42a79c4c};
test_bias[1369:1369] = '{32'hc2683773};
test_output[1369:1369] = '{32'hc610192d};
test_input[10960:10967] = '{32'h4286d746, 32'hc2801795, 32'h429c07b7, 32'h424981ce, 32'h42286918, 32'h3ff82d1d, 32'hc2a79780, 32'h41c63452};
test_weights[10960:10967] = '{32'h4219bddf, 32'h4209bd7b, 32'hc2981bee, 32'h42b672c5, 32'hc2b01e43, 32'h4243f937, 32'hc295f049, 32'h41a57efd};
test_bias[1370:1370] = '{32'hc1578f1c};
test_output[1370:1370] = '{32'h450a8bbe};
test_input[10968:10975] = '{32'h42b3c9a1, 32'hc2acbc91, 32'h427c07c2, 32'hc2837c60, 32'h42b10da2, 32'hbfbe5e12, 32'h4132ac35, 32'hc24a15eb};
test_weights[10968:10975] = '{32'hc0dafa5b, 32'h42397605, 32'h425a96ac, 32'h41c5c903, 32'h4222ef73, 32'hc2826bf9, 32'hc202f75a, 32'hc1b68949};
test_bias[1371:1371] = '{32'h421baff0};
test_output[1371:1371] = '{32'h44d7e777};
test_input[10976:10983] = '{32'hc1ecc888, 32'h429a6df5, 32'hc1a1def3, 32'hc2a78b14, 32'h42c4b363, 32'h4287234f, 32'h42455e83, 32'h41e2a973};
test_weights[10976:10983] = '{32'hc0a039d5, 32'hc2839287, 32'h424a5061, 32'hc189b841, 32'hc2c5bf5d, 32'hc2c16cf9, 32'h42b7df8b, 32'h423c04de};
test_bias[1372:1372] = '{32'hc241812d};
test_output[1372:1372] = '{32'hc669a023};
test_input[10984:10991] = '{32'h41c8dba5, 32'hc209ce11, 32'h420125d3, 32'h4228e0f6, 32'h409c34ab, 32'h41916d10, 32'hc12ca349, 32'h4030c59b};
test_weights[10984:10991] = '{32'h42196dab, 32'hc125db59, 32'h40be87e1, 32'h42519afd, 32'hc260f10e, 32'h42948682, 32'hc0c4d349, 32'h41a40266};
test_bias[1373:1373] = '{32'hc2402348};
test_output[1373:1373] = '{32'h4598597f};
test_input[10992:10999] = '{32'hc23c8f2e, 32'hc29a484b, 32'hc132649b, 32'hc2b27b3b, 32'hc2989398, 32'h41c0ef34, 32'h42492f7f, 32'h41ff329b};
test_weights[10992:10999] = '{32'h42455fe8, 32'hc1e76f1c, 32'h427594fe, 32'h428a0071, 32'hbf820251, 32'h42b7f6e1, 32'hc2766e79, 32'h42a6f59c};
test_bias[1374:1374] = '{32'h427bc598};
test_output[1374:1374] = '{32'hc59cac7f};
test_input[11000:11007] = '{32'hc2468b68, 32'h427a585e, 32'h423e30e6, 32'hc25ccf54, 32'hc229312d, 32'h4254c96c, 32'hc21bb188, 32'h42b44a81};
test_weights[11000:11007] = '{32'hc2ae0ac1, 32'h428513f9, 32'hc2b50ac2, 32'h42a169cf, 32'hc277fcfc, 32'h4235d27b, 32'h400b3ad5, 32'hc295ab60};
test_bias[1375:1375] = '{32'hc29e3f57};
test_output[1375:1375] = '{32'hc5060d67};
test_input[11008:11015] = '{32'hc2b0151e, 32'hc2a9562e, 32'h42aa7110, 32'hc2a03ccd, 32'h421e81f5, 32'hc21588c2, 32'h42aab65d, 32'hc1d7eda0};
test_weights[11008:11015] = '{32'hc23b3303, 32'hc219e3aa, 32'hc1aa422b, 32'hc198ee4b, 32'hc2a8c31a, 32'hc21a551e, 32'h42c58614, 32'h42592d7d};
test_bias[1376:1376] = '{32'h428c78f1};
test_output[1376:1376] = '{32'h463f13a2};
test_input[11016:11023] = '{32'h4279ddf2, 32'hc2b32ab8, 32'hc20bfe86, 32'hc2523c3b, 32'h42c2a87d, 32'hc0a9c9c8, 32'h42ae4e97, 32'hc264398b};
test_weights[11016:11023] = '{32'h42349504, 32'h4295b250, 32'hc191bdcf, 32'h42b6fe72, 32'h4225cd2c, 32'hc1e4bd1c, 32'hc29ff464, 32'hc2bdabbc};
test_bias[1377:1377] = '{32'h42c6b226};
test_output[1377:1377] = '{32'hc5a69366};
test_input[11024:11031] = '{32'hc2a01374, 32'h421407db, 32'hc2a139e2, 32'hc20c8a2d, 32'h409edc6e, 32'h424cf84f, 32'hc1bef042, 32'hc1fb3fbc};
test_weights[11024:11031] = '{32'h4292aec2, 32'hc2197b3a, 32'hc1b8c23b, 32'hc1f058cb, 32'h41592a71, 32'hc1499e8b, 32'h423d66aa, 32'hc2a8139a};
test_bias[1378:1378] = '{32'hc02efd7a};
test_output[1378:1378] = '{32'hc5574a66};
test_input[11032:11039] = '{32'h429c2432, 32'hc262018d, 32'hc2b31c4b, 32'hc1c375f2, 32'h42a99ddf, 32'hc2994735, 32'hc2c06794, 32'h41b66f1f};
test_weights[11032:11039] = '{32'h41964112, 32'h422e558e, 32'h420ac7f4, 32'hc2999ad7, 32'hc212208b, 32'h42b37275, 32'h4288a8e9, 32'h41566e33};
test_bias[1379:1379] = '{32'hc27025a8};
test_output[1379:1379] = '{32'hc690c2aa};
test_input[11040:11047] = '{32'hc200ad51, 32'hc2b594ae, 32'h42a2a99d, 32'hc0edfa6d, 32'h42616b8a, 32'h412b00fa, 32'h41f74831, 32'h4189626c};
test_weights[11040:11047] = '{32'h429195bd, 32'h40c3ef73, 32'hc273c635, 32'hc0e2699f, 32'hc28f6383, 32'hc1d1a501, 32'hc2b22140, 32'h410c04cd};
test_bias[1380:1380] = '{32'hc2a994d9};
test_output[1380:1380] = '{32'hc667661c};
test_input[11048:11055] = '{32'hc1aa8dfb, 32'hc20e12fe, 32'hc2ad2089, 32'hc2b8a5dd, 32'h421e5631, 32'hc1a96e49, 32'hc2b3b8ca, 32'h42bf0224};
test_weights[11048:11055] = '{32'h41d27ed4, 32'hc1d40079, 32'h42bdda97, 32'h428e2161, 32'h42595b33, 32'hc29975c4, 32'hc2115024, 32'hc1b4c32d};
test_bias[1381:1381] = '{32'h41efb208};
test_output[1381:1381] = '{32'hc61435a1};
test_input[11056:11063] = '{32'h4291b641, 32'h42c0ed46, 32'hc233df63, 32'h42adfbfc, 32'h4175ccdc, 32'h42409e84, 32'h41bff845, 32'h42ba1d8b};
test_weights[11056:11063] = '{32'h41bc1e43, 32'hc17fd370, 32'hc25914ad, 32'h422fc255, 32'hc23f67da, 32'hc2123041, 32'hc208a059, 32'hc2934794};
test_bias[1382:1382] = '{32'hc1273128};
test_output[1382:1382] = '{32'hc56a031b};
test_input[11064:11071] = '{32'h42c7886c, 32'h3d690200, 32'hc2c0047e, 32'hc1abb555, 32'h424a4582, 32'hc1e2ba06, 32'hc2960608, 32'hc20a5c3a};
test_weights[11064:11071] = '{32'hc27c4ea6, 32'h42c5dfe9, 32'h4205b8bb, 32'hc080ca9b, 32'hc283e151, 32'h4122fb73, 32'hc26b4bff, 32'hc26f1f91};
test_bias[1383:1383] = '{32'h427f9f38};
test_output[1383:1383] = '{32'hc5cacb9b};
test_input[11072:11079] = '{32'h42228033, 32'h4255cfc7, 32'h428f5aaf, 32'h41afe8a7, 32'hc2646563, 32'hc2acaaf8, 32'hc2603fdb, 32'h4251e2ee};
test_weights[11072:11079] = '{32'hc129f280, 32'hc2b22c3d, 32'h42224929, 32'h423ab298, 32'h412924e1, 32'hc2a5c8dd, 32'hbffd380e, 32'h41b79a11};
test_bias[1384:1384] = '{32'hc23a4af4};
test_output[1384:1384] = '{32'h45cd123a};
test_input[11080:11087] = '{32'hc10ece2d, 32'hc10205ce, 32'hc2948e9d, 32'h42bdee81, 32'h42c374f5, 32'h42a3a802, 32'hc2a7609b, 32'hc2075d69};
test_weights[11080:11087] = '{32'hc2a20e28, 32'hc23564e9, 32'h4257b90e, 32'h42911884, 32'hc2a07133, 32'h41d5a301, 32'hc248f924, 32'hc0ad7d19};
test_bias[1385:1385] = '{32'h40d8a9fc};
test_output[1385:1385] = '{32'h4529bbcf};
test_input[11088:11095] = '{32'h429f6107, 32'hc1a18dee, 32'h4221a669, 32'hc2bbdd35, 32'h4194bb4c, 32'hc2c0a09a, 32'hc12739b7, 32'h41c06a7b};
test_weights[11088:11095] = '{32'h42c0cc6f, 32'h422893d3, 32'h40e9b884, 32'h41b3f3fa, 32'h4199770f, 32'h429e0738, 32'h41b4f37e, 32'h4281a7b7};
test_bias[1386:1386] = '{32'h40b9dac2};
test_output[1386:1386] = '{32'hc463eb87};
test_input[11096:11103] = '{32'hc113dbbb, 32'h42bf05f1, 32'hc24a2e36, 32'h4280192d, 32'h427ae16e, 32'hc0dd4843, 32'hc1c11b05, 32'hc2bd05eb};
test_weights[11096:11103] = '{32'h42876309, 32'h424a81e0, 32'hc2256390, 32'h42935be1, 32'h4250607f, 32'h42748471, 32'hc24fb77b, 32'hc2beb626};
test_bias[1387:1387] = '{32'h423274ce};
test_output[1387:1387] = '{32'h46bcdbb3};
test_input[11104:11111] = '{32'hc203abb4, 32'h41bfd549, 32'h3f1096f4, 32'hc146a79f, 32'hc20831ee, 32'h411ef02f, 32'hc22e83b2, 32'hc24629bd};
test_weights[11104:11111] = '{32'hc11b5afe, 32'h42c6ac6e, 32'h4111e4d4, 32'hc2a29063, 32'hc1646f79, 32'h41cb8ca5, 32'hc2ac493c, 32'h4182ad9e};
test_bias[1388:1388] = '{32'h4186bf8a};
test_output[1388:1388] = '{32'h45e7e601};
test_input[11112:11119] = '{32'h42c5d104, 32'h421c1d17, 32'hc08914d9, 32'h40926214, 32'h428b6adc, 32'h4222cdb9, 32'h41994baf, 32'hc0dafcfa};
test_weights[11112:11119] = '{32'hc2bbf212, 32'hc117e556, 32'hbe9087be, 32'h41d67a3a, 32'hc294eaf5, 32'h42abae39, 32'h429d7d0f, 32'h4214d291};
test_bias[1389:1389] = '{32'hc2875813};
test_output[1389:1389] = '{32'hc61d0d97};
test_input[11120:11127] = '{32'hc2a453e6, 32'hc28cea51, 32'h42872f4c, 32'h40a830f7, 32'hc219848f, 32'h42b6e02f, 32'hc1ef62d5, 32'h42a9ec32};
test_weights[11120:11127] = '{32'hc29e731d, 32'h41041f43, 32'h42104d1d, 32'hc2a86ca1, 32'hc0c357c3, 32'hc1a9920a, 32'hc290deb9, 32'hc29b88b5};
test_bias[1390:1390] = '{32'hc2b10e9a};
test_output[1390:1390] = '{32'h44d36a3d};
test_input[11128:11135] = '{32'hc22ca766, 32'hc120c637, 32'h428c4759, 32'h42a619ed, 32'hc1ede1cd, 32'h40c03d16, 32'h42147599, 32'h41864941};
test_weights[11128:11135] = '{32'h42aa78e2, 32'h40c658d5, 32'h41d15dd7, 32'hc14fb199, 32'hc206be11, 32'hc250f8e2, 32'h42941be4, 32'hc250c82b};
test_bias[1391:1391] = '{32'h4258a4ac};
test_output[1391:1391] = '{32'hc3b8bee8};
test_input[11136:11143] = '{32'h42105a07, 32'hc0120608, 32'h423bec1c, 32'h416f6cdc, 32'hc2b4753f, 32'hc287ef86, 32'hc299007d, 32'hc28587a4};
test_weights[11136:11143] = '{32'hc1e8ec5a, 32'hc0b1984e, 32'hc21adb7b, 32'h41bc5271, 32'hc29295a2, 32'hc2bba6fc, 32'hbed76f83, 32'hc2436273};
test_bias[1392:1392] = '{32'h41aa6c03};
test_output[1392:1392] = '{32'h4657a153};
test_input[11144:11151] = '{32'hc1886b6d, 32'hc22bbdea, 32'hc20eae7c, 32'hc248c650, 32'hc21d1b73, 32'hc2a7f09d, 32'hc0d2de6d, 32'h41a665d1};
test_weights[11144:11151] = '{32'hc20d8ea9, 32'h428b44b3, 32'h42bcd6ee, 32'hc28f2fd4, 32'hc1e4a672, 32'h42b42cc9, 32'h42835521, 32'hc23eb01a};
test_bias[1393:1393] = '{32'hc296d348};
test_output[1393:1393] = '{32'hc61dda09};
test_input[11152:11159] = '{32'h42a88c44, 32'h409fb79c, 32'h428466c6, 32'hc1abe9ee, 32'hc28e6294, 32'hc01a53b5, 32'h408cbc8f, 32'hc2459fdb};
test_weights[11152:11159] = '{32'hc15c941d, 32'h42c316dd, 32'hc291aa98, 32'hc2b65ae8, 32'h4243b7e3, 32'h41b1e6ff, 32'hc2beacc1, 32'hc28e3340};
test_bias[1394:1394] = '{32'hc281f9ec};
test_output[1394:1394] = '{32'hc57cdc6d};
test_input[11160:11167] = '{32'h4240e18f, 32'h40eca213, 32'h42928805, 32'hc100fc06, 32'hc20a8522, 32'h41cc7ecc, 32'hc2743368, 32'h40438470};
test_weights[11160:11167] = '{32'hc1469033, 32'hc2a550f1, 32'hc2289f8a, 32'hc27f645e, 32'hc1891404, 32'h41a46624, 32'hc21ff2d6, 32'h3fa407eb};
test_bias[1395:1395] = '{32'hc290f313};
test_output[1395:1395] = '{32'hc39217f5};
test_input[11168:11175] = '{32'hc25cede8, 32'hc2951137, 32'h428054fe, 32'hc156e70b, 32'h428d24c3, 32'hc14ea9e8, 32'hc2c760b7, 32'h4243ac63};
test_weights[11168:11175] = '{32'h42232bae, 32'h42a414f9, 32'h41b69c91, 32'hc17553f4, 32'hc1ae8c4a, 32'hc2975a3b, 32'hc043f353, 32'h4242e840};
test_bias[1396:1396] = '{32'hc2a019bd};
test_output[1396:1396] = '{32'hc5915607};
test_input[11176:11183] = '{32'hc276c110, 32'h41d324d1, 32'h41eab3ac, 32'hc11c567a, 32'hc1296c59, 32'h41eb28f9, 32'hc28f2a14, 32'hc23502b1};
test_weights[11176:11183] = '{32'hc2805ada, 32'hc20dee99, 32'h423a2cff, 32'h42a22925, 32'hc124f489, 32'hc1e58059, 32'hc0afb5e6, 32'h41810458};
test_bias[1397:1397] = '{32'h4082ff9b};
test_output[1397:1397] = '{32'h451e101d};
test_input[11184:11191] = '{32'h42ae80da, 32'h420cb82a, 32'hc2961b8f, 32'h427db12c, 32'hc20a450a, 32'h42b60e20, 32'hc05b1b68, 32'hc29fcec2};
test_weights[11184:11191] = '{32'hc28ff2bb, 32'hc2c77630, 32'h4223b374, 32'hc2b8de2d, 32'hc14c47cd, 32'h425f4aba, 32'hc2321f24, 32'h41a35adf};
test_bias[1398:1398] = '{32'hc2b13149};
test_output[1398:1398] = '{32'hc666bd7a};
test_input[11192:11199] = '{32'hc180b1e8, 32'hc1661ba7, 32'hc17681af, 32'h4261ac3c, 32'h4295aa94, 32'hc19d5618, 32'h4293ba3d, 32'hc235711c};
test_weights[11192:11199] = '{32'hc28d221f, 32'h42810a19, 32'hc29b12a7, 32'hc2a9231e, 32'hc1885f1b, 32'hc182fe85, 32'h425a331c, 32'hc2a4cb08};
test_bias[1399:1399] = '{32'hc2bebae0};
test_output[1399:1399] = '{32'h455147ed};
test_input[11200:11207] = '{32'hc24fc36c, 32'hc25f7744, 32'hc1aaea11, 32'h429742e6, 32'h4168aa56, 32'h419ee4c5, 32'h425bb0b2, 32'h427c2a87};
test_weights[11200:11207] = '{32'h428e90c7, 32'hc2be62e6, 32'hc207ee1a, 32'hc199b3d2, 32'hc2a5517b, 32'hbf908e43, 32'h42573f3f, 32'h41a1d365};
test_bias[1400:1400] = '{32'h42b918c4};
test_output[1400:1400] = '{32'h457935fe};
test_input[11208:11215] = '{32'hc291e2f3, 32'hc22d80f1, 32'hc259dee4, 32'h42bd09e5, 32'h418e5042, 32'h3f90dee1, 32'hc11f9655, 32'h4164aa19};
test_weights[11208:11215] = '{32'h410d08a9, 32'h40a1267d, 32'hc24421d4, 32'h424764b4, 32'h42a951ee, 32'hc2023b12, 32'hc29bdf52, 32'h416b7ffc};
test_bias[1401:1401] = '{32'h423257d2};
test_output[1401:1401] = '{32'h460cf9aa};
test_input[11216:11223] = '{32'hc2971afe, 32'hc124beb3, 32'h40330052, 32'hc281f10e, 32'hc29c401b, 32'h42bc7a7e, 32'h42a83b88, 32'h4286bec3};
test_weights[11216:11223] = '{32'hc2b8be63, 32'h42af2ff4, 32'hc266c9e0, 32'hc278e996, 32'h42ae7ed4, 32'h422205ca, 32'h425952a9, 32'hc1d65ea2};
test_bias[1402:1402] = '{32'hc2a00010};
test_output[1402:1402] = '{32'h4616b1a8};
test_input[11224:11231] = '{32'hc2a47e25, 32'hc173586e, 32'hc285701e, 32'h4184c82b, 32'h42a91dd4, 32'h427fe441, 32'h415faa7c, 32'h427ddb4c};
test_weights[11224:11231] = '{32'h4285402d, 32'h41a74112, 32'h4278d9c0, 32'hc1bb0a8b, 32'h429aa22f, 32'h42b2342b, 32'hc23d7e8e, 32'h4284ef86};
test_bias[1403:1403] = '{32'hc29462f4};
test_output[1403:1403] = '{32'h45a83a3e};
test_input[11232:11239] = '{32'h4250ff7b, 32'hc0cc6b10, 32'h4138133b, 32'h42c1189b, 32'hc29bedeb, 32'h425aca5e, 32'h41cf3022, 32'hc1aa71d1};
test_weights[11232:11239] = '{32'hc25c9b22, 32'h421a9e35, 32'hc2c17a04, 32'hc162a903, 32'h42b14ab7, 32'h407e7845, 32'hc29747c2, 32'h4234fe37};
test_bias[1404:1404] = '{32'h42a2bc19};
test_output[1404:1404] = '{32'hc66ca293};
test_input[11240:11247] = '{32'hc1dc40b8, 32'hc22c1362, 32'h42170ef5, 32'hc103127f, 32'hc219f105, 32'hc2577c1e, 32'h41b9bbc8, 32'hc2597608};
test_weights[11240:11247] = '{32'hc2c5104c, 32'hc2b1882d, 32'hc24b6279, 32'h41e0c2d1, 32'h42b27830, 32'h428215e8, 32'hc2b0c616, 32'h428dfb4e};
test_bias[1405:1405] = '{32'h42a0588b};
test_output[1405:1405] = '{32'hc60311db};
test_input[11248:11255] = '{32'hc29512e5, 32'h42a3c5f7, 32'hc1b5e0ef, 32'hc287bd10, 32'hc201aedd, 32'hc283b4bc, 32'h42098c9b, 32'hc2ad5f2a};
test_weights[11248:11255] = '{32'hc1071f75, 32'hc17a4405, 32'hc1b97f9d, 32'h4204aa0d, 32'hc226d415, 32'hc28fa516, 32'h419b01e8, 32'h42753534};
test_bias[1406:1406] = '{32'h422044ae};
test_output[1406:1406] = '{32'hc4613ad7};
test_input[11256:11263] = '{32'hc1e3f496, 32'h424185c6, 32'h42940e9a, 32'h40ba7f7d, 32'h42801180, 32'hc2bd42c3, 32'hc29b574d, 32'hc2a12021};
test_weights[11256:11263] = '{32'h42851112, 32'h420d84dc, 32'h423faa71, 32'hc197704e, 32'hc2c53b0a, 32'h4195981e, 32'h42a99209, 32'hc2b891e2};
test_bias[1407:1407] = '{32'hc1a386c0};
test_output[1407:1407] = '{32'hc57a2922};
test_input[11264:11271] = '{32'hc2712e4e, 32'h422a0335, 32'hc213b0de, 32'h426526bd, 32'h42adb307, 32'h429b80fd, 32'h42b59a0f, 32'hc0cf5d82};
test_weights[11264:11271] = '{32'h425028ba, 32'h41f04455, 32'hc27b1539, 32'hc13f0ef7, 32'h4287c2c3, 32'h4197cf62, 32'hc26b55f5, 32'h420a19e4};
test_bias[1408:1408] = '{32'hc18d1395};
test_output[1408:1408] = '{32'h44c2f463};
test_input[11272:11279] = '{32'hc1bf0505, 32'hc1bf9e81, 32'hc25ac125, 32'hc21cf4e5, 32'h42853b74, 32'hc2696a91, 32'h42a3c0b7, 32'hc2329f0c};
test_weights[11272:11279] = '{32'hc0a85747, 32'h41d35125, 32'h428222a6, 32'h4114a0b9, 32'hc2824e5c, 32'hc28fc36e, 32'hc27ad3f4, 32'h3ef05b23};
test_bias[1409:1409] = '{32'hc197751c};
test_output[1409:1409] = '{32'hc6185743};
test_input[11280:11287] = '{32'hc201dc10, 32'hc1ef0cd0, 32'hc2ab0fa4, 32'hc169d9a0, 32'hc295b88b, 32'hc192b82b, 32'h4214a10a, 32'hc167de03};
test_weights[11280:11287] = '{32'hc1527d3b, 32'hc29bd1d5, 32'hc24e9166, 32'hc2c75542, 32'h42ada665, 32'hc205edf0, 32'h425557af, 32'h4121a6ee};
test_bias[1410:1410] = '{32'hc264617f};
test_output[1410:1410] = '{32'h458d4b33};
test_input[11288:11295] = '{32'h428d4fad, 32'h42836d45, 32'hc2a16405, 32'h42c21ac8, 32'hc108b85e, 32'hc24cf0b0, 32'h426d6a99, 32'hc2866d66};
test_weights[11288:11295] = '{32'hc20bbfc5, 32'h414e2d58, 32'h415ff4c7, 32'h4260b33b, 32'hc28c8eeb, 32'h42b69737, 32'h42ba670a, 32'hc218f5d0};
test_bias[1411:1411] = '{32'h424aceb1};
test_output[1411:1411] = '{32'h45d3c42e};
test_input[11296:11303] = '{32'h42bbf458, 32'h41ac6267, 32'h42af60b1, 32'h418dcaa0, 32'h428fcb01, 32'h42c35774, 32'hc22fb8cc, 32'h41d4e6e9};
test_weights[11296:11303] = '{32'h41993935, 32'hc14db4a2, 32'hc2b0855d, 32'h42b8e471, 32'hc10b2917, 32'hc19b3487, 32'hc292a245, 32'h42b57f8e};
test_bias[1412:1412] = '{32'hc2a428d3};
test_output[1412:1412] = '{32'hc4c10c90};
test_input[11304:11311] = '{32'h42b02886, 32'h4287dc68, 32'hc2135e8d, 32'hc1b598e2, 32'hc240a4fb, 32'hc2508b10, 32'hc2a2fc16, 32'hc27c6b8f};
test_weights[11304:11311] = '{32'hc153dd29, 32'hc285b085, 32'hc226a727, 32'h42b273b8, 32'h422b3ff5, 32'h3ee32253, 32'h427887af, 32'h428cafbe};
test_bias[1413:1413] = '{32'hc209ff46};
test_output[1413:1413] = '{32'hc68b36c5};
test_input[11312:11319] = '{32'h4298dc49, 32'hc2c317e7, 32'h4291dd6f, 32'h427e52a0, 32'h42622294, 32'hc2740e3a, 32'hc117acd1, 32'hc29fd623};
test_weights[11312:11319] = '{32'h410e809a, 32'h424d7990, 32'hc12763ad, 32'h4121415d, 32'h42ab70f5, 32'h40e98f86, 32'h42956dd2, 32'h416818e3};
test_bias[1414:1414] = '{32'hc1c2d169};
test_output[1414:1414] = '{32'hc4f2ef67};
test_input[11320:11327] = '{32'h41c7b74d, 32'hc223cf5a, 32'h426e4a74, 32'h42ba919a, 32'hc128bda1, 32'hc201e8a3, 32'h42423831, 32'h428cbcb2};
test_weights[11320:11327] = '{32'hc28adc2e, 32'hc18b2c16, 32'hc286f0b2, 32'h42689fca, 32'h42b18a7c, 32'h429dc1f8, 32'hc267f719, 32'h42a5ce84};
test_bias[1415:1415] = '{32'h420fa98c};
test_output[1415:1415] = '{32'hc26cce44};
test_input[11328:11335] = '{32'h4247c22d, 32'h425b73cd, 32'h42c5169d, 32'h4019f5c9, 32'h425e990f, 32'h42985d57, 32'hc2354aa2, 32'h41a9242d};
test_weights[11328:11335] = '{32'h421bee5f, 32'h4210adc2, 32'hc2bf1236, 32'hc0ad2d1c, 32'hc2b26085, 32'hc1f55ea6, 32'hc1ce17e6, 32'hc28468c8};
test_bias[1416:1416] = '{32'h42a966fb};
test_output[1416:1416] = '{32'hc64a3eaf};
test_input[11336:11343] = '{32'h42728190, 32'hc2a572ea, 32'hc28b91bf, 32'hc12e04ed, 32'h4247d273, 32'h41c505eb, 32'hc170201b, 32'h4249e916};
test_weights[11336:11343] = '{32'h422ae017, 32'h4062820b, 32'hc293d38d, 32'hc2bb7451, 32'hc2882900, 32'hc0b13abc, 32'hc1441228, 32'h42c0e9ee};
test_bias[1417:1417] = '{32'hc1a6c548};
test_output[1417:1417] = '{32'h461bc480};
test_input[11344:11351] = '{32'h423db3a1, 32'h41740bc4, 32'hc2aad028, 32'hc28b7548, 32'h40098d35, 32'h41f9a29e, 32'hc2ae46b1, 32'hc1cdf79d};
test_weights[11344:11351] = '{32'h42880ef3, 32'h424ab670, 32'hc0f80dc7, 32'hc2b270e0, 32'hc2473d4a, 32'hc18fa5c3, 32'hc2b43df4, 32'hc2897da8};
test_bias[1418:1418] = '{32'h41787a9a};
test_output[1418:1418] = '{32'h469b1b52};
test_input[11352:11359] = '{32'hc1ea0308, 32'h4209d0e3, 32'hc211f6f5, 32'h42200ecb, 32'h4233d537, 32'hc2aaaf62, 32'h423a1293, 32'h427d8b36};
test_weights[11352:11359] = '{32'h424e6730, 32'h41ce9c32, 32'h4293e7c3, 32'hc20b9649, 32'h41d9f620, 32'hc2821f67, 32'h4073fd1d, 32'hc1de1356};
test_bias[1419:1419] = '{32'hc2bc543a};
test_output[1419:1419] = '{32'h43c13835};
test_input[11360:11367] = '{32'h419156f0, 32'h3e6ad5ef, 32'h4283da32, 32'h420b4273, 32'hc24e26e5, 32'h42b3453b, 32'h4296a469, 32'h42423e5c};
test_weights[11360:11367] = '{32'h4296fd7c, 32'h428d5518, 32'h42c5823b, 32'hc1d3e3ba, 32'h41e094f5, 32'hc1887b1e, 32'h4281b5ac, 32'hc18e8fef};
test_bias[1420:1420] = '{32'hc2b771cc};
test_output[1420:1420] = '{32'h45f7bfe9};
test_input[11368:11375] = '{32'h42ac52c9, 32'h4139ca62, 32'hc1f2118c, 32'hc2a67a35, 32'hc200d73b, 32'hc28cbe9e, 32'h42046f5a, 32'hc292ce70};
test_weights[11368:11375] = '{32'h4239624f, 32'h425a20a7, 32'h4260eb1e, 32'h42b1e38b, 32'h40bc6c0a, 32'h4115aa93, 32'hc28c6c00, 32'h42a8aba5};
test_bias[1421:1421] = '{32'hc1e92086};
test_output[1421:1421] = '{32'hc658bae2};
test_input[11376:11383] = '{32'hc20f1436, 32'hc255129b, 32'h41a073b1, 32'h4222db2f, 32'hc24ad816, 32'hc1c4561a, 32'hc017e25e, 32'hc2aa9fb3};
test_weights[11376:11383] = '{32'h42a0e915, 32'h4285dfc6, 32'hc2b1f3c3, 32'h408973c1, 32'hc282f3ce, 32'h41c3d5b4, 32'h42a96b7f, 32'h42bfe8ec};
test_bias[1422:1422] = '{32'hc0b91089};
test_output[1422:1422] = '{32'hc65679de};
test_input[11384:11391] = '{32'hc251023c, 32'h42c56b28, 32'h424a5cad, 32'hc263073c, 32'h41ac2e28, 32'h425c638a, 32'hc2b9e82e, 32'h4247e0a4};
test_weights[11384:11391] = '{32'h42abff48, 32'hc248a62c, 32'h42ae2a1d, 32'h429b5732, 32'h4191a572, 32'h428a90f2, 32'hc22b0858, 32'h42b85cde};
test_bias[1423:1423] = '{32'h41cb700e};
test_output[1423:1423] = '{32'h455276ed};
test_input[11392:11399] = '{32'h42a0b470, 32'h42adb7fa, 32'h425b2f70, 32'h40e059d8, 32'hc2a0821d, 32'hc216e619, 32'h423a4a87, 32'h4244e42a};
test_weights[11392:11399] = '{32'h42036f54, 32'hc12036e6, 32'hc16d63fa, 32'h424314fd, 32'h419b45a8, 32'h426bd0c1, 32'hc10569af, 32'h42534d6c};
test_bias[1424:1424] = '{32'h418f2a09};
test_output[1424:1424] = '{32'hc37c7278};
test_input[11400:11407] = '{32'h42b80ed8, 32'h42c1e390, 32'hc18e922c, 32'h42b31943, 32'hc2c42d29, 32'hc292122f, 32'hc15f7097, 32'h4293159d};
test_weights[11400:11407] = '{32'hc0de0795, 32'hc27aee36, 32'hc20add86, 32'hc12bd477, 32'h3ee4f6af, 32'h4216f053, 32'h4284bb1c, 32'hc1bf7017};
test_bias[1425:1425] = '{32'hc26f71e7};
test_output[1425:1425] = '{32'hc64505dc};
test_input[11408:11415] = '{32'h4095f890, 32'hc1e6d8aa, 32'h42269282, 32'hc2b39fcb, 32'h418fb094, 32'hc2517b67, 32'h4276736d, 32'h429768ec};
test_weights[11408:11415] = '{32'hc25f26ce, 32'hc2a97555, 32'h42412d85, 32'hc2461206, 32'hc14ed2be, 32'hbf8f0b83, 32'hc2184a67, 32'hc0ff7e91};
test_bias[1426:1426] = '{32'hc1a53e9a};
test_output[1426:1426] = '{32'h45abcafd};
test_input[11416:11423] = '{32'h40c842e6, 32'hc1ada12e, 32'hc2a89f26, 32'h400d4e27, 32'h428033f6, 32'hc0ae570d, 32'h428ac889, 32'hc1d538d9};
test_weights[11416:11423] = '{32'hc28d1b96, 32'h42c662d4, 32'h42a21ce2, 32'h42166f0a, 32'hc296e067, 32'hc29bf4ab, 32'hc23073de, 32'h417449fd};
test_bias[1427:1427] = '{32'hc1767fd1};
test_output[1427:1427] = '{32'hc686af30};
test_input[11424:11431] = '{32'h40eff581, 32'hc220f219, 32'hc1ca579f, 32'h4272baf5, 32'h41a256ab, 32'h42c1e05b, 32'hc2aade6e, 32'hc27f4858};
test_weights[11424:11431] = '{32'h423e4636, 32'h428cdea6, 32'hc23bb88c, 32'h40771f44, 32'h420a2d37, 32'hc13a08d1, 32'hc2b93c77, 32'hc223b9a3};
test_bias[1428:1428] = '{32'hc2a1284f};
test_output[1428:1428] = '{32'h460c0927};
test_input[11432:11439] = '{32'hc0251c47, 32'hc2be21f2, 32'h42c71231, 32'h42257c18, 32'h422419b9, 32'h40491be8, 32'h414e72c5, 32'hc146fd5f};
test_weights[11432:11439] = '{32'h429bf4e2, 32'h42ac534b, 32'h427b84df, 32'hc2881b5b, 32'h4292c33a, 32'hc25ad42d, 32'hc274411d, 32'h40288b6f};
test_bias[1429:1429] = '{32'hc2163689};
test_output[1429:1429] = '{32'hc5398a99};
test_input[11440:11447] = '{32'h42c45667, 32'h428f5411, 32'hc18910a9, 32'h429a9b9a, 32'hc193fac6, 32'h412b4509, 32'h4274be34, 32'hc2a4292e};
test_weights[11440:11447] = '{32'hc2b588f1, 32'hc2af8032, 32'hc251dc68, 32'h3ed3ab57, 32'h40ba08ca, 32'hc1cb0975, 32'h42c0dc47, 32'hc21159a0};
test_bias[1430:1430] = '{32'hc130dd3a};
test_output[1430:1430] = '{32'hc5b47df4};
test_input[11448:11455] = '{32'hc21fb6ff, 32'hbf97db82, 32'hc2b0950d, 32'hc0d9e09b, 32'hc20cc3ab, 32'h41ce22bd, 32'h429c9b6a, 32'h4218810c};
test_weights[11448:11455] = '{32'h4281c87a, 32'h41ac86e8, 32'h42824018, 32'h40b082f4, 32'h42b91025, 32'h41ed25cb, 32'h4286dcab, 32'hc2212f42};
test_bias[1431:1431] = '{32'hc24cd2a6};
test_output[1431:1431] = '{32'hc5e1208b};
test_input[11456:11463] = '{32'hc1b36cf8, 32'hc21af22c, 32'h4239cf82, 32'h422590c9, 32'h42bc506f, 32'h420a014c, 32'h41da396d, 32'hc2492d18};
test_weights[11456:11463] = '{32'hc2306b3a, 32'hc1b3c7d4, 32'hc222303c, 32'hc15f3c42, 32'h429a8801, 32'h41d4b65d, 32'h4279c139, 32'hc1deb269};
test_bias[1432:1432] = '{32'h422a53b8};
test_output[1432:1432] = '{32'h4627c3df};
test_input[11464:11471] = '{32'hc0ba98d5, 32'h42b26085, 32'h3fa162af, 32'h422db880, 32'h42bac04a, 32'h42a08c58, 32'h42c44fd4, 32'h425ae92b};
test_weights[11464:11471] = '{32'h42a73902, 32'hc20215ca, 32'hc22977fc, 32'hc279ee28, 32'hc298e0af, 32'h40045cb3, 32'hc28a5a31, 32'h424758c0};
test_bias[1433:1433] = '{32'hc277ef52};
test_output[1433:1433] = '{32'hc686c66b};
test_input[11472:11479] = '{32'hc2abe7e1, 32'hc21578d6, 32'hc1fd174e, 32'h41876582, 32'h41c88bf3, 32'hc2a150fd, 32'h427a909b, 32'h4110c6fb};
test_weights[11472:11479] = '{32'hc0bb9b9d, 32'hc2ab7e7e, 32'h4288bb18, 32'hc0abd380, 32'hc1ee87c9, 32'h42759f4a, 32'h42766ffa, 32'hc1b35dfa};
test_bias[1434:1434] = '{32'hc24211cc};
test_output[1434:1434] = '{32'hc41f80b5};
test_input[11480:11487] = '{32'hc2876500, 32'hc2b714a8, 32'hc2028e20, 32'hc23527af, 32'h42a2bf86, 32'h42a0c0a3, 32'h42bfea2a, 32'h41d65c4c};
test_weights[11480:11487] = '{32'hc2127ffc, 32'hc161d120, 32'h42b3c02f, 32'hc26f63dd, 32'h414c31b6, 32'h403ee7ea, 32'hc2c494cc, 32'hc10c6d7c};
test_bias[1435:1435] = '{32'h422471fc};
test_output[1435:1435] = '{32'hc595f91f};
test_input[11488:11495] = '{32'hc2b6eb29, 32'hc29ffe1e, 32'h422edf35, 32'h42bf7202, 32'h41ff5e48, 32'hc2b10a16, 32'h4298e3c4, 32'hc2aa673c};
test_weights[11488:11495] = '{32'hc2192351, 32'h4214e751, 32'hc27e905f, 32'h42817584, 32'hc15fb1a4, 32'h4174d8c5, 32'h42c1cdfa, 32'h4290f183};
test_bias[1436:1436] = '{32'h42373072};
test_output[1436:1436] = '{32'h455573e6};
test_input[11496:11503] = '{32'hc1ecec44, 32'h42408f24, 32'h42a5abc2, 32'h4244439c, 32'hc19426ad, 32'h4197ae27, 32'h42aca98b, 32'h4182137f};
test_weights[11496:11503] = '{32'h428dc8da, 32'hc21fd565, 32'h42082da6, 32'hc2b2d75e, 32'h40f06f70, 32'hc1f73304, 32'h4272ce80, 32'h40c5e536};
test_bias[1437:1437] = '{32'h422baf59};
test_output[1437:1437] = '{32'hc468e626};
test_input[11504:11511] = '{32'hc288bbc3, 32'hc2c2deff, 32'h425e7184, 32'h3f885fa9, 32'h4281ae9c, 32'h41dab525, 32'h4014eea9, 32'hc217453b};
test_weights[11504:11511] = '{32'hc0e6727c, 32'hc199e89d, 32'hc228d59c, 32'h40d05e47, 32'hc2c672d7, 32'h4271cf6f, 32'hc0af27ae, 32'hc2a08c28};
test_bias[1438:1438] = '{32'h427bb8b8};
test_output[1438:1438] = '{32'hc4d09420};
test_input[11512:11519] = '{32'hc111bb37, 32'h4291e913, 32'h4254387e, 32'h4220f708, 32'hc22ea84f, 32'hc0d21083, 32'h41204a56, 32'hc15568ba};
test_weights[11512:11519] = '{32'h4268a2b6, 32'h420f0c0f, 32'hc29ace70, 32'hbfc95b93, 32'h429e8bb0, 32'h42496937, 32'h415074ce, 32'hc11f6476};
test_bias[1439:1439] = '{32'h3f690a1c};
test_output[1439:1439] = '{32'hc5af9254};
test_input[11520:11527] = '{32'h42b78a60, 32'h4240d286, 32'h4218c58b, 32'h42bce001, 32'h42a29b3e, 32'h42b8c343, 32'hc2afd784, 32'h4243b305};
test_weights[11520:11527] = '{32'h424122f8, 32'h42b5c11f, 32'hc1d99ada, 32'h427b5eb4, 32'hc17cb5be, 32'h41d8f2df, 32'hc2bb2669, 32'hc1eb3ba1};
test_bias[1440:1440] = '{32'hc248138f};
test_output[1440:1440] = '{32'h46a946bc};
test_input[11528:11535] = '{32'h425714ff, 32'h3fe0c839, 32'hc1a45324, 32'hc2c6a9be, 32'hc0cfe25c, 32'h42b16465, 32'hc277cd1e, 32'h428b9d26};
test_weights[11528:11535] = '{32'h424bb84f, 32'hc1bcd3af, 32'hc2926296, 32'h42bf5c2d, 32'hc29794d5, 32'hc2759022, 32'h42b2ef5f, 32'h42b30ad4};
test_bias[1441:1441] = '{32'h42783723};
test_output[1441:1441] = '{32'hc6143e5a};
test_input[11536:11543] = '{32'h3ef15e35, 32'hc1e7b8b7, 32'h4246147f, 32'hc2ba5aaf, 32'hc1efd470, 32'hc2467cc2, 32'h42906e4d, 32'hc2bb3ae7};
test_weights[11536:11543] = '{32'h4174bdc0, 32'hc040af17, 32'h42053a7a, 32'h429690a8, 32'h428b5699, 32'h429206e7, 32'hc288e304, 32'hc2bdee0e};
test_bias[1442:1442] = '{32'hc2a40be8};
test_output[1442:1442] = '{32'hc5de6833};
test_input[11544:11551] = '{32'h4235a0ae, 32'h42a452a8, 32'hc2769462, 32'h41a63273, 32'hc28aaa1b, 32'h428ba307, 32'hc2b15194, 32'hc2b0ecf6};
test_weights[11544:11551] = '{32'h423061bd, 32'hc218bb0f, 32'hc23d9477, 32'h412edff5, 32'h40d4a0be, 32'h4290445b, 32'h42bdce49, 32'hbfce519b};
test_bias[1443:1443] = '{32'hc1e78a88};
test_output[1443:1443] = '{32'hc4d5e031};
test_input[11552:11559] = '{32'h42bff6c0, 32'h4214201a, 32'hc1caf1cc, 32'hc2a59205, 32'h42279ff5, 32'hc20fb594, 32'hc2c7802e, 32'hc203fa38};
test_weights[11552:11559] = '{32'h4148e64b, 32'hc2be27df, 32'h412805ad, 32'hc1cc3cb7, 32'h418d93cf, 32'hc13f70e7, 32'h42bec2b1, 32'h409b0ea4};
test_bias[1444:1444] = '{32'hc2b844bc};
test_output[1444:1444] = '{32'hc60d9d60};
test_input[11560:11567] = '{32'h4272bd8f, 32'h4214c147, 32'h402157fa, 32'hc0c0fa6f, 32'h422b1eef, 32'h42965f5b, 32'h410a61bd, 32'h42475b8f};
test_weights[11560:11567] = '{32'hc2962e28, 32'h42c0198c, 32'h42313601, 32'hc0e98f92, 32'hc255a336, 32'h4079d6c1, 32'hc119e9ba, 32'h421fb12f};
test_bias[1445:1445] = '{32'h427e3b99};
test_output[1445:1445] = '{32'hc4549bc2};
test_input[11568:11575] = '{32'hc27e0226, 32'hc27a1fe5, 32'hc1120e01, 32'h425578b0, 32'h4281bc00, 32'h420247a2, 32'hc0804b7f, 32'h405969a3};
test_weights[11568:11575] = '{32'h42b8a1fe, 32'hc2bb7900, 32'hc296c1c7, 32'h42b160fd, 32'h42155c13, 32'hc2a0699c, 32'h41e501ee, 32'h40daacb9};
test_bias[1446:1446] = '{32'hc2aa1b43};
test_output[1446:1446] = '{32'h459decf8};
test_input[11576:11583] = '{32'hc194dd16, 32'h41f8a050, 32'h41c35922, 32'hc191ee2c, 32'h410da80b, 32'h42a7f09b, 32'h424871c6, 32'h4280996b};
test_weights[11576:11583] = '{32'h42a50826, 32'hc10a726d, 32'hbf6886e5, 32'h42c51920, 32'h426b6271, 32'hc1d402ce, 32'hc2b9ef5c, 32'h42a00188};
test_bias[1447:1447] = '{32'h4295dbe8};
test_output[1447:1447] = '{32'hc595012a};
test_input[11584:11591] = '{32'h42b564b3, 32'h429c6e7a, 32'hc02953fb, 32'hc21c674b, 32'hc297f7f9, 32'h424cdedb, 32'hc297bb9e, 32'hc18a0842};
test_weights[11584:11591] = '{32'h427c6de3, 32'hc252b0b9, 32'hc1be3156, 32'h42b7294b, 32'h428c33bd, 32'h42abecec, 32'hc223e0e8, 32'h402bf674};
test_bias[1448:1448] = '{32'hc231d4a2};
test_output[1448:1448] = '{32'h4333717c};
test_input[11592:11599] = '{32'hc29abd7f, 32'h42a264ef, 32'h412f05c8, 32'hc157a683, 32'h42493f90, 32'h428d8ac1, 32'h412b57ff, 32'hc2b08852};
test_weights[11592:11599] = '{32'h42542a89, 32'hc20776ed, 32'hc1f1b2af, 32'h41151cda, 32'h426c1156, 32'hc244f28c, 32'hc1c8941c, 32'h42bea46c};
test_bias[1449:1449] = '{32'h42c02ad1};
test_output[1449:1449] = '{32'hc6803631};
test_input[11600:11607] = '{32'hc2794f41, 32'h42816669, 32'h4231f256, 32'h3f040532, 32'h42b0ec20, 32'h42c3676b, 32'hc22b4c34, 32'h411c109f};
test_weights[11600:11607] = '{32'h428cdb4e, 32'hc135f49e, 32'hc22ae645, 32'hc2c6291c, 32'h41f5dd24, 32'h421eb5b5, 32'h41829ed6, 32'hc2967c92};
test_bias[1450:1450] = '{32'hc2b2d28f};
test_output[1450:1450] = '{32'hc4fa8fdf};
test_input[11608:11615] = '{32'hc2132174, 32'h4276bf67, 32'hc2a9ded8, 32'h42b0656d, 32'h42bb7fb8, 32'hc286809b, 32'hc27044de, 32'hc21c0118};
test_weights[11608:11615] = '{32'hc29e3ef7, 32'hc2a1e117, 32'hc295ec30, 32'h40209cae, 32'hc1bd26e4, 32'h42befc7f, 32'hc2aa997f, 32'h4138160f};
test_bias[1451:1451] = '{32'hc00a8b33};
test_output[1451:1451] = '{32'h4406f539};
test_input[11616:11623] = '{32'h424b0a8d, 32'hc26e0693, 32'hc2c2e1f6, 32'h41a108bc, 32'hc2b6c02d, 32'hc2c31227, 32'hc298a10f, 32'h42c1bb3b};
test_weights[11616:11623] = '{32'hc233dbc9, 32'h42a0e047, 32'hc1831e11, 32'h420e25df, 32'hc01cf48e, 32'hc2c73269, 32'hc118e4ef, 32'h41b613fc};
test_bias[1452:1452] = '{32'h423dd4cc};
test_output[1452:1452] = '{32'h45ff1986};
test_input[11624:11631] = '{32'hc24e55ed, 32'hc23bfc78, 32'h4266ab87, 32'hc2c0a5da, 32'hc29a7dd2, 32'h3f88d0aa, 32'h428b16dc, 32'hc2ab641b};
test_weights[11624:11631] = '{32'h4128374b, 32'hc290b12e, 32'hc234dd92, 32'h429c98b7, 32'hc263b86b, 32'h42142f54, 32'hc2b06e84, 32'h42ae344a};
test_bias[1453:1453] = '{32'h41f7894c};
test_output[1453:1453] = '{32'hc6804dc3};
test_input[11632:11639] = '{32'hc2b34f0e, 32'hc1e9fdcc, 32'h429c843c, 32'hc2797929, 32'hc12a67a3, 32'h429ab0cb, 32'hc2ae83b7, 32'h423d0ef3};
test_weights[11632:11639] = '{32'h4285dde4, 32'hc2492d21, 32'hc1a36bbf, 32'hc14f09c9, 32'h42176b28, 32'hc23ed5de, 32'hc012158f, 32'hc2b45244};
test_bias[1454:1454] = '{32'hc24ae235};
test_output[1454:1454] = '{32'hc6535e5f};
test_input[11640:11647] = '{32'hc228227b, 32'hc2b236f7, 32'hc29bae47, 32'hc1f8a2d2, 32'h40afac84, 32'hc1b72694, 32'hc28caf92, 32'hc2b998f9};
test_weights[11640:11647] = '{32'hc29b74b9, 32'hc2297fd8, 32'h4262564c, 32'hc28a1da7, 32'hc2255328, 32'h42833695, 32'hc21a7768, 32'h408400af};
test_bias[1455:1455] = '{32'h42b7b3a0};
test_output[1455:1455] = '{32'h45ab4b4c};
test_input[11648:11655] = '{32'h42664a48, 32'hc1d39250, 32'h427f8217, 32'hc2844927, 32'hc1e17c39, 32'hc21b3224, 32'hc248a5ec, 32'h42653d52};
test_weights[11648:11655] = '{32'h41825752, 32'h41fc283e, 32'hc28b2f00, 32'hc1fa68d1, 32'hc1e3e13f, 32'hc2bdb68e, 32'h42bc7faf, 32'h42a6921a};
test_bias[1456:1456] = '{32'h41da3ea8};
test_output[1456:1456] = '{32'h450ed46b};
test_input[11656:11663] = '{32'hc2147571, 32'hc2b036b2, 32'h4291304b, 32'hc2b12c80, 32'hc1e8ff0c, 32'hc29ecfaf, 32'hc285519b, 32'h42b7680e};
test_weights[11656:11663] = '{32'hc1f51a4e, 32'hc28ddc38, 32'hc023de48, 32'hc23cafa1, 32'h4273296d, 32'hc215e145, 32'h42984cef, 32'h42b0048f};
test_bias[1457:1457] = '{32'hc277c05d};
test_output[1457:1457] = '{32'h467273a9};
test_input[11664:11671] = '{32'h42416baf, 32'h42a1492b, 32'hc29ebaeb, 32'h42bbcff2, 32'hc2977ed6, 32'h428f04f8, 32'h4183dfe7, 32'h42825d7b};
test_weights[11664:11671] = '{32'hc23ef87f, 32'h426351b2, 32'hc2a13378, 32'h41b87889, 32'h40f11d69, 32'h42bb7872, 32'hc1f349dc, 32'h41c94cb1};
test_bias[1458:1458] = '{32'h4282fd9e};
test_output[1458:1458] = '{32'h468dfa3f};
test_input[11672:11679] = '{32'h42bc607b, 32'hc2508fc4, 32'h4230796d, 32'h41dd6867, 32'h427c9353, 32'hc2a51aa5, 32'h3fba4ffd, 32'h42b37fd8};
test_weights[11672:11679] = '{32'hc291111e, 32'h421bb8d1, 32'hc2164109, 32'h4259d9e9, 32'hc2a7629d, 32'hc241daf7, 32'hc23c06a6, 32'hc2009392};
test_bias[1459:1459] = '{32'h4213c827};
test_output[1459:1459] = '{32'hc64e6f8b};
test_input[11680:11687] = '{32'h4232da50, 32'hbf2f5539, 32'h42882115, 32'hc10537d9, 32'hc2616ad6, 32'h428d3c40, 32'h42aed766, 32'h42c08213};
test_weights[11680:11687] = '{32'h42b23d25, 32'h41df7a9f, 32'hc18d3d57, 32'hc268ec0d, 32'hc28c6ea2, 32'h40a9f8f0, 32'h42327966, 32'hc24c0235};
test_bias[1460:1460] = '{32'h42bc4257};
test_output[1460:1460] = '{32'h45d053ba};
test_input[11688:11695] = '{32'hc2a22606, 32'hc20c486f, 32'h42a2f636, 32'h3de6987d, 32'hc132b23e, 32'hc1f8743f, 32'h41e4e374, 32'h42ac1e7a};
test_weights[11688:11695] = '{32'h40a83705, 32'hc1d61f38, 32'hc2840e64, 32'hc1cac968, 32'hc216f72d, 32'h423dc577, 32'h418c7755, 32'hc10f432c};
test_bias[1461:1461] = '{32'h420e07fd};
test_output[1461:1461] = '{32'hc5c057f6};
test_input[11696:11703] = '{32'hc25f86cd, 32'h42b99dcf, 32'h429e49e5, 32'hc1dcacb2, 32'h428a1f41, 32'h413fe2b6, 32'h4102d064, 32'h42c20a5c};
test_weights[11696:11703] = '{32'h415122ab, 32'hc066b5d0, 32'h42c06adc, 32'hc291ddf0, 32'hc2a9a667, 32'h426a4922, 32'h428f5465, 32'hc0a65443};
test_bias[1462:1462] = '{32'h42b88db1};
test_output[1462:1462] = '{32'h455fb739};
test_input[11704:11711] = '{32'hc232fd28, 32'hc29b59f8, 32'h42c3a561, 32'h417656a5, 32'h3faf1b0a, 32'hc2b0c320, 32'hc2b6dc5a, 32'hc12cbb1b};
test_weights[11704:11711] = '{32'hc2c312df, 32'h418a275c, 32'hc287c69f, 32'hc1aa8d5e, 32'hc28e537a, 32'hc28f7cc2, 32'hc26b9060, 32'hc26bfcdd};
test_bias[1463:1463] = '{32'hc19b3ac1};
test_output[1463:1463] = '{32'h4601acf3};
test_input[11712:11719] = '{32'h41f651c4, 32'h42042c4a, 32'h414e03ed, 32'h422f65b9, 32'hc247b137, 32'h42853462, 32'hc1b75613, 32'hc2c5c70a};
test_weights[11712:11719] = '{32'hc2be00c0, 32'h4264cd87, 32'h428ad748, 32'hc1d77992, 32'hc29875d1, 32'hc289565f, 32'hc1b10ebb, 32'h4205b9ed};
test_bias[1464:1464] = '{32'h421a84c0};
test_output[1464:1464] = '{32'hc59791b8};
test_input[11720:11727] = '{32'h42ad4f03, 32'h4243f63d, 32'h41f1fda2, 32'h426fe633, 32'hc2a0f256, 32'h427a7dc9, 32'h42c69175, 32'hc2b0fd13};
test_weights[11720:11727] = '{32'hc26fcf17, 32'h42225631, 32'hc2409e00, 32'h42787b29, 32'h42b095cd, 32'h41f83210, 32'hc1b73d2a, 32'h428543db};
test_bias[1465:1465] = '{32'h4128fb14};
test_output[1465:1465] = '{32'hc65ed14e};
test_input[11728:11735] = '{32'hc29370a9, 32'h4258b20b, 32'hc2b955db, 32'h42b0f182, 32'h429f806a, 32'hc29222d0, 32'h4215189f, 32'hc2b47f55};
test_weights[11728:11735] = '{32'h42bf6a1f, 32'hc29e52a9, 32'h40f1fef9, 32'h4216d4a9, 32'hc28ec936, 32'hc2875776, 32'h42699ebe, 32'h42367b6d};
test_bias[1466:1466] = '{32'hc2610eb2};
test_output[1466:1466] = '{32'hc632f92e};
test_input[11736:11743] = '{32'hc24c22a2, 32'h415e93d9, 32'hc133e55f, 32'h42bd3bae, 32'hc2a13f1c, 32'h42aea9b9, 32'h416f9798, 32'hc23a64fb};
test_weights[11736:11743] = '{32'hc29c2f67, 32'hc27c6534, 32'h41c81ff5, 32'h40ef36fc, 32'hc275792e, 32'hc25a113b, 32'h42696578, 32'hc1306a18};
test_bias[1467:1467] = '{32'hc289a05e};
test_output[1467:1467] = '{32'h459d784a};
test_input[11744:11751] = '{32'hc1d3f088, 32'hc22ac5ba, 32'hc26c4ac3, 32'h427e4f27, 32'hc28ee035, 32'hc1a27e41, 32'h4200246a, 32'h414045ea};
test_weights[11744:11751] = '{32'hc1d6fdc1, 32'hc29b1d1b, 32'h42643a1f, 32'hc162ae05, 32'hc1f74c1c, 32'hc2a61659, 32'hc2c30df5, 32'h428d031a};
test_bias[1468:1468] = '{32'h417c2066};
test_output[1468:1468] = '{32'h44ad332b};
test_input[11752:11759] = '{32'h42920f66, 32'h42b47112, 32'h428da76c, 32'h424101e3, 32'h42ae683a, 32'h42854979, 32'h42b9e38d, 32'h42544c7e};
test_weights[11752:11759] = '{32'hc2a03753, 32'hc295fdfa, 32'hc20afb60, 32'hc203cbab, 32'hc2c40621, 32'hc290a29f, 32'h428af9ed, 32'hc24e8c25};
test_bias[1469:1469] = '{32'h41764721};
test_output[1469:1469] = '{32'hc6cd78e2};
test_input[11760:11767] = '{32'h4141f1ca, 32'h41eb0ccd, 32'h428f20d5, 32'hc26ce6df, 32'h428c6c47, 32'hc2bcf2f9, 32'h4253a7ab, 32'h429ce787};
test_weights[11760:11767] = '{32'hc118926e, 32'hc22ce663, 32'hc2ab24ed, 32'h42432b5a, 32'hc28233e8, 32'h420f92b4, 32'h425bc545, 32'h42a78a9d};
test_bias[1470:1470] = '{32'hc234ae77};
test_output[1470:1470] = '{32'hc60b7c34};
test_input[11768:11775] = '{32'h422b10bc, 32'hc20d997b, 32'h41ae7b89, 32'hc2bb3d8e, 32'hc21258cd, 32'h4295540d, 32'h42755ba3, 32'hc2b65c80};
test_weights[11768:11775] = '{32'h42336306, 32'h41f5cb14, 32'hc1fbcdea, 32'hc1fe6338, 32'h42749659, 32'hc1836ecb, 32'hc292d9bd, 32'h4165400e};
test_bias[1471:1471] = '{32'h4114a537};
test_output[1471:1471] = '{32'hc5c00090};
test_input[11776:11783] = '{32'h4211a807, 32'h41047666, 32'hc2b271aa, 32'hc1ae4cd0, 32'h4286c56e, 32'h3fe42a8f, 32'h3f765326, 32'hc2b219ca};
test_weights[11776:11783] = '{32'hc1ee9eb3, 32'h41be2cf3, 32'h412e496f, 32'h4226b3ee, 32'hc23f7629, 32'hc2b1122f, 32'h425f4e77, 32'hc003e2e4};
test_bias[1472:1472] = '{32'hc1823480};
test_output[1472:1472] = '{32'hc5b95c55};
test_input[11784:11791] = '{32'h42a524a2, 32'h42021d1e, 32'h41d0599b, 32'h404fc3ab, 32'h4050edbe, 32'h42474771, 32'hc2b58ba7, 32'hc28cfc86};
test_weights[11784:11791] = '{32'hc12ef393, 32'h42b796bf, 32'hc2979669, 32'h42325080, 32'h4249ab7e, 32'hc29134fa, 32'hc172d376, 32'h42258649};
test_bias[1473:1473] = '{32'h428ab8a1};
test_output[1473:1473] = '{32'hc591e64f};
test_input[11792:11799] = '{32'h42c0c310, 32'hc211d39d, 32'hc1f62754, 32'h42892379, 32'h42c5dd91, 32'hc29e767c, 32'h4259bae8, 32'hc23cc787};
test_weights[11792:11799] = '{32'h42b9dcf0, 32'h42ab9938, 32'hc1bfef5c, 32'hc2b726d5, 32'hc28101ec, 32'h42957363, 32'h42a5a8c6, 32'hc255b5d1};
test_bias[1474:1474] = '{32'hc2c7d9e4};
test_output[1474:1474] = '{32'hc59ee101};
test_input[11800:11807] = '{32'hc285b61a, 32'h4202010e, 32'hc28d084d, 32'hc07c8136, 32'hc2972da9, 32'hc234bb88, 32'hc2adf98b, 32'h41ffed0e};
test_weights[11800:11807] = '{32'hc2be6f43, 32'hc20a8b96, 32'h4293130c, 32'hc1fbe94f, 32'hc289009a, 32'hc1c22008, 32'h41c264af, 32'h428758b6};
test_bias[1475:1475] = '{32'h4149a031};
test_output[1475:1475] = '{32'h45cba756};
test_input[11808:11815] = '{32'hc27d3660, 32'hc1587939, 32'hc272d5f2, 32'h42a57abd, 32'hc2a90fd1, 32'h421cbbab, 32'h42b2cd26, 32'h4293fb68};
test_weights[11808:11815] = '{32'hc1b7915d, 32'hc0ac7a0e, 32'hbf9c2da9, 32'h42a1abd6, 32'h41e9626b, 32'h42589aeb, 32'h42b52d85, 32'h407b38ba};
test_bias[1476:1476] = '{32'hc2840785};
test_output[1476:1476] = '{32'h467e2b32};
test_input[11816:11823] = '{32'h4268f04f, 32'h421db29c, 32'h422b6342, 32'h420255e1, 32'hc22b7af6, 32'hc28f7d90, 32'hc2921c5a, 32'hc28a116c};
test_weights[11816:11823] = '{32'h42102799, 32'h404c3c71, 32'hc28cba03, 32'hc228ccd8, 32'h428bfbd1, 32'hc291c78c, 32'hc1aee439, 32'h42c7a131};
test_bias[1477:1477] = '{32'h41fa3118};
test_output[1477:1477] = '{32'hc5a27590};
test_input[11824:11831] = '{32'hc2627ee8, 32'h425a9f51, 32'h424412f7, 32'hc0955003, 32'hc1aa2461, 32'h429ea8b3, 32'h429876ff, 32'hc2c57d49};
test_weights[11824:11831] = '{32'hc2173bc7, 32'h4204c21f, 32'h4281f60e, 32'hc0559f86, 32'h427fe7fd, 32'hc23a5a33, 32'h429d124a, 32'h429a493f};
test_bias[1478:1478] = '{32'hc24a9117};
test_output[1478:1478] = '{32'h43d10bb5};
test_input[11832:11839] = '{32'hc1e7be3a, 32'h41b11775, 32'hc2b5fcc0, 32'h428b4e54, 32'hc2856065, 32'h41f8c9a9, 32'h3fa7b09d, 32'h4235cdf6};
test_weights[11832:11839] = '{32'h42afad8d, 32'hc1cd4953, 32'h429d2ccf, 32'h42181369, 32'h4146cba5, 32'hc2252f45, 32'hc29a3d50, 32'h42328101};
test_bias[1479:1479] = '{32'hc2bcb37e};
test_output[1479:1479] = '{32'hc5f6ba55};
test_input[11840:11847] = '{32'hc2958cce, 32'h4251a7b2, 32'h422e4e25, 32'hc2b5689b, 32'h425cf2df, 32'h4098308a, 32'hc00f8517, 32'hc2c339d5};
test_weights[11840:11847] = '{32'hc0b3813c, 32'hc22b6948, 32'hc22c8af7, 32'h4233a9dc, 32'h4258bb31, 32'hc2b3dc17, 32'hc0c4aeb0, 32'h41863c18};
test_bias[1480:1480] = '{32'hc293fae9};
test_output[1480:1480] = '{32'hc5d80a21};
test_input[11848:11855] = '{32'hc27c099f, 32'h41c36d21, 32'h42bd402b, 32'h42b8b8e0, 32'hc20a21b3, 32'h4289e04d, 32'h42b2bcc5, 32'hc252eda5};
test_weights[11848:11855] = '{32'hc25135ee, 32'h42a8440f, 32'hc198d10d, 32'hc2151894, 32'hc18d7a57, 32'h42c1620a, 32'h414adac5, 32'h420bed2a};
test_bias[1481:1481] = '{32'h428a3252};
test_output[1481:1481] = '{32'h45d2740a};
test_input[11856:11863] = '{32'hc27ff40f, 32'hc28a69fe, 32'h4285e7e8, 32'h42add810, 32'h42178a55, 32'h429e2d61, 32'h41eb9795, 32'hc183d497};
test_weights[11856:11863] = '{32'hc24f6fb1, 32'h426a4320, 32'h42c56585, 32'hc1eeeabf, 32'hc2986ea8, 32'h42303541, 32'hc2942ea3, 32'h414a17a3};
test_bias[1482:1482] = '{32'h429afe8e};
test_output[1482:1482] = '{32'h44c32f6a};
test_input[11864:11871] = '{32'hc28473b3, 32'h42aaa1c4, 32'hc23179ba, 32'h40f91f56, 32'hc257d3fb, 32'h41f1af9e, 32'h424d219c, 32'h42c618b9};
test_weights[11864:11871] = '{32'hc2b88559, 32'hc1212712, 32'hc287c907, 32'h426ca578, 32'hc22def18, 32'h4287986e, 32'h4292b903, 32'h42b855b6};
test_bias[1483:1483] = '{32'hc2bcf72c};
test_output[1483:1483] = '{32'h46ca759d};
test_input[11872:11879] = '{32'h42a6ecff, 32'hc1af4b61, 32'h41b7e426, 32'h42217d1a, 32'hc22661ab, 32'h42386cab, 32'hc21151a1, 32'h4245b015};
test_weights[11872:11879] = '{32'h42804c40, 32'hc1f7f780, 32'h429cb4ef, 32'h425c2331, 32'hc1b9d93a, 32'h4287fc83, 32'hc2250d61, 32'hc23ed02f};
test_bias[1484:1484] = '{32'h41af3898};
test_output[1484:1484] = '{32'h465022f9};
test_input[11880:11887] = '{32'hc2634fdc, 32'h429e3927, 32'hc2667625, 32'h42a57de2, 32'hc25641ee, 32'hc0aa4679, 32'h41ff575d, 32'h3ff9e9b7};
test_weights[11880:11887] = '{32'h428e6c9b, 32'hc27ea2f2, 32'hc1981141, 32'hc2a003d2, 32'hc2146d54, 32'h4160c20b, 32'h42961b70, 32'h42b0c03d};
test_bias[1485:1485] = '{32'hc2bcd291};
test_output[1485:1485] = '{32'hc61fb669};
test_input[11888:11895] = '{32'hc260955b, 32'hc1cbdcda, 32'hc0e86467, 32'h42993c1e, 32'h4261c37c, 32'h42b239f0, 32'h428ead99, 32'hc27f0428};
test_weights[11888:11895] = '{32'hc2c1d010, 32'hc27fc390, 32'hc2104207, 32'h4214d068, 32'h42b6342c, 32'h42c0faee, 32'hc2b51541, 32'h4252f40e};
test_bias[1486:1486] = '{32'h422d057c};
test_output[1486:1486] = '{32'h465d037f};
test_input[11896:11903] = '{32'h42b3396a, 32'h424512d2, 32'h41a762a4, 32'hc2305db0, 32'h41b6fbbb, 32'hc2a8952b, 32'h423a82a8, 32'h42c5f73a};
test_weights[11896:11903] = '{32'h41b43007, 32'h41e52e82, 32'hbff4f89f, 32'hc20dca71, 32'h3fe54ef8, 32'hbe86ee8b, 32'hc2167724, 32'hc29945ac};
test_bias[1487:1487] = '{32'h42068a11};
test_output[1487:1487] = '{32'hc58610c1};
test_input[11904:11911] = '{32'hc28643ec, 32'h42783d5d, 32'h4228a15a, 32'hc2b379fb, 32'h42500d1c, 32'h42953d96, 32'hbe757683, 32'hc25e849f};
test_weights[11904:11911] = '{32'h426091c7, 32'h42b0d08a, 32'h41c68217, 32'h41d1b15b, 32'hc0a0f432, 32'hc1c4a459, 32'hc1b4c8c5, 32'hc1041c65};
test_bias[1488:1488] = '{32'hc275b90c};
test_output[1488:1488] = '{32'hc4a020c9};
test_input[11912:11919] = '{32'h3fd32b0a, 32'hc2680f0c, 32'h429a079b, 32'hc2a7d843, 32'hc1a234c6, 32'hc10ce0bc, 32'h42be4f01, 32'hc2820c31};
test_weights[11912:11919] = '{32'hc1799b4c, 32'h4290975e, 32'hc20cb359, 32'h41bebb89, 32'h4247d945, 32'hc19cfacb, 32'hc2bcceeb, 32'h41a8a6a2};
test_bias[1489:1489] = '{32'h42371422};
test_output[1489:1489] = '{32'hc69cdc0d};
test_input[11920:11927] = '{32'h428881ad, 32'h4212ed01, 32'h404548cb, 32'hc23d7102, 32'hc1bcc25c, 32'h41afbd2a, 32'h4146292b, 32'h42ac949e};
test_weights[11920:11927] = '{32'hc20fe7e6, 32'hc276f8bd, 32'h4186b2b5, 32'hc2384c61, 32'h41ee380d, 32'hc29f8445, 32'hc294bc26, 32'hc1b5ed3d};
test_bias[1490:1490] = '{32'h41b6ecc5};
test_output[1490:1490] = '{32'hc5f3e498};
test_input[11928:11935] = '{32'h41ee4dfc, 32'hc2c22e3a, 32'hc224676e, 32'hc298dcbf, 32'h42a624e4, 32'h428c2aa3, 32'h40d91f2e, 32'h41d3797c};
test_weights[11928:11935] = '{32'hc2931ec3, 32'hc1d3a342, 32'h424a2e89, 32'hc29266da, 32'hc1eebf4a, 32'hc18ee482, 32'hc27ade59, 32'h414e5dfe};
test_bias[1491:1491] = '{32'h420231bd};
test_output[1491:1491] = '{32'h42df4bea};
test_input[11936:11943] = '{32'h415d761a, 32'h41ed060f, 32'hc113025a, 32'h42c59016, 32'h41e32483, 32'hc27da5cb, 32'hc28bb745, 32'h42c504e9};
test_weights[11936:11943] = '{32'hc2a381e0, 32'h3ee2b2d5, 32'hc24cc20e, 32'h42069205, 32'hc2654877, 32'h40886c2e, 32'hc2002b3c, 32'hc07f24a8};
test_bias[1492:1492] = '{32'h42b4f90a};
test_output[1492:1492] = '{32'h45299781};
test_input[11944:11951] = '{32'h42abbbf2, 32'hbfec5f05, 32'hc1e61aff, 32'h428f4cf3, 32'hc2bfe328, 32'hc1bfc7aa, 32'hc1566e4b, 32'hc2675b2a};
test_weights[11944:11951] = '{32'hc1e9964a, 32'hc1d59b61, 32'hc29836ef, 32'h41ba0d95, 32'hc2aed316, 32'h41eb3dbc, 32'hc2b16b92, 32'h42b9e7d6};
test_bias[1493:1493] = '{32'hc1b0c1f4};
test_output[1493:1493] = '{32'h45982e53};
test_input[11952:11959] = '{32'hc29d6bcd, 32'h418b598e, 32'hc1dc2dfa, 32'hc2c7ccb2, 32'h42ae6270, 32'h42b9f758, 32'h426e29c9, 32'hc2a70f49};
test_weights[11952:11959] = '{32'h42816ab9, 32'h42024a47, 32'h42ba0c62, 32'hc22c8de2, 32'hc243dcca, 32'h42bc5950, 32'h41de3c3a, 32'hc2913a9d};
test_bias[1494:1494] = '{32'hc1bdb0f3};
test_output[1494:1494] = '{32'h4612f997};
test_input[11960:11967] = '{32'h42854097, 32'h42b190ff, 32'hc2b117ce, 32'h4002d3b7, 32'hc292efe9, 32'h42544ab8, 32'h42333117, 32'h42447c1e};
test_weights[11960:11967] = '{32'hc2c67783, 32'h4283bc53, 32'hc0b5211b, 32'h42b83d22, 32'hc260c946, 32'hc1fbf535, 32'hc2a8950c, 32'h42a4393b};
test_bias[1495:1495] = '{32'hc29fd0b6};
test_output[1495:1495] = '{32'h4520089a};
test_input[11968:11975] = '{32'h428619a3, 32'h42a67989, 32'h417a7bd9, 32'h4242a8f7, 32'hc2334b3a, 32'hc29ee502, 32'h4273521f, 32'h416ab8da};
test_weights[11968:11975] = '{32'h40e46a68, 32'hc262ef77, 32'hc1ef4c3b, 32'hc26317f6, 32'h425f0286, 32'h420ca18b, 32'h42b1bf49, 32'hc22a0ce3};
test_bias[1496:1496] = '{32'h42702f42};
test_output[1496:1496] = '{32'hc5f7a47f};
test_input[11976:11983] = '{32'hc276ef36, 32'h42532e01, 32'hc1afe641, 32'h405adf5c, 32'hc29ae65e, 32'hc2270235, 32'hc2a29379, 32'hc2625393};
test_weights[11976:11983] = '{32'h41d66e6e, 32'hc17013b5, 32'hc19548e1, 32'hc229bb42, 32'h42a3bc0f, 32'hc2812a46, 32'h42016fa6, 32'hc29d9a7a};
test_bias[1497:1497] = '{32'hc2b09f60};
test_output[1497:1497] = '{32'hc57f5d6c};
test_input[11984:11991] = '{32'h42a8ba69, 32'h42a608e2, 32'h3fe6efe4, 32'hc1d821ad, 32'h41415d6f, 32'hc259cc14, 32'h413b0699, 32'hc2a79dc6};
test_weights[11984:11991] = '{32'h41aec8bb, 32'h41ac462b, 32'h41406111, 32'h40df557b, 32'h42a8d774, 32'hc2ae8c68, 32'hc1c46e9e, 32'h429aa099};
test_bias[1498:1498] = '{32'hc26e903c};
test_output[1498:1498] = '{32'h4516a257};
test_input[11992:11999] = '{32'h42a08e1e, 32'h423951a3, 32'h41a7ff01, 32'hc0cd6ae3, 32'h42c3da29, 32'hbf9513cf, 32'h429d3213, 32'h42c32192};
test_weights[11992:11999] = '{32'hc1b940ae, 32'h402bc895, 32'h418624ff, 32'hc08ead05, 32'hc295b689, 32'hc2b31b4c, 32'h4223e567, 32'h41b306e5};
test_bias[1499:1499] = '{32'h4235c666};
test_output[1499:1499] = '{32'hc543ab18};
test_input[12000:12007] = '{32'h3fbc7ac1, 32'hc18cbb52, 32'h42418877, 32'h42b16757, 32'hc2584a70, 32'h422ddf72, 32'hc27e767f, 32'h42a38bfe};
test_weights[12000:12007] = '{32'h41f2557e, 32'hc296e0a5, 32'hc1a6e857, 32'hc178fd53, 32'hc0f34bbc, 32'hc2825da7, 32'hc2a50e0c, 32'h42aaa8da};
test_bias[1500:1500] = '{32'h428a2cfb};
test_output[1500:1500] = '{32'h460a61c7};
test_input[12008:12015] = '{32'h423039d6, 32'hc28a3c72, 32'h41b2f587, 32'hc2bf616e, 32'h42176030, 32'h41dd997e, 32'h41e29f7d, 32'hc280eb0c};
test_weights[12008:12015] = '{32'h42a658c6, 32'hc2a2cd6e, 32'h42031f5c, 32'h41b45a0e, 32'h4246e7e6, 32'h41bf527d, 32'hc2a16f85, 32'hc2b99800};
test_bias[1501:1501] = '{32'h427ca9fd};
test_output[1501:1501] = '{32'h465d64b9};
test_input[12016:12023] = '{32'hc1d9a737, 32'h41c072b8, 32'h4082f584, 32'h429b153c, 32'h4295fd4a, 32'h42c034e6, 32'h4110bf55, 32'hc2a1f124};
test_weights[12016:12023] = '{32'hc28ee3dd, 32'h429e5e71, 32'hc0ca9062, 32'hc2c0831c, 32'hc24dcecd, 32'h4257fc21, 32'hc2275b8b, 32'h401c5fe8};
test_bias[1502:1502] = '{32'hc1a26ff3};
test_output[1502:1502] = '{32'hc535b29d};
test_input[12024:12031] = '{32'h416f4be7, 32'hc219f954, 32'hc2258c2b, 32'hc278a3d6, 32'hc13ac978, 32'hc15a21b4, 32'h4269cbdb, 32'hc1b77e06};
test_weights[12024:12031] = '{32'hc2c162cf, 32'h42435602, 32'hc21a476e, 32'hc18bc14d, 32'hc1982b4a, 32'h41df0d51, 32'h4225519f, 32'h42415e3a};
test_bias[1503:1503] = '{32'h424d465a};
test_output[1503:1503] = '{32'h440b18f4};
test_input[12032:12039] = '{32'h413615e7, 32'h42b17195, 32'hc225f855, 32'hc2c5581e, 32'h42a0a6c8, 32'h42b2ac12, 32'h4283f82b, 32'h40c2e4b9};
test_weights[12032:12039] = '{32'h423d97fc, 32'h423b4e76, 32'h421f5866, 32'h41711b61, 32'hc2877f40, 32'h418aa981, 32'h41b3de6f, 32'h40f95ac5};
test_bias[1504:1504] = '{32'h40b26f04};
test_output[1504:1504] = '{32'hc448b0ee};
test_input[12040:12047] = '{32'h42197075, 32'hc1911f5d, 32'h411027f3, 32'hc2ad9f37, 32'hc295f993, 32'hc2c1e816, 32'h41ba4d95, 32'hc242584d};
test_weights[12040:12047] = '{32'h42b1865c, 32'hc2a2e00e, 32'h4226b536, 32'h419a6846, 32'h426f5c83, 32'hc2b2275d, 32'hc2ab0f9a, 32'hc2c34958};
test_bias[1505:1505] = '{32'hc29ae61d};
test_output[1505:1505] = '{32'h46229833};
test_input[12048:12055] = '{32'h426ccac8, 32'h4291e0e2, 32'h4130ed52, 32'h42152d33, 32'h41d2997c, 32'h42354125, 32'hc2616937, 32'hc2709828};
test_weights[12048:12055] = '{32'h41fbcc97, 32'hc2b9ae9a, 32'h41c896fa, 32'h42bbc507, 32'hc2a5226c, 32'h42376218, 32'hc1c02c68, 32'h42a2575f};
test_bias[1506:1506] = '{32'hc202b8a5};
test_output[1506:1506] = '{32'hc5959a84};
test_input[12056:12063] = '{32'hc1989745, 32'hc2481c78, 32'hc1efc1c7, 32'h42901d6e, 32'h429385e9, 32'h42bd3a1b, 32'hc2c52df6, 32'hc2804c75};
test_weights[12056:12063] = '{32'hc243cb38, 32'hc2566a2f, 32'hc228db73, 32'h42a296bb, 32'hc2aef1fb, 32'h42ab4cbc, 32'h42bb1b4f, 32'h42c75633};
test_bias[1507:1507] = '{32'h4230b062};
test_output[1507:1507] = '{32'hc546f0ad};
test_input[12064:12071] = '{32'h4261cda8, 32'h42abe0fa, 32'h428e1d40, 32'h428b538c, 32'hc2a224a0, 32'hc28255a9, 32'h40d65e9b, 32'h40a51e40};
test_weights[12064:12071] = '{32'h42aa379b, 32'h42b1e506, 32'hc111c2ab, 32'h420d97a5, 32'h4241343b, 32'hc29421b8, 32'h4016c2e1, 32'hbf2f6363};
test_bias[1508:1508] = '{32'hc2890f1d};
test_output[1508:1508] = '{32'h466c46c6};
test_input[12072:12079] = '{32'h42b1685e, 32'h42adf22e, 32'h412352fa, 32'h427dbc1e, 32'h427b38f5, 32'h4207311d, 32'h41e41cd5, 32'hc0a449e2};
test_weights[12072:12079] = '{32'hc257c317, 32'hc21cc6fd, 32'hc2669738, 32'hc02f97d0, 32'hc2b78400, 32'hc1120fcb, 32'hc2932a4f, 32'hc043a447};
test_bias[1509:1509] = '{32'h4207482e};
test_output[1509:1509] = '{32'hc6856849};
test_input[12080:12087] = '{32'h400cd863, 32'h41f2703c, 32'hc21c5d36, 32'hc1a537d6, 32'h41e446e4, 32'hc2c544f4, 32'h42355ca1, 32'hc207d697};
test_weights[12080:12087] = '{32'hc2287889, 32'hc251b328, 32'h419cd7d3, 32'hc1e80ec8, 32'h423ea513, 32'hc289897d, 32'h41b52336, 32'h41e20eef};
test_bias[1510:1510] = '{32'h424e4609};
test_output[1510:1510] = '{32'h45c8663e};
test_input[12088:12095] = '{32'h42202724, 32'h4261ea83, 32'hc2b0e14c, 32'h40308826, 32'hc1948f34, 32'hc19196d0, 32'h414f7e28, 32'hc119c411};
test_weights[12088:12095] = '{32'hc0be16bf, 32'hc1ce5693, 32'h418675ed, 32'hc1f3ea4f, 32'hc296c4b0, 32'h423eddfd, 32'h41e59a07, 32'hc2876d1a};
test_bias[1511:1511] = '{32'hc24312ea};
test_output[1511:1511] = '{32'hc4dbee7e};
test_input[12096:12103] = '{32'h42be0d91, 32'hc1e21f60, 32'hc2a42aa1, 32'h41b5a2b9, 32'h41294346, 32'h3fb156ce, 32'h42c706c7, 32'h4254f981};
test_weights[12096:12103] = '{32'hc26164f1, 32'h41a94f79, 32'hc1aa417a, 32'hc20edf0f, 32'hc22bfd1a, 32'h41df75e9, 32'hc21fc861, 32'h42afa05d};
test_bias[1512:1512] = '{32'h40d645b5};
test_output[1512:1512] = '{32'hc593afba};
test_input[12104:12111] = '{32'h428def6e, 32'hc175b909, 32'h42a6ce7e, 32'h41dbe9ce, 32'h42531327, 32'h42bc6b46, 32'hc292bc7f, 32'h428902b9};
test_weights[12104:12111] = '{32'hc2b74320, 32'hc10be8ca, 32'h41a61530, 32'h42a62fa9, 32'h413d3de7, 32'hc2b86c8b, 32'h4266e761, 32'hc29b1ea2};
test_bias[1513:1513] = '{32'hc29e2b5d};
test_output[1513:1513] = '{32'hc69c973f};
test_input[12112:12119] = '{32'hc2b52e1c, 32'h42bee7df, 32'hc175211c, 32'h42afafae, 32'h42a38ff9, 32'hc29949fa, 32'h42813f30, 32'hc2943f5d};
test_weights[12112:12119] = '{32'h4287326f, 32'hc2813385, 32'hc010fcc0, 32'h425c7b9a, 32'h4104c3ca, 32'h42103442, 32'hc01ad70e, 32'hc085391d};
test_bias[1514:1514] = '{32'hc04bbfaa};
test_output[1514:1514] = '{32'hc6121354};
test_input[12120:12127] = '{32'hc250743c, 32'h40d8df2c, 32'h42a18a8b, 32'hc2071602, 32'hc1f98ad7, 32'hc0e40551, 32'h42c2f240, 32'h42087f90};
test_weights[12120:12127] = '{32'h421aca2d, 32'h4280a34f, 32'h42b43201, 32'h42837078, 32'hc230db51, 32'hc26e3ec7, 32'h409a8a53, 32'h429ac593};
test_bias[1515:1515] = '{32'hc28f9cdf};
test_output[1515:1515] = '{32'h46020136};
test_input[12128:12135] = '{32'hc25a0066, 32'hc24b351e, 32'h415b5c1d, 32'h42333c3d, 32'hc2bf442f, 32'hc2a7437a, 32'h419fd8e3, 32'h41d61b02};
test_weights[12128:12135] = '{32'h423c747f, 32'h42bbfac5, 32'h42bc683c, 32'h42a25502, 32'h415f8b75, 32'hc1fc72a6, 32'h429f7afa, 32'hc29cd2dc};
test_bias[1516:1516] = '{32'h42710e37};
test_output[1516:1516] = '{32'hc4c28508};
test_input[12136:12143] = '{32'hc29cd6db, 32'hc2b775c1, 32'h41e843cb, 32'h421673af, 32'hc2c037aa, 32'h41fb887b, 32'h429f0be7, 32'hc26cce8b};
test_weights[12136:12143] = '{32'h420f4225, 32'hc2197312, 32'hc285e1e3, 32'h41dd5161, 32'hc1ef9ded, 32'hc1454109, 32'hc0f92254, 32'hc232d9ad};
test_bias[1517:1517] = '{32'h42bad13d};
test_output[1517:1517] = '{32'h458a1eaf};
test_input[12144:12151] = '{32'h41ca40ba, 32'h40c5b350, 32'hc1bc9b86, 32'hc19dcf1f, 32'hc2abf45e, 32'hc2c62d0b, 32'hc21fe6dd, 32'h42c49fb6};
test_weights[12144:12151] = '{32'hc2213b34, 32'hc28e6cb0, 32'hc2c1593a, 32'hc2c202ae, 32'h42a9b984, 32'hc27db02d, 32'hc259b435, 32'h42aab55e};
test_bias[1518:1518] = '{32'hc0b2d0ce};
test_output[1518:1518] = '{32'h463fed38};
test_input[12152:12159] = '{32'hc2534a44, 32'h42935203, 32'h4261f57d, 32'hc1114f1f, 32'h42028c2c, 32'hc1c82d83, 32'hc215501c, 32'hc2840170};
test_weights[12152:12159] = '{32'h407539c3, 32'h423519ac, 32'h41ece30f, 32'hbf6affc7, 32'hc21d95d2, 32'h42a9afae, 32'h423813ed, 32'h42a5ce69};
test_bias[1519:1519] = '{32'h415ae802};
test_output[1519:1519] = '{32'hc5b458cf};
test_input[12160:12167] = '{32'h4101bb45, 32'hc2bac734, 32'hc2b15260, 32'h422f6825, 32'hc2a6d9c3, 32'hc2c4d872, 32'hbec36c1f, 32'h429f05af};
test_weights[12160:12167] = '{32'hbfc66995, 32'h4225107c, 32'h42175e0c, 32'h42b1171c, 32'h422c21c7, 32'h425cf7d5, 32'h3fc959b2, 32'h422331a3};
test_bias[1520:1520] = '{32'hc1754d36};
test_output[1520:1520] = '{32'hc60ec6e1};
test_input[12168:12175] = '{32'hc1bf8a85, 32'hc294afef, 32'h4138bd9e, 32'hc2b952ad, 32'h427ac0dc, 32'h41cbdfda, 32'hc11a5a68, 32'h42c2fc41};
test_weights[12168:12175] = '{32'hc29d7752, 32'hc28ae727, 32'hc27c145d, 32'hc0f17a21, 32'h40ee7964, 32'hc15999b7, 32'hc158ae64, 32'hc1eabc30};
test_bias[1521:1521] = '{32'h428355dc};
test_output[1521:1521] = '{32'h458be1c9};
test_input[12176:12183] = '{32'hc1efd9b8, 32'h4292a41c, 32'hc24e2d9d, 32'h3fe8c3b8, 32'h42a348ff, 32'hc1e8a7fc, 32'h420c27c4, 32'h42445a6d};
test_weights[12176:12183] = '{32'h42a329b3, 32'h42b642a8, 32'h41f3f81a, 32'h424cc9b7, 32'hc28dae16, 32'hc1fb7f22, 32'h428405cb, 32'h4210e9e7};
test_bias[1522:1522] = '{32'h411e9c85};
test_output[1522:1522] = '{32'h44f89e2b};
test_input[12184:12191] = '{32'h42ad3267, 32'h42b863e0, 32'hc272a99a, 32'h42576dc1, 32'h420a32aa, 32'hc24154d4, 32'hc2b28a76, 32'h42a7d135};
test_weights[12184:12191] = '{32'hc167fce1, 32'h40d5175c, 32'h4268e54f, 32'h42114562, 32'h41c556a4, 32'h41f8cad5, 32'h41d23bb2, 32'hc1b8bf48};
test_bias[1523:1523] = '{32'hc28cf415};
test_output[1523:1523] = '{32'hc5e1b75b};
test_input[12192:12199] = '{32'h419663b0, 32'hc2784892, 32'hc174e71c, 32'h4222d9b8, 32'h40f7424e, 32'h42abd4f9, 32'h412fb718, 32'h42a25bf4};
test_weights[12192:12199] = '{32'h40dbb37d, 32'hc1a6454b, 32'h42b56f7d, 32'h429fbe19, 32'hc1c52d28, 32'h3f7b4ab5, 32'h420ebb77, 32'hc295b866};
test_bias[1524:1524] = '{32'hc202d182};
test_output[1524:1524] = '{32'hc51edb5c};
test_input[12200:12207] = '{32'hc283602d, 32'h42bac45a, 32'h41fe587f, 32'hc1a1728c, 32'h4178e3ce, 32'hc250b676, 32'hc20e146e, 32'hc20eaea5};
test_weights[12200:12207] = '{32'hc299d0a9, 32'hc28c697f, 32'h409d940a, 32'h42686223, 32'hc2b99cdc, 32'hc25325aa, 32'h417af154, 32'h42776596};
test_bias[1525:1525] = '{32'h4203c5b2};
test_output[1525:1525] = '{32'hc5763c00};
test_input[12208:12215] = '{32'hc2b31691, 32'h4130c3df, 32'h4273133d, 32'h41c9ca26, 32'h4264d1a2, 32'hc29d11a9, 32'hc169f2ff, 32'h4234e796};
test_weights[12208:12215] = '{32'h416eab86, 32'hc139ed89, 32'hc2b4368c, 32'h40a65676, 32'h42939291, 32'hc286d7f3, 32'hbfb0fbcc, 32'h4218b93d};
test_bias[1526:1526] = '{32'hc107ed58};
test_output[1526:1526] = '{32'h458aeda4};
test_input[12216:12223] = '{32'hbe96ae85, 32'hc2294a58, 32'hc2202db5, 32'h42241937, 32'h429e6c4e, 32'h42123288, 32'h4280207f, 32'h41ab199f};
test_weights[12216:12223] = '{32'h41cdc917, 32'hc1b5d71e, 32'h41f68517, 32'h4288bd55, 32'hc20a58b6, 32'h42af2741, 32'hbf020734, 32'hbffd3e69};
test_bias[1527:1527] = '{32'h41ac81f7};
test_output[1527:1527] = '{32'h4537536b};
test_input[12224:12231] = '{32'hc18e88e1, 32'hc1f5bbb3, 32'hc1c55565, 32'hc152a58d, 32'h429130c1, 32'hc202d79c, 32'hc294ab31, 32'hc26e38a6};
test_weights[12224:12231] = '{32'hc1e023ba, 32'h4245db3c, 32'hc1929e13, 32'hc23aff52, 32'h422b8528, 32'hc2948a24, 32'h426acf2b, 32'hbffde797};
test_bias[1528:1528] = '{32'hc2418f45};
test_output[1528:1528] = '{32'h44a1f97a};
test_input[12232:12239] = '{32'h421192e2, 32'hc01aa0dd, 32'hc270167d, 32'h42adcbcb, 32'h42a73450, 32'hc182a75c, 32'hc28b4752, 32'h411e9d05};
test_weights[12232:12239] = '{32'hc29cb3a0, 32'hc2a712da, 32'hc2a1657c, 32'hc29eb0a2, 32'hc206db2a, 32'h4233fcfb, 32'hc2b5680f, 32'hc2b81823};
test_bias[1529:1529] = '{32'h423161a6};
test_output[1529:1529] = '{32'hc52f5f7d};
test_input[12240:12247] = '{32'h411ac7e6, 32'h3fc7ac16, 32'h42be0ded, 32'hc1f5ebfc, 32'h422f215c, 32'hc2b01a51, 32'h428df04d, 32'hc2311680};
test_weights[12240:12247] = '{32'h420e2171, 32'hc25a3f8a, 32'h42c72383, 32'hc2bc3e4c, 32'h422c5176, 32'h41ffc87d, 32'hc194065c, 32'hc2b76881};
test_bias[1530:1530] = '{32'h41818d5e};
test_output[1530:1530] = '{32'h4661be51};
test_input[12248:12255] = '{32'h426a51ce, 32'h429096a1, 32'h42b2d000, 32'hc26958a4, 32'h41d4314c, 32'h41abf8dc, 32'hc2c2997f, 32'h42bf14a7};
test_weights[12248:12255] = '{32'h425f9f52, 32'h42b84ab7, 32'hc1c84b2c, 32'hc244bcc3, 32'h4297bd44, 32'hc0c21297, 32'hbf92bb0e, 32'h428f54cb};
test_bias[1531:1531] = '{32'h4257562a};
test_output[1531:1531] = '{32'h46980b64};
test_input[12256:12263] = '{32'hc200e308, 32'hc258aa38, 32'hc292f94a, 32'h426e8d45, 32'hc2158796, 32'h422a4f13, 32'h42aec123, 32'hc29843d1};
test_weights[12256:12263] = '{32'hc283fb34, 32'h41b4969a, 32'h42bb8848, 32'h42b2f21c, 32'hc24f1f16, 32'h42a67cff, 32'h428bab0e, 32'h4213da71};
test_bias[1532:1532] = '{32'h4232c1c9};
test_output[1532:1532] = '{32'h45ff0bc3};
test_input[12264:12271] = '{32'h41a4801d, 32'h428e2033, 32'hc25ce00a, 32'hc26350b7, 32'hc199d1ef, 32'hc2afb8a6, 32'hc05290f6, 32'h422d0817};
test_weights[12264:12271] = '{32'hc2b6a10e, 32'hc28b1af7, 32'hc2bbea91, 32'hc20a0e21, 32'h420501c2, 32'hc29c06e0, 32'h42584b39, 32'hc23d975f};
test_bias[1533:1533] = '{32'hc29e8255};
test_output[1533:1533] = '{32'h458466a2};
test_input[12272:12279] = '{32'h42430dcb, 32'hc2b03975, 32'h416a7241, 32'h41ca57c7, 32'hc2980618, 32'hc27a9777, 32'h42132fe0, 32'h41d8be14};
test_weights[12272:12279] = '{32'hc2a598ed, 32'h41ffd457, 32'h42c3863d, 32'hc22e53c3, 32'hc2b891da, 32'h420fd761, 32'h3fc92be6, 32'hc1f698e4};
test_bias[1534:1534] = '{32'hc28dcfea};
test_output[1534:1534] = '{32'hc52335d9};
test_input[12280:12287] = '{32'hc1847ebf, 32'h42b4f581, 32'hc04edf87, 32'hc236f701, 32'h42ae3406, 32'h41cb34ea, 32'h412db888, 32'h420a3f8d};
test_weights[12280:12287] = '{32'h40fcbd5e, 32'hc2869561, 32'h41d25a3d, 32'hc147cb21, 32'h42104909, 32'hc1addc92, 32'h42976630, 32'h42800c8e};
test_bias[1535:1535] = '{32'hc289b6e3};
test_output[1535:1535] = '{32'hc3316f1f};
test_input[12288:12295] = '{32'hc2978e39, 32'hc1ccca9f, 32'hc28c714b, 32'h4298a78e, 32'hc224fe28, 32'h428f38b9, 32'hc109c633, 32'hc0ec273d};
test_weights[12288:12295] = '{32'hc2580edb, 32'hc2899db1, 32'hc2a79fb1, 32'h42bb6265, 32'hbfa20ed4, 32'hc1e1043e, 32'h429c61f1, 32'hc2b80ce0};
test_bias[1536:1536] = '{32'h42063fcd};
test_output[1536:1536] = '{32'h46849124};
test_input[12296:12303] = '{32'h41b267f0, 32'h425e9586, 32'hc1e0d08e, 32'h426af786, 32'hc22d95e5, 32'hc09230d0, 32'h42866c81, 32'h428f6055};
test_weights[12296:12303] = '{32'hc2b20a4b, 32'h41f0abb6, 32'hc1fed961, 32'h42a2f779, 32'h429cb2c4, 32'hc2c11978, 32'h426e6553, 32'hc28a6001};
test_bias[1537:1537] = '{32'hc2824b83};
test_output[1537:1537] = '{32'h44ae0715};
test_input[12304:12311] = '{32'h42b8a572, 32'hc28a2ff5, 32'h4229bab8, 32'h421aef35, 32'hc2423096, 32'hc17f5b73, 32'h421dfa90, 32'h425448da};
test_weights[12304:12311] = '{32'hc22291a0, 32'h4081072d, 32'h42bdc41a, 32'h41b1e54d, 32'hc2202c23, 32'hc13daa94, 32'h4216f607, 32'h42740bda};
test_bias[1538:1538] = '{32'hc28a51f3};
test_output[1538:1538] = '{32'h45ef090a};
test_input[12312:12319] = '{32'hc29f7788, 32'hc239d318, 32'hc285d8e0, 32'hc28c0192, 32'h42243a8b, 32'hbff47d58, 32'h420507a7, 32'h429aa2ec};
test_weights[12312:12319] = '{32'hc270c136, 32'hc18dbc3b, 32'h42abb696, 32'h420827da, 32'hc268dcba, 32'hc1371cf2, 32'h426b8033, 32'h41d6975e};
test_bias[1539:1539] = '{32'h42a9afa6};
test_output[1539:1539] = '{32'hc43d7fb9};
test_input[12320:12327] = '{32'hc26c497b, 32'hc234fc1e, 32'hc27594b4, 32'hc2201506, 32'hc2c26108, 32'hc2b9b300, 32'h41c13b2c, 32'hc1b17f4e};
test_weights[12320:12327] = '{32'hc1683319, 32'h42bc4ad8, 32'h42a6c00f, 32'hc1887018, 32'h42bfdb60, 32'h4215b4b7, 32'hc28807c9, 32'h401b9c2c};
test_bias[1540:1540] = '{32'h40965349};
test_output[1540:1540] = '{32'hc6ae7242};
test_input[12328:12335] = '{32'h426f71ed, 32'h420dec91, 32'hc280c5e1, 32'hbe2245fb, 32'hc25c9a35, 32'h4291e352, 32'hc01a39aa, 32'h42b90fe0};
test_weights[12328:12335] = '{32'h420bb34d, 32'h426635e9, 32'h42b1e8fa, 32'hc1b87b7d, 32'h40f60db7, 32'h429caa6b, 32'h42b185af, 32'h4256bf97};
test_bias[1541:1541] = '{32'hc28b52c4};
test_output[1541:1541] = '{32'h4602fb69};
test_input[12336:12343] = '{32'h41548f62, 32'hc206fd8b, 32'hc2a11229, 32'hc20d7698, 32'h427ac143, 32'h425ec111, 32'h429963ce, 32'h416fe3c9};
test_weights[12336:12343] = '{32'h42a6f7ae, 32'hc2acc417, 32'h42947157, 32'hc18c24ba, 32'hc0a88eae, 32'h423edd79, 32'hc248433d, 32'hc17c43a6};
test_bias[1542:1542] = '{32'hc25089c9};
test_output[1542:1542] = '{32'hc543ee15};
test_input[12344:12351] = '{32'h425387aa, 32'h42c07fcc, 32'h42008427, 32'h426247a7, 32'h428d25a4, 32'h4282e57e, 32'h41fcaa9f, 32'hc2970950};
test_weights[12344:12351] = '{32'hc2701492, 32'hc29e4b11, 32'h42b5bf3c, 32'hc2b32885, 32'h42c546d9, 32'h421500fc, 32'hc2c15239, 32'h42c25f51};
test_bias[1543:1543] = '{32'hc2867e2b};
test_output[1543:1543] = '{32'hc65abf43};
test_input[12352:12359] = '{32'h4224f9b7, 32'hc1c5f257, 32'h42c51dcd, 32'hc29093be, 32'hc22d936f, 32'hc2c7c9d9, 32'hc2a6b386, 32'hc14652ae};
test_weights[12352:12359] = '{32'h425bb65a, 32'hc289fd41, 32'h420b5912, 32'h4297f081, 32'h4211f1e2, 32'h42c0c768, 32'hc1a54fee, 32'h409b192b};
test_bias[1544:1544] = '{32'h4206c78e};
test_output[1544:1544] = '{32'hc5ed8dcd};
test_input[12360:12367] = '{32'hc23e8dca, 32'hc2781a22, 32'h3ff9274f, 32'hc1ac672a, 32'h41386ce6, 32'h42463962, 32'hc220d0b3, 32'h41d0a449};
test_weights[12360:12367] = '{32'hc296fdb0, 32'h4208de4b, 32'h429f7a08, 32'hc28637fd, 32'h42ae1be8, 32'hc20b3d36, 32'h4252ca63, 32'hc22717c5};
test_bias[1545:1545] = '{32'h428445af};
test_output[1545:1545] = '{32'hc444fd4a};
test_input[12368:12375] = '{32'hc29c9f4a, 32'h414f4dbf, 32'h42baedb5, 32'h421dba7a, 32'hc2682b1e, 32'h4084ede5, 32'hc23ffe18, 32'h426f9d9b};
test_weights[12368:12375] = '{32'hc1acd3f8, 32'h429cf966, 32'h4282a8d2, 32'h42694d8d, 32'hbfda2f72, 32'h4210ab51, 32'hc0e8b1dd, 32'hc23dc225};
test_bias[1546:1546] = '{32'h42bb35c3};
test_output[1546:1546] = '{32'h460c126d};
test_input[12376:12383] = '{32'hc1d18542, 32'hc18495ec, 32'hc2836737, 32'hbf89897a, 32'h4268d811, 32'hc21bc3e1, 32'h416b2353, 32'h41ae6973};
test_weights[12376:12383] = '{32'hc2665df1, 32'hc0e010af, 32'hc18e88b6, 32'hbfc19478, 32'hc1cd8e6d, 32'h41b6c94b, 32'hc1d80276, 32'h4281f597};
test_bias[1547:1547] = '{32'h419c0f92};
test_output[1547:1547] = '{32'h44b54fc5};
test_input[12384:12391] = '{32'h3fd82abb, 32'hc29bed37, 32'hc2869f46, 32'hc2bca852, 32'hc2a2804d, 32'h42c718e5, 32'hc0defd69, 32'hc22f32bc};
test_weights[12384:12391] = '{32'hc187bdb9, 32'h420708c5, 32'hc1b030c5, 32'hc1996813, 32'h42546988, 32'hc27161ad, 32'hc2b6e641, 32'hbf61a5d7};
test_bias[1548:1548] = '{32'hc244ae69};
test_output[1548:1548] = '{32'hc60da241};
test_input[12392:12399] = '{32'hc228b3cd, 32'hc23c55c7, 32'hc2833d34, 32'hc2ae2625, 32'hc22c607a, 32'hc26e69ad, 32'hc1f22de5, 32'h416b4d3b};
test_weights[12392:12399] = '{32'hc24e1bbb, 32'hc010fc8c, 32'h428c361b, 32'hc0282e41, 32'hc28150f2, 32'hc18c6861, 32'hc113a650, 32'h42aa3e6d};
test_bias[1549:1549] = '{32'h41d98b04};
test_output[1549:1549] = '{32'h454e33ae};
test_input[12400:12407] = '{32'h42252145, 32'h423870e6, 32'hc2c05c7e, 32'h41c92363, 32'h40358897, 32'hc26f3f35, 32'hc2810d1b, 32'hc2941853};
test_weights[12400:12407] = '{32'hc1d83932, 32'h428953cc, 32'hc296a4fd, 32'h41f9140f, 32'h411d007c, 32'h42b93a3e, 32'h41270b0e, 32'h42b98771};
test_bias[1550:1550] = '{32'hc2a7a115};
test_output[1550:1550] = '{32'hc53f45a2};
test_input[12408:12415] = '{32'h40b847e9, 32'hc2184c2f, 32'hbffe05a7, 32'h428c2c02, 32'h41bffd3f, 32'hc25c6fc7, 32'h42bb56cb, 32'h420e3da1};
test_weights[12408:12415] = '{32'h424a58a4, 32'h41ca8abf, 32'hc0f636f0, 32'hc04c5770, 32'h421a6ed3, 32'hc2ba42c1, 32'hc093f977, 32'hc22169eb};
test_bias[1551:1551] = '{32'hc2034bfd};
test_output[1551:1551] = '{32'h454ccca8};
test_input[12416:12423] = '{32'h42bc8c33, 32'h41f4256f, 32'h41610cc1, 32'h425a1dfc, 32'h421e7ce8, 32'h4285278f, 32'h4286cd4c, 32'hc24fb12c};
test_weights[12416:12423] = '{32'h416b1037, 32'hc2748bac, 32'hc2a4ebff, 32'h428cfda3, 32'h428fa12f, 32'h425afb11, 32'hc27794cd, 32'hc2c7f974};
test_bias[1552:1552] = '{32'hc2c2efae};
test_output[1552:1552] = '{32'h46164026};
test_input[12424:12431] = '{32'hc290eadd, 32'h41ade17a, 32'hc18b12a2, 32'h41e3d572, 32'h428450d8, 32'hc2b20fcb, 32'h41207bf5, 32'hc1fae05a};
test_weights[12424:12431] = '{32'hc271ebf6, 32'hc2816d6a, 32'h42b46a22, 32'hc280d3e4, 32'h4258c0a0, 32'hc1e9a28f, 32'h41fd17bf, 32'h426436f1};
test_bias[1553:1553] = '{32'hc287eb87};
test_output[1553:1553] = '{32'h4583d32a};
test_input[12432:12439] = '{32'h428c5ec1, 32'h41e80a8f, 32'h419e3f4f, 32'hc17106c9, 32'hc28ec105, 32'hc2b17367, 32'h4290d376, 32'hc1bc257d};
test_weights[12432:12439] = '{32'h41c43a82, 32'hc2163dc2, 32'h41a54cf4, 32'hc117b2b0, 32'hc1a778e1, 32'hc22b9ca8, 32'h42b46d95, 32'h4140a8e9};
test_bias[1554:1554] = '{32'hc1ec83cb};
test_output[1554:1554] = '{32'h4646816a};
test_input[12440:12447] = '{32'hc1879a6d, 32'h41baeafe, 32'hc2af10fe, 32'h42447bfb, 32'h42877daa, 32'hc1c44327, 32'h41d83b50, 32'h40c04579};
test_weights[12440:12447] = '{32'hc241b8ae, 32'hc1a7e0c5, 32'h41df9b85, 32'h4296b291, 32'h42025681, 32'hc29fb298, 32'h42bb3cb7, 32'hc101fca9};
test_bias[1555:1555] = '{32'h42c22fab};
test_output[1555:1555] = '{32'h460228fa};
test_input[12448:12455] = '{32'hc18d82af, 32'hbf829850, 32'hc2963a5c, 32'hc2963a81, 32'h3ff7091c, 32'h42ad05bd, 32'h409f0beb, 32'h42a4560d};
test_weights[12448:12455] = '{32'hbfd98ba5, 32'hc229279a, 32'hc07b878d, 32'hc166167e, 32'h42b5ff41, 32'h424f7529, 32'h422d509b, 32'h427f3523};
test_bias[1556:1556] = '{32'hc0ba3de8};
test_output[1556:1556] = '{32'h4634ac58};
test_input[12456:12463] = '{32'h42b82600, 32'h4112ce53, 32'hc2b489d3, 32'hc2807002, 32'hc28c5804, 32'hc093c8fd, 32'hc226bcb5, 32'hc2997163};
test_weights[12456:12463] = '{32'hc06bd7ff, 32'hc128015e, 32'hc088c54a, 32'hc0dc4528, 32'hc2b822c3, 32'hc1b77ec6, 32'h42bd2eca, 32'hc2828243};
test_bias[1557:1557] = '{32'h41f4edb9};
test_output[1557:1557] = '{32'h45fba649};
test_input[12464:12471] = '{32'hc2bc3766, 32'hc28485e2, 32'hc2c54a07, 32'h4294ad93, 32'hc2a1c179, 32'hc297f7d4, 32'hc1b66fd0, 32'hc233218f};
test_weights[12464:12471] = '{32'hc269cef8, 32'h4263453c, 32'h419aee1c, 32'h426ff0ae, 32'h42b0538a, 32'hc2a07f3a, 32'hbea2d9ea, 32'hc298c877};
test_bias[1558:1558] = '{32'h42ac289f};
test_output[1558:1558] = '{32'h45d372f1};
test_input[12472:12479] = '{32'h42bea419, 32'hc1c485c1, 32'h42a4fc6d, 32'hc2860183, 32'hc280f579, 32'h429b8197, 32'hc25ad061, 32'h41f837ac};
test_weights[12472:12479] = '{32'hc2beb94a, 32'h42a8a915, 32'h41df2df8, 32'hc285d3c5, 32'h4278ef7d, 32'hc2194bf7, 32'hc2a86b96, 32'h429af8f9};
test_bias[1559:1559] = '{32'h422ab230};
test_output[1559:1559] = '{32'hc586dfca};
test_input[12480:12487] = '{32'h413a6419, 32'hc240c401, 32'h41f0353b, 32'hc1df39c6, 32'hc24bfc0a, 32'h42595bfa, 32'h420190f0, 32'h418c2648};
test_weights[12480:12487] = '{32'hc255b895, 32'hc2454c83, 32'h4157d33a, 32'hc2219ea9, 32'h41cfb632, 32'hc240c815, 32'hc1ac35f2, 32'hc2844906};
test_bias[1560:1560] = '{32'h41abf7cb};
test_output[1560:1560] = '{32'hc51ba73e};
test_input[12488:12495] = '{32'hc282c210, 32'hc1fd5695, 32'h429baade, 32'h41558bbb, 32'h42239f95, 32'hc2683235, 32'h42898cea, 32'h426d5e51};
test_weights[12488:12495] = '{32'hc2965beb, 32'h42a6d136, 32'hc1b406d4, 32'h423b15fd, 32'h418815d2, 32'hc0cbeec9, 32'hc0a2f046, 32'hc1d48864};
test_bias[1561:1561] = '{32'hc0cfb310};
test_output[1561:1561] = '{32'h438b91d3};
test_input[12496:12503] = '{32'h40d8a526, 32'hc1eb0e1e, 32'hc231b06d, 32'h411ab3bc, 32'hc295f509, 32'h41e2e9cf, 32'h42a9f0d3, 32'h41ba68a0};
test_weights[12496:12503] = '{32'h4237c211, 32'h4237d3dc, 32'h423abde9, 32'hc1ae4d0d, 32'hc198a47b, 32'hc0f7e85c, 32'h424158c0, 32'hbf8ea1e6};
test_bias[1562:1562] = '{32'h409a4d64};
test_output[1562:1562] = '{32'h44f6a314};
test_input[12504:12511] = '{32'h4275ffa7, 32'hc1ea4451, 32'h42a45a75, 32'h42b8cd03, 32'hc1f4225a, 32'hc2af3ea7, 32'h42acdf59, 32'hc1c252bb};
test_weights[12504:12511] = '{32'h4203c919, 32'h4226b7b1, 32'h426c7ba8, 32'h41665536, 32'h41dc0f19, 32'hc2b142c9, 32'h40c9d882, 32'h42c331c6};
test_bias[1563:1563] = '{32'hc202190e};
test_output[1563:1563] = '{32'h463c7b28};
test_input[12512:12519] = '{32'hc2233147, 32'h42272ffc, 32'h423cd70e, 32'h427d1747, 32'hc200b656, 32'hc212ad38, 32'hc2a31c82, 32'h42beed8d};
test_weights[12512:12519] = '{32'h4295a3b9, 32'hc124959c, 32'h42a439cd, 32'h41cbce32, 32'h421e4938, 32'hc2ba5d25, 32'hc2c642d0, 32'hc201f68c};
test_bias[1564:1564] = '{32'hc23f550c};
test_output[1564:1564] = '{32'h460df2d5};
test_input[12520:12527] = '{32'h42a9a90d, 32'hc1d379dc, 32'hc2a71554, 32'hc21e06e8, 32'hc22ed26d, 32'h42bb0ad3, 32'hc2c56876, 32'hc0ac678c};
test_weights[12520:12527] = '{32'hc2b7387f, 32'h410226b6, 32'hc19ac8f2, 32'h424776b0, 32'h4138f914, 32'hc2194492, 32'h41a5a933, 32'h42ba36e1};
test_bias[1565:1565] = '{32'h42901217};
test_output[1565:1565] = '{32'hc668d903};
test_input[12528:12535] = '{32'hc259ec4a, 32'h42a5532d, 32'hc298bb29, 32'h4185c655, 32'hc2327975, 32'hc24051af, 32'h4194b59d, 32'hc12d9cbf};
test_weights[12528:12535] = '{32'h41956f97, 32'hc2c5bb13, 32'hc284ce81, 32'hc228b9e7, 32'hc2927a66, 32'h3f9be61e, 32'hc28fc6fa, 32'hc1a7a9fc};
test_bias[1566:1566] = '{32'hc2afc253};
test_output[1566:1566] = '{32'hc52fc129};
test_input[12536:12543] = '{32'h41b6eb8f, 32'hc17e3e74, 32'h41bbaba3, 32'h422edd66, 32'hc25ae522, 32'hc291fc14, 32'h428e67c9, 32'h414c6511};
test_weights[12536:12543] = '{32'hc19357f7, 32'hc2215f8a, 32'hc2363a2d, 32'hc29cf3e0, 32'h42c3797c, 32'hc176dd4c, 32'hc282ab33, 32'h42c2a7cf};
test_bias[1567:1567] = '{32'hc2740056};
test_output[1567:1567] = '{32'hc63b0dd9};
test_input[12544:12551] = '{32'h42278277, 32'hc19cac29, 32'hc214bc62, 32'hc2c56150, 32'hc29187e1, 32'hc240ace1, 32'h42bf8340, 32'h428408d8};
test_weights[12544:12551] = '{32'hc0fd4a9a, 32'h425b4960, 32'hc24499c8, 32'hc268d0ec, 32'h4204a710, 32'h41043fbb, 32'hc1a0a1cc, 32'h3f1e29e4};
test_bias[1568:1568] = '{32'h42a9022e};
test_output[1568:1568] = '{32'h44c2bf5b};
test_input[12552:12559] = '{32'hc22ab46f, 32'hc049d8d4, 32'hc2758d13, 32'h425fcd02, 32'hc1d65a4c, 32'hc233af27, 32'h40008d76, 32'h429f8a50};
test_weights[12552:12559] = '{32'hc29d7514, 32'hc1b72258, 32'hc142aa9e, 32'hc1a2ec67, 32'hc2a2087d, 32'h428bd2e1, 32'hc2638858, 32'hc0f1cc48};
test_bias[1569:1569] = '{32'hc0e5f3a6};
test_output[1569:1569] = '{32'h44a830b0};
test_input[12560:12567] = '{32'hc1c471ad, 32'h42907c14, 32'hc265827a, 32'hc2b7aa7c, 32'hc1839e88, 32'hc25150db, 32'hc0f26999, 32'h428634da};
test_weights[12560:12567] = '{32'h42809111, 32'h429aa526, 32'h42b541ab, 32'hc2b7bfae, 32'h425f6204, 32'hc2b7f6fa, 32'h4257a249, 32'h424fd08f};
test_bias[1570:1570] = '{32'hc1ea6795};
test_output[1570:1570] = '{32'h465daea5};
test_input[12568:12575] = '{32'h4035c371, 32'hc2a4c336, 32'hc23b60f2, 32'h42982540, 32'hc282d8b6, 32'hc17e55cc, 32'hc231f29e, 32'h40f011fa};
test_weights[12568:12575] = '{32'h3f9f73af, 32'hc2a80b1c, 32'h417cd55c, 32'hc13f60ef, 32'hc22e7c21, 32'h42195493, 32'h425de2de, 32'h41cf8c9b};
test_bias[1571:1571] = '{32'h421cbf14};
test_output[1571:1571] = '{32'h45a52e18};
test_input[12576:12583] = '{32'hc25d087f, 32'hc27ad3d8, 32'hc194436d, 32'h422af5ee, 32'h41e879d0, 32'h429e9c4c, 32'h42bff28d, 32'h42acb598};
test_weights[12576:12583] = '{32'h40b507c9, 32'hc2a6eb79, 32'hc23e3ef6, 32'hc27daaea, 32'hc260c8d0, 32'hc24baffa, 32'h4246d8ed, 32'h428a66d1};
test_bias[1572:1572] = '{32'hc27d728c};
test_output[1572:1572] = '{32'h45fd3fea};
test_input[12584:12591] = '{32'h40c0c076, 32'hc22542ac, 32'hc2780fd4, 32'h42a193be, 32'h40acd095, 32'h40ef60f6, 32'hc0bec620, 32'h4253f45c};
test_weights[12584:12591] = '{32'h42121813, 32'hc2b3cfc2, 32'h42807a4e, 32'h418e6677, 32'h40afe272, 32'h42b006ba, 32'hc2084cfc, 32'h42ada3aa};
test_bias[1573:1573] = '{32'hc1e2745a};
test_output[1573:1573] = '{32'h45d6208c};
test_input[12592:12599] = '{32'hc2a32846, 32'h42c262b8, 32'h429e775e, 32'h42866866, 32'h42ad9e19, 32'h40ccbcdc, 32'h429fba22, 32'h42b9b18d};
test_weights[12592:12599] = '{32'hc17589ae, 32'h42140909, 32'hc2838098, 32'h4268a56b, 32'hc219a10f, 32'hc25b0aab, 32'hc299284d, 32'h4252ce28};
test_bias[1574:1574] = '{32'hc1875fe7};
test_output[1574:1574] = '{32'hc4ac04d8};
test_input[12600:12607] = '{32'h42b3d884, 32'hc27b9bf3, 32'h428781dc, 32'h40a5f056, 32'h42a6d51e, 32'h41efc4c2, 32'h429a0503, 32'hc20d4c98};
test_weights[12600:12607] = '{32'hc18f80ec, 32'hc2bcf4a8, 32'h4104d7c6, 32'hc297fd9d, 32'hbf426561, 32'h429ad8ca, 32'h421603d4, 32'hc11b3cf1};
test_bias[1575:1575] = '{32'hc2058e92};
test_output[1575:1575] = '{32'h461b83ac};
test_input[12608:12615] = '{32'h42b675ff, 32'hc2b3e7a2, 32'hc24150ab, 32'h42c10cca, 32'h41e5acb8, 32'hc120f59b, 32'hc23c6609, 32'hc1b204ba};
test_weights[12608:12615] = '{32'hc18df931, 32'h429dbb1b, 32'h42496b02, 32'h4234825e, 32'h42368f81, 32'h4196ff7e, 32'hc212f4aa, 32'hc0e8a90c};
test_bias[1576:1576] = '{32'hc19076c6};
test_output[1576:1576] = '{32'hc56d44ad};
test_input[12616:12623] = '{32'h417d7b8f, 32'hc26b258e, 32'h419194d0, 32'h421231f1, 32'h40ef9279, 32'hc242cdfc, 32'hc1f3f5e0, 32'hc25c75d9};
test_weights[12616:12623] = '{32'hc0d3918a, 32'h42961bce, 32'hc1b29284, 32'hc28b15ea, 32'hc2bb9d9a, 32'h428b8540, 32'hc16dd3ff, 32'h422f4235};
test_bias[1577:1577] = '{32'hc2aba321};
test_output[1577:1577] = '{32'hc654afb9};
test_input[12624:12631] = '{32'h42a69943, 32'h42a6058f, 32'hc1baf864, 32'h41408fdc, 32'hc2017302, 32'hc1fc6949, 32'h428760b2, 32'hc2b6d401};
test_weights[12624:12631] = '{32'h4287d2ad, 32'hc077db90, 32'hc18b595b, 32'hbff846ef, 32'h41ff421d, 32'hc2b3648c, 32'h429611d9, 32'h41672182};
test_bias[1578:1578] = '{32'h42a4b27a};
test_output[1578:1578] = '{32'h46317628};
test_input[12632:12639] = '{32'hc29d9208, 32'hbfc62698, 32'h40f43095, 32'hc217626b, 32'h4216cbb2, 32'hc1148872, 32'hc2896183, 32'hc2504282};
test_weights[12632:12639] = '{32'hc18b4996, 32'h41e7115a, 32'h3e86111a, 32'hc2c47fd8, 32'h423b47b2, 32'hc2bdc9ae, 32'h42a4f2f7, 32'hc038c99b};
test_bias[1579:1579] = '{32'h4081bf33};
test_output[1579:1579] = '{32'h450868a2};
test_input[12640:12647] = '{32'hc282ea2b, 32'hc2bdf45d, 32'h4285e928, 32'h4273606a, 32'hc257e5ea, 32'h426ebc42, 32'hc21a080c, 32'hc2903f93};
test_weights[12640:12647] = '{32'h4197a6cb, 32'h418dc2b3, 32'h42b18824, 32'hc20972dc, 32'h3e4fcaa6, 32'hc25954aa, 32'h4299c45c, 32'h426b74bd};
test_bias[1580:1580] = '{32'h42691baf};
test_output[1580:1580] = '{32'hc6140348};
test_input[12648:12655] = '{32'hbf11a6b0, 32'hc1d20a71, 32'hc1719c12, 32'h423eb356, 32'hc2a4189e, 32'h426c842b, 32'hc1091a0a, 32'h427382d9};
test_weights[12648:12655] = '{32'h41cd335c, 32'h4121e1c1, 32'hc2b19db8, 32'h428147bc, 32'hc1e9436b, 32'hc2a3d21c, 32'h42634824, 32'hbddc308e};
test_bias[1581:1581] = '{32'h42b86c19};
test_output[1581:1581] = '{32'h44a14ca4};
test_input[12656:12663] = '{32'hc29ba4a2, 32'hc217291f, 32'hc2aaaa09, 32'hc223fc1c, 32'hc2c15e8a, 32'hc28d846b, 32'hc265d479, 32'h42bcc519};
test_weights[12656:12663] = '{32'hc1c23ab0, 32'h4269c2a0, 32'hc26fc14c, 32'hc116febe, 32'h4244223f, 32'h419b1e15, 32'h423e0598, 32'hc20c7b5c};
test_bias[1582:1582] = '{32'h427a04fc};
test_output[1582:1582] = '{32'hc5d800f4};
test_input[12664:12671] = '{32'hc2319b2d, 32'hc154368b, 32'hc29c6a48, 32'h42a21ee6, 32'h4153df0d, 32'h42ba6b67, 32'hc283e181, 32'hc2704888};
test_weights[12664:12671] = '{32'hc1218f00, 32'h42b745c8, 32'h4232ac92, 32'h4242a3dd, 32'h42b69766, 32'h4207adad, 32'h42ae3910, 32'hc26cc5f7};
test_bias[1583:1583] = '{32'h40d33fb5};
test_output[1583:1583] = '{32'h44ea1706};
test_input[12672:12679] = '{32'hc2ac85b4, 32'hc2b14cf5, 32'h41c7aa2f, 32'hc25017ec, 32'h42a89e1e, 32'h4204f6e6, 32'hc23a4d6c, 32'h41b8e50e};
test_weights[12672:12679] = '{32'h42c3ce3e, 32'h42be12df, 32'hc27f757b, 32'h42aa33fb, 32'h3deda9ec, 32'h42538ce8, 32'hc2931827, 32'h4203cbe1};
test_bias[1584:1584] = '{32'h4215e0cb};
test_output[1584:1584] = '{32'hc684064d};
test_input[12680:12687] = '{32'h42a43094, 32'hc268e7ed, 32'hc237e55b, 32'hc238102a, 32'h40937b6a, 32'hc23b4390, 32'hc29ef559, 32'hc16511a3};
test_weights[12680:12687] = '{32'h42b55d31, 32'h42803668, 32'h41bd5edf, 32'hbf63075a, 32'hc1f58f2d, 32'hc067a6a3, 32'h4290f847, 32'h41d4a5a4};
test_bias[1585:1585] = '{32'h41c7b8ff};
test_output[1585:1585] = '{32'hc5560419};
test_input[12688:12695] = '{32'h42b12c8d, 32'h423b7509, 32'h42bb674a, 32'hc22c6c55, 32'h4292add0, 32'h4084491b, 32'h420f2dc8, 32'hc2b1e659};
test_weights[12688:12695] = '{32'h42b2c01f, 32'h417fc926, 32'hc0c9699a, 32'h4284c5b5, 32'h41a9af8b, 32'hbfc63b76, 32'hc1f5a133, 32'hc21fc368};
test_bias[1586:1586] = '{32'hc2936fa8};
test_output[1586:1586] = '{32'h460ee1ce};
test_input[12696:12703] = '{32'h42c71d4f, 32'h42565124, 32'h42ae64e0, 32'h428f1855, 32'hc25b6ff6, 32'hc26fab83, 32'hc2b14580, 32'h4203da42};
test_weights[12696:12703] = '{32'hc2a9b1f6, 32'hc2148d7a, 32'h42c20c10, 32'h42ad8e2f, 32'hc27fcf8a, 32'hc28aa2df, 32'h429d3bef, 32'h41f0e328};
test_bias[1587:1587] = '{32'h418af51a};
test_output[1587:1587] = '{32'h45b97a36};
test_input[12704:12711] = '{32'h41d5dab0, 32'h426e6da9, 32'h42b02099, 32'hc2b596c8, 32'hc1f247e7, 32'h41bd3109, 32'h4296338c, 32'hc2b222bc};
test_weights[12704:12711] = '{32'hc2847ac2, 32'h4220fd48, 32'h42b9b3f6, 32'hc254f00c, 32'hc260cc86, 32'h41852a1c, 32'h421ced40, 32'hc19aa0d8};
test_bias[1588:1588] = '{32'h42bc888b};
test_output[1588:1588] = '{32'h46a020ba};
test_input[12712:12719] = '{32'h4293cd45, 32'hc2260e25, 32'h41cd1447, 32'hc1870660, 32'h425c3fc1, 32'h42b518af, 32'hc260aff1, 32'h42c769ef};
test_weights[12712:12719] = '{32'hc0730488, 32'h42b39857, 32'h427bdeec, 32'h412510d0, 32'h422083c2, 32'h42c5145d, 32'hc29338eb, 32'hbe34d887};
test_bias[1589:1589] = '{32'h42525a79};
test_output[1589:1589] = '{32'h4646f67d};
test_input[12720:12727] = '{32'hc2b122cb, 32'h4246e619, 32'hc0188f0c, 32'h415e6c67, 32'h415fbada, 32'hc2a30360, 32'hc1c2f70a, 32'h41ae1b2a};
test_weights[12720:12727] = '{32'h424afa22, 32'h418ece34, 32'hc1a3a036, 32'h42172e0b, 32'h42b9b6a8, 32'hc2b5ab6c, 32'h4176c107, 32'hc2a53ae2};
test_bias[1590:1590] = '{32'hc104baf0};
test_output[1590:1590] = '{32'h4559f699};
test_input[12728:12735] = '{32'h425fa7ab, 32'h42ac7d7b, 32'h42783135, 32'h42b2223f, 32'h418a6600, 32'hc293f1e7, 32'h428274f6, 32'h428b266f};
test_weights[12728:12735] = '{32'hc125843c, 32'hc2a2f924, 32'hc18ec139, 32'h421f1002, 32'h42a7e9a6, 32'h412e5262, 32'h42a208a2, 32'hc29eeb77};
test_bias[1591:1591] = '{32'hc2036b75};
test_output[1591:1591] = '{32'hc5960ea0};
test_input[12736:12743] = '{32'h425c07bd, 32'h427bc09e, 32'h426665e0, 32'hc2bfe052, 32'hc170de01, 32'hc2973663, 32'hc2becb03, 32'h429356d8};
test_weights[12736:12743] = '{32'h42a0c2fc, 32'hc08daf30, 32'h42ae4279, 32'h41be7e1d, 32'hc2607390, 32'hc22163d6, 32'h4284a510, 32'h42a4addc};
test_bias[1592:1592] = '{32'hc1cb5143};
test_output[1592:1592] = '{32'h4623d7b0};
test_input[12744:12751] = '{32'h4265046f, 32'h41d947a9, 32'h42c48c6c, 32'h42bccd16, 32'h41bf5a02, 32'hc1a7efdb, 32'hc1ab3b0c, 32'hc2c277a8};
test_weights[12744:12751] = '{32'hc2c5a354, 32'hc2b1b391, 32'hbf6630e9, 32'hc1a95b76, 32'hc297d813, 32'hc2ba8f6c, 32'h42990028, 32'hc196376f};
test_bias[1593:1593] = '{32'h41074957};
test_output[1593:1593] = '{32'hc6196b36};
test_input[12752:12759] = '{32'h4292dc13, 32'hc205f691, 32'hc2a2c498, 32'h42305a8a, 32'h410b3c9a, 32'hc2899617, 32'h40e21641, 32'h4211aaf6};
test_weights[12752:12759] = '{32'h429dd217, 32'h429e0b99, 32'h418bec85, 32'hc2244dd8, 32'hc23c0be2, 32'hc1fad794, 32'hc226c51e, 32'hc193f761};
test_bias[1594:1594] = '{32'hc29d4010};
test_output[1594:1594] = '{32'h4419a57f};
test_input[12760:12767] = '{32'h425b473e, 32'h424a42ec, 32'h41b6d138, 32'h4284b5fb, 32'hc211f293, 32'hc2439971, 32'hc1ab87b0, 32'h42b9bc71};
test_weights[12760:12767] = '{32'h420d31de, 32'hc2bd10a5, 32'hc28c9c82, 32'hc0d203c4, 32'hc20dba9f, 32'hc2a382be, 32'h420d1cd9, 32'hc2b8db05};
test_bias[1595:1595] = '{32'hc29ada2e};
test_output[1595:1595] = '{32'hc60cd7ae};
test_input[12768:12775] = '{32'h41fadcd6, 32'h4297999b, 32'h422b4063, 32'h425637f8, 32'h4204f1e8, 32'hc1b660b9, 32'hc2b19c04, 32'hc2602c34};
test_weights[12768:12775] = '{32'h417075a9, 32'h42bfcfbf, 32'h42acf895, 32'h422b936a, 32'h42131334, 32'hc2b32a55, 32'h425216f1, 32'h428e1532};
test_bias[1596:1596] = '{32'h42c6729f};
test_output[1596:1596] = '{32'h46042abc};
test_input[12776:12783] = '{32'hc1f6fbc7, 32'h41441399, 32'hc1c6595e, 32'hc1166633, 32'h4192a888, 32'h42946b89, 32'hc2979680, 32'h42c33621};
test_weights[12776:12783] = '{32'h42bf7188, 32'h42a066ee, 32'hc20f2516, 32'h41cf3778, 32'h403e2a8c, 32'hc111d4f8, 32'h418422f3, 32'hc29f60ae};
test_bias[1597:1597] = '{32'h42960ac3};
test_output[1597:1597] = '{32'hc62a65c8};
test_input[12784:12791] = '{32'hc299e184, 32'h428961f8, 32'h41c88f27, 32'hc2a4677b, 32'hc2c792c2, 32'hc19972d6, 32'h42834c89, 32'h419318ea};
test_weights[12784:12791] = '{32'h42978bf6, 32'h421eddac, 32'h416d1ac9, 32'hc17826b9, 32'hc28179f0, 32'hc1312792, 32'hc2b5656e, 32'hc2a55142};
test_bias[1598:1598] = '{32'hc23fab4b};
test_output[1598:1598] = '{32'hc51011e8};
test_input[12792:12799] = '{32'hc1655cc3, 32'h4018a8ab, 32'hc1e61b08, 32'h429c1c12, 32'hc2a9671c, 32'hc0c7e2a4, 32'h41f84635, 32'hc216a0b6};
test_weights[12792:12799] = '{32'hc23aa1bb, 32'hc26e069d, 32'hc2481e67, 32'hc2c089a2, 32'hc245a01a, 32'h418b1dad, 32'h426ccbc6, 32'hc1bd3811};
test_bias[1599:1599] = '{32'hc286ab24};
test_output[1599:1599] = '{32'h44948c2e};
test_input[12800:12807] = '{32'hc1d86950, 32'hc2b2ef64, 32'hc1a645ab, 32'hc1bf8e00, 32'h41a368b9, 32'h41d711c3, 32'h42784c71, 32'hc239977b};
test_weights[12800:12807] = '{32'h42580818, 32'h42931a38, 32'h406b776e, 32'hc1bfebe3, 32'hc242e53e, 32'h41a8d6d5, 32'hc2739f3f, 32'hc2507043};
test_bias[1600:1600] = '{32'h42223720};
test_output[1600:1600] = '{32'hc61136c8};
test_input[12808:12815] = '{32'hc18ff789, 32'hc2b19aaf, 32'hc201a868, 32'hc16ece0d, 32'h42a5de92, 32'h4288cace, 32'h41dbc0eb, 32'h42460dda};
test_weights[12808:12815] = '{32'h41bfa856, 32'h41b93615, 32'h42a5bd0b, 32'h42658936, 32'hc26ceb92, 32'h4199876a, 32'h3f02c59e, 32'hc2b2ea40};
test_bias[1601:1601] = '{32'h429b2030};
test_output[1601:1601] = '{32'hc65a3c34};
test_input[12816:12823] = '{32'hc2c6cc19, 32'h40d8e418, 32'hc1f6e586, 32'hc1d11df3, 32'h41c7380e, 32'h42bf1de1, 32'hc0f91335, 32'hc28f29fb};
test_weights[12816:12823] = '{32'h41640139, 32'h42996996, 32'hc2066ea2, 32'h411051b8, 32'h424752a7, 32'hc28df639, 32'h41a4fc43, 32'hc297ec52};
test_bias[1602:1602] = '{32'hc2ac8484};
test_output[1602:1602] = '{32'hc3df2b56};
test_input[12824:12831] = '{32'h429bc118, 32'h42c27a0c, 32'h41ba422e, 32'hc2a37767, 32'hc016454f, 32'hc1832add, 32'hc19ff8c9, 32'h4190565f};
test_weights[12824:12831] = '{32'hc2a26d2e, 32'hc1a382ab, 32'h421b86fd, 32'h41aac25e, 32'hc21c970f, 32'h42c68dda, 32'h414eb168, 32'hc2bd2e2d};
test_bias[1603:1603] = '{32'hc2ac1191};
test_output[1603:1603] = '{32'hc64708d6};
test_input[12832:12839] = '{32'hc22f3d03, 32'hc229d34a, 32'h40c8b078, 32'h42830695, 32'hc218e901, 32'hc2a93f35, 32'h42b22d24, 32'h41b46ebe};
test_weights[12832:12839] = '{32'h42b1c420, 32'hc20bf674, 32'hc236283b, 32'hc2b877d8, 32'hc2c3a0c2, 32'h42bbfaf1, 32'h42434843, 32'h3ed1e262};
test_bias[1604:1604] = '{32'h42c2feb2};
test_output[1604:1604] = '{32'hc604bbe6};
test_input[12840:12847] = '{32'h42a8d49a, 32'h42add332, 32'hc2903152, 32'hc0bd4839, 32'h42b31262, 32'hc29e49a5, 32'h42c07555, 32'hc29a9592};
test_weights[12840:12847] = '{32'hc1ed5454, 32'h4261926e, 32'h427f7190, 32'h41ac6e6d, 32'hc12346dd, 32'hc2b3eca3, 32'hc25ae590, 32'hc099dd09};
test_bias[1605:1605] = '{32'hc2149395};
test_output[1605:1605] = '{32'hc4847eca};
test_input[12848:12855] = '{32'h42c68bed, 32'h41e1edc8, 32'h4194bfc6, 32'h420169ac, 32'h4200d7f6, 32'hc1b0d24e, 32'hc21c281e, 32'hc29f6051};
test_weights[12848:12855] = '{32'h40429bd4, 32'hc2a9fbbb, 32'hc0dec2d9, 32'hc20d890b, 32'h41d2094b, 32'h42a0b748, 32'h4283b10c, 32'h40fec73a};
test_bias[1606:1606] = '{32'hc2a0474d};
test_output[1606:1606] = '{32'hc5ed21c2};
test_input[12856:12863] = '{32'h428a55a9, 32'hc1d61bf0, 32'h41417bda, 32'hc2884a4a, 32'hc28ee7b3, 32'hc21b2c7e, 32'h413213b3, 32'h42c3113e};
test_weights[12856:12863] = '{32'h42642827, 32'hc201c8d5, 32'hc2c1a040, 32'h419ae53a, 32'hc290913b, 32'hc24fd91d, 32'h42b659e6, 32'h428dde40};
test_bias[1607:1607] = '{32'h41d2ea45};
test_output[1607:1607] = '{32'h46886f67};
test_input[12864:12871] = '{32'h420fc09a, 32'hc1006faf, 32'hc2962c1f, 32'hc2b5f0e8, 32'hc225b8ba, 32'h421e7283, 32'hc25aef0c, 32'hc209cab4};
test_weights[12864:12871] = '{32'hc0cbca19, 32'hc20fdada, 32'h41aa5309, 32'hc2b3a223, 32'hc25f575a, 32'hc2c27c72, 32'h429ac118, 32'h42c1499b};
test_bias[1608:1608] = '{32'hc21d4f9c};
test_output[1608:1608] = '{32'hc51ce749};
test_input[12872:12879] = '{32'h42a81e23, 32'h419ab665, 32'h41ef74f2, 32'h41809898, 32'h413cf6c3, 32'hc050da5f, 32'hc1b5d5f2, 32'hc2650b7b};
test_weights[12872:12879] = '{32'h413db284, 32'h403bd400, 32'hc2294c88, 32'h40e460c7, 32'h420a350d, 32'hc2aad5fd, 32'h42b95d79, 32'h4281cb59};
test_bias[1609:1609] = '{32'h42aeee1f};
test_output[1609:1609] = '{32'hc5a0d9c3};
test_input[12880:12887] = '{32'hc2c0f85d, 32'h42c721f1, 32'hc0c3b802, 32'h42a7ced2, 32'hc2bf6847, 32'h426092b1, 32'hc2802bf5, 32'h40da355a};
test_weights[12880:12887] = '{32'h424ae0b5, 32'hc29ab18c, 32'h42b1b172, 32'hc174432a, 32'h42c07afa, 32'hc20fa560, 32'h4282718d, 32'hc2612dbd};
test_bias[1610:1610] = '{32'hc24b578d};
test_output[1610:1610] = '{32'hc6ec68b2};
test_input[12888:12895] = '{32'h429aa563, 32'h423ea460, 32'h42543ae8, 32'h42bc4ae9, 32'hc25ea378, 32'h4120b45e, 32'h422edbea, 32'hc204e572};
test_weights[12888:12895] = '{32'hc25ce95e, 32'hc10c56bd, 32'hc0206ac4, 32'hc28b9c8c, 32'hc19ee65a, 32'hc291ad38, 32'h429907ba, 32'h402f9fdb};
test_bias[1611:1611] = '{32'hc238a5e9};
test_output[1611:1611] = '{32'hc5f41f58};
test_input[12896:12903] = '{32'hc278b5ac, 32'hc2b9bb6d, 32'hc18bf06f, 32'h4171da48, 32'hc287a7b1, 32'h4288b89e, 32'h420457d7, 32'h4245b4c6};
test_weights[12896:12903] = '{32'hc28572ac, 32'h420ca773, 32'h41e73de1, 32'h4232749c, 32'hc1ab4436, 32'hc1d77abc, 32'hc2bc5def, 32'hbeca820e};
test_bias[1612:1612] = '{32'hc2ab85ca};
test_output[1612:1612] = '{32'hc51feae5};
test_input[12904:12911] = '{32'h42955b3a, 32'h42b1adbf, 32'h42938ab7, 32'hc23b1a42, 32'hc23fec7d, 32'h42256329, 32'hc2c6b639, 32'hc12d261e};
test_weights[12904:12911] = '{32'h41cdc861, 32'h4186b5e3, 32'hc227617a, 32'hc2859e18, 32'h4094f784, 32'hc28ff242, 32'hc2540c67, 32'h42b016ae};
test_bias[1613:1613] = '{32'h429a74d2};
test_output[1613:1613] = '{32'h459139c6};
test_input[12912:12919] = '{32'hc0b399af, 32'h40f1faf8, 32'hc2a230cf, 32'hc2ab4fb1, 32'h41aa3a1a, 32'hc1ff9873, 32'hc120aa2e, 32'h4228e852};
test_weights[12912:12919] = '{32'hc23b3862, 32'hc260bcae, 32'h42bb96e4, 32'hc26ccf3b, 32'h429fbbbc, 32'h413ca787, 32'h40d5a429, 32'h42c09e8b};
test_bias[1614:1614] = '{32'hc12504a9};
test_output[1614:1614] = '{32'h45236c2e};
test_input[12920:12927] = '{32'hc29e7946, 32'h429c1fc4, 32'h4277e1ef, 32'hc1ba30c9, 32'hc138bd74, 32'hc21e1346, 32'hc28c7d3a, 32'hc19d6587};
test_weights[12920:12927] = '{32'h42355651, 32'h427fd9fe, 32'hc2433f3f, 32'h4203278d, 32'hc1f20077, 32'h4251113a, 32'h41d75003, 32'hc2a7421b};
test_bias[1615:1615] = '{32'h42844d5a};
test_output[1615:1615] = '{32'hc585d30f};
test_input[12928:12935] = '{32'hc2c56bdd, 32'h42b86923, 32'hc2611edf, 32'hc1e03db1, 32'hc0002945, 32'hc10808d4, 32'h424ee89e, 32'hc144b79c};
test_weights[12928:12935] = '{32'hc286fee9, 32'hc1152acb, 32'h42914332, 32'hc2a5fbbd, 32'hc112da72, 32'hc03915bf, 32'h40df4fdf, 32'h423219ee};
test_bias[1616:1616] = '{32'h42c4155d};
test_output[1616:1616] = '{32'h4579c42d};
test_input[12936:12943] = '{32'hc28d8db3, 32'hc03c01da, 32'h4289a182, 32'hc198f0df, 32'hc17015b5, 32'h4240f1bb, 32'hc2841d2a, 32'hbea8624d};
test_weights[12936:12943] = '{32'hc2908055, 32'hc2889fbe, 32'h41a64089, 32'hc2a0bdbb, 32'h412b8093, 32'h42067ffa, 32'h41572f48, 32'hc1824da9};
test_bias[1617:1617] = '{32'hc2aa966a};
test_output[1617:1617] = '{32'h460916b8};
test_input[12944:12951] = '{32'hc29cbfc4, 32'hc251702c, 32'h42247967, 32'h40110915, 32'hc1744a24, 32'hc2948435, 32'h42a29739, 32'hc2a2218d};
test_weights[12944:12951] = '{32'h424c2ad8, 32'h42bff6f8, 32'hc011902e, 32'hc2a695df, 32'h42291283, 32'h3fb28955, 32'hbec048dc, 32'hc29cbeaa};
test_bias[1618:1618] = '{32'h42b38e0b};
test_output[1618:1618] = '{32'hc563ca27};
test_input[12952:12959] = '{32'hc29d5e6d, 32'h427e12f0, 32'h42354fa2, 32'h42b3ebb4, 32'hc286f3c2, 32'h3ed24173, 32'hc297e2f4, 32'hc2c1861c};
test_weights[12952:12959] = '{32'hc2060b87, 32'h42be49d2, 32'hc22242e3, 32'hc158f482, 32'hc28c09ea, 32'hc271b990, 32'hc1f2f26d, 32'hc27c29f5};
test_bias[1619:1619] = '{32'hc0bc14fb};
test_output[1619:1619] = '{32'h469243ac};
test_input[12960:12967] = '{32'h429cb7eb, 32'hc2b7083a, 32'h420cd4fe, 32'h421eca50, 32'h424c2c12, 32'hc07cd388, 32'h4123c95e, 32'hc2a67e66};
test_weights[12960:12967] = '{32'h42b78dbb, 32'h41dae537, 32'h4228ddb7, 32'h40941e5e, 32'h41e06c56, 32'hc279f9cc, 32'hc21210ca, 32'hc2ac061a};
test_bias[1620:1620] = '{32'h424260b0};
test_output[1620:1620] = '{32'h46685d9e};
test_input[12968:12975] = '{32'hc1b9f83a, 32'hc243d221, 32'hc2b55ef1, 32'h42b42417, 32'h42254a28, 32'hbffaa025, 32'h41b0e20a, 32'hc1d8cfbc};
test_weights[12968:12975] = '{32'h4277ff6f, 32'hc17f3720, 32'hc294e0d7, 32'h42255b1b, 32'h42190eeb, 32'h423a481d, 32'h424482c5, 32'hc1fd4ae7};
test_bias[1621:1621] = '{32'h4283d341};
test_output[1621:1621] = '{32'h46500743};
test_input[12976:12983] = '{32'hc160aa8d, 32'h4290a862, 32'h415a7d1d, 32'h4219ea27, 32'h42af0664, 32'hc1e44999, 32'hc29d4897, 32'hc19847d4};
test_weights[12976:12983] = '{32'hc27a32f0, 32'h42ba2b12, 32'h42be3708, 32'h41cfcb9f, 32'h42a11435, 32'h42c4cc8b, 32'h41e16faa, 32'h424517c2};
test_bias[1622:1622] = '{32'h42b41602};
test_output[1622:1622] = '{32'h462d3600};
test_input[12984:12991] = '{32'hc141bd58, 32'h40e6fc41, 32'h427a9b98, 32'hc1063000, 32'h42812917, 32'h42b37fa1, 32'hc28690a6, 32'hc28cdb78};
test_weights[12984:12991] = '{32'hc25c2ee1, 32'hc250d94a, 32'h429da354, 32'hc2020730, 32'h4222aefa, 32'h4273688f, 32'h421575f0, 32'h42848d46};
test_bias[1623:1623] = '{32'h425b5109};
test_output[1623:1623] = '{32'h45c9ebf1};
test_input[12992:12999] = '{32'h4251e466, 32'hc2b4807b, 32'hc1b385c3, 32'h4263108b, 32'hc28672e5, 32'h42b032af, 32'hc20fbc5b, 32'hc22ab997};
test_weights[12992:12999] = '{32'h4289116e, 32'hc29c7d33, 32'hc2a44b31, 32'h413257da, 32'hc2a9c3fd, 32'h417409eb, 32'h42ab8002, 32'h41884ef2};
test_bias[1624:1624] = '{32'h41c53e2e};
test_output[1624:1624] = '{32'h46801ff8};
test_input[13000:13007] = '{32'hc05aa9e0, 32'hc26eb96a, 32'h41688655, 32'hc2741845, 32'h4294770a, 32'h4269c034, 32'hc111d199, 32'hc2be1138};
test_weights[13000:13007] = '{32'hc28befb8, 32'h416ac278, 32'h4268b37d, 32'h41c3c5bc, 32'h42018e34, 32'h4198e1d0, 32'hc28e961c, 32'h42271e4c};
test_bias[1625:1625] = '{32'hc181e715};
test_output[1625:1625] = '{32'hc4898cf0};
test_input[13008:13015] = '{32'hc2bfd026, 32'hc20a3800, 32'h424077b9, 32'hc1e81a2e, 32'hc2653b25, 32'h42b1de96, 32'hc2c45762, 32'hc270de03};
test_weights[13008:13015] = '{32'hc2425b94, 32'hc2ac277c, 32'hc1f1fee6, 32'hc1d705d1, 32'hc2ab9a8f, 32'h4282db99, 32'h4262d335, 32'h4218c0ff};
test_bias[1626:1626] = '{32'hc2bdd008};
test_output[1626:1626] = '{32'h46181554};
test_input[13016:13023] = '{32'hc202e9c6, 32'hc2c3bfa5, 32'h423adb47, 32'h423f1d39, 32'hc28d5984, 32'hc25aece5, 32'h414f985c, 32'h42add8e9};
test_weights[13016:13023] = '{32'hc2146447, 32'hc25e925f, 32'h42935a49, 32'h4253f098, 32'h42b11232, 32'hc23f5a52, 32'hc206a017, 32'h403648d0};
test_bias[1627:1627] = '{32'hc28732ad};
test_output[1627:1627] = '{32'h460886fd};
test_input[13024:13031] = '{32'hc291bcd0, 32'hc2868c7c, 32'hc2b7e8b8, 32'h427c56ee, 32'hc195383d, 32'h41ddd54c, 32'h42c52381, 32'h427721a1};
test_weights[13024:13031] = '{32'hc1f683b2, 32'h429c8c90, 32'h42b761f8, 32'h41dfe471, 32'hc293ba27, 32'hc2027de3, 32'h40fde829, 32'h421f7f5c};
test_bias[1628:1628] = '{32'hc253bc85};
test_output[1628:1628] = '{32'hc5bc242a};
test_input[13032:13039] = '{32'hc11a8cac, 32'h41346b1d, 32'hc22c42c6, 32'h42120474, 32'h42151729, 32'h42b63edd, 32'hc28073f3, 32'hc196689e};
test_weights[13032:13039] = '{32'h4155f7ae, 32'hc2807ffb, 32'hc1efc85f, 32'hc2944f23, 32'hc1d41642, 32'h4165228a, 32'hc1a2a702, 32'h42430920};
test_bias[1629:1629] = '{32'h40c871f5};
test_output[1629:1629] = '{32'hc4c2b497};
test_input[13040:13047] = '{32'h425f6819, 32'h421b7abb, 32'h4280422b, 32'hc2a83a9a, 32'h426558d3, 32'hc2618a9f, 32'h426141c1, 32'h41d95c99};
test_weights[13040:13047] = '{32'h4294d6d4, 32'hc21dc8cd, 32'h428e7534, 32'hc212757e, 32'h422364af, 32'hc295fee9, 32'h4284cda3, 32'hc23d1748};
test_bias[1630:1630] = '{32'hc127407a};
test_output[1630:1630] = '{32'h4696ac87};
test_input[13048:13055] = '{32'h42263706, 32'hc2bd4458, 32'h428c97b7, 32'hc226ec6e, 32'h4297aff1, 32'hc1efba84, 32'hc2b0c09f, 32'hc0a70017};
test_weights[13048:13055] = '{32'hc2535b73, 32'hc23a826a, 32'hc28d281b, 32'h429d320a, 32'hc1bbcccf, 32'h42580a80, 32'hc100c7a6, 32'h421d3202};
test_bias[1631:1631] = '{32'h42bc155b};
test_output[1631:1631] = '{32'hc609dc97};
test_input[13056:13063] = '{32'hc09f0a84, 32'h42beced0, 32'h42c74e2e, 32'h42624357, 32'h42295234, 32'h4186ea41, 32'hc06561ea, 32'hc29e0c68};
test_weights[13056:13063] = '{32'h41bf5e48, 32'h3fcb5ffc, 32'hc1fd4765, 32'hc0c80eaf, 32'hc29de212, 32'hc27d8397, 32'h426c5cca, 32'h40433dc0};
test_bias[1632:1632] = '{32'hc2aeab46};
test_output[1632:1632] = '{32'hc603aa57};
test_input[13064:13071] = '{32'hc1a5f255, 32'hc15d7c47, 32'hc1c7b991, 32'h414835d3, 32'hc1daf613, 32'hc2b9473b, 32'h42342c26, 32'hc25d9b54};
test_weights[13064:13071] = '{32'hc1418e42, 32'h41d461ad, 32'h417f3890, 32'hc120aeb6, 32'hc2aeffef, 32'hc0af567a, 32'hbfcb7438, 32'hc2a6b979};
test_bias[1633:1633] = '{32'h4203844e};
test_output[1633:1633] = '{32'h45d5cdbf};
test_input[13072:13079] = '{32'hc2c5cf95, 32'h42bdb474, 32'h41346ec3, 32'hc2a3c166, 32'h42ab6a84, 32'h42a00f0d, 32'h420365f2, 32'hc205100c};
test_weights[13072:13079] = '{32'h423cc2dc, 32'hc2b90471, 32'hc20b9b75, 32'hc28d03aa, 32'h41c21657, 32'hc28d2f2c, 32'hc24d36c6, 32'h42a7f65a};
test_bias[1634:1634] = '{32'h4288caee};
test_output[1634:1634] = '{32'hc67aad6c};
test_input[13080:13087] = '{32'hc193ef57, 32'h40c98b9b, 32'hc2507654, 32'h421b2ff9, 32'h424db7f7, 32'hc1f347de, 32'h41f48b7c, 32'hc2baa42a};
test_weights[13080:13087] = '{32'h3f78cb82, 32'h4294f328, 32'h4195532f, 32'h422f842e, 32'hc22e5f7d, 32'h42806412, 32'h426fbccb, 32'h4290e77d};
test_bias[1635:1635] = '{32'hc1511ead};
test_output[1635:1635] = '{32'hc5f89dfe};
test_input[13088:13095] = '{32'hc2992849, 32'hbe2beb45, 32'hc2ae3186, 32'hc24eaf91, 32'hc2a2184a, 32'h429bbfdf, 32'hc24001c5, 32'h4240e339};
test_weights[13088:13095] = '{32'hc284ee32, 32'h4252cb4b, 32'hc238da00, 32'h42835704, 32'h429481d1, 32'h40570a0d, 32'hbfe54ea7, 32'h41fb1777};
test_bias[1636:1636] = '{32'h42858d48};
test_output[1636:1636] = '{32'h44cad2b2};
test_input[13096:13103] = '{32'hc21de578, 32'hc201e645, 32'hc2c43063, 32'hc2a37377, 32'hc222c3f4, 32'hc2c58b94, 32'hc28dec70, 32'hc28a6e4f};
test_weights[13096:13103] = '{32'hc27383a2, 32'hc297d296, 32'hc2957abf, 32'h42bfce67, 32'h427c2250, 32'hc1845349, 32'hc288870b, 32'hc20946c2};
test_bias[1637:1637] = '{32'hc29c356b};
test_output[1637:1637] = '{32'h462531ba};
test_input[13104:13111] = '{32'hc23af738, 32'h429ddee9, 32'h416d9bfe, 32'h42a08709, 32'h42506924, 32'hc286b1e2, 32'hc2821ab4, 32'h42852954};
test_weights[13104:13111] = '{32'hc2700291, 32'h42a8dd5f, 32'h424c6c9b, 32'hc231e99d, 32'h3e9318c7, 32'h41b86076, 32'hc1f6dee2, 32'h42774166};
test_bias[1638:1638] = '{32'hc2a27203};
test_output[1638:1638] = '{32'h462e6b9e};
test_input[13112:13119] = '{32'hc16b7323, 32'h42a9f409, 32'hc238ffcc, 32'hc14b9a8c, 32'hc1c68683, 32'h4242d2e3, 32'hc279dc54, 32'h41a5c5be};
test_weights[13112:13119] = '{32'h425a6105, 32'hc186a04a, 32'h418f5579, 32'hc29fd469, 32'hc23a86d8, 32'hc28bd555, 32'h4157ea52, 32'hc067d835};
test_bias[1639:1639] = '{32'hc2b3e44d};
test_output[1639:1639] = '{32'hc5a5a9e2};
test_input[13120:13127] = '{32'hc1f1215c, 32'h429b8365, 32'h41a9bae0, 32'hc28a4be2, 32'h420a722e, 32'hc27f3963, 32'h42b37668, 32'hc210d481};
test_weights[13120:13127] = '{32'hc29f8bf0, 32'hc2276504, 32'h42ad2ab8, 32'h42091134, 32'hc1f780a2, 32'hc2be1d1f, 32'hc1a8a869, 32'h41324ddf};
test_bias[1640:1640] = '{32'hc257f8ae};
test_output[1640:1640] = '{32'h449de3e9};
test_input[13128:13135] = '{32'h41ee4d22, 32'h4235c9f3, 32'hc20996fc, 32'h3fc0b48e, 32'h42999838, 32'hc14e87d5, 32'h40d4c335, 32'h40ac57c2};
test_weights[13128:13135] = '{32'h41d01a13, 32'h427cef6c, 32'hc2bd1483, 32'hc1d7eeb1, 32'h4295b871, 32'h429d21dd, 32'h41cb2194, 32'hc29b56ba};
test_bias[1641:1641] = '{32'h42244d8b};
test_output[1641:1641] = '{32'h4631e9e5};
test_input[13136:13143] = '{32'hc239e716, 32'hbf420eb7, 32'hc27bea10, 32'h41f7995a, 32'hc2a2a106, 32'h42a91fb9, 32'h42a8d2a3, 32'h42246745};
test_weights[13136:13143] = '{32'hbcc187f9, 32'h42288f52, 32'hc2784c22, 32'hc2aca98a, 32'h40d00be9, 32'h415ce028, 32'hc24326fb, 32'h41337bab};
test_bias[1642:1642] = '{32'hc29d197b};
test_output[1642:1642] = '{32'hc4ec4ff9};
test_input[13144:13151] = '{32'h423625b6, 32'h42ae84e6, 32'h41cc6cc8, 32'h4095a9b6, 32'hc2a133cc, 32'h4225257c, 32'hc29a8d16, 32'hc2a64b13};
test_weights[13144:13151] = '{32'h423b8663, 32'hc275156c, 32'hc206d8e6, 32'hc28d3f35, 32'hc21cacc1, 32'hc29b23b6, 32'hc2555264, 32'hc17586d0};
test_bias[1643:1643] = '{32'hc2317091};
test_output[1643:1643] = '{32'h4461f051};
test_input[13152:13159] = '{32'hc27014b5, 32'h428744ab, 32'hc246bddf, 32'hc2aea33e, 32'hc218f7a4, 32'h42911e47, 32'h42684763, 32'hc291157f};
test_weights[13152:13159] = '{32'hc24fa59b, 32'hc2604dec, 32'hc215da23, 32'hc294c360, 32'hc254eb90, 32'hc24a06a3, 32'hc2771c84, 32'hc254b87b};
test_bias[1644:1644] = '{32'h42c0758b};
test_output[1644:1644] = '{32'h45c88715};
test_input[13160:13167] = '{32'hc1ecfe6d, 32'hc249f11c, 32'h429d9762, 32'h4297bb8e, 32'hc27e0bc6, 32'h426cb7de, 32'hc1f87742, 32'hc22b89e1};
test_weights[13160:13167] = '{32'hc270f6fd, 32'hc264775d, 32'h419a844b, 32'hc2a5ff01, 32'h41f9dbfa, 32'h4262bae7, 32'hc2c1b047, 32'hc1a92f15};
test_bias[1645:1645] = '{32'h42b203d8};
test_output[1645:1645] = '{32'h45a49f07};
test_input[13168:13175] = '{32'hc2c5d8d5, 32'hc2a14581, 32'hc27d577e, 32'hc27eef2c, 32'hc2a395b6, 32'h426d9435, 32'h4211f212, 32'h403ff434};
test_weights[13168:13175] = '{32'h41ed34be, 32'h41ea7b62, 32'h423beb35, 32'h42532a21, 32'hc1a558e4, 32'hc1ed702b, 32'hc264a170, 32'h413a748f};
test_bias[1646:1646] = '{32'h42b4f3a5};
test_output[1646:1646] = '{32'hc655940a};
test_input[13176:13183] = '{32'h42931462, 32'h428f7d6b, 32'h42af653d, 32'h41f013d9, 32'h411969fc, 32'hc28c2104, 32'hc1db7e8b, 32'h42937a83};
test_weights[13176:13183] = '{32'h41f85012, 32'h4287d24d, 32'h42a8fd6c, 32'hc0870bb0, 32'hc2ac9daf, 32'h422fbe17, 32'h4221114f, 32'h4104fedb};
test_bias[1647:1647] = '{32'hc0d1fb43};
test_output[1647:1647] = '{32'h461cc7bb};
test_input[13184:13191] = '{32'hc18a19c8, 32'hc29f27e5, 32'hc2bb4d40, 32'hc1cc71ec, 32'h412bf741, 32'hc1d4512b, 32'hc221919a, 32'hc1aae697};
test_weights[13184:13191] = '{32'h427a7408, 32'h42895cd2, 32'hc2be4c90, 32'h42c0fb0b, 32'hc26e3e72, 32'h42b768e0, 32'hc0476453, 32'h403ac306};
test_bias[1648:1648] = '{32'h41b823b1};
test_output[1648:1648] = '{32'hc5410dc8};
test_input[13192:13199] = '{32'hc0551d3d, 32'hc11d07c5, 32'h42afbcf5, 32'h40cea0ce, 32'hc2590956, 32'hc2ab09ad, 32'hc29b612d, 32'hc25f070b};
test_weights[13192:13199] = '{32'hc22aca54, 32'h41a74572, 32'hc0b7e2cd, 32'h412868b5, 32'h42b1b641, 32'hc299b98c, 32'hc11b1f10, 32'hc1ef0f49};
test_bias[1649:1649] = '{32'h422c054c};
test_output[1649:1649] = '{32'h456824f5};
test_input[13200:13207] = '{32'h42742400, 32'h413b0a3d, 32'hc257d8f0, 32'hc2ae0595, 32'h42750733, 32'h4296dbc7, 32'hc1e4ea01, 32'hc1aff64f};
test_weights[13200:13207] = '{32'h42aefe62, 32'h42239fdd, 32'h3f4fc825, 32'h428bc981, 32'h4278b3c4, 32'hc22931fc, 32'hc2b87954, 32'hc1d70448};
test_bias[1650:1650] = '{32'hc18c817e};
test_output[1650:1650] = '{32'h455c44b8};
test_input[13208:13215] = '{32'hc2bd2ba9, 32'h42c1a697, 32'h42766772, 32'h41ae91a0, 32'hc1cf2146, 32'h41ecfbd1, 32'hc2ad550c, 32'h40d34b87};
test_weights[13208:13215] = '{32'h422e4bde, 32'hc1ee7620, 32'h4295cd39, 32'h403ee2b0, 32'h429cfe6b, 32'hc231bdc2, 32'h42796b3c, 32'hc09c0552};
test_bias[1651:1651] = '{32'h42a0639a};
test_output[1651:1651] = '{32'hc62c6524};
test_input[13216:13223] = '{32'h41c73246, 32'h417c4da5, 32'h424ad91b, 32'hc23ba419, 32'h4180f553, 32'h42320001, 32'hc28884ae, 32'h4204e3a0};
test_weights[13216:13223] = '{32'hc2b52799, 32'h425ac5bd, 32'hc23042c9, 32'h425ad289, 32'hc26e7812, 32'hc294670d, 32'hc20e63cf, 32'h42ac1d3e};
test_bias[1652:1652] = '{32'h428dd032};
test_output[1652:1652] = '{32'hc59f47c6};
test_input[13224:13231] = '{32'h40a00d08, 32'hc2c09fbf, 32'hc25a2f09, 32'h4264f20b, 32'hc21b8420, 32'h41f267b1, 32'hc1a7ceb5, 32'hc16083f6};
test_weights[13224:13231] = '{32'hc23671bd, 32'h423ab64b, 32'h42a81a3a, 32'h4295e18b, 32'h42ac4209, 32'hc2993893, 32'hc1da0d53, 32'h428fe04f};
test_bias[1653:1653] = '{32'hc200a1f7};
test_output[1653:1653] = '{32'hc62e5bca};
test_input[13232:13239] = '{32'h429ad7e2, 32'hc134e4a4, 32'hc1d97fd1, 32'hc268d0d2, 32'hc2202055, 32'h42c1c5d7, 32'hc1ac6e84, 32'hc0910239};
test_weights[13232:13239] = '{32'hc2bbbd99, 32'hc1edfcd3, 32'h4291690a, 32'hc24b38d6, 32'h42a525ed, 32'h41a82e61, 32'h42b4e5a8, 32'h40d36d36};
test_bias[1654:1654] = '{32'h424668e5};
test_output[1654:1654] = '{32'hc60ef5e4};
test_input[13240:13247] = '{32'h42c74770, 32'h42b8d6fe, 32'h423ebade, 32'h4289ed49, 32'hc21c2054, 32'h427afbe4, 32'hc24fc375, 32'hc2937cf6};
test_weights[13240:13247] = '{32'hc26f66a6, 32'h426026ec, 32'hc2361811, 32'h41e1c905, 32'hc2102842, 32'hc2b45b75, 32'hc229c80c, 32'h41a3e6b4};
test_bias[1655:1655] = '{32'hc14ee161};
test_output[1655:1655] = '{32'hc58f1c3d};
test_input[13248:13255] = '{32'h4200ed8d, 32'hc2b42a3d, 32'hc2b846bd, 32'hc1734e15, 32'hc1d306d7, 32'h4292b57c, 32'h41d62063, 32'h42143114};
test_weights[13248:13255] = '{32'h425f3f15, 32'h42728f46, 32'h416a04e7, 32'hc2a812cd, 32'hc2acf52f, 32'hc11d8021, 32'h3e51b7f6, 32'h41cf84a8};
test_bias[1656:1656] = '{32'hc2b8051e};
test_output[1656:1656] = '{32'hc4a27a77};
test_input[13256:13263] = '{32'hc1bdf201, 32'hc1edbc7d, 32'h4253a244, 32'h42a6af07, 32'hc1fb03dc, 32'hc1e3020f, 32'hc28073f4, 32'hc17a4124};
test_weights[13256:13263] = '{32'hc2b8460a, 32'hc2629648, 32'hc29a6317, 32'h42a72405, 32'hc2a59b81, 32'hc1b284bd, 32'hc1a7a51f, 32'hc158d7d7};
test_bias[1657:1657] = '{32'hc205a2e8};
test_output[1657:1657] = '{32'h4633ce0b};
test_input[13264:13271] = '{32'hbe5715c8, 32'h419ff9f8, 32'h42aeca91, 32'hc2be86c0, 32'h42a5cb36, 32'hc21205e5, 32'h42b5f27a, 32'h427c736c};
test_weights[13264:13271] = '{32'h41b80f2a, 32'h42a86223, 32'hc24cd638, 32'hc095aae6, 32'hc295cc88, 32'hc202016b, 32'h423c0653, 32'hc29a0afc};
test_bias[1658:1658] = '{32'h420da09b};
test_output[1658:1658] = '{32'hc5f79739};
test_input[13272:13279] = '{32'hc1dbe870, 32'hc2c43110, 32'hc1a01c29, 32'h415dc183, 32'hc244f754, 32'h420c5d89, 32'hc28b1a3b, 32'h4294c28f};
test_weights[13272:13279] = '{32'h41df8d65, 32'h41253069, 32'h41a43579, 32'hc1e21d63, 32'hc15d0f08, 32'h41aa5f73, 32'hc1e1d040, 32'hc2ae21e0};
test_bias[1659:1659] = '{32'hc1978e91};
test_output[1659:1659] = '{32'hc5b1bc2f};
test_input[13280:13287] = '{32'h40c28c2c, 32'h42c0a5cc, 32'hc0573ff5, 32'h4278bb6c, 32'hc2a53644, 32'h427f21bb, 32'hc1f4e042, 32'h42ba2dfc};
test_weights[13280:13287] = '{32'h40c96f30, 32'h4229f048, 32'hc15a6147, 32'hc243cf26, 32'hc0326076, 32'h417444ad, 32'h41c5dcfd, 32'h412438fb};
test_bias[1660:1660] = '{32'hc1f0ac88};
test_output[1660:1660] = '{32'h451c8c4f};
test_input[13288:13295] = '{32'h4278405c, 32'hc22d8717, 32'h428ad07a, 32'hc2408b75, 32'h422e2fd6, 32'h41d5f98a, 32'h42a07b69, 32'h42163a42};
test_weights[13288:13295] = '{32'hc25ba65c, 32'h425210d9, 32'h41a4440f, 32'hc282dfb3, 32'h429dd131, 32'h41851ece, 32'hc25b1a1a, 32'h42927775};
test_bias[1661:1661] = '{32'h42bfe41f};
test_output[1661:1661] = '{32'h4498a4ad};
test_input[13296:13303] = '{32'h4204b8e9, 32'h41d7c895, 32'h42304eda, 32'h41870f7f, 32'h419a3867, 32'h40b3a7f5, 32'h4155b79b, 32'h40f0bcb0};
test_weights[13296:13303] = '{32'hc15b4b05, 32'h429a5a9b, 32'hc2892d06, 32'h424cc78a, 32'h42ae1c23, 32'hc109649f, 32'h42be2b89, 32'hc1fb682b};
test_bias[1662:1662] = '{32'h42c7b9ec};
test_output[1662:1662] = '{32'h450b7986};
test_input[13304:13311] = '{32'h42960010, 32'hc27e0d96, 32'hc232635c, 32'hc2a31a89, 32'hc2a17b8a, 32'h425421d6, 32'h41c8e855, 32'h4284da85};
test_weights[13304:13311] = '{32'h40f1754b, 32'h42564898, 32'h41ead48a, 32'h42a1391a, 32'h42851a19, 32'h424275d5, 32'hc2b17983, 32'h416ac7ee};
test_bias[1663:1663] = '{32'hc1c7808a};
test_output[1663:1663] = '{32'hc6672640};
test_input[13312:13319] = '{32'hc23b0a65, 32'h41e18abc, 32'h429ac39c, 32'hc2b96acc, 32'h41fb7f8c, 32'h42a7478f, 32'h40827d19, 32'h4177d6ac};
test_weights[13312:13319] = '{32'hc2ad9a7e, 32'hc29de90f, 32'h42bb78b5, 32'h42a716ca, 32'hc2255332, 32'hc1b13d54, 32'hc244c250, 32'h42a77104};
test_bias[1664:1664] = '{32'hc21ceaa5};
test_output[1664:1664] = '{32'hc43c92c6};
test_input[13320:13327] = '{32'h401e4089, 32'hc2ba408e, 32'h419e147c, 32'hc2881b0a, 32'hc1f41bc3, 32'hc25e16dc, 32'hc1ab2828, 32'hc240920e};
test_weights[13320:13327] = '{32'hc16dc1ac, 32'hc2298f29, 32'hc1ae9977, 32'h4284ceb3, 32'hc187b008, 32'h422e1b3c, 32'h42044873, 32'hc2974f46};
test_bias[1665:1665] = '{32'hc178ab99};
test_output[1665:1665] = '{32'hc19b0c0c};
test_input[13328:13335] = '{32'hc0089ce2, 32'hc241358e, 32'h42936f17, 32'hc22d52e0, 32'hc2912ee1, 32'hc2b13ce8, 32'hc21a166d, 32'hc1cd5eaa};
test_weights[13328:13335] = '{32'h4234ab6b, 32'hc220a3dd, 32'hc145be2a, 32'hc1fdb10e, 32'hc0c6c7fd, 32'hc2a27f27, 32'hc0324aeb, 32'h429ed2d9};
test_bias[1666:1666] = '{32'h42682e62};
test_output[1666:1666] = '{32'h45fca22a};
test_input[13336:13343] = '{32'h42c200e7, 32'hbe81e9da, 32'hc1741254, 32'h40d0e8aa, 32'hc28f8b1d, 32'hc15c0822, 32'h40fbe80c, 32'h42c5b5cc};
test_weights[13336:13343] = '{32'h42077ee6, 32'hc15f055d, 32'h422ac28b, 32'h429532d6, 32'hc1c32aa2, 32'h41b8d28d, 32'h42b7b999, 32'h416ae836};
test_bias[1667:1667] = '{32'hc174429d};
test_output[1667:1667] = '{32'h45d1ed0a};
test_input[13344:13351] = '{32'h42a395c1, 32'h4242ff73, 32'h429c10d6, 32'hc2359690, 32'h42be1209, 32'hc294e1c1, 32'h41883e59, 32'hc229f2dd};
test_weights[13344:13351] = '{32'hc1e9d4de, 32'hc1e91c49, 32'h4203dcdb, 32'hc2af7738, 32'hbea8d19e, 32'hc2100a2d, 32'hc21cd2c2, 32'hc2ae37e6};
test_bias[1668:1668] = '{32'h42b17e9f};
test_output[1668:1668] = '{32'h46050d75};
test_input[13352:13359] = '{32'hc2890fae, 32'hc21973e4, 32'hc2c33a52, 32'h428885b9, 32'hc220faff, 32'h42201b40, 32'hc263c597, 32'hc06481e2};
test_weights[13352:13359] = '{32'hc21343f0, 32'h42c7e081, 32'hc287c433, 32'h420e0d79, 32'hc29103c2, 32'h429f7329, 32'h429a4ba9, 32'hc1a6f2e8};
test_bias[1669:1669] = '{32'h420b33dc};
test_output[1669:1669] = '{32'h4615744f};
test_input[13360:13367] = '{32'h42957adf, 32'hc21a1f7b, 32'h41d8f10b, 32'hc2b852e3, 32'hc2c680e0, 32'h414e2e12, 32'hc0f7ebfc, 32'hc195e282};
test_weights[13360:13367] = '{32'hc18fd380, 32'hc1e647cc, 32'hc2870256, 32'h42bb6fbe, 32'hc1e2ad83, 32'hc273f5db, 32'hc1539457, 32'hc2b7790d};
test_bias[1670:1670] = '{32'hc2618fcc};
test_output[1670:1670] = '{32'hc5d7fa2b};
test_input[13368:13375] = '{32'hc282a9c3, 32'hc24e06b8, 32'h4230a2f3, 32'h42c157dc, 32'h4293e270, 32'hc1dfa7e1, 32'h42914888, 32'h41024c36};
test_weights[13368:13375] = '{32'h420f1b24, 32'h41126e0d, 32'hc29aecbe, 32'hc2a29537, 32'hc2265af8, 32'hc22c7cac, 32'hc11685fb, 32'h42995115};
test_bias[1671:1671] = '{32'h4292dff5};
test_output[1671:1671] = '{32'hc6791d09};
test_input[13376:13383] = '{32'h4201a02c, 32'h42384ec3, 32'h429d52ba, 32'h429f4e34, 32'hc22b5400, 32'h41db3556, 32'hc29ecfab, 32'h429a2296};
test_weights[13376:13383] = '{32'hc260bc63, 32'h42ae39b1, 32'hc18d6a62, 32'hc2b07e1e, 32'h42abd824, 32'hc1c9c841, 32'h4232fdbe, 32'h40999e26};
test_bias[1672:1672] = '{32'hc237cc8b};
test_output[1672:1672] = '{32'hc6580bd1};
test_input[13384:13391] = '{32'h4173d3b2, 32'h4247680a, 32'hc2c3d49c, 32'hc24809ac, 32'h40bf9f17, 32'h3edb6a56, 32'h42370e2b, 32'h423d19f4};
test_weights[13384:13391] = '{32'h419c4ae3, 32'hc29a45d9, 32'hc29d7f93, 32'h42bb203f, 32'h4286a965, 32'h4207c667, 32'hc2b124bf, 32'h4258e6d4};
test_bias[1673:1673] = '{32'hc2675365};
test_output[1673:1673] = '{32'hc4cdbcb0};
test_input[13392:13399] = '{32'h407639df, 32'h42b83c92, 32'hbfa0287e, 32'h4297f068, 32'hc1f33cfd, 32'hc2c64f7b, 32'h40a6a442, 32'h410d3a62};
test_weights[13392:13399] = '{32'hc1fc8ed3, 32'hc208a30c, 32'h42b88e94, 32'hc2a26c36, 32'h410a8144, 32'h40cbec7e, 32'hc235c52c, 32'h429fbcc1};
test_bias[1674:1674] = '{32'h4285d28e};
test_output[1674:1674] = '{32'hc61ae41f};
test_input[13400:13407] = '{32'hc11c67f3, 32'h41923c94, 32'h4297e1bf, 32'h3e0b754c, 32'hc20db897, 32'hc2c6522e, 32'hc2c690e0, 32'hc2a9d3b8};
test_weights[13400:13407] = '{32'hc2999e07, 32'h42846522, 32'hc1914b1c, 32'h42b4a7d7, 32'hc251c565, 32'h42b14624, 32'h42592232, 32'h42944d05};
test_bias[1675:1675] = '{32'hc288091a};
test_output[1675:1675] = '{32'hc68d561b};
test_input[13408:13415] = '{32'h42b9b0d7, 32'hc2a3283e, 32'h42a4a1b3, 32'h41b7f998, 32'h4208a0bc, 32'hc2c65f23, 32'hc26cb625, 32'h41920e7a};
test_weights[13408:13415] = '{32'h3e997b82, 32'h421fc9b3, 32'hc2ab8238, 32'h42a2feb7, 32'hc124b523, 32'h3ffd34a7, 32'hc1d2499c, 32'h4291ab91};
test_bias[1676:1676] = '{32'hc26f6f1e};
test_output[1676:1676] = '{32'hc5bfd0f4};
test_input[13416:13423] = '{32'h416681a0, 32'h422b9389, 32'h42c0b743, 32'h42a7ce92, 32'h42b278f5, 32'hc2a88686, 32'hc2c50aa9, 32'hc2891a26};
test_weights[13416:13423] = '{32'h40596cb7, 32'h424222ef, 32'hc2bae6b0, 32'h417dc58b, 32'h42b54935, 32'h42123f41, 32'hc29987d8, 32'hc1a6166e};
test_bias[1677:1677] = '{32'h40ef688e};
test_output[1677:1677] = '{32'h46042951};
test_input[13424:13431] = '{32'h416fe04b, 32'hbfc03a63, 32'h4201009b, 32'h42525761, 32'h41e5a0cd, 32'hc124a465, 32'h42834192, 32'h42a4a2c1};
test_weights[13424:13431] = '{32'h42aab2be, 32'h42a088e4, 32'h41fba78f, 32'hc19a14b8, 32'hc2301487, 32'h4234160f, 32'h429185bd, 32'h424825ea};
test_bias[1678:1678] = '{32'h425d354b};
test_output[1678:1678] = '{32'h4602fd63};
test_input[13432:13439] = '{32'h41a7a8ae, 32'hc298017b, 32'h421512cf, 32'h4220816e, 32'hc1974d0c, 32'hc03d6b94, 32'hc245bccf, 32'hc1dfbe61};
test_weights[13432:13439] = '{32'hc24adebd, 32'h42833a2f, 32'hc2676c53, 32'h4275054c, 32'h41544819, 32'h42a3c62b, 32'hc28ff09e, 32'h40809e14};
test_bias[1679:1679] = '{32'hc28f99b7};
test_output[1679:1679] = '{32'hc5333ae0};
test_input[13440:13447] = '{32'hc25cd6f4, 32'h425a9316, 32'h42b9fe04, 32'hc24a0737, 32'h4291d660, 32'h42863068, 32'h4223e6cf, 32'h428176b6};
test_weights[13440:13447] = '{32'h41c8c301, 32'hc2a3b008, 32'hc2c509be, 32'h41fc110a, 32'hc1d63123, 32'h42159f2a, 32'h42161958, 32'hc28596d6};
test_bias[1680:1680] = '{32'h420825be};
test_output[1680:1680] = '{32'hc692eb87};
test_input[13448:13455] = '{32'h429a9221, 32'hc211e193, 32'h420177a7, 32'h428259e2, 32'hc29ce82c, 32'hc26c06d4, 32'h42c7a92d, 32'hc0d319e2};
test_weights[13448:13455] = '{32'hc2bc5c8b, 32'h4293eccd, 32'h4250c49b, 32'h429260a2, 32'h4282dbd3, 32'hc2b8e61a, 32'h42123045, 32'hbef684e1};
test_bias[1681:1681] = '{32'hc2a06b9b};
test_output[1681:1681] = '{32'h43bc50c9};
test_input[13456:13463] = '{32'h42bc383e, 32'h42a36222, 32'h416a1aae, 32'h4228406d, 32'hc2332a1a, 32'h42b08e67, 32'h4134c400, 32'h4143f75d};
test_weights[13456:13463] = '{32'hc2b5d636, 32'hc230731f, 32'hc1853cd4, 32'hc249f0e5, 32'hc04d19e8, 32'hc215d7e4, 32'h42b97589, 32'h41937309};
test_bias[1682:1682] = '{32'hc2c66da0};
test_output[1682:1682] = '{32'hc68108db};
test_input[13464:13471] = '{32'h42a66f1b, 32'hbfec8f95, 32'h41aa5aed, 32'h42639376, 32'hc2954ee2, 32'hc2b4f772, 32'hc10f43ee, 32'hc2827135};
test_weights[13464:13471] = '{32'hc28afb72, 32'hc28528f1, 32'h4214c3b4, 32'hc25fb7da, 32'h42924a48, 32'h41cfea51, 32'hc275c0f7, 32'h41c1e01c};
test_bias[1683:1683] = '{32'hc290f67e};
test_output[1683:1683] = '{32'hc6848a0c};
test_input[13472:13479] = '{32'h42a9c54e, 32'h4003ccd7, 32'h42908b21, 32'hc27af739, 32'hc27e9c35, 32'hc27672f1, 32'hc206086e, 32'hc23ff3fb};
test_weights[13472:13479] = '{32'h417d3abe, 32'hc21fc55d, 32'h41de20b1, 32'h427cf75e, 32'hc241987f, 32'h42bf3bb9, 32'h420171ad, 32'h4269d3b0};
test_bias[1684:1684] = '{32'h4282dc57};
test_output[1684:1684] = '{32'hc5e53490};
test_input[13480:13487] = '{32'h4298e531, 32'hbf62484d, 32'hc194ff8d, 32'hc28f0a33, 32'hc222d0f6, 32'h402eae0b, 32'h42994da1, 32'h41a281d2};
test_weights[13480:13487] = '{32'hc2c4efc7, 32'h4071b72d, 32'h420d8fab, 32'hc25a2386, 32'hc11b3235, 32'hc2a9566e, 32'h40d04431, 32'hc0f095cb};
test_bias[1685:1685] = '{32'hc2c254d0};
test_output[1685:1685] = '{32'hc57251d8};
test_input[13488:13495] = '{32'hc0ea84be, 32'hc2c57617, 32'h41aef36c, 32'hc112f172, 32'h420f7060, 32'hc24eaf4b, 32'hc2b04ff8, 32'hc29d32f2};
test_weights[13488:13495] = '{32'h414aaaa3, 32'hc2c088c4, 32'hc12118d8, 32'h429741a9, 32'h421b9d18, 32'h42b1f7eb, 32'hc1214630, 32'h41116249};
test_bias[1686:1686] = '{32'hc19dfb26};
test_output[1686:1686] = '{32'h45aa45bf};
test_input[13496:13503] = '{32'h421131c9, 32'h41a0fb67, 32'hc224baaf, 32'hc23790d5, 32'h4266c161, 32'h426d9b9b, 32'h42905350, 32'h42809a2c};
test_weights[13496:13503] = '{32'hc2b1873c, 32'h428ec9a4, 32'h42423746, 32'hc29e8e20, 32'h4184ced0, 32'hc2bfd4a0, 32'hc20039f6, 32'hc1b12d48};
test_bias[1687:1687] = '{32'hc2c62bdf};
test_output[1687:1687] = '{32'hc6084c69};
test_input[13504:13511] = '{32'h4234dc07, 32'h4017f1a8, 32'h4010df00, 32'h4225fb12, 32'hc2837171, 32'h4281527c, 32'hbf991242, 32'hc255ada6};
test_weights[13504:13511] = '{32'hc2c12b31, 32'hc114fe8d, 32'hc18ed919, 32'h4207b179, 32'h42007588, 32'h41e6d242, 32'h426fea83, 32'h42a936e3};
test_bias[1688:1688] = '{32'hc2c126f8};
test_output[1688:1688] = '{32'hc5f89729};
test_input[13512:13519] = '{32'h419b2fa2, 32'h422a8f27, 32'h40fa683a, 32'h41b79c8a, 32'hc2c73fa8, 32'h421a9d3d, 32'hc2039725, 32'hc15c6620};
test_weights[13512:13519] = '{32'h4238bef0, 32'h41a9629b, 32'hc238a48c, 32'hc29fdbff, 32'h4109273a, 32'h41cea23d, 32'h426284b9, 32'hc20b46d8};
test_bias[1689:1689] = '{32'h41c830cc};
test_output[1689:1689] = '{32'hc4c95c3a};
test_input[13520:13527] = '{32'hc256cb32, 32'hc2c0c3bc, 32'hc282ab7e, 32'h42a767d9, 32'h4218933b, 32'h4270de18, 32'h428b62c7, 32'h41ac9a0f};
test_weights[13520:13527] = '{32'hc1f7f410, 32'h422fd2fc, 32'h42af2e66, 32'hc2b50cf3, 32'hc2342a41, 32'h424760e0, 32'hc275b282, 32'h41c1a08e};
test_bias[1690:1690] = '{32'h42948d68};
test_output[1690:1690] = '{32'hc68ec240};
test_input[13528:13535] = '{32'h423ecedc, 32'h42558d56, 32'h429f5ba9, 32'h4253557c, 32'hc2ab9f0d, 32'hc0c418f7, 32'h41a2f0e9, 32'hc287633c};
test_weights[13528:13535] = '{32'hc297fd2d, 32'h414b5e35, 32'h42ba8972, 32'h42949b9b, 32'h4246dfeb, 32'h42b0e677, 32'hc283163a, 32'hbfa9569e};
test_bias[1691:1691] = '{32'hc285c8b1};
test_output[1691:1691] = '{32'h450f20de};
test_input[13536:13543] = '{32'hc2686660, 32'h42993d78, 32'hc2a468a2, 32'hc25325ed, 32'h41a3b721, 32'hc250d5f1, 32'hc27998ac, 32'h4295c15a};
test_weights[13536:13543] = '{32'hc2b3e7b8, 32'hc25a9cf7, 32'hc2be1a85, 32'h42908eeb, 32'h4205b508, 32'h423b671e, 32'h413da924, 32'h4282d1ef};
test_bias[1692:1692] = '{32'hc25666ed};
test_output[1692:1692] = '{32'h45e69bf0};
test_input[13544:13551] = '{32'hc2c4d0b8, 32'h42603ed1, 32'h42419645, 32'hc1aaf13a, 32'hc225b370, 32'hbf883ec6, 32'h4258681a, 32'h40571f50};
test_weights[13544:13551] = '{32'hc2967581, 32'h41f86b7b, 32'hc2b5ee18, 32'h403a1e1c, 32'h424fb66c, 32'h428f63f5, 32'h4280baab, 32'h42441cea};
test_bias[1693:1693] = '{32'h41c5a1cf};
test_output[1693:1693] = '{32'h45bf5de2};
test_input[13552:13559] = '{32'hc241d71f, 32'h4292b9f5, 32'h42900517, 32'h42bc8eed, 32'h41fbb73c, 32'hc281a8cb, 32'h42be920d, 32'h3f49dbec};
test_weights[13552:13559] = '{32'hc0d47762, 32'hc19bd81b, 32'hc28d86ea, 32'h42439b1f, 32'h422e0725, 32'hc183d4cd, 32'hc2142e4f, 32'h4252983c};
test_bias[1694:1694] = '{32'hc1d31b67};
test_output[1694:1694] = '{32'hc526e2d1};
test_input[13560:13567] = '{32'h41dc73bf, 32'h42170843, 32'hc2462f50, 32'hc1ec2615, 32'hc19b72d3, 32'hc2553643, 32'h420d2fc2, 32'hc2c1ed5f};
test_weights[13560:13567] = '{32'hc1ecf81d, 32'h41d1e24f, 32'h42514a02, 32'hc24c42ec, 32'hc29e0318, 32'h41d264f0, 32'h42a6cbc4, 32'hc2a5fcd4};
test_bias[1695:1695] = '{32'h42ba8ba0};
test_output[1695:1695] = '{32'h46210c10};
test_input[13568:13575] = '{32'hc221777f, 32'h4212e2ea, 32'hc0c06b55, 32'hc106965e, 32'h42bad19c, 32'h40f34869, 32'hc14d58b8, 32'h42710e43};
test_weights[13568:13575] = '{32'hc225fa26, 32'hc22280d7, 32'hc2b02ddf, 32'h42c673b3, 32'hc287b6c1, 32'h42582c30, 32'hc21ebc09, 32'hc2b472f8};
test_bias[1696:1696] = '{32'h4198faa9};
test_output[1696:1696] = '{32'hc62b392a};
test_input[13576:13583] = '{32'h412458cf, 32'h42418e1d, 32'h4193176a, 32'h42945944, 32'hc1c7b371, 32'h41afda4a, 32'hc2531b24, 32'h4245a004};
test_weights[13576:13583] = '{32'hc12a7274, 32'hc22ea4f4, 32'h42a6d5d0, 32'hc26c233c, 32'h42c44a20, 32'hc1865746, 32'hc1fda3aa, 32'hc2c73833};
test_bias[1697:1697] = '{32'h428ae0e1};
test_output[1697:1697] = '{32'hc62ce3b7};
test_input[13584:13591] = '{32'hc2be060c, 32'h42122d96, 32'h40caf20f, 32'hc2ba5054, 32'h42b42c65, 32'h42507528, 32'hc0e08799, 32'hc21316e1};
test_weights[13584:13591] = '{32'h42b57438, 32'hc0cc44bd, 32'hc233f621, 32'hc27330a8, 32'hc121d929, 32'hc2b3569b, 32'h41df29bc, 32'hc1fee04d};
test_bias[1698:1698] = '{32'hc1f8fb7b};
test_output[1698:1698] = '{32'hc5fd955a};
test_input[13592:13599] = '{32'h42a717ef, 32'hc2535262, 32'h4251f5d3, 32'hc2805120, 32'hc2ae4190, 32'h416f99fd, 32'h42a5c1db, 32'hbf4c5713};
test_weights[13592:13599] = '{32'hc298e6e4, 32'h423113a6, 32'h42845115, 32'h41ca3900, 32'hc2011dc9, 32'h42b08d98, 32'h418c51e2, 32'h41c90fb0};
test_bias[1699:1699] = '{32'h423b9b02};
test_output[1699:1699] = '{32'hc49d873d};
test_input[13600:13607] = '{32'hc229725d, 32'hc299b645, 32'h41674e85, 32'h41c8667a, 32'h42398524, 32'hc2a253ee, 32'hc2b0d1b9, 32'hc2857175};
test_weights[13600:13607] = '{32'h422f702f, 32'h428538f3, 32'h3f9021e9, 32'h42913162, 32'h428b5544, 32'h42373847, 32'h4294b459, 32'hc2a558b4};
test_bias[1700:1700] = '{32'hc2b70778};
test_output[1700:1700] = '{32'hc5d3d084};
test_input[13608:13615] = '{32'h41fc9fc1, 32'hc1036422, 32'h42bad711, 32'h42be158f, 32'hc2a77696, 32'hc1b7b768, 32'hc281fb5d, 32'hc2b6fc1f};
test_weights[13608:13615] = '{32'h42c438eb, 32'hc22990e8, 32'hc1994b12, 32'hc2c598f9, 32'h42930a35, 32'h42b7adb8, 32'hc2c5cad7, 32'hc2a9cb63};
test_bias[1701:1701] = '{32'hc251138c};
test_output[1701:1701] = '{32'hc4e809c5};
test_input[13616:13623] = '{32'hc2754cd1, 32'hc1e0488a, 32'hc2a79f6d, 32'hc235c1bc, 32'h42982f08, 32'hc2b54844, 32'h41dc498a, 32'h42160b37};
test_weights[13616:13623] = '{32'h4209791f, 32'hc201c2a3, 32'hc29abc09, 32'hc13acdfb, 32'hc2be9cd2, 32'hbf49853a, 32'hc2385fb6, 32'h42068989};
test_bias[1702:1702] = '{32'hc29b4fb5};
test_output[1702:1702] = '{32'hc4b52996};
test_input[13624:13631] = '{32'hc0e6e4ab, 32'hc29b58f8, 32'h42b1176e, 32'h42267f42, 32'hc2ae9fee, 32'h41dafe3d, 32'hc2a87877, 32'hc2c625be};
test_weights[13624:13631] = '{32'hc27bddc8, 32'h41a95849, 32'hc2a0b35c, 32'h42abef0e, 32'hc20df341, 32'h4240600b, 32'h4270f2b1, 32'hc29336a9};
test_bias[1703:1703] = '{32'h40efad1e};
test_output[1703:1703] = '{32'h44ef55f8};
test_input[13632:13639] = '{32'h411b224e, 32'h42c598bc, 32'hc2ae04b9, 32'hbf5b4a84, 32'h42450063, 32'h42a6fd76, 32'hc2abd4b2, 32'h41b16905};
test_weights[13632:13639] = '{32'h42be637f, 32'h429de07e, 32'h418c875a, 32'hc2b5a887, 32'h411382c2, 32'h4283bde2, 32'hc2b6a1a6, 32'hc1c379e4};
test_bias[1704:1704] = '{32'hc29717ff};
test_output[1704:1704] = '{32'h469fcaad};
test_input[13640:13647] = '{32'hc288bf8d, 32'h426daea2, 32'hc208df3f, 32'hc24d3d5e, 32'hc29a5186, 32'h40134787, 32'hc02eba2e, 32'h4116068d};
test_weights[13640:13647] = '{32'hc2830ea0, 32'h3f2eacb0, 32'hc25bbc2a, 32'h42a6343f, 32'hc23a498d, 32'h41a701cd, 32'hc28e29d8, 32'hc29fba51};
test_bias[1705:1705] = '{32'h4288d0fe};
test_output[1705:1705] = '{32'h45a55ef7};
test_input[13648:13655] = '{32'hc1ec15be, 32'h419c310a, 32'h42c44760, 32'h41a0e1e3, 32'h428ec237, 32'h41dbbb7d, 32'h4220e46f, 32'h42b95038};
test_weights[13648:13655] = '{32'h4130b9c8, 32'h421aa42e, 32'hc1e02969, 32'h426c76f8, 32'hc170d036, 32'h42b2ab9b, 32'h42759233, 32'hc2b3cdb8};
test_bias[1706:1706] = '{32'hc2c31a25};
test_output[1706:1706] = '{32'hc5b27777};
test_input[13656:13663] = '{32'h42531fa1, 32'h4265fe84, 32'h428cf5dd, 32'h42be09cb, 32'hc284431f, 32'hc2aea7aa, 32'h41a07ecd, 32'h42301fb0};
test_weights[13656:13663] = '{32'hc2a34448, 32'hc09ddda6, 32'h42866ed8, 32'hc214ce78, 32'h416b7072, 32'hc1cd3753, 32'hc2846739, 32'h428993e6};
test_bias[1707:1707] = '{32'hc278d2a9};
test_output[1707:1707] = '{32'hc3f22198};
test_input[13664:13671] = '{32'h42509da7, 32'hc28d3d22, 32'h42c7cae9, 32'hc253a493, 32'h42a46254, 32'h41b296ba, 32'h428006ec, 32'h42736cf1};
test_weights[13664:13671] = '{32'hc2a7c1b4, 32'h42b0ae0f, 32'hc28c024c, 32'h41c8c91f, 32'hc26e7e39, 32'h42373534, 32'hc007d146, 32'hc204e57e};
test_bias[1708:1708] = '{32'hc2152d40};
test_output[1708:1708] = '{32'hc6c35ec7};
test_input[13672:13679] = '{32'h42129912, 32'hc2aa6444, 32'hc2102c4f, 32'hc0eeda8b, 32'hc26a2b2e, 32'h4125436f, 32'hc29e896a, 32'hc24bb967};
test_weights[13672:13679] = '{32'h428fae04, 32'hc226a2cf, 32'hc2855507, 32'h42b66f2b, 32'hc0fae72d, 32'hc29d3366, 32'h42243ec0, 32'h42c3d8e4};
test_bias[1709:1709] = '{32'hc22687e1};
test_output[1709:1709] = '{32'hc4372812};
test_input[13680:13687] = '{32'hc2217f7f, 32'h4270353f, 32'hc136c353, 32'hc232d766, 32'h41827353, 32'hc18c8ca7, 32'hc1b32f91, 32'h428e4256};
test_weights[13680:13687] = '{32'hc2c44457, 32'hc24da8d0, 32'hc29a70ef, 32'h4205b6b9, 32'h425aa8c0, 32'hc18c528e, 32'h42a46688, 32'hc1ff1e7b};
test_bias[1710:1710] = '{32'hc2312508};
test_output[1710:1710] = '{32'hc5284340};
test_input[13688:13695] = '{32'hc20ee20d, 32'hc2bbb2d8, 32'hc26948b2, 32'h429b7ee4, 32'hc28adbbd, 32'hc2af1f93, 32'h422d37d0, 32'h42259efd};
test_weights[13688:13695] = '{32'hc12b8496, 32'hc0bbcf5d, 32'hc08d4aa9, 32'hc2a8ab8a, 32'hc18beac8, 32'hc1d15d6b, 32'hc1cdbd2d, 32'hc09dfa7a};
test_bias[1711:1711] = '{32'h42accaa6};
test_output[1711:1711] = '{32'hc54137cc};
test_input[13696:13703] = '{32'h4295273a, 32'hc24f29a2, 32'h42019ff4, 32'hc0f4220d, 32'h424ded56, 32'h42b7abe5, 32'h42c4c5b1, 32'h424cd386};
test_weights[13696:13703] = '{32'hc12ee88c, 32'hc251b0b2, 32'h41defbf1, 32'h41ec7936, 32'h42a2adb0, 32'h42bfd185, 32'hc29e8552, 32'h42a1f88e};
test_bias[1712:1712] = '{32'hc2ad9936};
test_output[1712:1712] = '{32'h4638ebc1};
test_input[13704:13711] = '{32'h40ac420a, 32'h419da0aa, 32'hc12f6c8b, 32'hc145ccf7, 32'h4295285c, 32'hc2c56407, 32'hc14018dd, 32'h42b2606f};
test_weights[13704:13711] = '{32'h4270338d, 32'hc27cfc73, 32'hc1a28f1d, 32'hc1bcc2b9, 32'hc21902f7, 32'h412986bc, 32'hc299863d, 32'h42c6a33f};
test_bias[1713:1713] = '{32'h414a58ad};
test_output[1713:1713] = '{32'h45ab6aa6};
test_input[13712:13719] = '{32'hc2c2bcdc, 32'hc17a7dc1, 32'hc26eb8a4, 32'h41fffa37, 32'hc2841f71, 32'h42883051, 32'h42157e50, 32'h426f5b2f};
test_weights[13712:13719] = '{32'h3fdf950a, 32'hc2645650, 32'hc2be1e75, 32'h41d46cb1, 32'hc2a2afd8, 32'hc2432e84, 32'h41dd3aaf, 32'h419c45ee};
test_bias[1714:1714] = '{32'hc2933f48};
test_output[1714:1714] = '{32'h463288b9};
test_input[13720:13727] = '{32'hc2a18cf0, 32'hc25c9264, 32'hc2c20637, 32'hc2b9e51f, 32'hc281c7f9, 32'h422f1ca7, 32'hc154cf8b, 32'h41a99327};
test_weights[13720:13727] = '{32'hc29c997f, 32'hc18c6205, 32'h40d44875, 32'h420ffc37, 32'hc201cbc5, 32'hc24b836a, 32'h42651471, 32'hc086d1d4};
test_bias[1715:1715] = '{32'hc2c7a10b};
test_output[1715:1715] = '{32'h450b66ec};
test_input[13728:13735] = '{32'h42c4cef9, 32'h424891fa, 32'hc29f270a, 32'h4280274f, 32'h417594a5, 32'h42bf2055, 32'hc120815b, 32'h41e0a616};
test_weights[13728:13735] = '{32'hc291d79e, 32'hc2077870, 32'h4271648a, 32'hc298774f, 32'hc2abd141, 32'h4228547b, 32'hc232067d, 32'hbf1879f7};
test_bias[1716:1716] = '{32'h4205ab0f};
test_output[1716:1716] = '{32'hc6708b9d};
test_input[13736:13743] = '{32'h4203dd14, 32'hc2b88db7, 32'h429b7fe7, 32'hc1353f46, 32'h42ae8cfe, 32'hc16cd9d8, 32'hc1c75624, 32'h406b0b1c};
test_weights[13736:13743] = '{32'h41b0cac3, 32'h417f528b, 32'h425dfb65, 32'h4206da31, 32'h420bcada, 32'h421d6c12, 32'h42640f56, 32'hc2a21cee};
test_bias[1717:1717] = '{32'h422b981a};
test_output[1717:1717] = '{32'h4578cf26};
test_input[13744:13751] = '{32'hc1d74559, 32'h421bfb70, 32'h42816d2e, 32'h4112a522, 32'h4092a5cb, 32'h412798b2, 32'hc1969d40, 32'h42816621};
test_weights[13744:13751] = '{32'h4227ac35, 32'h41522ad8, 32'hc2c3430a, 32'h42c53c26, 32'h40a9a5a2, 32'h418c4f47, 32'hc2c4239e, 32'hc1a5c231};
test_bias[1718:1718] = '{32'h4213163f};
test_output[1718:1718] = '{32'hc5a4fac4};
test_input[13752:13759] = '{32'h41bf25df, 32'hc2b26436, 32'hc2a1070c, 32'h424b9a2b, 32'hc2b135ed, 32'h4267bc70, 32'hc1e0b4c6, 32'h41ce6e3e};
test_weights[13752:13759] = '{32'hc2ad1a5e, 32'hc2b63ec4, 32'hbf9bbfee, 32'h422af1c3, 32'hc2c3d229, 32'h4214324f, 32'h4275cded, 32'h42516207};
test_bias[1719:1719] = '{32'h4067318f};
test_output[1719:1719] = '{32'h4692be1e};
test_input[13760:13767] = '{32'hc13511b3, 32'h4261ee75, 32'hc1bc0d5b, 32'hc2b01735, 32'hc274cd5d, 32'h4251b6d6, 32'h42101b48, 32'hc27dca1b};
test_weights[13760:13767] = '{32'hc219ca84, 32'h42b2e99b, 32'hc1a1482d, 32'hc2734488, 32'hc060939a, 32'h429ac0ec, 32'h422c7b4a, 32'h428548e4};
test_bias[1720:1720] = '{32'hc216b0f4};
test_output[1720:1720] = '{32'h46492db8};
test_input[13768:13775] = '{32'h42b0675d, 32'h4226b255, 32'hc259dc5c, 32'h41b93cd4, 32'hc2b70e7f, 32'hc2487cec, 32'hc2a7e8bf, 32'hc1e84144};
test_weights[13768:13775] = '{32'hc0395d30, 32'hc237398d, 32'h429bb4c8, 32'h42ba7f98, 32'h42af2306, 32'h42a2e120, 32'h42898fb8, 32'hc2b18529};
test_bias[1721:1721] = '{32'h428e2151};
test_output[1721:1721] = '{32'hc69819e6};
test_input[13776:13783] = '{32'hc27f53d0, 32'h42bd9b33, 32'hc24bd000, 32'hc1796b8a, 32'h42850dd1, 32'hc27b88fe, 32'h42ba3a8e, 32'hc2bf9a1a};
test_weights[13776:13783] = '{32'hc224bfd2, 32'hc2626797, 32'h4216486a, 32'h420df168, 32'hc19385d3, 32'h42213b00, 32'hc1195bb7, 32'h40f98da0};
test_bias[1722:1722] = '{32'hc28c6304};
test_output[1722:1722] = '{32'hc626cec8};
test_input[13784:13791] = '{32'h4281f05d, 32'hc294b67c, 32'hc21fb9d5, 32'h41f2791d, 32'hc29282a2, 32'h418c6965, 32'h428e9ad0, 32'h41f92eb5};
test_weights[13784:13791] = '{32'h4217ce29, 32'hc29956fa, 32'h4285ab51, 32'hc2907a8d, 32'h4253456b, 32'hc27eab2a, 32'h42c6cbbd, 32'h41db022b};
test_bias[1723:1723] = '{32'h422bc666};
test_output[1723:1723] = '{32'h45c504b1};
test_input[13792:13799] = '{32'hc1c4524c, 32'h4233c9e6, 32'hc2c458c0, 32'hc2700e82, 32'hc2ba161a, 32'hc2c0663e, 32'hc28d6166, 32'h422f747a};
test_weights[13792:13799] = '{32'hc2c47c37, 32'hc10e6c7c, 32'hc2985ab9, 32'h423f4194, 32'hc14fd5e8, 32'hc2560ce4, 32'hc294dcd0, 32'h41c2d2f3};
test_bias[1724:1724] = '{32'h3ea4dccf};
test_output[1724:1724] = '{32'h4696d4e3};
test_input[13800:13807] = '{32'hc2b4458b, 32'h427e9cb9, 32'h41658dbf, 32'h4265b868, 32'h42a5cb75, 32'h418ac542, 32'h41d15a0e, 32'h42706d67};
test_weights[13800:13807] = '{32'hc004060d, 32'hc25e4aef, 32'h429793ba, 32'hc1501fe4, 32'hc15356ae, 32'h42985953, 32'h428e59c2, 32'hc10725bf};
test_bias[1725:1725] = '{32'h425b1249};
test_output[1725:1725] = '{32'hc4abe404};
test_input[13808:13815] = '{32'hc2a80a57, 32'hc1908450, 32'h42ae5872, 32'h40e7be66, 32'h42b96510, 32'h422354e2, 32'h42c5d3ed, 32'h41dfea18};
test_weights[13808:13815] = '{32'hc1fb9be1, 32'h42772868, 32'hc2a6af47, 32'h429a9d3d, 32'hc29e3bc1, 32'h424353ab, 32'hc28552c0, 32'h42a34647};
test_bias[1726:1726] = '{32'h42be1a79};
test_output[1726:1726] = '{32'hc66632d6};
test_input[13816:13823] = '{32'hc2384f21, 32'h42704a1f, 32'h4235b16e, 32'h41797ae1, 32'h427f196e, 32'hc20a7394, 32'hc24036cd, 32'h4171fbf5};
test_weights[13816:13823] = '{32'hc20e2b77, 32'hbfb4ea3d, 32'h42a90cec, 32'hc212e8ef, 32'hc24cc866, 32'hc2a550bc, 32'hc0e4350f, 32'h42c6fd84};
test_bias[1727:1727] = '{32'h420dc17f};
test_output[1727:1727] = '{32'h45c4d39e};
test_input[13824:13831] = '{32'h4257743d, 32'hc29488a0, 32'h429cebf6, 32'h41a3fe9a, 32'hc1e05ce2, 32'h42503fcd, 32'h42b6befd, 32'hc19e4180};
test_weights[13824:13831] = '{32'h4210c77f, 32'h423cec55, 32'hc2814416, 32'hc26eaaac, 32'hc2bb39ac, 32'h41ca1677, 32'h4299f3f5, 32'hc0d87465};
test_bias[1728:1728] = '{32'hc14c048d};
test_output[1728:1728] = '{32'h454aaca0};
test_input[13832:13839] = '{32'h427ca0dd, 32'hc27e892c, 32'h40b9f778, 32'h42866437, 32'h428acc33, 32'hc19605ca, 32'h41b17aae, 32'hc1d4761f};
test_weights[13832:13839] = '{32'h42c1717d, 32'hc2812eb4, 32'h4283bd64, 32'h405608bd, 32'h41d8a149, 32'h4231b19d, 32'h42c579fb, 32'hc29a2516};
test_bias[1729:1729] = '{32'hbf29d8db};
test_output[1729:1729] = '{32'h467bb4f9};
test_input[13840:13847] = '{32'hc209f31b, 32'hc2950177, 32'h4201b2eb, 32'h42aa68a0, 32'hc1742d9b, 32'hc29653ed, 32'h42471891, 32'h42a9c0a8};
test_weights[13840:13847] = '{32'h4282156d, 32'hc21218c9, 32'hc25ffae5, 32'h4284cc89, 32'h41e7fc95, 32'hc23995eb, 32'hc2a4c779, 32'h3e861a19};
test_bias[1730:1730] = '{32'h3fb72baa};
test_output[1730:1730] = '{32'h454d7865};
test_input[13848:13855] = '{32'h42c2522a, 32'h422f9617, 32'h40b3cb6c, 32'hc2269a48, 32'hc1f108df, 32'hc26a7bd0, 32'h4260b421, 32'h42afb47e};
test_weights[13848:13855] = '{32'h4282037e, 32'h41804056, 32'hc2a4845f, 32'hc0fc2efe, 32'h42b5f50e, 32'hc269c898, 32'h41ad0e98, 32'hbf1933d9};
test_bias[1731:1731] = '{32'hc25286be};
test_output[1731:1731] = '{32'h4607a39d};
test_input[13856:13863] = '{32'hc2a4ea52, 32'h41a0e83e, 32'hc1f8475e, 32'hc19a7e25, 32'hc201ca2b, 32'hc247c3cf, 32'h4196bb03, 32'hbf85b6b0};
test_weights[13856:13863] = '{32'hc205aed9, 32'hc275876f, 32'h426b9e3d, 32'hc20294e5, 32'hc2006a4f, 32'h41f6d092, 32'hc28bd48b, 32'h42315b3c};
test_bias[1732:1732] = '{32'hc1ae2054};
test_output[1732:1732] = '{32'hc4c31df9};
test_input[13864:13871] = '{32'h424befae, 32'h4126ba64, 32'hc1bae121, 32'h427d1fbe, 32'hc2421089, 32'hc2960b3a, 32'hc24422da, 32'h42329e4a};
test_weights[13864:13871] = '{32'hc28b5de3, 32'hc28ed64b, 32'h42bdc5fa, 32'hc133d550, 32'hc28caba6, 32'h4135ed56, 32'h4285e9c3, 32'h4287768e};
test_bias[1733:1733] = '{32'hc285bf55};
test_output[1733:1733] = '{32'hc59bf726};
test_input[13872:13879] = '{32'h428c4852, 32'h4211b28a, 32'hc23ff31f, 32'h411196d7, 32'hc2bdf051, 32'h42344777, 32'h402e7e8a, 32'h41984749};
test_weights[13872:13879] = '{32'h41d4e7c4, 32'hc20d96a5, 32'hc2659c89, 32'hc2c243ba, 32'hc26a1aaa, 32'hc2bbd372, 32'h42450f05, 32'h42c1e8fe};
test_bias[1734:1734] = '{32'h41e3afde};
test_output[1734:1734] = '{32'h45b4afe1};
test_input[13880:13887] = '{32'h42af03aa, 32'h42a2455c, 32'h429f86eb, 32'h42c30a81, 32'hc2799ea4, 32'h42bb9887, 32'hc261513d, 32'hc2aade4d};
test_weights[13880:13887] = '{32'hc297cdaa, 32'hc29d93ef, 32'hc236ccab, 32'hc08ceee3, 32'hc28362e1, 32'h428bef4b, 32'h4221bae6, 32'hc2415291};
test_bias[1735:1735] = '{32'hc1ed608a};
test_output[1735:1735] = '{32'hc5908799};
test_input[13888:13895] = '{32'h4233e202, 32'hc193ab87, 32'hc2111ae2, 32'h429eca6f, 32'hc21146f5, 32'hc2966379, 32'h428b90a3, 32'h428f7c1d};
test_weights[13888:13895] = '{32'hc13eb386, 32'hc2a7373c, 32'hc1a6e237, 32'hc2716b99, 32'hc27ab395, 32'h42b5cebf, 32'hc274c67c, 32'hc2c52aaa};
test_bias[1736:1736] = '{32'hc23dbe9a};
test_output[1736:1736] = '{32'hc6944297};
test_input[13896:13903] = '{32'h416bf3a8, 32'h42193f03, 32'h4228048a, 32'h424656a6, 32'hc1339341, 32'hc27fb773, 32'h40e49086, 32'hc2af3b6b};
test_weights[13896:13903] = '{32'h41a85b2a, 32'h4224e3f0, 32'hc280d99a, 32'h42a4c06c, 32'hc25d032e, 32'h429b54ae, 32'hc214b572, 32'hc28e0372};
test_bias[1737:1737] = '{32'hc155a031};
test_output[1737:1737] = '{32'h45980c84};
test_input[13904:13911] = '{32'hc275d369, 32'h42605a94, 32'hc2ad8bdc, 32'h41e64256, 32'hc280f6c7, 32'h428ba32b, 32'hc109e6f6, 32'hc2bc6e22};
test_weights[13904:13911] = '{32'h420fc49b, 32'hc2789b2f, 32'h42bf1484, 32'h42bbb0a0, 32'hc270513a, 32'h400f7f29, 32'h423d731e, 32'h41cd65b0};
test_bias[1738:1738] = '{32'hc1dae40c};
test_output[1738:1738] = '{32'hc61df013};
test_input[13912:13919] = '{32'h4195fd08, 32'h429df8ae, 32'hc202428c, 32'h40e36eca, 32'h423ea9a2, 32'h428b6f64, 32'h4252cd3d, 32'hc2aaa3d3};
test_weights[13912:13919] = '{32'hc2a56919, 32'hc27e774e, 32'h4287a2fa, 32'h420245cc, 32'hc2a61dc1, 32'h40ddb186, 32'h420f5251, 32'h4263fcbd};
test_bias[1739:1739] = '{32'hc10c5762};
test_output[1739:1739] = '{32'hc66a8fa7};
test_input[13920:13927] = '{32'h42c3b72a, 32'hc2a885f3, 32'hc2970bd7, 32'h425a45bd, 32'hc20965ac, 32'h427b914c, 32'h42a7c0aa, 32'hc1ccf661};
test_weights[13920:13927] = '{32'hc29a740a, 32'hc240e29f, 32'hc1fb3035, 32'h425a90d6, 32'hc290d9f7, 32'h40c36697, 32'h4238deaf, 32'hc25af5a0};
test_bias[1740:1740] = '{32'hc1fbb722};
test_output[1740:1740] = '{32'h461be949};
test_input[13928:13935] = '{32'h42431c7d, 32'h3f196de0, 32'h429d1ba9, 32'h420b72e5, 32'h4281b286, 32'hc21b14a8, 32'hc2be4788, 32'hc2a5747b};
test_weights[13928:13935] = '{32'hc2999cfd, 32'hc2276a91, 32'hc1e047b3, 32'hc214e9e3, 32'hc232413f, 32'h4282e802, 32'hc18c4213, 32'hc1b82cc0};
test_bias[1741:1741] = '{32'hc1bd6094};
test_output[1741:1741] = '{32'hc60ef944};
test_input[13936:13943] = '{32'h429b755f, 32'hc2b6343a, 32'hc2bd08f3, 32'hc1b3a42a, 32'hc29c8237, 32'hc2603a51, 32'h42954fec, 32'hc1acc58e};
test_weights[13936:13943] = '{32'h42926419, 32'hc18e424d, 32'h41f8c5ce, 32'hc2143ca0, 32'h42c5e47e, 32'hc29343d4, 32'hc291ecf6, 32'hc2716227};
test_bias[1742:1742] = '{32'h42c37761};
test_output[1742:1742] = '{32'hc519b0cc};
test_input[13944:13951] = '{32'hc14518dc, 32'hc25271a6, 32'h41ed1826, 32'h4246d100, 32'h429ab330, 32'hc28c521d, 32'hc23cf1e1, 32'h42af9418};
test_weights[13944:13951] = '{32'h4245b6c6, 32'h41afe887, 32'hc2917973, 32'hc20552fd, 32'hc29caba3, 32'h3fe7bbc5, 32'h4166b9d1, 32'h423b0d79};
test_bias[1743:1743] = '{32'hc2c34926};
test_output[1743:1743] = '{32'hc603d777};
test_input[13952:13959] = '{32'h41dce249, 32'hc2194562, 32'hc25b128f, 32'hc0b14a68, 32'h4278ef6c, 32'h42a10b74, 32'hc28fec80, 32'h428c9ca3};
test_weights[13952:13959] = '{32'hc00bab09, 32'h42b3747d, 32'hc2bef0eb, 32'hc28819fe, 32'h41a1e509, 32'hc0c2d404, 32'hc2b70ad1, 32'h42272a19};
test_bias[1744:1744] = '{32'h42b52782};
test_output[1744:1744] = '{32'h46432d2d};
test_input[13960:13967] = '{32'h428a9d5e, 32'hc22da938, 32'h42a238e5, 32'h428912f3, 32'hc20df5f1, 32'hc1fabba2, 32'h411eecb9, 32'h40a7d3b8};
test_weights[13960:13967] = '{32'h4259b74a, 32'hc29f95eb, 32'hc22f8d6d, 32'h429e9a94, 32'hc1206bb7, 32'hc2c57b7e, 32'h414e65a9, 32'h427c9130};
test_bias[1745:1745] = '{32'h413a94ea};
test_output[1745:1745] = '{32'h464ba562};
test_input[13968:13975] = '{32'hc0f16ca9, 32'hc0bb0851, 32'h412bf437, 32'h422159b3, 32'hc1fabb65, 32'h42a0879c, 32'h42a64043, 32'h42701827};
test_weights[13968:13975] = '{32'h42bc1526, 32'h3e77085f, 32'hc28b61df, 32'h406deb02, 32'hc23938b3, 32'hc279d4c0, 32'h42a4d112, 32'hc1115242};
test_bias[1746:1746] = '{32'hc24aff99};
test_output[1746:1746] = '{32'h44acd009};
test_input[13976:13983] = '{32'hc2b2f366, 32'h417528d2, 32'hc2b62d7f, 32'hc276d54a, 32'hc22e181c, 32'hc2812ec2, 32'h42c1f40f, 32'h3f4653e6};
test_weights[13976:13983] = '{32'h41db1cbd, 32'h41471d7a, 32'hc299e2af, 32'h418a9139, 32'hc2a212f4, 32'h4254155b, 32'hc284517f, 32'h415e592e};
test_bias[1747:1747] = '{32'hc2139b45};
test_output[1747:1747] = '{32'hc5263e0f};
test_input[13984:13991] = '{32'h42104cdc, 32'h418f0930, 32'h4296ea5b, 32'hc27a164b, 32'h4254cf60, 32'hc2745878, 32'hc28e142c, 32'h423952f5};
test_weights[13984:13991] = '{32'h42b4060d, 32'h400e3f5d, 32'h40d76f65, 32'h42c0ddcc, 32'hc2a9c868, 32'h40eef3e3, 32'hc1abe8fe, 32'h429f86a4};
test_bias[1748:1748] = '{32'h42540bfa};
test_output[1748:1748] = '{32'hc4f178ae};
test_input[13992:13999] = '{32'hc21035b2, 32'hc13ecf56, 32'hc030a9c4, 32'hc2c6a8ee, 32'h4266f182, 32'hc16aaecf, 32'h42b7f4a6, 32'hc22e2285};
test_weights[13992:13999] = '{32'hc1cc7c6e, 32'hc2995144, 32'h42c6c64f, 32'hc2a938b8, 32'hc2ba6cab, 32'h42a3de7e, 32'h429836dd, 32'h42688861};
test_bias[1749:1749] = '{32'hc1c62df4};
test_output[1749:1749] = '{32'h45f4977f};
test_input[14000:14007] = '{32'h42b98c8b, 32'hc16dd6c1, 32'h410b20c0, 32'h41ba1bb4, 32'h427c588f, 32'hc201d03c, 32'h4154a8e7, 32'h41981bb9};
test_weights[14000:14007] = '{32'h4104678c, 32'hc2878823, 32'hc0fbda00, 32'h41374b4c, 32'h41f30706, 32'h4202ed12, 32'hc19f4d22, 32'h42c454ed};
test_bias[1750:1750] = '{32'h42b01ec2};
test_output[1750:1750] = '{32'h458d29e2};
test_input[14008:14015] = '{32'hc2b79107, 32'h41bac7ee, 32'hc1aa22ad, 32'hc28dd9ad, 32'hc2aedcd9, 32'hc1ee719c, 32'hc2592b58, 32'hc1d4843f};
test_weights[14008:14015] = '{32'h428ca291, 32'h41a5cdc9, 32'h42b30b04, 32'hc2bac5d8, 32'h421d2a60, 32'hc20e2973, 32'hc1badca4, 32'hc298a1d0};
test_bias[1751:1751] = '{32'hc2c1b336};
test_output[1751:1751] = '{32'hc3d5f0c7};
test_input[14016:14023] = '{32'h41f60651, 32'hc294b122, 32'hc21dc3aa, 32'hc2080779, 32'h40e222cf, 32'h42565772, 32'h425aafb7, 32'hc1fd1d12};
test_weights[14016:14023] = '{32'h424757e7, 32'hc21d543d, 32'hc29ef4d5, 32'hc191472f, 32'h42600606, 32'hc1ba711f, 32'hc1ee5aba, 32'h421a605c};
test_bias[1752:1752] = '{32'h42a574e9};
test_output[1752:1752] = '{32'h458f6629};
test_input[14024:14031] = '{32'hc2046443, 32'hc2b59c4a, 32'h42197cab, 32'h41876f42, 32'h41835023, 32'h421d83bf, 32'h42894a7f, 32'hc1f539c7};
test_weights[14024:14031] = '{32'hc204c575, 32'h425312bd, 32'h41e7e5e6, 32'hc220d607, 32'hc25f1086, 32'hc17867a4, 32'h429ffd2a, 32'hc25e2ece};
test_bias[1753:1753] = '{32'hc210539a};
test_output[1753:1753] = '{32'h45141ab7};
test_input[14032:14039] = '{32'h42747293, 32'h42bfc554, 32'hc278fab9, 32'h4215b514, 32'hc2c0946a, 32'hc2b19f2f, 32'hc2156aae, 32'h4204779c};
test_weights[14032:14039] = '{32'hc28484dd, 32'hc213ea13, 32'hc10d3eb2, 32'hbfff6a2f, 32'h423fc66e, 32'h410351bc, 32'h3f830379, 32'h41650eb9};
test_bias[1754:1754] = '{32'h3ff1d5f9};
test_output[1754:1754] = '{32'hc63bef33};
test_input[14040:14047] = '{32'h4193c201, 32'hc1b31616, 32'hc232fe15, 32'hc2b24b46, 32'hc2203f73, 32'h40d61713, 32'hc221eeed, 32'h40659054};
test_weights[14040:14047] = '{32'h42c41352, 32'h416699b7, 32'h412b016d, 32'h428e890b, 32'hc2833974, 32'h428bb122, 32'hc20d03bd, 32'hc219859b};
test_bias[1755:1755] = '{32'hc14a17b0};
test_output[1755:1755] = '{32'hc472af02};
test_input[14048:14055] = '{32'hc290298d, 32'hc191b091, 32'h4151c4ae, 32'h4149367a, 32'h42bcc3c3, 32'hc1795475, 32'hc2a5e06d, 32'hc25ac655};
test_weights[14048:14055] = '{32'hc28afc48, 32'hc1259b52, 32'h426993e7, 32'h41c1679f, 32'h42c2b953, 32'hc21183d3, 32'h41ce29ea, 32'hc288eaec};
test_bias[1756:1756] = '{32'hc213e883};
test_output[1756:1756] = '{32'h46897296};
test_input[14056:14063] = '{32'h403ba0d3, 32'hc27c3d87, 32'hc1bc77c6, 32'h4236a83c, 32'hc2207ac5, 32'hc282740f, 32'hc2aefff8, 32'h414c8aeb};
test_weights[14056:14063] = '{32'h42af1602, 32'h41dd931b, 32'hc2a017b7, 32'h422d81de, 32'hc27828ff, 32'hc1df5d29, 32'hc26be3d7, 32'h428371e3};
test_bias[1757:1757] = '{32'hc171f831};
test_output[1757:1757] = '{32'h4645ffef};
test_input[14064:14071] = '{32'hc2610701, 32'h42a4874b, 32'hc2890b18, 32'h42b0c76b, 32'hc20b0d95, 32'h4173fabf, 32'hc29a0c9d, 32'h423ca20d};
test_weights[14064:14071] = '{32'hc29477ca, 32'hc265b83a, 32'h42c269ed, 32'hc1a0404d, 32'hc29fde3f, 32'hc22f3bda, 32'hc1a691b7, 32'h410c46f8};
test_bias[1758:1758] = '{32'hc29ecba9};
test_output[1758:1758] = '{32'hc59a187b};
test_input[14072:14079] = '{32'h4038e0d1, 32'h42031f39, 32'h42b6264c, 32'hc1acb2d3, 32'hc29d109c, 32'hc2217692, 32'h423e18c1, 32'h423521da};
test_weights[14072:14079] = '{32'hc294c607, 32'h425d842e, 32'hc28fa684, 32'hc158c4d3, 32'hc2ac2ffb, 32'h42bd6d14, 32'hc2616e64, 32'h425324e3};
test_bias[1759:1759] = '{32'h42976d89};
test_output[1759:1759] = '{32'hc4f05c2a};
test_input[14080:14087] = '{32'h4274bc32, 32'hc26c27e0, 32'h406583c0, 32'hc2a0d314, 32'h426e1532, 32'h420824bb, 32'h4280c730, 32'hbf35070b};
test_weights[14080:14087] = '{32'hc11b974e, 32'h42c0c91b, 32'h41cc229e, 32'h42a5216d, 32'hc257b850, 32'h4231c3c8, 32'h41a918e5, 32'h42545170};
test_bias[1760:1760] = '{32'hc2c5ebfd};
test_output[1760:1760] = '{32'hc64fea0a};
test_input[14088:14095] = '{32'h42a17126, 32'h42b8447e, 32'h4285c478, 32'hc247bad8, 32'hc1afc14f, 32'h428ae3f2, 32'h424199af, 32'hc1f67deb};
test_weights[14088:14095] = '{32'h42439472, 32'hc234cba3, 32'h4282d3d5, 32'hc1c6e3a4, 32'hc0a41d98, 32'hc103db43, 32'h411b5845, 32'hc2c4da72};
test_bias[1761:1761] = '{32'hc1cd8ffc};
test_output[1761:1761] = '{32'h46038113};
test_input[14096:14103] = '{32'hc2854a9a, 32'hc2b33df4, 32'h4273fa37, 32'h428d50fd, 32'h422df9ed, 32'hc1d4a83e, 32'hc13330f3, 32'h41bc108b};
test_weights[14096:14103] = '{32'hc2210365, 32'hc2ad62fb, 32'hc2a7945f, 32'h429372f8, 32'hc124e6b8, 32'hc2ab1449, 32'h4222b98d, 32'h4056847a};
test_bias[1762:1762] = '{32'hc28da031};
test_output[1762:1762] = '{32'h463a62eb};
test_input[14104:14111] = '{32'h4205165a, 32'hc214f19f, 32'h41b3c361, 32'h418370e8, 32'hc2af822c, 32'hc1e28a3d, 32'h42809284, 32'h41f9aafb};
test_weights[14104:14111] = '{32'h42bdd2f4, 32'hc1e130ec, 32'h41b668fc, 32'hc194ea60, 32'h428899bd, 32'h42483e84, 32'h41e75561, 32'h42b5d5e5};
test_bias[1763:1763] = '{32'h42c63de3};
test_output[1763:1763] = '{32'h44e09949};
test_input[14112:14119] = '{32'hc05a1796, 32'h4224137f, 32'h42c2ff7f, 32'hc27448d9, 32'hc24223de, 32'h428f0ed2, 32'hc1edbc20, 32'h3e47ba0b};
test_weights[14112:14119] = '{32'hc296c531, 32'hc00b7bcf, 32'hc12e7eef, 32'hc256f1c9, 32'hc2235b18, 32'hbfe88039, 32'hc19798df, 32'hc2238c01};
test_bias[1764:1764] = '{32'hc23ec6a7};
test_output[1764:1764] = '{32'h45944c57};
test_input[14120:14127] = '{32'h42820ef1, 32'h429cbe08, 32'h4280b3e0, 32'h425ec351, 32'hbf9d9633, 32'hc1dd1280, 32'h4257db1e, 32'hc10f0af3};
test_weights[14120:14127] = '{32'hc2b8f7c7, 32'h3f33c96a, 32'hc296d9a4, 32'hc28996d0, 32'hc113de1b, 32'h429d3dea, 32'hc1343459, 32'hc25aacd3};
test_bias[1765:1765] = '{32'h42020fb9};
test_output[1765:1765] = '{32'hc683f797};
test_input[14128:14135] = '{32'h429099ec, 32'hc2ae8224, 32'hc21c266c, 32'hc1d3a604, 32'hc2535c02, 32'hc2a8ce13, 32'hc25a2e0b, 32'h428ec404};
test_weights[14128:14135] = '{32'h420da92a, 32'h3f99071b, 32'h42b69983, 32'h427582d5, 32'hc2adf58c, 32'hc1a31832, 32'h40fd6632, 32'h42ab2883};
test_bias[1766:1766] = '{32'h42c6db8c};
test_output[1766:1766] = '{32'h46124574};
test_input[14136:14143] = '{32'h412ea950, 32'hc24169e3, 32'hc25c3936, 32'hc2920348, 32'hc151af2e, 32'hc2951a71, 32'h42b6cb9e, 32'hc23aa7e7};
test_weights[14136:14143] = '{32'h427e4238, 32'h4246fd24, 32'h40ab7a42, 32'hc2b6b7c1, 32'h428874c0, 32'h42928f84, 32'hc2a1c50b, 32'hc2863b94};
test_bias[1767:1767] = '{32'hc26d6142};
test_output[1767:1767] = '{32'hc5bbf1cf};
test_input[14144:14151] = '{32'h42ad956b, 32'h41ba31c2, 32'hc04c238e, 32'h4242cba4, 32'hc2b75966, 32'hc2941103, 32'h428a7d4b, 32'h412b83bf};
test_weights[14144:14151] = '{32'hbeb4f427, 32'hc2235249, 32'hc2484f77, 32'hc20fbb70, 32'hc1fa08aa, 32'h41456604, 32'h42571969, 32'h42941d35};
test_bias[1768:1768] = '{32'hc194d51a};
test_output[1768:1768] = '{32'h4572795f};
test_input[14152:14159] = '{32'h426bc545, 32'hc1e9dca4, 32'h42b85718, 32'hc1e58060, 32'h42810080, 32'h429b1eeb, 32'hc1d357bd, 32'h41d67db6};
test_weights[14152:14159] = '{32'h42a6d9bf, 32'hc28934c6, 32'h41d7da67, 32'h41bec939, 32'h422ee026, 32'hc297adca, 32'hc2a5bcec, 32'hc2a52ca4};
test_bias[1769:1769] = '{32'h42b8ce43};
test_output[1769:1769] = '{32'h45b31512};
test_input[14160:14167] = '{32'h4282c01a, 32'h428af27f, 32'hc2a8c643, 32'hc2bf22ed, 32'h427f021c, 32'h409bf39e, 32'hc21f5ae6, 32'hc20dea52};
test_weights[14160:14167] = '{32'h42b4996f, 32'h42440314, 32'hc2ac94ec, 32'hc1ed57dc, 32'h41cd6a96, 32'h4213c437, 32'h42a3d5a3, 32'h4221497c};
test_bias[1770:1770] = '{32'h42a1c9af};
test_output[1770:1770] = '{32'h4681e98b};
test_input[14168:14175] = '{32'h42c78d85, 32'h42aa6728, 32'h42a626ca, 32'hc267ece9, 32'hc222e7ac, 32'hc23adaf5, 32'h426928f8, 32'hc1b0d125};
test_weights[14168:14175] = '{32'h425ac247, 32'h422f29dc, 32'h4272ab24, 32'h413f5da7, 32'h41f19fda, 32'h41efd644, 32'hc2901f82, 32'h405c8cff};
test_bias[1771:1771] = '{32'h426dce12};
test_output[1771:1771] = '{32'h45d0f4a0};
test_input[14176:14183] = '{32'hc2c1822e, 32'hc1e25be7, 32'h425df6f7, 32'hc1bfb92d, 32'hc283166a, 32'hc2b3108f, 32'h427c637f, 32'h428dc28b};
test_weights[14176:14183] = '{32'hc22c61c1, 32'hc1403e32, 32'h40c9ea5b, 32'hc1b58671, 32'h429a48e0, 32'h429c799f, 32'hc2b5a15d, 32'h406f3d1b};
test_bias[1772:1772] = '{32'hc2547bf7};
test_output[1772:1772] = '{32'hc63e3f0e};
test_input[14184:14191] = '{32'hc133d75a, 32'h4181d0e4, 32'h42ba8161, 32'hc2a21af8, 32'h41edad18, 32'hc26f2091, 32'h4299d36f, 32'h41a06d8c};
test_weights[14184:14191] = '{32'hc2a490f6, 32'h42b86375, 32'hc27949d2, 32'hc2647c93, 32'hc2134fa5, 32'h4212fb1c, 32'h427618b6, 32'h4298c9a4};
test_bias[1773:1773] = '{32'h423d9210};
test_output[1773:1773] = '{32'h45851cbd};
test_input[14192:14199] = '{32'h3e866353, 32'h4295cbe5, 32'hc29b2df1, 32'hc1867ab2, 32'h41f978b2, 32'hc2693198, 32'h40da06b2, 32'hc2a1aafd};
test_weights[14192:14199] = '{32'hc2a48853, 32'hc13c94e1, 32'hc2777159, 32'h423bbf42, 32'hc1c642a2, 32'hc020a766, 32'h42942046, 32'hc2ab2d6a};
test_bias[1774:1774] = '{32'h413dbfe6};
test_output[1774:1774] = '{32'h461aeb6a};
test_input[14200:14207] = '{32'hc0cf38cf, 32'hc253f5af, 32'h42b32b88, 32'h42b12eef, 32'hc12f901a, 32'h4285ea8f, 32'h42c709e5, 32'h4219dd7a};
test_weights[14200:14207] = '{32'h4268db00, 32'hc2109ece, 32'hc16f18d2, 32'hc2ad6fcb, 32'hc2b43c49, 32'hc2b69e45, 32'h426ddfa1, 32'h429e5c18};
test_bias[1775:1775] = '{32'h42acb73a};
test_output[1775:1775] = '{32'hc55e50c6};
test_input[14208:14215] = '{32'hc28c2606, 32'h42a25be3, 32'hc23b5850, 32'hc2a5f1f8, 32'hc2b45905, 32'hc28fadb1, 32'h42627854, 32'hc21daa30};
test_weights[14208:14215] = '{32'hc242c28b, 32'h419efe8e, 32'hc0627e5e, 32'h40a65562, 32'h42b38643, 32'h426f2499, 32'h418fc454, 32'h42b45928};
test_bias[1776:1776] = '{32'hc1b3206c};
test_output[1776:1776] = '{32'hc61f329a};
test_input[14216:14223] = '{32'h41d9741f, 32'hc2363f8a, 32'hc2291ad2, 32'h42ad318b, 32'h402ca49a, 32'h42acfffe, 32'hc27bf697, 32'h42715fde};
test_weights[14216:14223] = '{32'h420251f1, 32'h424a0f11, 32'hbede60ec, 32'h4276b99f, 32'h4005695a, 32'hc1c1b5c2, 32'h4050346d, 32'hc24ac277};
test_bias[1777:1777] = '{32'h425ebf8d};
test_output[1777:1777] = '{32'hc4a92408};
test_input[14224:14231] = '{32'hc1317094, 32'hc24b3a38, 32'hc1bca8aa, 32'h42a79d53, 32'hc29157d3, 32'hc2c4b475, 32'hc1cca5bc, 32'hc1acab59};
test_weights[14224:14231] = '{32'hc266c20c, 32'hc22c2d02, 32'hc257090c, 32'h42b2c9fb, 32'h42b43bf7, 32'hc2b44e2a, 32'hc2b3fc9c, 32'h42b5a4f4};
test_bias[1778:1778] = '{32'hc192bc8c};
test_output[1778:1778] = '{32'h465e4e9f};
test_input[14232:14239] = '{32'h42a9303b, 32'hc231d2d9, 32'hc289d0d4, 32'hc228cf2a, 32'hc26d1bc6, 32'h421abd20, 32'hc20580b1, 32'hc24d30bc};
test_weights[14232:14239] = '{32'h42851a16, 32'hc1def486, 32'hc2ab8a27, 32'hc2a0f3ab, 32'h4299ccbc, 32'h41eae637, 32'hc2a9d1e9, 32'h41d8cf62};
test_bias[1779:1779] = '{32'hc25e6ce7};
test_output[1779:1779] = '{32'h465cf356};
test_input[14240:14247] = '{32'hc1447217, 32'h42b63443, 32'h42190d2f, 32'h40bdacd3, 32'h429ffe99, 32'h42649c41, 32'hc2535dbf, 32'h41943f09};
test_weights[14240:14247] = '{32'h42c29d6b, 32'h429b10c2, 32'h42c473cf, 32'h40ea34be, 32'h42337561, 32'hc2681f35, 32'h4171417c, 32'h42266142};
test_bias[1780:1780] = '{32'h4185b332};
test_output[1780:1780] = '{32'h461b3699};
test_input[14248:14255] = '{32'h420cd781, 32'hc09b477c, 32'h40906a37, 32'hc23ac911, 32'h42a062dc, 32'hc1f44619, 32'hc23385ad, 32'hc0ec1473};
test_weights[14248:14255] = '{32'h4201b2c0, 32'h422279be, 32'hc26a2e66, 32'hc1b7e075, 32'hc29344c3, 32'h418bd096, 32'hc124465a, 32'hc14d390f};
test_bias[1781:1781] = '{32'h42b4c74c};
test_output[1781:1781] = '{32'hc57c7203};
test_input[14256:14263] = '{32'h412cd356, 32'hc28298f5, 32'h42b1e487, 32'h41a98f6d, 32'h41da8ab5, 32'h424a7d10, 32'hc28d8091, 32'hc19169fb};
test_weights[14256:14263] = '{32'hc22709c1, 32'hc1b56b20, 32'h41e86554, 32'h4260ee24, 32'hc299cce5, 32'hc24c1cfc, 32'hc2a02efd, 32'h425116bb};
test_bias[1782:1782] = '{32'hc29a3382};
test_output[1782:1782] = '{32'h4594c6f3};
test_input[14264:14271] = '{32'h423a9d34, 32'hc2775cbb, 32'hc2af7cca, 32'hc26a5daa, 32'h42b72237, 32'h419bf107, 32'h420e0f5c, 32'h41518a3c};
test_weights[14264:14271] = '{32'hc2376751, 32'hc2af2de7, 32'hc0b5b896, 32'hc105474d, 32'h4244e773, 32'hc2c3c7cd, 32'hc2b80a4d, 32'h41cc3ae8};
test_bias[1783:1783] = '{32'hc249e4c5};
test_output[1783:1783] = '{32'h45726eab};
test_input[14272:14279] = '{32'hc2bffbd9, 32'h411035dc, 32'hc2720d43, 32'hc1fa867b, 32'h408b1b83, 32'h4236b063, 32'h4295216c, 32'h41b7ea1b};
test_weights[14272:14279] = '{32'hc24a49ce, 32'h4294d2a5, 32'h41383f46, 32'h42a187d9, 32'h41db0577, 32'hc199b63a, 32'h41b87ca1, 32'hc236121e};
test_bias[1784:1784] = '{32'h4296da2b};
test_output[1784:1784] = '{32'h450f1264};
test_input[14280:14287] = '{32'hc1f02cb2, 32'hc2ab255d, 32'hc1df09ec, 32'h42529673, 32'hc13aefa7, 32'hc1c28c01, 32'hc2abfefe, 32'h42506af3};
test_weights[14280:14287] = '{32'hc2b3fbb0, 32'h428fa90c, 32'hc215f7a4, 32'hc2a1a8b7, 32'hc2a2c254, 32'h41e54e6d, 32'h4110a96e, 32'hc1ffa923};
test_bias[1785:1785] = '{32'h426892c6};
test_output[1785:1785] = '{32'hc60947c5};
test_input[14288:14295] = '{32'h42bef613, 32'h427833f5, 32'hc234bfc9, 32'hc296e4af, 32'hc194676e, 32'h429b6a62, 32'hc241cc2c, 32'h42944451};
test_weights[14288:14295] = '{32'h41b03860, 32'h428ab8ad, 32'hc2023690, 32'hc1ecbb7f, 32'h41f61b32, 32'hc1a13e1f, 32'h420e7a1a, 32'h423dbae3};
test_bias[1786:1786] = '{32'h42b88dcd};
test_output[1786:1786] = '{32'h461a0293};
test_input[14296:14303] = '{32'h42697fde, 32'h42b1eb2c, 32'hc2acdebd, 32'hc1f58e6c, 32'hc13d4e55, 32'h42a5802c, 32'h42a16150, 32'h4195f7cb};
test_weights[14296:14303] = '{32'hc1e99a28, 32'h41a67b93, 32'hc2a0dae8, 32'h4299ecfb, 32'hbf010603, 32'hc1c22cc0, 32'h427f3076, 32'hc1027a51};
test_bias[1787:1787] = '{32'h423b25b0};
test_output[1787:1787] = '{32'h45f2fa85};
test_input[14304:14311] = '{32'h42934fee, 32'h428af9ba, 32'hc202fbfa, 32'hc2adb700, 32'h4299ba30, 32'hc28a4825, 32'hc07b0cff, 32'hc1f4f975};
test_weights[14304:14311] = '{32'hc1134030, 32'h42a0a0d8, 32'hc285bf28, 32'h42aa4a43, 32'hc287f764, 32'hc29cd42e, 32'h42ade2dd, 32'h42990744};
test_bias[1788:1788] = '{32'h423ca855};
test_output[1788:1788] = '{32'hc52b756c};
test_input[14312:14319] = '{32'hbf30bdde, 32'hc2887666, 32'h4227236c, 32'h41dfc752, 32'hc288b0b7, 32'hc25fecd1, 32'hc297a8f9, 32'h42c4c15b};
test_weights[14312:14319] = '{32'hc239e20a, 32'h42520991, 32'hc209aa09, 32'h42a3108f, 32'hc28f27b2, 32'hc2bbe09f, 32'hc229ff47, 32'hc144d392};
test_bias[1789:1789] = '{32'hc19437d0};
test_output[1789:1789] = '{32'h461372aa};
test_input[14320:14327] = '{32'hc1e77370, 32'hc229f5d5, 32'hc23b2e4d, 32'hc29f9cd1, 32'hc1fc8b3c, 32'h42b3750f, 32'h41192132, 32'hc14f5491};
test_weights[14320:14327] = '{32'h40dfd2fc, 32'hc2a2c89d, 32'hc2be78a9, 32'h42b1c0e0, 32'h4177e85a, 32'h429a3f8e, 32'hc211b8f8, 32'hc1933838};
test_bias[1790:1790] = '{32'hc23986c8};
test_output[1790:1790] = '{32'h45d77167};
test_input[14328:14335] = '{32'h427e5ed4, 32'hc2bb4ddf, 32'h41a692b5, 32'h41e9ef64, 32'hc2506eae, 32'h416390c7, 32'h423c792e, 32'h4279372d};
test_weights[14328:14335] = '{32'hc25e976d, 32'hbff47c96, 32'h423a79c8, 32'hc1d0918d, 32'hc2773da0, 32'hc2a26ece, 32'h42561c23, 32'hc2832abf};
test_bias[1791:1791] = '{32'h42afcfbc};
test_output[1791:1791] = '{32'hc5201fdb};
test_input[14336:14343] = '{32'hc15b04d8, 32'h42a96b99, 32'h42525e92, 32'h427168ba, 32'h40fbf067, 32'hc261eef7, 32'h4200e07c, 32'h42c2c6a6};
test_weights[14336:14343] = '{32'hbc77fe9e, 32'h420655f8, 32'hc299a1ef, 32'hc22664c2, 32'hc2bf0f4b, 32'h42bf645e, 32'h42146f52, 32'hc106e1b8};
test_bias[1792:1792] = '{32'h423d44f2};
test_output[1792:1792] = '{32'hc613833b};
test_input[14344:14351] = '{32'h4218de1e, 32'hc2201fff, 32'hc2abadc6, 32'hc2c305cb, 32'hbf936b0b, 32'hc2b42698, 32'hc287dc86, 32'h42c063c1};
test_weights[14344:14351] = '{32'h4129b91a, 32'h42726e0f, 32'hc0d3cbe4, 32'hc2a95e31, 32'hc274b8b3, 32'h42c50439, 32'h417eb5b3, 32'hc0c438d4};
test_bias[1793:1793] = '{32'h424dd5aa};
test_output[1793:1793] = '{32'hc5621895};
test_input[14352:14359] = '{32'h429f633b, 32'h42beaf10, 32'hc0fbba10, 32'hc18a3271, 32'h41de56fd, 32'h419d2a5b, 32'hc2a861b7, 32'h42b8171c};
test_weights[14352:14359] = '{32'hc28c0ca1, 32'hc2602f85, 32'hc21b4fe6, 32'h42402c3f, 32'hc2315f75, 32'hc2bf70a0, 32'h42b96341, 32'h42244964};
test_bias[1794:1794] = '{32'h42802277};
test_output[1794:1794] = '{32'hc690b1e4};
test_input[14360:14367] = '{32'h4299830b, 32'hc20bd4fd, 32'hc231f487, 32'h42889c04, 32'h4285c556, 32'h4267ff71, 32'hc25df1f2, 32'h429e83f1};
test_weights[14360:14367] = '{32'h42531793, 32'hc21b712d, 32'hc195cc8c, 32'h420b08a8, 32'hc2b99522, 32'h41952d06, 32'h425a00cf, 32'h411e301d};
test_bias[1795:1795] = '{32'hc24577c2};
test_output[1795:1795] = '{32'h44963531};
test_input[14368:14375] = '{32'hc28cbc81, 32'hc2a5209b, 32'h410c7bd9, 32'hc0bbeb45, 32'hc11838db, 32'hc1189b98, 32'h426a5ce0, 32'hc1b5c1bd};
test_weights[14368:14375] = '{32'hc24f06df, 32'hc1873c2f, 32'hc284766a, 32'hc2ad0745, 32'hc273cca3, 32'hbfe15a35, 32'h42c27415, 32'hc1dffd2c};
test_bias[1796:1796] = '{32'h42578e03};
test_output[1796:1796] = '{32'h463aadf4};
test_input[14376:14383] = '{32'hc292f536, 32'hc20c94cb, 32'hc0ffdf24, 32'hc20b247e, 32'h4206e8c6, 32'h3f7afb11, 32'h4234e745, 32'hc2b51d11};
test_weights[14376:14383] = '{32'hc1fd119b, 32'h42aadc6d, 32'hc252e27d, 32'h42240071, 32'h429f5dd2, 32'h40d4af2f, 32'hc2c1c933, 32'h4118341a};
test_bias[1797:1797] = '{32'hc2b95a03};
test_output[1797:1797] = '{32'hc587274d};
test_input[14384:14391] = '{32'hc1f074bd, 32'h42389b5d, 32'hc2c3c7bd, 32'h42915462, 32'h40408bd8, 32'hc287d7bb, 32'h428a1f2d, 32'h425a86a1};
test_weights[14384:14391] = '{32'h423c2d57, 32'hc29fccd9, 32'h4235e4d1, 32'h4217fbef, 32'hc2a661f9, 32'hc203c6db, 32'hc1ebcebf, 32'hc2a35164};
test_bias[1798:1798] = '{32'h408ab21b};
test_output[1798:1798] = '{32'hc6308457};
test_input[14392:14399] = '{32'hc1faa821, 32'hc10bcb70, 32'hc2891a81, 32'hc1dc7d3e, 32'h41071484, 32'hc28e31e2, 32'hc21a41a2, 32'h429e86f3};
test_weights[14392:14399] = '{32'h425324c5, 32'h42304303, 32'hc2838571, 32'hc20f2dc2, 32'hc1265027, 32'h42290b32, 32'hc2b8fa15, 32'h42acda3c};
test_bias[1799:1799] = '{32'hc2c0796b};
test_output[1799:1799] = '{32'h4626f0cb};
test_input[14400:14407] = '{32'h427eb25f, 32'h42ad1521, 32'h4287cb58, 32'hc2aacd64, 32'h4119eb59, 32'hc2a10332, 32'h42c0906e, 32'hc1fae560};
test_weights[14400:14407] = '{32'h42b03d3c, 32'h4204f294, 32'hc2b96f3b, 32'h421ac349, 32'hc13a16f4, 32'h425c0c80, 32'h428af6b6, 32'hc1c3a702};
test_bias[1800:1800] = '{32'h4179af8a};
test_output[1800:1800] = '{32'h44e3731a};
test_input[14408:14415] = '{32'h41bd87d4, 32'hc22564ca, 32'h41ef49d5, 32'hc281a430, 32'h42a7656c, 32'hc2ba9643, 32'hc254c12b, 32'h42670a6c};
test_weights[14408:14415] = '{32'hc1977a26, 32'h4208c5c9, 32'h40ec4dfa, 32'h42bbc4b5, 32'h42bfd5d8, 32'h42c557a9, 32'hc23e4e35, 32'hc239904d};
test_bias[1801:1801] = '{32'hc23292d4};
test_output[1801:1801] = '{32'hc60e2868};
test_input[14416:14423] = '{32'h42020cad, 32'hc2a3df20, 32'hc0f1356c, 32'hc1e95ea4, 32'h41dcbadb, 32'hc08f203d, 32'hc29dba42, 32'hc2a7c4c9};
test_weights[14416:14423] = '{32'h41f0dc3b, 32'hc22019cc, 32'h41dfa51e, 32'hc24e5d94, 32'hc17f0548, 32'h41b40d92, 32'hc1909a5d, 32'hc13f90e4};
test_bias[1802:1802] = '{32'hc1216729};
test_output[1802:1802] = '{32'h45e83f6e};
test_input[14424:14431] = '{32'h42a8fe59, 32'h42a48e18, 32'hc2a1a2b6, 32'h420a3318, 32'h413b9a8e, 32'hc1457f8c, 32'h4251d082, 32'hc21e91f6};
test_weights[14424:14431] = '{32'h42ba7a93, 32'hc2acddfe, 32'h429f036e, 32'hc116429f, 32'h41b3fac4, 32'h424d38b1, 32'h420615b8, 32'hc28c30d2};
test_bias[1803:1803] = '{32'hc29dae39};
test_output[1803:1803] = '{32'hc4eccd51};
test_input[14432:14439] = '{32'hc28d4cab, 32'h42aa9a2d, 32'h428f66dd, 32'hc11d47f6, 32'hc29cb9c0, 32'hc11bb64c, 32'hc258e0d5, 32'h41f37019};
test_weights[14432:14439] = '{32'h4221ab5e, 32'hc27966b9, 32'h42ad662d, 32'hc2051d00, 32'h421db4ec, 32'h4256623d, 32'hc241f6e1, 32'hc186d922};
test_bias[1804:1804] = '{32'hc2726674};
test_output[1804:1804] = '{32'hc5472008};
test_input[14440:14447] = '{32'h41a69e0e, 32'h4281c083, 32'h423f4f94, 32'hc2b4bebd, 32'h40d0fc56, 32'hc2b64295, 32'hc0a0bb78, 32'hc20d2277};
test_weights[14440:14447] = '{32'hc2bab045, 32'h42b17aab, 32'hc2a44454, 32'h42938219, 32'hc2c17896, 32'hbfc88336, 32'hc2a6fbc9, 32'h42a5699f};
test_bias[1805:1805] = '{32'h429be8a1};
test_output[1805:1805] = '{32'hc61769f6};
test_input[14448:14455] = '{32'hc2a2b55f, 32'h40b57425, 32'hc1f6b36d, 32'hc1754d07, 32'h4297976a, 32'h42c4aaa7, 32'h42918a3c, 32'h4108031b};
test_weights[14448:14455] = '{32'h4277ed03, 32'h427a8620, 32'hc0d0d20e, 32'h42247c6f, 32'h42968980, 32'h425ca7e8, 32'hbffdf49d, 32'hc2b63c10};
test_bias[1806:1806] = '{32'hc089dc51};
test_output[1806:1806] = '{32'h459f0dbe};
test_input[14456:14463] = '{32'h429f84e9, 32'h42c13bb7, 32'hc2c13011, 32'hc16b5f52, 32'hc158f53e, 32'hc2938dc3, 32'hc1e62fcc, 32'hc155469d};
test_weights[14456:14463] = '{32'h428bdac3, 32'hc224873d, 32'hc21c04e9, 32'hc262ee97, 32'hc0e72264, 32'h42a6f89f, 32'hc2917ee7, 32'h41ef9f75};
test_bias[1807:1807] = '{32'hc29aadcb};
test_output[1807:1807] = '{32'h44dc18ad};
test_input[14464:14471] = '{32'hc2ad3c2a, 32'hc0c9d4ea, 32'hc1dcdc0c, 32'h41937275, 32'hc294184b, 32'h4248d70b, 32'hc2841fe0, 32'hc142369e};
test_weights[14464:14471] = '{32'hc26a6b67, 32'hc212715d, 32'hc260919f, 32'hc2abfa24, 32'hc1d8a4bf, 32'hc289f454, 32'h429322a2, 32'hc12ceb44};
test_bias[1808:1808] = '{32'h4235b240};
test_output[1808:1808] = '{32'hc45954ce};
test_input[14472:14479] = '{32'hc22ead45, 32'hc275897f, 32'hc294b06a, 32'hc277b50c, 32'hc21edcfc, 32'h42099a58, 32'h41858bc8, 32'h409d97f1};
test_weights[14472:14479] = '{32'hc129af28, 32'hc27023bf, 32'hc262051b, 32'h422ee003, 32'h42a3c918, 32'h424d7531, 32'hc2aaba43, 32'h415b93cc};
test_bias[1809:1809] = '{32'h429b0cc2};
test_output[1809:1809] = '{32'h4533c727};
test_input[14480:14487] = '{32'h426f1cd8, 32'h4274f966, 32'hc04a223a, 32'hc15aa17e, 32'hc2b92c54, 32'hc16e2b47, 32'h4176a8bf, 32'h41b4119b};
test_weights[14480:14487] = '{32'hc0c62a36, 32'hc201fb8d, 32'hc2302ba3, 32'hc2adfad9, 32'h426638a4, 32'h42b675b0, 32'h422c7724, 32'hc1b18298};
test_bias[1810:1810] = '{32'hc20c8be7};
test_output[1810:1810] = '{32'hc5ed2a77};
test_input[14488:14495] = '{32'h412f0ef9, 32'hc21782c2, 32'hc22dd204, 32'hc2be36a1, 32'hc2b71a0c, 32'hc2aff697, 32'h42abd71e, 32'hc283f4b7};
test_weights[14488:14495] = '{32'h41808438, 32'h423f237d, 32'h42912968, 32'h3ed2da9d, 32'h42afd8e7, 32'hc0e85c83, 32'hc2956b4b, 32'h42b92528};
test_bias[1811:1811] = '{32'hc2326a72};
test_output[1811:1811] = '{32'hc6c1d2d7};
test_input[14496:14503] = '{32'h42c38617, 32'hc2ad80dc, 32'hc29f2403, 32'h42795d9f, 32'h42b93cc2, 32'hc25a0d9a, 32'hbf32aef0, 32'hc108b54b};
test_weights[14496:14503] = '{32'hc2c071df, 32'h42928572, 32'h41e75c36, 32'h40a97a26, 32'hc2728c8a, 32'h42c6a8ec, 32'h42bc829c, 32'hc2bb1426};
test_bias[1812:1812] = '{32'hc2c7aba2};
test_output[1812:1812] = '{32'hc6dbc56d};
test_input[14504:14511] = '{32'hc2bc3715, 32'h41f5c254, 32'h418c6842, 32'h42aaa3b3, 32'hc2a50091, 32'h423052dd, 32'hc1acf83c, 32'hc19afde3};
test_weights[14504:14511] = '{32'hc0fee725, 32'hc2a0453a, 32'hc1528760, 32'h415eee83, 32'h413c7067, 32'hc2a63f29, 32'hc28c7cec, 32'hc27b2196};
test_bias[1813:1813] = '{32'h42ada26b};
test_output[1813:1813] = '{32'hc520824c};
test_input[14512:14519] = '{32'hc27618c2, 32'hc2829a90, 32'h4268dc8a, 32'hc24e823e, 32'h4280c053, 32'h42b3cf80, 32'h428132ec, 32'h42b9a677};
test_weights[14512:14519] = '{32'hc202488a, 32'h42aaa362, 32'h42265300, 32'h41c45d89, 32'h401f2bc4, 32'hc20ae7dd, 32'h42ac242d, 32'h419cc24b};
test_bias[1814:1814] = '{32'h420e708f};
test_output[1814:1814] = '{32'h44fecefc};
test_input[14520:14527] = '{32'hc26a6286, 32'hc215e0c3, 32'h4184fdcc, 32'hc29fb7fc, 32'hc2a19d0b, 32'h41aefb83, 32'h41e199bd, 32'hc25473ca};
test_weights[14520:14527] = '{32'hc18d2707, 32'hc26e2331, 32'h42528df7, 32'hc205851b, 32'hc065ad73, 32'h40faa887, 32'h421e9d4d, 32'hc02b9c2c};
test_bias[1815:1815] = '{32'hc26b4bb8};
test_output[1815:1815] = '{32'h4604520e};
test_input[14528:14535] = '{32'hbc5169a5, 32'hc2521853, 32'h42a07cc1, 32'hc2a4d30e, 32'hc1c0b164, 32'h4200ebe0, 32'hc280cda0, 32'h42b498a2};
test_weights[14528:14535] = '{32'hc285ec62, 32'h423cad5c, 32'h41aed8d6, 32'hc2c25534, 32'hc23c4e7a, 32'h4299938b, 32'h428efa3b, 32'h424a875d};
test_bias[1816:1816] = '{32'h42172f1d};
test_output[1816:1816] = '{32'h462a4dde};
test_input[14536:14543] = '{32'hc26777f5, 32'hc2a2b629, 32'hc2bd4603, 32'hc240706e, 32'h41423623, 32'hc292cd25, 32'hc2c1ab11, 32'h41ec1eef};
test_weights[14536:14543] = '{32'hc23b2e42, 32'h428f0fa5, 32'hc1a3b4b4, 32'hc2a90743, 32'hc1cec363, 32'hc1297bc2, 32'hc25f0394, 32'hc2bf93eb};
test_bias[1817:1817] = '{32'hbf8f77d7};
test_output[1817:1817] = '{32'h45b92a76};
test_input[14544:14551] = '{32'h4178842f, 32'hc245421c, 32'hc28ef33a, 32'hc1cb11e2, 32'hc2664858, 32'h420687d3, 32'h42505bed, 32'hc208b0b6};
test_weights[14544:14551] = '{32'h42ac836b, 32'hc280e235, 32'hc08c9351, 32'hc236a01a, 32'h4200a280, 32'h425ffb28, 32'hc28bdcb5, 32'h4069632c};
test_bias[1818:1818] = '{32'hc2196b1e};
test_output[1818:1818] = '{32'h450a8ce7};
test_input[14552:14559] = '{32'hc2bf83b8, 32'h4295ab14, 32'h424455d2, 32'h4197c2c3, 32'h42a34ecd, 32'h41c90efd, 32'h42c29e29, 32'h41a128ac};
test_weights[14552:14559] = '{32'h42b82caf, 32'hc2c04121, 32'h413fef0d, 32'hc094c7cd, 32'h427c24a1, 32'hc29b74a8, 32'h42bb0b18, 32'h40e1efe4};
test_bias[1819:1819] = '{32'h41d1ab74};
test_output[1819:1819] = '{32'hc53e872f};
test_input[14560:14567] = '{32'hc127b04a, 32'h42859550, 32'hc294a859, 32'h3f50d733, 32'hc12c72f0, 32'hc2af80e0, 32'h4269e3e3, 32'h42483565};
test_weights[14560:14567] = '{32'hc124cefd, 32'h4281f055, 32'h40172937, 32'h42af88f4, 32'hc1f1f3de, 32'hc253a29a, 32'hc207a6e6, 32'hc27914b9};
test_bias[1820:1820] = '{32'hc2b42f8b};
test_output[1820:1820] = '{32'h4580d31c};
test_input[14568:14575] = '{32'hc203f2e0, 32'hc037fddb, 32'hc0def26c, 32'h42a502bc, 32'hc262a0e5, 32'h4285e2a5, 32'h4294b1aa, 32'h4289c133};
test_weights[14568:14575] = '{32'hc29aa72a, 32'h41d29138, 32'h427b4b2d, 32'h422be055, 32'h3f3b2c2a, 32'hc21c8b6f, 32'hc1b93259, 32'hc23cca3e};
test_bias[1821:1821] = '{32'hc297c887};
test_output[1821:1821] = '{32'hc504e8a6};
test_input[14576:14583] = '{32'h41fb3b7b, 32'hc2a3a392, 32'hc2833b60, 32'h41586b20, 32'h42970043, 32'hc2909534, 32'hc2ae54e2, 32'hc21b49a7};
test_weights[14576:14583] = '{32'h4294a9e3, 32'h421a8eed, 32'h423a71c9, 32'h40b37724, 32'h42ba4c86, 32'hc2bf8d32, 32'h4225baf4, 32'hc1878d50};
test_bias[1822:1822] = '{32'h40a4a73b};
test_output[1822:1822] = '{32'h45e0f282};
test_input[14584:14591] = '{32'hc2a4b6f4, 32'h413989cc, 32'hc271eec4, 32'h42625bb2, 32'hc14d8884, 32'hc282353f, 32'h42b5186d, 32'hc19698b1};
test_weights[14584:14591] = '{32'h42a1af77, 32'h41c9b6c8, 32'h42af4e95, 32'hc2a5f8ee, 32'hc0421ab1, 32'hbf9ef267, 32'hc27082f4, 32'hc1ad957e};
test_bias[1823:1823] = '{32'h42c6d7e8};
test_output[1823:1823] = '{32'hc6a57826};
test_input[14592:14599] = '{32'h429915b4, 32'hc2bdb4fb, 32'h410760d6, 32'hc2849831, 32'hc215b642, 32'hc26d4892, 32'hc27c688f, 32'h3ffce6e0};
test_weights[14592:14599] = '{32'hc2ace10b, 32'hc1a11a06, 32'h42a4b903, 32'hc27451b6, 32'hc208f3c7, 32'h42676b27, 32'hc2b5cda9, 32'hc2180903};
test_bias[1824:1824] = '{32'hc167873f};
test_output[1824:1824] = '{32'h455d0214};
test_input[14600:14607] = '{32'hc2053982, 32'hc1dcb255, 32'hc1f9397e, 32'hc2ab004d, 32'h4298f784, 32'hc22902c8, 32'hc2c70486, 32'hc187b7e4};
test_weights[14600:14607] = '{32'hc2a788ff, 32'h429a4c7d, 32'hc29b08e6, 32'h42462617, 32'h42761f39, 32'h42b034e3, 32'h408cce39, 32'h42a8773c};
test_bias[1825:1825] = '{32'hc2b75729};
test_output[1825:1825] = '{32'hc5055f72};
test_input[14608:14615] = '{32'h42be29d8, 32'hc2085e5b, 32'hc0cba10c, 32'h42ac8693, 32'hc236f766, 32'h42383015, 32'hc2a80e80, 32'hc1e7ef03};
test_weights[14608:14615] = '{32'hc1853fd5, 32'h4235a7a4, 32'h41bec0fc, 32'hc23d9cc9, 32'hc29064d0, 32'h421f4f90, 32'h420e6e6d, 32'h41848859};
test_bias[1826:1826] = '{32'hc2856f94};
test_output[1826:1826] = '{32'hc5b47c4d};
test_input[14616:14623] = '{32'hc2b0f317, 32'hc281c9f6, 32'h4258a66e, 32'h42937f32, 32'h42b44343, 32'h42680430, 32'h41d2c3ab, 32'hc25124a0};
test_weights[14616:14623] = '{32'hc2c22a0c, 32'hc215ebef, 32'h41d641ad, 32'h42742949, 32'hc22fb5b0, 32'h418ab5ff, 32'hc2aedcd0, 32'hc20be230};
test_bias[1827:1827] = '{32'h42bb8756};
test_output[1827:1827] = '{32'h46551c6f};
test_input[14624:14631] = '{32'hc275936a, 32'h41a25b3e, 32'h4299e65d, 32'hc25a2751, 32'hc289f667, 32'h40d6aa2b, 32'h429702c4, 32'hc23bd719};
test_weights[14624:14631] = '{32'hc1442101, 32'h42732aad, 32'hc288dbf3, 32'hc1651532, 32'h42940855, 32'hc251fdf5, 32'hc29d27ae, 32'h41cc495a};
test_bias[1828:1828] = '{32'h41fd4ee8};
test_output[1828:1828] = '{32'hc66b43a4};
test_input[14632:14639] = '{32'h412a50cc, 32'hc1eb3c4a, 32'hc2aa159b, 32'hc29622f2, 32'h42969ec9, 32'h4207b520, 32'hc2137eba, 32'hc0064b09};
test_weights[14632:14639] = '{32'h4139734e, 32'h4291eb09, 32'hc2b9b3e1, 32'hc28dba18, 32'h428f29cf, 32'hc206cba6, 32'h42c4c31c, 32'h3e764459};
test_bias[1829:1829] = '{32'hc0c1e49d};
test_output[1829:1829] = '{32'h46387ce0};
test_input[14640:14647] = '{32'h42c2c3b9, 32'hc1e81366, 32'hc15506bd, 32'hc1d81d2d, 32'h42b022e7, 32'h4237e326, 32'h413bdc49, 32'hc26417e5};
test_weights[14640:14647] = '{32'hc20d94c2, 32'hc227d611, 32'hc1a144a1, 32'h420ea060, 32'hc29b0452, 32'hc2c610b7, 32'hc18fc6bd, 32'hc2a6e85b};
test_bias[1830:1830] = '{32'h428894ce};
test_output[1830:1830] = '{32'hc6175c9c};
test_input[14648:14655] = '{32'hc29b9cd7, 32'hc1a18945, 32'hc1a85fb4, 32'h41f66471, 32'h42c53001, 32'h41e16a11, 32'hc1d98a16, 32'hc20d578f};
test_weights[14648:14655] = '{32'h40baf340, 32'h4248e617, 32'hc0505fdf, 32'hc2a3a926, 32'hc21391da, 32'h429fcf62, 32'h42c38ea3, 32'h425149ab};
test_bias[1831:1831] = '{32'hc21b5c70};
test_output[1831:1831] = '{32'hc619f376};
test_input[14656:14663] = '{32'h42010026, 32'hc2822bf4, 32'h41ab8cca, 32'hc1832dbb, 32'h4196f68c, 32'hc226faae, 32'hc1d6210e, 32'h4289c194};
test_weights[14656:14663] = '{32'h42afa6ba, 32'h414e2316, 32'h3f787191, 32'h421bb7d2, 32'h42971752, 32'h421da7b2, 32'h420d3ba0, 32'hc2a5981c};
test_bias[1832:1832] = '{32'hc2af6258};
test_output[1832:1832] = '{32'hc5ae58b0};
test_input[14664:14671] = '{32'hc1ebb7ea, 32'h428e089a, 32'h42395e33, 32'h426a5c49, 32'hc2b1d211, 32'h42c68a9e, 32'h429b4e0f, 32'h42992ee2};
test_weights[14664:14671] = '{32'h40d3b1d3, 32'h425488d5, 32'h4202fdb9, 32'hc0fc2fd2, 32'hc2604ea5, 32'h425ed2d0, 32'h4224aacb, 32'hc296bac6};
test_bias[1833:1833] = '{32'hc1a47b1b};
test_output[1833:1833] = '{32'h464427ab};
test_input[14672:14679] = '{32'hc2541e78, 32'h42155170, 32'h41de7d25, 32'h42a62aa6, 32'h40c94ee1, 32'h4218d288, 32'hc29ebce8, 32'hc2b2056b};
test_weights[14672:14679] = '{32'hc2a99211, 32'h421d7e42, 32'hc18d3cef, 32'h42946953, 32'hc1e131c1, 32'h4241f118, 32'h4264e97f, 32'h429fae7d};
test_bias[1834:1834] = '{32'h4180e406};
test_output[1834:1834] = '{32'h44d25a68};
test_input[14680:14687] = '{32'h427354f5, 32'hc2614f79, 32'h411a3f44, 32'hc2617e85, 32'h42b1cc27, 32'hc2693f3f, 32'h42aa9de9, 32'hc28538f4};
test_weights[14680:14687] = '{32'hbe7af287, 32'h4215ad57, 32'h42822986, 32'h41d6836a, 32'h42a8f374, 32'h40da96f8, 32'h4286e8ef, 32'h415a8dbe};
test_bias[1835:1835] = '{32'h4226e8b0};
test_output[1835:1835] = '{32'h460c7ba8};
test_input[14688:14695] = '{32'hc2882622, 32'hc22487f8, 32'hc21c6b6c, 32'h41d78f85, 32'h4205f2f5, 32'hc2b5be8b, 32'h4239e127, 32'hc2534488};
test_weights[14688:14695] = '{32'h422e82f7, 32'h420e02ca, 32'hc15f61d9, 32'hc1af2351, 32'h428ca0e2, 32'hc2414ed3, 32'hc2af4b3a, 32'hc21863b2};
test_bias[1836:1836] = '{32'h42171c2b};
test_output[1836:1836] = '{32'h437906f8};
test_input[14696:14703] = '{32'h428dcc82, 32'hc26062f9, 32'hc1d57ce2, 32'h428149f7, 32'hc2b76267, 32'h424cca1d, 32'h4151bada, 32'hc2afb053};
test_weights[14696:14703] = '{32'hc2bcff31, 32'h429ecfa9, 32'hc2aab4cd, 32'hc258ab5b, 32'h426c3c50, 32'hc192d46b, 32'h42c376eb, 32'h429ab815};
test_bias[1837:1837] = '{32'h418627f6};
test_output[1837:1837] = '{32'hc6bd4d9c};
test_input[14704:14711] = '{32'h42b35e5c, 32'h41deae4e, 32'hc0001510, 32'hc238f827, 32'h421f03d8, 32'h42a7942d, 32'hc12d648b, 32'h4280dcc4};
test_weights[14704:14711] = '{32'h42307ad3, 32'hc18980fb, 32'h41f8c304, 32'h429ab510, 32'h424156dd, 32'hc1976e20, 32'h42b04164, 32'h428f6781};
test_bias[1838:1838] = '{32'h42433535};
test_output[1838:1838] = '{32'h45730443};
test_input[14712:14719] = '{32'h3f3f2e6d, 32'hc0f4f760, 32'h427cfa1b, 32'hc1c85bbf, 32'hc206e976, 32'h422caba0, 32'h42612dbb, 32'h429fb18a};
test_weights[14712:14719] = '{32'h4143140c, 32'hc2c761c5, 32'hc1074d8d, 32'hc1326856, 32'hc2c69094, 32'h42392973, 32'hc2503c8f, 32'hc1f81e93};
test_bias[1839:1839] = '{32'h42451ab7};
test_output[1839:1839] = '{32'h43fcdd0f};
test_input[14720:14727] = '{32'h42869033, 32'h42155a8e, 32'h41fce7d5, 32'h419744f6, 32'hc1cf3e47, 32'hc2624879, 32'hc26d1e7b, 32'h42bedb55};
test_weights[14720:14727] = '{32'hc0d9b884, 32'h41629198, 32'h4280d7a9, 32'h4255fed7, 32'hc2c18346, 32'hc26dde46, 32'h4180e916, 32'hc12e4261};
test_bias[1840:1840] = '{32'h42a23b7e};
test_output[1840:1840] = '{32'h45dd2256};
test_input[14728:14735] = '{32'h42a5f773, 32'hc2344507, 32'hc2949109, 32'h422ae5c7, 32'hc28d30d9, 32'hc2ace8af, 32'h42bbc096, 32'h41bb1f8c};
test_weights[14728:14735] = '{32'hc2277154, 32'h42ac1eaa, 32'hc1011fea, 32'h41e06885, 32'hc00a0793, 32'h41472929, 32'hc1e9b465, 32'h4213eed7};
test_bias[1841:1841] = '{32'hc0a453da};
test_output[1841:1841] = '{32'hc602a2ac};
test_input[14736:14743] = '{32'h423270a5, 32'hc1f552d9, 32'hc1921635, 32'h4262cdf4, 32'hc24d7c68, 32'hbf57965c, 32'h41a285f8, 32'h429dbfab};
test_weights[14736:14743] = '{32'hc22e699e, 32'h42b9d596, 32'hc2316c92, 32'hc28dcd31, 32'hc2a00e58, 32'h429b8890, 32'h41a74dd0, 32'h41a0d285};
test_bias[1842:1842] = '{32'h42186c30};
test_output[1842:1842] = '{32'hc4eecddd};
test_input[14744:14751] = '{32'h418074dd, 32'hc192e3ba, 32'hc21e9731, 32'hc2bea1d6, 32'h42c29d7a, 32'h416220dd, 32'hc215d8bc, 32'hc2752869};
test_weights[14744:14751] = '{32'hc29221c2, 32'h42bb761f, 32'hc1e77e56, 32'h429a7c6b, 32'h4174291d, 32'h42b4b54a, 32'h40b62be6, 32'hc2c3a9f7};
test_bias[1843:1843] = '{32'h429ab6e8};
test_output[1843:1843] = '{32'hc3f3b402};
test_input[14752:14759] = '{32'hc20f6e14, 32'h42548ecf, 32'hc21e6b29, 32'h41fc4664, 32'hc23983af, 32'h4275bd84, 32'h426be848, 32'hc2c5db04};
test_weights[14752:14759] = '{32'hc1f9da79, 32'hc26128eb, 32'hc2837ed7, 32'h4223fd0d, 32'h4239a8a3, 32'hc1fb6ab4, 32'hc29d0034, 32'h42bad41a};
test_bias[1844:1844] = '{32'hc272c876};
test_output[1844:1844] = '{32'hc679d688};
test_input[14760:14767] = '{32'hc2178ad2, 32'h41ebb964, 32'h429b2e46, 32'hc2a049ac, 32'hc0cd27a8, 32'hc001b72e, 32'h41b244c7, 32'hc2648df8};
test_weights[14760:14767] = '{32'hc28602ba, 32'hc2af34fe, 32'hc2c04ef4, 32'hc2133da8, 32'hc2aee147, 32'h423b7aa5, 32'hc27b2aa7, 32'hc1050fd2};
test_bias[1845:1845] = '{32'hc2bec32d};
test_output[1845:1845] = '{32'hc59f98d7};
test_input[14768:14775] = '{32'hc18acfbf, 32'h425e2f51, 32'hc2988e89, 32'hc27fadb2, 32'h420aaef9, 32'hc25931b5, 32'h41d6e8c3, 32'h429c6b6f};
test_weights[14768:14775] = '{32'h4113cd72, 32'h427f85c5, 32'hc12c9c19, 32'hc288c49b, 32'hc2998e16, 32'hc1c06893, 32'h412dedbd, 32'hc1abbfa4};
test_bias[1846:1846] = '{32'h423516e7};
test_output[1846:1846] = '{32'h45b7e209};
test_input[14776:14783] = '{32'h41a33a82, 32'h424bf734, 32'hbfe7c7e1, 32'hc2aafcdd, 32'h41bd2f96, 32'hbf8c20c8, 32'h42831cbf, 32'hc17d47af};
test_weights[14776:14783] = '{32'h42b260a8, 32'hc1dcbcb0, 32'hc15d429c, 32'hc290e0fc, 32'h42015e0f, 32'hc2970490, 32'hc238283d, 32'hc272e69b};
test_bias[1847:1847] = '{32'hc1e1b3e1};
test_output[1847:1847] = '{32'h45a88b00};
test_input[14784:14791] = '{32'h41816772, 32'h40b1fe65, 32'hc217e4f8, 32'h3ff3a659, 32'h41469806, 32'h41009232, 32'h41ae91c9, 32'hc2a14682};
test_weights[14784:14791] = '{32'hc12c8172, 32'h423db09b, 32'hc15c69a2, 32'h413df2ae, 32'hc282893f, 32'hc280f2d8, 32'h4155d1c2, 32'h42ac3142};
test_bias[1848:1848] = '{32'h4271f5a3};
test_output[1848:1848] = '{32'hc5e39ceb};
test_input[14792:14799] = '{32'hc229b782, 32'hc2b8724a, 32'h42b0fdbf, 32'h42513d9f, 32'h428e92f5, 32'hc2a74c0e, 32'hc21241d6, 32'hc2ba7251};
test_weights[14792:14799] = '{32'hc2c00eec, 32'h408e88f9, 32'h426d5a3e, 32'hc20c488e, 32'h42ab8ea8, 32'h41a064fe, 32'hc242114b, 32'hc1a70681};
test_bias[1849:1849] = '{32'h4211ad39};
test_output[1849:1849] = '{32'h466eab35};
test_input[14800:14807] = '{32'hbfc8c475, 32'hc2ad2620, 32'hc2ba49a8, 32'hc21bc8fa, 32'h429d85be, 32'hbd8891a6, 32'hc263d133, 32'hc14e9e08};
test_weights[14800:14807] = '{32'h41b3ca12, 32'h423a49b0, 32'h42a9e3b5, 32'h3ff81976, 32'hc1aaa72f, 32'hc13b9cec, 32'hc2881bc7, 32'h422f3d58};
test_bias[1850:1850] = '{32'hc2666229};
test_output[1850:1850] = '{32'hc623c5c5};
test_input[14808:14815] = '{32'hc1194e51, 32'h429538d8, 32'h4224c736, 32'h4256c604, 32'hc07f200f, 32'h4299df8a, 32'hc2345844, 32'hbfc04749};
test_weights[14808:14815] = '{32'hc0cb62ff, 32'hc03bcff9, 32'hc2997842, 32'hc1e0704b, 32'h42472784, 32'hc21e14d7, 32'h42b9f66d, 32'hc2b2061d};
test_bias[1851:1851] = '{32'h422a6300};
test_output[1851:1851] = '{32'hc63cc17a};
test_input[14816:14823] = '{32'h429bfe6b, 32'h412c1e24, 32'h428f2ae1, 32'hc2717725, 32'hc288e85e, 32'h417d79d3, 32'h42853579, 32'h41034ff8};
test_weights[14816:14823] = '{32'hc250c3bc, 32'h4125c20a, 32'hc222ef49, 32'hc2912a23, 32'h4278c12d, 32'hc224160c, 32'hc19d9259, 32'hc2c3cba7};
test_bias[1852:1852] = '{32'hc2be705e};
test_output[1852:1852] = '{32'hc6162c70};
test_input[14824:14831] = '{32'hc156aab4, 32'hc29314a5, 32'hc2aa4aa5, 32'hc2990ddf, 32'hc298a750, 32'hc2b33161, 32'h42086f23, 32'hc2698367};
test_weights[14824:14831] = '{32'h3e518219, 32'hc27c0e3e, 32'h42553bca, 32'hc2b1fe7c, 32'hc2022eec, 32'hc2b6065f, 32'h3e15ac56, 32'hc20db1fd};
test_bias[1853:1853] = '{32'h42b6d0e7};
test_output[1853:1853] = '{32'h4699f3cf};
test_input[14832:14839] = '{32'hc2616fe2, 32'hc2842d32, 32'hc101af2e, 32'hc22fadd9, 32'h40b6dadf, 32'h42b6554c, 32'hc2b425a2, 32'h41c9af9b};
test_weights[14832:14839] = '{32'hc2a541e8, 32'h429ca79b, 32'h4271de55, 32'h429d5f2a, 32'hc280a442, 32'h4218528f, 32'hc1310ed7, 32'h42b06c3f};
test_bias[1854:1854] = '{32'hc22f641a};
test_output[1854:1854] = '{32'h44e2eac8};
test_input[14840:14847] = '{32'hc2889016, 32'hc2973280, 32'h42a859ee, 32'hc13a564f, 32'h4299727a, 32'h4208bc57, 32'hbff56527, 32'hc2a4c24f};
test_weights[14840:14847] = '{32'h4224d908, 32'hc23aa4e0, 32'hc24e4273, 32'h41104b28, 32'h425b1096, 32'h41e06038, 32'h42732a7a, 32'h42acb7bd};
test_bias[1855:1855] = '{32'h42802201};
test_output[1855:1855] = '{32'hc5b350d3};
test_input[14848:14855] = '{32'h416e2fb9, 32'h411d2199, 32'hc1970b87, 32'hc18c5e79, 32'h405d2ebf, 32'hc182559d, 32'hc25ccc10, 32'h42844d49};
test_weights[14848:14855] = '{32'hc23462d7, 32'h420f8047, 32'h428312f5, 32'hc1fc2d7e, 32'hc1f3cc7c, 32'h427c527e, 32'hc2afba33, 32'h40d0a7d1};
test_bias[1856:1856] = '{32'hc2b06184};
test_output[1856:1856] = '{32'h453f0d67};
test_input[14856:14863] = '{32'h4274b9d2, 32'h41abb724, 32'hc24e39e0, 32'hc23f599b, 32'hc23f5f4c, 32'h42c5bd20, 32'hc0e24998, 32'hc215461e};
test_weights[14856:14863] = '{32'h429db823, 32'h4281aadb, 32'h42821f1a, 32'h414acb8d, 32'hc29350ca, 32'h41bc24db, 32'hc05cdfd4, 32'hc2c3e46b};
test_bias[1857:1857] = '{32'hc2a2b168};
test_output[1857:1857] = '{32'h4636dcdf};
test_input[14864:14871] = '{32'hc2868c15, 32'h3fcff064, 32'h42a30b4f, 32'h42a494d0, 32'hc28af44d, 32'h42200f0a, 32'h4227829d, 32'hc214ea5a};
test_weights[14864:14871] = '{32'hbfe21382, 32'hc1e48ac0, 32'hc1b28a21, 32'hc2ad97b4, 32'h429c5cc0, 32'h428d8a2a, 32'h429c1fa1, 32'hc28d194f};
test_bias[1858:1858] = '{32'hc26f2438};
test_output[1858:1858] = '{32'hc5b0adc6};
test_input[14872:14879] = '{32'hc15d0ff1, 32'hc212f0d2, 32'h4210c6b0, 32'h425745c0, 32'h42ae8bd7, 32'hc2b5818a, 32'h3fa46ab7, 32'hc1b65dcb};
test_weights[14872:14879] = '{32'hc2b04651, 32'h42471055, 32'h417c8561, 32'h4283d7bf, 32'h41ac8b02, 32'hbf03bf3a, 32'hc2426f95, 32'h426b4d00};
test_bias[1859:1859] = '{32'hc28e8252};
test_output[1859:1859] = '{32'h4577aeb1};
test_input[14880:14887] = '{32'hc2155e22, 32'h4127757f, 32'h41d9428c, 32'hc2886c01, 32'h40d88e21, 32'hc2a8e8d0, 32'hc2aff062, 32'h424038da};
test_weights[14880:14887] = '{32'h42ab3bfe, 32'hc29b8afe, 32'h423aeb40, 32'hc1106b4b, 32'hc298d2fb, 32'hc279d2c8, 32'h3fe7faee, 32'hc2aa5c2d};
test_bias[1860:1860] = '{32'hc2ab6c11};
test_output[1860:1860] = '{32'hc4d5686c};
test_input[14888:14895] = '{32'h42c7e202, 32'hc2bae2bc, 32'h420bd5ea, 32'h426843cd, 32'h426b8e50, 32'hc2530d1a, 32'h428525fc, 32'h41b6fc82};
test_weights[14888:14895] = '{32'hc27a528b, 32'h42192150, 32'hc2c2b5e7, 32'hc2b9deb4, 32'h418012b8, 32'h4206e55c, 32'hc19f68bd, 32'h42803f98};
test_bias[1861:1861] = '{32'hc28e1d8c};
test_output[1861:1861] = '{32'hc6978de2};
test_input[14896:14903] = '{32'hc16a9f23, 32'h41dfd873, 32'h4204a362, 32'hc25cce02, 32'hc263b9af, 32'hc1eea343, 32'hc2a09a02, 32'hc1c297d3};
test_weights[14896:14903] = '{32'h4285d69b, 32'hc2a88d8a, 32'hc101aa0e, 32'hc257180f, 32'hc2833929, 32'hc1300e3d, 32'hc2a22a66, 32'h419b8c59};
test_bias[1862:1862] = '{32'h42a76d7d};
test_output[1862:1862] = '{32'h46152665};
test_input[14904:14911] = '{32'h42c74669, 32'h42606efd, 32'h4141aa81, 32'h429bc954, 32'hc237720d, 32'hc2445271, 32'hc179c503, 32'hc2ad83fd};
test_weights[14904:14911] = '{32'h41289e98, 32'h42c32c2c, 32'hc1680249, 32'hc23554eb, 32'hc23bb7c4, 32'hc26908af, 32'h4234eb2e, 32'h4226cbbb};
test_bias[1863:1863] = '{32'h402a9fb8};
test_output[1863:1863] = '{32'h455b550f};
test_input[14912:14919] = '{32'h40d675bd, 32'h4214c7b1, 32'hc2a426a9, 32'hbeefd928, 32'h42213f3c, 32'hc1c3258f, 32'h4200330e, 32'hc297ecd0};
test_weights[14912:14919] = '{32'hc22e2ee2, 32'h424bc39a, 32'h41234ca8, 32'h420e71be, 32'h4056aa01, 32'h42826cbd, 32'hc25a753e, 32'hc180e6a5};
test_bias[1864:1864] = '{32'hbfb5b941};
test_output[1864:1864] = '{32'hc49a5aca};
test_input[14920:14927] = '{32'h4255f460, 32'hc285a84b, 32'hc2c05775, 32'hc1c0f6e0, 32'h42c41d97, 32'h40db88b9, 32'h4294e2bf, 32'h42058c15};
test_weights[14920:14927] = '{32'h42283ebf, 32'h4276559b, 32'hc11d5d54, 32'hc2812464, 32'h41aa46b1, 32'hc2c70ba0, 32'h415034b8, 32'h424eb61f};
test_bias[1865:1865] = '{32'h4271e9b8};
test_output[1865:1865] = '{32'h4595e402};
test_input[14928:14935] = '{32'hc1a4f7ae, 32'hc1c69eca, 32'h42274023, 32'hc1978ad9, 32'h4292e954, 32'h411752a1, 32'h408999c0, 32'hc17812ab};
test_weights[14928:14935] = '{32'h423f1cc0, 32'hc2520034, 32'h423f3677, 32'hc1b6ea1f, 32'hc1e167fa, 32'h424d1193, 32'h42875bf1, 32'h413c148b};
test_bias[1866:1866] = '{32'hc2929b62};
test_output[1866:1866] = '{32'h449618be};
test_input[14936:14943] = '{32'h4121ea13, 32'hc2ab48b3, 32'hc2a4dd8a, 32'hc1caab88, 32'h416ea84d, 32'h42bb460a, 32'h42ae1677, 32'h420d112d};
test_weights[14936:14943] = '{32'hc23559df, 32'hc2415207, 32'hc20d0b9b, 32'h42a4b7e1, 32'h4174d65a, 32'hc18b9cd0, 32'h41cf162a, 32'h41f91dd9};
test_bias[1867:1867] = '{32'hc290d34b};
test_output[1867:1867] = '{32'h45c72d08};
test_input[14944:14951] = '{32'h42b7e53a, 32'h42443493, 32'hc267a82d, 32'h4270c67a, 32'hc262c19b, 32'hc203a7b1, 32'hc1d1ad78, 32'h42541682};
test_weights[14944:14951] = '{32'h4221a53d, 32'hc2b764e2, 32'h42b31731, 32'h428b9602, 32'hc2a06c27, 32'h424cdbb1, 32'h4201e125, 32'h423d0962};
test_bias[1868:1868] = '{32'hc2a2d7fd};
test_output[1868:1868] = '{32'h4526bcb0};
test_input[14952:14959] = '{32'hc2093196, 32'h42894104, 32'hc21c1864, 32'hc21ba488, 32'hc18d401c, 32'h41e18ee4, 32'hc163ca86, 32'h42a0ba82};
test_weights[14952:14959] = '{32'hc1d4846c, 32'hc0c17534, 32'h4281b0bf, 32'hc2513ab5, 32'h428b371c, 32'hc2a084ff, 32'h4285aeb5, 32'h417858aa};
test_bias[1869:1869] = '{32'hc29f84ee};
test_output[1869:1869] = '{32'hc54cadd5};
test_input[14960:14967] = '{32'hc2054efb, 32'hc1d5d065, 32'hc297df14, 32'hc19bc348, 32'h3fec09fc, 32'hc2c5afb3, 32'h424df851, 32'h4248cc2b};
test_weights[14960:14967] = '{32'hc286a4bd, 32'hc28a4333, 32'h42533ffb, 32'hc246ab89, 32'h42983e1d, 32'hc2077271, 32'h4270866c, 32'h4292f74f};
test_bias[1870:1870] = '{32'h429cf1c8};
test_output[1870:1870] = '{32'h46321bc7};
test_input[14968:14975] = '{32'h423e5248, 32'h41fe06bc, 32'h42988c8a, 32'h41ebdac4, 32'h429e28b6, 32'hc1282262, 32'h42893e35, 32'hc2c473a2};
test_weights[14968:14975] = '{32'h4202c0a1, 32'h40cbdfc4, 32'h410cccfd, 32'h42a3506c, 32'hc27e6d2b, 32'h417647ca, 32'h42c6aafb, 32'hc296a760};
test_bias[1871:1871] = '{32'hc290960d};
test_output[1871:1871] = '{32'h46576ecf};
test_input[14976:14983] = '{32'hc28d3ab9, 32'hc255b02d, 32'h425134bc, 32'hc1b8b734, 32'hc1d3658c, 32'hc19174c8, 32'h42ba7056, 32'hc0b796fe};
test_weights[14976:14983] = '{32'h4214b96d, 32'hc2b9ff7b, 32'hc1bca5a2, 32'hc203bdc7, 32'h408e060e, 32'hc286bf4e, 32'hc1872d68, 32'h42b2d2f8};
test_bias[1872:1872] = '{32'hc06c03f8};
test_output[1872:1872] = '{32'h445d6db8};
test_input[14984:14991] = '{32'h4295dc24, 32'h40e4bbf7, 32'h42a83df2, 32'hc2558215, 32'hc1331769, 32'h4293471e, 32'h42a38bc6, 32'hc2c19ef2};
test_weights[14984:14991] = '{32'hc295034a, 32'hc28dfc29, 32'hc285dc2b, 32'h429639da, 32'hc25765b7, 32'h4209aa17, 32'h42292afd, 32'hc294f83b};
test_bias[1873:1873] = '{32'h41843e92};
test_output[1873:1873] = '{32'hc4ee5b34};
test_input[14992:14999] = '{32'hc085f53f, 32'h42318b4b, 32'h42c572c2, 32'hc2299462, 32'h42c57a52, 32'hc29c5faf, 32'h42324335, 32'hc16f9639};
test_weights[14992:14999] = '{32'h421a9ece, 32'h42c32800, 32'h42c22435, 32'hc2a0861c, 32'h429402c8, 32'hc1a3c595, 32'hc13748ab, 32'hc183f2e6};
test_bias[1874:1874] = '{32'hc2a71496};
test_output[1874:1874] = '{32'h46c8e7e8};
test_input[15000:15007] = '{32'h428d2d1d, 32'hc198b9aa, 32'hc1a3d285, 32'hc2247913, 32'h41c568fa, 32'h42b37358, 32'h42bc51d6, 32'h42affa4f};
test_weights[15000:15007] = '{32'hc2c55876, 32'hc209d2f4, 32'hc2557ae7, 32'hc289335e, 32'hc2aa5faf, 32'hc1b27d63, 32'h424bf55e, 32'hc237f0c8};
test_bias[1875:1875] = '{32'h423cc604};
test_output[1875:1875] = '{32'hc5b1fbff};
test_input[15008:15015] = '{32'h428c4a7b, 32'h4249b4d1, 32'h41d6da4b, 32'h4212dcc9, 32'h420c0d03, 32'h412843d3, 32'hc25b07b9, 32'h4295b786};
test_weights[15008:15015] = '{32'h42ab5966, 32'h4174d118, 32'h425b0478, 32'hc2653af8, 32'h42126be9, 32'hc1c581aa, 32'h4198e2f3, 32'hc24b64c6};
test_bias[1876:1876] = '{32'hc267bc0a};
test_output[1876:1876] = '{32'h450d2e30};
test_input[15016:15023] = '{32'h4165e7b4, 32'h42b9b2f1, 32'h4176292c, 32'h41d51997, 32'h419611d3, 32'hc251895c, 32'hc1d6673f, 32'hc2a70ec7};
test_weights[15016:15023] = '{32'hc2431d8b, 32'h4297c520, 32'h42044537, 32'h41d4e96b, 32'h4163723c, 32'h42050909, 32'hc2bf5081, 32'hc2892714};
test_bias[1877:1877] = '{32'h421c0da4};
test_output[1877:1877] = '{32'h46614768};
test_input[15024:15031] = '{32'h41fbee74, 32'hc20c2a83, 32'hc1ae41fd, 32'h42a5e4cb, 32'h42a7e51f, 32'hc2504eb3, 32'hc27adc2d, 32'hc19aa3da};
test_weights[15024:15031] = '{32'h42c54221, 32'hc19bb679, 32'h41d16fc2, 32'h42779aa5, 32'h42c520dc, 32'hc2b0c192, 32'h427d61f4, 32'h424dbcd3};
test_bias[1878:1878] = '{32'hc26f8d1f};
test_output[1878:1878] = '{32'h467d2867};
test_input[15032:15039] = '{32'h41fcbf2d, 32'hc1c032ac, 32'hc1ae5c9b, 32'hc1730e15, 32'hc24a83d8, 32'h41a53e38, 32'hc1c45b6c, 32'h41ff23a1};
test_weights[15032:15039] = '{32'h42a2572a, 32'hc28e5f1f, 32'h41298d57, 32'h428cca26, 32'h42932589, 32'hc240f828, 32'hc2ae098f, 32'h42993620};
test_bias[1879:1879] = '{32'h413de966};
test_output[1879:1879] = '{32'h4531bcb7};
test_input[15040:15047] = '{32'h42b1ebce, 32'hc19a8045, 32'h41448886, 32'hc21dc6f6, 32'h4000b5bf, 32'hc22da455, 32'h4250bdc0, 32'hc2b14586};
test_weights[15040:15047] = '{32'h42bed20a, 32'hc1890b39, 32'h3f1fb415, 32'h4250851e, 32'hc269c851, 32'hc22aab46, 32'h42706f90, 32'h41957631};
test_bias[1880:1880] = '{32'hc001ebfa};
test_output[1880:1880] = '{32'h461bfdfd};
test_input[15048:15055] = '{32'h4273f0c6, 32'h4243b445, 32'h42ae4510, 32'hc28fcae7, 32'hc2157c87, 32'hc231cfa7, 32'hc2a25be8, 32'h41f456a3};
test_weights[15048:15055] = '{32'hc2b0822c, 32'h42acc535, 32'h4056c32c, 32'hc29783f4, 32'h42c0f89f, 32'h41d179ba, 32'hc17496df, 32'hc1ad5c08};
test_bias[1881:1881] = '{32'h427a9236};
test_output[1881:1881] = '{32'h43e3ae23};
test_input[15056:15063] = '{32'h414b3b36, 32'hc26fe1d4, 32'hc2ac4d92, 32'hc10a1bc1, 32'h42c4ad72, 32'h423eecd1, 32'hc1c299da, 32'hbe99e47c};
test_weights[15056:15063] = '{32'h42a555f4, 32'hc2b07c0b, 32'h4271210f, 32'hc1eb365b, 32'h41ceb204, 32'hc1f22741, 32'hc21b0927, 32'hc20444ca};
test_bias[1882:1882] = '{32'hc28e9f3c};
test_output[1882:1882] = '{32'h45533c9a};
test_input[15064:15071] = '{32'h429f0429, 32'h42a11767, 32'hc222c178, 32'h41d1984a, 32'h4164e5f4, 32'h42c69c31, 32'hc2b7f240, 32'hc1c4a8f3};
test_weights[15064:15071] = '{32'hc246958c, 32'h42261088, 32'h41fea356, 32'hc266eb12, 32'hc184338c, 32'hc284f108, 32'hc20e709e, 32'hc2a33a8e};
test_bias[1883:1883] = '{32'h414eff5e};
test_output[1883:1883] = '{32'hc59ace98};
test_input[15072:15079] = '{32'h4290d8a1, 32'hc2984b9e, 32'h42b79432, 32'hc2a78579, 32'hc2ae2d1c, 32'h4296a4a5, 32'hc1c9d263, 32'hc266a52a};
test_weights[15072:15079] = '{32'hc2b19278, 32'hc20cf7fe, 32'hc2a1e961, 32'hc27980a2, 32'hc04d269f, 32'h428d23b8, 32'h423214a4, 32'hc2bae975};
test_bias[1884:1884] = '{32'hc2c5bc58};
test_output[1884:1884] = '{32'h456e08cb};
test_input[15080:15087] = '{32'hc2996d34, 32'h4248197f, 32'h429fce2b, 32'h425709e3, 32'hc2aaf2e3, 32'hbf957a2b, 32'hc2c63b2c, 32'h41a4e2fb};
test_weights[15080:15087] = '{32'h426770d8, 32'h42a974cd, 32'hc1b541ec, 32'hc23ee4f9, 32'hc2c642ed, 32'h429d80a2, 32'hc1c9059c, 32'hc25d1ad2};
test_bias[1885:1885] = '{32'h42912f6f};
test_output[1885:1885] = '{32'h45a36760};
test_input[15088:15095] = '{32'hc2c5e713, 32'hc268b481, 32'hc2838ecd, 32'h42726652, 32'hc2237b5d, 32'h422af3a8, 32'hc204af96, 32'h417d0b27};
test_weights[15088:15095] = '{32'hc20233df, 32'hc28061ef, 32'hc2bb4747, 32'hc2c79813, 32'hc1b71996, 32'hc00043c4, 32'h4292424a, 32'h426768b4};
test_bias[1886:1886] = '{32'hc160917e};
test_output[1886:1886] = '{32'h45c7c004};
test_input[15096:15103] = '{32'hc17b8a5b, 32'h40eef3a8, 32'hc24a3fa9, 32'h4292831e, 32'h42a1d5d4, 32'hc288f9fe, 32'h42b25e6f, 32'hc2881c35};
test_weights[15096:15103] = '{32'hbec6d6c5, 32'h41cc5446, 32'hc29b496d, 32'h4286d482, 32'hc1fe3733, 32'hc1ce33f3, 32'hc155765f, 32'hc19c3bcd};
test_bias[1887:1887] = '{32'hc214cb84};
test_output[1887:1887] = '{32'h460294e3};
test_input[15104:15111] = '{32'h41c069bf, 32'h42a674d9, 32'h429adb1e, 32'h4224e2bc, 32'hc26953c2, 32'hbe1a3c3d, 32'hc0eb8967, 32'h42b6e9cc};
test_weights[15104:15111] = '{32'h422d4755, 32'hc189c7ca, 32'hc0c95d97, 32'hc2119bad, 32'h42067277, 32'h42875e6c, 32'h41d4c810, 32'hc2b3d6db};
test_bias[1888:1888] = '{32'hc2c0dd2a};
test_output[1888:1888] = '{32'hc6490832};
test_input[15112:15119] = '{32'h41faabeb, 32'hbff8412d, 32'h428410dd, 32'hc0944f40, 32'hc208f272, 32'h42a66115, 32'hc2817487, 32'h429b52fd};
test_weights[15112:15119] = '{32'hc1cf8fbe, 32'hc2173c7e, 32'h428861f5, 32'hc24f0725, 32'hc1f19fda, 32'hc1b28f4e, 32'h419876fd, 32'hc2a66c5c};
test_bias[1889:1889] = '{32'hc27b15eb};
test_output[1889:1889] = '{32'hc58f12ec};
test_input[15120:15127] = '{32'h429f8183, 32'h41c0313c, 32'h41bcf168, 32'h421b4fa3, 32'hc2c0c8ec, 32'hc22f039a, 32'hc1125f5e, 32'h41f8e679};
test_weights[15120:15127] = '{32'hc209ee12, 32'h428b1b71, 32'h41f7adee, 32'h3e84b1b5, 32'hc1068559, 32'h408d35e3, 32'h401af1b7, 32'h41b1bfc1};
test_bias[1890:1890] = '{32'h42b07849};
test_output[1890:1890] = '{32'h44819b92};
test_input[15128:15135] = '{32'hc19f8ba7, 32'hc2447088, 32'hc2105648, 32'hc2b27e73, 32'hc21888fb, 32'h42b94439, 32'h412e3bc7, 32'hc280ae8d};
test_weights[15128:15135] = '{32'h42024686, 32'hc134c74e, 32'hc26800fa, 32'hc239a97e, 32'h40e09e92, 32'h42bf3e1b, 32'h42915372, 32'hc2b93036};
test_bias[1891:1891] = '{32'h42bc5ba1};
test_output[1891:1891] = '{32'h46a88b97};
test_input[15136:15143] = '{32'hc197bc1d, 32'hc0c0d125, 32'h41477c5f, 32'h4268f74d, 32'h42062f2a, 32'hc205a25f, 32'hc27a83ab, 32'h418b176d};
test_weights[15136:15143] = '{32'hc127694b, 32'h42960bc0, 32'hc2114879, 32'h3fa69a5e, 32'h41cfb2d4, 32'h420b2c31, 32'hc26878ca, 32'hc0bce8fd};
test_bias[1892:1892] = '{32'h4217eabf};
test_output[1892:1892] = '{32'h4525d17f};
test_input[15144:15151] = '{32'h4281cfe5, 32'hc2ab7f9c, 32'h42b85e0c, 32'h41bd7867, 32'hc1f64fc3, 32'h40f8fc43, 32'hc22409c4, 32'h42b9355a};
test_weights[15144:15151] = '{32'hc2970a5c, 32'hc1232755, 32'hc2b91ea0, 32'hc27d761b, 32'hc2c2768e, 32'h42a85433, 32'hc2375c8f, 32'hc149e63a};
test_bias[1893:1893] = '{32'h417b5ec6};
test_output[1893:1893] = '{32'hc61753ec};
test_input[15152:15159] = '{32'hc2c7eeed, 32'h42963117, 32'h426b758d, 32'hc28897e5, 32'hc2a66148, 32'hc24b7c2f, 32'hbf498525, 32'hc212ee39};
test_weights[15152:15159] = '{32'h4265837d, 32'h42b0f012, 32'h429befca, 32'h4180f5b3, 32'h41a7ef8d, 32'h41d01085, 32'h4283127c, 32'hc202942c};
test_bias[1894:1894] = '{32'hc174d3b0};
test_output[1894:1894] = '{32'h4519b38c};
test_input[15160:15167] = '{32'hc2aa74d0, 32'h428bb6d7, 32'hc2ad70d2, 32'hc0f4edb7, 32'h42b6ff51, 32'h4281533d, 32'h423acc07, 32'hc2bab486};
test_weights[15160:15167] = '{32'h42346bc8, 32'h4120880b, 32'hc1c74e1a, 32'hc2115b65, 32'hc1e7042c, 32'h42296b7e, 32'h4299f6ff, 32'h4182b0bc};
test_bias[1895:1895] = '{32'hc230c007};
test_output[1895:1895] = '{32'h44b13476};
test_input[15168:15175] = '{32'h41e1dd6f, 32'hc192ebf9, 32'hc23eccaf, 32'h42919f59, 32'hc28af779, 32'hc2b7c293, 32'h429984b2, 32'h41c3d41b};
test_weights[15168:15175] = '{32'h40f6e25c, 32'h42831823, 32'hc2219748, 32'hc29c18c2, 32'hc138d974, 32'hc2689b14, 32'hc1d54ad5, 32'hc1931cae};
test_bias[1896:1896] = '{32'hc2afa2e6};
test_output[1896:1896] = '{32'hc4939208};
test_input[15176:15183] = '{32'h429addbb, 32'h429dc1b0, 32'hc2bcd08b, 32'hc2b4e847, 32'hc28ff3c7, 32'hc2ac28c3, 32'hc13969dd, 32'hc2aaa6cd};
test_weights[15176:15183] = '{32'hc2af2767, 32'h42b89819, 32'h42b61a71, 32'hc206e33c, 32'h40ed797a, 32'h4212519b, 32'hc20bbf6d, 32'hc2464534};
test_bias[1897:1897] = '{32'hc2c533de};
test_output[1897:1897] = '{32'hc5831054};
test_input[15184:15191] = '{32'h42ae0593, 32'h42116099, 32'hc236efdf, 32'hc1e94877, 32'h41e94432, 32'h424caba3, 32'hc2aea8e4, 32'h424e28a6};
test_weights[15184:15191] = '{32'hc1d80d0e, 32'h428f8939, 32'h42188725, 32'h427fe4d5, 32'h413bf422, 32'hc11b9a22, 32'h423e8b35, 32'hc213724e};
test_bias[1898:1898] = '{32'h4117f54c};
test_output[1898:1898] = '{32'hc6155188};
test_input[15192:15199] = '{32'h42b584d8, 32'hc2c0f5f7, 32'h42bf5587, 32'h3f98dd9e, 32'hc2be49a6, 32'h417bcc5a, 32'hc11707b3, 32'h429c62fd};
test_weights[15192:15199] = '{32'hc20ca68f, 32'hc03e79e6, 32'hc23e3350, 32'h414b20a5, 32'h42973008, 32'hc1bada65, 32'hbefd563e, 32'hc2b9ce49};
test_bias[1899:1899] = '{32'h40402cd5};
test_output[1899:1899] = '{32'hc6addd2e};
test_input[15200:15207] = '{32'h41ed4e96, 32'hc2a3de01, 32'h4240591c, 32'hc2171df8, 32'h42575aad, 32'hc14690f9, 32'hc22c29ce, 32'hc0ec6049};
test_weights[15200:15207] = '{32'h42aa48be, 32'h42a160c3, 32'hc2810966, 32'hc1a4ac17, 32'h42ae0ed0, 32'h41cde48f, 32'hc24adba3, 32'hc2c75ad8};
test_bias[1900:1900] = '{32'hc26d8371};
test_output[1900:1900] = '{32'h444bdbb6};
test_input[15208:15215] = '{32'hc206918e, 32'h423221d2, 32'hc23437e5, 32'h41eeb84b, 32'hc2914dda, 32'h42729c21, 32'h4223306b, 32'h3f9c7e02};
test_weights[15208:15215] = '{32'h4271b82a, 32'h421cf67d, 32'hc2581a43, 32'h40b4d7b1, 32'hc2c41616, 32'h41a20c1b, 32'h42b648c9, 32'hc254df56};
test_bias[1901:1901] = '{32'hc260f502};
test_output[1901:1901] = '{32'h465ee7a6};
test_input[15216:15223] = '{32'h42b0fccd, 32'h41ba8bdd, 32'h42ae7159, 32'hc2279a2d, 32'hc2070cb8, 32'h42c79a8d, 32'hc2c1dba6, 32'hc2a7d92b};
test_weights[15216:15223] = '{32'h418b33cf, 32'h41c8ff2b, 32'hc2b80bb0, 32'hc1c53bcf, 32'hc2476a5d, 32'hc2896a9b, 32'hc29b8f12, 32'hc1f94102};
test_bias[1902:1902] = '{32'h42a4024a};
test_output[1902:1902] = '{32'h434237a1};
test_input[15224:15231] = '{32'h429ef916, 32'hc29b42c8, 32'h4203bc37, 32'h41158aa3, 32'hc22d8cfd, 32'hc1f26b6c, 32'hc2ad49ac, 32'h426fe091};
test_weights[15224:15231] = '{32'hc19bedc9, 32'hc29d321b, 32'h4154cce8, 32'hc07ebb1a, 32'h4210cc05, 32'hc17c9ed5, 32'h40ce7f5c, 32'h42994eb2};
test_bias[1903:1903] = '{32'h41587e75};
test_output[1903:1903] = '{32'h45f741fa};
test_input[15232:15239] = '{32'h41e05f7b, 32'h42438420, 32'h41e0800b, 32'h41fecff5, 32'h42320a95, 32'hc16d9cb8, 32'hc186c9c0, 32'hc2b72f58};
test_weights[15232:15239] = '{32'hc1f1f4fe, 32'hc2c7bdc2, 32'h4262f423, 32'h42c69731, 32'hc2b666a7, 32'h42c1e97b, 32'h42199778, 32'hc26a7ad9};
test_bias[1904:1904] = '{32'h4299ba44};
test_output[1904:1904] = '{32'hc4d16287};
test_input[15240:15247] = '{32'h429bcc83, 32'h4134c955, 32'h4120d51b, 32'hc1d21ba3, 32'hc228f6c3, 32'hc262f9fa, 32'h42af5bf6, 32'hc29b44fb};
test_weights[15240:15247] = '{32'hc233b1f4, 32'hc22e005a, 32'h41debc16, 32'hc2a6d513, 32'h4297f485, 32'hc1cf53b9, 32'h4272545d, 32'hc2183904};
test_bias[1905:1905] = '{32'h4195b460};
test_output[1905:1905] = '{32'h459d0e84};
test_input[15248:15255] = '{32'hc26b9cf3, 32'h4202d957, 32'hc28b8813, 32'h426c275b, 32'hc1aed10d, 32'h428544a6, 32'hc08c33c1, 32'h417178df};
test_weights[15248:15255] = '{32'h42154c6e, 32'hc1901bfd, 32'h41a54fcb, 32'hc28deafb, 32'h41c3649a, 32'h421fe754, 32'h41e70e4a, 32'hc1f8ff62};
test_bias[1906:1906] = '{32'hc28af3a1};
test_output[1906:1906] = '{32'hc5d953b7};
test_input[15256:15263] = '{32'hc248bc55, 32'hc15c92a5, 32'hc1af1ce0, 32'h42b935e1, 32'hc26d6c05, 32'h41058b52, 32'hbfdd7d14, 32'hc21ce941};
test_weights[15256:15263] = '{32'hc1044295, 32'h42942a40, 32'h42ab5902, 32'hc2a33472, 32'hc2341db0, 32'h417f06db, 32'h40d8ef34, 32'hc2834a41};
test_bias[1907:1907] = '{32'h427a56ef};
test_output[1907:1907] = '{32'hc58ff6f9};
test_input[15264:15271] = '{32'h429efffb, 32'hc2a8d9ac, 32'h419213e2, 32'hc2318aa0, 32'h427cffd1, 32'h42961212, 32'hc2950d83, 32'hc1ceae56};
test_weights[15264:15271] = '{32'h408df63c, 32'h41c29c0e, 32'hc25ff440, 32'h42aa85f8, 32'hc2c28754, 32'hc2b91ec0, 32'hc2a1a231, 32'hc265e68b};
test_bias[1908:1908] = '{32'hbfc8d055};
test_output[1908:1908] = '{32'hc63d0ac3};
test_input[15272:15279] = '{32'h4162dd9b, 32'h42b6d616, 32'h428ebaf6, 32'h423bc842, 32'h429f4794, 32'h42a2b818, 32'h41d00f84, 32'hc1862be1};
test_weights[15272:15279] = '{32'hc280c16b, 32'h418bbb6a, 32'hc139fc1e, 32'hc1904f41, 32'h413e5e26, 32'hc2ac4e4f, 32'hc2c495d3, 32'hc27ea347};
test_bias[1909:1909] = '{32'h4286af3d};
test_output[1909:1909] = '{32'hc6046e76};
test_input[15280:15287] = '{32'h4223e1d6, 32'hc1bf9e36, 32'hc08d717f, 32'hc2bdb9c4, 32'h415b9c7c, 32'hc209ec99, 32'h429eae3d, 32'hc1ef61f7};
test_weights[15280:15287] = '{32'h4229e983, 32'hc2947895, 32'h40dae5ea, 32'hc2603998, 32'hc23496a5, 32'h40bb6cb9, 32'hc1c75693, 32'h420c03e7};
test_bias[1910:1910] = '{32'hc004cced};
test_output[1910:1910] = '{32'h459aee78};
test_input[15288:15295] = '{32'hc08a39cf, 32'h42820761, 32'hc1a117ed, 32'h42592fde, 32'hc23478ed, 32'hc273fd4d, 32'h42a789c4, 32'hc22368af};
test_weights[15288:15295] = '{32'h42946c0e, 32'hc21bea43, 32'h4202346e, 32'hc220811b, 32'hc1aa2fd7, 32'hc244b8ab, 32'h4271cd6d, 32'hc26cb505};
test_bias[1911:1911] = '{32'hc2c2f8e9};
test_output[1911:1911] = '{32'h45b0b54f};
test_input[15296:15303] = '{32'h41de4a87, 32'hc2857991, 32'h4286d14d, 32'h42536612, 32'h42af37d6, 32'h421a09c5, 32'hc21d0ee3, 32'hc2a34915};
test_weights[15296:15303] = '{32'h42b4557c, 32'hc29769ec, 32'h41a4ccc6, 32'h3ed099ae, 32'h42a25d9a, 32'h421a19e2, 32'h42bcda09, 32'h42c15cef};
test_bias[1912:1912] = '{32'hc0e6648f};
test_output[1912:1912] = '{32'h45ba1ee0};
test_input[15304:15311] = '{32'h410029ea, 32'hc2998f2c, 32'hc1f55f27, 32'h409c7f9f, 32'h4248e9a0, 32'h411f1e56, 32'h425c070a, 32'hc231f494};
test_weights[15304:15311] = '{32'h4238f1f4, 32'hc228e706, 32'hc17e371c, 32'hc251bb60, 32'hc1ef2d94, 32'hc2144736, 32'hc2a5a701, 32'hc2a71dc9};
test_bias[1913:1913] = '{32'h404aef46};
test_output[1913:1913] = '{32'h448e31c7};
test_input[15312:15319] = '{32'h417d6053, 32'h4117ffdf, 32'hc281707a, 32'hc28a236b, 32'h42850116, 32'h40c1dc6e, 32'hc13ecfbc, 32'h42660d19};
test_weights[15312:15319] = '{32'h41a6b285, 32'h42a30937, 32'hc00eb79a, 32'h42321845, 32'hc28427a7, 32'hc22f6299, 32'hc10eafa9, 32'h421eabbf};
test_bias[1914:1914] = '{32'h425cf52a};
test_output[1914:1914] = '{32'hc57cb6c2};
test_input[15320:15327] = '{32'hc09a649f, 32'h42bbebbb, 32'h4289d231, 32'hc1d51d6e, 32'h41ed9550, 32'hc28fd58e, 32'hc283bf84, 32'hbf36ba28};
test_weights[15320:15327] = '{32'hc17fee38, 32'hc1e5122d, 32'h414f7e75, 32'h4113342f, 32'h4088dfa7, 32'h4286a467, 32'h413ba20e, 32'h42c70af6};
test_bias[1915:1915] = '{32'h3fcd4c54};
test_output[1915:1915] = '{32'hc5eb0946};
test_input[15328:15335] = '{32'h42b1941a, 32'hc249ebe2, 32'h40fc2529, 32'hc2245887, 32'h426e19da, 32'h41091740, 32'hc2643c79, 32'hc2349930};
test_weights[15328:15335] = '{32'h429ef6ec, 32'hc1624270, 32'hc181f1e2, 32'h4109e29e, 32'hc1a27540, 32'h41ab28ea, 32'hc23b678e, 32'hc1babd00};
test_bias[1916:1916] = '{32'h40b8eecc};
test_output[1916:1916] = '{32'h461c31c1};
test_input[15336:15343] = '{32'h40eb023f, 32'h41a6e31d, 32'h42999322, 32'hc2a25544, 32'h419b8a06, 32'hc1d1ff1f, 32'hc11abeb8, 32'hc234d3ab};
test_weights[15336:15343] = '{32'hc1584142, 32'hc2aa8505, 32'hc250cad3, 32'hc23dba17, 32'h42b86885, 32'h429a1bb3, 32'hc1e9d3ed, 32'hc26bec48};
test_bias[1917:1917] = '{32'hc174af2d};
test_output[1917:1917] = '{32'h4426e6fd};
test_input[15344:15351] = '{32'h4233814e, 32'hc25cbe45, 32'hc2685ac0, 32'h42585cab, 32'hc2a9bf51, 32'hc119ef7a, 32'hc241bc66, 32'h414951d7};
test_weights[15344:15351] = '{32'h41558fc9, 32'h42510d5a, 32'h429f7aeb, 32'h42a840de, 32'h422c4472, 32'h429783d3, 32'h424d84f4, 32'h42c2c4bd};
test_bias[1918:1918] = '{32'h42304ab1};
test_output[1918:1918] = '{32'hc5f90f92};
test_input[15352:15359] = '{32'h4298f337, 32'hc25ab4f1, 32'hc27cfe3e, 32'h42c58cb2, 32'h40db0b7e, 32'hc2649d53, 32'hc239ee10, 32'h4271577a};
test_weights[15352:15359] = '{32'hc228f316, 32'h427da5e5, 32'h42a60c45, 32'hc2b2770a, 32'hc2210066, 32'h40207767, 32'h42840d31, 32'h41f56e1c};
test_bias[1919:1919] = '{32'h408588f4};
test_output[1919:1919] = '{32'hc6aef5f7};
test_input[15360:15367] = '{32'h426fcd48, 32'hc21a178b, 32'h42c49796, 32'hc2b064a5, 32'hbfa8b11f, 32'h41a875aa, 32'h41fe76af, 32'hc25afcb9};
test_weights[15360:15367] = '{32'h42b9a524, 32'hc289ad73, 32'h42b833f1, 32'hc2a27347, 32'hc2ad7a7d, 32'h42baf30a, 32'h428faffb, 32'hc2599fb0};
test_bias[1920:1920] = '{32'h42c5615b};
test_output[1920:1920] = '{32'h46f90d6e};
test_input[15368:15375] = '{32'h4196704b, 32'h424ac556, 32'h42529c95, 32'h423b235c, 32'hc036c96e, 32'hc1876359, 32'hc2aac0dc, 32'h42a6c92e};
test_weights[15368:15375] = '{32'h41694788, 32'hc1ca5dd6, 32'h42312094, 32'h42860167, 32'hc1b651bb, 32'hc231a665, 32'hc0744de7, 32'h419c5506};
test_bias[1921:1921] = '{32'h41d5e4e1};
test_output[1921:1921] = '{32'h45e2c8b4};
test_input[15376:15383] = '{32'hc21e0999, 32'h40e7125f, 32'h422d57b2, 32'h41743e9f, 32'h423da014, 32'hc26a98ac, 32'h42a6c18f, 32'hc2a4def7};
test_weights[15376:15383] = '{32'h42a5d054, 32'h42a180f2, 32'hc24d64ad, 32'h4261080b, 32'hc21b0623, 32'hc2b3f8cc, 32'hc28f4ceb, 32'hc22b5872};
test_bias[1922:1922] = '{32'h41d030b0};
test_output[1922:1922] = '{32'hc53db647};
test_input[15384:15391] = '{32'h4272ae72, 32'h42615684, 32'hc2b2dd72, 32'hc0a1ce5b, 32'hc2a05470, 32'h4294772c, 32'h42ac90cb, 32'hc18761b5};
test_weights[15384:15391] = '{32'h424fe4c0, 32'h425af410, 32'h42b936e5, 32'hc2979714, 32'h406fff89, 32'hc1862baf, 32'hc28b828c, 32'h425c08bb};
test_bias[1923:1923] = '{32'hc1ec1e87};
test_output[1923:1923] = '{32'hc61f2a69};
test_input[15392:15399] = '{32'hc0f10258, 32'hc2b1c5c2, 32'hc235dd1c, 32'hc2b2eaa0, 32'hc195ab51, 32'hc2a407e1, 32'h41ce58c9, 32'h4146a5ce};
test_weights[15392:15399] = '{32'h41bb2b62, 32'hc2b64b35, 32'h41a38629, 32'hc240ee36, 32'h40517669, 32'hc28ea688, 32'h41858ff8, 32'hc2807d5b};
test_bias[1924:1924] = '{32'h42aba3e5};
test_output[1924:1924] = '{32'h4683649f};
test_input[15400:15407] = '{32'hc28692ed, 32'h42b94474, 32'hc28bbb46, 32'hc29f32d5, 32'h4273c1c2, 32'hc23363e7, 32'hc2a1f925, 32'hc0bcee4e};
test_weights[15400:15407] = '{32'hc1e4a5f3, 32'hc2ac74e4, 32'h41a721b9, 32'h42b732b6, 32'hc21af311, 32'h4264881a, 32'h41fcb28d, 32'h424df984};
test_bias[1925:1925] = '{32'hc1e87bd3};
test_output[1925:1925] = '{32'hc6b0cae7};
test_input[15408:15415] = '{32'hbf5fa659, 32'h425f5ab7, 32'hc2bc998d, 32'h42444d2b, 32'h42c399c8, 32'h427d80d9, 32'hc2a3b8fd, 32'hc269aabf};
test_weights[15408:15415] = '{32'hc189ba7c, 32'hc28d24eb, 32'hc20c5626, 32'h42b754cd, 32'h40caa734, 32'hc2a5018f, 32'hc285d47f, 32'h41cd878b};
test_bias[1926:1926] = '{32'hc1b3136b};
test_output[1926:1926] = '{32'h4549a950};
test_input[15416:15423] = '{32'h4289d6a6, 32'hc2b0e84a, 32'hc1916dc9, 32'hc111b957, 32'hc0db2fb0, 32'h418dc216, 32'h4283a0b5, 32'hc100d6b4};
test_weights[15416:15423] = '{32'h419b86ad, 32'hc1628b82, 32'hc1f0dd8e, 32'h413ec135, 32'h41fbdc22, 32'hc1e530bb, 32'h42bb9465, 32'hc205260d};
test_bias[1927:1927] = '{32'hc2a2af3d};
test_output[1927:1927] = '{32'h46076c58};
test_input[15424:15431] = '{32'h42989a85, 32'h421abeac, 32'h4261f17c, 32'hc279137e, 32'hc19ba291, 32'h42373888, 32'hc254f1dc, 32'hc1dafe31};
test_weights[15424:15431] = '{32'h40d06eef, 32'h428d9c18, 32'h42c7ad9d, 32'h418052d8, 32'hc2163118, 32'h42c7c55a, 32'h4298e826, 32'h42a4da2f};
test_bias[1928:1928] = '{32'hc2c42754};
test_output[1928:1928] = '{32'h45d33096};
test_input[15432:15439] = '{32'hc283e7c2, 32'h42ae18f0, 32'hc2912720, 32'h41419238, 32'h412c6f78, 32'hc1075c2a, 32'h4160e285, 32'h42c7e7b6};
test_weights[15432:15439] = '{32'hc2b6ebc6, 32'hc2c60893, 32'hc2a9f554, 32'hc2a3c65c, 32'hbf943a29, 32'h41ba5d24, 32'hc24dbc5d, 32'h42ba0c4f};
test_bias[1929:1929] = '{32'hc25258ec};
test_output[1929:1929] = '{32'h462a59ff};
test_input[15440:15447] = '{32'h4253f7a9, 32'h429e2df3, 32'h419b81ff, 32'hc13a80ec, 32'hc1d4fb6c, 32'h4286e9cc, 32'h427a52c1, 32'hc28b4887};
test_weights[15440:15447] = '{32'hc2b589a7, 32'h42c650b2, 32'h42b8ef9e, 32'h42444632, 32'h419f2ee2, 32'hc2891cc0, 32'h41d923f2, 32'h428a5be9};
test_bias[1930:1930] = '{32'hc2bc979f};
test_output[1930:1930] = '{32'hc5806fb5};
test_input[15448:15455] = '{32'h425c235c, 32'h422876f4, 32'hc2715dc1, 32'h4246dda6, 32'h42874f42, 32'h41df62e9, 32'hc1d3d513, 32'h42add667};
test_weights[15448:15455] = '{32'hc2ba967b, 32'hc2c6543e, 32'hc19821da, 32'hc2ae83d9, 32'hc29457c5, 32'hc18de8b3, 32'hc23c187c, 32'hc20ab81a};
test_bias[1931:1931] = '{32'h4268d680};
test_output[1931:1931] = '{32'hc69a1b9c};
test_input[15456:15463] = '{32'hc1dae0b1, 32'h41561e37, 32'h42aa1bdd, 32'h42ae896b, 32'hc284155c, 32'hc223842d, 32'hc225aada, 32'h42798191};
test_weights[15456:15463] = '{32'h411a7911, 32'h4213452b, 32'h41066b75, 32'hc0d07b67, 32'hc2a516dc, 32'h4233a2e7, 32'h4130b748, 32'h4291f84d};
test_bias[1932:1932] = '{32'hc2c32beb};
test_output[1932:1932] = '{32'h45f99d17};
test_input[15464:15471] = '{32'hc286d2bd, 32'h42b3e237, 32'hc1f21dad, 32'hc1a2455e, 32'hc2b8a9dc, 32'hc2c74d79, 32'h428e9e54, 32'hc1acf4c2};
test_weights[15464:15471] = '{32'hc20c857b, 32'h4281138e, 32'hc13b08f2, 32'h422aa642, 32'hc2355d62, 32'hc0822f24, 32'hbff4751b, 32'hc26015a0};
test_bias[1933:1933] = '{32'hc28b7023};
test_output[1933:1933] = '{32'h464f2986};
test_input[15472:15479] = '{32'h428ccc6f, 32'h422c4169, 32'h429393e9, 32'h41f21dd5, 32'h42278b82, 32'hc159a1bb, 32'h413d09f0, 32'hc2bd2753};
test_weights[15472:15479] = '{32'hc22dff8d, 32'h418c576c, 32'h421b1e82, 32'h408e7d40, 32'hc18f1827, 32'h405ce77a, 32'h4213e5a9, 32'h42868a3d};
test_bias[1934:1934] = '{32'hc1906ba5};
test_output[1934:1934] = '{32'hc5bd112e};
test_input[15480:15487] = '{32'h41c26764, 32'h426b44d7, 32'hc2abd8d3, 32'h3f825a0d, 32'hc21efea7, 32'hc2836ede, 32'h42630785, 32'h429471c8};
test_weights[15480:15487] = '{32'h424c60fc, 32'h42b139d3, 32'hc1f509ca, 32'h417005f6, 32'h4296026f, 32'hc2966cd7, 32'h41ea70f9, 32'h3f884164};
test_bias[1935:1935] = '{32'hc2bee6fe};
test_output[1935:1935] = '{32'h46469399};
test_input[15488:15495] = '{32'h4298cb11, 32'h4287a18b, 32'hc2b2f649, 32'hc195e56b, 32'h42909a46, 32'hc1bb7fad, 32'h42139d2d, 32'h41510e36};
test_weights[15488:15495] = '{32'h41ab077e, 32'hc10e3fb8, 32'h424f4cdd, 32'hc28f5946, 32'hc2bd3087, 32'h41f9102a, 32'hc2b2857f, 32'hc23c54af};
test_bias[1936:1936] = '{32'h41e7ba6c};
test_output[1936:1936] = '{32'hc6564537};
test_input[15496:15503] = '{32'hc2808d82, 32'hc2598358, 32'hc1253149, 32'h41e9e306, 32'h42c29161, 32'hc181ab2b, 32'hc1360b9a, 32'hc2b18416};
test_weights[15496:15503] = '{32'h4294ad34, 32'hc28ee55d, 32'hc09932f5, 32'hc2c6d279, 32'h42ae1678, 32'h428f928f, 32'hbff844ab, 32'h426951f1};
test_bias[1937:1937] = '{32'hc295109d};
test_output[1937:1937] = '{32'hc4d166f6};
test_input[15504:15511] = '{32'hc1f0891b, 32'hc275b451, 32'h42bae140, 32'h414b8936, 32'h4246691d, 32'hc2969b5b, 32'h4244c678, 32'h41f3bf40};
test_weights[15504:15511] = '{32'h418b2157, 32'hc23a5526, 32'h4284ade3, 32'h3f9799c6, 32'hc29c8927, 32'hc2564561, 32'hc2aee30b, 32'hc27a263b};
test_bias[1938:1938] = '{32'h42c3b962};
test_output[1938:1938] = '{32'h45222ab8};
test_input[15512:15519] = '{32'h42bd52c8, 32'hc255210a, 32'h424dcf48, 32'h42a564bb, 32'h4256ee2a, 32'h4182bcf5, 32'h4249625e, 32'hc08ae05e};
test_weights[15512:15519] = '{32'hc2c56a31, 32'h42049f32, 32'hc21d36ba, 32'h42159bb5, 32'hc249d8f2, 32'h42556e93, 32'hc26e8328, 32'hc0b37c53};
test_bias[1939:1939] = '{32'hc29970e1};
test_output[1939:1939] = '{32'hc669560a};
test_input[15520:15527] = '{32'hc1c7433a, 32'h4093c400, 32'hc23d9d71, 32'hc2b1f675, 32'h4283daa6, 32'hc22d1fca, 32'h4204e891, 32'hc14149dc};
test_weights[15520:15527] = '{32'h429ddc17, 32'hc2c60889, 32'h427db719, 32'h42c7e299, 32'hc298c52c, 32'hc2864040, 32'h41c8c88c, 32'hc0812574};
test_bias[1940:1940] = '{32'hc28f5e39};
test_output[1940:1940] = '{32'hc6746a46};
test_input[15528:15535] = '{32'h4223d770, 32'h429d57c7, 32'h41839a6a, 32'h428014b2, 32'h42bccc99, 32'h425d541b, 32'hc23e8ff7, 32'h42830c1c};
test_weights[15528:15535] = '{32'hc26e9327, 32'hc257f866, 32'h425cb857, 32'hc1d949e9, 32'hc23021df, 32'hc225affe, 32'h4296fc48, 32'h422dabae};
test_bias[1941:1941] = '{32'hc1c7c640};
test_output[1941:1941] = '{32'hc6666e99};
test_input[15536:15543] = '{32'hc174c156, 32'hc22a1c06, 32'h41d4d3d4, 32'h42948377, 32'h42a87e53, 32'hc2c071c7, 32'hc280407c, 32'hc278e784};
test_weights[15536:15543] = '{32'hc20bfd6a, 32'h41dac43d, 32'h41d2e8bd, 32'hc2584526, 32'h4298fff0, 32'h42845410, 32'hc24b7f10, 32'hc21c7440};
test_bias[1942:1942] = '{32'h422e99dc};
test_output[1942:1942] = '{32'h44eaa5d3};
test_input[15544:15551] = '{32'hc2aabdef, 32'hc1c35ab2, 32'hc255f991, 32'h3e996c6f, 32'hc28d0a43, 32'h42c25f98, 32'hc2a5490e, 32'hc1ce6030};
test_weights[15544:15551] = '{32'h425b4460, 32'hc12ab4f2, 32'hc0ff5ce1, 32'h4145db8d, 32'h41d7f069, 32'h4290ebed, 32'hc206098a, 32'hc2acf8d9};
test_bias[1943:1943] = '{32'hc1f37ec8};
test_output[1943:1943] = '{32'h45bf4032};
test_input[15552:15559] = '{32'h42b4c09b, 32'hc2363a3c, 32'hc0d1faef, 32'h42201263, 32'hc1ce7881, 32'h42c789bb, 32'h40c6aa7e, 32'hc2af7091};
test_weights[15552:15559] = '{32'h4293a002, 32'hbf0534ac, 32'h4247a00f, 32'hc25bff18, 32'h3f99f35d, 32'h4168247f, 32'h41b2ad78, 32'h42047ee2};
test_bias[1944:1944] = '{32'hc2c4247f};
test_output[1944:1944] = '{32'h4529da13};
test_input[15560:15567] = '{32'h3e42abe6, 32'hc247ec17, 32'hc19976de, 32'hc20cf64f, 32'hc22fbc09, 32'h41379e39, 32'h42c72e94, 32'h421800e3};
test_weights[15560:15567] = '{32'h429ab092, 32'hc2c15f64, 32'hc28a6014, 32'h4194f9cc, 32'h41b3d2d5, 32'hc22b820e, 32'hc2bf7366, 32'hc2b6e5e9};
test_bias[1945:1945] = '{32'h41bc199e};
test_output[1945:1945] = '{32'hc60bc9f9};
test_input[15568:15575] = '{32'hc2ad7334, 32'h425b4324, 32'h4158b82a, 32'hc281ce70, 32'h429f0996, 32'h428e1c59, 32'h42b0d655, 32'hc10328d3};
test_weights[15568:15575] = '{32'hc1d81d60, 32'h3f54ca49, 32'h42628b4b, 32'h42726c0f, 32'hc0b98ed9, 32'h40769b45, 32'h42bec029, 32'hc28685e0};
test_bias[1946:1946] = '{32'h42255971};
test_output[1946:1946] = '{32'h45fbe301};
test_input[15576:15583] = '{32'h426fba88, 32'h42515530, 32'h41eabe66, 32'hc240d6cf, 32'h41fd529c, 32'hc22e1c22, 32'hc2397b8a, 32'hc2a3827b};
test_weights[15576:15583] = '{32'h423befac, 32'hc12b9c89, 32'h420b4d10, 32'h4228f7fe, 32'h4251df19, 32'h42c2aed1, 32'h42bc64ee, 32'h40dc3926};
test_bias[1947:1947] = '{32'h4258a095};
test_output[1947:1947] = '{32'hc5c2211c};
test_input[15584:15591] = '{32'hc2c5704e, 32'h4030ac8e, 32'h412a4a85, 32'h40807d29, 32'hc2492dc8, 32'hc2868374, 32'h4238ec1c, 32'h426aefc9};
test_weights[15584:15591] = '{32'h4205e121, 32'hc29908b7, 32'hbfb04283, 32'hc2b35b14, 32'hc234ba26, 32'h42490162, 32'hc2a0a1e0, 32'hc2417909};
test_bias[1948:1948] = '{32'hc26394ab};
test_output[1948:1948] = '{32'hc63560fe};
test_input[15592:15599] = '{32'hc14709ff, 32'hc2728b93, 32'h425f0071, 32'h4277ddc4, 32'hc2c12ebe, 32'h42af4e2b, 32'h4202eecd, 32'h429066a8};
test_weights[15592:15599] = '{32'hc2b52a04, 32'h42a1026c, 32'h404f94c4, 32'hc2c08b11, 32'hc2bc02c6, 32'hc284f7e7, 32'h42840efa, 32'h42092b90};
test_bias[1949:1949] = '{32'hc234a526};
test_output[1949:1949] = '{32'hc4d3d830};
test_input[15600:15607] = '{32'h41c80169, 32'h42a62dab, 32'hc21a69ef, 32'h41c836d9, 32'h4201382d, 32'h42ab48a3, 32'hc24aeafd, 32'h42a04585};
test_weights[15600:15607] = '{32'hc1aee93c, 32'h41fffab6, 32'h42934ac8, 32'hc1d8f78f, 32'h429b171c, 32'h428a1039, 32'h4264016a, 32'hc0c2d5c0};
test_bias[1950:1950] = '{32'h42b90ad2};
test_output[1950:1950] = '{32'h4568854c};
test_input[15608:15615] = '{32'hc138ecba, 32'hc0920362, 32'hc1861b5c, 32'hc2a409f9, 32'h41b98c54, 32'hc2886208, 32'h402914cd, 32'hc261dd47};
test_weights[15608:15615] = '{32'hc1a663c5, 32'h4283f152, 32'h415e4281, 32'h42302d50, 32'hc0c479ad, 32'h42c5e1d8, 32'h405b9f35, 32'h42c3e0b5};
test_bias[1951:1951] = '{32'hc2b7f98b};
test_output[1951:1951] = '{32'hc68030f4};
test_input[15616:15623] = '{32'h4284e967, 32'hc2a151b1, 32'hc29392d9, 32'hc2c7d2ae, 32'h41c24767, 32'h41a9e16e, 32'hc1684e24, 32'hc2a4a9c2};
test_weights[15616:15623] = '{32'h41e59f88, 32'h42153cc6, 32'hc23f4301, 32'hc22dd11d, 32'h4196b229, 32'h4263a9e2, 32'h42bd2d5e, 32'h40e901f2};
test_bias[1952:1952] = '{32'hc28fb796};
test_output[1952:1952] = '{32'h45c7a9bb};
test_input[15624:15631] = '{32'h421e169a, 32'hc1be0f6c, 32'hc2a71629, 32'hc262f86d, 32'h40ae2ae4, 32'hc29ec143, 32'h415c9dd2, 32'h4247f03f};
test_weights[15624:15631] = '{32'hc2648df1, 32'hc11ca995, 32'h42b616f1, 32'h42a9deb8, 32'h42b81685, 32'h42a291df, 32'h42b74a2a, 32'hc211995b};
test_bias[1953:1953] = '{32'hc240c03b};
test_output[1953:1953] = '{32'hc6a41cd6};
test_input[15632:15639] = '{32'h4067b574, 32'h42a87b2b, 32'h42a71504, 32'hc29987a6, 32'hc299aebc, 32'hc294519f, 32'h4282ceec, 32'hc298c3e9};
test_weights[15632:15639] = '{32'h42b48ee3, 32'h42841364, 32'hc287b994, 32'h4185b3bd, 32'h41cbc349, 32'hc23affdb, 32'h42aaa811, 32'hc299ae91};
test_bias[1954:1954] = '{32'h4283bfa9};
test_output[1954:1954] = '{32'h463aedc4};
test_input[15640:15647] = '{32'h428537cb, 32'hc2b22c82, 32'h3ffd2cf1, 32'h42a55fb7, 32'h42b0a780, 32'h421cde62, 32'hc1b1c3e6, 32'h42964b0a};
test_weights[15640:15647] = '{32'h4237e771, 32'hc261a104, 32'h409f49e0, 32'h41e35e95, 32'h42338964, 32'h42415b51, 32'hc18e5a43, 32'hc18e5040};
test_bias[1955:1955] = '{32'hc28a7088};
test_output[1955:1955] = '{32'h466f0444};
test_input[15648:15655] = '{32'h427005e2, 32'hc1336c88, 32'hc2899327, 32'h422aa311, 32'h40914fb3, 32'h4281182f, 32'h42be86d9, 32'h40f3cd69};
test_weights[15648:15655] = '{32'h4299a496, 32'h428c19c6, 32'h428abbac, 32'h42497a83, 32'h42b78af4, 32'hc2329fb4, 32'h41286794, 32'h4258100b};
test_bias[1956:1956] = '{32'hc2281f85};
test_output[1956:1956] = '{32'h42d7b9d7};
test_input[15656:15663] = '{32'h40b0bb40, 32'hc2265439, 32'hc2add81f, 32'h425c61eb, 32'h4238ec2d, 32'h422c1258, 32'h4275a779, 32'hc2202315};
test_weights[15656:15663] = '{32'h428753ee, 32'hc266b60f, 32'hc2212e2c, 32'h41fd1b20, 32'h42213ab8, 32'h429397a0, 32'h426f8983, 32'hc0c7fc60};
test_bias[1957:1957] = '{32'hc1d62843};
test_output[1957:1957] = '{32'h468479b7};
test_input[15664:15671] = '{32'hc2bff101, 32'hc02cd30b, 32'hc1eb9fb6, 32'h40dc946b, 32'hc2b455d1, 32'hc2ace5f5, 32'hc1633945, 32'h4295b969};
test_weights[15664:15671] = '{32'hc1b687c5, 32'hc238a4d1, 32'h42be7f16, 32'h420c39eb, 32'h4128a662, 32'h42449eb2, 32'h42b7498f, 32'h42a2242a};
test_bias[1958:1958] = '{32'hc0362286};
test_output[1958:1958] = '{32'hc42b180f};
test_input[15672:15679] = '{32'h4183937e, 32'hc2875020, 32'hc28742b9, 32'hc24eaecc, 32'h4251b94f, 32'hc28640b8, 32'hc2b17da5, 32'hc25b5071};
test_weights[15672:15679] = '{32'h41a01235, 32'hc2bb3f60, 32'hc2962c74, 32'hc175c321, 32'h428e535f, 32'hc26fad68, 32'hc1f3359b, 32'hc20433b1};
test_bias[1959:1959] = '{32'h41c23ea3};
test_output[1959:1959] = '{32'h46c1eda3};
test_input[15680:15687] = '{32'hc2a1845d, 32'hc207f880, 32'hc1c34a68, 32'hc224f0c3, 32'h4288591e, 32'h4213f5d1, 32'h426ac21e, 32'h42b876ab};
test_weights[15680:15687] = '{32'h42c5b51b, 32'h41d278ec, 32'h41d097f8, 32'h414b9477, 32'h41d4bc09, 32'hc2898d63, 32'hc23eaed7, 32'hc204790c};
test_bias[1960:1960] = '{32'h4250a88b};
test_output[1960:1960] = '{32'hc681742e};
test_input[15688:15695] = '{32'h41c3dd25, 32'h419b64a3, 32'h41411e74, 32'h42c11721, 32'hc0d278a8, 32'h42a995dd, 32'h3f98bf20, 32'h418490ac};
test_weights[15688:15695] = '{32'hc0d772bd, 32'hc2a5a2fa, 32'h4239ac6f, 32'h4218d1b9, 32'hc2266aa8, 32'h421e58f1, 32'hc2377f30, 32'h42a08b2e};
test_bias[1961:1961] = '{32'hc2bca783};
test_output[1961:1961] = '{32'h45e3b52c};
test_input[15696:15703] = '{32'hc28026a0, 32'h40c18d2d, 32'hc1295b70, 32'h4292cec8, 32'h424b196f, 32'h41dcfa23, 32'hc29eed71, 32'hc1c0d965};
test_weights[15696:15703] = '{32'h42a44156, 32'h41e5d6af, 32'hc243bfe7, 32'hc257aa12, 32'h427e8b6e, 32'h417512e9, 32'hc09db41b, 32'h42b3ae73};
test_bias[1962:1962] = '{32'h3fbfdda1};
test_output[1962:1962] = '{32'hc5cfb519};
test_input[15704:15711] = '{32'h42a2e2bc, 32'hc25fd2e6, 32'hc28eedc1, 32'h4239fd4a, 32'h425b5fb3, 32'hc21a0e76, 32'h42180803, 32'hc12a13eb};
test_weights[15704:15711] = '{32'hc197c577, 32'hc289902e, 32'hc2041ce5, 32'hc28c96f0, 32'h42ac35fd, 32'h42a46329, 32'hc1a907a8, 32'hc1c05476};
test_bias[1963:1963] = '{32'h4213b22d};
test_output[1963:1963] = '{32'h4518998e};
test_input[15712:15719] = '{32'hc23c04eb, 32'hc0353ef9, 32'hc286d04d, 32'h41ee04c4, 32'hc2b22e8b, 32'hc2aca14f, 32'hc1922fba, 32'h41eb9218};
test_weights[15712:15719] = '{32'hc21f8d9b, 32'hc1776f47, 32'h42ab059c, 32'h40086256, 32'hc2aa8e3b, 32'hc22901df, 32'hc29163c3, 32'h4243ff93};
test_bias[1964:1964] = '{32'h42875290};
test_output[1964:1964] = '{32'h4620f5d2};
test_input[15720:15727] = '{32'hc2901eb1, 32'hc2bb4489, 32'hc28fd2cd, 32'h3f50c437, 32'hc1bf878c, 32'h409e32b1, 32'hc29325a8, 32'h42ba9633};
test_weights[15720:15727] = '{32'h42a585af, 32'h4281c3e2, 32'h4216889c, 32'h42a4a25e, 32'hc2b0f54c, 32'hc1bda5a8, 32'hc1854542, 32'hc23890b0};
test_bias[1965:1965] = '{32'h419f79be};
test_output[1965:1965] = '{32'hc675e076};
test_input[15728:15735] = '{32'h41a0823a, 32'h42c5258f, 32'h42ac8fab, 32'hc1d2592f, 32'h42c14c33, 32'h420b0dca, 32'hc1924622, 32'h421d42c4};
test_weights[15728:15735] = '{32'hc2943bf6, 32'h42132248, 32'h428547da, 32'hc21b49c0, 32'hc09475d5, 32'hc2878e7f, 32'hc20e075a, 32'hc1e554a6};
test_bias[1966:1966] = '{32'h429f44da};
test_output[1966:1966] = '{32'h45b254b2};
test_input[15736:15743] = '{32'hc2b6e26f, 32'h413de893, 32'h41ea0f53, 32'hc116b872, 32'h42a95de9, 32'h42c440b7, 32'hc288b93f, 32'h42547900};
test_weights[15736:15743] = '{32'hc1f89579, 32'hc214c4e4, 32'h425b0ca4, 32'hc2c06956, 32'h42a1699d, 32'h422cdb07, 32'hc20419f3, 32'h4204b673};
test_bias[1967:1967] = '{32'hc2baf7b7};
test_output[1967:1967] = '{32'h469b8bbc};
test_input[15744:15751] = '{32'h418cc099, 32'hc1f7afe1, 32'h42aa4367, 32'h428b3f26, 32'hc29c82d7, 32'h42b33f63, 32'hc2858f2a, 32'h41d2d0db};
test_weights[15744:15751] = '{32'h41d88583, 32'hc284df66, 32'hc28f26ab, 32'hc20f1b8c, 32'hc2b28f10, 32'h42bba29a, 32'h41ffa67c, 32'hc2b90f2b};
test_bias[1968:1968] = '{32'hc251f78c};
test_output[1968:1968] = '{32'h45937738};
test_input[15752:15759] = '{32'hc239d553, 32'h41dd35c5, 32'h403c5177, 32'hc2bdb952, 32'hc299c0a9, 32'h3f947efd, 32'hc29e529d, 32'h427cb331};
test_weights[15752:15759] = '{32'hc28be5cb, 32'hc2651113, 32'h40627387, 32'h42760059, 32'h42c0e01a, 32'h4203a605, 32'hc2959244, 32'hc2416eaa};
test_bias[1969:1969] = '{32'hc2221753};
test_output[1969:1969] = '{32'hc60811ae};
test_input[15760:15767] = '{32'hc237396f, 32'h40c61a3f, 32'hc2c06330, 32'h427c81b0, 32'h4195b137, 32'hc2c1f343, 32'hc253221f, 32'h42685ade};
test_weights[15760:15767] = '{32'h4226248e, 32'h41a855a2, 32'h429caa08, 32'hc21c1920, 32'hc1ae762d, 32'hc28971db, 32'h42018c4f, 32'hc2c23021};
test_bias[1970:1970] = '{32'hc2c08a5b};
test_output[1970:1970] = '{32'hc64a8195};
test_input[15768:15775] = '{32'hbfd7467f, 32'hc19b7c22, 32'hc2346b8d, 32'h4268f218, 32'h416dcc10, 32'hc15324d9, 32'hc06aa109, 32'h42c3f99a};
test_weights[15768:15775] = '{32'h41dd5cd8, 32'hc29a94a4, 32'h428558f3, 32'h42c3828e, 32'h42b52528, 32'h40838f71, 32'h4142c12f, 32'h4280f1f3};
test_bias[1971:1971] = '{32'h4282792c};
test_output[1971:1971] = '{32'h4637ecd6};
test_input[15776:15783] = '{32'h42999a71, 32'hc1bc23fd, 32'hc071980c, 32'h411cd50b, 32'hc2844d74, 32'hc192469a, 32'hc2768b8b, 32'hc25caefb};
test_weights[15776:15783] = '{32'hc1c6375b, 32'hc23dbdb8, 32'hc2afe6c8, 32'h41ca2fe2, 32'hc2aab82f, 32'hc2632a3a, 32'h428436fa, 32'h4225dd04};
test_bias[1972:1972] = '{32'hc28e4f31};
test_output[1972:1972] = '{32'h422fd7c0};
test_input[15784:15791] = '{32'h41e0cd24, 32'hc28cc053, 32'h41062850, 32'hc2a3b045, 32'hc0f0c577, 32'h4236d463, 32'hc2a7c72c, 32'h42792c9c};
test_weights[15784:15791] = '{32'hc287f909, 32'hc29c8030, 32'h3ff96449, 32'h42aa8bea, 32'h4235b900, 32'h41d11f5e, 32'h4241333b, 32'hc0d2e190};
test_bias[1973:1973] = '{32'hc2222ae2};
test_output[1973:1973] = '{32'hc5db41c6};
test_input[15792:15799] = '{32'h421b5958, 32'h421ff40f, 32'hc2a26e30, 32'hc0062f20, 32'h422bf8cd, 32'h4211843c, 32'hc28cea89, 32'h404afb14};
test_weights[15792:15799] = '{32'h41b2284c, 32'h42728a07, 32'h41b2daed, 32'hc0218116, 32'hc2b94348, 32'hc23fbec1, 32'h42baf8d5, 32'hbf4c84e0};
test_bias[1974:1974] = '{32'hc2a7d8ec};
test_output[1974:1974] = '{32'hc62aa221};
test_input[15800:15807] = '{32'h422200f6, 32'hc236d07e, 32'hc22ae087, 32'hc23b7e57, 32'h40e8250b, 32'h425e01ff, 32'h42077c0b, 32'hc21f1ffc};
test_weights[15800:15807] = '{32'h424d0b7a, 32'hc24561e5, 32'hbf3270d9, 32'hc2bdc0f4, 32'h41f00b19, 32'hc1c61e06, 32'hc290c29a, 32'hc259a513};
test_bias[1975:1975] = '{32'h41750825};
test_output[1975:1975] = '{32'h45e69e9c};
test_input[15808:15815] = '{32'hc2a1cb5f, 32'h429562f2, 32'hc2461a7b, 32'hc2021f7d, 32'h423ea57a, 32'hc23ae64c, 32'h41d8fcd5, 32'hc2aa0022};
test_weights[15808:15815] = '{32'h4280729f, 32'hc2b79fe0, 32'hc2515aca, 32'hc278f1b8, 32'hc2b0cf2d, 32'h4293d5de, 32'h42329c04, 32'h423c02ee};
test_bias[1976:1976] = '{32'hc21e8029};
test_output[1976:1976] = '{32'hc68c0f49};
test_input[15816:15823] = '{32'h422edd2c, 32'hc25581da, 32'h423f8851, 32'hc2b653bb, 32'h42b36517, 32'hc1f6e027, 32'hc2ade363, 32'hc29ed717};
test_weights[15816:15823] = '{32'hc095b60b, 32'hc11f4b08, 32'h3f9fc250, 32'h426c1121, 32'h41c05af6, 32'h41c2b37b, 32'h41206cba, 32'h42b4ff4e};
test_bias[1977:1977] = '{32'h3ff25690};
test_output[1977:1977] = '{32'hc635f475};
test_input[15824:15831] = '{32'h429b385e, 32'h41cfabee, 32'h427a0226, 32'hc20c9945, 32'hc1e68ec8, 32'h4223923d, 32'hc1ef2908, 32'h40668647};
test_weights[15824:15831] = '{32'h40dcbca1, 32'hc18c739e, 32'hc2a9d88d, 32'h425ed782, 32'h42b3fc2b, 32'h42b02778, 32'h4201db70, 32'hc2704a55};
test_bias[1978:1978] = '{32'hc253dd15};
test_output[1978:1978] = '{32'hc5e7d14d};
test_input[15832:15839] = '{32'h42b3734a, 32'h4263d710, 32'h42864230, 32'hc0bc526b, 32'h424e63cc, 32'h420566cf, 32'hc18c1e3c, 32'hc2c5b929};
test_weights[15832:15839] = '{32'hc2a77596, 32'h40a0de99, 32'h425b0ab3, 32'hc186850e, 32'hc05fddfb, 32'hc25307bc, 32'hc25a7cc5, 32'hc0c884c4};
test_bias[1979:1979] = '{32'hc1022f8a};
test_output[1979:1979] = '{32'hc56ef412};
test_input[15840:15847] = '{32'h427170a8, 32'h41b1958c, 32'h4048cc4d, 32'hc26b566b, 32'h426fadb3, 32'h41a19aa0, 32'hc18d3790, 32'hc26ee0d6};
test_weights[15840:15847] = '{32'hc057c2fd, 32'hc2590a07, 32'h42abe07b, 32'h3ee9fc49, 32'h425a70e3, 32'hc1383a67, 32'hc2a5e505, 32'h4287723d};
test_bias[1980:1980] = '{32'hc294c858};
test_output[1980:1980] = '{32'hc4430ab7};
test_input[15848:15855] = '{32'hc218f68f, 32'hc1286aa2, 32'h41a11988, 32'hc2ba3ae7, 32'hc2aa3393, 32'h425afb59, 32'hc26e3a7c, 32'h429e1463};
test_weights[15848:15855] = '{32'hc283d7a5, 32'h41ac3417, 32'hc19feba5, 32'hc255ed63, 32'h42a6cdbe, 32'hc2825b9c, 32'h42372a92, 32'h42740b93};
test_bias[1981:1981] = '{32'hc2c40370};
test_output[1981:1981] = '{32'hc4e09fc8};
test_input[15856:15863] = '{32'hc182d592, 32'hc12e355d, 32'h42190dd5, 32'hc03934b3, 32'h418cf3bd, 32'h41d097d0, 32'hc28032e2, 32'h41fb7152};
test_weights[15856:15863] = '{32'h41a8a75e, 32'hc2403537, 32'hc2843b8b, 32'h41a14b0c, 32'h422a4018, 32'h42a21803, 32'hc28dba5f, 32'hc164555e};
test_bias[1982:1982] = '{32'h42c6cba9};
test_output[1982:1982] = '{32'h45913487};
test_input[15864:15871] = '{32'h42502452, 32'hc258a6bb, 32'h423495b2, 32'hc12827fc, 32'hc292e18c, 32'hc009128f, 32'hc269d699, 32'hc2c66f08};
test_weights[15864:15871] = '{32'hc286035f, 32'h41a74735, 32'hc2b13913, 32'h42411f77, 32'hc27e234e, 32'hc2b17233, 32'h41d974d4, 32'h41760b3b};
test_bias[1983:1983] = '{32'hc1f6eaed};
test_output[1983:1983] = '{32'hc5e7c611};
test_input[15872:15879] = '{32'h429c6af9, 32'hc2bc7aec, 32'h425d2646, 32'hc2a48b83, 32'h3e7107ea, 32'h4227dd68, 32'h418b5ac5, 32'h42b8a852};
test_weights[15872:15879] = '{32'hc09ece22, 32'hc143e580, 32'hc2a4fad7, 32'hc28f1ed1, 32'hc282100f, 32'hc204f49e, 32'h4247ec60, 32'hc1ddc688};
test_bias[1984:1984] = '{32'hc0d37910};
test_output[1984:1984] = '{32'hc47d4f1b};
test_input[15880:15887] = '{32'hc2a923ce, 32'hc29633b2, 32'hc21481c0, 32'hc27f8cea, 32'hc23ecd29, 32'hc2986e40, 32'h415b70ca, 32'h4281f0c6};
test_weights[15880:15887] = '{32'hc2a93a62, 32'h4288da0a, 32'hc2142067, 32'h419df2e5, 32'hc2b99c68, 32'hc215cdc5, 32'hc0574fcc, 32'hc29dd4ef};
test_bias[1985:1985] = '{32'hc2bc67e9};
test_output[1985:1985] = '{32'h458180dc};
test_input[15888:15895] = '{32'hc2b969a8, 32'hc2c19b5c, 32'h41cb2ec4, 32'h4196a681, 32'hbff962a7, 32'h42701a7a, 32'h42b14ace, 32'h4287ed84};
test_weights[15888:15895] = '{32'hc22b841e, 32'h4284dbba, 32'h41dff595, 32'hc2ac959a, 32'hc219a2c3, 32'h427bf8e1, 32'hc00dadca, 32'hc1182e73};
test_bias[1986:1986] = '{32'h4235f034};
test_output[1986:1986] = '{32'hc39b446a};
test_input[15896:15903] = '{32'hc0709d66, 32'h4251270f, 32'h41f9723b, 32'hbec575f5, 32'h429222ea, 32'h4257c8e9, 32'h41930bdd, 32'hc281e828};
test_weights[15896:15903] = '{32'hc2bc9252, 32'hc2a54a65, 32'hc27d0555, 32'h4230fe7c, 32'hc20f9a96, 32'h41f5c665, 32'h42a41a5b, 32'h4289abe9};
test_bias[1987:1987] = '{32'hc1fd403c};
test_output[1987:1987] = '{32'hc61af330};
test_input[15904:15911] = '{32'hc1feef41, 32'h41f65956, 32'h42c229c5, 32'hc0acea82, 32'h40af9bc8, 32'h40378fa7, 32'h4149971a, 32'h4299f6b4};
test_weights[15904:15911] = '{32'h4232d050, 32'h42c06a9c, 32'h4242321b, 32'h429392cd, 32'hc2851768, 32'hc2c1ce4a, 32'hc286c09c, 32'hc20b4128};
test_bias[1988:1988] = '{32'hc1f25373};
test_output[1988:1988] = '{32'h44ce46ae};
test_input[15912:15919] = '{32'h41f82e7a, 32'h42107876, 32'h4294d7ce, 32'hc2a8dd27, 32'h423dd391, 32'hc21b585d, 32'hc2528e65, 32'h421824ee};
test_weights[15912:15919] = '{32'hc2be24f8, 32'h41cc8e21, 32'hc270182e, 32'h42c0c0da, 32'hc187651b, 32'h42a2fa6b, 32'hc247786e, 32'h42ae26e9};
test_bias[1989:1989] = '{32'h42c1a161};
test_output[1989:1989] = '{32'hc6445124};
test_input[15920:15927] = '{32'hc1d50b2b, 32'h421af7ee, 32'h425ddb46, 32'hc2af085c, 32'hc22b9c41, 32'h406e042a, 32'h4298f4df, 32'hc295eb6c};
test_weights[15920:15927] = '{32'h42877115, 32'hc1861b74, 32'hc29ff210, 32'h4209b316, 32'hc1a62f78, 32'hc283346a, 32'h41107e5c, 32'hc2444daf};
test_bias[1990:1990] = '{32'h42c0e960};
test_output[1990:1990] = '{32'hc595a14f};
test_input[15928:15935] = '{32'hc26fa2b7, 32'hc2265ff3, 32'hc242d0d5, 32'hc1dd723e, 32'hc2a91e82, 32'hc2c50eb5, 32'h4290eba9, 32'h42b7312c};
test_weights[15928:15935] = '{32'hc185fee2, 32'h42426d0f, 32'h3de317eb, 32'hc28d6ade, 32'hc23a5211, 32'h42a35372, 32'h42c64cbf, 32'hc2174b0c};
test_bias[1991:1991] = '{32'hc287144c};
test_output[1991:1991] = '{32'h43ef54f2};
test_input[15936:15943] = '{32'h412946a8, 32'h42a3025b, 32'h42adbdbd, 32'hc24f8749, 32'hc2b05cd8, 32'hc143aae5, 32'hc221b856, 32'h41c33f4b};
test_weights[15936:15943] = '{32'h425212bd, 32'h428c1950, 32'hc14dd445, 32'hc190cf86, 32'h424f4413, 32'hc2bf5be7, 32'h4206c0c3, 32'hc21c71f1};
test_bias[1992:1992] = '{32'hc2a0d778};
test_output[1992:1992] = '{32'h439138a5};
test_input[15944:15951] = '{32'hc12496cf, 32'h4295a90f, 32'hbf5e9bb6, 32'h4107817a, 32'hc2969485, 32'h41180652, 32'hc25495d2, 32'hc2839340};
test_weights[15944:15951] = '{32'h4241a7a0, 32'hc1a2bca6, 32'hc289da2e, 32'h42973468, 32'hc2675e55, 32'h41027de6, 32'hc26d2ef2, 32'h419be9bc};
test_bias[1993:1993] = '{32'h428aa69d};
test_output[1993:1993] = '{32'h459dd7b0};
test_input[15952:15959] = '{32'h42128222, 32'h425f1d72, 32'h42a56a4e, 32'h41a979b0, 32'h4141b1bd, 32'hc1c752b7, 32'h42c5ff99, 32'hc17d7be2};
test_weights[15952:15959] = '{32'hbdb0e0fb, 32'hc23cd22f, 32'h41f2d983, 32'h41b884f9, 32'hc2b21c73, 32'h42096b59, 32'hc10299a1, 32'hc1b4c843};
test_bias[1994:1994] = '{32'h42bca23c};
test_output[1994:1994] = '{32'hc4f0d71a};
test_input[15960:15967] = '{32'h41c92734, 32'h419eea8d, 32'hc29b3e06, 32'h428d961c, 32'hc264aa7a, 32'h42bb4d4b, 32'hc2033d31, 32'hc2a1be6d};
test_weights[15960:15967] = '{32'h4298d4cb, 32'hc2bd691f, 32'h41163d9f, 32'h4163999a, 32'hc266e574, 32'hc2bbc7d9, 32'h427366d2, 32'hc2010204};
test_bias[1995:1995] = '{32'hc257d442};
test_output[1995:1995] = '{32'hc5904741};
test_input[15968:15975] = '{32'hc1a4f278, 32'hc0103d0a, 32'h42baada4, 32'hc0b00376, 32'h42216b4c, 32'h41861216, 32'h42beda4d, 32'hc2824afc};
test_weights[15968:15975] = '{32'hc2beea65, 32'hc18b2f97, 32'h42776ba3, 32'hc20d1655, 32'h41b11ea5, 32'hbfa9aa34, 32'hc215d36f, 32'h42c5b5f8};
test_bias[1996:1996] = '{32'hc27825df};
test_output[1996:1996] = '{32'hc499c9a9};
test_input[15976:15983] = '{32'h423ec55e, 32'hbdce4374, 32'hc2a9e8e2, 32'hc225ec60, 32'h422e375b, 32'h42389fce, 32'h4295ffe3, 32'h42c52de5};
test_weights[15976:15983] = '{32'h423b19d2, 32'hc1c6a5fb, 32'h42167376, 32'h41c1593a, 32'h41ffe2f2, 32'h42370a14, 32'hc2b55850, 32'hc0ea2a36};
test_bias[1997:1997] = '{32'hc270d1d6};
test_output[1997:1997] = '{32'hc5bccb83};
test_input[15984:15991] = '{32'hc28055b5, 32'h42af6274, 32'hc2c4704e, 32'hc2af0cdc, 32'hc236b089, 32'hc18585a9, 32'hc062b220, 32'hc1d3b103};
test_weights[15984:15991] = '{32'h41acf679, 32'hc1bd401d, 32'hc220155f, 32'hc25b563d, 32'hc26f696d, 32'hc158a6e8, 32'hc2a9317d, 32'h4219bb23};
test_bias[1998:1998] = '{32'h42b35ed4};
test_output[1998:1998] = '{32'h45ed8301};
test_input[15992:15999] = '{32'h4156e211, 32'h42bcde3b, 32'h412b5dc9, 32'hbeed4fed, 32'hc2b10ae8, 32'hc2a13ef5, 32'hc22c0fbb, 32'h420a7238};
test_weights[15992:15999] = '{32'hc27f71e8, 32'h4111a37a, 32'hc2a705b2, 32'hc1b6eddd, 32'h428929bb, 32'hc1b44e7b, 32'h42bb0c1a, 32'hc200d4b8};
test_bias[1999:1999] = '{32'hc28d7e81};
test_output[1999:1999] = '{32'hc621a0d4};
test_input[16000:16007] = '{32'h42906024, 32'hc2148979, 32'h400d8e0d, 32'hc262cee3, 32'hc29e7fa8, 32'hc2b9e588, 32'hc262a739, 32'hc280af0b};
test_weights[16000:16007] = '{32'h422831a9, 32'h40ce0f24, 32'hc2722378, 32'h42a498c6, 32'hbf406efe, 32'h4289e55e, 32'hc1876efa, 32'h4287d7e0};
test_bias[2000:2000] = '{32'hc092107c};
test_output[2000:2000] = '{32'hc637e292};
test_input[16008:16015] = '{32'h41868c58, 32'h426b4561, 32'hc2bd8503, 32'hc28095ae, 32'hc211ceee, 32'h403475ef, 32'h425142a1, 32'h3f4a9e70};
test_weights[16008:16015] = '{32'hc1475fa9, 32'h42afb9d1, 32'hc202d42a, 32'h4038a2f6, 32'hc23dabcd, 32'h41083921, 32'hc2b131f8, 32'h42c7c9f9};
test_bias[2001:2001] = '{32'hc2a70b40};
test_output[2001:2001] = '{32'h459bc9ae};
test_input[16016:16023] = '{32'hbfcf386a, 32'h40a10275, 32'hc29793d0, 32'hc03b01be, 32'hc29de271, 32'hc21d5713, 32'hc20117d0, 32'h425fb6a7};
test_weights[16016:16023] = '{32'hc287978f, 32'hc2091750, 32'hc2b77b26, 32'hc259d7e9, 32'h424f0627, 32'h422e6c28, 32'hc26f02c0, 32'h41ac75dd};
test_bias[2002:2002] = '{32'hc2756dc6};
test_output[2002:2002] = '{32'h458708df};
test_input[16024:16031] = '{32'hc2912705, 32'h42725eb9, 32'h41e83c30, 32'h4288e8f9, 32'hc2a4913e, 32'h40777a50, 32'hc24274de, 32'h42869bdf};
test_weights[16024:16031] = '{32'h428270d1, 32'h4181c522, 32'hc28426cb, 32'hc2aab056, 32'h41fe550f, 32'h4278ebd1, 32'hc2a86e60, 32'h42b2bb9a};
test_bias[2003:2003] = '{32'h4228d806};
test_output[2003:2003] = '{32'hc5697353};
test_input[16032:16039] = '{32'h42b05a19, 32'h41bc1e48, 32'hc20ec21f, 32'hc2c0c81c, 32'h428f758e, 32'hc11ed514, 32'hc05bade1, 32'hc2b03fde};
test_weights[16032:16039] = '{32'h42b0cdc3, 32'h4128cae6, 32'hc2222cf1, 32'h42bdd067, 32'hc1c27331, 32'hc2a466cf, 32'h42703fa8, 32'h425e462d};
test_bias[2004:2004] = '{32'h41dd8e74};
test_output[2004:2004] = '{32'hc5b0e8a7};
test_input[16040:16047] = '{32'hc175880a, 32'hc2c195c2, 32'h41c008ed, 32'h42808f30, 32'hc23c5798, 32'h41efbab8, 32'hc078547d, 32'hc29c01cc};
test_weights[16040:16047] = '{32'hc25323f2, 32'h42a43a5e, 32'h42620e33, 32'h41c3aec7, 32'hc1ce3009, 32'hc218580f, 32'h429004c9, 32'hc1e8c0e4};
test_bias[2005:2005] = '{32'hc242fb60};
test_output[2005:2005] = '{32'hc50938d1};
test_input[16048:16055] = '{32'hc280f143, 32'h42a2c11e, 32'hc23d8b7a, 32'hc22cdd2d, 32'hc16e15af, 32'h42496142, 32'h41e9beac, 32'h428aa107};
test_weights[16048:16055] = '{32'h42880889, 32'hc1d1ac40, 32'h42743de1, 32'hc22793e2, 32'h42224ca3, 32'hc19b0805, 32'h41d7e730, 32'hc13419c5};
test_bias[2006:2006] = '{32'hc1e13011};
test_output[2006:2006] = '{32'hc60fc05a};
test_input[16056:16063] = '{32'hc29afb73, 32'h42928d37, 32'h3f947efb, 32'hc25dc5fc, 32'hc2719311, 32'hc28d912a, 32'h4181c223, 32'hc1f06cef};
test_weights[16056:16063] = '{32'hc0b428bb, 32'hc0df74ef, 32'h429148af, 32'h42b57872, 32'hc17e20d8, 32'hc260a508, 32'hc2823afe, 32'h42a8c47e};
test_bias[2007:2007] = '{32'hc2166ae8};
test_output[2007:2007] = '{32'hc56850c8};
test_input[16064:16071] = '{32'hc2992bca, 32'h42b899fa, 32'hc2c09da7, 32'h40a9e663, 32'hc17690c9, 32'h3fae0a28, 32'hc238c6bb, 32'hc2048e4c};
test_weights[16064:16071] = '{32'h4207a6d7, 32'hc105b249, 32'h42817033, 32'h4293348a, 32'h42a7f9f3, 32'hc0f22c70, 32'h41923ba0, 32'h42a68080};
test_bias[2008:2008] = '{32'h404e5c98};
test_output[2008:2008] = '{32'hc65c8d1d};
test_input[16072:16079] = '{32'hc269274f, 32'h414430d9, 32'h42a3019c, 32'hc2b88c21, 32'hc263e7e7, 32'hc067a75a, 32'h4297ee80, 32'h412495bf};
test_weights[16072:16079] = '{32'hc21e0dc6, 32'hc2aa68b9, 32'h4212851c, 32'h428827b0, 32'h41c7a272, 32'h42c473e9, 32'hc1c5f7bb, 32'h4272aa7f};
test_bias[2009:2009] = '{32'h412b2d4c};
test_output[2009:2009] = '{32'hc59e22c9};
test_input[16080:16087] = '{32'h427dcb53, 32'hc2632c5b, 32'hc25a8d57, 32'hc263329d, 32'h42bb1672, 32'hc1bf20df, 32'h427aed11, 32'h42c7465f};
test_weights[16080:16087] = '{32'hc2924d18, 32'h420511ab, 32'h41a2c9e7, 32'hc2b9e8d1, 32'hc133c4a7, 32'hc1dd7640, 32'hc2a6740e, 32'h41edc503};
test_bias[2010:2010] = '{32'hc21714db};
test_output[2010:2010] = '{32'hc59dcd89};
test_input[16088:16095] = '{32'h42be2ba3, 32'h42a87975, 32'hc2bf84e8, 32'hc2900cc5, 32'h42913def, 32'h42b1011e, 32'hc2821518, 32'hc2099b73};
test_weights[16088:16095] = '{32'hc26cd51c, 32'h419f9ce3, 32'h42b7ce5e, 32'hc2be36b3, 32'h425d3474, 32'hc2212320, 32'h42a61777, 32'hc294e4bc};
test_bias[2011:2011] = '{32'hc2beb8f3};
test_output[2011:2011] = '{32'hc6030241};
test_input[16096:16103] = '{32'h4281586b, 32'h40f58207, 32'h41472ced, 32'h4286e9e0, 32'hc2812b9f, 32'hc21c65f7, 32'h42466850, 32'hc136cc94};
test_weights[16096:16103] = '{32'h42717ed0, 32'h411a62e2, 32'h4226d0a1, 32'hc258b851, 32'h4213fec9, 32'h42a8f609, 32'h428d78e6, 32'h420128e5};
test_bias[2012:2012] = '{32'hc2a26f7c};
test_output[2012:2012] = '{32'hc4dfe9d0};
test_input[16104:16111] = '{32'hc25a1e3a, 32'h42a431fc, 32'hc2702204, 32'hc1e93c9c, 32'hc2246443, 32'hc0d46557, 32'hc2c2d202, 32'h41c0ffc5};
test_weights[16104:16111] = '{32'hc194c45a, 32'h41aaa8aa, 32'hc2ba7f1e, 32'hc29d3be6, 32'h41236d45, 32'h4112ab30, 32'h4028120a, 32'h42a3ac1e};
test_bias[2013:2013] = '{32'hc1991d4a};
test_output[2013:2013] = '{32'h46398876};
test_input[16112:16119] = '{32'h4281932b, 32'hc2c78236, 32'h4278c538, 32'h41fbda8c, 32'hc179f904, 32'hc1ea19d2, 32'h428f5359, 32'h428751f3};
test_weights[16112:16119] = '{32'h42648c5d, 32'hc26449dd, 32'h4241633b, 32'h42851717, 32'hc2c751e6, 32'h4067aa5a, 32'h40b9463c, 32'hc08f02d6};
test_bias[2014:2014] = '{32'hc1672aa7};
test_output[2014:2014] = '{32'h467ab7a4};
test_input[16120:16127] = '{32'h41c29eeb, 32'h42b6af4c, 32'hc16533b6, 32'hc1b86730, 32'hc24d17dd, 32'hc286e972, 32'h42929fb4, 32'h42a72d7c};
test_weights[16120:16127] = '{32'hc2b7b8ef, 32'h41cb2ef9, 32'h425ee9d1, 32'h416a9209, 32'hc2500e59, 32'h429ca3ea, 32'hc1d5edb0, 32'h3fa667e3};
test_bias[2015:2015] = '{32'hbf6fe9fc};
test_output[2015:2015] = '{32'hc5ac8050};
test_input[16128:16135] = '{32'h422a0132, 32'h42c76f53, 32'h418bd2f3, 32'h41ab9a09, 32'hc278009f, 32'h40ea356e, 32'hbfee5720, 32'h429c7c85};
test_weights[16128:16135] = '{32'h41a5ca0e, 32'h42339ec6, 32'h4289c418, 32'h42abed28, 32'h423a3fc1, 32'hc1b53888, 32'h420f53e6, 32'hc20cd361};
test_bias[2016:2016] = '{32'h4247ab7c};
test_output[2016:2016] = '{32'h452164ff};
test_input[16136:16143] = '{32'hc207593b, 32'h41e3ea76, 32'hc24b28f8, 32'hc2773618, 32'h42c3be38, 32'hc2095154, 32'h42896cd4, 32'h42014e9d};
test_weights[16136:16143] = '{32'h42851cdc, 32'h4291bc30, 32'hc22192b4, 32'hc14818e9, 32'hc106fae4, 32'h4214b808, 32'h413c7b26, 32'hc209ea49};
test_bias[2017:2017] = '{32'h4188db15};
test_output[2017:2017] = '{32'h4381261b};
test_input[16144:16151] = '{32'h42036229, 32'h40a10fd0, 32'h41acfa69, 32'hc288457c, 32'hc28e9d10, 32'hc2b35acc, 32'hc2030da9, 32'h410a9228};
test_weights[16144:16151] = '{32'hc2763c0b, 32'hc225c47a, 32'h42250b33, 32'h42bd69ef, 32'h418a95d3, 32'h42a55946, 32'hc1b605bf, 32'hc2a19e4f};
test_bias[2018:2018] = '{32'h3fbac3be};
test_output[2018:2018] = '{32'hc6801309};
test_input[16152:16159] = '{32'h42b108be, 32'hc003b70f, 32'hc2767b45, 32'hc013dcae, 32'h41b03130, 32'hc2456693, 32'h42aaee9f, 32'hc2a4f2c9};
test_weights[16152:16159] = '{32'hc0930857, 32'hc27cc3bc, 32'hc29c9e9d, 32'h418563b5, 32'hc27388b4, 32'h42824097, 32'h42c44d7a, 32'h41fa3177};
test_bias[2019:2019] = '{32'h42223dcb};
test_output[2019:2019] = '{32'h45b56a1a};
test_input[16160:16167] = '{32'hc1dad1d1, 32'h414753c6, 32'hc15fcad9, 32'hc2bfe63c, 32'hc091db56, 32'hc2c654d9, 32'h41f315bb, 32'h42947ef3};
test_weights[16160:16167] = '{32'h42a33585, 32'hc2ad15dd, 32'h4253327a, 32'h42b3d29d, 32'h42b64276, 32'h416273b9, 32'h424315dd, 32'hc276bfdd};
test_bias[2020:2020] = '{32'h42349138};
test_output[2020:2020] = '{32'hc6891752};
test_input[16168:16175] = '{32'hc290ab3a, 32'hc23e3a72, 32'hc1bbde25, 32'h4257b2b0, 32'h42b63182, 32'hc28f08ad, 32'h422bca93, 32'hc260a24b};
test_weights[16168:16175] = '{32'hc1b11586, 32'h42573e9a, 32'h4282b8f5, 32'h42b53b59, 32'h42b04c5c, 32'h40ea9d77, 32'h4289294d, 32'hc134ed96};
test_bias[2021:2021] = '{32'h42c03274};
test_output[2021:2021] = '{32'h46541f67};
test_input[16176:16183] = '{32'h419cde88, 32'hc18ebd81, 32'hc158ced6, 32'hc2a9eb00, 32'hbf0cce42, 32'h4185f866, 32'hc193d49f, 32'hc131c72c};
test_weights[16176:16183] = '{32'hc152c782, 32'h426a1859, 32'hc20b90c2, 32'h427e7080, 32'hc1d9c8f5, 32'hc0af43cd, 32'h41d5d2d5, 32'hc2a6312d};
test_bias[2022:2022] = '{32'h413d7712};
test_output[2022:2022] = '{32'hc5b76bd8};
test_input[16184:16191] = '{32'hc0cc60a0, 32'h419e93c8, 32'hc0bf1e1f, 32'h40cee76f, 32'h421b3e26, 32'hc2aaa226, 32'hc1b63c2b, 32'hc1d02dbb};
test_weights[16184:16191] = '{32'h42654d50, 32'h426b91bf, 32'hc1917e6e, 32'hc1a85b14, 32'hc2af6c33, 32'hc1f4973a, 32'hc2c7bb0d, 32'h4188da5e};
test_bias[2023:2023] = '{32'hc1422159};
test_output[2023:2023] = '{32'h44e0767b};
test_input[16192:16199] = '{32'hc2a8c44b, 32'hc2371f6b, 32'h42c53c35, 32'h41ef027a, 32'hc26310e0, 32'h41f5504e, 32'hc29595a7, 32'h421c1af0};
test_weights[16192:16199] = '{32'h41b571ae, 32'hc215f430, 32'hc2b96948, 32'hc1c6f3d1, 32'hc1818508, 32'h42a7517b, 32'h42c629da, 32'h42ade900};
test_bias[2024:2024] = '{32'hc21ec935};
test_output[2024:2024] = '{32'hc6267d54};
test_input[16200:16207] = '{32'hc29a26e3, 32'h4116585d, 32'hc28bcddc, 32'h428d94b3, 32'h423aac58, 32'hc2817b2c, 32'hc1b2533b, 32'h42a12247};
test_weights[16200:16207] = '{32'h3f044a0f, 32'h42865e50, 32'h41a60c14, 32'hc1ec6d6d, 32'h41c5da74, 32'hc2a0097f, 32'h42965fcd, 32'hc29b0f86};
test_bias[2025:2025] = '{32'hc27ecbbc};
test_output[2025:2025] = '{32'hc58fd768};
test_input[16208:16215] = '{32'hc2a8296e, 32'h40b4e7ad, 32'h427a3d85, 32'h423e8521, 32'hc0ea7596, 32'h425cb5b2, 32'h42a284f7, 32'hc2072aba};
test_weights[16208:16215] = '{32'hc1c3e8c1, 32'h42b0c7cb, 32'h4287f173, 32'hc29c41aa, 32'h42b1c775, 32'hc1a74ba6, 32'hc2adc993, 32'h41a20b1b};
test_bias[2026:2026] = '{32'h41f8e2de};
test_output[2026:2026] = '{32'hc5c8ed6c};
test_input[16216:16223] = '{32'h41f60cb4, 32'h424fc8c6, 32'h42940293, 32'hc22d99eb, 32'h41efd645, 32'hc2668d65, 32'h42130757, 32'hc2c66a73};
test_weights[16216:16223] = '{32'hc2c3a67b, 32'hc0dbb012, 32'hc1da4628, 32'hc1d48990, 32'h42b83728, 32'h422d0bc1, 32'hc225ee24, 32'hc2ac4e2e};
test_bias[2027:2027] = '{32'h42bd426f};
test_output[2027:2027] = '{32'h4545138c};
test_input[16224:16231] = '{32'hc2afcf12, 32'hc2b55e24, 32'h421a2aca, 32'hc2bf4a41, 32'hc2c1d04d, 32'hc2952d3d, 32'h41f16698, 32'hc21c30ac};
test_weights[16224:16231] = '{32'h420e77f3, 32'h4082e145, 32'hc219755c, 32'h42512f02, 32'hc23098e8, 32'h4280af6a, 32'h42a8490b, 32'hc29397fc};
test_bias[2028:2028] = '{32'h41a54879};
test_output[2028:2028] = '{32'hc59e2eec};
test_input[16232:16239] = '{32'h42181d57, 32'h429284dc, 32'h408c3bf1, 32'h42475a05, 32'hc230b5ba, 32'h420901de, 32'hc206523b, 32'hc2695cfd};
test_weights[16232:16239] = '{32'h417a3939, 32'hc283adef, 32'h426aa94e, 32'h42737cdc, 32'hc24d8a86, 32'hc2603274, 32'hc2a81015, 32'hc2c25555};
test_bias[2029:2029] = '{32'h4051a385};
test_output[2029:2029] = '{32'h45f71270};
test_input[16240:16247] = '{32'h42c01f24, 32'hc21bc48a, 32'hc2826c6b, 32'h42607359, 32'hc1099dfe, 32'h4275f2f6, 32'hc0a6b483, 32'h42009ced};
test_weights[16240:16247] = '{32'hc2b1b917, 32'hc2a36dfb, 32'h429ae062, 32'h4251582f, 32'hc1920efe, 32'hc28a6fcc, 32'hc277d0d3, 32'h429e4dde};
test_bias[2030:2030] = '{32'hc2c66a20};
test_output[2030:2030] = '{32'hc6097678};
test_input[16248:16255] = '{32'h3fb733b1, 32'hc1bbead6, 32'hc183a67b, 32'hc2096aa8, 32'h418fe2f6, 32'hc1d978f8, 32'h4206d4ee, 32'h41cd07f3};
test_weights[16248:16255] = '{32'h421fca17, 32'hc1c0a391, 32'hc2bc0385, 32'h42302faa, 32'h42a2f89c, 32'h42c08fec, 32'h40ee07b3, 32'h427b10f4};
test_bias[2031:2031] = '{32'h425bf70b};
test_output[2031:2031] = '{32'h44b1685a};
test_input[16256:16263] = '{32'hc24f91fc, 32'hc1ef4eb3, 32'h41d80a49, 32'h418a6b1f, 32'h41f8cd4b, 32'h42c012e1, 32'h41ef897a, 32'hc1d3cbc1};
test_weights[16256:16263] = '{32'h42174067, 32'h42c1a443, 32'h428465c2, 32'hc1fb2ffb, 32'hc1da3d13, 32'h41808882, 32'hbfb98a99, 32'hc26f32f8};
test_bias[2032:2032] = '{32'hc1b01104};
test_output[2032:2032] = '{32'hc4af35ae};
test_input[16264:16271] = '{32'h428fe3c6, 32'h41a6fbe5, 32'hc17961d4, 32'hc1eb7ae1, 32'hc2c1c387, 32'hc275fbe9, 32'h409624fb, 32'hc2a80f1f};
test_weights[16264:16271] = '{32'h41316bdc, 32'hc2b6bb7f, 32'hc2402120, 32'hc1e1062a, 32'hc2c00884, 32'h4143ec0a, 32'h4252af7d, 32'h42a9488f};
test_bias[2033:2033] = '{32'h41838d13};
test_output[2033:2033] = '{32'h45077b7d};
test_input[16272:16279] = '{32'hc19931a0, 32'hc29e54d1, 32'h41d31806, 32'h42aa9c89, 32'hc247ae58, 32'hc27553b6, 32'h42002fe8, 32'hc1c37841};
test_weights[16272:16279] = '{32'hc25f5e59, 32'hc24edc27, 32'hc244b931, 32'h425fdcb9, 32'h41c0d0ab, 32'h42a091a0, 32'hc0a298a4, 32'hc28951a1};
test_bias[2034:2034] = '{32'h4104eb3f};
test_output[2034:2034] = '{32'h457c3c48};
test_input[16280:16287] = '{32'h429ea8fd, 32'hc247af5e, 32'hc291283a, 32'hc20ec0eb, 32'hc2bfbe59, 32'hc234cdd2, 32'hc26d2963, 32'h42aaad10};
test_weights[16280:16287] = '{32'hc2bb6ba0, 32'h423ad94a, 32'hbf00775e, 32'hc290d842, 32'h41439c9a, 32'hc21884a3, 32'hc2a2d471, 32'h4265766e};
test_bias[2035:2035] = '{32'h40fb29d1};
test_output[2035:2035] = '{32'h45440ed4};
test_input[16288:16295] = '{32'h42702171, 32'hc2569505, 32'h41dd9729, 32'h42047181, 32'h416425a3, 32'h406f9656, 32'hc1132143, 32'h427efeb1};
test_weights[16288:16295] = '{32'h414cae8f, 32'h42c7d4f6, 32'hc2bc160e, 32'hc22dd8ef, 32'h42335548, 32'hc26d530b, 32'hc1c82955, 32'h42c717d6};
test_bias[2036:2036] = '{32'hc2b060e6};
test_output[2036:2036] = '{32'hc4d85f52};
test_input[16296:16303] = '{32'hc2b2ed55, 32'h42c4933f, 32'h4020e06c, 32'hc22f4738, 32'h42381743, 32'hc293a4c1, 32'h42b541b2, 32'h42b7cce6};
test_weights[16296:16303] = '{32'h41d35b89, 32'h42bd57d3, 32'hc26fcdd0, 32'h423d5fce, 32'hc28ccb40, 32'hc288e8bc, 32'h41d944ea, 32'hc137c88d};
test_bias[2037:2037] = '{32'h42622a4a};
test_output[2037:2037] = '{32'h45f9c025};
test_input[16304:16311] = '{32'hc27da964, 32'hc2795fd2, 32'hc051a43e, 32'hc1b59f37, 32'hc28629ba, 32'hc24598f5, 32'h4090c485, 32'hc2ab8231};
test_weights[16304:16311] = '{32'hc24ae0d1, 32'hc1b70c19, 32'hc189c47f, 32'h4216cb74, 32'hc225fd1b, 32'hc1f8a3cf, 32'hc0cb6fc7, 32'hc22012de};
test_bias[2038:2038] = '{32'h41bb69ff};
test_output[2038:2038] = '{32'h46351377};
test_input[16312:16319] = '{32'hc1e9468a, 32'hc21fb359, 32'h40516578, 32'hc210352a, 32'h41136f1a, 32'hc20de3d4, 32'h42412c3e, 32'hc27df645};
test_weights[16312:16319] = '{32'hc21b9e2c, 32'h4112cdce, 32'hc25e4f2d, 32'hc23abcff, 32'hc24a31e5, 32'hc27bb27b, 32'hbff256e2, 32'h420c3a27};
test_bias[2039:2039] = '{32'h41f71979};
test_output[2039:2039] = '{32'h44daaa14};
test_input[16320:16327] = '{32'h429f9e36, 32'hc2292cf8, 32'hc2302e13, 32'h42c17583, 32'hc1e79974, 32'h418a392a, 32'hc2a77cec, 32'h42c77b3a};
test_weights[16320:16327] = '{32'hc216ddc1, 32'h4230b8f0, 32'h4258fb1f, 32'hc2a3d225, 32'hc1d84fc6, 32'h42b6d81b, 32'hc010dc01, 32'h41a120a7};
test_bias[2040:2040] = '{32'hc27838d4};
test_output[2040:2040] = '{32'hc627116e};
test_input[16328:16335] = '{32'hc28c196c, 32'h41a96326, 32'hc2621d7f, 32'h4265667d, 32'hc295da02, 32'h4290548e, 32'h42abea9a, 32'hc1ed2573};
test_weights[16328:16335] = '{32'hc2981a06, 32'hc2403106, 32'hc2385dc6, 32'hc2861812, 32'hc29b322b, 32'h42858cf0, 32'hc22952f0, 32'hc29a3978};
test_bias[2041:2041] = '{32'h428a0934};
test_output[2041:2041] = '{32'h46420ddd};
test_input[16336:16343] = '{32'hc286fd48, 32'hc2aee441, 32'hc0f64b03, 32'h40b3b795, 32'hc26c448e, 32'h421d1082, 32'h4229ae5d, 32'hc2121f39};
test_weights[16336:16343] = '{32'h41aab0aa, 32'hc2848bf4, 32'h4296c03c, 32'h4127f7ce, 32'h4201e1fb, 32'h42788e91, 32'hc29cd975, 32'h4261f662};
test_bias[2042:2042] = '{32'hc24cd564};
test_output[2042:2042] = '{32'hc487b1ae};
test_input[16344:16351] = '{32'hc29e47b4, 32'h427cd60f, 32'hc1f04f61, 32'hc21fbde3, 32'h42613524, 32'hc148f0b6, 32'hc2b95825, 32'hc2aeba9a};
test_weights[16344:16351] = '{32'h3fb44a38, 32'hc29d0999, 32'h424cee67, 32'hc1097e22, 32'h4099f4dd, 32'hc2c1f574, 32'hc2b00bf2, 32'h40ba74b5};
test_bias[2043:2043] = '{32'hc266db7e};
test_output[2043:2043] = '{32'h452f901e};
test_input[16352:16359] = '{32'hc12c6e2c, 32'h42b29e93, 32'hc28a4e35, 32'h4214095e, 32'h42bb6f63, 32'h42b4a79a, 32'h429501f7, 32'h42abc01b};
test_weights[16352:16359] = '{32'h429b54bb, 32'hc26ac80d, 32'h42a33583, 32'hc2070ad5, 32'hc2c3cfad, 32'h418dac31, 32'h427d2d58, 32'h41da90f5};
test_bias[2044:2044] = '{32'h40d3373e};
test_output[2044:2044] = '{32'hc6529c68};
test_input[16360:16367] = '{32'hc23371ef, 32'h41c7826e, 32'h4220cf55, 32'hc1a92941, 32'hc23a63d2, 32'hc23252e1, 32'h42abeb45, 32'h4201732f};
test_weights[16360:16367] = '{32'hc228ff25, 32'h429bcd05, 32'h4023a319, 32'hc20bad3d, 32'hc281a390, 32'h413a57fd, 32'h424f27c6, 32'hc287fb73};
test_bias[2045:2045] = '{32'hc285caa4};
test_output[2045:2045] = '{32'h461253c9};
test_input[16368:16375] = '{32'hc249d6c4, 32'h414ba28c, 32'hc2a6cc35, 32'hc23eb286, 32'h42811e06, 32'hc2c7a0e1, 32'hc1cf4444, 32'hc2bae83c};
test_weights[16368:16375] = '{32'hc1cc2386, 32'h424824b9, 32'hc190fb1b, 32'hc1eaa30d, 32'hc1ce3a45, 32'h426bd054, 32'h42743a9a, 32'h3eda4e9e};
test_bias[2046:2046] = '{32'hc1bb0ef7};
test_output[2046:2046] = '{32'hc5883d2a};
test_input[16376:16383] = '{32'h41c79dfc, 32'hc29ece25, 32'h40f578d1, 32'h428b22c5, 32'h4231f379, 32'h4223c0f4, 32'h41b5a496, 32'h42922c8a};
test_weights[16376:16383] = '{32'hc26ddf16, 32'hc27b8fd9, 32'hc23fdec4, 32'h42948f65, 32'h42020108, 32'h42c100cd, 32'h42692d67, 32'h41ab5cb9};
test_bias[2047:2047] = '{32'hc2c44d8b};
test_output[2047:2047] = '{32'h4680e1c0};
test_input[16384:16391] = '{32'hc1cdef57, 32'hc288be26, 32'hc1f6b83f, 32'h40c5ffb6, 32'h42316769, 32'hc1639344, 32'h403bfd87, 32'hc2330798};
test_weights[16384:16391] = '{32'h42026232, 32'hc2785281, 32'h41f6e3a3, 32'hc18bdb37, 32'h42010cc2, 32'hc29f3d01, 32'h42a2c45a, 32'h41234b8f};
test_bias[2048:2048] = '{32'hc27bba6a};
test_output[2048:2048] = '{32'h4590a182};
test_input[16392:16399] = '{32'hc2761d75, 32'hc2357fdc, 32'hc280ee55, 32'hc2aa6fef, 32'h42b28685, 32'h428b3e6e, 32'h4102204f, 32'hc2b0b5dd};
test_weights[16392:16399] = '{32'hc299d141, 32'h41c2f6b2, 32'hc1e206cf, 32'h42304471, 32'h429a50be, 32'h402a0b4f, 32'h4254d911, 32'hc1f16432};
test_bias[2049:2049] = '{32'h42963930};
test_output[2049:2049] = '{32'h463a8a20};
test_input[16400:16407] = '{32'h42b29062, 32'hbfc33132, 32'h4214f622, 32'hc1ecea3c, 32'h41491ee2, 32'hc27b4fdb, 32'hc2c2d383, 32'h42865bc6};
test_weights[16400:16407] = '{32'hc1a8535d, 32'hc2b3de27, 32'hc28b96c3, 32'hc21516be, 32'h422d24b2, 32'h41ac796a, 32'hc25119cc, 32'hc16da6ef};
test_bias[2050:2050] = '{32'hc28004e4};
test_output[2050:2050] = '{32'hc1861a91};
test_input[16408:16415] = '{32'hc29c0eed, 32'h42c2b443, 32'hc2c58b8c, 32'h422400ce, 32'hc229c4e7, 32'hc25d91d1, 32'hc285a2d1, 32'hc19b7a7f};
test_weights[16408:16415] = '{32'hc21c9788, 32'hc1ef2ca9, 32'hc2af3823, 32'hc25f17ca, 32'hc21038ea, 32'h42a9d445, 32'h42220ce1, 32'h4201e743};
test_bias[2051:2051] = '{32'hc2c5ec53};
test_output[2051:2051] = '{32'hc2c72b8b};
test_input[16416:16423] = '{32'h42595cfb, 32'hc2c07e23, 32'hc2a81e3b, 32'hc298f3d4, 32'hc272b89d, 32'hc2c1127a, 32'hc0cd3739, 32'h41367fc1};
test_weights[16416:16423] = '{32'hc2a73970, 32'h426428b4, 32'hc28258e6, 32'hbf01eb42, 32'h420814af, 32'h42ab3c7d, 32'h41adde12, 32'hc1d6c3ac};
test_bias[2052:2052] = '{32'hc2b137b0};
test_output[2052:2052] = '{32'hc6704fda};
test_input[16424:16431] = '{32'hc0a29061, 32'hc2c117eb, 32'hc2ab673f, 32'hc20fc076, 32'h42b7affc, 32'h42606a81, 32'h4243bbb0, 32'hc1eba209};
test_weights[16424:16431] = '{32'h42bd3a6e, 32'hc1de4068, 32'h41e40e25, 32'hc2ad7ae3, 32'h421fbe36, 32'h42a02882, 32'h41824d68, 32'hc278cf4b};
test_bias[2053:2053] = '{32'hc24add41};
test_output[2053:2053] = '{32'h4654bb00};
test_input[16432:16439] = '{32'h41af6acc, 32'h42b00527, 32'h4265259e, 32'hc2a260b4, 32'hc22b13ee, 32'h4225a9b1, 32'hc2bef7ca, 32'hc2b9a789};
test_weights[16432:16439] = '{32'h42b3ea5d, 32'h42061692, 32'hc203b21f, 32'h42bbc1de, 32'hc2931b05, 32'h426a70a7, 32'hc288f5d2, 32'hc1e2e968};
test_bias[2054:2054] = '{32'h42bc9398};
test_output[2054:2054] = '{32'h462037dc};
test_input[16440:16447] = '{32'h409ac1e1, 32'hc1feea9e, 32'h427f8358, 32'h426a3516, 32'h42384d2a, 32'hc25faa42, 32'h42ab0329, 32'hc257b838};
test_weights[16440:16447] = '{32'hc2c109a6, 32'h40a74adc, 32'hc2b683f5, 32'h41972277, 32'hc25f6d6f, 32'h4254a8f4, 32'h41a92737, 32'hc2a26e90};
test_bias[2055:2055] = '{32'hc03a5cd0};
test_output[2055:2055] = '{32'hc5937003};
test_input[16448:16455] = '{32'hc209d71a, 32'h42608569, 32'h418b4a1f, 32'hc2868ea1, 32'h42c79c09, 32'h42268cf0, 32'hc27c50cc, 32'h421376c1};
test_weights[16448:16455] = '{32'h428d027a, 32'h42aba81c, 32'h4293ea4f, 32'hc21fa02b, 32'hc24cf10f, 32'h42694efc, 32'h422a7bd8, 32'h42bc518d};
test_bias[2056:2056] = '{32'h41153438};
test_output[2056:2056] = '{32'h458b9d81};
test_input[16456:16463] = '{32'hc2b04b82, 32'h42216fde, 32'hc2809bc5, 32'h428f275b, 32'hc26c03da, 32'hc2197532, 32'hc10795ad, 32'h41e57c1b};
test_weights[16456:16463] = '{32'h3fbd389b, 32'hc2a66fa7, 32'h409d5958, 32'hc1e2b0bc, 32'hc2b29bbb, 32'h429bb01b, 32'hbfa5ac03, 32'hbf89ddd4};
test_bias[2057:2057] = '{32'hc2988356};
test_output[2057:2057] = '{32'hc563eb00};
test_input[16464:16471] = '{32'h40f18630, 32'hc2361b00, 32'h42b5bea2, 32'h4200c3b1, 32'hc1ab6373, 32'hc28ca1a4, 32'h4243f692, 32'hc247b28a};
test_weights[16464:16471] = '{32'hc2c490fa, 32'hc2497213, 32'h41e5e16d, 32'hc22a63b3, 32'hc2808901, 32'hc2aaa9c8, 32'h4237ac6d, 32'hc2256320};
test_bias[2058:2058] = '{32'h42666660};
test_output[2058:2058] = '{32'h46632d43};
test_input[16472:16479] = '{32'h42a995ea, 32'h4299371e, 32'hc1b2a6cb, 32'h41a87b12, 32'hc2166609, 32'h428bfc5a, 32'hc2941ae0, 32'h426f25a1};
test_weights[16472:16479] = '{32'h418d8d61, 32'h41de8531, 32'h41c413c9, 32'h411d769e, 32'hc0bcab9f, 32'h42588ee8, 32'hc21df196, 32'hc2b66830};
test_bias[2059:2059] = '{32'hc2675fff};
test_output[2059:2059] = '{32'h45935cbf};
test_input[16480:16487] = '{32'hc2ac1c94, 32'hc2b21d70, 32'hc2b2cbe7, 32'hc1ada8a4, 32'hc0bde69c, 32'hc203f4fb, 32'h427f3224, 32'h3fc9cded};
test_weights[16480:16487] = '{32'h42c18218, 32'h42611b8a, 32'hc2b71c91, 32'h4250b550, 32'hc255b758, 32'h421fd995, 32'h4228585d, 32'h40d06dc6};
test_bias[2060:2060] = '{32'hc29d1aef};
test_output[2060:2060] = '{32'hc591f283};
test_input[16488:16495] = '{32'hc29518ca, 32'h428a1663, 32'hc2a6166a, 32'h40e6aae5, 32'h422b0527, 32'hc28a7467, 32'hc282183f, 32'hc1cabe8a};
test_weights[16488:16495] = '{32'hc2aa6a11, 32'hc2430e6e, 32'h4263d5bf, 32'hc176c7a7, 32'hc18d7cbf, 32'h42a508d5, 32'hc286c707, 32'hc216c53d};
test_bias[2061:2061] = '{32'h425cf55b};
test_output[2061:2061] = '{32'hc5372b63};
test_input[16496:16503] = '{32'h4259dc72, 32'hc2c40997, 32'h41edcb95, 32'h426291d6, 32'hc19ff378, 32'hc2a46836, 32'h421daef6, 32'hc1f624c4};
test_weights[16496:16503] = '{32'hc1fe0f4c, 32'hc2c40425, 32'h42002584, 32'hc1b07984, 32'h42890e97, 32'h4160579e, 32'h4182c617, 32'h41eadcbd};
test_bias[2062:2062] = '{32'h40621f58};
test_output[2062:2062] = '{32'h45960cfd};
test_input[16504:16511] = '{32'hc2c68e96, 32'h41b1e85b, 32'h4212efcd, 32'h3fcc8d96, 32'hc1871719, 32'hc15161ff, 32'h4197f1b3, 32'hc29a8b01};
test_weights[16504:16511] = '{32'h42c3e8eb, 32'h4086e998, 32'hc2a3302a, 32'h428dd0f0, 32'h428a9b0d, 32'h4294ad3a, 32'h4163ea3a, 32'h416971b7};
test_bias[2063:2063] = '{32'hc1c11822};
test_output[2063:2063] = '{32'hc672cc7d};
test_input[16512:16519] = '{32'hc1e1a0b2, 32'h4294f090, 32'h42614c7b, 32'h4020788f, 32'h3f96a048, 32'h42027256, 32'h41972575, 32'hc27c4128};
test_weights[16512:16519] = '{32'hc29d6479, 32'h42a0d998, 32'hc1c24e2a, 32'hc219fffa, 32'hc27cceec, 32'hc223b37b, 32'hc297c1bc, 32'h426d5285};
test_bias[2064:2064] = '{32'h41181cf6};
test_output[2064:2064] = '{32'h43297bd9};
test_input[16520:16527] = '{32'hc2b7311f, 32'h4117c275, 32'h4290ca14, 32'h41d5f4c6, 32'h42c0809b, 32'h4289f313, 32'h42c21313, 32'hc207eafe};
test_weights[16520:16527] = '{32'hc1e4ca90, 32'hc2978c07, 32'hc214eaea, 32'h42303f33, 32'hc2b89e38, 32'h4271536f, 32'hc289a9ba, 32'h427f64f4};
test_bias[2065:2065] = '{32'h42b058ca};
test_output[2065:2065] = '{32'hc64cb03e};
test_input[16528:16535] = '{32'hc2425963, 32'hc2866b7f, 32'hc11446ed, 32'hc21fbe61, 32'h40df635c, 32'hc241ae6d, 32'h428cab26, 32'hc262540b};
test_weights[16528:16535] = '{32'h42a13339, 32'hc19ba868, 32'h41aabd89, 32'hc20ed7b6, 32'hc24aa41a, 32'hc266d771, 32'h4018b2bd, 32'h40c35f42};
test_bias[2066:2066] = '{32'hc29cd5fb};
test_output[2066:2066] = '{32'h444924aa};
test_input[16536:16543] = '{32'hc29b89aa, 32'h427d314e, 32'h42a9aafe, 32'h4297213d, 32'hc1ede499, 32'h3f1c3d28, 32'hc2367279, 32'hbfb7e741};
test_weights[16536:16543] = '{32'h428ddc76, 32'hc208bce5, 32'hc1efb11d, 32'h41563796, 32'h410b6be9, 32'h41611bf7, 32'h4250bd33, 32'h3e262045};
test_bias[2067:2067] = '{32'hc2bffecc};
test_output[2067:2067] = '{32'hc63a8439};
test_input[16544:16551] = '{32'hc18fe653, 32'h427c5904, 32'hc2ba23c7, 32'h41a2c42e, 32'h41d170ee, 32'hc24ce8eb, 32'h41b5c154, 32'h4293f33f};
test_weights[16544:16551] = '{32'h42946f24, 32'h42a8b4d2, 32'hc25ec162, 32'h41a4aca7, 32'h423aac64, 32'h4039f42b, 32'hc1ad9a27, 32'hc27d3be5};
test_bias[2068:2068] = '{32'h42aa5aaa};
test_output[2068:2068] = '{32'h45ae11b7};
test_input[16552:16559] = '{32'hc256ecca, 32'hc20d932b, 32'hc2935070, 32'hc201148b, 32'h4230b50c, 32'hc2476781, 32'h42273c61, 32'h40007f1e};
test_weights[16552:16559] = '{32'hc270a023, 32'h419b4871, 32'hc2963c95, 32'h41536972, 32'hc05f508d, 32'hc258fed8, 32'h427eb948, 32'hc0ffbf49};
test_bias[2069:2069] = '{32'hc28d35c9};
test_output[2069:2069] = '{32'h4647a784};
test_input[16560:16567] = '{32'h41985a1e, 32'h42bcbbbb, 32'hc1130f5c, 32'hc1234821, 32'h422e0e5c, 32'hc26d95dc, 32'h412c652b, 32'hc2933df9};
test_weights[16560:16567] = '{32'hc20b0127, 32'h42a0db6f, 32'hc15109eb, 32'hc24abeb9, 32'h42c4358b, 32'h3e1109b7, 32'hc24bbb98, 32'hc192c4b4};
test_bias[2070:2070] = '{32'h4176a96c};
test_output[2070:2070] = '{32'h46458c72};
test_input[16568:16575] = '{32'hc2be8175, 32'hc25e8c15, 32'hc1273a76, 32'hc1b15d02, 32'hc1bd0471, 32'hc2c585ad, 32'hc2aa560b, 32'hc1a09b75};
test_weights[16568:16575] = '{32'hc2c21a64, 32'h423b2359, 32'h424638db, 32'hc2bd6311, 32'h4261b8d8, 32'hc13f9f85, 32'h428ede43, 32'hc2545b8d};
test_bias[2071:2071] = '{32'h41ec400e};
test_output[2071:2071] = '{32'h4540be79};
test_input[16576:16583] = '{32'hc22dd302, 32'h41ebcca9, 32'hc188c6fd, 32'hc1ce6e1f, 32'h420b9ad6, 32'h4227868a, 32'h421150a5, 32'hc0171bbb};
test_weights[16576:16583] = '{32'h42c2552e, 32'hc0caf473, 32'hc22a0b81, 32'h42ac3db3, 32'hc254e42c, 32'hc2780423, 32'hc28e78c6, 32'hc2b46c18};
test_bias[2072:2072] = '{32'h41a61c72};
test_output[2072:2072] = '{32'hc646a551};
test_input[16584:16591] = '{32'hc04149bf, 32'h42969e26, 32'hc2946a97, 32'hc29e1eb8, 32'h41ae59c3, 32'h4224c8da, 32'hc19a9e56, 32'hc1a9f2bc};
test_weights[16584:16591] = '{32'hc2706eca, 32'h4285de1a, 32'h41fb0094, 32'h425c5b41, 32'hc22b5480, 32'h423bbf0f, 32'h42815b73, 32'h422b7ca1};
test_bias[2073:2073] = '{32'hc2a43c89};
test_output[2073:2073] = '{32'hc5290362};
test_input[16592:16599] = '{32'h42aa6819, 32'h41d096cf, 32'h420163e8, 32'hc28a9749, 32'h42450772, 32'h42a358c0, 32'hc08793dd, 32'hc1c5a3c1};
test_weights[16592:16599] = '{32'hc04ebdc5, 32'hc296f774, 32'h4271de61, 32'h42bdb143, 32'hc28ce49c, 32'h42a4f179, 32'hc20f03ca, 32'h41957344};
test_bias[2074:2074] = '{32'hc15a021c};
test_output[2074:2074] = '{32'hc574dbdc};
test_input[16600:16607] = '{32'hc1e0fb83, 32'h41e4701f, 32'h40880a6f, 32'hc17f8474, 32'hc205e8b6, 32'h4275e857, 32'h412f413b, 32'hc29e49c7};
test_weights[16600:16607] = '{32'h40b1bfdf, 32'h42ba7d57, 32'hc19a5f4d, 32'hc2778722, 32'hc264f122, 32'hc21a16e7, 32'h42b0239a, 32'hc0c22020};
test_bias[2075:2075] = '{32'hc0851b2c};
test_output[2075:2075] = '{32'h45898872};
test_input[16608:16615] = '{32'hc152da2f, 32'h41cff22e, 32'h42951462, 32'hc18a886c, 32'h418358d5, 32'hc2b67628, 32'hc291e9ff, 32'h4293c091};
test_weights[16608:16615] = '{32'h425042b3, 32'h4283694a, 32'hc21abc18, 32'hc2712b68, 32'h42c6d588, 32'hc1991d07, 32'h42aa74e0, 32'hc20a2250};
test_bias[2076:2076] = '{32'hc251f003};
test_output[2076:2076] = '{32'hc5c3a7d3};
test_input[16616:16623] = '{32'hc18ed660, 32'hc101d466, 32'h41c5eca6, 32'hc2ac8f9b, 32'h405d863d, 32'hc2ab58e7, 32'hc2c67b1e, 32'h42a80181};
test_weights[16616:16623] = '{32'hc25d0750, 32'hc24316c7, 32'h421c77f0, 32'h40133406, 32'h42a0b999, 32'h42c6664a, 32'hc2994836, 32'hc2c0bc33};
test_bias[2077:2077] = '{32'hc2a15c21};
test_output[2077:2077] = '{32'hc5cf7746};
test_input[16624:16631] = '{32'hc22e784c, 32'h428bf3e0, 32'hc10bef16, 32'h4231ec50, 32'hc2bef58f, 32'h40964dc0, 32'h42a4ee0b, 32'h4183f68b};
test_weights[16624:16631] = '{32'hc2893d12, 32'hc2af5ea4, 32'h41df966e, 32'h4286dae2, 32'hc12d12a4, 32'hc19e0d0c, 32'h40216396, 32'h42846e75};
test_bias[2078:2078] = '{32'h42a2260c};
test_output[2078:2078] = '{32'h44f1a72a};
test_input[16632:16639] = '{32'hc1220b1c, 32'h41402364, 32'h424c00d1, 32'h428c10b9, 32'hc1d33dea, 32'h429973c3, 32'hc275d6e3, 32'hc1a3235a};
test_weights[16632:16639] = '{32'hc26e8f6d, 32'h41c77bd8, 32'h40ad366e, 32'hc2a06844, 32'hc24ab1d4, 32'h42c6b9c3, 32'h42451835, 32'h40c0b170};
test_bias[2079:2079] = '{32'hc138f85d};
test_output[2079:2079] = '{32'h44aa36b7};
test_input[16640:16647] = '{32'hc1ee6286, 32'hc2c5da6a, 32'h42ab01bb, 32'hc1a3fba1, 32'h42af58ec, 32'h420bafef, 32'h4193ec5b, 32'hc2885773};
test_weights[16640:16647] = '{32'h42ba6930, 32'hc2bfd6ad, 32'h42ac3420, 32'h419885eb, 32'h429a82cb, 32'h4218d8fe, 32'hbfcadc4e, 32'hc2b386b4};
test_bias[2080:2080] = '{32'h41446160};
test_output[2080:2080] = '{32'h46d9e96b};
test_input[16648:16655] = '{32'h4235e97b, 32'hc193e4b2, 32'hc1c06793, 32'hc2695d87, 32'h429d427a, 32'h42724319, 32'h41a63c28, 32'h4198c36d};
test_weights[16648:16655] = '{32'hc26932f6, 32'h42790d7f, 32'h429ce62c, 32'h419d3597, 32'hc29a53e0, 32'h41a0fe54, 32'hc2997fec, 32'h42b4bcb3};
test_bias[2081:2081] = '{32'hc2a1c8a5};
test_output[2081:2081] = '{32'hc635c905};
test_input[16656:16663] = '{32'hc29fac3f, 32'hc2811675, 32'h42610f77, 32'hc1c417fe, 32'h424c074c, 32'h424a5266, 32'h417e728e, 32'hc22917bb};
test_weights[16656:16663] = '{32'h428f9826, 32'h426650ec, 32'hc285431a, 32'h42634d9e, 32'h41c82bac, 32'h42c16dc0, 32'h42bb87db, 32'hc203d7a1};
test_bias[2082:2082] = '{32'h418cba54};
test_output[2082:2082] = '{32'hc5ac80bf};
test_input[16664:16671] = '{32'hc28c371e, 32'h41ea1b69, 32'h3ff9ef5f, 32'h4110bea7, 32'hc21e6a99, 32'h418c298f, 32'hc15a3248, 32'h42b433a1};
test_weights[16664:16671] = '{32'hc2b84b71, 32'hc2c3d4a2, 32'hc29a627b, 32'hc1eedc04, 32'hc29192b9, 32'hc20446cf, 32'h420af90e, 32'h425c144c};
test_bias[2083:2083] = '{32'h4217963f};
test_output[2083:2083] = '{32'h461c3b08};
test_input[16672:16679] = '{32'hc2796ec7, 32'hc25a22e6, 32'hc2965488, 32'h42c24a53, 32'h41cc5dda, 32'hc1efc1bc, 32'h410b04e3, 32'hc106401e};
test_weights[16672:16679] = '{32'hc0ef00b4, 32'hc19c4dca, 32'hc27f98d1, 32'h42533892, 32'hc1947388, 32'h41cc41f7, 32'hc22e9fb3, 32'hc1d9761a};
test_bias[2084:2084] = '{32'hc21e47b1};
test_output[2084:2084] = '{32'h461cc7db};
test_input[16680:16687] = '{32'h42ae8c08, 32'hc297a46d, 32'h42091cbc, 32'hc1f729dc, 32'h4245a7be, 32'hc20153dc, 32'hc14bb13c, 32'hc1891e33};
test_weights[16680:16687] = '{32'h40f45874, 32'hc29c1a7a, 32'hc254f72b, 32'hc212bee6, 32'h42a60f85, 32'hc2b056bf, 32'h4292463c, 32'hc2bae1c3};
test_bias[2085:2085] = '{32'h4028fc65};
test_output[2085:2085] = '{32'h46533dbd};
test_input[16688:16695] = '{32'hc28a9305, 32'h429d7ea6, 32'h421b1cd2, 32'hc20b3dcb, 32'hc2706bf4, 32'h42b36a7b, 32'hc2447292, 32'hc2166fdf};
test_weights[16688:16695] = '{32'h42b48ca2, 32'hc1faf47c, 32'hc2b092d5, 32'h42840cc0, 32'h411b6b4f, 32'h422023ec, 32'hc1a547bc, 32'h418cac5c};
test_bias[2086:2086] = '{32'h42b0a6db};
test_output[2086:2086] = '{32'hc62bd739};
test_input[16696:16703] = '{32'h42b286f7, 32'hc2afe30d, 32'hc283a0c9, 32'hc2b129b7, 32'h41498819, 32'h42c5c3a4, 32'hc207d1cf, 32'h421b03fd};
test_weights[16696:16703] = '{32'hc1d4077d, 32'hc204fbfd, 32'h42c6672f, 32'hc216a60a, 32'hc236f99d, 32'h40fcfae2, 32'hc29a77ea, 32'hbef279d3};
test_bias[2087:2087] = '{32'hc0d79376};
test_output[2087:2087] = '{32'h43283786};
test_input[16704:16711] = '{32'hc22a51f9, 32'hc26b702b, 32'hc26dcd02, 32'hc2aafad1, 32'h40d3f49c, 32'h42b41978, 32'h41c77b77, 32'hc2aff0e6};
test_weights[16704:16711] = '{32'hc204c9f3, 32'h422b2e09, 32'h41b2b699, 32'h427217c6, 32'hc10d29d9, 32'hc263f5d3, 32'hc2b0ee67, 32'h42ac4126};
test_bias[2088:2088] = '{32'hc1ec2087};
test_output[2088:2088] = '{32'hc6b0a405};
test_input[16712:16719] = '{32'h42a2890d, 32'h4250e558, 32'hc22d97cd, 32'h4246fd98, 32'h4250eac6, 32'hc2c3d651, 32'hc2344c2d, 32'hc29c3cbc};
test_weights[16712:16719] = '{32'h41e95503, 32'h41691929, 32'hc1250a02, 32'hc06b63d1, 32'h42b1526b, 32'h429e5c1a, 32'hc23f9d46, 32'hc2b57755};
test_bias[2089:2089] = '{32'h4261fc6a};
test_output[2089:2089] = '{32'h4615a3f2};
test_input[16720:16727] = '{32'h42b86972, 32'hc2a6dfc1, 32'hc28b177f, 32'h4258d5e1, 32'h428747fd, 32'hc19dcb51, 32'hc16d8404, 32'h42187d2e};
test_weights[16720:16727] = '{32'h41a9aea7, 32'hc291967a, 32'h42819c0d, 32'h42350cc9, 32'h42c215f4, 32'h41e705a6, 32'hc29d9d8c, 32'h42adb950};
test_bias[2090:2090] = '{32'hc2a58e44};
test_output[2090:2090] = '{32'h467fc43f};
test_input[16728:16735] = '{32'h42a54c89, 32'h42811536, 32'h4206def3, 32'h428e901a, 32'h414e6b51, 32'h428d7d74, 32'h4256d9d5, 32'h423d5ffd};
test_weights[16728:16735] = '{32'hc29f2904, 32'h423fea8d, 32'hbf115354, 32'hc29be557, 32'hc2329fe5, 32'h42c485e1, 32'hc254cfa5, 32'h42a2cd4b};
test_bias[2091:2091] = '{32'h427d0484};
test_output[2091:2091] = '{32'hc4caa627};
test_input[16736:16743] = '{32'hc1a4f451, 32'h42a2b914, 32'hc2977f05, 32'hc25afc5a, 32'hc2c75a3f, 32'h42235843, 32'hc2c227aa, 32'hc1b50127};
test_weights[16736:16743] = '{32'hc29496d8, 32'hc2ab5e5d, 32'hbf9f6a4d, 32'hc10077a6, 32'hc2bcf12a, 32'h41d6e6ea, 32'h42443d06, 32'hc2850a52};
test_bias[2092:2092] = '{32'h42a17b88};
test_output[2092:2092] = '{32'h4517f1e2};
test_input[16744:16751] = '{32'hc23d3145, 32'hc264be36, 32'h42515bdb, 32'h42a10c5f, 32'hc1e1b52f, 32'hc2c79d60, 32'h42545678, 32'h4286eb02};
test_weights[16744:16751] = '{32'hc2788655, 32'hc2c454e1, 32'h424ab390, 32'hc29e486b, 32'h3f9478c9, 32'h42893a30, 32'h42a56a43, 32'hc2c50a18};
test_bias[2093:2093] = '{32'hc24c4f09};
test_output[2093:2093] = '{32'hc5881cd1};
test_input[16752:16759] = '{32'hc2721806, 32'hc1ee0fbd, 32'h41413734, 32'h429fd424, 32'h42083671, 32'hc23c91e7, 32'hc2a65691, 32'h42c4b251};
test_weights[16752:16759] = '{32'h4286c491, 32'hc0acd071, 32'h42aebb1a, 32'h4180ab13, 32'h4235d79d, 32'h421c3c0a, 32'hc29321fe, 32'h42bc7a88};
test_bias[2094:2094] = '{32'h4251a619};
test_output[2094:2094] = '{32'h46540276};
test_input[16760:16767] = '{32'h421f65c3, 32'h40b31373, 32'hc2a608ad, 32'h42c0e124, 32'hc2c2be57, 32'hc2b5489f, 32'hc29e7195, 32'hc2c4f26d};
test_weights[16760:16767] = '{32'hc2a4c87e, 32'hc224f937, 32'h41e9c878, 32'hc20e136b, 32'h42aa3d97, 32'h41de13ba, 32'hc195a73e, 32'h42024f45};
test_bias[2095:2095] = '{32'h42b9a438};
test_output[2095:2095] = '{32'hc6aa5667};
test_input[16768:16775] = '{32'hc22bcb9c, 32'hc295ed06, 32'h41721030, 32'h42af77b1, 32'h410c7493, 32'hc22054d3, 32'hc20861f2, 32'h42bc5f98};
test_weights[16768:16775] = '{32'hc2be0c5f, 32'hc1ae1971, 32'hc2652149, 32'hc23a8a1f, 32'h42409425, 32'h41ace686, 32'h42aecb1d, 32'hc21170a3};
test_bias[2096:2096] = '{32'hc1cc4beb};
test_output[2096:2096] = '{32'hc5bf3990};
test_input[16776:16783] = '{32'h419a332e, 32'hc26fdf14, 32'h42a58029, 32'hc277909e, 32'h41b425b2, 32'h3bc75af3, 32'h426e0bfc, 32'hc124d30c};
test_weights[16776:16783] = '{32'h42702ceb, 32'h4264192f, 32'hc2827329, 32'hc00aa172, 32'h41c32310, 32'hc251e150, 32'hc007a472, 32'h4182c847};
test_bias[2097:2097] = '{32'h42637fbd};
test_output[2097:2097] = '{32'hc5e1729e};
test_input[16784:16791] = '{32'h41444ccb, 32'h42970d80, 32'hc2c2e0ed, 32'hc1b831e6, 32'h42419647, 32'h40f0fce8, 32'hc27d621b, 32'h42a54cce};
test_weights[16784:16791] = '{32'hc2b5a82b, 32'hc242177d, 32'h42209a46, 32'hc26f3efa, 32'h42946e0d, 32'h401cbeb7, 32'hc239a410, 32'hc2206fa3};
test_bias[2098:2098] = '{32'h424d9212};
test_output[2098:2098] = '{32'hc57bbc32};
test_input[16792:16799] = '{32'hc234a822, 32'h4285eeb7, 32'hc2508bf7, 32'hc254389c, 32'h42b775c4, 32'h42b3a32e, 32'hc2afdfe3, 32'hc281b6b0};
test_weights[16792:16799] = '{32'h42764ca0, 32'hc28ba04a, 32'h42a8c6dc, 32'h42539068, 32'h42853a30, 32'h4187990c, 32'hc265a87c, 32'h424f9c0e};
test_bias[2099:2099] = '{32'h42233d7b};
test_output[2099:2099] = '{32'hc5a5cd1a};
test_input[16800:16807] = '{32'h4272144e, 32'h4290fd96, 32'hc28d4fd6, 32'hc249b295, 32'hc2728527, 32'h41e5c852, 32'hc1a334fe, 32'hc180908b};
test_weights[16800:16807] = '{32'h42c20295, 32'hc28dbf97, 32'h42908459, 32'hc29cb25a, 32'h4270320b, 32'hc2a73d84, 32'h41ebf7dd, 32'h42afed05};
test_bias[2100:2100] = '{32'h42375045};
test_output[2100:2100] = '{32'hc603c8f8};
test_input[16808:16815] = '{32'h428edc6e, 32'h42051fbd, 32'hc089aef0, 32'h42961688, 32'hc2639257, 32'hc0e5d3f0, 32'h42b59935, 32'h422f3fc1};
test_weights[16808:16815] = '{32'hc120bd3a, 32'h42bb6987, 32'hc12b4930, 32'h420db546, 32'h429bd9b6, 32'h40090e5c, 32'hc2a76f2b, 32'h425a91ab};
test_bias[2101:2101] = '{32'hc2b8328a};
test_output[2101:2101] = '{32'hc591152d};
test_input[16816:16823] = '{32'hc22b14dd, 32'h4187c8cf, 32'h42a49eed, 32'hc2a2960a, 32'h422997ed, 32'h42184870, 32'h426119e4, 32'hc21fb260};
test_weights[16816:16823] = '{32'hc276f73e, 32'hc2b152ea, 32'hc2b1cb3d, 32'hc1aef84c, 32'h42409bdd, 32'h42983d6b, 32'hc2a237b4, 32'h4244d931};
test_bias[2102:2102] = '{32'h42902073};
test_output[2102:2102] = '{32'hc5b90753};
test_input[16824:16831] = '{32'h42abc6e2, 32'h4227518a, 32'hc29a87c2, 32'h427b8903, 32'hc287a1aa, 32'h420d3a1a, 32'hc192b51b, 32'hc28fe511};
test_weights[16824:16831] = '{32'hc117adc4, 32'hc2815bc0, 32'h40bace3d, 32'h422c6b0c, 32'h41000943, 32'h425ddd95, 32'h418699c0, 32'hc1d10067};
test_bias[2103:2103] = '{32'h429dec9c};
test_output[2103:2103] = '{32'h44e1b0a3};
test_input[16832:16839] = '{32'h42bbc81c, 32'hc180dd52, 32'hc1e24072, 32'h418fbc2b, 32'h4241e844, 32'h40487aa5, 32'hc28b2391, 32'h42a48966};
test_weights[16832:16839] = '{32'h42b570b3, 32'hc2ab3446, 32'hc2ba64a6, 32'h42152a19, 32'h4292995e, 32'hc25cd940, 32'hc264fe4f, 32'hc24a7c76};
test_bias[2104:2104] = '{32'hc2425a51};
test_output[2104:2104] = '{32'h467f818e};
test_input[16840:16847] = '{32'hc26ddb6c, 32'hc1a42258, 32'hc2903344, 32'h4010c97b, 32'hc1929ea5, 32'hc2059985, 32'h41b9b0b0, 32'hc2328737};
test_weights[16840:16847] = '{32'hc2c75b79, 32'hc2328028, 32'h4279c048, 32'hc19df707, 32'hc17c7103, 32'h422f0908, 32'hc1a2f1bc, 32'h414b2b72};
test_bias[2105:2105] = '{32'hc0fa685b};
test_output[2105:2105] = '{32'h42997481};
test_input[16848:16855] = '{32'h420f35b2, 32'h42a2792d, 32'hc1e41266, 32'hc24c477d, 32'h421453e7, 32'h4294b116, 32'h42c62ee5, 32'h42c00cf8};
test_weights[16848:16855] = '{32'hc22074be, 32'hc191945a, 32'h42447897, 32'hc0a740db, 32'h42084d7b, 32'h42bc7596, 32'hc0a0d20c, 32'h42a0d281};
test_bias[2106:2106] = '{32'hc208f364};
test_output[2106:2106] = '{32'h46324a63};
test_input[16856:16863] = '{32'h4186a12f, 32'hc211ea6a, 32'hc1325711, 32'hc1f5f40c, 32'hc282fb4d, 32'hc28b44ad, 32'hc28f32eb, 32'h3d502c5c};
test_weights[16856:16863] = '{32'h42c44f84, 32'h420162e8, 32'h429d1fcd, 32'hc2b95d33, 32'hc1e724c7, 32'hc1f01095, 32'hc006c404, 32'hc0c1b8c6};
test_bias[2107:2107] = '{32'h42c31b4c};
test_output[2107:2107] = '{32'h45d09b87};
test_input[16864:16871] = '{32'h42a248a1, 32'hc22341ac, 32'hc2b8c36d, 32'hc29ab866, 32'hc1b8d3d9, 32'h40eb73ba, 32'h422698d0, 32'hc1722d5f};
test_weights[16864:16871] = '{32'h42328a7b, 32'hc26ebe87, 32'hc29a5dde, 32'hc2c790ce, 32'hc23c15e4, 32'h428f4fca, 32'h41e5c8bc, 32'hc283990d};
test_bias[2108:2108] = '{32'h4223e742};
test_output[2108:2108] = '{32'h46c16451};
test_input[16872:16879] = '{32'h42539819, 32'h4192d982, 32'h428d704e, 32'hc2929684, 32'h411a2ce9, 32'hbf5e5225, 32'hc23c274d, 32'h42a297b6};
test_weights[16872:16879] = '{32'hc1d706c4, 32'hc17a1e02, 32'hc21f7a6d, 32'hc18bb645, 32'h4142f465, 32'hc26a3473, 32'hc293e4cb, 32'h41a63cc7};
test_bias[2109:2109] = '{32'hc11dd3b5};
test_output[2109:2109] = '{32'h4501dbb2};
test_input[16880:16887] = '{32'h428de47e, 32'hc2536a7b, 32'h4296fdbf, 32'h42c02e32, 32'hc104740f, 32'h40e6b15e, 32'h4233c686, 32'hc120995a};
test_weights[16880:16887] = '{32'hc2891661, 32'h42441ce8, 32'hc2453aec, 32'hc21b5d1f, 32'h427fe9b4, 32'hc1aa3e2c, 32'h420f141c, 32'h41a4514d};
test_bias[2110:2110] = '{32'hc1692ef4};
test_output[2110:2110] = '{32'hc65df49f};
test_input[16888:16895] = '{32'h41dea198, 32'h4291535d, 32'hc276e5e2, 32'h426ce73b, 32'hc21c4787, 32'hc2b0daf9, 32'h4245cd75, 32'h41022be3};
test_weights[16888:16895] = '{32'hc2917f1a, 32'h419001e3, 32'hc28c47fd, 32'hc046cae3, 32'h426c3b63, 32'h429d389e, 32'hc0608ee1, 32'h41ab9c96};
test_bias[2111:2111] = '{32'hc1d87230};
test_output[2111:2111] = '{32'hc5b6feda};
test_input[16896:16903] = '{32'hc17e3401, 32'hc1c25310, 32'h4295ba30, 32'hc246c8dd, 32'hc2487788, 32'hc1c13fc0, 32'hc250b28e, 32'h429dbc92};
test_weights[16896:16903] = '{32'h41b9c762, 32'hc2c28cfb, 32'h42928ea8, 32'hc1788aa5, 32'h41818c4f, 32'hc00bf273, 32'h42244fdc, 32'hc2a30978};
test_bias[2112:2112] = '{32'h426a826e};
test_output[2112:2112] = '{32'hc47f3098};
test_input[16904:16911] = '{32'h3f99f2bb, 32'hc1255640, 32'hc28785fe, 32'h42bffc90, 32'h418d8722, 32'hc26e380f, 32'h424ee8f5, 32'h42856ec4};
test_weights[16904:16911] = '{32'hc1c67db7, 32'h410a7840, 32'hc1f056c9, 32'hc21c3123, 32'hc261d082, 32'hc26e670b, 32'hc20fcdd5, 32'h42901e34};
test_bias[2113:2113] = '{32'h42a97459};
test_output[2113:2113] = '{32'h456a7785};
test_input[16912:16919] = '{32'hc2523170, 32'h423d334b, 32'h42c604da, 32'hc1c1a8ea, 32'hc14ba14d, 32'hc0b1f1b6, 32'h42641cec, 32'hc2b85a14};
test_weights[16912:16919] = '{32'h4282dcb1, 32'hc29d4153, 32'hc2703b3c, 32'h4287f429, 32'hc2823892, 32'h41b70812, 32'h42411c79, 32'h3f952017};
test_bias[2114:2114] = '{32'h42a68d7a};
test_output[2114:2114] = '{32'hc630dad7};
test_input[16920:16927] = '{32'h4200239b, 32'hc1c78e65, 32'hbf832742, 32'h42197825, 32'hc2c3e1ff, 32'hc2282635, 32'hc2609d2e, 32'hc29f10a7};
test_weights[16920:16927] = '{32'hc048ad72, 32'h428f6ebd, 32'hc2a54fb0, 32'h41b7855f, 32'h42839432, 32'hc2871aab, 32'h42111b8e, 32'h4294abd7};
test_bias[2115:2115] = '{32'hc21a1a8a};
test_output[2115:2115] = '{32'hc6439026};
test_input[16928:16935] = '{32'h40d8d1ba, 32'hc281ec1b, 32'hc22f26ec, 32'hc2926251, 32'hc13066e7, 32'hc2ba8ec7, 32'hc2b7df71, 32'h4241dffa};
test_weights[16928:16935] = '{32'hc0a19a73, 32'hc10541ca, 32'hc2c7d102, 32'hc0da91d3, 32'hc2a58198, 32'h42b7ea34, 32'h423c3f30, 32'h42b8ada8};
test_bias[2116:2116] = '{32'h42b459e8};
test_output[2116:2116] = '{32'hc4ff97e5};
test_input[16936:16943] = '{32'hc2a335cc, 32'h426b9716, 32'hc0996650, 32'h41538f28, 32'hc2c52d78, 32'h429fc0fd, 32'hc26efdee, 32'hc2b09fbf};
test_weights[16936:16943] = '{32'h42af0ebf, 32'hc2962dee, 32'hc2272f47, 32'h3fdb187a, 32'h42a65d18, 32'h42aef5b3, 32'hc21b1f3a, 32'hc1d8416a};
test_bias[2117:2117] = '{32'h41c497eb};
test_output[2117:2117] = '{32'hc5f49596};
test_input[16944:16951] = '{32'h424f2dec, 32'h426cf75b, 32'hc252ca77, 32'h4285f851, 32'hc19bda6a, 32'hc27290d6, 32'h4285e08b, 32'hc2a2ef3d};
test_weights[16944:16951] = '{32'hc1e28617, 32'hc15597c4, 32'h414592be, 32'h4281ccce, 32'hc27c2c9b, 32'h42a2b2c2, 32'h416d7e8b, 32'h41da0e6f};
test_bias[2118:2118] = '{32'hc28f6f8d};
test_output[2118:2118] = '{32'hc55ec760};
test_input[16952:16959] = '{32'h428de1cd, 32'hc258beb2, 32'hc2807a76, 32'hc21eb185, 32'hc289ef86, 32'hc25274e5, 32'h41d8096f, 32'h4278b605};
test_weights[16952:16959] = '{32'h42b2f8d7, 32'hc2be22c3, 32'h419f5111, 32'hc2c15491, 32'hc2990dba, 32'h419e07b8, 32'hc29cf80d, 32'h42923762};
test_bias[2119:2119] = '{32'hc09773e8};
test_output[2119:2119] = '{32'h46a1d6d7};
test_input[16960:16967] = '{32'h428357ae, 32'hc2ac5820, 32'h428fab94, 32'hc188fe58, 32'h41836fe5, 32'h41063ee3, 32'h4277c6fd, 32'h4012d5d4};
test_weights[16960:16967] = '{32'h426b1c96, 32'hc28eaa5d, 32'hc1e06acc, 32'hc28b7250, 32'hc250ffd7, 32'hc28174d0, 32'hc2420aa5, 32'hc2aba881};
test_bias[2120:2120] = '{32'hc2784302};
test_output[2120:2120] = '{32'h458d422f};
test_input[16968:16975] = '{32'hbf519858, 32'hc25b444f, 32'hc1138e5a, 32'h42518f5d, 32'hc14efe42, 32'h42990587, 32'hc1363715, 32'hc245a55c};
test_weights[16968:16975] = '{32'h424ef623, 32'hc2459ac1, 32'hc286f856, 32'h42847872, 32'hc23c34fa, 32'h412b24d4, 32'h412106c9, 32'h423a49de};
test_bias[2121:2121] = '{32'hc28b9ec9};
test_output[2121:2121] = '{32'h45b21c7a};
test_input[16976:16983] = '{32'h41904269, 32'h424fe6da, 32'hc2a71df7, 32'h40d04c9c, 32'hc1a954ca, 32'hc2813c10, 32'hc117780e, 32'hc225ded4};
test_weights[16976:16983] = '{32'h421cdbe2, 32'h42a7287d, 32'h41e08c6f, 32'h41c589ed, 32'h4288d265, 32'hc295c660, 32'h42bc406f, 32'hc29779c4};
test_bias[2122:2122] = '{32'hc2b1ea99};
test_output[2122:2122] = '{32'h460388d5};
test_input[16984:16991] = '{32'h4182e259, 32'h4115d5e7, 32'hc21223f5, 32'h3ee68fff, 32'hc2c6997f, 32'hc2bde958, 32'hc2059cc8, 32'h42b4f822};
test_weights[16984:16991] = '{32'hc2872585, 32'hc1a099ce, 32'h428597be, 32'h4240c376, 32'h41f6cd4f, 32'h4247a275, 32'h3f90bf40, 32'hc2928d34};
test_bias[2123:2123] = '{32'hbfab7075};
test_output[2123:2123] = '{32'hc68e1074};
test_input[16992:16999] = '{32'hc2c013f3, 32'h41a2cb03, 32'hc28123f6, 32'h41d38369, 32'h40674b55, 32'hc1805b00, 32'h42a6361b, 32'hc1965ae8};
test_weights[16992:16999] = '{32'hc23baf43, 32'hc0246718, 32'hc2b6e91d, 32'hc1fa783b, 32'h4235fc60, 32'h41a22e8c, 32'h417aaf3d, 32'hc11b8923};
test_bias[2124:2124] = '{32'h4188e936};
test_output[2124:2124] = '{32'h4629e238};
test_input[17000:17007] = '{32'h424d6ff9, 32'h401e17c9, 32'h41f83496, 32'hc29a5ef6, 32'h41e44d2c, 32'h41be8e0e, 32'hc287392e, 32'h3fba2d8e};
test_weights[17000:17007] = '{32'hc1def8be, 32'hc0dac439, 32'hc1a259b1, 32'h42c0ed7e, 32'hc211f691, 32'h4270601c, 32'h42b5a22f, 32'hc195b34e};
test_bias[2125:2125] = '{32'h428c1e93};
test_output[2125:2125] = '{32'hc66dfbec};
test_input[17008:17015] = '{32'h421f838f, 32'h4228ae2d, 32'hc2ad406a, 32'h42315cea, 32'h40f8593d, 32'hc1b112e3, 32'h42b08004, 32'hc18ef42e};
test_weights[17008:17015] = '{32'hc22c9230, 32'h4282b869, 32'hc1f3ebec, 32'h42040edc, 32'hc2bf4161, 32'hc28ca603, 32'h4290cf15, 32'h429e6945};
test_bias[2126:2126] = '{32'hc2b22632};
test_output[2126:2126] = '{32'h46296263};
test_input[17016:17023] = '{32'hc280c1e8, 32'h42acc7a6, 32'h42022684, 32'hc149ac2d, 32'hc206b320, 32'h4299a432, 32'h41f223a1, 32'h42885cd8};
test_weights[17016:17023] = '{32'hc1522437, 32'h403b3019, 32'h425174a1, 32'h41b20411, 32'hc2414446, 32'h41ce4222, 32'h42065c63, 32'h41c7f467};
test_bias[2127:2127] = '{32'hc242cbf4};
test_output[2127:2127] = '{32'h46098561};
test_input[17024:17031] = '{32'h42396090, 32'hc02f2663, 32'hc29dbb9d, 32'hc2ba3354, 32'h42917af1, 32'hc19f226b, 32'h417f8642, 32'hc2c56499};
test_weights[17024:17031] = '{32'hc2961cca, 32'hc218dcaa, 32'h42665796, 32'hc103aa9d, 32'hc2143107, 32'h42b4e443, 32'hc29c62f0, 32'hc24838bd};
test_bias[2128:2128] = '{32'h424f1f9c};
test_output[2128:2128] = '{32'hc5f6dfb8};
test_input[17032:17039] = '{32'hc2692426, 32'h42c636c6, 32'h3f8ddc34, 32'hc28efa6f, 32'hc2c4d0a0, 32'hc20dc5d0, 32'h41f3b438, 32'h41fb205b};
test_weights[17032:17039] = '{32'h416a7cde, 32'h42157744, 32'hc2263993, 32'hc1c18d0f, 32'h4286ac8d, 32'hc1fdf9c4, 32'h42bf316f, 32'hc24310cb};
test_bias[2129:2129] = '{32'h41578f25};
test_output[2129:2129] = '{32'h43d51777};
test_input[17040:17047] = '{32'hc25bb3e6, 32'hc2ae1a46, 32'h417a8fb6, 32'h423c1b62, 32'h4268f09d, 32'hc277da5e, 32'hc1db8e5f, 32'hc2c522d2};
test_weights[17040:17047] = '{32'hc2060520, 32'hc25c097b, 32'hc2763a66, 32'h40b93dfe, 32'hc29ab099, 32'h429e16c4, 32'h427e2bea, 32'hc2960278};
test_bias[2130:2130] = '{32'h42931dda};
test_output[2130:2130] = '{32'h450d1da7};
test_input[17048:17055] = '{32'h425d6c51, 32'h423ec09e, 32'h4010c3b9, 32'hc2ac7f7b, 32'h42a90b55, 32'h4291a77b, 32'h42aa8535, 32'hc23ea934};
test_weights[17048:17055] = '{32'h423e8326, 32'hc287d1cb, 32'h420791f7, 32'hc24d4719, 32'h4101148f, 32'hc1fe3f14, 32'h42af36fd, 32'h404b7fdf};
test_bias[2131:2131] = '{32'h426819fd};
test_output[2131:2131] = '{32'h4616b0ba};
test_input[17056:17063] = '{32'h420bf797, 32'hc2c55a49, 32'h423d38e7, 32'hc2573701, 32'h427054ea, 32'h42a0e8a7, 32'hbf3508bd, 32'hbfefcbd2};
test_weights[17056:17063] = '{32'h42677e56, 32'hc2acee6e, 32'h4004fd23, 32'hc2bf9ac6, 32'hc2c0e16e, 32'h426de2f0, 32'hc2034d16, 32'hc1ffb5e3};
test_bias[2132:2132] = '{32'hc1f0c031};
test_output[2132:2132] = '{32'h46681578};
test_input[17064:17071] = '{32'h4289e088, 32'hc2b44ccf, 32'hc1e57f63, 32'hbfa82261, 32'h422f68a5, 32'h41c65278, 32'hc1b3b17d, 32'h42c3ccf7};
test_weights[17064:17071] = '{32'h4281ca0b, 32'h428e8ebe, 32'h429d7b24, 32'hc2a2e3a6, 32'hc1b6ca78, 32'hc256c291, 32'h42ac787d, 32'h4215045e};
test_bias[2133:2133] = '{32'h419185a8};
test_output[2133:2133] = '{32'hc59323b7};
test_input[17072:17079] = '{32'hc28e2530, 32'hc19a00b1, 32'hc133e5c4, 32'h42beee8d, 32'h416256f1, 32'hc252bee3, 32'hc289cc8b, 32'hc1a52ee8};
test_weights[17072:17079] = '{32'hc2a60272, 32'hbf4c2719, 32'h3fb31c2e, 32'h40bbf12c, 32'hc0e85fb6, 32'h42b3f0b1, 32'hc1d71047, 32'hc2ae1cfd};
test_bias[2134:2134] = '{32'hc245eaae};
test_output[2134:2134] = '{32'h45a30839};
test_input[17080:17087] = '{32'hc1b3e55d, 32'h42978f63, 32'hc1aadb5b, 32'hc22b6a11, 32'hc2b2ace2, 32'h428eddf3, 32'h429d8b1c, 32'h42ab0349};
test_weights[17080:17087] = '{32'hc2144647, 32'hc2a03dbe, 32'h42adfb16, 32'h428d1778, 32'hc212177b, 32'h422cbcc0, 32'hc1a6f801, 32'hc2be3d03};
test_bias[2135:2135] = '{32'h418abd20};
test_output[2135:2135] = '{32'hc6536d41};
test_input[17088:17095] = '{32'h3fb321f9, 32'h41da5196, 32'hc0f2d22c, 32'hc2743642, 32'h4280fd8d, 32'h418e0aa8, 32'hc267543e, 32'hc2a3a61d};
test_weights[17088:17095] = '{32'h41724c8e, 32'h41f3b090, 32'h42775f44, 32'hc1cc7676, 32'hc202840b, 32'h42a4c10c, 32'hc27e5f98, 32'h429ded62};
test_bias[2136:2136] = '{32'hc1ec05a9};
test_output[2136:2136] = '{32'hc4bce3c2};
test_input[17096:17103] = '{32'h41e8d2c8, 32'hc2bb3360, 32'h42869a7e, 32'hc17d9025, 32'h41f468a7, 32'h40dc269b, 32'h420acbf1, 32'hc20a6e8e};
test_weights[17096:17103] = '{32'h4283016e, 32'h41d8c897, 32'h41423617, 32'h4178aa2f, 32'hc2683ccb, 32'hc211a54d, 32'h42a6f149, 32'hc1eafd88};
test_bias[2137:2137] = '{32'h41b43a67};
test_output[2137:2137] = '{32'h44e778af};
test_input[17104:17111] = '{32'h42bb4367, 32'hc1bdf171, 32'hc2afbe36, 32'h429c6af6, 32'hc1af4fb7, 32'h42276e54, 32'hc1c0cffb, 32'hc2209b39};
test_weights[17104:17111] = '{32'h4002d0c7, 32'hc225c5ff, 32'hc22cc0ec, 32'h42a94c95, 32'h42a94025, 32'h4231541c, 32'hc1a7f22e, 32'hc25bfeaf};
test_bias[2138:2138] = '{32'hc0dbeca7};
test_output[2138:2138] = '{32'h465f6d35};
test_input[17112:17119] = '{32'hc295637b, 32'h4291e194, 32'h42628a77, 32'hc0149a25, 32'hc24bc262, 32'hc2a2e266, 32'h418deba4, 32'hc29bf1c1};
test_weights[17112:17119] = '{32'hc1c6aeb7, 32'h429899fb, 32'hc29fdda9, 32'hc13770af, 32'h42ae65a0, 32'hc1b702b3, 32'h42b8abb0, 32'hc294b6b1};
test_bias[2139:2139] = '{32'hc29b0d0c};
test_output[2139:2139] = '{32'h45f09c93};
test_input[17120:17127] = '{32'h4255d570, 32'hc265ea1d, 32'h429554b9, 32'hc1c6433a, 32'h41bdd73f, 32'h42adae5f, 32'h423b5e8b, 32'hc2364f46};
test_weights[17120:17127] = '{32'h429bf877, 32'hc2223d30, 32'h42aedcf9, 32'hc2182597, 32'hc1deb8f2, 32'hc2b8cdd4, 32'h42986cb1, 32'hc20f9e88};
test_bias[2140:2140] = '{32'h411544c5};
test_output[2140:2140] = '{32'h462417a5};
test_input[17128:17135] = '{32'hc2a570c4, 32'h41b19ff2, 32'hc28af523, 32'h42a6bcae, 32'h427fe53f, 32'hc24c85dd, 32'hc2a5d173, 32'hc15b8f2c};
test_weights[17128:17135] = '{32'hc2a9ebb9, 32'hc282367d, 32'hc2949803, 32'h428a524a, 32'hc1def7a2, 32'h42370144, 32'h42c61fd8, 32'h42aaf667};
test_bias[2141:2141] = '{32'h4159f011};
test_output[2141:2141] = '{32'h453c76a0};
test_input[17136:17143] = '{32'h42880c14, 32'h3ee9fb8d, 32'hc1aec4fc, 32'h42bc194c, 32'h42bcb759, 32'h427e3f79, 32'h4169e43b, 32'hc1b26bb4};
test_weights[17136:17143] = '{32'hc267b6ff, 32'h41b55738, 32'h4207f507, 32'hc28be072, 32'h4267e8a1, 32'h40f41bca, 32'hc21cfa40, 32'h42ba3ede};
test_bias[2142:2142] = '{32'hc2bb6ee2};
test_output[2142:2142] = '{32'hc5fb3929};
test_input[17144:17151] = '{32'hc18b9808, 32'hc28860a1, 32'h4278e3ec, 32'hc2b8e5c5, 32'h40fbc04d, 32'h42a5698d, 32'hc29d5f4e, 32'h427a8dec};
test_weights[17144:17151] = '{32'h414aab70, 32'hc225ef5b, 32'hc192a9a6, 32'h421c5dbd, 32'hc28b945e, 32'hc25953d3, 32'h42ade804, 32'hc2b20ed8};
test_bias[2143:2143] = '{32'h40359c72};
test_output[2143:2143] = '{32'hc6992ae0};
test_input[17152:17159] = '{32'h41bdd8de, 32'hc24d1d80, 32'hc221265f, 32'hc20001f7, 32'h42b98257, 32'hc0831828, 32'h40df5cbe, 32'h4201b7f3};
test_weights[17152:17159] = '{32'h4195a887, 32'h41f1bcb5, 32'h41920c56, 32'hc183e967, 32'hc2b62890, 32'h428cac6c, 32'hc19a6fe5, 32'hc2a04fd4};
test_bias[2144:2144] = '{32'h420758fa};
test_output[2144:2144] = '{32'hc647377a};
test_input[17160:17167] = '{32'hc2baf219, 32'h419288b3, 32'hc1804b0b, 32'h422fd453, 32'hc1265366, 32'h41ee0ffd, 32'h41d9974a, 32'hc1afd99c};
test_weights[17160:17167] = '{32'hc292321f, 32'h41dfb5c4, 32'hc222e753, 32'h41f4f6ab, 32'h41d58876, 32'hc1ccd99b, 32'hc261e7c6, 32'hc26629de};
test_bias[2145:2145] = '{32'h41c882af};
test_output[2145:2145] = '{32'h45fbd27b};
test_input[17168:17175] = '{32'h41621588, 32'hc176db2d, 32'hc2a4f1d9, 32'hc19b1db8, 32'h414981ac, 32'hc2b0ec16, 32'h41d7cb4b, 32'hc03ec4c1};
test_weights[17168:17175] = '{32'h408b0f0d, 32'hc24da2cb, 32'hc2b4ee6a, 32'hc19815ee, 32'hc19808e2, 32'h42aa4367, 32'h42680395, 32'h41294540};
test_bias[2146:2146] = '{32'hc227fae0};
test_output[2146:2146] = '{32'h45164fb1};
test_input[17176:17183] = '{32'h429256f9, 32'hc182e952, 32'h42481312, 32'hc2a9b1b0, 32'h41893d88, 32'hc23afbf1, 32'h428f1562, 32'h42bd6804};
test_weights[17176:17183] = '{32'hc284aa00, 32'hc209056a, 32'hc24e5980, 32'h40b61f6a, 32'h40e3f351, 32'h42b80ab9, 32'hc25bfb01, 32'h42bd943f};
test_bias[2147:2147] = '{32'h4243a0d9};
test_output[2147:2147] = '{32'hc5c96217};
test_input[17184:17191] = '{32'h40f422af, 32'h41831275, 32'h4264ab2a, 32'hbfd8faf2, 32'hc2beec77, 32'hc2bd841e, 32'h4124b694, 32'hc0ac76c1};
test_weights[17184:17191] = '{32'h40cb97eb, 32'h3f27cd53, 32'h42aaf706, 32'hc24ffa02, 32'h424e07b2, 32'h41e2be6c, 32'h41b05fdb, 32'hc045cef8};
test_bias[2148:2148] = '{32'hc224b4bf};
test_output[2148:2148] = '{32'hc513e13e};
test_input[17192:17199] = '{32'h41ce6ae5, 32'hc162536b, 32'h4299ede8, 32'hc22424f0, 32'hc1ac15b1, 32'h42b18d21, 32'h41f73f69, 32'h42c358bc};
test_weights[17192:17199] = '{32'hc11ceeab, 32'h422971b6, 32'h42031c63, 32'h42bb3d45, 32'h42882ddd, 32'hc1cf9837, 32'h42a9f324, 32'hc2a7ddc2};
test_bias[2149:2149] = '{32'h428822c0};
test_output[2149:2149] = '{32'hc632cd8b};
test_input[17200:17207] = '{32'hc2b30ba4, 32'hc20aac9a, 32'hc23be623, 32'h420e8037, 32'hc2c5efce, 32'h4204ad20, 32'hc22910f6, 32'h420f6e80};
test_weights[17200:17207] = '{32'hc068e0be, 32'hc223b527, 32'h425b8972, 32'h42a21e9b, 32'hc18d962b, 32'hc1141296, 32'hc2a0a2da, 32'hc2bf9a65};
test_bias[2150:2150] = '{32'h424d7d95};
test_output[2150:2150] = '{32'h455b5bb5};
test_input[17208:17215] = '{32'hc25ebb5a, 32'hc2a7c35e, 32'hc2c7beda, 32'h42af66c0, 32'hc2883371, 32'hc21a7c06, 32'h4221cfaf, 32'hc2c2068c};
test_weights[17208:17215] = '{32'hc05b7354, 32'hc1659de2, 32'hc20467e7, 32'h413316d7, 32'hc2ac82ad, 32'hc2bb67f4, 32'h41c7c984, 32'h4230d063};
test_bias[2151:2151] = '{32'hc25377b6};
test_output[2151:2151] = '{32'h46391139};
test_input[17216:17223] = '{32'hc1bb8eb7, 32'hc2b18ee7, 32'hc00ef407, 32'h42b135f3, 32'h42778fb9, 32'h42c4c577, 32'hc2942cbb, 32'hc1c1ef30};
test_weights[17216:17223] = '{32'hc20fd0ea, 32'h4214a075, 32'h42b53132, 32'h42024c0e, 32'hc2a7b0e8, 32'h42b612f1, 32'h42ba2ca8, 32'hc289ecdd};
test_bias[2152:2152] = '{32'hc20866b7};
test_output[2152:2152] = '{32'hc49dea0b};
test_input[17224:17231] = '{32'h41a9d53d, 32'h429f51d4, 32'hc1eb3361, 32'h42bca253, 32'hc26d99bd, 32'hc261b1c8, 32'h42b5d759, 32'hc2be4797};
test_weights[17224:17231] = '{32'hc28b84c2, 32'hc199ec37, 32'h42c35b78, 32'h420b3405, 32'hc0c2e432, 32'hc28c532d, 32'h4241ea3e, 32'h42825b9b};
test_bias[2153:2153] = '{32'h421cd548};
test_output[2153:2153] = '{32'hc212a489};
test_input[17232:17239] = '{32'hc204eeed, 32'hc2b483e2, 32'hc11012a5, 32'hc1d7b501, 32'hc2ab9e29, 32'hc217faea, 32'hc2438d27, 32'h4296e04a};
test_weights[17232:17239] = '{32'hc0c08edb, 32'h428f7669, 32'hc2076a62, 32'h423ea277, 32'h414151aa, 32'hc2806484, 32'hc0ad242e, 32'h41ef6cda};
test_bias[2154:2154] = '{32'h429b6dda};
test_output[2154:2154] = '{32'hc54b432d};
test_input[17240:17247] = '{32'h4130d7ed, 32'h42046b65, 32'hc2a7643f, 32'hc14823c0, 32'hc2bd862d, 32'h42886944, 32'hc18351f4, 32'h42c37901};
test_weights[17240:17247] = '{32'hc23fc4c3, 32'hc2a03a4e, 32'h42aa396d, 32'h42a02441, 32'h42c05cf6, 32'hc206fe10, 32'h422764c2, 32'h42653a24};
test_bias[2155:2155] = '{32'hc280626f};
test_output[2155:2155] = '{32'hc68ba309};
test_input[17248:17255] = '{32'hc16e2678, 32'hc2b0c75f, 32'h42172ddf, 32'h42b55c42, 32'h420925ab, 32'h429a6fce, 32'hc2584402, 32'hc20d3a4e};
test_weights[17248:17255] = '{32'h42379fe7, 32'hc2429be4, 32'hc18ac467, 32'h42249bb5, 32'h42403cfe, 32'h3fe340dd, 32'hc233f2bc, 32'hc2704fd6};
test_bias[2156:2156] = '{32'h42212ba2};
test_output[2156:2156] = '{32'h464c3f34};
test_input[17256:17263] = '{32'h42c63b36, 32'hc1eb7ff5, 32'hc224f1a1, 32'hc21a7b96, 32'h4215b249, 32'hc2898468, 32'h428fd9de, 32'hc24d69ee};
test_weights[17256:17263] = '{32'h4285ea6c, 32'hc22827c1, 32'h418c0c03, 32'h40fc9171, 32'h425c7e59, 32'h420ce82f, 32'hc20effea, 32'hc1b615a4};
test_bias[2157:2157] = '{32'hc2c59767};
test_output[2157:2157] = '{32'h459bd736};
test_input[17264:17271] = '{32'h42538594, 32'hc18fa66b, 32'hc2806d9f, 32'hc1e83205, 32'hc292cc84, 32'h422710e9, 32'h422b42ce, 32'h42442f8f};
test_weights[17264:17271] = '{32'h42a1693a, 32'hc291d158, 32'h429cb4b8, 32'h42197a78, 32'hc2171eba, 32'hc21c1681, 32'hc247f555, 32'hc2b7813f};
test_bias[2158:2158] = '{32'hc21a9993};
test_output[2158:2158] = '{32'hc5bebfdd};
test_input[17272:17279] = '{32'hc23856a8, 32'h42bfb41c, 32'hc1514e9c, 32'h4267e578, 32'h4293d569, 32'h42638064, 32'h423e4fd3, 32'hc28f58c2};
test_weights[17272:17279] = '{32'h42a0ed64, 32'hc27c792d, 32'hc292f65c, 32'h41a2d8c3, 32'h42c7bc31, 32'hc27ca43b, 32'h41288848, 32'hc2b2f271};
test_bias[2159:2159] = '{32'hc1b9a154};
test_output[2159:2159] = '{32'h453f7a9c};
test_input[17280:17287] = '{32'hc2948b56, 32'hc23c516e, 32'hc2330b30, 32'h3f28bff2, 32'h42b569cf, 32'h41a43397, 32'h42bc3f92, 32'h427ff1d8};
test_weights[17280:17287] = '{32'h4279fb23, 32'h427fab2c, 32'hc2bc341d, 32'hbf8d860c, 32'h426caba9, 32'h428eca3d, 32'h42b04ceb, 32'h42686601};
test_bias[2160:2160] = '{32'hc2551d57};
test_output[2160:2160] = '{32'h466fe8a7};
test_input[17288:17295] = '{32'h42221956, 32'hc2a296ff, 32'h426059a6, 32'h42424bf3, 32'h413213d1, 32'hc20399c9, 32'h42b1a037, 32'h4257efd7};
test_weights[17288:17295] = '{32'hc27b118c, 32'h41d8f9c0, 32'hc29730ba, 32'h42881391, 32'hc09819c2, 32'hc2c13af2, 32'hc1f20d67, 32'h420d4fe1};
test_bias[2161:2161] = '{32'hc2277ab4};
test_output[2161:2161] = '{32'hc5533ae1};
test_input[17296:17303] = '{32'hc2c4eda9, 32'hc2a52ebf, 32'hc1e8e6bc, 32'h425f6e39, 32'hc18b1533, 32'hc21e4f16, 32'h4294ed62, 32'hc29027e9};
test_weights[17296:17303] = '{32'hc24123b9, 32'h42373b8b, 32'hc0eee590, 32'hc0a16e83, 32'h42be4d4c, 32'hc24c47b1, 32'hc252f7e9, 32'h429415ce};
test_bias[2162:2162] = '{32'h4294b1c4};
test_output[2162:2162] = '{32'hc5f762cf};
test_input[17304:17311] = '{32'hc0fef394, 32'hc28390d3, 32'hc2b9ac6c, 32'h40e8b805, 32'h4294407b, 32'hc066d6dd, 32'h419f70c8, 32'h41a55765};
test_weights[17304:17311] = '{32'h4220c731, 32'h42b791a1, 32'hc29100f4, 32'h417226d1, 32'hc1286474, 32'h4267e1bb, 32'h429eefcf, 32'hc2b4f234};
test_bias[2163:2163] = '{32'hc1d3b528};
test_output[2163:2163] = '{32'hc44cbb94};
test_input[17312:17319] = '{32'hc2781790, 32'h420f43fd, 32'hc1fb151b, 32'h42b7494a, 32'hc2a5b755, 32'hc2b195ed, 32'h41697670, 32'h411671a5};
test_weights[17312:17319] = '{32'h42a2924c, 32'h41f6220e, 32'h4232e7f6, 32'hc24447bc, 32'hc254546b, 32'hc2b475a4, 32'hc1c61c86, 32'h4215ab39};
test_bias[2164:2164] = '{32'hc2afe894};
test_output[2164:2164] = '{32'h451a8448};
test_input[17320:17327] = '{32'h42b673a2, 32'hc2b9bdac, 32'h414513ea, 32'h419c0481, 32'h41a87cb1, 32'hc20f82d7, 32'h41856c4b, 32'h42829d62};
test_weights[17320:17327] = '{32'hc196312a, 32'hc27be561, 32'hc1829435, 32'hc282deca, 32'hc28fcc5f, 32'h425ee6c5, 32'hc2a91073, 32'hc29b7463};
test_bias[2165:2165] = '{32'h4199ec4e};
test_output[2165:2165] = '{32'hc5e4cdde};
test_input[17328:17335] = '{32'h420eaa6d, 32'h412ac2f3, 32'h4283497c, 32'hc2a5832a, 32'hc238cb61, 32'hbec98359, 32'h3fb920e6, 32'hc29fea9e};
test_weights[17328:17335] = '{32'h4293b234, 32'h40a3fd8a, 32'h4281dab9, 32'h40b1a54e, 32'h423ce55a, 32'h428c7561, 32'h4297faaf, 32'hc1574ad8};
test_bias[2166:2166] = '{32'h422d232d};
test_output[2166:2166] = '{32'h45ac37ef};
test_input[17336:17343] = '{32'hc111b009, 32'hc29fa886, 32'h42c646a8, 32'h41e20493, 32'h42a41ae4, 32'hc1efe791, 32'h426b8dbb, 32'hc28991f9};
test_weights[17336:17343] = '{32'hc28b863b, 32'h41cea28d, 32'h42a7ebd9, 32'hc2bc1151, 32'hc1b597b3, 32'hc28150b3, 32'h42b27ce7, 32'h42ab5cbf};
test_bias[2167:2167] = '{32'hc22d89e4};
test_output[2167:2167] = '{32'h4563335c};
test_input[17344:17351] = '{32'hc0040153, 32'hc201427b, 32'h423f979a, 32'hc231e123, 32'hc2b66672, 32'h42aa9ba9, 32'h42b8bc10, 32'h423f57d2};
test_weights[17344:17351] = '{32'h428a6327, 32'h41cd91da, 32'hc1b305f9, 32'hc2b4a710, 32'h42494a21, 32'h3e3dc9ea, 32'hc091a920, 32'h429ce996};
test_bias[2168:2168] = '{32'hc20293ab};
test_output[2168:2168] = '{32'h442e8b4f};
test_input[17352:17359] = '{32'h4205e423, 32'h421da610, 32'h423ef12e, 32'hc013e72c, 32'h4215dc9d, 32'h420cfda0, 32'h422689aa, 32'hc0f91ab8};
test_weights[17352:17359] = '{32'hc256a517, 32'h42756ae2, 32'h40dc2334, 32'h4245a996, 32'h4219e469, 32'hc1c327fe, 32'hc2573dfb, 32'h3fff479d};
test_bias[2169:2169] = '{32'h429f566f};
test_output[2169:2169] = '{32'hc43da3ec};
test_input[17360:17367] = '{32'h42925f94, 32'h42666322, 32'h428e800d, 32'h42076d29, 32'hc2574697, 32'hc1d8557e, 32'hc2073f8e, 32'hc1a10da1};
test_weights[17360:17367] = '{32'hc2b4c3d6, 32'hc0e51211, 32'h42610b41, 32'hc1e446d5, 32'h3eb8d54b, 32'h4165c36b, 32'hc1e04797, 32'hc222abca};
test_bias[2170:2170] = '{32'hc1f47360};
test_output[2170:2170] = '{32'hc5260430};
test_input[17368:17375] = '{32'h42bb6a91, 32'hc28b823d, 32'h41f335f6, 32'h42690c27, 32'h42003a24, 32'h42acf3cb, 32'hc21e1339, 32'hc28902e3};
test_weights[17368:17375] = '{32'hc28ec8dd, 32'hc0b6ba6a, 32'h41812af8, 32'h42544413, 32'hc29a6f9f, 32'hc224e150, 32'h42186c07, 32'hc265a2a1};
test_bias[2171:2171] = '{32'h4217fdff};
test_output[2171:2171] = '{32'hc5c460a5};
test_input[17376:17383] = '{32'hbf1d0f27, 32'hc298f1d7, 32'hc2b52ad9, 32'hc2adcd8b, 32'hc19f2c3f, 32'h41e59ef7, 32'h42ae3692, 32'hc285edf9};
test_weights[17376:17383] = '{32'h41edcdac, 32'h42152687, 32'h4258ee18, 32'hc29722a8, 32'h4233a9e5, 32'hc0d5f807, 32'hc2aec254, 32'h41d3e659};
test_bias[2172:2172] = '{32'h42147004};
test_output[2172:2172] = '{32'hc6360395};
test_input[17384:17391] = '{32'h42684b6e, 32'h422bfb44, 32'h409ec240, 32'hc10a1ed1, 32'hc105eaa7, 32'h42ba6961, 32'hc29eaea5, 32'h425b9414};
test_weights[17384:17391] = '{32'hc2c5cca3, 32'h428f525d, 32'h42ade009, 32'hc20cf431, 32'h428bc16a, 32'h41664bca, 32'hc1d39ec5, 32'h426b0329};
test_bias[2173:2173] = '{32'hc2bc9965};
test_output[2173:2173] = '{32'h457db875};
test_input[17392:17399] = '{32'h424a936c, 32'hc2b25e62, 32'hc265c6ec, 32'h4242d87d, 32'hc2728315, 32'h4047e3fb, 32'hc2ac3d2c, 32'hbf73100e};
test_weights[17392:17399] = '{32'hc221f714, 32'hc2468bd2, 32'h412ef726, 32'h42611be3, 32'hc263bc13, 32'h42a39111, 32'hc18b59b2, 32'hc295caeb};
test_bias[2174:2174] = '{32'hc2323296};
test_output[2174:2174] = '{32'h4617eccf};
test_input[17400:17407] = '{32'hc25a108e, 32'h425c365c, 32'hc2c428c1, 32'h42513844, 32'h42574dff, 32'h42831f49, 32'h42acd47f, 32'hc211de18};
test_weights[17400:17407] = '{32'h425f5508, 32'hc0b990e6, 32'hc27aa27b, 32'h42b2d9ec, 32'h413e8c73, 32'h41920ed4, 32'h42818ec7, 32'hc2ab7410};
test_bias[2175:2175] = '{32'h40cfad1a};
test_output[2175:2175] = '{32'h468cd8da};
test_input[17408:17415] = '{32'h42b18888, 32'hc213b4cd, 32'hc28e87db, 32'h42506ebd, 32'hc1d2b11e, 32'h4289d427, 32'h42087bbd, 32'h4288ccc1};
test_weights[17408:17415] = '{32'h42ae2527, 32'h40ec6bff, 32'h425f67b5, 32'hc280afb9, 32'hc17a68c7, 32'hc298cd1d, 32'h42973601, 32'hc2944847};
test_bias[2176:2176] = '{32'h419f4a7c};
test_output[2176:2176] = '{32'hc5e10a3a};
test_input[17416:17423] = '{32'h423a2f66, 32'h4189c3fd, 32'h425b0998, 32'h42b6bfe9, 32'hc2ba184b, 32'h425270bf, 32'hc24b0dc9, 32'hc2696cfc};
test_weights[17416:17423] = '{32'h428acf30, 32'h41e467af, 32'h4232a7ac, 32'hc29b826a, 32'hc2b737d9, 32'h41595c4d, 32'hc268a5c9, 32'hc1f7dc72};
test_bias[2177:2177] = '{32'hc28a9143};
test_output[2177:2177] = '{32'h464b0451};
test_input[17424:17431] = '{32'h411801ed, 32'h42600185, 32'hc299494f, 32'h41af3a1b, 32'h42c7b901, 32'hc24d69c6, 32'h42525774, 32'h42b8a0b7};
test_weights[17424:17431] = '{32'hc24f14bf, 32'hc131536b, 32'h4185e438, 32'h42806d71, 32'h417e15cc, 32'hc2af4497, 32'hc147869f, 32'hc2bc66ed};
test_bias[2178:2178] = '{32'h429113a6};
test_output[2178:2178] = '{32'hc582af2c};
test_input[17432:17439] = '{32'h425eb408, 32'hc23d0062, 32'h420e0ca3, 32'hc2580dc1, 32'hc22f3476, 32'hc2732e3c, 32'h42394833, 32'hc1cde924};
test_weights[17432:17439] = '{32'hc1030b89, 32'h424bae4a, 32'h42b53cbb, 32'h42af1de2, 32'hc1b2c760, 32'h42be855f, 32'h428a24e2, 32'hc2b290dd};
test_bias[2179:2179] = '{32'h42924456};
test_output[2179:2179] = '{32'hc561f290};
test_input[17440:17447] = '{32'hc1b71977, 32'h422a79bb, 32'hc29f81fe, 32'hc0bc532c, 32'hc2101dd9, 32'h41b4d2c5, 32'hc23262da, 32'hc27f00b6};
test_weights[17440:17447] = '{32'hc2ad08bf, 32'hc26052de, 32'h42b17c19, 32'hc0d3dc57, 32'h428eb5df, 32'h41ec86f1, 32'h41beee37, 32'h4191ef03};
test_bias[2180:2180] = '{32'hc26b319a};
test_output[2180:2180] = '{32'hc635d4d2};
test_input[17448:17455] = '{32'h420ff645, 32'hc29b8d7a, 32'hc238351a, 32'h425695b0, 32'h428d151d, 32'hc2bbeba9, 32'h421bf866, 32'h42b3f915};
test_weights[17448:17455] = '{32'hc1282341, 32'h42a08909, 32'h42a8baf2, 32'h429906a4, 32'hc24aff1a, 32'h42a3bff3, 32'hc264a05e, 32'hc20802cc};
test_bias[2181:2181] = '{32'hc21fc8e7};
test_output[2181:2181] = '{32'hc6b3b5f8};
test_input[17456:17463] = '{32'h417a6093, 32'h422f2319, 32'hc243b3fa, 32'hc1e8377c, 32'h4266098b, 32'h41f0adb6, 32'hc2264e4a, 32'hc1f8e401};
test_weights[17456:17463] = '{32'h429cbd7c, 32'h42ad5c19, 32'hc2c3fbec, 32'hc1c0263f, 32'hc245d0c7, 32'hc221c4b8, 32'h4290ec5f, 32'h41857b7c};
test_bias[2182:2182] = '{32'h42762c40};
test_output[2182:2182] = '{32'h453a61cd};
test_input[17464:17471] = '{32'h42a6faba, 32'hc2326cdb, 32'hc208320c, 32'hc2801623, 32'hc2327710, 32'h41c4d874, 32'hc13826ca, 32'hc18fb338};
test_weights[17464:17471] = '{32'h420ae873, 32'h42160332, 32'hc1f7bd9a, 32'h42985169, 32'hc2b89d49, 32'hc20dde65, 32'h42a8d453, 32'h42a3e878};
test_bias[2183:2183] = '{32'h42ba85b4};
test_output[2183:2183] = '{32'hc4d4a922};
test_input[17472:17479] = '{32'hc293d6e6, 32'h428c9e14, 32'hc2a9359e, 32'hc0af5b45, 32'hc20fd337, 32'h424d496b, 32'h42a9cfaa, 32'hc0ca3f82};
test_weights[17472:17479] = '{32'h40e862f9, 32'hc294b21d, 32'hc17a95a6, 32'hc167db2b, 32'hc1eb0e51, 32'h426772d6, 32'hc1efe120, 32'h4262698b};
test_bias[2184:2184] = '{32'hc18fc1d6};
test_output[2184:2184] = '{32'hc54b738b};
test_input[17480:17487] = '{32'h422e6241, 32'h41334ba5, 32'hc2575b5b, 32'h4189069f, 32'hc226435c, 32'hc25f5e32, 32'h4067953b, 32'hc1c41dfa};
test_weights[17480:17487] = '{32'h4258a7ad, 32'hc28f9e7e, 32'h42a462ae, 32'hc268630c, 32'h41a36535, 32'hc099cbfb, 32'h428ef261, 32'h428fa638};
test_bias[2185:2185] = '{32'hc29441b7};
test_output[2185:2185] = '{32'hc5bc23f0};
test_input[17488:17495] = '{32'hc28e5587, 32'h42817433, 32'hc2c5ca16, 32'hc2a7669f, 32'h420e5658, 32'hc297c9f9, 32'h41365bac, 32'h425bf41a};
test_weights[17488:17495] = '{32'h42c054d4, 32'h41a8e3fe, 32'h416ca259, 32'hc1ec0f23, 32'hc20fabf5, 32'h42b57e1d, 32'hc1ff8194, 32'hc28dc905};
test_bias[2186:2186] = '{32'h40c56b33};
test_output[2186:2186] = '{32'hc683f720};
test_input[17496:17503] = '{32'hc2391f30, 32'hc2a9bfc0, 32'h4298da2f, 32'h418ad60d, 32'h4283daf6, 32'hc299e603, 32'h412fed60, 32'h42129b22};
test_weights[17496:17503] = '{32'h42abc38e, 32'hbe59d4f5, 32'hc238fefe, 32'hc23f4451, 32'hc2923f22, 32'hc2855f99, 32'hc11ed6f4, 32'h4293c44e};
test_bias[2187:2187] = '{32'h4291d83b};
test_output[2187:2187] = '{32'hc5a6d5c9};
test_input[17504:17511] = '{32'hc2960583, 32'hc1a75bc0, 32'hc13dff0b, 32'hc25aff83, 32'hc0d4231c, 32'h41ffade5, 32'h42bb653f, 32'hc290ed96};
test_weights[17504:17511] = '{32'h42bbea93, 32'hc02b05a2, 32'hc20ea035, 32'hc26af0fb, 32'h41e29039, 32'h424a82bf, 32'h42bc6a03, 32'h405ba968};
test_bias[2188:2188] = '{32'hc1d7e13b};
test_output[2188:2188] = '{32'h45cf2634};
test_input[17512:17519] = '{32'hc25cd7eb, 32'h42c29854, 32'hc2bb4a03, 32'h429226ed, 32'hc18aba12, 32'h424023f3, 32'hc2c7cf80, 32'hc29e14de};
test_weights[17512:17519] = '{32'hc263dd08, 32'hc2bdf1f4, 32'hc29bd23a, 32'hc26af899, 32'hc0daba33, 32'h406d8578, 32'h4297206e, 32'h429cf81b};
test_bias[2189:2189] = '{32'hc2b7d3df};
test_output[2189:2189] = '{32'hc6820009};
test_input[17520:17527] = '{32'h42679d2c, 32'hc115bfb1, 32'hc299d9bf, 32'hc095c6e2, 32'h424cbc97, 32'h42ace6b3, 32'h428e626a, 32'hc15f6373};
test_weights[17520:17527] = '{32'hc2385818, 32'hc289785a, 32'hc26e3ce8, 32'hc29355f9, 32'h426244f9, 32'hc1a1474b, 32'hc2a12300, 32'hc2414438};
test_bias[2190:2190] = '{32'h427a4ca8};
test_output[2190:2190] = '{32'hc46c3cb6};
test_input[17528:17535] = '{32'h429ed6d3, 32'h425d6346, 32'h42864709, 32'h410f377f, 32'hc23581e9, 32'hc269f82a, 32'hc28bdd41, 32'h41b3e206};
test_weights[17528:17535] = '{32'hc1ca8fe5, 32'h42c79401, 32'hc2c01443, 32'h428cd2f3, 32'hc2441ab0, 32'h42895c2e, 32'hc2c2c195, 32'h4247a696};
test_bias[2191:2191] = '{32'hc25c7687};
test_output[2191:2191] = '{32'h456c2d23};
test_input[17536:17543] = '{32'hc2633e94, 32'hbfeed9ad, 32'h42792469, 32'h42b80372, 32'h42b4cc39, 32'h41b3df42, 32'hc25dd996, 32'hbffed4e3};
test_weights[17536:17543] = '{32'hc10719bb, 32'h411717a4, 32'h41fc5fef, 32'h41d434d8, 32'h42749526, 32'hc1cdd233, 32'hc25327c7, 32'hc0779196};
test_bias[2192:2192] = '{32'h4223adc1};
test_output[2192:2192] = '{32'h4647e403};
test_input[17544:17551] = '{32'h42c0f7c6, 32'hc2c43a5d, 32'h424f3318, 32'h41558939, 32'hc0be52bf, 32'hc1fd7d39, 32'hc18b1e1d, 32'hc284a08a};
test_weights[17544:17551] = '{32'hc29adccd, 32'hc259f44c, 32'hc2a614d0, 32'h42754ae2, 32'h42ba6cba, 32'h42ac858c, 32'hc2930e33, 32'hc213c3a3};
test_bias[2193:2193] = '{32'h41b5b2c9};
test_output[2193:2193] = '{32'hc5a0c3ef};
test_input[17552:17559] = '{32'h425c5beb, 32'hc2a04293, 32'hc2bf7eaf, 32'h4125eaca, 32'h429001e4, 32'h429a9b6f, 32'h428377cb, 32'hc2b6c098};
test_weights[17552:17559] = '{32'h42a127f9, 32'h42a6d7b7, 32'hc2197c76, 32'h4225d573, 32'hc2b405ab, 32'hc25d5b8a, 32'hc1e45c8e, 32'h42604650};
test_bias[2194:2194] = '{32'hc2891bc8};
test_output[2194:2194] = '{32'hc67983e9};
test_input[17560:17567] = '{32'h426a91ff, 32'hc25626c1, 32'hc2b47dbc, 32'hc0c28830, 32'h4227c35d, 32'hc28ffa70, 32'h428d95ab, 32'h41b7df8a};
test_weights[17560:17567] = '{32'hc20400a3, 32'hc2b16223, 32'hc28b5f94, 32'hc1b1efaa, 32'hc1c91140, 32'hc16934dc, 32'h4232eedf, 32'h421d2226};
test_bias[2195:2195] = '{32'h428436b4};
test_output[2195:2195] = '{32'h4650e0b3};
test_input[17568:17575] = '{32'h42c0a95e, 32'hc24472c5, 32'hc202263f, 32'h422ae5d9, 32'h4086688c, 32'h42c207cc, 32'h41e278d9, 32'h4278d9e5};
test_weights[17568:17575] = '{32'hc2840e45, 32'h41df1653, 32'h42855aef, 32'h42b7f216, 32'h42ab6cca, 32'hc23b4294, 32'h42932d9b, 32'hc26adf14};
test_bias[2196:2196] = '{32'h4261b16b};
test_output[2196:2196] = '{32'hc63644b3};
test_input[17576:17583] = '{32'h42639fb3, 32'hc249372c, 32'h405e4094, 32'hc2495efd, 32'h42289145, 32'h41d6144c, 32'hc1ecce03, 32'hc1d3f10f};
test_weights[17576:17583] = '{32'h4242c5e6, 32'h41bfcf07, 32'hc2a9da76, 32'h40962cb1, 32'hc2bd4592, 32'hc20a7b65, 32'hc1f56f63, 32'h419f810e};
test_bias[2197:2197] = '{32'h42976e62};
test_output[2197:2197] = '{32'hc556146c};
test_input[17584:17591] = '{32'hc2c2cd20, 32'h42ba1b7e, 32'hc29b33c2, 32'h42890bee, 32'h4213a1c8, 32'hc1cc3dd2, 32'h41c52664, 32'hc2aa6a8e};
test_weights[17584:17591] = '{32'h3fa82015, 32'h427e204e, 32'h41d540b6, 32'hc2545a9e, 32'h421f0212, 32'hc23817fd, 32'h42a04de3, 32'hc29de2c2};
test_bias[2198:2198] = '{32'hc2895bf2};
test_output[2198:2198] = '{32'h46316351};
test_input[17592:17599] = '{32'h41ee6bb3, 32'h4185dc30, 32'hc22ffe87, 32'h427bf0a9, 32'hc2b47a88, 32'hc1675420, 32'h41a82a2b, 32'hc2964900};
test_weights[17592:17599] = '{32'h421bb756, 32'hc1985ada, 32'hc2854d1c, 32'h42b7fb05, 32'h421ceab7, 32'h4247df7a, 32'hc285de1e, 32'h42756cbf};
test_bias[2199:2199] = '{32'hc280e5c0};
test_output[2199:2199] = '{32'hc44212d6};
test_input[17600:17607] = '{32'hc0da77ec, 32'hc280fd9f, 32'h4296ba52, 32'hc1ca8e23, 32'hc0c68089, 32'hc1bb7ce9, 32'hc2a2bfa9, 32'h40c81feb};
test_weights[17600:17607] = '{32'hc22ccb4d, 32'hc26242bf, 32'hc2445c63, 32'h427cd660, 32'hc28aad77, 32'h4136dcd6, 32'hc2960ebf, 32'h424d797e};
test_bias[2200:2200] = '{32'h42affcf8};
test_output[2200:2200] = '{32'h45a64001};
test_input[17608:17615] = '{32'hc2018aac, 32'hc1aef0e5, 32'h429b208c, 32'h429f81d6, 32'hc26acaa8, 32'h40a3376e, 32'hc2b787e4, 32'hc2c644bf};
test_weights[17608:17615] = '{32'hc2189454, 32'h42a953f5, 32'hc081a5d2, 32'hc1eb388a, 32'hc1c1a9e8, 32'hc27afaf5, 32'hc2789561, 32'h429209dc};
test_bias[2201:2201] = '{32'hc2bc287a};
test_output[2201:2201] = '{32'hc56dc4c2};
test_input[17616:17623] = '{32'hc26252ec, 32'hc2205215, 32'h4292e7a9, 32'h4211d08d, 32'hc260edaf, 32'h4270b053, 32'hc22c3e46, 32'hc1d143a9};
test_weights[17616:17623] = '{32'hc2334cf1, 32'hc22f820d, 32'h42049a9b, 32'h42c33156, 32'h41af2caf, 32'h423af850, 32'h411ddde4, 32'h42799594};
test_bias[2202:2202] = '{32'hc2784734};
test_output[2202:2202] = '{32'h4618573f};
test_input[17624:17631] = '{32'hc1eff880, 32'h41448ef1, 32'hc20e6a80, 32'hc28d68ec, 32'hc2330220, 32'hc2b51000, 32'hc24af486, 32'h41d4d6fb};
test_weights[17624:17631] = '{32'h419f55dc, 32'hc278c7aa, 32'h41139631, 32'hc1b78ce6, 32'h42649759, 32'hc2459fba, 32'h42900aa8, 32'hc28ac939};
test_bias[2203:2203] = '{32'hc2be96c6};
test_output[2203:2203] = '{32'hc56a41ca};
test_input[17632:17639] = '{32'hc2c6d699, 32'hc20b5dc1, 32'hc2a78012, 32'hc12d95f2, 32'h4280094b, 32'hc23299a8, 32'hc28c724f, 32'h4204ad78};
test_weights[17632:17639] = '{32'hc2733cfe, 32'hc2502826, 32'h428b8e29, 32'hc26aef1c, 32'hc1f5b474, 32'h428323a1, 32'hc287327a, 32'hc2815007};
test_bias[2204:2204] = '{32'h41480eec};
test_output[2204:2204] = '{32'h43ba8a89};
test_input[17640:17647] = '{32'hc234d179, 32'hc20b4bde, 32'hc2a975c0, 32'hc1ec3ce0, 32'hc23af016, 32'h41976a46, 32'h3ec9c9be, 32'h424bf95d};
test_weights[17640:17647] = '{32'h42b52d16, 32'h42a32714, 32'h4264a597, 32'h42aee764, 32'h423ca6cb, 32'h42afe212, 32'h428c26c4, 32'hc2539248};
test_bias[2205:2205] = '{32'h42c1f10d};
test_output[2205:2205] = '{32'hc68883aa};
test_input[17648:17655] = '{32'hc28a7754, 32'hc2a4a1a0, 32'hc2c04749, 32'h4281165e, 32'h4187b1ff, 32'hc29fbe84, 32'hc2373943, 32'hc187d6e4};
test_weights[17648:17655] = '{32'h428d061c, 32'hc23e5c0b, 32'hc2818666, 32'h41a2bd76, 32'h4239c44d, 32'h427cce88, 32'h42719f2b, 32'h41d9663c};
test_bias[2206:2206] = '{32'hc27bc809};
test_output[2206:2206] = '{32'hc47431d6};
test_input[17656:17663] = '{32'h42a263a7, 32'hc2acda66, 32'h42968e16, 32'hc2b0256f, 32'hc186ec4d, 32'h41645b53, 32'hc24f8c3a, 32'hc2b7bd16};
test_weights[17656:17663] = '{32'h42423140, 32'h426883d2, 32'hc292e29a, 32'hc199b15a, 32'hc2a98ae3, 32'hc2aebe24, 32'h42ba246d, 32'h41dec061};
test_bias[2207:2207] = '{32'hc2896562};
test_output[2207:2207] = '{32'hc63e7ef6};
test_input[17664:17671] = '{32'hc2845c27, 32'h42b29c9d, 32'h41e13079, 32'hc22a1fab, 32'hc1f1b8a3, 32'hc1101d1a, 32'h3d575223, 32'h420c0fc2};
test_weights[17664:17671] = '{32'h428647a4, 32'hc2bb36b2, 32'hc1ae6363, 32'h3fa86707, 32'hc29af484, 32'hc2ad4851, 32'hc11a57c1, 32'h42c38492};
test_bias[2208:2208] = '{32'hc20f6125};
test_output[2208:2208] = '{32'hc5d9a355};
test_input[17672:17679] = '{32'hc28843b4, 32'hbe940d3b, 32'hc1fa226b, 32'h42b54b3b, 32'h408ff6c2, 32'hc2c6adba, 32'h42904760, 32'h4219c54c};
test_weights[17672:17679] = '{32'h422c13d3, 32'hc1af2e60, 32'hc0db17f2, 32'hc293ac02, 32'h428c39f6, 32'h3dc6bec8, 32'h4266a63b, 32'h422033b3};
test_bias[2209:2209] = '{32'h4298a25f};
test_output[2209:2209] = '{32'hc54fa1f0};
test_input[17680:17687] = '{32'hc2bceed9, 32'hc0f39fbd, 32'h406c9d09, 32'hc28381b2, 32'hc2a6e897, 32'h4290d714, 32'hc21804b2, 32'h421cae2b};
test_weights[17680:17687] = '{32'hc1e6f4d5, 32'hc1f521e4, 32'h4188b5bd, 32'h42acd00f, 32'hc292cbb7, 32'hc222b639, 32'hc1066238, 32'hc14f3bce};
test_bias[2210:2210] = '{32'h41917c5d};
test_output[2210:2210] = '{32'h43afd6cd};
test_input[17688:17695] = '{32'hc2b29296, 32'h42999786, 32'hc18f57df, 32'hc2b1f45e, 32'hc291b80c, 32'hc2107652, 32'h42948e45, 32'h42bdfb69};
test_weights[17688:17695] = '{32'h3fbdbff6, 32'hc1d86e52, 32'h4124d92a, 32'h41e4a433, 32'hc25f057d, 32'hc086a428, 32'hc2850707, 32'hc2526a62};
test_bias[2211:2211] = '{32'h404c777f};
test_output[2211:2211] = '{32'hc6268613};
test_input[17696:17703] = '{32'h411dc0c5, 32'hc2958f34, 32'hc217266a, 32'hc28c97f9, 32'hc28e6ab0, 32'h42c64e8c, 32'h42400b2c, 32'h42ba9733};
test_weights[17696:17703] = '{32'hc1a3fd91, 32'hc224b33e, 32'h41c57416, 32'h42711551, 32'hc250d72c, 32'hc2098263, 32'h420becd5, 32'h41dcc638};
test_bias[2212:2212] = '{32'h3ef59db2};
test_output[2212:2212] = '{32'h450df395};
test_input[17704:17711] = '{32'hc19a8420, 32'hc1d6031b, 32'h425f6433, 32'hc2853b4b, 32'h41c10a6b, 32'h42a1c742, 32'hc2ad4a67, 32'hc0ffd1f8};
test_weights[17704:17711] = '{32'hc109081f, 32'h426da792, 32'h42a3e440, 32'h428ac4ca, 32'hc20f179e, 32'hc1e6f2be, 32'hc2a4e287, 32'h429d3962};
test_bias[2213:2213] = '{32'h423015f0};
test_output[2213:2213] = '{32'h44ec5c02};
test_input[17712:17719] = '{32'h428688cc, 32'hc245f7cd, 32'h428ce6f2, 32'hc12a86c7, 32'h42a79a35, 32'hc118599b, 32'hc0b33d2b, 32'h42a52421};
test_weights[17712:17719] = '{32'h4070e81e, 32'h420d0db0, 32'h429a21be, 32'h3ed7a5c0, 32'h416a377e, 32'hc1d768fc, 32'hc2c06e27, 32'h42c4e392};
test_bias[2214:2214] = '{32'h42c06a6e};
test_output[2214:2214] = '{32'h465d8ecb};
test_input[17720:17727] = '{32'hc2c5d994, 32'hc2b6c053, 32'hc14d2054, 32'hc2b7d5a1, 32'h42bca74e, 32'hc26d2b79, 32'hc241ddc9, 32'h42719d05};
test_weights[17720:17727] = '{32'hc2a84ce6, 32'h4180997c, 32'hc2441880, 32'h429c67f4, 32'hc05389cb, 32'hc2a9e13f, 32'hc28a9a5b, 32'h422c28ce};
test_bias[2215:2215] = '{32'h42b675c5};
test_output[2215:2215] = '{32'h462cf935};
test_input[17728:17735] = '{32'h42199fc9, 32'hc29f4ab4, 32'h42c41e67, 32'h42030505, 32'h421c1dab, 32'hc2ae3c8b, 32'hc244208f, 32'h42a9fb8a};
test_weights[17728:17735] = '{32'h4104b770, 32'h4158f105, 32'h41151cd3, 32'h419fbffb, 32'h42936b94, 32'hc2843d12, 32'h4257e351, 32'h42b79985};
test_bias[2216:2216] = '{32'hc0e5001c};
test_output[2216:2216] = '{32'h46640146};
test_input[17736:17743] = '{32'hc28ee9ba, 32'hc11f55a0, 32'h42bcd847, 32'hc23069f5, 32'hc27abcd6, 32'h42c58eff, 32'hc03f45a9, 32'h42906d0a};
test_weights[17736:17743] = '{32'h422a0a80, 32'hc1887b64, 32'h41e5f1c9, 32'h42ac375a, 32'hc2b8256d, 32'hc24a742b, 32'h42a5d1d7, 32'h40146693};
test_bias[2217:2217] = '{32'h42c34cdb};
test_output[2217:2217] = '{32'hc545a1f6};
test_input[17744:17751] = '{32'h408af907, 32'h41e2d8f4, 32'h41b30d17, 32'hc051c194, 32'hc2ab5536, 32'h42bb09cd, 32'h418973b6, 32'h40d20943};
test_weights[17744:17751] = '{32'hc2893d96, 32'hc247def1, 32'hc2c4465a, 32'hc2599435, 32'h429e5cea, 32'hc28e23a1, 32'hc046e8e7, 32'h426ebba8};
test_bias[2218:2218] = '{32'h42690bed};
test_output[2218:2218] = '{32'hc682fc0e};
test_input[17752:17759] = '{32'h42b521ef, 32'hc27f2f85, 32'h42a0614e, 32'hc201762a, 32'h422a999a, 32'h3f25eab0, 32'hc20c3101, 32'hc2a0098c};
test_weights[17752:17759] = '{32'hc284fbad, 32'hc2a8f2fd, 32'hc2839474, 32'h429af7ad, 32'h42ad7b34, 32'hc2c428d9, 32'h42a9184b, 32'hc2a80df4};
test_bias[2219:2219] = '{32'hc06320f7};
test_output[2219:2219] = '{32'hc47fd2e7};
test_input[17760:17767] = '{32'hc1b5df24, 32'hc14df9ad, 32'h41ab5965, 32'h428c2220, 32'hc248041b, 32'hc28893c6, 32'hc1bf2411, 32'h42250a0c};
test_weights[17760:17767] = '{32'hc2ae5d63, 32'h42825d52, 32'hc2378167, 32'hc2c458db, 32'h41288acc, 32'h401c3503, 32'hc207c7d6, 32'h42a7dcf8};
test_bias[2220:2220] = '{32'hc29bfa08};
test_output[2220:2220] = '{32'hc548fc83};
test_input[17768:17775] = '{32'h4144e282, 32'hc21f2230, 32'hc2a309dc, 32'hc1273876, 32'hc2bf05c6, 32'hc25156d6, 32'h41baddf3, 32'hc2a62cc1};
test_weights[17768:17775] = '{32'hc2ae8fc7, 32'h42bc4d0b, 32'hc2373bf0, 32'h427df8af, 32'hc2b30c02, 32'hc201b074, 32'h41fa2592, 32'h424edf1e};
test_bias[2221:2221] = '{32'hc1d97bc7};
test_output[2221:2221] = '{32'h459943a7};
test_input[17776:17783] = '{32'hc209660f, 32'h42417a09, 32'hc2c5f179, 32'hc284026d, 32'hc28b99fc, 32'hc1cb69e6, 32'hc2a51cbb, 32'h42026348};
test_weights[17776:17783] = '{32'h41528d08, 32'hc2697d16, 32'hc14fc710, 32'hc1cda9fa, 32'hc214ba6a, 32'hc2b8f576, 32'hc274ae6b, 32'h409d052c};
test_bias[2222:2222] = '{32'hc2c042a3};
test_output[2222:2222] = '{32'h46189d06};
test_input[17784:17791] = '{32'h429388b5, 32'hc274c7a8, 32'hc253e9cc, 32'h4118383d, 32'h42262316, 32'h4275a783, 32'hc1efb492, 32'h42bc54e7};
test_weights[17784:17791] = '{32'hc20a001e, 32'hc2924fc4, 32'hc217b842, 32'h42843e2e, 32'hc2818c3b, 32'hc296e5b3, 32'h42688213, 32'h42912aac};
test_bias[2223:2223] = '{32'h42272cbf};
test_output[2223:2223] = '{32'h4514d68e};
test_input[17792:17799] = '{32'hc2828f90, 32'hc2b5c76e, 32'h417d3eb7, 32'h428451c5, 32'hc25b6e2c, 32'h42992c1c, 32'hc10d1fb1, 32'h42540eaf};
test_weights[17792:17799] = '{32'h4280b066, 32'hc1a09c3f, 32'h42a64118, 32'h428b3ea1, 32'h42b6cee5, 32'h42baa159, 32'h42a3e11f, 32'hc2704123};
test_bias[2224:2224] = '{32'h41e407f2};
test_output[2224:2224] = '{32'h44e105e1};
test_input[17800:17807] = '{32'h41901f89, 32'hc227c253, 32'h42418164, 32'h41211bb1, 32'hc18a3632, 32'hc2408682, 32'hc124b394, 32'hc1ce5b65};
test_weights[17800:17807] = '{32'hc2aad04e, 32'h4068353a, 32'h429f7d3d, 32'h42885c30, 32'h40eb8995, 32'hc26a5d6e, 32'h4229ed5f, 32'h42982986};
test_bias[2225:2225] = '{32'hc2a1e3b4};
test_output[2225:2225] = '{32'h453f9a70};
test_input[17808:17815] = '{32'h41b0f2b0, 32'hc285baf4, 32'hc29331d1, 32'h429e52d2, 32'hc0db625b, 32'hc2ad615e, 32'h42c673c5, 32'h42128140};
test_weights[17808:17815] = '{32'h42192280, 32'hc1c0611d, 32'hc19c5f42, 32'hbfc8dda9, 32'hc1fcbcce, 32'hc2a12ca6, 32'h42232fbd, 32'h41dc1c0d};
test_bias[2226:2226] = '{32'h42aaafd3};
test_output[2226:2226] = '{32'h467bc3ad};
test_input[17816:17823] = '{32'h42bdeb54, 32'hc0849485, 32'h42a5417b, 32'hc297f6d5, 32'hbe4bacf9, 32'hc26def90, 32'hc2bf7fd2, 32'hc1459f59};
test_weights[17816:17823] = '{32'hc249cf0f, 32'h4247c657, 32'hc2264820, 32'hc2a14316, 32'hc15675ee, 32'h42052279, 32'hc295a7fa, 32'hc2a2e81d};
test_bias[2227:2227] = '{32'hc1ae3a94};
test_output[2227:2227] = '{32'h45719a93};
test_input[17824:17831] = '{32'h41cac9a3, 32'hc1736c19, 32'hc2810f53, 32'h42c0f6ce, 32'h4186f548, 32'hc20088d7, 32'h427c229e, 32'h41147600};
test_weights[17824:17831] = '{32'hc2a751e6, 32'h414ddda5, 32'hc13c2309, 32'h424d7eb0, 32'h41f98a27, 32'hc26c9774, 32'h427a43ab, 32'h42752de5};
test_bias[2228:2228] = '{32'hc2c4511a};
test_output[2228:2228] = '{32'h462000e9};
test_input[17832:17839] = '{32'h424abcf2, 32'h4271bbfc, 32'hc2912e77, 32'h42908774, 32'h42c464fa, 32'h42b1e4fc, 32'h419a61c4, 32'h40c910da};
test_weights[17832:17839] = '{32'h42510a6b, 32'hc281b30c, 32'h420bb17b, 32'hc27d442c, 32'h422fd160, 32'hc0db5663, 32'hc151eff4, 32'hc2b25837};
test_bias[2229:2229] = '{32'h4207a47a};
test_output[2229:2229] = '{32'hc5aa703d};
test_input[17840:17847] = '{32'hc0beb76d, 32'h428c4c1c, 32'hc28a6c9e, 32'hc29e379f, 32'hc2acf725, 32'h4243024d, 32'hc186d1ee, 32'hc1f758c5};
test_weights[17840:17847] = '{32'hc1c507a0, 32'hc28dc8e8, 32'h41b980ab, 32'hc2a451a1, 32'hc1c8977c, 32'hc21fc188, 32'hc054e1ca, 32'h429a70df};
test_bias[2230:2230] = '{32'hc2980f9f};
test_output[2230:2230] = '{32'hc5045bbe};
test_input[17848:17855] = '{32'h42722f8e, 32'h427626a1, 32'h42348e5e, 32'hc226cbe5, 32'hc2829644, 32'h4285b34a, 32'hc2241cb3, 32'hc293b993};
test_weights[17848:17855] = '{32'h415f600a, 32'h421ce696, 32'h42a30919, 32'h42361142, 32'h42b8da2f, 32'h41afce9b, 32'h4242cb4b, 32'hc27e2e44};
test_bias[2231:2231] = '{32'hc2693518};
test_output[2231:2231] = '{32'h454284c5};
test_input[17856:17863] = '{32'h4247ecbf, 32'hc1e976da, 32'h42031a07, 32'hc2b6c002, 32'hc1cb2847, 32'hc299d98e, 32'h42c69b7c, 32'h41ac0c8c};
test_weights[17856:17863] = '{32'hc0cf6fc0, 32'hc23b66d5, 32'hc2662e5f, 32'h41b2e160, 32'hc20f4b99, 32'h42840dfc, 32'h427f9ce4, 32'h4286de77};
test_bias[2232:2232] = '{32'h42940219};
test_output[2232:2232] = '{32'h444bac3f};
test_input[17864:17871] = '{32'h429c9212, 32'hc17014a3, 32'h4190e0cf, 32'h419ec00c, 32'h40857d30, 32'h41e3f2e6, 32'hc00f17d8, 32'hc1c960c7};
test_weights[17864:17871] = '{32'hc13dc35d, 32'hc29050c3, 32'h41bf434f, 32'hc1ff48c3, 32'hc2623b48, 32'h42c16728, 32'hc2611f67, 32'h428207d0};
test_bias[2233:2233] = '{32'h41f21999};
test_output[2233:2233] = '{32'h44783ca6};
test_input[17872:17879] = '{32'hc2597d7e, 32'hc2a03367, 32'h419747df, 32'h42996699, 32'hc25838e8, 32'hc18aafe4, 32'hc21e6ed5, 32'h42baffa7};
test_weights[17872:17879] = '{32'hc1ba8630, 32'h428a231b, 32'hc2bf6405, 32'h42bbef25, 32'hc220f861, 32'h4218ea8c, 32'h416aae92, 32'h42c65e42};
test_bias[2234:2234] = '{32'hc264ef4d};
test_output[2234:2234] = '{32'h4630443f};
test_input[17880:17887] = '{32'hc275f792, 32'h42a28018, 32'hc21363a5, 32'h42469409, 32'hc1ccc147, 32'hc12ab045, 32'h418d268e, 32'h42b817ec};
test_weights[17880:17887] = '{32'hc29be907, 32'h42601e5f, 32'h42bddd38, 32'hc23a814e, 32'hc2206455, 32'hc2266d4d, 32'hc2bc52e8, 32'hc1487b9e};
test_bias[2235:2235] = '{32'hc2020705};
test_output[2235:2235] = '{32'h4506c2fb};
test_input[17888:17895] = '{32'hc1c61ae5, 32'h42818af2, 32'h42c63ba5, 32'h42503def, 32'h428b1e35, 32'hc2071829, 32'h428df655, 32'h42b177df};
test_weights[17888:17895] = '{32'h4188a99b, 32'hc1a5e958, 32'h4201537c, 32'h42a2c9a4, 32'h41315e68, 32'hc15affd4, 32'h41df5e67, 32'hc13e60a2};
test_bias[2236:2236] = '{32'h4293ec2d};
test_output[2236:2236] = '{32'h45f72891};
test_input[17896:17903] = '{32'h418c2db4, 32'h42c438d9, 32'h42231c16, 32'hc203e406, 32'h42845ad7, 32'hc2801eb4, 32'h429d8901, 32'h40dc3675};
test_weights[17896:17903] = '{32'h42371999, 32'hc23fac98, 32'h42c7975e, 32'h418423c2, 32'hc26cfacf, 32'hc29bc227, 32'h3fd75ad1, 32'hc2910158};
test_bias[2237:2237] = '{32'hc2c422b7};
test_output[2237:2237] = '{32'h43654f72};
test_input[17904:17911] = '{32'h4118e306, 32'h40d1af28, 32'hc275b64e, 32'h426260a0, 32'h41e39e08, 32'h42bc8b29, 32'h42a70160, 32'h41a91b79};
test_weights[17904:17911] = '{32'hc29b5aa7, 32'h4292f53a, 32'hc2b782cb, 32'hc1beacab, 32'h41e672d8, 32'hc2a42d5d, 32'h42528751, 32'h40d8ee23};
test_bias[2238:2238] = '{32'hc2b04d6f};
test_output[2238:2238] = '{32'h44c2b7b7};
test_input[17912:17919] = '{32'hc1f01e88, 32'hc27f55cd, 32'hc2a36cce, 32'hc1e80da9, 32'h42bdadc7, 32'hc2a5c95e, 32'h42233702, 32'h415acf31};
test_weights[17912:17919] = '{32'h42ae5748, 32'hc23ec8da, 32'h42a365fd, 32'h411a4d23, 32'hc06b530a, 32'hc23fdb52, 32'hc267c914, 32'h4191df59};
test_bias[2239:2239] = '{32'hc2a0e3b8};
test_output[2239:2239] = '{32'hc59f3d87};
test_input[17920:17927] = '{32'hc2188e38, 32'h42a895d1, 32'hc2c43e5b, 32'h42481d49, 32'hc2061ce5, 32'h4225131a, 32'h42a1e960, 32'hc1c26e40};
test_weights[17920:17927] = '{32'hc2899500, 32'h42272e71, 32'h42118af6, 32'h41adbaf8, 32'h417fb979, 32'h400669ce, 32'hc113d415, 32'hc1fcb2f3};
test_bias[2240:2240] = '{32'h42c1c711};
test_output[2240:2240] = '{32'h45502440};
test_input[17928:17935] = '{32'hc20e8f20, 32'hc29b3e57, 32'hc1e89fbc, 32'h426a4b44, 32'hc296c696, 32'hc1d96c41, 32'hc1d8d3f9, 32'hc2c74846};
test_weights[17928:17935] = '{32'h42af3c73, 32'hc0be6c4c, 32'h426e061f, 32'hc29eb1ed, 32'hc19167e8, 32'hc1eecef3, 32'hc20b5f49, 32'hc1d2de2a};
test_bias[2241:2241] = '{32'hc20dd693};
test_output[2241:2241] = '{32'hc54f9f15};
test_input[17936:17943] = '{32'hc1d930db, 32'hc279f6b3, 32'h42bcef66, 32'h42632715, 32'h413939fa, 32'h423b6f2c, 32'h424c3004, 32'hc0a50672};
test_weights[17936:17943] = '{32'hc2b28145, 32'hc2b33a45, 32'h4137002a, 32'h4282df3f, 32'hc266d2c5, 32'hc1911aca, 32'hc27c6e63, 32'hc1568fa2};
test_bias[2242:2242] = '{32'hc27b2e76};
test_output[2242:2242] = '{32'h45fcb47a};
test_input[17944:17951] = '{32'hc27c6e26, 32'h4289da82, 32'h401c1edd, 32'hc1156c88, 32'hc2c6d545, 32'hc1c134e1, 32'h42a7429c, 32'h42533625};
test_weights[17944:17951] = '{32'h415e73a1, 32'h4217c8c2, 32'h426d950c, 32'hc1dd2cc5, 32'hc19c46ed, 32'hc29a25eb, 32'h4169d05f, 32'hc2c5449d};
test_bias[2243:2243] = '{32'hc24353ed};
test_output[2243:2243] = '{32'h44eeb8d6};
test_input[17952:17959] = '{32'hc2659b55, 32'hc0206666, 32'hc23edcc3, 32'hc20e9344, 32'hc21e5f47, 32'hc2c3b20d, 32'hc06891af, 32'h4212fda8};
test_weights[17952:17959] = '{32'hc29a2fef, 32'h42927633, 32'h42baba59, 32'h42641fdc, 32'h42acdc2a, 32'hc2bdf35b, 32'hc2c1ffe2, 32'hc298b819};
test_bias[2244:2244] = '{32'h427bef5a};
test_output[2244:2244] = '{32'h449a5244};
test_input[17960:17967] = '{32'h41d364f1, 32'h42c0d435, 32'hc2874f7e, 32'hc21e4da1, 32'hc2821e21, 32'h3e1bd94c, 32'hc2384e3e, 32'hc06aa735};
test_weights[17960:17967] = '{32'hc28fc653, 32'h41cb6f1d, 32'hc1bfcc95, 32'hc26b0b74, 32'h42bd4e8c, 32'h4265cf08, 32'hc28d62e9, 32'h3fbe48a8};
test_bias[2245:2245] = '{32'h424ce695};
test_output[2245:2245] = '{32'h44ceafad};
test_input[17968:17975] = '{32'hc1b9dee0, 32'hc25e3687, 32'h4210384f, 32'hc232293b, 32'h429ead53, 32'hc271cfd5, 32'h422b6a07, 32'hc20982ec};
test_weights[17968:17975] = '{32'h42c278e2, 32'h42c7f40b, 32'h422160dd, 32'h42341e59, 32'h4131aad7, 32'hc1a67d53, 32'hc13cabe8, 32'hc254987d};
test_bias[2246:2246] = '{32'h42bfc4a2};
test_output[2246:2246] = '{32'hc5963b49};
test_input[17976:17983] = '{32'hc28c29a8, 32'hc2c1af92, 32'hc273855c, 32'h42a6fe7c, 32'hc28fcb5e, 32'h4264e104, 32'h4288f1b6, 32'h4274ba7e};
test_weights[17976:17983] = '{32'hc15ecdcb, 32'h42a99dac, 32'h4255351d, 32'hc2849d17, 32'hc147d1d3, 32'hc13c213e, 32'hc23ed75a, 32'h4258905e};
test_bias[2247:2247] = '{32'hc23330b3};
test_output[2247:2247] = '{32'hc676c2a0};
test_input[17984:17991] = '{32'hc1c3b33a, 32'h3fbaaaa4, 32'hc09cd7c5, 32'h429592f9, 32'hc22b45e3, 32'hc1045155, 32'hc28e34cd, 32'h42831787};
test_weights[17984:17991] = '{32'h427ad71f, 32'h41bd98df, 32'hc2125881, 32'hc19f6b84, 32'h42808f7c, 32'hc2348295, 32'hc290f52e, 32'hc175a5e4};
test_bias[2248:2248] = '{32'hc25e5f52};
test_output[2248:2248] = '{32'hc4894315};
test_input[17992:17999] = '{32'h41e061aa, 32'h40a3892e, 32'h42bc5f90, 32'hc219803a, 32'h42a5f35b, 32'h422c6b84, 32'hc1bfa8ce, 32'hc0fbca66};
test_weights[17992:17999] = '{32'h41ca00b9, 32'hc23eb62a, 32'hc2bae94f, 32'h42823590, 32'hc2bef170, 32'h42915d40, 32'hc2b8faaa, 32'hc288b11d};
test_bias[2249:2249] = '{32'hc28452ae};
test_output[2249:2249] = '{32'hc64a2610};
test_input[18000:18007] = '{32'hc2a2e779, 32'hc2ab8827, 32'hc28b8c21, 32'h42b369c9, 32'hc2b94655, 32'hc283f045, 32'hc1f1762e, 32'hc1f0b94c};
test_weights[18000:18007] = '{32'hc20eacb0, 32'hc20989ab, 32'hc19595a2, 32'hc1c73f3b, 32'hc1ffa43e, 32'h42b7c7e4, 32'h414ca9b1, 32'h42c38c44};
test_bias[2250:2250] = '{32'hc262c1c7};
test_output[2250:2250] = '{32'hc4c33a54};
test_input[18008:18015] = '{32'h4290995c, 32'h4254be87, 32'h4292720e, 32'hc2c03263, 32'h41a34389, 32'hc183fa27, 32'h41dfb2c8, 32'hc256b697};
test_weights[18008:18015] = '{32'h41860cd9, 32'hc08f9488, 32'h429220e8, 32'hc1ce2810, 32'h411e687d, 32'hc05b1181, 32'h429f0263, 32'hc25255fe};
test_bias[2251:2251] = '{32'hc299844e};
test_output[2251:2251] = '{32'h465b2ae6};
test_input[18016:18023] = '{32'hc2a2c8d1, 32'h417831b8, 32'hc1e52aaa, 32'h42bc518e, 32'hc235630b, 32'h41919972, 32'h41576d1d, 32'h41a80dcd};
test_weights[18016:18023] = '{32'h4291b942, 32'h42010415, 32'hc17727d9, 32'hc1295962, 32'h40f4b78b, 32'hc29aa7bc, 32'hc2be820d, 32'hc0ca47f4};
test_bias[2252:2252] = '{32'hbfbe350a};
test_output[2252:2252] = '{32'hc60f0c68};
test_input[18024:18031] = '{32'h42892001, 32'h419a885b, 32'hc2abc4dd, 32'h42085b86, 32'hc241ce60, 32'h42c6556e, 32'hc27bd6a3, 32'h4281ebe9};
test_weights[18024:18031] = '{32'hc25df0e7, 32'h42971dec, 32'h4061e682, 32'hc17d6e15, 32'h428bc581, 32'hc2c6e2d0, 32'h41c6c286, 32'hc2ae89df};
test_bias[2253:2253] = '{32'h41e62363};
test_output[2253:2253] = '{32'hc6b8afae};
test_input[18032:18039] = '{32'hc250acae, 32'hc2680d8a, 32'h42a1ea1c, 32'hc28fa5b7, 32'hc14fd544, 32'h42a6f944, 32'hc15b3c0d, 32'h42746dd7};
test_weights[18032:18039] = '{32'h42be61cc, 32'hc2256aac, 32'h420db536, 32'h42b1bcc6, 32'hc28a09d7, 32'h423de55b, 32'h42c6db5a, 32'h41ca1691};
test_bias[2254:2254] = '{32'h4292a346};
test_output[2254:2254] = '{32'hc471c9cb};
test_input[18040:18047] = '{32'hc25c4218, 32'h42a1bd03, 32'hc265f3be, 32'h41fb7cb3, 32'h42a1b44e, 32'hc29342f0, 32'hc23fea60, 32'hc21a88d1};
test_weights[18040:18047] = '{32'hc2192f0b, 32'hc1dfb55e, 32'h426e35e0, 32'h41a3719c, 32'hc2476e3d, 32'hc12fed72, 32'h40644356, 32'h42267f8e};
test_bias[2255:2255] = '{32'h420df275};
test_output[2255:2255] = '{32'hc5f6d986};
test_input[18048:18055] = '{32'hc2ab0f9e, 32'hc28db3d4, 32'hc27a74f8, 32'hc0848ee9, 32'h42b5ccb2, 32'h428ca178, 32'hc2c4b903, 32'h42c377b1};
test_weights[18048:18055] = '{32'hc2a0fd8f, 32'hc21a16ec, 32'hc28e5d14, 32'hc2c0ba73, 32'hc200d0e4, 32'h4202e059, 32'h42420375, 32'h414b9166};
test_bias[2256:2256] = '{32'hc24c77af};
test_output[2256:2256] = '{32'h46206492};
test_input[18056:18063] = '{32'hc223a961, 32'hc28a0996, 32'h42b0c641, 32'hc1e4d6b7, 32'hc28bed5c, 32'hc1f6a856, 32'hc239de38, 32'hc242a68f};
test_weights[18056:18063] = '{32'h40971b6f, 32'h415f30f7, 32'hc228f022, 32'hc13cebd4, 32'hc21caf9b, 32'h42c58dfa, 32'h4286ea68, 32'hc299042c};
test_bias[2257:2257] = '{32'h42178657};
test_output[2257:2257] = '{32'hc5842e03};
test_input[18064:18071] = '{32'h41af8417, 32'hc2b07bba, 32'hc2825260, 32'hc27a7736, 32'h42ab600b, 32'h4245d3ee, 32'hc2a14034, 32'h408b70e9};
test_weights[18064:18071] = '{32'h4223cb48, 32'hc2adbdc2, 32'hc1d70d34, 32'hc275befb, 32'h42b2737f, 32'hc1d46c02, 32'h4208965b, 32'hc26011c7};
test_bias[2258:2258] = '{32'hc2194c21};
test_output[2258:2258] = '{32'h468866aa};
test_input[18072:18079] = '{32'h422d8137, 32'h42b2f314, 32'h42509721, 32'hc2ab551a, 32'h42694a2d, 32'hc0897820, 32'hc2920abf, 32'hc18178f3};
test_weights[18072:18079] = '{32'h42b394c7, 32'h4287bd00, 32'h41b211a1, 32'hc229bd46, 32'hc2af77f7, 32'h42a0c158, 32'h428db76e, 32'hc29c6628};
test_bias[2259:2259] = '{32'h42c7ee92};
test_output[2259:2259] = '{32'h45aba466};
test_input[18080:18087] = '{32'hc078472b, 32'h424044d1, 32'hc1db251e, 32'hc2a0b947, 32'hc08aacab, 32'hc12b4f18, 32'h428399b9, 32'hc19e7ca3};
test_weights[18080:18087] = '{32'hc28d3c82, 32'hc212ef1e, 32'hc2ae58cd, 32'h42801d42, 32'hc2c50f91, 32'hc251799c, 32'h42966291, 32'hc2bbaab1};
test_bias[2260:2260] = '{32'hc2569cfd};
test_output[2260:2260] = '{32'h455a11e8};
test_input[18088:18095] = '{32'hc12079a4, 32'hc2b3fb00, 32'hc25b1c0d, 32'h424eeaf4, 32'hc0279fc6, 32'hc28ebcf6, 32'hc1f29043, 32'hc2204a36};
test_weights[18088:18095] = '{32'h423ac2b2, 32'hc18deb37, 32'hc21e6f52, 32'h423fc511, 32'h4241ea4e, 32'h421b5004, 32'hc2a3a967, 32'hc2a11b11};
test_bias[2261:2261] = '{32'h426ca1be};
test_output[2261:2261] = '{32'h46071fed};
test_input[18096:18103] = '{32'h41c55de6, 32'hc213ebb7, 32'hc22644dd, 32'h42066ac4, 32'hc11fdfd7, 32'h4237de17, 32'hc2b8fad5, 32'h42913295};
test_weights[18096:18103] = '{32'hc1aee3e1, 32'h42a980b8, 32'h4290e125, 32'h41dca033, 32'hc2281a0b, 32'h42be1aff, 32'hc2b80ebe, 32'h41ac5fa6};
test_bias[2262:2262] = '{32'h429ad4d5};
test_output[2262:2262] = '{32'h460f8322};
test_input[18104:18111] = '{32'h42a49d9e, 32'h41cebc61, 32'h42abde93, 32'h421d0722, 32'h41ccf63f, 32'hc2527cf3, 32'hc200a13c, 32'h42668584};
test_weights[18104:18111] = '{32'hc2bba43d, 32'hc1bd9911, 32'hc2bc3069, 32'h42739477, 32'h42008720, 32'h4217e5a9, 32'hc1dddf3a, 32'hc24b3b54};
test_bias[2263:2263] = '{32'hc29dec13};
test_output[2263:2263] = '{32'hc68750a0};
test_input[18112:18119] = '{32'hc2c48b41, 32'h42aaa124, 32'hbfbbb6de, 32'h40ff032c, 32'hc27fbcf8, 32'h42b85b68, 32'hc25daddb, 32'h427797a5};
test_weights[18112:18119] = '{32'h4148f306, 32'h42085dbb, 32'hc1bb890f, 32'h4254f010, 32'h42aa6790, 32'h420f53d2, 32'hc18a66eb, 32'h42c19436};
test_bias[2264:2264] = '{32'hc255eb2a};
test_output[2264:2264] = '{32'h45d726a4};
test_input[18120:18127] = '{32'h41af4702, 32'h418b7b16, 32'hc222332f, 32'hc270819a, 32'h41bef924, 32'h418e38c8, 32'hc2b42b81, 32'hc0c5cf76};
test_weights[18120:18127] = '{32'h42294991, 32'h429aa9ec, 32'hc1d6b4de, 32'hc185f4e3, 32'h42644f09, 32'hc0ac223d, 32'hc26ffd56, 32'hc2b676c3};
test_bias[2265:2265] = '{32'h42be4808};
test_output[2265:2265] = '{32'h4636d5f8};
test_input[18128:18135] = '{32'h4295b121, 32'hc1c38901, 32'h4250da69, 32'h42660c6f, 32'h4114f4e1, 32'h41a50982, 32'hc2533580, 32'h4225d6f7};
test_weights[18128:18135] = '{32'h42a7e0c3, 32'h428a5668, 32'hc26e8b9b, 32'hc27547e4, 32'hc276ff43, 32'hc222536d, 32'hc2c1e096, 32'hc078e78a};
test_bias[2266:2266] = '{32'hc21d3cb7};
test_output[2266:2266] = '{32'h44b62c4f};
test_input[18136:18143] = '{32'hc2251f59, 32'hc23d5a4f, 32'h4279ee0c, 32'h41285f45, 32'hc2b1d215, 32'h41d915ea, 32'h4276db05, 32'hc2bfcdcf};
test_weights[18136:18143] = '{32'h42824470, 32'h42a626df, 32'hc20e70d0, 32'h424157a4, 32'hc2816209, 32'hc1aff213, 32'hc237eb6e, 32'h42bd7678};
test_bias[2267:2267] = '{32'h416fae39};
test_output[2267:2267] = '{32'hc66bc992};
test_input[18144:18151] = '{32'hc190db7c, 32'hc209337c, 32'h41d5ce55, 32'h4107b487, 32'h41eb6f35, 32'h41f5b5d4, 32'hc1884332, 32'h415addbd};
test_weights[18144:18151] = '{32'h4191f2c5, 32'hc1d772cb, 32'hc2aa3e10, 32'h41497299, 32'hc13be8d7, 32'h429c4596, 32'h41ea67d3, 32'hc29d126b};
test_bias[2268:2268] = '{32'hc2bc3461};
test_output[2268:2268] = '{32'hc4947fdc};
test_input[18152:18159] = '{32'h41f0ff78, 32'h40f66bac, 32'hc1878df9, 32'hc1a049b0, 32'hc241205c, 32'h42b7845e, 32'h42a3c5c3, 32'h42872b6c};
test_weights[18152:18159] = '{32'h4221c7ba, 32'h411a1e1d, 32'hc1914984, 32'h41be3fb8, 32'hc0fbf0e0, 32'hc00fcc24, 32'hc2639599, 32'hc27c6c4a};
test_bias[2269:2269] = '{32'h42862ad1};
test_output[2269:2269] = '{32'hc5ec3912};
test_input[18160:18167] = '{32'h428b4543, 32'hc2ad97bc, 32'h42b3b5e4, 32'h426d337d, 32'hc201ab89, 32'h42262368, 32'h42b2f13e, 32'hc1342b59};
test_weights[18160:18167] = '{32'h418f8560, 32'hc2782f95, 32'hc296489c, 32'hc2ad896e, 32'h429638f8, 32'h41b1b43c, 32'h425607ad, 32'h427b4658};
test_bias[2270:2270] = '{32'h419d0f33};
test_output[2270:2270] = '{32'hc5273487};
test_input[18168:18175] = '{32'h41cf0e7f, 32'h423f795e, 32'hc297995e, 32'hc1eaf4d7, 32'h4212b3cc, 32'h42c17b19, 32'hc2b4156e, 32'hc2befe5b};
test_weights[18168:18175] = '{32'hc21dda01, 32'hc26f8d64, 32'h419a5d0d, 32'hc2b35891, 32'hc29e4c60, 32'hc014c134, 32'hc2bd8054, 32'h41db1c6d};
test_bias[2271:2271] = '{32'h4026b91b};
test_output[2271:2271] = '{32'h4293a2dc};
test_input[18176:18183] = '{32'h42bee00d, 32'hc23f3a25, 32'hc23ec9d4, 32'h40e2ef22, 32'hc02a2b1e, 32'hc22f3a5e, 32'hc18a7846, 32'h41f18f5e};
test_weights[18176:18183] = '{32'hbf2a9ea0, 32'h42a6ecf7, 32'hc259c946, 32'h428b71cd, 32'h40f36ec8, 32'h42b1a2e5, 32'h42a06cce, 32'h3fd27aec};
test_bias[2272:2272] = '{32'hc232be77};
test_output[2272:2272] = '{32'hc5c38665};
test_input[18184:18191] = '{32'hc29004d2, 32'hc299d297, 32'hc1f64f2e, 32'hc29f5383, 32'h414efb6f, 32'hc1100e26, 32'h422f67f9, 32'h422b33a6};
test_weights[18184:18191] = '{32'h41c16546, 32'h42c663ce, 32'hc2aa7372, 32'h42a52772, 32'hc206fbf5, 32'h42965e78, 32'h41b54ecb, 32'h410524c9};
test_bias[2273:2273] = '{32'h42937add};
test_output[2273:2273] = '{32'hc64b586d};
test_input[18192:18199] = '{32'h420bbd0b, 32'hc2b62001, 32'hc2220f12, 32'h4246dcb9, 32'h42a026fb, 32'hc28d67c2, 32'hc2a9f07f, 32'h4281ee83};
test_weights[18192:18199] = '{32'hc2be1cb2, 32'h42267d0f, 32'h421dcd47, 32'h3f6d4667, 32'h3fbca022, 32'h428d0758, 32'h424c47b0, 32'h41b516ae};
test_bias[2274:2274] = '{32'hc2c31ae1};
test_output[2274:2274] = '{32'hc680e248};
test_input[18200:18207] = '{32'hc2c7dfb1, 32'hc127a2e3, 32'h428e3bd7, 32'hc2b001c1, 32'h422b1480, 32'hc2411521, 32'hc285c6b2, 32'hc29c7af2};
test_weights[18200:18207] = '{32'hc2a51f61, 32'hbe34f631, 32'hc0983f80, 32'h4247ff99, 32'hc24426b4, 32'hc1150f59, 32'h40507812, 32'hc1b41249};
test_bias[2275:2275] = '{32'h428fbddc};
test_output[2275:2275] = '{32'h45599ba1};
test_input[18208:18215] = '{32'hc27d1d8b, 32'h4283eb6c, 32'h428b5b5e, 32'h41258b7e, 32'h41854f62, 32'hc2aff1cd, 32'h420fc896, 32'h4236dec5};
test_weights[18208:18215] = '{32'h41b3cf8c, 32'hc1ffd5c2, 32'h421a788b, 32'h4232f886, 32'hc29bf3a1, 32'h42b24a48, 32'h41ab04ec, 32'h4221118c};
test_bias[2276:2276] = '{32'h426df19b};
test_output[2276:2276] = '{32'hc5d615af};
test_input[18216:18223] = '{32'hc22a2eeb, 32'h42478d5e, 32'hc262740d, 32'hc1e9233c, 32'h42a6a49c, 32'hc2b7bba8, 32'hc27fc739, 32'h420da265};
test_weights[18216:18223] = '{32'h429a7a2f, 32'hc2414254, 32'hc26544c0, 32'h423a7d34, 32'hc255606a, 32'hc28536bb, 32'hc29c5ead, 32'hc26f1de6};
test_bias[2277:2277] = '{32'hc23da0ff};
test_output[2277:2277] = '{32'h442ed669};
test_input[18224:18231] = '{32'h4204c988, 32'h41406dc1, 32'h41c29622, 32'hc22510ef, 32'hc2c26412, 32'h419a120a, 32'hc2c3cd2d, 32'h4291f0d2};
test_weights[18224:18231] = '{32'h425740b6, 32'h411f0742, 32'hc260dfdc, 32'h420afd68, 32'h42b307dc, 32'h422bdc30, 32'hc1abcedb, 32'hc29b0172};
test_bias[2278:2278] = '{32'hc24662eb};
test_output[2278:2278] = '{32'hc6414b8a};
test_input[18232:18239] = '{32'hc29ed89e, 32'hc2985c05, 32'h42b9a390, 32'hc293bedf, 32'h42260832, 32'h42941341, 32'hc242d3a5, 32'hc2524a53};
test_weights[18232:18239] = '{32'hc1975f67, 32'hc2c0d655, 32'hc2287f91, 32'h41ee7de4, 32'hc2b56015, 32'hc29ca2df, 32'h4200f314, 32'hc2abb0f8};
test_bias[2279:2279] = '{32'hc2636cb6};
test_output[2279:2279] = '{32'hc5764efc};
test_input[18240:18247] = '{32'hc1b71ed7, 32'hc08f8809, 32'hc13f5bec, 32'hc294ea5e, 32'h42807fbd, 32'h428aae9a, 32'hc062e483, 32'hc23192d2};
test_weights[18240:18247] = '{32'hc2371d1a, 32'hc20262b3, 32'h407b6d7c, 32'h42a0d5ce, 32'h3fae0ab5, 32'h4184773d, 32'hc2a011da, 32'h421ab4c4};
test_bias[2280:2280] = '{32'h422d9179};
test_output[2280:2280] = '{32'hc59c1794};
test_input[18248:18255] = '{32'h427f5766, 32'h4008f6f5, 32'h400f4f9b, 32'h4271b6bf, 32'h429a2d01, 32'h41dead33, 32'h42974bd4, 32'hc24b19e1};
test_weights[18248:18255] = '{32'hc29eb5e8, 32'h41c65e46, 32'h419b463c, 32'hc1dee7a4, 32'h42a8f54a, 32'h428d0409, 32'h42136a00, 32'h42b95b69};
test_bias[2281:2281] = '{32'h42b1a1ab};
test_output[2281:2281] = '{32'hc0e2033e};
test_input[18256:18263] = '{32'h420a7886, 32'hc21398bb, 32'h420adb65, 32'hc1c37378, 32'h41aa6c59, 32'h424ede76, 32'hc24357f9, 32'h42a02e8a};
test_weights[18256:18263] = '{32'h4294f09d, 32'h41ea5f4c, 32'h413a2b2a, 32'h421f8bc7, 32'h42bd1d47, 32'hc23d8298, 32'hc25f71b0, 32'h4226373b};
test_bias[2282:2282] = '{32'h42b74937};
test_output[2282:2282] = '{32'h45cf721c};
test_input[18264:18271] = '{32'hc20beb1a, 32'h40807eaa, 32'h4263dbd4, 32'h429a7243, 32'h40ae163b, 32'h42aa7c6a, 32'hc00954ef, 32'h42acea8b};
test_weights[18264:18271] = '{32'hc13bb602, 32'h42b26163, 32'h4233d721, 32'hc20cc474, 32'hc20f4d81, 32'hc1a494c1, 32'h422ad84f, 32'h4233ffbd};
test_bias[2283:2283] = '{32'h41f88985};
test_output[2283:2283] = '{32'h451bd774};
test_input[18272:18279] = '{32'hc1ed08f7, 32'hbd1e245b, 32'h42b31c27, 32'h42433161, 32'h41881ee9, 32'hc1f02183, 32'h421548f9, 32'h429fd021};
test_weights[18272:18279] = '{32'hc29b8092, 32'hc2164bbb, 32'hc1a0dfc8, 32'h42ab238b, 32'hc28d52f7, 32'h41e19b25, 32'hc07483b4, 32'hc20fdc28};
test_bias[2284:2284] = '{32'h42500757};
test_output[2284:2284] = '{32'hc3a6a6e8};
test_input[18280:18287] = '{32'hc19af791, 32'h42b23410, 32'h42a15069, 32'hc1b9286c, 32'hc267edb3, 32'h42875e68, 32'h429377d7, 32'h41fb52a0};
test_weights[18280:18287] = '{32'hc1bc21ce, 32'h41caf009, 32'h427a564a, 32'hc17c7482, 32'hc1e388f7, 32'h42a9ecdd, 32'h425ddeef, 32'h4264401d};
test_bias[2285:2285] = '{32'hc27e7b60};
test_output[2285:2285] = '{32'h46a6c6fb};
test_input[18288:18295] = '{32'hc29b4312, 32'hc2ae49e8, 32'h429b5f5c, 32'hc14646d2, 32'hc2127f6c, 32'hc0b8c290, 32'hc2b1e3a6, 32'h4200f16a};
test_weights[18288:18295] = '{32'h4268cec3, 32'hc0562d37, 32'h42309dfe, 32'hc2c29600, 32'hc2393f09, 32'hc11846f4, 32'hc2b69436, 32'h41c7fa68};
test_bias[2286:2286] = '{32'h41ce0774};
test_output[2286:2286] = '{32'h462d9e4b};
test_input[18296:18303] = '{32'hc27a95d0, 32'hc28d944a, 32'h4104df1d, 32'h4188664b, 32'hc24801a5, 32'hc2a58ba2, 32'h426b742c, 32'h4298bb96};
test_weights[18296:18303] = '{32'h413c007b, 32'hc289aba5, 32'hc03540fb, 32'h42783fb9, 32'h42865ff5, 32'hc22eba32, 32'h422fe16f, 32'h421c4c4f};
test_bias[2287:2287] = '{32'hc21ec507};
test_output[2287:2287] = '{32'h462b4043};
test_input[18304:18311] = '{32'h42501a54, 32'h42669904, 32'h427e1beb, 32'hc1caa102, 32'h41048988, 32'hc2a6c79a, 32'hc143d185, 32'hc29564ba};
test_weights[18304:18311] = '{32'hc2b6d845, 32'h40b50d3f, 32'h42349d8f, 32'hc2bbc0fc, 32'h423e646e, 32'h429868c8, 32'hc21d8fca, 32'h41a9216b};
test_bias[2288:2288] = '{32'h400dbcc3};
test_output[2288:2288] = '{32'hc5c2f957};
test_input[18312:18319] = '{32'h410ad6d0, 32'hc1c524ad, 32'hc1822796, 32'h41e3e13e, 32'h3fe655d3, 32'hc0be5bb0, 32'hc2bb6fab, 32'hc10c03bc};
test_weights[18312:18319] = '{32'h42790a83, 32'hc257934a, 32'h412b909d, 32'h42b24a7a, 32'hc2af6345, 32'h4276409d, 32'hc182d2c2, 32'h42918b88};
test_bias[2289:2289] = '{32'hc258a0cf};
test_output[2289:2289] = '{32'h458e362b};
test_input[18320:18327] = '{32'hc1c6e268, 32'h410c8e30, 32'hc28aa1a9, 32'hc203a816, 32'hc25b3af4, 32'h421b81de, 32'hc201bf9b, 32'h4229ad2c};
test_weights[18320:18327] = '{32'hc2acc102, 32'hc2a263cc, 32'hc11a0b2c, 32'hc2150b9a, 32'h405798b3, 32'hc1e7fe53, 32'hc2734ff3, 32'hc04bd62c};
test_bias[2290:2290] = '{32'h41b00387};
test_output[2290:2290] = '{32'h45723d7d};
test_input[18328:18335] = '{32'h4290da3d, 32'h42b63e37, 32'h422f8acf, 32'hc2864fe2, 32'hc2910cee, 32'hc1585e91, 32'h41d2e57b, 32'h4120563c};
test_weights[18328:18335] = '{32'hc29c76ef, 32'hbf819add, 32'h3f09f01d, 32'h420bae98, 32'h41e8ba39, 32'h406ea83b, 32'hc0c9880a, 32'hbf4300c8};
test_bias[2291:2291] = '{32'hc28aa7d8};
test_output[2291:2291] = '{32'hc623cc35};
test_input[18336:18343] = '{32'h429c786f, 32'h3e80eb2d, 32'hc2968948, 32'h4299ccfa, 32'h4195d4a1, 32'h42567919, 32'hc270250c, 32'h42ae76f7};
test_weights[18336:18343] = '{32'h4193bd36, 32'hc2903d09, 32'h41a1cfb7, 32'h42a3c424, 32'hc2a70b86, 32'h42bcc06a, 32'h42580341, 32'h42b233e1};
test_bias[2292:2292] = '{32'h42673489};
test_output[2292:2292] = '{32'h465f34f3};
test_input[18344:18351] = '{32'hc07c3a19, 32'h42aec24d, 32'hc2a80a8c, 32'h41c44692, 32'h4192e111, 32'hc25abf27, 32'hc1b71e2f, 32'hc17459c4};
test_weights[18344:18351] = '{32'hc26bc4cd, 32'h42b37a1b, 32'hc23522ac, 32'h421705e0, 32'h42af915a, 32'hc1d9e2f1, 32'h42531902, 32'hc280a764};
test_bias[2293:2293] = '{32'h420eeb4d};
test_output[2293:2293] = '{32'h46758fda};
test_input[18352:18359] = '{32'h42a88528, 32'hc214ff4c, 32'h42ba090c, 32'hc2bddfc7, 32'h4198f8a6, 32'h42a81043, 32'hc25d747e, 32'hc1cdd80f};
test_weights[18352:18359] = '{32'hc22f18d7, 32'hc2a75b07, 32'h428c4aed, 32'h4202afc5, 32'hc29d87b0, 32'hc11b7c93, 32'h41b52bba, 32'hc2237feb};
test_bias[2294:2294] = '{32'h42a8a4d4};
test_output[2294:2294] = '{32'h43cd95fa};
test_input[18360:18367] = '{32'hc133a6a1, 32'h3f90d175, 32'hc2bd3b65, 32'h42a6a542, 32'h421a5c08, 32'hc29e5212, 32'hc1ba975e, 32'hc2a52dfc};
test_weights[18360:18367] = '{32'hc28df92d, 32'hc20f3ca0, 32'h42a98967, 32'h426e1bb6, 32'hc192eb4d, 32'hc2ad3a38, 32'h41e4edcb, 32'h40b1f3a1};
test_bias[2295:2295] = '{32'hc257b1da};
test_output[2295:2295] = '{32'h45267138};
test_input[18368:18375] = '{32'hc0c84bf8, 32'hc04f572a, 32'hc1da5954, 32'h4279d144, 32'hc18dd8c6, 32'hc2c78e53, 32'h422c22b2, 32'h41e4d3e0};
test_weights[18368:18375] = '{32'h4264e8ee, 32'hc1c9fbf6, 32'hc2bd00ec, 32'hc29e828f, 32'hc1fb4254, 32'hc28f673c, 32'hc27956c2, 32'h42040ed4};
test_bias[2296:2296] = '{32'h42721b57};
test_output[2296:2296] = '{32'h4553a8ac};
test_input[18376:18383] = '{32'h41023811, 32'hc2862535, 32'hc27fafc7, 32'h42b99faa, 32'hc27dea76, 32'h41ce7a2d, 32'hc25f269b, 32'h4213ac46};
test_weights[18376:18383] = '{32'hc23b94e1, 32'h41e91505, 32'h42717b4b, 32'hc191167e, 32'h429c3bf0, 32'hc0fb291a, 32'hc2aad7bc, 32'hc2a2219e};
test_bias[2297:2297] = '{32'h418af14a};
test_output[2297:2297] = '{32'hc62fc593};
test_input[18384:18391] = '{32'hc29fe1b4, 32'h42364d93, 32'h42487642, 32'h41dbf33e, 32'h428da325, 32'hc1f3e495, 32'hc2b5b4e3, 32'hc0d7b547};
test_weights[18384:18391] = '{32'hc1c88544, 32'hc23acca5, 32'hc29eb0fa, 32'hc0f55d30, 32'h422e6b39, 32'hc20387ba, 32'h4258b072, 32'h42c6292c};
test_bias[2298:2298] = '{32'hc279ee2a};
test_output[2298:2298] = '{32'hc5b78c23};
test_input[18392:18399] = '{32'hc26c7799, 32'hbf160a52, 32'hc1b357aa, 32'h4188e050, 32'h41c508e2, 32'h424d1349, 32'h42ac4a22, 32'h41072c66};
test_weights[18392:18399] = '{32'hc1718c6d, 32'h42001e51, 32'h428e837d, 32'hc2b792b9, 32'hc03df578, 32'h42536f6a, 32'hc269c04d, 32'h41ae5c4c};
test_bias[2299:2299] = '{32'hc22b7cd0};
test_output[2299:2299] = '{32'hc58e30b8};
test_input[18400:18407] = '{32'h413bdb83, 32'h41a38873, 32'h422c7c9d, 32'hbd468d9d, 32'h4080dd9e, 32'hc256a6ac, 32'h41a8d084, 32'hc140592e};
test_weights[18400:18407] = '{32'h429384b9, 32'hc2b42850, 32'hc1925ecc, 32'h42651ce0, 32'hc2b2e237, 32'hc2bcfb3e, 32'hbf26361e, 32'hc2c5ada5};
test_bias[2300:2300] = '{32'h42981154};
test_output[2300:2300] = '{32'h45830f53};
test_input[18408:18415] = '{32'hc1a6c79e, 32'h426298a2, 32'hbf226f75, 32'h42a156b3, 32'hc28777d5, 32'hc230d27f, 32'hc1a33bd0, 32'hc2b1f84f};
test_weights[18408:18415] = '{32'h4193aeef, 32'h4299d374, 32'hc2135f4e, 32'hc2929987, 32'hc2c29318, 32'hc1ddfc40, 32'h42980e1c, 32'h3ff7a06e};
test_bias[2301:2301] = '{32'h4259f6a8};
test_output[2301:2301] = '{32'h45842ef1};
test_input[18416:18423] = '{32'h42a0af17, 32'hc1edcc2d, 32'h428e71f5, 32'h429ad892, 32'hc22340c9, 32'h41225c84, 32'h420db6a5, 32'h3f53480f};
test_weights[18416:18423] = '{32'h425d999c, 32'hbe3f2e73, 32'hc0858e8f, 32'h4291e70c, 32'hc2be6737, 32'hc2b2e917, 32'h42940078, 32'h42a92efc};
test_bias[2302:2302] = '{32'h429170e4};
test_output[2302:2302] = '{32'h4672f55e};
test_input[18424:18431] = '{32'h4188d02b, 32'hc2024b26, 32'h42c78ac2, 32'hc220b976, 32'hc13c5c19, 32'hc1ff44a9, 32'hc2667be4, 32'h42a6e907};
test_weights[18424:18431] = '{32'hc1a8793b, 32'hc2a8ab8e, 32'h42888994, 32'hc242c0c2, 32'hbfe01985, 32'h412e9a98, 32'h42bef350, 32'h4200cf45};
test_bias[2303:2303] = '{32'h426df0f5};
test_output[2303:2303] = '{32'h45fc43e1};
test_input[18432:18439] = '{32'h42c185fa, 32'hc1959bf2, 32'h42baa067, 32'hc29df370, 32'hc1b6df2c, 32'hc28f1609, 32'h40d5cc91, 32'hc20ab772};
test_weights[18432:18439] = '{32'hc11fc0b8, 32'hc1c6d622, 32'h3efe98f5, 32'h42a959ec, 32'hc2c48823, 32'hc2862a65, 32'hc2b706f0, 32'h429727c9};
test_bias[2304:2304] = '{32'h422ead38};
test_output[2304:2304] = '{32'hc54d55e4};
test_input[18440:18447] = '{32'h420a5e08, 32'hc297500a, 32'hc2916d2c, 32'h41b09c51, 32'h4296e951, 32'h418cbeeb, 32'hc24e2f63, 32'h420a9220};
test_weights[18440:18447] = '{32'h421f1843, 32'hc2615cb0, 32'h42c47f78, 32'h41eb080b, 32'h3fd8c2d8, 32'h421086ea, 32'h42b4955f, 32'hc23b619d};
test_bias[2305:2305] = '{32'hc1f26130};
test_output[2305:2305] = '{32'hc5c807a2};
test_input[18448:18455] = '{32'h4288fb8d, 32'hc20994ff, 32'hc29e18ba, 32'hc2c45e7d, 32'hc2877925, 32'h428661cf, 32'h415ee4fe, 32'h4205bf04};
test_weights[18448:18455] = '{32'hc2bb9a5d, 32'h429da14b, 32'h423bd2ed, 32'hc176dec9, 32'h4280d210, 32'h41c6bf0f, 32'h42c4d1f5, 32'h42b50aaa};
test_bias[2306:2306] = '{32'h419353c8};
test_output[2306:2306] = '{32'hc61627d6};
test_input[18456:18463] = '{32'h42be9de9, 32'h425d2623, 32'h42c2943e, 32'hc2608b37, 32'hc192a9af, 32'hc2345c1a, 32'hc268f697, 32'hc2350833};
test_weights[18456:18463] = '{32'h41a1ede5, 32'h424e74c5, 32'h40f5fc93, 32'h41f3d924, 32'hc120a690, 32'h414cc310, 32'hc1cf8c55, 32'hc254d8e6};
test_bias[2307:2307] = '{32'hc2ad3a0a};
test_output[2307:2307] = '{32'h45e2d986};
test_input[18464:18471] = '{32'hc2199ba0, 32'h42103c77, 32'hc0b26222, 32'h4231e0b6, 32'h414686e2, 32'h41d5332e, 32'hc262662a, 32'hc267f040};
test_weights[18464:18471] = '{32'hc2ba9ae0, 32'hc2314a43, 32'hc20275e2, 32'hc09f9978, 32'hc189d098, 32'hc26ab1e8, 32'h42a5c58e, 32'hc16219a0};
test_bias[2308:2308] = '{32'h420488be};
test_output[2308:2308] = '{32'hc565766b};
test_input[18472:18479] = '{32'hc24e241e, 32'hc1e73286, 32'hc22c7cef, 32'hc1f8691a, 32'h425a76d6, 32'h41a0ed09, 32'h4287bd0d, 32'h4215b40f};
test_weights[18472:18479] = '{32'hc1f5dd68, 32'h42167bf8, 32'h428bb6e0, 32'h4227dd04, 32'hc1b986a2, 32'h42906435, 32'hc2aea35c, 32'hc0eef3e6};
test_bias[2309:2309] = '{32'h41ff0903};
test_output[2309:2309] = '{32'hc6193c3b};
test_input[18480:18487] = '{32'h41c809ad, 32'h41f79986, 32'hc29281c5, 32'h42afca1d, 32'h4261ec9d, 32'hc2110ff7, 32'h418fbdcd, 32'hc271c50d};
test_weights[18480:18487] = '{32'hc1ab45b1, 32'h428affd3, 32'hbeca5d53, 32'hc2b5a1c4, 32'h42917bb1, 32'hc0adc3d4, 32'hc2779964, 32'h42506e0c};
test_bias[2310:2310] = '{32'hc230dd1d};
test_output[2310:2310] = '{32'hc5c61090};
test_input[18488:18495] = '{32'hc2a958e1, 32'hc1d927c6, 32'hc12735ec, 32'hc234e2e7, 32'hc24b1548, 32'h419a08bb, 32'hc2a57ae3, 32'hc27ec2dd};
test_weights[18488:18495] = '{32'hc299be8f, 32'hc20c6441, 32'h42aaeca1, 32'hc28ec250, 32'h42a2c844, 32'hc2bed6f5, 32'hc1784519, 32'h424eab94};
test_bias[2311:2311] = '{32'h41953cb1};
test_output[2311:2311] = '{32'h44e5d90a};
test_input[18496:18503] = '{32'hc1d42489, 32'hc267cb8d, 32'h42a91ccb, 32'h425ba3fd, 32'h4078e2fe, 32'hc2a04779, 32'h42611c98, 32'hc2925875};
test_weights[18496:18503] = '{32'hc29c4582, 32'hc25b61ae, 32'h4297b4f1, 32'hc22c626f, 32'hc2b85017, 32'hc1cf2172, 32'h402234bb, 32'h4225b8c4};
test_bias[2312:2312] = '{32'hc2bc3d0f};
test_output[2312:2312] = '{32'h45faf937};
test_input[18504:18511] = '{32'hc23d5085, 32'h4231725f, 32'h412b379a, 32'hc1654748, 32'hc287d6ac, 32'h424e2400, 32'hc24f5cf6, 32'hc1b907c4};
test_weights[18504:18511] = '{32'h42079f52, 32'hc294a913, 32'h425c51ef, 32'hc12ae693, 32'hc2415af5, 32'h42be97a8, 32'hc2a7997d, 32'h4293e1e9};
test_bias[2313:2313] = '{32'hc211f9d6};
test_output[2313:2313] = '{32'h45cf4173};
test_input[18512:18519] = '{32'hc2a6e276, 32'h42a88050, 32'h4215c7c9, 32'hc15596e5, 32'hc292aa31, 32'h423cf260, 32'hc144db27, 32'h421a77ec};
test_weights[18512:18519] = '{32'hc220aefd, 32'h42291ed7, 32'hc2894ad9, 32'h42bf7649, 32'h4278c681, 32'h428ad6b0, 32'h42c534ff, 32'h41764fb8};
test_bias[2314:2314] = '{32'hc111dcf9};
test_output[2314:2314] = '{32'h449085f4};
test_input[18520:18527] = '{32'h4063db14, 32'hc2b46c37, 32'hc13d0f9c, 32'h41f3ba61, 32'h41a960aa, 32'h3ff0ed13, 32'h425c6067, 32'h424e21e5};
test_weights[18520:18527] = '{32'hc221e715, 32'hc252e6ff, 32'h42221685, 32'hc2248aa9, 32'h3f9a8ad4, 32'h423de122, 32'hc21a2d36, 32'h40835275};
test_bias[2315:2315] = '{32'hc25200c1};
test_output[2315:2315] = '{32'h4480d413};
test_input[18528:18535] = '{32'hc2a24382, 32'h4285c34a, 32'h42b915b1, 32'hc204ae52, 32'h4255f233, 32'h42b9ba18, 32'hc2c5a174, 32'h3f6146b6};
test_weights[18528:18535] = '{32'hc284b78b, 32'h423b5079, 32'hc281fbe0, 32'h42bddcd9, 32'h40af4ff2, 32'h428d39c5, 32'hc1acf7f7, 32'h42ad2c50};
test_bias[2316:2316] = '{32'hc20a2d6d};
test_output[2316:2316] = '{32'h4602f37a};
test_input[18536:18543] = '{32'h420e475a, 32'h429512e4, 32'h429969aa, 32'hc1f19f8a, 32'h416fa69d, 32'hc186775d, 32'h40b63367, 32'h42b7ab34};
test_weights[18536:18543] = '{32'hc22c26c7, 32'hc2b3b27b, 32'h42892e5e, 32'h423f5eb8, 32'hc2b369b8, 32'h41b7ec79, 32'h42a901ec, 32'hc2686f7d};
test_bias[2317:2317] = '{32'h417528d6};
test_output[2317:2317] = '{32'hc62b9617};
test_input[18544:18551] = '{32'h41121c4d, 32'hc29b5c43, 32'h41d06379, 32'h4237ed1a, 32'h406a6631, 32'h424a2287, 32'h426c502a, 32'h426c6d57};
test_weights[18544:18551] = '{32'hc24bd0fc, 32'h428568c4, 32'hc2916fbd, 32'h3f9e0420, 32'h426c7cdb, 32'hc0eb076b, 32'h426e7808, 32'h4131dcad};
test_bias[2318:2318] = '{32'hc29fb47f};
test_output[2318:2318] = '{32'hc55d3b6c};
test_input[18552:18559] = '{32'h4288b647, 32'hc29feb06, 32'hc13e11db, 32'hc29cb5d7, 32'hc2247a32, 32'hc040fe1d, 32'h41df1547, 32'hc236fc66};
test_weights[18552:18559] = '{32'hbfdaca8b, 32'h421b8559, 32'hc2385842, 32'hc2627966, 32'h42950d9e, 32'h42aea55b, 32'h429df84a, 32'h42b3ee80};
test_bias[2319:2319] = '{32'h428a18c8};
test_output[2319:2319] = '{32'hc5555b05};
test_input[18560:18567] = '{32'h4190bc20, 32'hc2254264, 32'h42286a12, 32'h42af1bb6, 32'h420a2bd0, 32'h41fb2a7d, 32'h42825dd9, 32'hc2b5ccdc};
test_weights[18560:18567] = '{32'h41ce654d, 32'h4284b2cc, 32'h42a75d09, 32'h429274fd, 32'h419cfeca, 32'h42046411, 32'hc24086c8, 32'hc2b1a628};
test_bias[2320:2320] = '{32'hc24b3d6b};
test_output[2320:2320] = '{32'h465edd2a};
test_input[18568:18575] = '{32'hc2bb7216, 32'h423ff322, 32'hc1c9ef44, 32'h41d81114, 32'h42920440, 32'hc1e3f3af, 32'h4106ffa5, 32'hc209bef9};
test_weights[18568:18575] = '{32'h413ee3b0, 32'h421ff866, 32'hc2423b59, 32'h4234afae, 32'hc19d29cf, 32'hc298122c, 32'h427f46b1, 32'hc2b0244f};
test_bias[2321:2321] = '{32'hc2c0f3f5};
test_output[2321:2321] = '{32'h45e8ee5a};
test_input[18576:18583] = '{32'h42acc6e9, 32'h429eed81, 32'h423ebe35, 32'hc28a818d, 32'hc23c77a7, 32'hc2b7cdea, 32'h42b88c33, 32'h42210291};
test_weights[18576:18583] = '{32'h423c5282, 32'h428aafd4, 32'hc19d6bde, 32'hc1610e43, 32'h421fbdde, 32'hc1ddfef1, 32'h42a8abc8, 32'hc2b0f87d};
test_bias[2322:2322] = '{32'hc250a655};
test_output[2322:2322] = '{32'h4661c7ba};
test_input[18584:18591] = '{32'hc299e3e8, 32'hc18079ef, 32'h41d523d9, 32'hc2a62578, 32'hc2222c5a, 32'h422898bc, 32'h4118839b, 32'hc1ba9ff8};
test_weights[18584:18591] = '{32'h422650fa, 32'h41b1d0b1, 32'hc26f083c, 32'hc2b8d107, 32'h4181ce4a, 32'h42158c89, 32'h42ad7a1c, 32'hc1d1e46d};
test_bias[2323:2323] = '{32'hc221c610};
test_output[2323:2323] = '{32'h4597657e};
test_input[18592:18599] = '{32'h42c5b7a8, 32'h422fd4cd, 32'h411616e1, 32'h42957b9b, 32'hc2c1bcbf, 32'h41aed185, 32'h4207f17f, 32'hc21e852d};
test_weights[18592:18599] = '{32'hc0484782, 32'hc18c2006, 32'hc2bf7e1f, 32'h4114f6a3, 32'h41c4efbe, 32'hc105e299, 32'h4023924b, 32'h4002f18b};
test_bias[2324:2324] = '{32'hc2a57ca3};
test_output[2324:2324] = '{32'hc57560e0};
test_input[18600:18607] = '{32'hc2ab1ea5, 32'hc2b579a4, 32'hc2650dd2, 32'hc28b7777, 32'hc1afee71, 32'h42c53476, 32'hc2821ae9, 32'hc26d6c8a};
test_weights[18600:18607] = '{32'hc1fb8bee, 32'h428c8efe, 32'hc2beb82e, 32'h41a05fe8, 32'hc2baf13e, 32'hc1d70cde, 32'h4200fe49, 32'h41c532ea};
test_bias[2325:2325] = '{32'hc2bf294c};
test_output[2325:2325] = '{32'hc5723840};
test_input[18608:18615] = '{32'h42a42e6c, 32'h42044306, 32'hc189df66, 32'h421b229a, 32'h428d66d7, 32'hc2735d2f, 32'h42a1bdd1, 32'hc169c215};
test_weights[18608:18615] = '{32'h4267d154, 32'h428cb5ab, 32'hc133dbb8, 32'hc2850883, 32'h4205abb6, 32'h41149180, 32'h421832d0, 32'h40c292a4};
test_bias[2326:2326] = '{32'hc2b9a84e};
test_output[2326:2326] = '{32'h4612bbcf};
test_input[18616:18623] = '{32'hc242b61e, 32'h4293e51b, 32'h41174244, 32'hc2a170ed, 32'h42c30ade, 32'hc260a725, 32'hc214f553, 32'hc0174a50};
test_weights[18616:18623] = '{32'h42101a63, 32'hc2afa6d9, 32'h424aeda8, 32'hc1e39e04, 32'h40a44c63, 32'hc13132ce, 32'hc0b52cf1, 32'h421010f3};
test_bias[2327:2327] = '{32'h42400d09};
test_output[2327:2327] = '{32'hc5827bab};
test_input[18624:18631] = '{32'h4205cf67, 32'h42983ccc, 32'h42a3d0f8, 32'h4132e6eb, 32'h41659ae9, 32'h426c4cf4, 32'h427de714, 32'h425bdade};
test_weights[18624:18631] = '{32'h426f1924, 32'h422632eb, 32'hc1d77a9f, 32'h42aca884, 32'h42c4a788, 32'h42b9e31f, 32'hc122aaac, 32'hc187d715};
test_bias[2328:2328] = '{32'hc105823a};
test_output[2328:2328] = '{32'h4610508a};
test_input[18632:18639] = '{32'h42adac2c, 32'h420adc63, 32'hc29b0895, 32'hc15f864f, 32'h429437d2, 32'h427c8449, 32'hc2337412, 32'h42377efe};
test_weights[18632:18639] = '{32'hc2a54efa, 32'hc1f99c99, 32'h429e84d7, 32'hc29e78ec, 32'hc29ba528, 32'h4203ffb8, 32'hc2648fcd, 32'hc141889d};
test_bias[2329:2329] = '{32'h424d1d8d};
test_output[2329:2329] = '{32'hc66926f7};
test_input[18640:18647] = '{32'hc23dc62d, 32'hc28d7098, 32'hc210e84a, 32'hbe0c3ca2, 32'h4223bf3d, 32'h412dc200, 32'hc23778bd, 32'h4100c83c};
test_weights[18640:18647] = '{32'hc2bff736, 32'h41986117, 32'hc2ab30d2, 32'h416359ec, 32'h428764dc, 32'h4224ad54, 32'h428fc873, 32'h417c575f};
test_bias[2330:2330] = '{32'h428885f7};
test_output[2330:2330] = '{32'h45c8adb9};
test_input[18648:18655] = '{32'hc25f6b8f, 32'hbf87b23b, 32'hc25b8532, 32'h4263dd47, 32'hc244e309, 32'hc28d03da, 32'hc1f715ba, 32'h412d7a3a};
test_weights[18648:18655] = '{32'hc24e1f0c, 32'h3efd6a94, 32'hc2548bae, 32'hc25a3dea, 32'h42851520, 32'hc152e9d7, 32'hc2a5f75c, 32'h408b23db};
test_bias[2331:2331] = '{32'h426bc4d0};
test_output[2331:2331] = '{32'h453c0f7f};
test_input[18656:18663] = '{32'h429051b7, 32'hc15da462, 32'h42186766, 32'h42afb0a7, 32'h4253a06f, 32'hc2855d54, 32'h421cb819, 32'h4202f646};
test_weights[18656:18663] = '{32'h40ba9327, 32'h41f4b339, 32'hc140ac5a, 32'h42802683, 32'hc2bdc0e0, 32'hc2b7933e, 32'hc2237ca3, 32'h41bea124};
test_bias[2332:2332] = '{32'h4212d122};
test_output[2332:2332] = '{32'h45ab5b2e};
test_input[18664:18671] = '{32'hc2994e9b, 32'hc1f1c8af, 32'h427d69fe, 32'hc289184e, 32'hc2c506b1, 32'hc2bc53af, 32'h40d712ec, 32'hc2abef91};
test_weights[18664:18671] = '{32'h408887a3, 32'hc1b46619, 32'h42ad936a, 32'h42b46902, 32'h40f5116c, 32'hc2a87eb0, 32'h4284687d, 32'h42ac19d3};
test_bias[2333:2333] = '{32'h42b17fda};
test_output[2333:2333] = '{32'hc17d2270};
test_input[18672:18679] = '{32'hc2bf9dff, 32'h400025b5, 32'h42a7c39d, 32'h428ae919, 32'h429f2215, 32'hc263883c, 32'hc28feac4, 32'hc0cfeacb};
test_weights[18672:18679] = '{32'h42b4497b, 32'hc28da5e9, 32'hc2bdc5b0, 32'hc1bb9136, 32'h41ccc35b, 32'h421be8a6, 32'h424578f8, 32'h420c49fe};
test_bias[2334:2334] = '{32'h42ae71b3};
test_output[2334:2334] = '{32'hc6adbf79};
test_input[18680:18687] = '{32'h425d2958, 32'h4201ee3f, 32'h42aa8a2d, 32'h41e6dea9, 32'h411676ea, 32'hc195f612, 32'h424747f5, 32'h4299cfb5};
test_weights[18680:18687] = '{32'hc295a61c, 32'hc2c54135, 32'h421010aa, 32'h4217ce63, 32'hc2a7b657, 32'h427c9716, 32'hc2c0402f, 32'hc2b7bf82};
test_bias[2335:2335] = '{32'hc236dfc6};
test_output[2335:2335] = '{32'hc6852e1d};
test_input[18688:18695] = '{32'hc1d1f206, 32'hc28ae079, 32'h4240adb9, 32'h41c69183, 32'h429f3890, 32'h423cfd54, 32'h428cd135, 32'h427e09a1};
test_weights[18688:18695] = '{32'hc1b9dfdf, 32'hc2bf89ff, 32'hc29fc87e, 32'h42b12327, 32'hc29e1390, 32'h420237a1, 32'h414cf722, 32'h41c401e2};
test_bias[2336:2336] = '{32'hc0829bd2};
test_output[2336:2336] = '{32'h454ed98e};
test_input[18696:18703] = '{32'hc0ed4cc8, 32'hc2c22d3f, 32'h42aba95f, 32'h4206cac8, 32'h3fcdfd5c, 32'hc2b07364, 32'hc279398b, 32'hc2b30a61};
test_weights[18696:18703] = '{32'h418e846c, 32'hc07d5f9e, 32'h42888478, 32'hc2c4559f, 32'hc200314f, 32'hc2bdc605, 32'h4253b6c8, 32'h4297af95};
test_bias[2337:2337] = '{32'h41f07991};
test_output[2337:2337] = '{32'h44853255};
test_input[18704:18711] = '{32'hc29c7c8c, 32'h4269adff, 32'hc2408658, 32'h41f29d72, 32'hc28bb637, 32'h42222014, 32'h4179823f, 32'hc1110a46};
test_weights[18704:18711] = '{32'hc2abd3ba, 32'h41dcdcee, 32'hc2a010ac, 32'h426cc560, 32'h426462cc, 32'hc28fdf08, 32'h41a9a853, 32'hc0d68dbf};
test_bias[2338:2338] = '{32'h423c6715};
test_output[2338:2338] = '{32'h45eae4f2};
test_input[18712:18719] = '{32'h41e76ca4, 32'hc29f428c, 32'h42a03327, 32'hc28fddd0, 32'hc2a63418, 32'hc27c6839, 32'h421ea514, 32'h414e4edf};
test_weights[18712:18719] = '{32'hc202be25, 32'h40bd52db, 32'hc26fb8f4, 32'h418e1136, 32'hc1de2db1, 32'hc2c36b27, 32'hc251b166, 32'hc24ac8dc};
test_bias[2339:2339] = '{32'hc27ac3e1};
test_output[2339:2339] = '{32'hc4e31010};
test_input[18720:18727] = '{32'hc289bab1, 32'hc2aec2a0, 32'h41339bf2, 32'hc2449383, 32'h40af1cfe, 32'h4100bc17, 32'h4287c647, 32'hc2636513};
test_weights[18720:18727] = '{32'h42c7b4c3, 32'hc1442216, 32'h41867c62, 32'h42ad199c, 32'h42a92249, 32'hc1c67949, 32'hc19e97da, 32'hc29a9eb4};
test_bias[2340:2340] = '{32'h427875d6};
test_output[2340:2340] = '{32'hc5cafbd1};
test_input[18728:18735] = '{32'h424f2035, 32'hc1952087, 32'h428088dd, 32'h42c253cc, 32'h404a3534, 32'h41f42cba, 32'h41001256, 32'h4226b107};
test_weights[18728:18735] = '{32'h42927760, 32'h421870a8, 32'h42a6eccd, 32'hc2a5a5b2, 32'hc240b36b, 32'h42c05d81, 32'hc21281bf, 32'h4272bc11};
test_bias[2341:2341] = '{32'h42c07820};
test_output[2341:2341] = '{32'h45ac4c7b};
test_input[18736:18743] = '{32'h4203192e, 32'hc2a08360, 32'hc1cc01c6, 32'h40fd196e, 32'hc2b6abc3, 32'h3f483055, 32'h424ca029, 32'h41d481db};
test_weights[18736:18743] = '{32'hc119fe8d, 32'hc2779533, 32'h41d24483, 32'h41b1d43b, 32'hc29a1829, 32'h42afa577, 32'h4273cc84, 32'hc2b66cd5};
test_bias[2342:2342] = '{32'hc249e40f};
test_output[2342:2342] = '{32'h463a1038};
test_input[18744:18751] = '{32'h4257a9c9, 32'h41f23ee9, 32'h42c3778f, 32'hc2958ccc, 32'h42648dfa, 32'h42a5db8d, 32'h42bd2945, 32'hc2a2c836};
test_weights[18744:18751] = '{32'h42c35a3f, 32'h4139038d, 32'h42847909, 32'hc24cbabb, 32'hc1b2c910, 32'h419b5f35, 32'h41c76341, 32'h4149acfa};
test_bias[2343:2343] = '{32'hc21db267};
test_output[2343:2343] = '{32'h46890d6d};
test_input[18752:18759] = '{32'h40bc7a6f, 32'hc291e54e, 32'h4285e86c, 32'h41a5d894, 32'hc2abcbcc, 32'h407c61e7, 32'hc1aebe15, 32'hc2928eca};
test_weights[18752:18759] = '{32'hc1e0c94f, 32'hc296d6fc, 32'hc297e09f, 32'h40a6208a, 32'h424bdc08, 32'h428e59f4, 32'hc20e6c8a, 32'h4254f170};
test_bias[2344:2344] = '{32'h42608576};
test_output[2344:2344] = '{32'hc5d4a6c7};
test_input[18760:18767] = '{32'h414473b9, 32'hc291c355, 32'hc21632b1, 32'h422d3c35, 32'hc28811d8, 32'hc2b04e18, 32'h42a6fe01, 32'h429d4ded};
test_weights[18760:18767] = '{32'hc1911416, 32'hc2c34e2d, 32'h42451e67, 32'h42b42cbf, 32'h4281c316, 32'hc20c4897, 32'hc14b1de9, 32'hc2b7a058};
test_bias[2345:2345] = '{32'hc19ab9ce};
test_output[2345:2345] = '{32'hc42968f6};
test_input[18768:18775] = '{32'h4200d5a6, 32'hc27490e9, 32'h41950d39, 32'hc2c27b7d, 32'hc1a736b1, 32'h427f7282, 32'hc21874b0, 32'h427b3f75};
test_weights[18768:18775] = '{32'hc2a2b947, 32'hbfaff58e, 32'hc2055469, 32'hc1a60d89, 32'h42b0e310, 32'hc28eb5f9, 32'h42850c93, 32'hc1ded774};
test_bias[2346:2346] = '{32'h42a5c046};
test_output[2346:2346] = '{32'hc6378bb3};
test_input[18776:18783] = '{32'h40982828, 32'h4192f9cc, 32'h41e73f2b, 32'h4206173a, 32'h4267dad2, 32'h423b82ba, 32'hc1eecdda, 32'hc27b5138};
test_weights[18776:18783] = '{32'hc2c4b137, 32'hc2725246, 32'h4284f47a, 32'h42729586, 32'hbb8288c7, 32'hc229c7ff, 32'h3f671cf5, 32'hc2b3946d};
test_bias[2347:2347] = '{32'hc09a5b4e};
test_output[2347:2347] = '{32'h45bb4d92};
test_input[18784:18791] = '{32'hc231059b, 32'hc258a32f, 32'h428a7736, 32'h42970550, 32'h4136970e, 32'hc2604ccb, 32'hc296c6e6, 32'h42b66c08};
test_weights[18784:18791] = '{32'hc13ff3a4, 32'h420873d4, 32'hc2bc5460, 32'h40e8c4fe, 32'hc299266b, 32'hc2c56fa4, 32'hc1b00864, 32'h429c129a};
test_bias[2348:2348] = '{32'h422ac5cc};
test_output[2348:2348] = '{32'h45c1936b};
test_input[18792:18799] = '{32'hc28a4dbb, 32'hc1d1520a, 32'h3ff56574, 32'h3fd58332, 32'h42b39093, 32'hc2c74add, 32'hc27aaa62, 32'hc236ee71};
test_weights[18792:18799] = '{32'h428de41e, 32'hc1eb81ed, 32'h42967b76, 32'h41c33c24, 32'h4163c7b6, 32'hc2848178, 32'hc2ac844f, 32'h42257cef};
test_bias[2349:2349] = '{32'hc116ced4};
test_output[2349:2349] = '{32'h45e849dd};
test_input[18800:18807] = '{32'hc2785e0a, 32'h41f9eaf9, 32'h42aecd1d, 32'hc1730a6a, 32'hc22cc2e3, 32'hc159a1ee, 32'hc24b26dc, 32'hc2428505};
test_weights[18800:18807] = '{32'h429e76d1, 32'hc2170e0e, 32'h42531239, 32'hc170d661, 32'hc20e1ac0, 32'h4275a710, 32'hc1d5c688, 32'h41abc62c};
test_bias[2350:2350] = '{32'h40b2aca3};
test_output[2350:2350] = '{32'hc37133d0};
test_input[18808:18815] = '{32'hc290168a, 32'hc21b9612, 32'h42421918, 32'hc2c6bbec, 32'h42bbcdb6, 32'hc128b7ce, 32'h422b23f9, 32'hc29f29de};
test_weights[18808:18815] = '{32'hc20a6bca, 32'hc21ee63a, 32'h4251ce7b, 32'h4194855b, 32'hc208063d, 32'hc1fbaa3c, 32'hc1e6fad1, 32'hc20bd94c};
test_bias[2351:2351] = '{32'h424e7fd8};
test_output[2351:2351] = '{32'h45593d8d};
test_input[18816:18823] = '{32'h42155547, 32'hc2bf2f00, 32'h3fa4a4a0, 32'hc1f40cbf, 32'h42c3baaf, 32'h425521cb, 32'hc2b26796, 32'h40f82d55};
test_weights[18816:18823] = '{32'h42a9e18e, 32'hc2a0d09e, 32'h42b43312, 32'h41773279, 32'hc1b452f0, 32'hc23abbbb, 32'h423e2a49, 32'hc1a6993e};
test_bias[2352:2352] = '{32'h42a6d8af};
test_output[2352:2352] = '{32'h44ba3830};
test_input[18824:18831] = '{32'h4284041c, 32'hc154b402, 32'h42a0102c, 32'hc1041139, 32'hc2794549, 32'h41a55674, 32'hc0e486f5, 32'h429f2e36};
test_weights[18824:18831] = '{32'h3ec6c4df, 32'h415febf2, 32'hc2c02607, 32'hc2a52a6a, 32'hc2ba254d, 32'h42263143, 32'hc2a32314, 32'hc2773eb1};
test_bias[2353:2353] = '{32'h426075c7};
test_output[2353:2353] = '{32'hc595af53};
test_input[18832:18839] = '{32'hc2749334, 32'h421c1c9d, 32'h41809f58, 32'h42c7f15f, 32'h4270ce6e, 32'hc112c457, 32'h41567177, 32'hc2902855};
test_weights[18832:18839] = '{32'hc184ac14, 32'h419c8d5a, 32'hc21d3073, 32'hbfac21e9, 32'hc2c4f971, 32'hc29bbfbb, 32'hc1de8456, 32'hc137d5af};
test_bias[2354:2354] = '{32'hc1d9fea2};
test_output[2354:2354] = '{32'hc56bf225};
test_input[18840:18847] = '{32'hc2b69515, 32'h42ada423, 32'h42428c19, 32'hc1bca38d, 32'h428d915a, 32'h412ad7cc, 32'h42a6b5c9, 32'h41fe7c11};
test_weights[18840:18847] = '{32'hc2408f7c, 32'h422ac931, 32'h429db2f7, 32'h40da4609, 32'h40d4bd31, 32'h4286e42e, 32'h42b68046, 32'hc08cb847};
test_bias[2355:2355] = '{32'h41fad574};
test_output[2355:2355] = '{32'h469fe082};
test_input[18848:18855] = '{32'hc2b8ae78, 32'h4274afbb, 32'h41da8fdd, 32'h417a9741, 32'h42082d05, 32'h4269930e, 32'hc2058269, 32'h421da829};
test_weights[18848:18855] = '{32'hc1906996, 32'hc1ef897d, 32'h42c10ae8, 32'hc08b22e5, 32'h42106f35, 32'h42b5da0d, 32'h426c339f, 32'hc2863487};
test_bias[2356:2356] = '{32'hc15ee01b};
test_output[2356:2356] = '{32'h4586ca2c};
test_input[18856:18863] = '{32'h42952597, 32'h427bb21f, 32'hc09acead, 32'hc28ce43c, 32'hc25c3454, 32'hc2a075b6, 32'hc2becf42, 32'hc21a221f};
test_weights[18856:18863] = '{32'h4287ed1a, 32'hc27e4974, 32'hc2af94b1, 32'h42180c70, 32'h41cd26c6, 32'h42625232, 32'hc2714ba0, 32'h410d7bc4};
test_bias[2357:2357] = '{32'hc28da9b5};
test_output[2357:2357] = '{32'hc4e01267};
test_input[18864:18871] = '{32'hc2913bb7, 32'h42c03005, 32'h4121dab8, 32'hc2b2cf41, 32'hc185bffb, 32'h421cb355, 32'hc1389125, 32'hc208d991};
test_weights[18864:18871] = '{32'hc1c8c489, 32'h4213f318, 32'hc27b637a, 32'hc2691166, 32'hc2a493f9, 32'h41407799, 32'h4293d538, 32'hc1b5252f};
test_bias[2358:2358] = '{32'hc11f2d60};
test_output[2358:2358] = '{32'h4636f549};
test_input[18872:18879] = '{32'hc20b2ac9, 32'hc1f06058, 32'hc2a4cae9, 32'h42aa9101, 32'h3e93be67, 32'hc05bc15b, 32'hc24984e9, 32'hc26838c8};
test_weights[18872:18879] = '{32'hc285750b, 32'hc28c6c6a, 32'hc1ac8931, 32'hc15d79d1, 32'hc28a1f1e, 32'hc2bd142f, 32'hc289b843, 32'hc2b77ae5};
test_bias[2359:2359] = '{32'h42c2811d};
test_output[2359:2359] = '{32'h465e438f};
test_input[18880:18887] = '{32'hc1d16204, 32'hc278b28e, 32'h422dc710, 32'hc284a579, 32'hc288b110, 32'hc0f2827c, 32'hc2833232, 32'h42b92591};
test_weights[18880:18887] = '{32'hbfcd9438, 32'h41e3c6fb, 32'h42a40ca1, 32'h41a17841, 32'hc20e6ced, 32'h42c0f6ef, 32'h42c48b4f, 32'h411e20c0};
test_bias[2360:2360] = '{32'h42ad11ca};
test_output[2360:2360] = '{32'hc54adfed};
test_input[18888:18895] = '{32'h4118f0b0, 32'h42a48d11, 32'hc2b95d39, 32'hc2062745, 32'hc296d204, 32'h41462d1d, 32'h4210f56c, 32'h429e024d};
test_weights[18888:18895] = '{32'h428bd57b, 32'hc2c18b7e, 32'h428c2516, 32'hc1a4b8f5, 32'h42159da7, 32'h429cf4ca, 32'hc0328887, 32'h41ea6a19};
test_bias[2361:2361] = '{32'h424941d5};
test_output[2361:2361] = '{32'hc64627f7};
test_input[18896:18903] = '{32'hc2727ae0, 32'hc1c2d97d, 32'h4177a603, 32'h41d38492, 32'h42bbab72, 32'h40dd3f37, 32'hc25aa832, 32'h41194da3};
test_weights[18896:18903] = '{32'h42b0f57c, 32'h4171539b, 32'h422376a6, 32'hc2407521, 32'h42a100a0, 32'hc1882a35, 32'hc221c54a, 32'hc205de0e};
test_bias[2362:2362] = '{32'hc1b0d59f};
test_output[2362:2362] = '{32'h453758c3};
test_input[18904:18911] = '{32'hc20b93ff, 32'h42c6c54c, 32'h415e0bc8, 32'hc1c28804, 32'h42916ad7, 32'h42271f98, 32'h4240c31a, 32'h41cd5f16};
test_weights[18904:18911] = '{32'h4264a957, 32'hc2c5be20, 32'hc1ac84fc, 32'h42747d51, 32'hc198082a, 32'hc1cf1a09, 32'hc1cb7193, 32'hc2c14ff5};
test_bias[2363:2363] = '{32'hc23a064c};
test_output[2363:2363] = '{32'hc69adeb5};
test_input[18912:18919] = '{32'hc2020a3a, 32'hc284ea79, 32'h423e4da7, 32'h4282966d, 32'h42946670, 32'h41aecb14, 32'hc22b844f, 32'hc28ea400};
test_weights[18912:18919] = '{32'h40ab290d, 32'h4211d09a, 32'h41cbd576, 32'h42016d87, 32'hc1cd4e99, 32'h41a011ba, 32'hc2b45f25, 32'h4204ee93};
test_bias[2364:2364] = '{32'hc16c9a65};
test_output[2364:2364] = '{32'h4439dc9f};
test_input[18920:18927] = '{32'hc26b24f4, 32'h41de91ce, 32'h41f06ceb, 32'hc2979c0c, 32'h3f762afc, 32'h429b49d3, 32'h42b9d6dc, 32'hc20c02bb};
test_weights[18920:18927] = '{32'h429db772, 32'h428e47a7, 32'hc2a947cd, 32'h4238b8f3, 32'hc015eb55, 32'hc2ac76d6, 32'hc0ba7c3c, 32'h41478501};
test_bias[2365:2365] = '{32'hc09ebc62};
test_output[2365:2365] = '{32'hc67ff674};
test_input[18928:18935] = '{32'hc2c4a4a0, 32'h421cdb55, 32'h42902b88, 32'hc115b119, 32'h41ad4679, 32'h41f9a359, 32'h42878b05, 32'h42475c63};
test_weights[18928:18935] = '{32'hc25c6705, 32'h3feb8761, 32'h4285e4a0, 32'hc1cf48c2, 32'h41ed99c5, 32'hc1e7637f, 32'hc23a8a53, 32'hbf3d6dd2};
test_bias[2366:2366] = '{32'h42854195};
test_output[2366:2366] = '{32'h45dfff82};
test_input[18936:18943] = '{32'h41fc5434, 32'hc2c17a20, 32'h429565e7, 32'hc1f13379, 32'hc216dd44, 32'h42bc2b28, 32'hc16a0189, 32'hc2940082};
test_weights[18936:18943] = '{32'hc209a904, 32'h4149e158, 32'hc2938e30, 32'h42b4a69b, 32'hc2a56ea7, 32'h42bbb1e2, 32'h4285b97d, 32'hc12f317a};
test_bias[2367:2367] = '{32'hc1ed7e5b};
test_output[2367:2367] = '{32'h44976ef5};
test_input[18944:18951] = '{32'hc12799cf, 32'h4157ac20, 32'h423be753, 32'h4108afca, 32'h425fc12d, 32'h41d5e3a5, 32'h411f7a4a, 32'h42ab6c2e};
test_weights[18944:18951] = '{32'hc0985357, 32'hc29ff174, 32'h428805bb, 32'h42bc4e0b, 32'h4291f455, 32'h4135bd3a, 32'h40b85615, 32'h4122651b};
test_bias[2368:2368] = '{32'h42b5cab0};
test_output[2368:2368] = '{32'h4602dd31};
test_input[18952:18959] = '{32'h42a39193, 32'h423b678c, 32'h41b63175, 32'h42b089d2, 32'hc2bfd429, 32'hc1e3f720, 32'h4045acb3, 32'h41c5b2b6};
test_weights[18952:18959] = '{32'h42297195, 32'hc2708021, 32'h42a20a27, 32'h42445016, 32'hc29563a1, 32'hbe2ea96b, 32'h423708fe, 32'h42a357f6};
test_bias[2369:2369] = '{32'h412c9d65};
test_output[2369:2369] = '{32'h467c915f};
test_input[18960:18967] = '{32'h4255f2a5, 32'h422924ce, 32'hc2315433, 32'hc1ab4585, 32'hc24e361f, 32'hc1ff664d, 32'hc20652b0, 32'hc2bc6902};
test_weights[18960:18967] = '{32'h422b7532, 32'hc28ee38d, 32'hc2873a22, 32'hc2badbd7, 32'h42af10c7, 32'hc24bef48, 32'hc29c04d6, 32'h42a97e73};
test_bias[2370:2370] = '{32'hc1e9d099};
test_output[2370:2370] = '{32'hc57a8d7f};
test_input[18968:18975] = '{32'hc282c3bf, 32'h42c3a508, 32'h427c7309, 32'h42a4d898, 32'hc0d0c302, 32'hc1078731, 32'hc1d1e6ad, 32'hc2862e8f};
test_weights[18968:18975] = '{32'h41966205, 32'h42b094f3, 32'h42a71276, 32'hc24c0a61, 32'h420e0537, 32'hc269f4ae, 32'h42a6986a, 32'hc29f644a};
test_bias[2371:2371] = '{32'hc2ba382d};
test_output[2371:2371] = '{32'h46387e34};
test_input[18976:18983] = '{32'h412fbd8a, 32'hc210895e, 32'h42930070, 32'hc268c39b, 32'h42c5aeba, 32'hc274356f, 32'hc26bbd99, 32'h42b2d358};
test_weights[18976:18983] = '{32'hc2b25c06, 32'hc2a47c22, 32'h425f4b45, 32'h424d2c8c, 32'h40697e1e, 32'h4214a9d7, 32'h42439864, 32'h4212eb06};
test_bias[2372:2372] = '{32'hc22836d8};
test_output[2372:2372] = '{32'h44c346a6};
test_input[18984:18991] = '{32'hc286ec47, 32'hc1c1e06b, 32'hc25f207b, 32'hc2950e9b, 32'h4297032b, 32'h41febb6b, 32'h42ba26f5, 32'hc22fd86d};
test_weights[18984:18991] = '{32'h41a06903, 32'h41a3c3cc, 32'h423eecf5, 32'hc29feec4, 32'h4290ce20, 32'hc2580de8, 32'hc040ae7b, 32'h42a26a49};
test_bias[2373:2373] = '{32'h40482652};
test_output[2373:2373] = '{32'h44a88a91};
test_input[18992:18999] = '{32'hc28e730d, 32'hc0e98c41, 32'h42a495e7, 32'h425d8783, 32'h42429915, 32'h42bb97f5, 32'h3e58d36f, 32'hc20bb30d};
test_weights[18992:18999] = '{32'h42aa4627, 32'hc1463c52, 32'h4263047d, 32'hc297d2b2, 32'hc203abfc, 32'hc2bba825, 32'hc2801264, 32'h419adac4};
test_bias[2374:2374] = '{32'hc2959f9b};
test_output[2374:2374] = '{32'hc6824388};
test_input[19000:19007] = '{32'hc2a5c1e9, 32'hc074ab66, 32'hc2af2657, 32'hc29b2007, 32'h4297694a, 32'h428d651c, 32'hc1c49655, 32'hc28b6b36};
test_weights[19000:19007] = '{32'hc245e9b2, 32'h424008db, 32'hc1d3810a, 32'hc2855abc, 32'hc1e62ee3, 32'hc273b71b, 32'hc1fca65d, 32'hc202b93b};
test_bias[2375:2375] = '{32'hc245bdf1};
test_output[2375:2375] = '{32'h45f798f8};
test_input[19008:19015] = '{32'hc2b65fa5, 32'hc2bf539e, 32'h42b57297, 32'h4293a7f9, 32'h3ff88f03, 32'hc2490346, 32'h422dc782, 32'h3ffb2768};
test_weights[19008:19015] = '{32'hc296bce1, 32'hc22d12df, 32'h42c32ba9, 32'hc29cd9cc, 32'hbf290553, 32'hc2447c42, 32'hc23c6f9d, 32'h42ae70fd};
test_bias[2376:2376] = '{32'hc27b4d8a};
test_output[2376:2376] = '{32'h4664303b};
test_input[19016:19023] = '{32'h42973390, 32'h42aa934c, 32'hc2437ef0, 32'hc1a370bb, 32'h41b05bbc, 32'hc2ae8ee2, 32'hc24fbc2c, 32'h4289a08d};
test_weights[19016:19023] = '{32'hc28931d5, 32'h42c3bae9, 32'hc26a5e0a, 32'h42b5ac98, 32'h4287bda4, 32'h42571ae8, 32'hc258f022, 32'h42a1daaa};
test_bias[2377:2377] = '{32'hc2c3a5ae};
test_output[2377:2377] = '{32'h4610ab2c};
test_input[19024:19031] = '{32'h4223330f, 32'h4264d8d3, 32'h420a47c4, 32'hc205edc2, 32'h42728bfa, 32'hc264d77f, 32'hc20a98e9, 32'h409630a1};
test_weights[19024:19031] = '{32'h41cd6dc1, 32'h419670ba, 32'hc1c64c93, 32'h41e308f9, 32'hc25cb5f1, 32'hc2a0ac8c, 32'h42b74d40, 32'h42533093};
test_bias[2378:2378] = '{32'h420654ba};
test_output[2378:2378] = '{32'hc4a5ef95};
test_input[19032:19039] = '{32'hc26a3ba4, 32'hc23276e5, 32'hc223b806, 32'h40f2325f, 32'h42c5df44, 32'hc2912536, 32'hc2809ad0, 32'hc2bcc9cc};
test_weights[19032:19039] = '{32'h423e4bc2, 32'hc1190d01, 32'hc1d36b8d, 32'h41eb27f5, 32'h42ab657b, 32'hc26d766a, 32'hc1c2e1f1, 32'h424a8e5c};
test_bias[2379:2379] = '{32'hc2acd064};
test_output[2379:2379] = '{32'h4603c029};
test_input[19040:19047] = '{32'hc1c867cb, 32'h42c2859e, 32'hc21cef0e, 32'h40cd5d33, 32'h42a58553, 32'hc28107ba, 32'hc2b7f1e1, 32'hc2314ec1};
test_weights[19040:19047] = '{32'hc27a2278, 32'h42a3b712, 32'h413ffb7b, 32'hc214a17e, 32'h42bda580, 32'h42295112, 32'hc1afd433, 32'h42211704};
test_bias[2380:2380] = '{32'h42928b12};
test_output[2380:2380] = '{32'h465e9477};
test_input[19048:19055] = '{32'hc27b51ec, 32'h428356ce, 32'hc2b5b5bf, 32'h421d5f22, 32'h3fe0e3c4, 32'h42887462, 32'h41f39564, 32'h4272e4b8};
test_weights[19048:19055] = '{32'hc2a70237, 32'hc1d9c4c9, 32'hc289878c, 32'h42240b23, 32'h41ca67e6, 32'hc2378448, 32'hc2106bfe, 32'hc1b9961b};
test_bias[2381:2381] = '{32'h42a58e51};
test_output[2381:2381] = '{32'h45b588b3};
test_input[19056:19063] = '{32'hc2398797, 32'hc0b34239, 32'h425385f2, 32'h40b6e9c9, 32'hc173b5ef, 32'hbfe18c8a, 32'h4295a7cc, 32'h409d2276};
test_weights[19056:19063] = '{32'hc2ac345c, 32'hc0f14125, 32'hc24f85c0, 32'hc298666f, 32'h424f188f, 32'h41ca0c3a, 32'hc27ef4f9, 32'hc21035b4};
test_bias[2382:2382] = '{32'hc2a0de16};
test_output[2382:2382] = '{32'hc59c59e6};
test_input[19064:19071] = '{32'h424ba43b, 32'hc297d578, 32'h41bef535, 32'h42468901, 32'h428ed296, 32'h425fe988, 32'h42aee725, 32'hc24418d9};
test_weights[19064:19071] = '{32'hc2b233d5, 32'h42a47de3, 32'hc1463430, 32'h42a4fd6e, 32'hc2ac69d5, 32'h419047b5, 32'hc2c24cec, 32'hc1ea82ae};
test_bias[2383:2383] = '{32'hc2884185};
test_output[2383:2383] = '{32'hc6966d72};
test_input[19072:19079] = '{32'hc1d53a64, 32'hc1adb275, 32'hc2678dd8, 32'h4280cdc7, 32'h4278cfce, 32'h423a26dc, 32'h42c26f8c, 32'h4202cee4};
test_weights[19072:19079] = '{32'h426b68fd, 32'h42a7fb2c, 32'h40b45ea2, 32'hc10c584c, 32'hc144c433, 32'hc2a1b996, 32'hc0d4005f, 32'h429e7a21};
test_bias[2384:2384] = '{32'h41d6683c};
test_output[2384:2384] = '{32'hc5d5acb2};
test_input[19080:19087] = '{32'hc296d404, 32'h42b8bc59, 32'h41621a88, 32'h42009129, 32'h4205160a, 32'h40996177, 32'hc2c066b4, 32'h425e8163};
test_weights[19080:19087] = '{32'h412635f6, 32'h42682ed3, 32'h42a5cf32, 32'h429565bb, 32'h422c155c, 32'h409e99e8, 32'hc2b28660, 32'h4293d180};
test_bias[2385:2385] = '{32'h42b368f2};
test_output[2385:2385] = '{32'h46aef3c6};
test_input[19088:19095] = '{32'h42a67818, 32'h42b6503e, 32'h42b12caa, 32'h4266c73e, 32'h42be9aa3, 32'h41329c12, 32'hc210fd2e, 32'hc173c951};
test_weights[19088:19095] = '{32'hc1f4b69c, 32'h419ce04f, 32'hc20ba19d, 32'h427a111c, 32'hc1bd441e, 32'h422c6688, 32'hc2c5a6f9, 32'hc2be8f46};
test_bias[2386:2386] = '{32'hc14d8e0a};
test_output[2386:2386] = '{32'h453bb79c};
test_input[19096:19103] = '{32'hc248e633, 32'hc08c48c1, 32'hc1dbeda5, 32'h41a4f270, 32'hc27efe95, 32'hc28048a0, 32'h421c0ede, 32'h41cd8773};
test_weights[19096:19103] = '{32'hc2bb620b, 32'h42a49d7c, 32'hc2b53cfe, 32'h429407a2, 32'h42549f1f, 32'h42430124, 32'h42c0b400, 32'hc25d6855};
test_bias[2387:2387] = '{32'hc28d24b6};
test_output[2387:2387] = '{32'h4580880f};
test_input[19104:19111] = '{32'h42ae442c, 32'h424cf558, 32'h423c881d, 32'hc08871cc, 32'hc247c81b, 32'h42833d63, 32'hc151e0ca, 32'hc298c6b0};
test_weights[19104:19111] = '{32'hc20cabd2, 32'h414d410e, 32'hc01243cb, 32'hc2b0bede, 32'hc26d14f2, 32'h4286d3b0, 32'h41dc9429, 32'hc26576ea};
test_bias[2388:2388] = '{32'h42bb3e15};
test_output[2388:2388] = '{32'h46124079};
test_input[19112:19119] = '{32'hc122c880, 32'hc21afa8a, 32'hc2a04777, 32'h421b5f62, 32'hc2a84102, 32'h42b71edf, 32'h4102d226, 32'hc2c0ad25};
test_weights[19112:19119] = '{32'hc1986bc5, 32'h42a475d8, 32'h417f6b9a, 32'h42205e02, 32'hc21fdc33, 32'h429b0c3a, 32'hc2b7d661, 32'h42060562};
test_bias[2389:2389] = '{32'h42428989};
test_output[2389:2389] = '{32'h456e7500};
test_input[19120:19127] = '{32'hc1181183, 32'h4199074b, 32'hc2ada850, 32'h42a8311a, 32'hc0b3eda0, 32'hc220b5e3, 32'h42c4032b, 32'h420f4d56};
test_weights[19120:19127] = '{32'h41b30871, 32'h42bb2fc2, 32'h42805864, 32'hc2b0b3f9, 32'h42b0cb6c, 32'hc29467e7, 32'hc267a900, 32'hc2623b24};
test_bias[2390:2390] = '{32'h4279bcdc};
test_output[2390:2390] = '{32'hc68187f0};
test_input[19128:19135] = '{32'h42c1ba3f, 32'h4295ec80, 32'hc10315a4, 32'hc260b243, 32'h42806f85, 32'h429c0580, 32'hc1c89897, 32'hc26674a5};
test_weights[19128:19135] = '{32'h428e9234, 32'hc22e2cf5, 32'h423c3a11, 32'h41b75cb2, 32'h42ab8d79, 32'hc2990a1e, 32'h42bc022c, 32'h42473479};
test_bias[2391:2391] = '{32'h4290ac43};
test_output[2391:2391] = '{32'hc563f361};
test_input[19136:19143] = '{32'hc2b06093, 32'hc19c7a9f, 32'hc2a7a47d, 32'hc1f27b24, 32'h3f31e909, 32'hc10dbe9f, 32'h42a84d8c, 32'h42075d00};
test_weights[19136:19143] = '{32'h4192100b, 32'hc1e9660f, 32'h4090fedf, 32'hc250ece9, 32'h41173523, 32'h42bd75a0, 32'h42adae87, 32'hc24d63b2};
test_bias[2392:2392] = '{32'h42566332};
test_output[2392:2392] = '{32'h459ad7a9};
test_input[19144:19151] = '{32'hc2263874, 32'hc2348deb, 32'hc2585ca5, 32'h42af8a5c, 32'hc1289a73, 32'h419dfad2, 32'hc1b3a28a, 32'h426c616c};
test_weights[19144:19151] = '{32'hc20a03c7, 32'hc13601ca, 32'h419261fc, 32'hc2b1af8f, 32'h42ae6b74, 32'hc2bb1283, 32'hc2a3b37c, 32'h4188507e};
test_bias[2393:2393] = '{32'hc1ee7291};
test_output[2393:2393] = '{32'hc5d43a42};
test_input[19152:19159] = '{32'h42902ec0, 32'hc27ae72a, 32'hc15220d3, 32'hc29b8291, 32'hbd1689e5, 32'hc2a91f17, 32'h42689cd5, 32'h4230c560};
test_weights[19152:19159] = '{32'h42220408, 32'hc14903b7, 32'h41a701b6, 32'h42a505c0, 32'h3f31e1f0, 32'hc1eccebb, 32'h415dbe57, 32'hc17732e2};
test_bias[2394:2394] = '{32'hc1761166};
test_output[2394:2394] = '{32'hc3b979fa};
test_input[19160:19167] = '{32'hc18a58be, 32'hc0bbbea0, 32'hc242e5c4, 32'h41888661, 32'h42b0832b, 32'hc285800d, 32'hc294bb55, 32'h429cba30};
test_weights[19160:19167] = '{32'h414663ab, 32'hc18c121f, 32'h42a1f464, 32'h4286cbc2, 32'h421e79ce, 32'hc1813e61, 32'hc216b2eb, 32'h42022d23};
test_bias[2395:2395] = '{32'h40ddef6a};
test_output[2395:2395] = '{32'h45db96ae};
test_input[19168:19175] = '{32'h42b5025c, 32'h420fe0db, 32'hc1cea3d3, 32'h423d0db9, 32'hc25de299, 32'hb9c4679c, 32'h3fea027b, 32'h428a019e};
test_weights[19168:19175] = '{32'h41f41480, 32'hc295e317, 32'h42b4df67, 32'hc274bc5d, 32'h40b1a035, 32'h42b3647a, 32'h426cd4de, 32'h4298603a};
test_bias[2396:2396] = '{32'hc2603457};
test_output[2396:2396] = '{32'hc320aa30};
test_input[19176:19183] = '{32'h42450a73, 32'h42b180e5, 32'hc21a4e97, 32'h42c4c3fc, 32'h42bb39e3, 32'hc270027e, 32'hc211bc5d, 32'h412baded};
test_weights[19176:19183] = '{32'h42a67939, 32'h40e5f2ef, 32'hc2ab8070, 32'hc1c58f5c, 32'hc25d15f7, 32'hc2b89f7e, 32'h42603db4, 32'h41e0a34d};
test_bias[2397:2397] = '{32'hc1796b06};
test_output[2397:2397] = '{32'h4584038c};
test_input[19184:19191] = '{32'hc209ea8c, 32'hc1c44887, 32'hc28fed73, 32'hc24b2402, 32'h42998bb5, 32'h42abbfcb, 32'h42ae3a6e, 32'h42808b07};
test_weights[19184:19191] = '{32'hc2b2677a, 32'h42b89f0b, 32'hc1b3657e, 32'h42182613, 32'h42a2d5cb, 32'h42896e11, 32'h4293c818, 32'h41d4b729};
test_bias[2398:2398] = '{32'h428e19dd};
test_output[2398:2398] = '{32'h46a2fa6d};
test_input[19192:19199] = '{32'h426e4b1e, 32'h42b787f1, 32'h42816353, 32'hc271a81a, 32'hc2bbfa8d, 32'hbf9f0b1a, 32'h41ba89fc, 32'h42b8e21d};
test_weights[19192:19199] = '{32'h42a8247e, 32'hc2a4f719, 32'h4268d865, 32'h429919c1, 32'h415affc1, 32'h41fda98c, 32'hc2c5e5d8, 32'h4201f88a};
test_bias[2399:2399] = '{32'hc0dd81bb};
test_output[2399:2399] = '{32'hc57d7cb1};
test_input[19200:19207] = '{32'h41c439b8, 32'hbfe2e0f4, 32'h425b543b, 32'hc213fd15, 32'hc1639b6c, 32'hc28f9df4, 32'hbf840dfd, 32'hc0856c77};
test_weights[19200:19207] = '{32'h41bd7250, 32'h42be3d55, 32'h40d83650, 32'h41cc7116, 32'hc2684517, 32'h42a9c3ce, 32'h42af9ea8, 32'h42c4d1ca};
test_bias[2400:2400] = '{32'h4127a065};
test_output[2400:2400] = '{32'hc5b91359};
test_input[19208:19215] = '{32'hc29c87c8, 32'hc1bedea2, 32'h429c5945, 32'hc284cc77, 32'hc214033b, 32'h42496623, 32'h42004a22, 32'h4117d6df};
test_weights[19208:19215] = '{32'hc2abfa8e, 32'h4203f639, 32'h40e6336f, 32'h429eab77, 32'hc17e6946, 32'hc17332ef, 32'h41739b82, 32'h42ba547c};
test_bias[2401:2401] = '{32'h4286e328};
test_output[2401:2401] = '{32'h451c467d};
test_input[19216:19223] = '{32'h414cf61f, 32'h42a2a183, 32'h42b56970, 32'h42735353, 32'hc2b21c02, 32'h429e3d20, 32'hbf4ddf21, 32'h40d83796};
test_weights[19216:19223] = '{32'h426f04f9, 32'hc2991fcb, 32'hc294651c, 32'h41878e49, 32'h4226bd82, 32'hc0a8d01a, 32'h421d2e2b, 32'h429514b5};
test_bias[2402:2402] = '{32'hc2a8f8d2};
test_output[2402:2402] = '{32'hc668d6bb};
test_input[19224:19231] = '{32'h3fe91f9e, 32'hbef3d96c, 32'hc209ce1f, 32'h42c30ef1, 32'h429c2a9e, 32'hc2be1f80, 32'h4287c6c9, 32'hc1a1591f};
test_weights[19224:19231] = '{32'hc26886f5, 32'hc1d25980, 32'h42b04a23, 32'hc24b625e, 32'h42c3a170, 32'hc14cb14c, 32'hc1c5019d, 32'hc2822b4d};
test_bias[2403:2403] = '{32'h42a456a5};
test_output[2403:2403] = '{32'h43f3f11f};
test_input[19232:19239] = '{32'hc1489832, 32'hc2928391, 32'hc10fbe75, 32'hc1ee0f3e, 32'hc2a53919, 32'h41f94445, 32'h42939529, 32'hbf864629};
test_weights[19232:19239] = '{32'hc1b38974, 32'h42b43f70, 32'hc29ae171, 32'h3f16b595, 32'hc2417502, 32'hc281fc6a, 32'h42b63f98, 32'hc002264f};
test_bias[2404:2404] = '{32'h4237c470};
test_output[2404:2404] = '{32'h4541bfc7};
test_input[19240:19247] = '{32'hc11a5fa2, 32'hc2bc149e, 32'h3f9b6f4f, 32'hc28800ab, 32'hc290db14, 32'h41a5e4e2, 32'hc1ba59cf, 32'hc28f3207};
test_weights[19240:19247] = '{32'h42b23bb9, 32'h41396343, 32'h41d135e0, 32'hc26f9df8, 32'hc256d5cc, 32'hc26dbc7a, 32'hc1a59fbf, 32'h42a9bbc8};
test_bias[2405:2405] = '{32'h4256914f};
test_output[2405:2405] = '{32'hc435bcd7};
test_input[19248:19255] = '{32'h427c34a2, 32'h41e1d2fe, 32'h423d0fb5, 32'hc259b27f, 32'h429567da, 32'hc210d081, 32'h4272d03c, 32'hc1e77b9f};
test_weights[19248:19255] = '{32'hc299e8d3, 32'h42b6e5a2, 32'hc2856ed3, 32'h42b98800, 32'h4206f190, 32'h4082acef, 32'hc1ad4b08, 32'h417414f7};
test_bias[2406:2406] = '{32'h419aaabc};
test_output[2406:2406] = '{32'hc619b5d8};
test_input[19256:19263] = '{32'h42085f15, 32'hc286211e, 32'h42574af4, 32'h42961282, 32'hc1a2174e, 32'hc2752f38, 32'hc28b6b89, 32'hc2688eb1};
test_weights[19256:19263] = '{32'h42786c24, 32'h4007c4f6, 32'h408b09ab, 32'hc28d07db, 32'h41a72f46, 32'hc2a55d82, 32'hc2017e39, 32'hc19a58e7};
test_bias[2407:2407] = '{32'hc168ca36};
test_output[2407:2407] = '{32'h4599f2be};
test_input[19264:19271] = '{32'hc200c5d0, 32'h41f2df32, 32'hc28d8c81, 32'h42378315, 32'h427d83e7, 32'h42962265, 32'h42a3ed27, 32'hc2c33577};
test_weights[19264:19271] = '{32'hc2b59196, 32'h428aae7c, 32'hc29a365a, 32'hc1296162, 32'h42b330b1, 32'hc2419f77, 32'hc0c67a67, 32'h42be19cd};
test_bias[2408:2408] = '{32'h42a9ed68};
test_output[2408:2408] = '{32'h4512738a};
test_input[19272:19279] = '{32'hc20df5f2, 32'h41e9a445, 32'hc2815de0, 32'h41636d12, 32'hc1bb0af2, 32'hc2afc78e, 32'hc19875c3, 32'hc1c7fafa};
test_weights[19272:19279] = '{32'h4245d7a2, 32'hc27306ab, 32'h42b0f69b, 32'hc2b6edd7, 32'h42b6a055, 32'hc25a9bfa, 32'hc2bddecc, 32'hc29a84b6};
test_bias[2409:2409] = '{32'hc2008a60};
test_output[2409:2409] = '{32'hc5828293};
test_input[19280:19287] = '{32'h418602ab, 32'hc169a53a, 32'hc20ef611, 32'h4247beb3, 32'hc229ca4f, 32'h4219543a, 32'h42200fa6, 32'hc1da1c85};
test_weights[19280:19287] = '{32'h41cbc2c9, 32'h41f7e090, 32'hc20b9e75, 32'h42544b1d, 32'hc295ccbc, 32'hc281d279, 32'h42bfa22f, 32'hc24fb700};
test_bias[2410:2410] = '{32'h42a130ff};
test_output[2410:2410] = '{32'h461a967e};
test_input[19288:19295] = '{32'hc0e0e853, 32'hc103e23c, 32'hc127d9b4, 32'h42469330, 32'h4264ebc4, 32'h41ca2e61, 32'hc278d5dd, 32'h4221448c};
test_weights[19288:19295] = '{32'h4299a52c, 32'hc280268f, 32'h42821211, 32'h41b8ba33, 32'h4287fe24, 32'h42b6e631, 32'h426969c9, 32'h41324c15};
test_bias[2411:2411] = '{32'hc2c1add4};
test_output[2411:2411] = '{32'h455313da};
test_input[19296:19303] = '{32'h42bccc9f, 32'hc2b85466, 32'hc29fed02, 32'h408905c3, 32'h420cd4d1, 32'h420fd16d, 32'hc10873b4, 32'h40e647c6};
test_weights[19296:19303] = '{32'hc1227f30, 32'hc28d8e7a, 32'hc1818b2e, 32'h408b518b, 32'h412586f9, 32'hc287a44f, 32'hc1df849d, 32'hc1d25cfd};
test_bias[2412:2412] = '{32'hc2ab678b};
test_output[2412:2412] = '{32'h4594f91a};
test_input[19304:19311] = '{32'hc2779d38, 32'h428c5fc8, 32'h428af9d0, 32'hc1e97677, 32'h415a793c, 32'h425290f3, 32'hc28fda4c, 32'hc17250fc};
test_weights[19304:19311] = '{32'hc23a4d62, 32'h42b0454c, 32'h4236030a, 32'hc296d498, 32'h40e2e1ee, 32'hc1dc4c50, 32'hc274c3f1, 32'h42649124};
test_bias[2413:2413] = '{32'h42b7007b};
test_output[2413:2413] = '{32'h468284f2};
test_input[19312:19319] = '{32'hc15e81fe, 32'hc2494bac, 32'hc0e9fcd3, 32'hc2730248, 32'hc25edb1f, 32'hc284159a, 32'hc272692c, 32'h42a57a81};
test_weights[19312:19319] = '{32'hc21002d6, 32'hc2390591, 32'h429b16ba, 32'hc1c58106, 32'hc2ae4913, 32'h42828677, 32'hc229f3fc, 32'h412bd815};
test_bias[2414:2414] = '{32'hc1a04c9e};
test_output[2414:2414] = '{32'h45f22e18};
test_input[19320:19327] = '{32'h42771fc6, 32'hc248fe73, 32'hbfa75ebb, 32'hc2be5403, 32'h423fdeb6, 32'hc2b73fa5, 32'h4294acf4, 32'hc21d1d7f};
test_weights[19320:19327] = '{32'hc24724d3, 32'h421ad1da, 32'hc247730a, 32'h4094c13d, 32'h4288f7ae, 32'hc0dace55, 32'h42300c80, 32'hc29e0aa9};
test_bias[2415:2415] = '{32'hc2855756};
test_output[2415:2415] = '{32'h4596b482};
test_input[19328:19335] = '{32'hc25e5951, 32'h42428f9e, 32'hc1707a63, 32'h42577876, 32'h41e870ab, 32'h42866eb7, 32'h42afd4cf, 32'h4280c051};
test_weights[19328:19335] = '{32'hc1d755b5, 32'h426045a3, 32'h428b1155, 32'hc1d8f828, 32'hc27964ea, 32'h417ed795, 32'h40a7edb9, 32'h42110f5a};
test_bias[2416:2416] = '{32'h418e8c18};
test_output[2416:2416] = '{32'h456ce2ca};
test_input[19336:19343] = '{32'hc03b5688, 32'hc299228e, 32'h422cfb5f, 32'hc1c82895, 32'hc28835fb, 32'hc2af8126, 32'h42a357c8, 32'hc26f5515};
test_weights[19336:19343] = '{32'hc1a68224, 32'hc2209b8b, 32'h42b95d93, 32'h4218f60d, 32'hc2c4310f, 32'h42c4f58e, 32'h41e56322, 32'h4284693d};
test_bias[2417:2417] = '{32'hc2bb3a34};
test_output[2417:2417] = '{32'h451d08e2};
test_input[19344:19351] = '{32'hc2324c33, 32'h4274a673, 32'hc29b9d00, 32'hc15afede, 32'h41b2e412, 32'hc2517efd, 32'h40ee8b2a, 32'hc24a1467};
test_weights[19344:19351] = '{32'hc2758c34, 32'hc15a0fe2, 32'h429577c4, 32'h41eb05a1, 32'hc1d8f5ac, 32'hc163d316, 32'h429cf4bb, 32'h429784ba};
test_bias[2418:2418] = '{32'hc1222a71};
test_output[2418:2418] = '{32'hc5e81abe};
test_input[19352:19359] = '{32'h41f6acc4, 32'h42a1dc64, 32'hc1b84f27, 32'hc2547d00, 32'hc29fd0f6, 32'h421a5b02, 32'hc053c21e, 32'h40d1a3d8};
test_weights[19352:19359] = '{32'hc2a70c2b, 32'hc22cb0dd, 32'hc15b2d07, 32'hc23ab265, 32'hc1b81773, 32'hbed20e49, 32'hc1e71dc8, 32'h429bb6f5};
test_bias[2419:2419] = '{32'hc242cb8b};
test_output[2419:2419] = '{32'hc45f9c47};
test_input[19360:19367] = '{32'h4126a2b0, 32'hc255f798, 32'hc2559e2d, 32'hc2a6d951, 32'hc16eb1cc, 32'h42736650, 32'h42a3c115, 32'h40d4a98c};
test_weights[19360:19367] = '{32'h42778a32, 32'hc2a8e2e4, 32'h4235d94a, 32'h42964861, 32'hc2751bf4, 32'h41f1b687, 32'hc29fcdf2, 32'hc2853348};
test_bias[2420:2420] = '{32'hc2590dd3};
test_output[2420:2420] = '{32'hc5f46aa0};
test_input[19368:19375] = '{32'hc22f3ee7, 32'h42bf3d70, 32'h4102f2a4, 32'h41fafa1d, 32'h420e058a, 32'h41a55f84, 32'hc20d9246, 32'h424db343};
test_weights[19368:19375] = '{32'h428ff335, 32'hc26d9b06, 32'h41d4def7, 32'h41c2a2a7, 32'h4268b094, 32'hc2a273c9, 32'hc25a09cf, 32'hc21a78a4};
test_bias[2421:2421] = '{32'hc223ee9e};
test_output[2421:2421] = '{32'hc5ec5c63};
test_input[19376:19383] = '{32'h41f7763e, 32'hc24d3f67, 32'h42bd0d95, 32'hc2c28dd1, 32'h42bef27b, 32'hc180c3ad, 32'h42b0687f, 32'h426afd74};
test_weights[19376:19383] = '{32'hbf663ec4, 32'h422512f7, 32'hc29f76ff, 32'h401e00e6, 32'h42c7347f, 32'h41fa3369, 32'hc2263cfc, 32'h426e7ef9};
test_bias[2422:2422] = '{32'hc28e5eac};
test_output[2422:2422] = '{32'hc48fcff5};
test_input[19384:19391] = '{32'hc15dcc8f, 32'hc1c98485, 32'h410e7ed4, 32'hc2735ca4, 32'h41be7324, 32'hbf42f8b4, 32'h424d8e9f, 32'hc2aeb566};
test_weights[19384:19391] = '{32'hc289294b, 32'h42a44a18, 32'h421d0d2a, 32'h41884d3e, 32'hc1edd3d0, 32'h429305de, 32'hc2155b31, 32'h42bfa333};
test_bias[2423:2423] = '{32'h42ad6b62};
test_output[2423:2423] = '{32'hc6478dae};
test_input[19392:19399] = '{32'hc1d8cdf6, 32'h401a5fe0, 32'h42116aab, 32'hc127fc28, 32'hc282c5dd, 32'h42c07dc3, 32'h42715d02, 32'h41a1aa34};
test_weights[19392:19399] = '{32'h42517dec, 32'h428d029f, 32'h41c58062, 32'hc25f7846, 32'hc248b60d, 32'hc2721384, 32'hc2a05cdc, 32'h42338b93};
test_bias[2424:2424] = '{32'h40cb857b};
test_output[2424:2424] = '{32'hc5c2cdf8};
test_input[19400:19407] = '{32'h412bdb07, 32'hc29533c2, 32'hc2ad399d, 32'h429e7d9d, 32'hc243ec57, 32'h42b268d9, 32'hc250cfec, 32'h4109bfca};
test_weights[19400:19407] = '{32'h40af12de, 32'h4284b4be, 32'h419f7e73, 32'h42a5c7a0, 32'hc21b6883, 32'hc2bf9414, 32'hc253b0ce, 32'hc1ed0fb9};
test_bias[2425:2425] = '{32'h429c5531};
test_output[2425:2425] = '{32'hc5804ba2};
test_input[19408:19415] = '{32'h42beae20, 32'hc27860a0, 32'h4283c2c5, 32'h4284bc3a, 32'hc252abfc, 32'hc1b97244, 32'h410fb1bf, 32'h426b3205};
test_weights[19408:19415] = '{32'h3fda927e, 32'h4272e8fc, 32'hc2a43228, 32'hc29855e1, 32'hc22681dd, 32'h429c760d, 32'h41d772f4, 32'h420ff462};
test_bias[2426:2426] = '{32'h4244bc2e};
test_output[2426:2426] = '{32'hc63056a4};
test_input[19416:19423] = '{32'hc2c7a9a2, 32'h41e3c452, 32'h42817abe, 32'h4285f445, 32'hc1a9d597, 32'h42a1ae15, 32'hc2b7c1c5, 32'hc265640e};
test_weights[19416:19423] = '{32'h425c3d85, 32'h420bafb4, 32'hc29ad1e3, 32'hc26184a3, 32'hc1dc87bc, 32'h423b6503, 32'hc2a933cc, 32'h42bc4179};
test_bias[2427:2427] = '{32'hc1934f70};
test_output[2427:2427] = '{32'hc5cd0876};
test_input[19424:19431] = '{32'hc29360c1, 32'hc051466c, 32'hc2be2ab0, 32'hc2a61ecf, 32'hc28ed405, 32'hc290f980, 32'hc133fcf2, 32'h42afbda9};
test_weights[19424:19431] = '{32'hc2ab50f0, 32'hc291467e, 32'h41a0fc1b, 32'hc2b34e36, 32'h428a31f3, 32'h42924219, 32'hc2c5c472, 32'hc07b33d8};
test_bias[2428:2428] = '{32'hc237b62a};
test_output[2428:2428] = '{32'h45208d9a};
test_input[19432:19439] = '{32'hc284ada2, 32'h41946506, 32'h41392358, 32'h41c62d75, 32'h4282b296, 32'hc2942741, 32'hc22cbf49, 32'hc2659213};
test_weights[19432:19439] = '{32'h4207ec0d, 32'h42860e0e, 32'h41cbdd14, 32'hc2562b27, 32'h42adbfc6, 32'h403b70fd, 32'h42b4e409, 32'hc116c229};
test_bias[2429:2429] = '{32'h429d561d};
test_output[2429:2429] = '{32'h43032db2};
test_input[19440:19447] = '{32'h427bba7b, 32'hc28be35d, 32'hc1532b72, 32'h4248d737, 32'hc2842600, 32'hc15b151d, 32'hc24d1682, 32'hc118dd04};
test_weights[19440:19447] = '{32'hc127f7cb, 32'h4280356e, 32'h42595275, 32'h4293bc0c, 32'h424f8ce4, 32'hc2a5e68d, 32'h426ad90a, 32'hc2b474ef};
test_bias[2430:2430] = '{32'hc2529498};
test_output[2430:2430] = '{32'hc5cfb078};
test_input[19448:19455] = '{32'h4200f81a, 32'hc2c0ccb4, 32'hc23a99e0, 32'h41446564, 32'h42be7ed4, 32'hc2b5a78c, 32'hc2c1fef4, 32'h419a0d0c};
test_weights[19448:19455] = '{32'h41a103a5, 32'h41436071, 32'hc23c5221, 32'hc1b7d118, 32'h42ac2e79, 32'h429bf0f9, 32'h428b9625, 32'hc2becbd4};
test_bias[2431:2431] = '{32'hc270802f};
test_output[2431:2431] = '{32'hc5c0966b};
test_input[19456:19463] = '{32'hc0b6aa00, 32'h42a431f0, 32'hc1b6f196, 32'h418d8136, 32'hbd17ab89, 32'hc2aacd23, 32'h4285d897, 32'h4196c255};
test_weights[19456:19463] = '{32'h4222ead2, 32'h42b4bbb5, 32'h410d9291, 32'h42c4219c, 32'hc16e163e, 32'h41fd2f72, 32'h42b16121, 32'h412b029d};
test_bias[2432:2432] = '{32'hc187dd60};
test_output[2432:2432] = '{32'h463da0eb};
test_input[19464:19471] = '{32'h40ff003c, 32'hc1ee62de, 32'h4224cf75, 32'hc0cdc26b, 32'hc28e100d, 32'hc292b6a4, 32'h4281f46f, 32'hc28a0991};
test_weights[19464:19471] = '{32'hc27e37b6, 32'hc297719e, 32'h42b4c1ab, 32'h420afacf, 32'h428fe065, 32'h418afe68, 32'h42369465, 32'h4295d3f7};
test_bias[2433:2433] = '{32'hc2836739};
test_output[2433:2433] = '{32'hc554c539};
test_input[19472:19479] = '{32'hc20f431f, 32'h42bf6e26, 32'hc25d5161, 32'h4260a939, 32'hc2ab295a, 32'h426aba5d, 32'h42329c5d, 32'h41907270};
test_weights[19472:19479] = '{32'hc1e2cffa, 32'hc28b9537, 32'h42bc5695, 32'hc2b19a33, 32'hc2332375, 32'h428b96d2, 32'h42bdca4b, 32'h420a291e};
test_bias[2434:2434] = '{32'hc1c97839};
test_output[2434:2434] = '{32'hc541a5bf};
test_input[19480:19487] = '{32'hc0a0a92b, 32'hc0b60e0b, 32'hc2c4f4a9, 32'hc194101c, 32'hc2c6df97, 32'hc2a8af58, 32'hc1b4e82c, 32'hc28df129};
test_weights[19480:19487] = '{32'hc13c675e, 32'h428ba437, 32'h429e4cd1, 32'hc29889ac, 32'h41192ae0, 32'hc29aeab3, 32'hc1d5ce1d, 32'hc28b7ada};
test_bias[2435:2435] = '{32'hc2aa3475};
test_output[2435:2435] = '{32'h458746b9};
test_input[19488:19495] = '{32'h42779c86, 32'hc1fb1220, 32'hc2543987, 32'hc210b842, 32'h426c4e62, 32'h427cfba9, 32'hc2a0eace, 32'h406dbdc7};
test_weights[19488:19495] = '{32'h4231e958, 32'hc181b4a8, 32'hc243ca95, 32'hc2be0bac, 32'hc14048d7, 32'hc22a80bb, 32'h42a1576a, 32'h3f69ab03};
test_bias[2436:2436] = '{32'hc289f080};
test_output[2436:2436] = '{32'hc4264373};
test_input[19496:19503] = '{32'hc2c7b07f, 32'hc2a35c60, 32'hc2a7f17b, 32'hc1da5875, 32'hc29b012f, 32'hc15bd82a, 32'h420e140c, 32'hc0037d17};
test_weights[19496:19503] = '{32'hc147fe89, 32'h42189ad8, 32'h41a515fd, 32'hc221696c, 32'hc1f1e6e6, 32'h42718207, 32'hc217037f, 32'hc1536ccd};
test_bias[2437:2437] = '{32'hc2ae30c2};
test_output[2437:2437] = '{32'hc5152ac6};
test_input[19504:19511] = '{32'hc20feed6, 32'h42ab2d04, 32'h42c3acc8, 32'hc298a624, 32'hc1e36b05, 32'h42438b76, 32'hc0893346, 32'h4132dc0b};
test_weights[19504:19511] = '{32'hbed670f3, 32'h42a07899, 32'h42383fc2, 32'h42ae358c, 32'hc2478919, 32'hc2986773, 32'h427f8de4, 32'hc29c8362};
test_bias[2438:2438] = '{32'h41c90f8a};
test_output[2438:2438] = '{32'h44a3bcd0};
test_input[19512:19519] = '{32'h4227cac5, 32'h42c41ebb, 32'hc255b6f0, 32'hc29a0b00, 32'h4027b935, 32'hc24e0703, 32'hc1a4c75e, 32'h425b6433};
test_weights[19512:19519] = '{32'h4215dee0, 32'hc275d84b, 32'hc2b4794c, 32'h418d5c00, 32'hc0e8c7ea, 32'hc186f90d, 32'h42442df5, 32'h41116791};
test_bias[2439:2439] = '{32'h40a3aca1};
test_output[2439:2439] = '{32'hc422e77f};
test_input[19520:19527] = '{32'hc2322967, 32'h418543fd, 32'h41fd6edd, 32'h41db2c17, 32'h413be864, 32'h42079085, 32'h42c570c6, 32'h41479221};
test_weights[19520:19527] = '{32'hc23b658f, 32'hc2604d5d, 32'hbfaf7633, 32'hc28d87b8, 32'h42a2fdb8, 32'h4286623f, 32'hc2c682e8, 32'hc27a8c52};
test_bias[2440:2440] = '{32'hc2825e45};
test_output[2440:2440] = '{32'hc600c11e};
test_input[19528:19535] = '{32'hc245c43b, 32'h410d5784, 32'hc15108a1, 32'h42aef10a, 32'h4277e8f3, 32'hc237b8b1, 32'h4258e465, 32'h427ca216};
test_weights[19528:19535] = '{32'h40a156d2, 32'h4250f218, 32'hc28cc6ee, 32'hc1a3cdae, 32'hc24a8a0a, 32'hc21e8b83, 32'h40f680bf, 32'h40e81760};
test_bias[2441:2441] = '{32'hc1c958f6};
test_output[2441:2441] = '{32'hc48ccae7};
test_input[19536:19543] = '{32'h419ed2d3, 32'h40855550, 32'hc1e3d722, 32'h41773c1f, 32'hc1608e14, 32'h422fb639, 32'h41f76116, 32'h4291b0fe};
test_weights[19536:19543] = '{32'h42879d7c, 32'h429ad7ee, 32'h42a4f6bc, 32'h42bfcb3f, 32'hc1ab7020, 32'h4266f6c3, 32'hc1ea25d4, 32'hc231309c};
test_bias[2442:2442] = '{32'h425b76bf};
test_output[2442:2442] = '{32'hc3db2e86};
test_input[19544:19551] = '{32'h427bbe0f, 32'hc2812da9, 32'hc269c1ff, 32'hc28a21d9, 32'hc1a7e8b3, 32'h41173d54, 32'hc226aca1, 32'hc27d7475};
test_weights[19544:19551] = '{32'h429cd333, 32'hc272ccc7, 32'h3f6f9ae0, 32'hc2a604fe, 32'hc2142557, 32'hc20c9dde, 32'hc23643ab, 32'h428f2a87};
test_bias[2443:2443] = '{32'hc21e07db};
test_output[2443:2443] = '{32'h464039a4};
test_input[19552:19559] = '{32'hc29e0abf, 32'hc2a13f32, 32'hc2c48ce9, 32'h42aaf006, 32'hc19107e0, 32'hc2c4b7b3, 32'h429dfe82, 32'h42ba0f7c};
test_weights[19552:19559] = '{32'h42a8200e, 32'hc2195702, 32'hc2aaff2a, 32'h42a0fbef, 32'h42194fc5, 32'h42adc740, 32'h4262efd9, 32'hc2a60909};
test_bias[2444:2444] = '{32'hc1535cd2};
test_output[2444:2444] = '{32'hc43f709f};
test_input[19560:19567] = '{32'hc1b12b10, 32'h41aa1e80, 32'h41788051, 32'h42ac3c69, 32'hc23655c9, 32'h42972afe, 32'h42aeac68, 32'hc1c60ff2};
test_weights[19560:19567] = '{32'hc2bc6dd0, 32'hc225dc39, 32'hc203cd75, 32'h42ae2831, 32'h42500281, 32'h428e7568, 32'h42a3c718, 32'hc2091ef3};
test_bias[2445:2445] = '{32'h4206b692};
test_output[2445:2445] = '{32'h46964f31};
test_input[19568:19575] = '{32'hc1bfec12, 32'h4014557f, 32'hc2ba69b7, 32'hc2c61642, 32'hc29eab1c, 32'h4260e523, 32'h41ce1ce0, 32'h4246a029};
test_weights[19568:19575] = '{32'h41c8acd6, 32'hc2889c65, 32'hc077a223, 32'h4129690b, 32'h427ef614, 32'hc137bfdc, 32'hc2667609, 32'hc2aad132};
test_bias[2446:2446] = '{32'h42b9e148};
test_output[2446:2446] = '{32'hc647bcac};
test_input[19576:19583] = '{32'hc1a7714d, 32'h42c2463a, 32'h42a6e5b5, 32'hc20f30f9, 32'hc2abc64e, 32'hc18ba4cd, 32'h41d12139, 32'hc2a68d2c};
test_weights[19576:19583] = '{32'h42018f6a, 32'h40d1d49e, 32'h40f6c09a, 32'hc1eae51a, 32'hc27b9a4e, 32'hc17d4f16, 32'h42b6ff2e, 32'hc1d94dcc};
test_bias[2447:2447] = '{32'hc2680063};
test_output[2447:2447] = '{32'h463a60cb};
test_input[19584:19591] = '{32'h429a6b63, 32'h42a67a7f, 32'hc11e6121, 32'hc0bab300, 32'hc1177f9a, 32'h42265ea0, 32'hc1b8e2da, 32'hc0cb6332};
test_weights[19584:19591] = '{32'hc18b9d7b, 32'hc250fb86, 32'h4184b574, 32'h42984bb4, 32'h42be5f73, 32'h4281213c, 32'hc2afd823, 32'h4289c7bc};
test_bias[2448:2448] = '{32'h4235ca97};
test_output[2448:2448] = '{32'hc534128c};
test_input[19592:19599] = '{32'h423ee5e6, 32'h412d8965, 32'hc1adc037, 32'hc21ddf73, 32'hc2809665, 32'hc2093b29, 32'h42438e6d, 32'hc2a8aefd};
test_weights[19592:19599] = '{32'hc14a04e9, 32'h41b3c998, 32'h42a4a4b4, 32'hc2690709, 32'h429d2cbc, 32'h41127fd6, 32'h414084ae, 32'hc2a472c1};
test_bias[2449:2449] = '{32'hc212e5a7};
test_output[2449:2449] = '{32'h450e02e9};
test_input[19600:19607] = '{32'h428bcc51, 32'h428965ba, 32'hc28dc36c, 32'h42c1a56d, 32'hc2142438, 32'h42034d31, 32'h4229e5c4, 32'hc2bae2e6};
test_weights[19600:19607] = '{32'h411c4c60, 32'hc17db297, 32'hc2c2ae43, 32'hc2a8808d, 32'hc1ae554c, 32'hc2c0d694, 32'hc1c39588, 32'h424812c1};
test_bias[2450:2450] = '{32'hc29114e1};
test_output[2450:2450] = '{32'hc6193c20};
test_input[19608:19615] = '{32'hc2272cca, 32'h41c17b99, 32'hc1babaac, 32'hc2965106, 32'hc0fa4bda, 32'h41a44763, 32'h4052d66c, 32'h41b8a2aa};
test_weights[19608:19615] = '{32'h4230e04e, 32'h428b8923, 32'hc2795ea8, 32'h42b89458, 32'hc15b5a66, 32'h42b9c2f3, 32'h42b87203, 32'hc2a36b7e};
test_bias[2451:2451] = '{32'h41fce32b};
test_output[2451:2451] = '{32'hc5a1ce3c};
test_input[19616:19623] = '{32'h42c6ced9, 32'hc2be26da, 32'hc2685915, 32'hc22006dd, 32'hc1e6a372, 32'h42ab039b, 32'h42b2abd5, 32'hc2ac3616};
test_weights[19616:19623] = '{32'h40821c0b, 32'hc2bed5e3, 32'hc2230017, 32'hc163aa20, 32'h42c0fc11, 32'hc142c39d, 32'hc2c1b3cd, 32'h42a662c7};
test_bias[2452:2452] = '{32'h42019a5f};
test_output[2452:2452] = '{32'hc5e0cc5f};
test_input[19624:19631] = '{32'hc2222599, 32'h428818b1, 32'hc0c41efa, 32'h4196627e, 32'hc272a865, 32'hc0f96823, 32'h41307fad, 32'h41bbe31c};
test_weights[19624:19631] = '{32'hc1a2a049, 32'hc2327c8f, 32'h42c671c3, 32'h429a51e8, 32'h4277fff3, 32'h429a77c3, 32'hc2904974, 32'hc21c84d7};
test_bias[2453:2453] = '{32'hc2844804};
test_output[2453:2453] = '{32'hc5ead130};
test_input[19632:19639] = '{32'h4281d740, 32'hc2a1dc05, 32'hc10bc92d, 32'hbfd0bb2d, 32'h425ea0f1, 32'h42b8f0d2, 32'hc18091ae, 32'h42c66539};
test_weights[19632:19639] = '{32'h42ab14af, 32'h42b416bb, 32'hc1aaf87a, 32'hc281e0e5, 32'h42b4c07a, 32'hc2881051, 32'h4273a94a, 32'h40e44788};
test_bias[2454:2454] = '{32'hc278e037};
test_output[2454:2454] = '{32'hc53dbc00};
test_input[19640:19647] = '{32'h42c6cb6a, 32'h4188c10b, 32'h41973099, 32'hc2023eeb, 32'h429d2924, 32'hc1c3cd56, 32'hc1b1ba54, 32'hc25311fc};
test_weights[19640:19647] = '{32'hc0175cdb, 32'hc2a391bc, 32'h42058167, 32'h401b9c39, 32'h426cb4c6, 32'h4209f84c, 32'h428e3e9b, 32'h42999e63};
test_bias[2455:2455] = '{32'hc2208a87};
test_output[2455:2455] = '{32'hc5384da9};
test_input[19648:19655] = '{32'hc1acb742, 32'h42aa56f9, 32'hc252d62c, 32'h41ba29c6, 32'h3f904dd1, 32'hc153f17d, 32'hc1f2b34f, 32'h42b65c9c};
test_weights[19648:19655] = '{32'h42b88452, 32'hc26d71f9, 32'hc287bff8, 32'h42901b77, 32'h3fe4db6c, 32'hc2c1e41b, 32'h422e7bf5, 32'hc239ffbe};
test_bias[2456:2456] = '{32'h41fb29e5};
test_output[2456:2456] = '{32'hc5bcb741};
test_input[19656:19663] = '{32'hc2a9add1, 32'hc0219ef2, 32'h429d4946, 32'hc1ef1a74, 32'hc27af5ad, 32'h42313e47, 32'hc1673299, 32'hc2892263};
test_weights[19656:19663] = '{32'hc21b034f, 32'hc21bf358, 32'hc2802bd5, 32'h416b7aca, 32'hc2a68ca6, 32'h424366d1, 32'hc2aaf59d, 32'h42834f6a};
test_bias[2457:2457] = '{32'hc105b350};
test_output[2457:2457] = '{32'h44fc98b9};
test_input[19664:19671] = '{32'h41d170cd, 32'hc24f7837, 32'h3fa455de, 32'hc20d8038, 32'hc2b28778, 32'hc2b96dde, 32'hc1ebfc33, 32'hc0a9ca4b};
test_weights[19664:19671] = '{32'hc1988606, 32'h413c9723, 32'hc0ec5ab7, 32'hc244b606, 32'hc2666260, 32'h425ddbcd, 32'h42aa4a5f, 32'h42a8df38};
test_bias[2458:2458] = '{32'hc1a16f80};
test_output[2458:2458] = '{32'hc5139362};
test_input[19672:19679] = '{32'hc1a1ed40, 32'hc2717b37, 32'h41758762, 32'hc2965567, 32'h4270c24c, 32'hc20c896a, 32'hc2975c30, 32'h421becf0};
test_weights[19672:19679] = '{32'hc29ffe38, 32'h420a018c, 32'h4250e22b, 32'hc29a61ef, 32'hc1f387df, 32'hc2918d50, 32'hc1500ca0, 32'h3f689c3c};
test_bias[2459:2459] = '{32'h42980a82};
test_output[2459:2459] = '{32'h45f8c0bd};
test_input[19680:19687] = '{32'hc27ab1bb, 32'h421d4467, 32'h429b0752, 32'hc2143bb0, 32'h419ef044, 32'hc060e61c, 32'hc26425ae, 32'h42869acb};
test_weights[19680:19687] = '{32'hc24ecf29, 32'hc26c84b1, 32'h42bebc2b, 32'hc2190dc5, 32'h420abe75, 32'hc2b083e2, 32'h426a8479, 32'hc287a29c};
test_bias[2460:2460] = '{32'hc17190e3};
test_output[2460:2460] = '{32'h452f1c0b};
test_input[19688:19695] = '{32'h41b866eb, 32'h426aa08e, 32'hc20c9e62, 32'hc20fc3c3, 32'h426b6bd0, 32'h42b77f12, 32'h42c4ac47, 32'h4188bbc7};
test_weights[19688:19695] = '{32'hc1858421, 32'hc2904479, 32'hc257a079, 32'h42362753, 32'h404c5ac7, 32'h418483ab, 32'hc23601af, 32'h4292c5d1};
test_bias[2461:2461] = '{32'h41a552c8};
test_output[2461:2461] = '{32'hc5b6ca67};
test_input[19696:19703] = '{32'h42a8eb49, 32'hc0d13175, 32'hc1418e08, 32'h429013ce, 32'h4208735d, 32'h42b5a5fe, 32'h3ffce883, 32'hc1e62949};
test_weights[19696:19703] = '{32'h42856795, 32'h41729e09, 32'h422ed8ec, 32'hc2a22f75, 32'h429032ee, 32'h429734e6, 32'h42af0003, 32'hc23e7cb9};
test_bias[2462:2462] = '{32'hc166d75c};
test_output[2462:2462] = '{32'h461c8a51};
test_input[19704:19711] = '{32'h4293cbcd, 32'h3f3d1c0a, 32'h420ff373, 32'hc1dea3f1, 32'h42b7d33b, 32'hc2c2caed, 32'h410128b0, 32'h3ef7713e};
test_weights[19704:19711] = '{32'hc20dd8f5, 32'hc1478722, 32'hc139dee6, 32'hc271981e, 32'hc2a8da97, 32'hc2a9624c, 32'hc26a8ddd, 32'h42762166};
test_bias[2463:2463] = '{32'h42a485c2};
test_output[2463:2463] = '{32'hc49af052};
test_input[19712:19719] = '{32'hc26f47f0, 32'h4295c172, 32'h423f96ff, 32'h42c5041d, 32'h42b29025, 32'hc1da9fb8, 32'h4109924e, 32'h418e1d73};
test_weights[19712:19719] = '{32'h42a64e01, 32'hc04ec387, 32'h42714528, 32'hc1aeeb37, 32'h42adef7d, 32'h429873a9, 32'h427793dd, 32'h429a94c5};
test_bias[2464:2464] = '{32'hc2b28f02};
test_output[2464:2464] = '{32'h453c886b};
test_input[19720:19727] = '{32'h4287485c, 32'hc1d36743, 32'hc2a5f5ac, 32'h417c6209, 32'h429c7290, 32'hc123f2a5, 32'h419f5877, 32'h422e3e6b};
test_weights[19720:19727] = '{32'hc222e822, 32'h40f23294, 32'h420f4a6f, 32'h413d435a, 32'h3fdbe387, 32'hc2add3ed, 32'h4191e532, 32'hc1c5eaee};
test_bias[2465:2465] = '{32'h4243c15a};
test_output[2465:2465] = '{32'hc5a82a92};
test_input[19728:19735] = '{32'h42409d59, 32'hc261b44d, 32'hc22e85e9, 32'hc2b74101, 32'hc2324dd4, 32'hc2329ba2, 32'h412633c1, 32'h42bab2d8};
test_weights[19728:19735] = '{32'hbfd7c3e3, 32'h42a5ecbd, 32'h42c6f326, 32'h42bc2f23, 32'h41c0fd0f, 32'h4221d6c8, 32'hbf4045ba, 32'hc21aae11};
test_bias[2466:2466] = '{32'hc247edd3};
test_output[2466:2466] = '{32'hc6bda2fa};
test_input[19736:19743] = '{32'h41700146, 32'h428d7cf9, 32'hc24c06c8, 32'hbffe1b02, 32'h42ac83c7, 32'h42c7bc34, 32'hc2617da6, 32'h4221f198};
test_weights[19736:19743] = '{32'hc29983d9, 32'h4233b640, 32'hc281f57c, 32'h4237964a, 32'h4248429f, 32'hc29e3ae8, 32'hc272225a, 32'h426c572c};
test_bias[2467:2467] = '{32'h41c7ddef};
test_output[2467:2467] = '{32'h45ea4a18};
test_input[19744:19751] = '{32'h420bda1e, 32'h41c0c848, 32'hc29d2f45, 32'hc2b6ddf9, 32'hc1685b4f, 32'h42632fa4, 32'hc26acd64, 32'hc033e86c};
test_weights[19744:19751] = '{32'hc29be7b9, 32'hc1a359f1, 32'hc22e395f, 32'h418bcb68, 32'hc1a15c6f, 32'hc2842595, 32'hc25ac5df, 32'h41b1f960};
test_bias[2468:2468] = '{32'hc20b6ca7};
test_output[2468:2468] = '{32'hc4d95899};
test_input[19752:19759] = '{32'hc1c88c19, 32'hc22e69da, 32'h429f6da4, 32'h422b9b48, 32'h423b23d0, 32'h41fab70b, 32'h4110f371, 32'h429769aa};
test_weights[19752:19759] = '{32'hc299258c, 32'h3ef98e07, 32'hbfe3a606, 32'hc2bfa31a, 32'h41f3a33b, 32'h429342b6, 32'h42b8a302, 32'hc28ae316};
test_bias[2469:2469] = '{32'h413c4559};
test_output[2469:2469] = '{32'hc53d7133};
test_input[19760:19767] = '{32'h427db050, 32'hc032cb7c, 32'hc2bbbb15, 32'hc2b7e738, 32'hc2be97dc, 32'h42c0be14, 32'hc258740e, 32'hc12a9055};
test_weights[19760:19767] = '{32'hc2a89d0c, 32'h42ad9674, 32'hc29c36ed, 32'h4206f6ad, 32'h40104f89, 32'hc2b72f97, 32'h41346856, 32'hc1869863};
test_bias[2470:2470] = '{32'hc11b7b19};
test_output[2470:2470] = '{32'hc6296ab3};
test_input[19768:19775] = '{32'hc2b6b678, 32'hc0d96f0b, 32'hc2a3297a, 32'hc1f89dad, 32'h40fd9854, 32'hc285423e, 32'hc28c63d9, 32'h428159e6};
test_weights[19768:19775] = '{32'hc2a6701e, 32'h42071051, 32'h411db554, 32'h407d316d, 32'h429f82d9, 32'h42958a94, 32'hc21f031b, 32'hc2bd05cc};
test_bias[2471:2471] = '{32'h42529cde};
test_output[2471:2471] = '{32'hc492a7ee};
test_input[19776:19783] = '{32'hc2483bc3, 32'hc281caae, 32'hc2983406, 32'hc23d439d, 32'h42557f0c, 32'hc26458bf, 32'hc29c8f8d, 32'hc265d7d3};
test_weights[19776:19783] = '{32'hc2ad6268, 32'hc224294a, 32'hc293b22a, 32'hc1d59974, 32'h42afc35c, 32'hc0de25e8, 32'hc1f7434d, 32'hc1dce118};
test_bias[2472:2472] = '{32'hc292c2a1};
test_output[2472:2472] = '{32'h46b2f392};
test_input[19784:19791] = '{32'h41841378, 32'h421aadb6, 32'h412bca29, 32'hc27a5dd4, 32'h422430f5, 32'hc294c2db, 32'hc226d4e1, 32'h421da90d};
test_weights[19784:19791] = '{32'h428d538b, 32'hc2abf353, 32'h41fffe41, 32'hc227c6ce, 32'h41fbc7d5, 32'hc2660fe4, 32'hc25f3084, 32'hc2b7f882};
test_bias[2473:2473] = '{32'hc29d3086};
test_output[2473:2473] = '{32'h459c5e75};
test_input[19792:19799] = '{32'h41ad538f, 32'hc21f0881, 32'hc20b5df0, 32'hc067ab7d, 32'hc145b1df, 32'h410ce618, 32'hc220c03a, 32'h42c113a8};
test_weights[19792:19799] = '{32'hc1d89561, 32'h427da57e, 32'hc186989e, 32'h4100a756, 32'h42a3b985, 32'hc2a2bb66, 32'hc2bc2446, 32'h42734e59};
test_bias[2474:2474] = '{32'hc2b88fee};
test_output[2474:2474] = '{32'h45a50d87};
test_input[19800:19807] = '{32'hc2c7c9d6, 32'h42915607, 32'hc2a88aae, 32'h42b118cc, 32'h409c5334, 32'hc2b780dc, 32'hc292abfb, 32'hc2181c5a};
test_weights[19800:19807] = '{32'hc262dd7b, 32'hc2c66966, 32'hc19eff8d, 32'h41b166dd, 32'hc1efd33f, 32'h41d347ed, 32'hc2419a7e, 32'hc11d7b40};
test_bias[2475:2475] = '{32'h427ded71};
test_output[2475:2475] = '{32'h455b8a7d};
test_input[19808:19815] = '{32'hbfc73e47, 32'hc2ba9f64, 32'h4298ba44, 32'hbf916bc6, 32'h429273b8, 32'hc2c32bff, 32'h42486337, 32'h42588fbe};
test_weights[19808:19815] = '{32'h40cf9c6c, 32'hc1a780e0, 32'hc2c43cab, 32'h41bb0a87, 32'hc20bb737, 32'h42248bef, 32'hc23715f7, 32'hc287f8b7};
test_bias[2476:2476] = '{32'hc23aba33};
test_output[2476:2476] = '{32'hc68df04a};
test_input[19816:19823] = '{32'hc2a9128a, 32'hc2b6824d, 32'h42a2c0f6, 32'hc28e4d1b, 32'h42268731, 32'h3f6c4957, 32'hc29757fe, 32'h42a6eac9};
test_weights[19816:19823] = '{32'hc229c67a, 32'h425abe79, 32'hc17f9892, 32'hbda58776, 32'hc29b33c4, 32'hc0b5455c, 32'h420cea77, 32'hc1b9e511};
test_bias[2477:2477] = '{32'hc232c9f7};
test_output[2477:2477] = '{32'hc6255934};
test_input[19824:19831] = '{32'h41d7c5c1, 32'h4084b5e6, 32'h429e1d38, 32'h4283daf4, 32'hc245bfb1, 32'hc2644488, 32'h429fcbee, 32'h42637fa2};
test_weights[19824:19831] = '{32'hc257a4d9, 32'hc1eca50e, 32'h428addde, 32'h42626645, 32'h4221bf6b, 32'h41ab8327, 32'h412bd75b, 32'hc24d5bff};
test_bias[2478:2478] = '{32'h422f897c};
test_output[2478:2478] = '{32'h45163779};
test_input[19832:19839] = '{32'h4128382c, 32'hc268769a, 32'h423a32f4, 32'hc22c6bc4, 32'hc293d429, 32'h421ba1df, 32'h419597c7, 32'h420c769d};
test_weights[19832:19839] = '{32'h418253ff, 32'hc28092c8, 32'h41fc7e77, 32'hc2c22f91, 32'h427b557e, 32'hc29d0d16, 32'hc2ab286a, 32'h42b0b5a1};
test_bias[2479:2479] = '{32'hc234082d};
test_output[2479:2479] = '{32'h454f792c};
test_input[19840:19847] = '{32'h42180a27, 32'h4208eb50, 32'hc2417865, 32'hc2684257, 32'hc1abe05a, 32'h4259fedf, 32'h42c6a649, 32'h4298149b};
test_weights[19840:19847] = '{32'h42be27ee, 32'h42593511, 32'hc236d1c6, 32'hc242e095, 32'h4065b9b0, 32'h421cfccd, 32'h42970914, 32'h4105c461};
test_bias[2480:2480] = '{32'hc2c0827f};
test_output[2480:2480] = '{32'h46a10c6a};
test_input[19848:19855] = '{32'h3faa37e6, 32'hc25cddba, 32'hc284ec22, 32'h429932b4, 32'h42244735, 32'h429dbcd0, 32'h42ad667c, 32'hc2bc500c};
test_weights[19848:19855] = '{32'hc12e1c30, 32'hc14645a0, 32'h425c5256, 32'h41cd22c7, 32'h40b1f519, 32'h421c8c7f, 32'hc206f0b5, 32'hc12985e8};
test_bias[2481:2481] = '{32'hc2060756};
test_output[2481:2481] = '{32'h43a3c951};
test_input[19856:19863] = '{32'h40b6ca21, 32'h42ba5026, 32'h42c3896d, 32'hc29ae861, 32'h414bdaad, 32'hc2b2d751, 32'hc254ba35, 32'hc2b6df20};
test_weights[19856:19863] = '{32'h42af5695, 32'h4225b251, 32'hc21f21c6, 32'hc20023c3, 32'h42bcd070, 32'h42126604, 32'h427e1408, 32'h41dd940d};
test_bias[2482:2482] = '{32'hc28ee99a};
test_output[2482:2482] = '{32'hc59f649a};
test_input[19864:19871] = '{32'hc2c49e8a, 32'h42a8b23e, 32'h4210ecdf, 32'hc282374c, 32'hc27e598a, 32'hc2919965, 32'hc093fddc, 32'hc2c78a75};
test_weights[19864:19871] = '{32'hc2bdfbe9, 32'hc2c64f1d, 32'h418de4b6, 32'h415ef38c, 32'hc0d483bc, 32'hc1addcbe, 32'hc207b9aa, 32'h4087dda0};
test_bias[2483:2483] = '{32'h41d71c69};
test_output[2483:2483] = '{32'h451ab253};
test_input[19872:19879] = '{32'h42116d2e, 32'hc1d640cc, 32'hc24de8c6, 32'hc28591cc, 32'h42c2444e, 32'h42a690c7, 32'hc23ae668, 32'hc13edeae};
test_weights[19872:19879] = '{32'hbe0c87f8, 32'h4298c649, 32'h420a1dfd, 32'hc1fa002c, 32'hc135e7da, 32'h412f9792, 32'h42161e20, 32'hc1a8150e};
test_bias[2484:2484] = '{32'hbe26ecca};
test_output[2484:2484] = '{32'hc556aa16};
test_input[19880:19887] = '{32'h41f48b4b, 32'hc2c14ee5, 32'h42a17545, 32'hc24fb197, 32'h420affc3, 32'h422c3fd5, 32'h42a72d8b, 32'hc1c080a5};
test_weights[19880:19887] = '{32'h429ce505, 32'h4280ef07, 32'hc272878c, 32'hc2240e31, 32'hc148dd30, 32'h428c3103, 32'h42a0c448, 32'hc292c2da};
test_bias[2485:2485] = '{32'hc2b4d755};
test_output[2485:2485] = '{32'h4588d402};
test_input[19888:19895] = '{32'h427d00ac, 32'h41a35bfe, 32'h42c2b607, 32'h42b38370, 32'h418121c7, 32'hc29a8301, 32'h42826a3d, 32'h41ead2b5};
test_weights[19888:19895] = '{32'hc2b58495, 32'h41c21a8c, 32'hc20f3ff2, 32'h42125fce, 32'hc2a65496, 32'h42645260, 32'h41bddcd0, 32'h421c3a09};
test_bias[2486:2486] = '{32'hc29b6f9a};
test_output[2486:2486] = '{32'hc6061c53};
test_input[19896:19903] = '{32'h41a3bc02, 32'h41817cff, 32'h4188cce2, 32'hc2bf112b, 32'hc2b185ac, 32'hc299791c, 32'h420862c9, 32'hc264106d};
test_weights[19896:19903] = '{32'h420a0e73, 32'h421a7845, 32'h41ac25e4, 32'hc2acf205, 32'h428910f7, 32'h41a0f1fe, 32'hc2ac930b, 32'h429b3472};
test_bias[2487:2487] = '{32'hc2ad6690};
test_output[2487:2487] = '{32'hc59ffe3d};
test_input[19904:19911] = '{32'h4287ad62, 32'hc1904b99, 32'hc2880293, 32'h425d0ae6, 32'h42bdd8e7, 32'hc29f92f5, 32'hc293b71a, 32'h422287e2};
test_weights[19904:19911] = '{32'hc26829fa, 32'h42774d77, 32'hc2924ebf, 32'hc1f71b95, 32'hc206513b, 32'hc24aae9d, 32'hc0a63300, 32'h42510808};
test_bias[2488:2488] = '{32'hc29487aa};
test_output[2488:2488] = '{32'h44bbedcd};
test_input[19912:19919] = '{32'hc25f8343, 32'hc2029e7d, 32'h4281f220, 32'h4272c7e5, 32'hc2595545, 32'h425e8873, 32'hc2a8e9ba, 32'h42a3c742};
test_weights[19912:19919] = '{32'h426444ba, 32'hc2bb3169, 32'hc28a5aa9, 32'h427aa1de, 32'hc29b9532, 32'h4015c3f8, 32'h428dae55, 32'h42464646};
test_bias[2489:2489] = '{32'hc20d20da};
test_output[2489:2489] = '{32'h44c4b786};
test_input[19920:19927] = '{32'hc2029cd6, 32'h42466282, 32'h42abf466, 32'hc1c31f53, 32'hc1b0cb90, 32'h428db717, 32'hc04e4455, 32'h429f16a8};
test_weights[19920:19927] = '{32'hc29865b8, 32'h429bdce7, 32'hc292f0c5, 32'hc2c17e3c, 32'hc2022ddf, 32'hc245711d, 32'h42a3d709, 32'hc19bab49};
test_bias[2490:2490] = '{32'hc1cdd6a6};
test_output[2490:2490] = '{32'hc50abc94};
test_input[19928:19935] = '{32'hc2892d60, 32'h424285ba, 32'h41c68499, 32'h429ada1b, 32'h42b6f659, 32'hc1bede9e, 32'hc212eca5, 32'hc098b4f7};
test_weights[19928:19935] = '{32'hc1f5ff0a, 32'h42aeeb04, 32'hc12bc88d, 32'h416a6a50, 32'hc27793b6, 32'h424e813b, 32'h42a06264, 32'hc25ff3ed};
test_bias[2491:2491] = '{32'hc1e96c51};
test_output[2491:2491] = '{32'hc51433dc};
test_input[19936:19943] = '{32'hc2110111, 32'hc0c7dbb4, 32'hc2648620, 32'h42c72896, 32'hc1634a63, 32'hc2a54e17, 32'h42ab1428, 32'h423dcf52};
test_weights[19936:19943] = '{32'h422931b4, 32'hc11d050d, 32'h42c6cddf, 32'h42b604ab, 32'h429b0f0b, 32'hc2c67718, 32'h41c88f93, 32'h4265400e};
test_bias[2492:2492] = '{32'h4260a1e8};
test_output[2492:2492] = '{32'h4659b15a};
test_input[19944:19951] = '{32'hc19fb62f, 32'h42a0142a, 32'hc2bdea7b, 32'h42427d35, 32'hc2998c2f, 32'hc26b733c, 32'hc29f9c00, 32'hc22880e7};
test_weights[19944:19951] = '{32'hc2b7e27f, 32'h4268b337, 32'h42c4dbe7, 32'h426b0b60, 32'hc0b93148, 32'hc128553e, 32'hc258144a, 32'h42c0cf8d};
test_bias[2493:2493] = '{32'hc1bd941f};
test_output[2493:2493] = '{32'h44a180e6};
test_input[19952:19959] = '{32'h4071680a, 32'hc26660c0, 32'hc2c033d2, 32'hc29edff5, 32'hc2a4da19, 32'h426f48f6, 32'h4182652f, 32'hc2128591};
test_weights[19952:19959] = '{32'h42ba1076, 32'h425f196c, 32'hc2ab367a, 32'h42b93497, 32'hc2ba4e23, 32'hc2165092, 32'hc2a1b431, 32'hc260a69b};
test_bias[2494:2494] = '{32'hc250ae9b};
test_output[2494:2494] = '{32'h4580f660};
test_input[19960:19967] = '{32'hc1f54749, 32'hc20725b8, 32'h428bbf87, 32'h41e5ad59, 32'hc23324c9, 32'hc2099a4f, 32'h405e8d0d, 32'h4140b850};
test_weights[19960:19967] = '{32'hc218d9e8, 32'hc2611afa, 32'hc03221c1, 32'hc24e4a44, 32'hc2942ed4, 32'hc22d12f7, 32'hc18227ac, 32'hc249ad67};
test_bias[2495:2495] = '{32'h4208ed66};
test_output[2495:2495] = '{32'h45ae37b8};
test_input[19968:19975] = '{32'h41d8e7d3, 32'h426a28d5, 32'hc24d8efc, 32'hc2c3025e, 32'hc2200a49, 32'hc287973a, 32'h4275382f, 32'h4295437b};
test_weights[19968:19975] = '{32'h41a0c7cf, 32'hc2382922, 32'h42410e26, 32'h421d11d8, 32'h42862372, 32'h423ddbb0, 32'hc22bfb64, 32'hc258487b};
test_bias[2496:2496] = '{32'h4271b4a4};
test_output[2496:2496] = '{32'hc6a3d6d5};
test_input[19976:19983] = '{32'hc286a659, 32'hc09add40, 32'h4246e8f8, 32'h4272ea26, 32'h41e65f31, 32'h429ea439, 32'h42615c24, 32'hc1f25b5f};
test_weights[19976:19983] = '{32'h422b1ef4, 32'hc1338d7e, 32'hc04bb66b, 32'hc29b8d93, 32'hc26f33cf, 32'hc219dd83, 32'h42be088c, 32'hc185b0fc};
test_bias[2497:2497] = '{32'hc22c7df4};
test_output[2497:2497] = '{32'hc5d04207};
test_input[19984:19991] = '{32'hc285d027, 32'h41c513c6, 32'h417f73d3, 32'h42bdb59b, 32'h40a3252f, 32'h42a5cec2, 32'h422e5080, 32'hc22ec238};
test_weights[19984:19991] = '{32'h4204e9d5, 32'h41ebbb46, 32'h426f08d3, 32'h42a4372a, 32'hc0261268, 32'hc21e350a, 32'h4132ed50, 32'h42b173b6};
test_bias[2498:2498] = '{32'h4261210e};
test_output[2498:2498] = '{32'h441b056e};
test_input[19992:19999] = '{32'h4208cb27, 32'h4294d477, 32'hc2907466, 32'h3fc872fb, 32'h406f293a, 32'hbfdfe35a, 32'h422cf8aa, 32'h416f35f2};
test_weights[19992:19999] = '{32'h42bc2215, 32'h4117066e, 32'hc1bc4967, 32'h421fc736, 32'h41b59bd0, 32'hc2c377ee, 32'h42b0d78d, 32'hc20e27c5};
test_bias[2499:2499] = '{32'hc29f77de};
test_output[2499:2499] = '{32'h460ef870};
test_input[20000:20007] = '{32'hc2bcab2b, 32'h4285aebe, 32'hc201abfd, 32'h41d57afa, 32'h420ce1a6, 32'h3f63f6d0, 32'h4260a444, 32'hc2c0ff85};
test_weights[20000:20007] = '{32'hc238db0a, 32'h4125ffd7, 32'hc26ee705, 32'h423a350c, 32'h4254d714, 32'hc240afb3, 32'hc2c0b1c0, 32'hc11b40d5};
test_bias[2500:2500] = '{32'hc25b5835};
test_output[2500:2500] = '{32'h45acea18};
test_input[20008:20015] = '{32'hc28717a7, 32'hc28b1051, 32'h42083069, 32'h40fac8f6, 32'hc207b3d3, 32'hc2b9e508, 32'h42b2ed4f, 32'hc27e6fa0};
test_weights[20008:20015] = '{32'h42993593, 32'h416a7b5c, 32'h428e3f89, 32'h42b708ee, 32'h411cc129, 32'h4256741c, 32'h4224af2a, 32'h42331d64};
test_bias[2501:2501] = '{32'hc236a870};
test_output[2501:2501] = '{32'hc5ece69b};
test_input[20016:20023] = '{32'h41430426, 32'hc24e1b94, 32'hbf9c764f, 32'h416ddfaf, 32'hc2b04e6b, 32'h4260f730, 32'h4251cdb3, 32'h4271db35};
test_weights[20016:20023] = '{32'hc2609d62, 32'hc221efd7, 32'h429881ca, 32'hc29608b8, 32'hc28b8195, 32'h428c9178, 32'h41df3a3d, 32'hc2a0ce46};
test_bias[2502:2502] = '{32'h4268fcec};
test_output[2502:2502] = '{32'h45d95a0b};
test_input[20024:20031] = '{32'hc25b8095, 32'hc1899dd0, 32'h41f558d7, 32'hc291419b, 32'h420c44e6, 32'hc2be346b, 32'h42846b2a, 32'hc1889a67};
test_weights[20024:20031] = '{32'h42911821, 32'hc21be1d3, 32'hc273cea1, 32'hc29cb2a1, 32'hc2808cba, 32'h4296fe79, 32'h410e69a2, 32'h42811223};
test_bias[2503:2503] = '{32'h42875fe4};
test_output[2503:2503] = '{32'hc6126207};
test_input[20032:20039] = '{32'h4116b314, 32'h4209d3c5, 32'h42c0d788, 32'hc28e7587, 32'hc2044854, 32'h411cdbd3, 32'hc1dece0c, 32'h419575f3};
test_weights[20032:20039] = '{32'h42a6b5be, 32'h4227cd90, 32'h41732cb2, 32'h42524006, 32'hc24bc460, 32'h42066105, 32'hc2430306, 32'hc268d5b0};
test_bias[2504:2504] = '{32'hc2a8b383};
test_output[2504:2504] = '{32'h4506803c};
test_input[20040:20047] = '{32'hc161fca5, 32'hc2a51354, 32'hc2a6ccd1, 32'hbe8df936, 32'h42453d45, 32'h42a11f21, 32'h426fa6ed, 32'hc2c3cd16};
test_weights[20040:20047] = '{32'h42b7ce9c, 32'h42a6b87c, 32'hc234522f, 32'hc2a3acfd, 32'h42c3d422, 32'h3eb80fee, 32'hc23a0e70, 32'hc137fcc5};
test_bias[2505:2505] = '{32'h4240c246};
test_output[2505:2505] = '{32'hc48ff8ed};
test_input[20048:20055] = '{32'h403ec492, 32'h42786aac, 32'h42916802, 32'hc22c85e0, 32'hc285ba53, 32'hc210d6a0, 32'hc2ae6368, 32'h40084b5b};
test_weights[20048:20055] = '{32'hc296a8f5, 32'hc2240a58, 32'hc2a8ac2e, 32'h4255aea1, 32'h4270c823, 32'h421a0861, 32'h42458d63, 32'hc188e75c};
test_bias[2506:2506] = '{32'h4274a530};
test_output[2506:2506] = '{32'hc6a357d7};
test_input[20056:20063] = '{32'h4295a2ca, 32'hc23620cc, 32'h42ab4202, 32'h421c323a, 32'h4152ccb1, 32'h42afbaf1, 32'hc2a3e54b, 32'h4181d221};
test_weights[20056:20063] = '{32'hc20cb5eb, 32'hc287113d, 32'h42778176, 32'hc269e6ac, 32'hc28fdb4f, 32'hc2c1cffb, 32'h42c4528c, 32'h42900f9a};
test_bias[2507:2507] = '{32'hc2c13085};
test_output[2507:2507] = '{32'hc64ac071};
test_input[20064:20071] = '{32'hc095e219, 32'h42710e86, 32'hc1cf8abd, 32'h41e81816, 32'hc17ed091, 32'h42bece03, 32'h41dca7ac, 32'hc2c7c991};
test_weights[20064:20071] = '{32'h42a5968c, 32'hc2060837, 32'h427d2551, 32'hc1633907, 32'hc2561b54, 32'h42a0e2f1, 32'hc19b6133, 32'hc299d6d2};
test_bias[2508:2508] = '{32'h4275939c};
test_output[2508:2508] = '{32'h46302dc5};
test_input[20072:20079] = '{32'h4215e107, 32'hc292228e, 32'h422cc151, 32'h4276915d, 32'h4284ea14, 32'hbf7f30b6, 32'h4270e89c, 32'hc2620cd6};
test_weights[20072:20079] = '{32'h417ef91e, 32'h42886dff, 32'hc2477750, 32'h42045a54, 32'h42009db2, 32'h42b881aa, 32'hc286ebb5, 32'hc08e009d};
test_bias[2509:2509] = '{32'h42a6cb16};
test_output[2509:2509] = '{32'hc5c148c4};
test_input[20080:20087] = '{32'hc261c4bc, 32'hc2478498, 32'h421bd2f1, 32'hc1c84158, 32'hc2c3abb9, 32'h4226ef9f, 32'h40f4bf75, 32'hc2025360};
test_weights[20080:20087] = '{32'hc15fa414, 32'h4276b883, 32'h42acb49c, 32'hc192f9a1, 32'hc29ed4f6, 32'h423bc15c, 32'hc2a23ee0, 32'h41849122};
test_bias[2510:2510] = '{32'hc14283ec};
test_output[2510:2510] = '{32'h461db13a};
test_input[20088:20095] = '{32'hc1fc4d5a, 32'hc191ab01, 32'h41b1ab1b, 32'h42970fd0, 32'hc2b8502b, 32'h42c3b9ba, 32'h42865073, 32'hc207380d};
test_weights[20088:20095] = '{32'hc297facf, 32'hc11997b6, 32'hc0f9d447, 32'hc2440231, 32'hc2acf3fc, 32'hc2bef2b5, 32'h42986db0, 32'hc19087ef};
test_bias[2511:2511] = '{32'hc282ed52};
test_output[2511:2511] = '{32'h453aa687};
test_input[20096:20103] = '{32'h42423920, 32'h4290f9b5, 32'h41d4e5d9, 32'hc193ccf2, 32'hc16aec66, 32'h42474df6, 32'h42ac77af, 32'h429f0718};
test_weights[20096:20103] = '{32'h418f1263, 32'hc21d5bba, 32'hc2b5b194, 32'h4164d8b2, 32'hc2b819e3, 32'hc28500c9, 32'hc202bb8a, 32'hc2917cb5};
test_bias[2512:2512] = '{32'h41f1f5f7};
test_output[2512:2512] = '{32'hc66d7d83};
test_input[20104:20111] = '{32'h41fa84a9, 32'h40c3b415, 32'h424522d6, 32'h428361b4, 32'hc25430e6, 32'hc12277f7, 32'h42186387, 32'hc28e0945};
test_weights[20104:20111] = '{32'h4290494b, 32'h42649296, 32'hc2876176, 32'hc22fb3b8, 32'hc1cb61e6, 32'h407a0849, 32'h428474b6, 32'hc2504961};
test_bias[2513:2513] = '{32'hc2b95a47};
test_output[2513:2513] = '{32'h456f0781};
test_input[20112:20119] = '{32'hc2691796, 32'hc1edd771, 32'h41f47ed9, 32'h3fe2115b, 32'hc1db1049, 32'h42a5c737, 32'h428c4dea, 32'h42a6bc81};
test_weights[20112:20119] = '{32'hc1eeea46, 32'hbf61e351, 32'h417e20b1, 32'h423f3989, 32'hc2018245, 32'hc0271e27, 32'h42a9af17, 32'h405d2220};
test_bias[2514:2514] = '{32'hc2c7271e};
test_output[2514:2514] = '{32'h460eeb5b};
test_input[20120:20127] = '{32'h40d22520, 32'hc1c6726f, 32'hc276a679, 32'h4225380d, 32'hc2a29e6f, 32'h428b0423, 32'hc2ac77f3, 32'h4202944a};
test_weights[20120:20127] = '{32'h42b3cb08, 32'h42bdae34, 32'h428c555a, 32'hc06a67b9, 32'hc235d1bb, 32'hc2b13cbd, 32'hc2797748, 32'h42113303};
test_bias[2515:2515] = '{32'hc227feee};
test_output[2515:2515] = '{32'hc5086dbc};
test_input[20128:20135] = '{32'hc27af30b, 32'h42084ed2, 32'hc1dae999, 32'hc29ddc3c, 32'hc18089ff, 32'h4229bfb8, 32'hc13a33f4, 32'h4211e8f5};
test_weights[20128:20135] = '{32'h42832379, 32'h41314352, 32'hc2a5ab51, 32'hc2b4a9d4, 32'h4215075b, 32'hc2362bcd, 32'hc1972bb9, 32'h41bf99de};
test_bias[2516:2516] = '{32'h4244a5df};
test_output[2516:2516] = '{32'h45857eda};
test_input[20136:20143] = '{32'hc2644189, 32'h42b8e700, 32'h4286245e, 32'h41e266cd, 32'h4224b303, 32'h42bac06b, 32'h42611b74, 32'h41b0934a};
test_weights[20136:20143] = '{32'hc2505dc0, 32'h42bedc44, 32'h42c72baa, 32'h42047688, 32'hc284bcc1, 32'h41248d8f, 32'hc2b048c9, 32'h425f9049};
test_bias[2517:2517] = '{32'hc2a8be7f};
test_output[2517:2517] = '{32'h465810a0};
test_input[20144:20151] = '{32'hc29e4e4d, 32'h429d8b17, 32'hc1c63fe6, 32'hc1ac5a52, 32'h42817a50, 32'hc18d0462, 32'h41e57f1c, 32'h42a25be0};
test_weights[20144:20151] = '{32'h41f8650c, 32'hc0ecd3e2, 32'h425a5e85, 32'hc24d0c80, 32'hc22bb678, 32'h413bbb2c, 32'h42479520, 32'h425f8823};
test_bias[2518:2518] = '{32'hc1ad4cd1};
test_output[2518:2518] = '{32'hc3a4656e};
test_input[20152:20159] = '{32'hc21ad6d5, 32'h418cb64c, 32'h41dba179, 32'h41c0ed36, 32'h41ef4805, 32'h4232b137, 32'hc23926d8, 32'h419e2c27};
test_weights[20152:20159] = '{32'hc104e71f, 32'hc1f4bb67, 32'hc20d672d, 32'h4259c571, 32'hbfebe24d, 32'h41647166, 32'h4293b644, 32'h422d2232};
test_bias[2519:2519] = '{32'hc1e65a65};
test_output[2519:2519] = '{32'hc4eb61fd};
test_input[20160:20167] = '{32'hc281d4a1, 32'h42456787, 32'h421eb9b5, 32'hc2a092fb, 32'hc2a6915e, 32'h429ef2b4, 32'h4234d25e, 32'hc29dac33};
test_weights[20160:20167] = '{32'h42082b23, 32'hc2163c2a, 32'hc2b2848a, 32'h4264bb63, 32'h42aa99c4, 32'hc2aac984, 32'h4292df6a, 32'hc219a46b};
test_bias[2520:2520] = '{32'hc2c67a1c};
test_output[2520:2520] = '{32'hc69afcf2};
test_input[20168:20175] = '{32'h42671422, 32'hc2bd88bb, 32'hc0acd1ee, 32'h4253e268, 32'hc290cbac, 32'h4160685c, 32'hc28bd651, 32'hc2bb7ce8};
test_weights[20168:20175] = '{32'hc28cbb1a, 32'hc221f382, 32'hc2526e14, 32'hc20f6fcf, 32'hc20e8c88, 32'hc2bdeca7, 32'h42c494bc, 32'h42888667};
test_bias[2521:2521] = '{32'hc2c777ce};
test_output[2521:2521] = '{32'hc65a3a3f};
test_input[20176:20183] = '{32'hc210b0b8, 32'hc22e22eb, 32'hbf1f3ee6, 32'hc29ee24d, 32'h4297099d, 32'hc14e7b85, 32'hc2842b3a, 32'h42ac827c};
test_weights[20176:20183] = '{32'hbe2d72e3, 32'hc2c664fd, 32'h42736a70, 32'hc1f8b809, 32'hc2afa6b3, 32'h41db807c, 32'h42a76c28, 32'hc255ea6d};
test_bias[2522:2522] = '{32'h42960b2a};
test_output[2522:2522] = '{32'hc620ef31};
test_input[20184:20191] = '{32'h4189ce36, 32'h4250a8e5, 32'hc1fa3209, 32'hc2436efd, 32'h419249fd, 32'h4228ff7e, 32'h428d98b3, 32'h429baf24};
test_weights[20184:20191] = '{32'h428994fe, 32'hc1dcc372, 32'h419aa157, 32'h42ada088, 32'hc2b8b48b, 32'hc27db54b, 32'hc2b062db, 32'hc29b1c6e};
test_bias[2523:2523] = '{32'hc2b5648e};
test_output[2523:2523] = '{32'hc6aaa1ab};
test_input[20192:20199] = '{32'h4245695d, 32'h42a13c68, 32'h41b410f4, 32'hc207ec6f, 32'hc2a073fe, 32'h428a5a89, 32'h42bc4461, 32'h4277a42f};
test_weights[20192:20199] = '{32'hc2343c03, 32'hc0ee16cd, 32'h422892b3, 32'h4249c7ff, 32'hc29fd33b, 32'h421caace, 32'h4241ab71, 32'hc2139821};
test_bias[2524:2524] = '{32'h429a2b5b};
test_output[2524:2524] = '{32'h45f64ddd};
test_input[20200:20207] = '{32'hc2b88925, 32'h424bd0e5, 32'h41b01725, 32'h42366ade, 32'h42aa4c27, 32'h425a753b, 32'h422ed3fe, 32'h426c2ab5};
test_weights[20200:20207] = '{32'h429493af, 32'hc292fd51, 32'h4244473f, 32'hc2659ab1, 32'h423c0875, 32'h428afb0a, 32'h41daf2bf, 32'hc2bac190};
test_bias[2525:2525] = '{32'h41e1e5e6};
test_output[2525:2525] = '{32'hc606cf58};
test_input[20208:20215] = '{32'hc29ece02, 32'hc20ecf0b, 32'h42bed6b5, 32'h42882d72, 32'h4275e4b8, 32'h404cc947, 32'hc169978d, 32'hc18c55f7};
test_weights[20208:20215] = '{32'h429cbc6e, 32'hc296d2d9, 32'hc2af43b2, 32'h4231b9bf, 32'hc2b65ce6, 32'h42902135, 32'hc2a86b7a, 32'h4285701c};
test_bias[2526:2526] = '{32'hc20516ec};
test_output[2526:2526] = '{32'hc65e1e8e};
test_input[20216:20223] = '{32'hc00ca756, 32'h41d9c642, 32'h415167db, 32'hc2878bd3, 32'hc23fd0fd, 32'h40f916ea, 32'h41859cc8, 32'hc1dd5569};
test_weights[20216:20223] = '{32'h41cf2202, 32'h41d1f39e, 32'hc2088a85, 32'hc25f60d7, 32'hc276c86a, 32'hc279ee64, 32'h42574341, 32'h420de8f8};
test_bias[2527:2527] = '{32'hc28b3ed7};
test_output[2527:2527] = '{32'h45c55ab3};
test_input[20224:20231] = '{32'hc253d133, 32'hc15f6472, 32'hc14c8572, 32'h3e256ac6, 32'h42a996fc, 32'h4284d3ef, 32'hc086c8cc, 32'h42ab1ccd};
test_weights[20224:20231] = '{32'h42b6b3a4, 32'h41adda7c, 32'hc2332114, 32'h42465c2b, 32'h42b38f89, 32'h429d40ad, 32'h4190d81e, 32'h42bec6d1};
test_bias[2528:2528] = '{32'hc1eb32de};
test_output[2528:2528] = '{32'h467f273c};
test_input[20232:20239] = '{32'hc2afe0b1, 32'hc28e5b5c, 32'h4059d4f6, 32'hc2a6dd72, 32'h42a4e4c8, 32'h428a8640, 32'hc269c74f, 32'hc10c4882};
test_weights[20232:20239] = '{32'h42078f5b, 32'hc2805465, 32'h41fbe921, 32'hc29ea5b5, 32'hc1c64b5d, 32'h41b4e4f8, 32'h42b1ec8e, 32'hc0fad1dd};
test_bias[2529:2529] = '{32'hc25a8b2e};
test_output[2529:2529] = '{32'h45259893};
test_input[20240:20247] = '{32'h40aa8326, 32'hc2531def, 32'h429d58ca, 32'h429aa527, 32'h4222ff12, 32'hc2c48e1b, 32'h429b20ec, 32'h428b04d9};
test_weights[20240:20247] = '{32'hc258fb8d, 32'h40e3109f, 32'hc2b4adfa, 32'h425317a8, 32'h41e047a7, 32'h41d2c84f, 32'hc2ba920f, 32'h427ac6f6};
test_bias[2530:2530] = '{32'h42af408b};
test_output[2530:2530] = '{32'hc5f7bbd3};
test_input[20248:20255] = '{32'h42476602, 32'h42aa1e05, 32'h416793b7, 32'hc2356242, 32'h4216725c, 32'h40ebd791, 32'hc2be0d07, 32'hc2129b1a};
test_weights[20248:20255] = '{32'h4181b641, 32'hc0e7d5ed, 32'hc243a1a2, 32'h41327e7a, 32'h42c7cffa, 32'h429d1539, 32'hc2203332, 32'h429563a4};
test_bias[2531:2531] = '{32'h42935f44};
test_output[2531:2531] = '{32'h458b447e};
test_input[20256:20263] = '{32'h41ac26dc, 32'h426f8af2, 32'hc2c0148c, 32'hc2bb4392, 32'hc2590d05, 32'hc25a3eea, 32'h4114e148, 32'hc0d6e7ab};
test_weights[20256:20263] = '{32'h42450d08, 32'h429c2fd6, 32'h42553c0f, 32'h42628d63, 32'hc10108da, 32'hc26213fa, 32'hc119be4d, 32'h421e383a};
test_bias[2532:2532] = '{32'h425ee2d6};
test_output[2532:2532] = '{32'hc4b70283};
test_input[20264:20271] = '{32'hc2064d55, 32'h4216fbf4, 32'hc2121571, 32'hc0948371, 32'h415aa110, 32'hc2abd20a, 32'h4293136e, 32'h42c3a036};
test_weights[20264:20271] = '{32'hc1e420b9, 32'hc28fd553, 32'h42653109, 32'h428769f1, 32'h40d51fa2, 32'h42845fdf, 32'h429310fa, 32'h410c1d4d};
test_bias[2533:2533] = '{32'hc29810c8};
test_output[2533:2533] = '{32'hc55f3151};
test_input[20272:20279] = '{32'h41d96615, 32'hc2030146, 32'hc2bc0adb, 32'h420a08ee, 32'hc12284ec, 32'h4265b389, 32'h411974db, 32'hc298df33};
test_weights[20272:20279] = '{32'hc289499d, 32'h42122c98, 32'hc2beb77c, 32'h42bc6126, 32'hc04a6099, 32'hc29752f5, 32'hc19419cd, 32'h424a40fe};
test_bias[2534:2534] = '{32'h4187657c};
test_output[2534:2534] = '{32'h444be350};
test_input[20280:20287] = '{32'hc0a3ab35, 32'h429169bf, 32'hc2b103d8, 32'h41b35398, 32'hc2180983, 32'h42174780, 32'hc1c7eb6a, 32'h3ef6d390};
test_weights[20280:20287] = '{32'hc2913975, 32'h4298b4e9, 32'hc2988f9c, 32'hc23be6b9, 32'hc0eaad33, 32'h42c0c154, 32'h42b9bc79, 32'h40e0af77};
test_bias[2535:2535] = '{32'h4290495a};
test_output[2535:2535] = '{32'h464fceac};
test_input[20288:20295] = '{32'hc2a73e46, 32'hc2a398af, 32'hc29bf280, 32'hc29aaf6f, 32'h41d0f60b, 32'h42b593e7, 32'hc2917b2f, 32'hc2b12655};
test_weights[20288:20295] = '{32'h426f48e1, 32'hc1b88718, 32'h429fd0a4, 32'hc2b33e39, 32'h4292fd56, 32'h41fda88d, 32'hc2c5cdbb, 32'hc2a0c6ce};
test_bias[2536:2536] = '{32'hc2a25212};
test_output[2536:2536] = '{32'h4681d21f};
test_input[20296:20303] = '{32'h4239e505, 32'h427754c4, 32'h4271bceb, 32'hc287cd8b, 32'hc23cc884, 32'hc255521d, 32'hc29bd8a3, 32'h42a27039};
test_weights[20296:20303] = '{32'h42a7744d, 32'h4159fea0, 32'h41d335e3, 32'hc2c2b113, 32'h4242b273, 32'h4110688c, 32'hc2117715, 32'hc292c130};
test_bias[2537:2537] = '{32'h41b019f0};
test_output[2537:2537] = '{32'h45dc84f2};
test_input[20304:20311] = '{32'hc2a2567b, 32'hc29b061b, 32'h41d43d7c, 32'h421d1ab1, 32'h423cfb24, 32'hc0e253c1, 32'hc1a80c6d, 32'h41f61684};
test_weights[20304:20311] = '{32'h4226cda6, 32'hc2c2f40e, 32'h42c7ff8f, 32'h4215db27, 32'h422d2c38, 32'h418af73b, 32'h42357fd2, 32'h42963c8c};
test_bias[2538:2538] = '{32'hc2163dfe};
test_output[2538:2538] = '{32'h46344707};
test_input[20312:20319] = '{32'hc28c627b, 32'hc1c04957, 32'h4287b6ca, 32'hc14e471a, 32'hc1ae56de, 32'h418838a7, 32'h423c08f9, 32'hc2516e34};
test_weights[20312:20319] = '{32'h427cd8f1, 32'hc29cb462, 32'hc2c71c5b, 32'h413e26b6, 32'hc2c74095, 32'h42a7e451, 32'h42a4ec3f, 32'hc259d9a4};
test_bias[2539:2539] = '{32'h4203f5e1};
test_output[2539:2539] = '{32'h4460bcc2};
test_input[20320:20327] = '{32'hc294356d, 32'h42a5947e, 32'hc1e2e90b, 32'hc2010ed5, 32'hc2822ec3, 32'h42672963, 32'h4188fb11, 32'hc2aacf27};
test_weights[20320:20327] = '{32'h4289abce, 32'h4276f239, 32'hc29f7d26, 32'hc2a0d2ed, 32'hc039d6d7, 32'h42bbee9b, 32'h422e9843, 32'h42b851af};
test_bias[2540:2540] = '{32'hc28c5942};
test_output[2540:2540] = '{32'h454dc295};
test_input[20328:20335] = '{32'h41b1a362, 32'h42777adc, 32'h4181a7ed, 32'hc0eeacfe, 32'hc2c70ab5, 32'hc252957e, 32'hc22d0abd, 32'h4252b290};
test_weights[20328:20335] = '{32'hc2c03a6e, 32'h4184513d, 32'hc2b1baa4, 32'h42046e39, 32'hc1b6730d, 32'hc25e76e9, 32'h42008e6c, 32'hc2b3dcbf};
test_bias[2541:2541] = '{32'hc0c4a8c1};
test_output[2541:2541] = '{32'hc5695f4a};
test_input[20336:20343] = '{32'hc2b9faca, 32'hc2bf2743, 32'h3fcfff32, 32'h4275748c, 32'h425d1e8d, 32'h41cf6889, 32'h3f922cbe, 32'h42b488e0};
test_weights[20336:20343] = '{32'h42ad7477, 32'h42779715, 32'h42447373, 32'hc2849424, 32'h4258a62a, 32'h40ac1af9, 32'h4280d641, 32'h41f2b560};
test_bias[2542:2542] = '{32'hc28460e2};
test_output[2542:2542] = '{32'hc63ce4de};
test_input[20344:20351] = '{32'h42b26473, 32'h4118ad12, 32'h428fec40, 32'h41e4c275, 32'hc2003553, 32'h42208c74, 32'h427435d4, 32'hc2080fe4};
test_weights[20344:20351] = '{32'h41268a23, 32'hc2620abc, 32'h42312dc4, 32'h41b26e78, 32'hc1f28648, 32'hc28aea58, 32'hc1c692b8, 32'hc1cc422c};
test_bias[2543:2543] = '{32'h429a3d67};
test_output[2543:2543] = '{32'h44e49013};
test_input[20352:20359] = '{32'h427f1e17, 32'hc18a8a36, 32'h426388a6, 32'hc28421f2, 32'h42388b4c, 32'hc2623233, 32'hc27e021c, 32'hc2b24ed9};
test_weights[20352:20359] = '{32'h424294f7, 32'hc130e1a5, 32'h423a97c2, 32'hc086e4ce, 32'h424c32ef, 32'h42bb0362, 32'hc114f5c7, 32'h41f23747};
test_bias[2544:2544] = '{32'hc217d403};
test_output[2544:2544] = '{32'h448f6fb3};
test_input[20360:20367] = '{32'hc282be80, 32'hc2852bff, 32'h42bf6d2a, 32'hc2396f19, 32'hc17a4e5a, 32'hc26b51cf, 32'hc2b39512, 32'h428a46cb};
test_weights[20360:20367] = '{32'h42700c9a, 32'h4239a4fb, 32'hc241daf9, 32'hc2beebc2, 32'h42b87462, 32'h42823e00, 32'h41db73bc, 32'hc211cbb6};
test_bias[2545:2545] = '{32'h3f8bb78f};
test_output[2545:2545] = '{32'hc6889532};
test_input[20368:20375] = '{32'h41298993, 32'h42b40347, 32'hc274000d, 32'hc2aa9335, 32'h41585e35, 32'h42057379, 32'hc2b20844, 32'h420bab1e};
test_weights[20368:20375] = '{32'h41cd448b, 32'h41f7d01a, 32'h4281c280, 32'hc2be0a24, 32'hc0886068, 32'h418abc3d, 32'h421ab3b7, 32'hc20225d2};
test_bias[2546:2546] = '{32'hc29ad2f3};
test_output[2546:2546] = '{32'h453fefd7};
test_input[20376:20383] = '{32'h4115effc, 32'h409e55fd, 32'hc27ede1d, 32'h41a86bd8, 32'h424d0a0e, 32'hc29cb866, 32'hc2a30bf4, 32'hc1e9f905};
test_weights[20376:20383] = '{32'h41091dcd, 32'hc2bc176d, 32'h421c09c0, 32'hc24d4614, 32'hc1c4a07e, 32'h41a206cc, 32'h42c7975b, 32'hc1ccaeb6};
test_bias[2547:2547] = '{32'h42b87252};
test_output[2547:2547] = '{32'hc65c3459};
test_input[20384:20391] = '{32'h42c694cf, 32'hc2b4e396, 32'h41b54379, 32'hc2791322, 32'h4281b08f, 32'hc149c9d2, 32'h42413582, 32'hc2a2fe8d};
test_weights[20384:20391] = '{32'h41bb0946, 32'h41fbe23e, 32'h423c49d1, 32'hc2c1a492, 32'h42a374b2, 32'hc29e1ad0, 32'h424740b3, 32'h427ad4a6};
test_bias[2548:2548] = '{32'hc2bf09e0};
test_output[2548:2548] = '{32'h461d4783};
test_input[20392:20399] = '{32'hc2a6f9b8, 32'hc29ce095, 32'hc20fa417, 32'hc1034388, 32'hc23b00ac, 32'hc244586b, 32'h42aa8614, 32'hc27bcc49};
test_weights[20392:20399] = '{32'h429f1087, 32'h42235cfb, 32'h42c71603, 32'h4296ac94, 32'hc1fb44de, 32'hc27fcb64, 32'h4293c8fd, 32'hc25cbcd6};
test_bias[2549:2549] = '{32'h4206c560};
test_output[2549:2549] = '{32'h43bd7ccb};
test_input[20400:20407] = '{32'h42b2e95c, 32'hc266ec17, 32'hc2b76762, 32'h41225527, 32'hc25a940f, 32'hc2bd3efa, 32'h41741a1d, 32'h3f90bb52};
test_weights[20400:20407] = '{32'hc2038666, 32'h42ae1083, 32'h42978e91, 32'hc2b493b5, 32'hc2695687, 32'h428642b5, 32'h4232f327, 32'h42a17cc8};
test_bias[2550:2550] = '{32'h4290cb27};
test_output[2550:2550] = '{32'hc68dca30};
test_input[20408:20415] = '{32'h425040cd, 32'hc20dc7a1, 32'hc2a737d0, 32'h4189d3d8, 32'hc1a1ee33, 32'hc2a1cd42, 32'hc218c0b0, 32'hc28665fb};
test_weights[20408:20415] = '{32'hc299ff3c, 32'hc270df38, 32'hc1af8a71, 32'h41cdf008, 32'h41047848, 32'hc2930869, 32'hc196d10e, 32'h414f694b};
test_bias[2551:2551] = '{32'hc22c502a};
test_output[2551:2551] = '{32'h45bb2b54};
test_input[20416:20423] = '{32'hc24402ee, 32'hc20749ee, 32'h41917eef, 32'h42a92784, 32'h42af4388, 32'h429e6f40, 32'h4254e703, 32'h40d4d978};
test_weights[20416:20423] = '{32'hc2118f93, 32'h40f75431, 32'hc286e491, 32'hc262b681, 32'hc277762e, 32'h41bcb249, 32'hc1d6d862, 32'hc2429133};
test_bias[2552:2552] = '{32'h425cdea1};
test_output[2552:2552] = '{32'hc618548a};
test_input[20424:20431] = '{32'h42bf7b83, 32'h42ad5c3d, 32'hc240e25d, 32'h4288d3ba, 32'h40a89a79, 32'h42872c22, 32'hc121b559, 32'hc0755596};
test_weights[20424:20431] = '{32'hc218b01a, 32'h4264a2cf, 32'h41f34a8c, 32'h42856025, 32'h422c1fc3, 32'hc297f8c4, 32'hc1f9c9b9, 32'hc2bffc76};
test_bias[2553:2553] = '{32'h42c34adf};
test_output[2553:2553] = '{32'h43860e86};
test_input[20432:20439] = '{32'hc15cd4a5, 32'hc24a8ec8, 32'hc254f51a, 32'hc264be7c, 32'h40e5f502, 32'h424b06f2, 32'hc215d50b, 32'h42a5671c};
test_weights[20432:20439] = '{32'hc1d767fd, 32'hc2c29d30, 32'h4229eba6, 32'hc2821b8b, 32'hc26e3bff, 32'hc23cd1ef, 32'hc23e1ef7, 32'hc29e7167};
test_bias[2554:2554] = '{32'h42873c80};
test_output[2554:2554] = '{32'hc4407c1b};
test_input[20440:20447] = '{32'hc27463dc, 32'h428eff39, 32'hc2091438, 32'hc1645a23, 32'hc1bea02e, 32'h429fce3a, 32'h41ad6af4, 32'hc2b3c806};
test_weights[20440:20447] = '{32'hc0e65b35, 32'h42630fb9, 32'h42a11878, 32'hc1df865c, 32'hc288e1e0, 32'h41af373c, 32'hc205aa52, 32'hc2189adb};
test_bias[2555:2555] = '{32'hc18d4975};
test_output[2555:2555] = '{32'h4600348c};
test_input[20448:20455] = '{32'h41bd58dc, 32'hc18f84ad, 32'h428cdb10, 32'h42912e0e, 32'h411dd360, 32'h41002a5c, 32'h41ef9fd6, 32'h42a46ec1};
test_weights[20448:20455] = '{32'h4228d6d4, 32'h428c9fee, 32'hc153eccf, 32'h42aa25ed, 32'hc28ba3a1, 32'hc2882b71, 32'h4112639a, 32'h42b8db53};
test_bias[2556:2556] = '{32'h42839010};
test_output[2556:2556] = '{32'h463694c6};
test_input[20456:20463] = '{32'h42696b75, 32'h429f61df, 32'hc276b630, 32'hc2819e3f, 32'hc2815841, 32'hc288ab91, 32'hc098f17d, 32'hc2c07b15};
test_weights[20456:20463] = '{32'hc1cdec75, 32'h4223e3e4, 32'hc18af4de, 32'h40c358b2, 32'h41ecbf75, 32'hc1b03877, 32'h422a453a, 32'h425e6d2f};
test_bias[2557:2557] = '{32'h427866ec};
test_output[2557:2557] = '{32'hc5586d34};
test_input[20464:20471] = '{32'h425bbe3e, 32'hbef2b4bb, 32'h41bd8718, 32'hc0e265d4, 32'h422e2b8f, 32'h42b0b3c5, 32'hc29cde36, 32'hc2a999a2};
test_weights[20464:20471] = '{32'h4278a68b, 32'hc29c1e1f, 32'hc1c90bc2, 32'h42a1159f, 32'hc26993ee, 32'h41dd133c, 32'h42c7fee4, 32'hc22f5acc};
test_bias[2558:2558] = '{32'h41a0b482};
test_output[2558:2558] = '{32'hc4efff62};
test_input[20472:20479] = '{32'hc1b275cc, 32'hc227f48b, 32'hc23cfc3d, 32'h42928db0, 32'h420034d5, 32'hbf4958fa, 32'h41a94658, 32'hc257c2f1};
test_weights[20472:20479] = '{32'h411e6a48, 32'h4231b9e8, 32'h425dcf58, 32'hc281c8e5, 32'hc2a48049, 32'h4290a569, 32'h42a71149, 32'hc280b74f};
test_bias[2559:2559] = '{32'h41130f46};
test_output[2559:2559] = '{32'hc5d7d3ab};
test_input[20480:20487] = '{32'h41ede42b, 32'hc196b7c4, 32'h42846bcc, 32'hc25c652e, 32'h429c3064, 32'h425481dd, 32'h40d080ff, 32'hc2651a04};
test_weights[20480:20487] = '{32'h428ba51e, 32'hc245208f, 32'h427ea0db, 32'h426bbc1d, 32'h4237614a, 32'hc139d6f3, 32'h41e866eb, 32'hc2a043ee};
test_bias[2560:2560] = '{32'h426ab8a9};
test_output[2560:2560] = '{32'h4637f45e};
test_input[20488:20495] = '{32'h4264d779, 32'h42209845, 32'hc257288d, 32'hc25edc18, 32'hc2c1434a, 32'hc26c9e87, 32'h42c38029, 32'hc21784a6};
test_weights[20488:20495] = '{32'hc24ddf78, 32'h41ef1313, 32'h429b650c, 32'hc20f9159, 32'h42160406, 32'hc20b59bb, 32'hc1412391, 32'hc251871d};
test_bias[2561:2561] = '{32'hc166dd1a};
test_output[2561:2561] = '{32'hc592cdd2};
test_input[20496:20503] = '{32'h41661b8c, 32'hc1cf5d3a, 32'hc13dee85, 32'hc2bcab59, 32'hc24840e6, 32'h426db9b9, 32'hc2703fbb, 32'h4246657d};
test_weights[20496:20503] = '{32'h4245037d, 32'hc29b031b, 32'hc24e2f6b, 32'h4292005c, 32'hc20f0032, 32'h421946a2, 32'hc29d7a63, 32'hc2051a78};
test_bias[2562:2562] = '{32'hc2a9fb45};
test_output[2562:2562] = '{32'h455afaaa};
test_input[20504:20511] = '{32'h41084a5f, 32'hc1e89ba2, 32'hc2561668, 32'hc291d667, 32'h42c7c086, 32'h42834a5f, 32'h42a4fdc0, 32'h42b4f871};
test_weights[20504:20511] = '{32'hc1dee149, 32'h420f4f9d, 32'hc186c84d, 32'hc2997d59, 32'hc1ceae52, 32'h41cbe452, 32'hc25a5b8f, 32'hc15f36f0};
test_bias[2563:2563] = '{32'hc2bdbca4};
test_output[2563:2563] = '{32'hc4c1a0eb};
test_input[20512:20519] = '{32'hc1b7025d, 32'hc2804f74, 32'h41fd6d49, 32'hc1fb8997, 32'hc1a14f2a, 32'h42b8c728, 32'h4297dbc6, 32'h41dfeb0c};
test_weights[20512:20519] = '{32'hc2b95070, 32'hc2a88fe3, 32'h42a4d6a4, 32'hc262316c, 32'h427a36a7, 32'h423f2ef8, 32'hc2c343d0, 32'h42195619};
test_bias[2564:2564] = '{32'h4258fa53};
test_output[2564:2564] = '{32'h460940a8};
test_input[20520:20527] = '{32'h42be6b57, 32'h41f9a360, 32'h41f85fed, 32'hc212ea97, 32'hc289fc71, 32'h4223e8ff, 32'hc2c526ce, 32'hc2071b94};
test_weights[20520:20527] = '{32'h403b9782, 32'h42ac73b7, 32'hc16a68e9, 32'h4299e9df, 32'hc23999b2, 32'hc29d2ba0, 32'h42a33974, 32'hc1f4aa4e};
test_bias[2565:2565] = '{32'h42b62bd9};
test_output[2565:2565] = '{32'hc5e29c21};
test_input[20528:20535] = '{32'hc19c0584, 32'h427051bd, 32'h42bd1efa, 32'h41e6fecd, 32'hc26991ae, 32'hc291cee3, 32'h42b2f9b7, 32'hc21ea6f8};
test_weights[20528:20535] = '{32'hc11f903d, 32'hc28e577d, 32'hc28ff07f, 32'h420d5448, 32'h40e366d8, 32'h42231f3a, 32'hc21c5c14, 32'h428fe4f4};
test_bias[2566:2566] = '{32'hc2a7af2e};
test_output[2566:2566] = '{32'hc699d49c};
test_input[20536:20543] = '{32'hc2551181, 32'hc2bbf034, 32'hc281d2bf, 32'hc0eae4ce, 32'h41db0680, 32'hc29e71bf, 32'hc11934d2, 32'hc21b86a0};
test_weights[20536:20543] = '{32'hc2b1d1b5, 32'h42907ec1, 32'h40011c46, 32'h42aaadc3, 32'hc271cc27, 32'hc28eb468, 32'hc2c780bd, 32'h42487b61};
test_bias[2567:2567] = '{32'hc081bb45};
test_output[2567:2567] = '{32'h433d93d5};
test_input[20544:20551] = '{32'h40627b2f, 32'h428d8cb4, 32'hc2b7f8af, 32'h42c1f6e7, 32'h41a65823, 32'hc2bcfa62, 32'hc27f524e, 32'hc1de4010};
test_weights[20544:20551] = '{32'h42a5ec32, 32'hc2471dc6, 32'hc2a6d838, 32'hc2bc99b0, 32'h41014439, 32'h420bc021, 32'hc124f2f2, 32'hc2a034a1};
test_bias[2568:2568] = '{32'hc2a8dcb7};
test_output[2568:2568] = '{32'hc59d5c81};
test_input[20552:20559] = '{32'h42a56dc8, 32'h42bd62e8, 32'hc28ba42d, 32'h42aba94e, 32'h42b55a6f, 32'hc2102a84, 32'h42026914, 32'h4197494b};
test_weights[20552:20559] = '{32'hc29e9f36, 32'hc1745026, 32'h429ad3ef, 32'hc224c52b, 32'hc28957a2, 32'hc28a4237, 32'h42aab66a, 32'hc0a93142};
test_bias[2569:2569] = '{32'h423f6d86};
test_output[2569:2569] = '{32'hc68c3eca};
test_input[20560:20567] = '{32'h41216941, 32'h4238ce90, 32'hc20edd1c, 32'h4222657b, 32'hc28bcf3f, 32'hc284fcd8, 32'h42078562, 32'hc25df3f4};
test_weights[20560:20567] = '{32'h41b1d859, 32'h41cd1ad5, 32'hc117643e, 32'h4203f5fa, 32'h41bba7f4, 32'hc2208c2a, 32'hc1a6f98d, 32'h3fb17a82};
test_bias[2570:2570] = '{32'hc2bb0ac8};
test_output[2570:2570] = '{32'h454a59aa};
test_input[20568:20575] = '{32'h42b69247, 32'h411246d9, 32'hc209ed8e, 32'h424bb3a5, 32'h4291a8d0, 32'h42a181df, 32'h41a16e30, 32'h421bd302};
test_weights[20568:20575] = '{32'h422705a7, 32'h42ad1467, 32'h429aad96, 32'hc1a9f531, 32'hbf8a9a4a, 32'hc22582d4, 32'hc2be9c52, 32'hc1eb847e};
test_bias[2571:2571] = '{32'hc2a04663};
test_output[2571:2571] = '{32'hc5b2a206};
test_input[20576:20583] = '{32'h42a620f2, 32'hc2bb621a, 32'hc076abd2, 32'h429f8e33, 32'h429f0db6, 32'hc22deda0, 32'h4154b89b, 32'hc1c6dd18};
test_weights[20576:20583] = '{32'h41ee0d9f, 32'h4296856e, 32'hc20c5dcc, 32'h415ac9f2, 32'hc2bfbe92, 32'h4210d58d, 32'h426497e1, 32'h41b9369a};
test_bias[2572:2572] = '{32'h42a1bf81};
test_output[2572:2572] = '{32'hc63ffc54};
test_input[20584:20591] = '{32'h424f5f3c, 32'hc26f4023, 32'h420899dd, 32'hc2a8e8ed, 32'h426b3bb3, 32'hc21bd5bc, 32'h41bf83e5, 32'h41c79a89};
test_weights[20584:20591] = '{32'hc27e857a, 32'h4258964d, 32'h40e23379, 32'h41e2f934, 32'hc2c75a04, 32'hc1a89b41, 32'hc2a8cd9e, 32'hc25e7556};
test_bias[2573:2573] = '{32'hc22de4b0};
test_output[2573:2573] = '{32'hc68640ed};
test_input[20592:20599] = '{32'h4296c38e, 32'hc2548713, 32'h429912ca, 32'h4241afc2, 32'h42c5d39c, 32'h3f8a8ed1, 32'h42aaf56d, 32'h414e6e2d};
test_weights[20592:20599] = '{32'hc2553f85, 32'hc2b58082, 32'hc20ce2fb, 32'h4201a446, 32'hc1b9c89c, 32'hc26136d3, 32'h42ba0d89, 32'h428aebee};
test_bias[2574:2574] = '{32'h4147ac57};
test_output[2574:2574] = '{32'h45c118e8};
test_input[20600:20607] = '{32'hc29b67da, 32'h42ace018, 32'h4289986e, 32'hc2692f91, 32'h42024148, 32'h400b1502, 32'hc2959cd1, 32'hc2b6133d};
test_weights[20600:20607] = '{32'h42862b51, 32'h4270aa04, 32'hc14c724b, 32'h40d7bf13, 32'h42bda2ad, 32'hc18b3357, 32'h42c7f396, 32'h42b79fcc};
test_bias[2575:2575] = '{32'hc28ca085};
test_output[2575:2575] = '{32'hc65cf769};
test_input[20608:20615] = '{32'h41c60254, 32'h424d3e75, 32'hc26a9210, 32'h421f6d96, 32'h41dee5c7, 32'hc12f1011, 32'hc11b65e6, 32'hc1922cbd};
test_weights[20608:20615] = '{32'h42afc0df, 32'hc1026513, 32'hc2b20f95, 32'hc21dbcea, 32'h428ae2b1, 32'h40b7df6a, 32'hc256e64d, 32'hc2bdea37};
test_bias[2576:2576] = '{32'h427b1014};
test_output[2576:2576] = '{32'h4615f6c0};
test_input[20616:20623] = '{32'hc225f31c, 32'hc142032e, 32'h424e3375, 32'h4280d078, 32'hc19b7f8c, 32'h4135f39a, 32'h425f8a51, 32'h42728fe7};
test_weights[20616:20623] = '{32'hc185a0fd, 32'hc292b2c2, 32'hc118ea6b, 32'hc283753e, 32'hc233d29b, 32'h42bf4754, 32'h426c40bd, 32'h40896180};
test_bias[2577:2577] = '{32'hc2859124};
test_output[2577:2577] = '{32'h451080a6};
test_input[20624:20631] = '{32'h405984a3, 32'hc2b1544c, 32'h41b64d05, 32'hc2458e5c, 32'h41a99d84, 32'hc1d2d3a2, 32'h42af8ef4, 32'hc2aded0e};
test_weights[20624:20631] = '{32'hc2b1fea9, 32'hc2093fe2, 32'h4296d06a, 32'hc2617f96, 32'hc12c3de0, 32'h42bb2693, 32'hc2876f9f, 32'h42b2c377};
test_bias[2578:2578] = '{32'h42935cd6};
test_output[2578:2578] = '{32'hc60e1d16};
test_input[20632:20639] = '{32'h4233fe10, 32'h41f7d285, 32'h423c3677, 32'h42a6f2c4, 32'hc2629b87, 32'h429a23fd, 32'hc1506963, 32'h42b5642c};
test_weights[20632:20639] = '{32'hc262b84c, 32'hc25cc857, 32'h42ad14eb, 32'h422bd160, 32'hc2719cbe, 32'hc2019702, 32'h42ab980f, 32'hc28b2dbd};
test_bias[2579:2579] = '{32'hc1c4233e};
test_output[2579:2579] = '{32'hc543b30b};
test_input[20640:20647] = '{32'h42a529c7, 32'h41dd7210, 32'h42b4642e, 32'hc1945315, 32'h41d136fa, 32'hc1b840f7, 32'h42b39327, 32'hc189b72b};
test_weights[20640:20647] = '{32'h4102c1da, 32'h42b56a0a, 32'h41dc2a47, 32'h41aa46b1, 32'h40f6496d, 32'h41c9ec41, 32'hc285f2fb, 32'h4299a126};
test_bias[2580:2580] = '{32'hc1eaab62};
test_output[2580:2580] = '{32'hc51a7d8c};
test_input[20648:20655] = '{32'h4265c372, 32'hc2b21b71, 32'h42c172fc, 32'h42c69594, 32'hc28849e4, 32'h4285aa60, 32'h4233f3ab, 32'hc2975c0a};
test_weights[20648:20655] = '{32'hc23b7afd, 32'h428505d1, 32'h42af771f, 32'h4201b99e, 32'h429c88e5, 32'hc24dd165, 32'hc2c314b5, 32'h42ba1e62};
test_bias[2581:2581] = '{32'hc239d7a3};
test_output[2581:2581] = '{32'hc6860dcb};
test_input[20656:20663] = '{32'hc0f9ef3a, 32'hc17797ac, 32'h40fed8ea, 32'hc2814b6a, 32'h42216ecc, 32'hc2b4ad96, 32'hc1b97c68, 32'h42045457};
test_weights[20656:20663] = '{32'hc16e758d, 32'h41d49d1f, 32'hc2c527fa, 32'hc0fe8d71, 32'h424be25c, 32'h41fae7df, 32'hc16804bb, 32'h418126cd};
test_bias[2582:2582] = '{32'hc2b09442};
test_output[2582:2582] = '{32'hc40bf8ef};
test_input[20664:20671] = '{32'hc03aaa38, 32'h41c378fa, 32'hc1e89495, 32'hc28cf6d8, 32'hc296c9e1, 32'h41243233, 32'hc21c48be, 32'hc28d7ae1};
test_weights[20664:20671] = '{32'hc2061e40, 32'hc21166c6, 32'h429459c0, 32'hc26445b2, 32'hc24e5385, 32'h42c09f9b, 32'hc2b3e874, 32'hc29186fc};
test_bias[2583:2583] = '{32'hc2bd9ba0};
test_output[2583:2583] = '{32'h4662df5f};
test_input[20672:20679] = '{32'h429a21b9, 32'h4200f53c, 32'h42a7e16b, 32'hc27c0b7e, 32'h41a0f4a1, 32'hc1a3bf2f, 32'h42821a23, 32'hc134b3ca};
test_weights[20672:20679] = '{32'h42b3e980, 32'h426be411, 32'hc28fd82e, 32'h4238f9d6, 32'h41aa3e9a, 32'h42b47199, 32'h41abcbce, 32'h41bafdf2};
test_bias[2584:2584] = '{32'h400b6f32};
test_output[2584:2584] = '{32'hc3c8565b};
test_input[20680:20687] = '{32'h429a0a6e, 32'hc2888739, 32'h42846273, 32'h4202fd6e, 32'hc1007018, 32'h429291ee, 32'h41f452db, 32'hc2a66743};
test_weights[20680:20687] = '{32'h42213e67, 32'h429787e8, 32'h41e1d867, 32'hc241be8f, 32'hc16dcf10, 32'h41e80cdf, 32'hc281ebcd, 32'h423b9a9c};
test_bias[2585:2585] = '{32'hc2b143b2};
test_output[2585:2585] = '{32'hc5ac5487};
test_input[20688:20695] = '{32'h411f9781, 32'h42c0d171, 32'hc2b13f04, 32'hc1e150da, 32'hc28c631b, 32'h426d2280, 32'h42c44a54, 32'h416a9423};
test_weights[20688:20695] = '{32'h423712a8, 32'hc2b4d2e0, 32'hc2948fad, 32'hc2b2ec72, 32'h40c276d7, 32'hc29e9440, 32'hc28717c6, 32'h4236ff23};
test_bias[2586:2586] = '{32'hc28f71d9};
test_output[2586:2586] = '{32'hc6212b7f};
test_input[20696:20703] = '{32'h41c9311c, 32'hc203ebad, 32'hc2b89f13, 32'hc265ed29, 32'h41117357, 32'h418b72f6, 32'hc29ecd24, 32'hc21b859f};
test_weights[20696:20703] = '{32'h4207ce4f, 32'h4284f599, 32'h425f11c5, 32'h42948bb8, 32'hc2918f6f, 32'h42427140, 32'hc1af008a, 32'h42220d84};
test_bias[2587:2587] = '{32'hc2173790};
test_output[2587:2587] = '{32'hc623390c};
test_input[20704:20711] = '{32'hc2be93df, 32'hc173872c, 32'h424265b8, 32'h4227b058, 32'h42332d89, 32'hc2a80ba7, 32'hc24e2e0a, 32'h420582e0};
test_weights[20704:20711] = '{32'h409cfc82, 32'h41e60da0, 32'h42c1fa75, 32'h41154062, 32'hc2c7cfaf, 32'h42288050, 32'h42273c97, 32'h42b6765d};
test_bias[2588:2588] = '{32'hc217a751};
test_output[2588:2588] = '{32'hc5393109};
test_input[20712:20719] = '{32'h413a7999, 32'h4089f5fe, 32'h428aceca, 32'hc2a4f9fa, 32'h4285c1a9, 32'h42a43492, 32'h415e6178, 32'h42aadb97};
test_weights[20712:20719] = '{32'h42b84103, 32'h427667f9, 32'h42057214, 32'hc1a95fd2, 32'h42280b04, 32'h4272e41d, 32'hc287142b, 32'hc2c2ff76};
test_bias[2589:2589] = '{32'h42087512};
test_output[2589:2589] = '{32'h4577a67f};
test_input[20720:20727] = '{32'h428f5412, 32'h42a39670, 32'h410691c2, 32'hc08ac998, 32'hc2c72aec, 32'h41794f41, 32'hc209d708, 32'h3d7ce9be};
test_weights[20720:20727] = '{32'h42b8b65d, 32'h4261ed1a, 32'h42886435, 32'hc201483a, 32'hc2845fe0, 32'h42ad7f53, 32'h40fd8155, 32'hc29db9bc};
test_bias[2590:2590] = '{32'hc1d96edd};
test_output[2590:2590] = '{32'h46990c1f};
test_input[20728:20735] = '{32'h41c31454, 32'h40a3c428, 32'hc290991b, 32'h41ae9c74, 32'hc2494a2b, 32'hc233eeaa, 32'h425cdfcb, 32'h425e2f07};
test_weights[20728:20735] = '{32'h418ef068, 32'h42ac05bd, 32'hc2768d1c, 32'hc270f0b3, 32'h4286e119, 32'hc22222a1, 32'h42a0554e, 32'hc28e4b69};
test_bias[2591:2591] = '{32'h422d06b8};
test_output[2591:2591] = '{32'h453951ef};
test_input[20736:20743] = '{32'hc29f49c7, 32'h422dcf0b, 32'hc2bbf98c, 32'h4268b541, 32'h41ca4c78, 32'hc2957b1e, 32'hc1455018, 32'hc1ec26a3};
test_weights[20736:20743] = '{32'hc107887c, 32'h4296029f, 32'hc1bf3c4e, 32'h42c0ea11, 32'hc28234f3, 32'h42832cfa, 32'hc2a516df, 32'h41048c0a};
test_bias[2592:2592] = '{32'h42a13d5f};
test_output[2592:2592] = '{32'h45be8e17};
test_input[20744:20751] = '{32'h41f80176, 32'hc236ed13, 32'hc0a525f0, 32'h421bfb62, 32'hc27901b8, 32'h42c6c685, 32'h403eab11, 32'h413290e3};
test_weights[20744:20751] = '{32'h4204da58, 32'hc293c969, 32'hc117e318, 32'hc2b356ef, 32'h424423c1, 32'hc10b10fe, 32'hc1f48631, 32'h41ce59e0};
test_bias[2593:2593] = '{32'hc28bd419};
test_output[2593:2593] = '{32'hc530c4a5};
test_input[20752:20759] = '{32'h4263ece7, 32'h42790793, 32'h42aad291, 32'hc29e3dd5, 32'h414b571c, 32'h421dd647, 32'hc274c0b3, 32'h429c51fd};
test_weights[20752:20759] = '{32'hbf8ded87, 32'hc26cf84e, 32'hc2710c28, 32'hc27c8736, 32'hc20c5399, 32'h42b178cf, 32'h420f67be, 32'h41d39834};
test_bias[2594:2594] = '{32'h40d92c1a};
test_output[2594:2594] = '{32'hc471dcbb};
test_input[20760:20767] = '{32'h428874b7, 32'hc2be996f, 32'hc2be2244, 32'h42890163, 32'hc2087fb1, 32'h4293f1cf, 32'hc2a96cb1, 32'hc2035047};
test_weights[20760:20767] = '{32'hc20abdd9, 32'h4284533c, 32'h41949921, 32'h41817e6d, 32'h42c6a5a5, 32'h4134b2da, 32'hc184b345, 32'h423baf10};
test_bias[2595:2595] = '{32'hc240712d};
test_output[2595:2595] = '{32'hc63c882f};
test_input[20768:20775] = '{32'hc185605a, 32'hc2a25590, 32'h42b2427a, 32'h41eedf64, 32'h4240e11b, 32'h425b5c13, 32'h42c3bcd0, 32'h4263ccf9};
test_weights[20768:20775] = '{32'h4176ff3a, 32'h41098ae4, 32'hc28bf62e, 32'h422b4153, 32'h42b88ba9, 32'hc279a3cc, 32'hc2bc0fb7, 32'h41e9d52b};
test_bias[2596:2596] = '{32'hc1a2479b};
test_output[2596:2596] = '{32'hc6427697};
test_input[20776:20783] = '{32'h41d3ad7f, 32'hc1c1c04d, 32'h4127eda3, 32'h42800695, 32'h428107db, 32'h41ad5bd7, 32'hc26ad5c0, 32'h425a7d38};
test_weights[20776:20783] = '{32'hc2b7b9b7, 32'hc240d777, 32'hc2153c69, 32'hc258fd0a, 32'h41c44c1a, 32'h423fceb5, 32'h41a3889b, 32'h4223dd6f};
test_bias[2597:2597] = '{32'h4239cca7};
test_output[2597:2597] = '{32'hc4b1a011};
test_input[20784:20791] = '{32'hc23e6891, 32'h4185f11e, 32'h427ff2b2, 32'h425aad72, 32'h428e1b50, 32'hc2622a8b, 32'hc21fe1e3, 32'hc1c4da7e};
test_weights[20784:20791] = '{32'hc13b0fec, 32'hc2ac3c6b, 32'hc108bc6a, 32'hc2c0d7dc, 32'h42bcbbf7, 32'h4013b4a6, 32'h41343047, 32'hc2831d04};
test_bias[2598:2598] = '{32'h411ea2d6};
test_output[2598:2598] = '{32'h448281c8};
test_input[20792:20799] = '{32'hc27b6cb4, 32'hc2b154b8, 32'hc2902cca, 32'h42174290, 32'h42b6488a, 32'hbe8ae9ce, 32'h41c4514f, 32'h423968ef};
test_weights[20792:20799] = '{32'hc25539ef, 32'h428b324a, 32'h42671d05, 32'hc218f8f6, 32'hc2649e3f, 32'hc2941d3d, 32'hc2081e00, 32'h4268b90c};
test_bias[2599:2599] = '{32'h424ad0c6};
test_output[2599:2599] = '{32'hc636f0bc};
test_input[20800:20807] = '{32'h42b8e226, 32'h413ed56b, 32'h42c0468e, 32'h4254470b, 32'hc0bfe67e, 32'hc2655cf6, 32'hc1b716db, 32'h42951da8};
test_weights[20800:20807] = '{32'hc2a708f7, 32'hc2aacc8d, 32'hc1af0f71, 32'hc26a0d9d, 32'h41375f93, 32'hc2668a1e, 32'hc12e82ca, 32'h429beb89};
test_bias[2600:2600] = '{32'h409acbfa};
test_output[2600:2600] = '{32'hc59127d6};
test_input[20808:20815] = '{32'h41658c83, 32'hc2000b8b, 32'h42c1dcd9, 32'hc272356f, 32'hc29e76df, 32'h41328f15, 32'h42c68ffe, 32'hc29be8ae};
test_weights[20808:20815] = '{32'hc216eed4, 32'hc2508fb4, 32'hc20ae1c0, 32'hc112a5c1, 32'h4223d371, 32'hc27cae68, 32'hc2c47429, 32'hc2200934};
test_bias[2601:2601] = '{32'hc2a45e4c};
test_output[2601:2601] = '{32'hc640f0e4};
test_input[20816:20823] = '{32'h42b01265, 32'h426b9dc5, 32'hc1a3af2d, 32'h42742fa1, 32'h411b2ef9, 32'h4240a5a0, 32'h42b43c17, 32'hc0e944e2};
test_weights[20816:20823] = '{32'hc2a80920, 32'h41ed84e3, 32'hc0ff0178, 32'h42b20c64, 32'hc266ad91, 32'h41a2a7ef, 32'h426df4cb, 32'hc29184db};
test_bias[2602:2602] = '{32'h42922fae};
test_output[2602:2602] = '{32'h45c5f272};
test_input[20824:20831] = '{32'h429cf0b4, 32'h4200d334, 32'hc259d326, 32'hc29f9310, 32'h4223518d, 32'h42063351, 32'h42b3b1a1, 32'hc1bf71df};
test_weights[20824:20831] = '{32'hc227dbba, 32'hc2180e2b, 32'h4249a93b, 32'h42ac0fb3, 32'hc1804446, 32'h42a0f52e, 32'hc1837db9, 32'h4145f968};
test_bias[2603:2603] = '{32'hc20f58ed};
test_output[2603:2603] = '{32'hc6590852};
test_input[20832:20839] = '{32'hc2b3e150, 32'hc257d98a, 32'hc142705f, 32'hc13781cb, 32'h40a45813, 32'hc2642b21, 32'hc2867b00, 32'hc01a625d};
test_weights[20832:20839] = '{32'hc22267af, 32'hc296ad7b, 32'hc2b9bbcd, 32'hc0b07643, 32'h4249f9d1, 32'hc183c83d, 32'h41fc10c7, 32'hc1919bce};
test_bias[2604:2604] = '{32'hc28e1336};
test_output[2604:2604] = '{32'h45f8d155};
test_input[20840:20847] = '{32'h416717fc, 32'h423b278b, 32'hc109e327, 32'h407f4ee8, 32'h4220a699, 32'h42b94981, 32'hc26ebaf1, 32'hc29e4334};
test_weights[20840:20847] = '{32'h428fa817, 32'h423074b0, 32'hc27b09c3, 32'hc2777d24, 32'h42bc0d04, 32'hc10d541d, 32'h428985ef, 32'hc2b68ecb};
test_bias[2605:2605] = '{32'hc1e90fad};
test_output[2605:2605] = '{32'h46138e0f};
test_input[20848:20855] = '{32'h42934682, 32'hc1e2594c, 32'h42a2ef0d, 32'hc22679b5, 32'hc27fb177, 32'hc250f1f7, 32'hc19941d3, 32'h416c9ede};
test_weights[20848:20855] = '{32'h420fb362, 32'h42a99b30, 32'hc2365fa0, 32'hc26775c6, 32'hc2759b6a, 32'hc241638a, 32'h4211a8cb, 32'hc25275ae};
test_bias[2606:2606] = '{32'h42930446};
test_output[2606:2606] = '{32'h45794436};
test_input[20856:20863] = '{32'h421c9246, 32'hc28fdf9f, 32'hc22b62b6, 32'hc1221527, 32'hc25efa1d, 32'h42570e18, 32'hc2b94a52, 32'hc0fcbfe1};
test_weights[20856:20863] = '{32'h428a4dc6, 32'hc2537f17, 32'hc17f481e, 32'h41004662, 32'h421d33e2, 32'h42bd6dad, 32'h40424d8e, 32'hc26c4993};
test_bias[2607:2607] = '{32'h429e7cbf};
test_output[2607:2607] = '{32'h46209b03};
test_input[20864:20871] = '{32'h42bf87c9, 32'h410a6dc8, 32'h4225a23d, 32'hc2459ace, 32'h428a79de, 32'h423e7ee9, 32'h4264be54, 32'hc236572f};
test_weights[20864:20871] = '{32'h4119d880, 32'hc297c68d, 32'hc27246a9, 32'h40f5cde8, 32'hc282f715, 32'h42b80113, 32'h42835350, 32'h41f89375};
test_bias[2608:2608] = '{32'hc2a440d2};
test_output[2608:2608] = '{32'hc401cf39};
test_input[20872:20879] = '{32'hc10ceced, 32'h4181bf89, 32'hc08c31fc, 32'hc224192b, 32'h422bcb3c, 32'h4296fc8e, 32'h401be76a, 32'hc0b7c269};
test_weights[20872:20879] = '{32'h42643530, 32'hc2c7d610, 32'hc20088b3, 32'h42c0d227, 32'hc27c8722, 32'hc201ab02, 32'h42c573c8, 32'h42981bdc};
test_bias[2609:2609] = '{32'h429fa40b};
test_output[2609:2609] = '{32'hc62f323a};
test_input[20880:20887] = '{32'h414b3ae3, 32'h423b89ac, 32'h3f979b57, 32'h42691a79, 32'h40fc8409, 32'h415f3b2c, 32'h41d225a3, 32'h426dd986};
test_weights[20880:20887] = '{32'h4182fe05, 32'hc296ebe0, 32'h42667c44, 32'h4216a1d2, 32'h4276d9f0, 32'hc156fbad, 32'hc2c282c7, 32'h422a9dc7};
test_bias[2610:2610] = '{32'h42c1d2e7};
test_output[2610:2610] = '{32'hc42c495d};
test_input[20888:20895] = '{32'hc0a58340, 32'h40a43aca, 32'h42c65c09, 32'hc10d5a7d, 32'h411433e1, 32'hc186e299, 32'hc14e63d4, 32'h4186c5c2};
test_weights[20888:20895] = '{32'hc21da4b0, 32'h42c74a9d, 32'h426db60a, 32'hc281b7d5, 32'hc1f5d7ad, 32'h4299cc1a, 32'h421632df, 32'h41708ffa};
test_bias[2611:2611] = '{32'h429ae9d4};
test_output[2611:2611] = '{32'h45aa3ba0};
test_input[20896:20903] = '{32'hc2886b62, 32'hc1acce32, 32'hc23bef4d, 32'hc21f9eae, 32'hc282facc, 32'h407b3057, 32'hc2bb231a, 32'hc2ac6639};
test_weights[20896:20903] = '{32'h428aa4c4, 32'h41a41d00, 32'h414b190a, 32'h41214986, 32'h426cbce0, 32'hc2325061, 32'h42b967fe, 32'h40ae40e8};
test_bias[2612:2612] = '{32'h40f439e7};
test_output[2612:2612] = '{32'hc69739fe};
test_input[20904:20911] = '{32'hc2bf267b, 32'h42846c03, 32'hc12d101f, 32'hc2c21abd, 32'hc299f4f7, 32'hc00602b5, 32'h42176855, 32'hc251fd86};
test_weights[20904:20911] = '{32'hc2802e50, 32'h421dfb03, 32'h4285cb35, 32'h418c6132, 32'h4238406b, 32'h42656dda, 32'h41cf02fd, 32'h42665513};
test_bias[2613:2613] = '{32'hc2638432};
test_output[2613:2613] = '{32'h4408e1cb};
test_input[20912:20919] = '{32'h42a61af5, 32'hc21a8dbb, 32'h42bfb84f, 32'hc2988186, 32'hc2467ae5, 32'hc2a12a82, 32'hc208e170, 32'h429166dd};
test_weights[20912:20919] = '{32'hc1a49524, 32'h41cd63d0, 32'h4214f4f0, 32'hc2b68d47, 32'hc19b3636, 32'hc2a18ccc, 32'hc005e23a, 32'h423101a2};
test_bias[2614:2614] = '{32'hc25358e0};
test_output[2614:2614] = '{32'h4690d1bb};
test_input[20920:20927] = '{32'h41bd6aad, 32'h424f7c25, 32'h42455747, 32'hc284b33e, 32'hc1ecd81e, 32'h41d79898, 32'h42205e2d, 32'h42407274};
test_weights[20920:20927] = '{32'h421c2bb1, 32'h41b8012a, 32'h4208e7ea, 32'hc23e0d73, 32'h428d6059, 32'h4220d08f, 32'h4292a9e3, 32'h428d9cc9};
test_bias[2615:2615] = '{32'h41f4661c};
test_output[2615:2615] = '{32'h464099c7};
test_input[20928:20935] = '{32'h424c0ce0, 32'hc28986f4, 32'h422eb0b6, 32'hc21993d4, 32'h3f80517a, 32'h42a306b9, 32'h423702fa, 32'h410bfd5b};
test_weights[20928:20935] = '{32'h40fc6d0a, 32'h41efbc44, 32'h42317391, 32'hc2310c04, 32'hc18a3598, 32'hc1e2c52c, 32'h428f58ed, 32'hc152e0f3};
test_bias[2616:2616] = '{32'h429ef48c};
test_output[2616:2616] = '{32'h4534e23b};
test_input[20936:20943] = '{32'h42b1d78d, 32'h410a0af9, 32'hc2b32fbf, 32'h4202feb0, 32'hc1887d83, 32'hc2c34034, 32'hc1c44217, 32'h42a03c53};
test_weights[20936:20943] = '{32'h4282e7ef, 32'hc2ac5ead, 32'hc1bafcdd, 32'hc1bad2e2, 32'hc1359307, 32'h4291e297, 32'hc2c68fe6, 32'hc28e65ff};
test_bias[2617:2617] = '{32'hc21ce8a8};
test_output[2617:2617] = '{32'hc56f57f1};
test_input[20944:20951] = '{32'hc28d7635, 32'hc2124b1d, 32'h421e84ed, 32'h423dca2f, 32'h427446cb, 32'h424fd25e, 32'h41b04918, 32'h428cbd4a};
test_weights[20944:20951] = '{32'h42027aa8, 32'hc250a709, 32'hc27c7d4a, 32'h42582e8c, 32'hc246adc1, 32'h417f30b0, 32'hc20b2da1, 32'hc1182217};
test_bias[2618:2618] = '{32'h42b050ef};
test_output[2618:2618] = '{32'hc5730f14};
test_input[20952:20959] = '{32'h42c35bca, 32'hc0eaf5ff, 32'h420f9116, 32'h42397f2a, 32'h41dc3ca4, 32'hc2074002, 32'h42b443b3, 32'hc1ac97c2};
test_weights[20952:20959] = '{32'hbf02eb27, 32'hc0fcd492, 32'h42b822f6, 32'h4265a7a3, 32'hc28d68d7, 32'hc252f10a, 32'h424102a8, 32'h42002f99};
test_bias[2619:2619] = '{32'hc1d4c8c3};
test_output[2619:2619] = '{32'h46138b5e};
test_input[20960:20967] = '{32'h42157000, 32'h42beac32, 32'hc2c520d7, 32'hc2c5622b, 32'h426c8296, 32'hc1b60b55, 32'hc13e9528, 32'hc2991fdb};
test_weights[20960:20967] = '{32'h41beeec2, 32'h41650b4b, 32'hc1f9265f, 32'h424b89f4, 32'hc2273dad, 32'hc001cc7f, 32'h423f462d, 32'hc2ad2b85};
test_bias[2620:2620] = '{32'h4130e7f0};
test_output[2620:2620] = '{32'h4576cc8c};
test_input[20968:20975] = '{32'h420e5ed3, 32'hc27f71c4, 32'hc15f2521, 32'hc2733fe7, 32'h428e6a54, 32'h41c1ebc1, 32'hc28acba5, 32'hc0d2bdcf};
test_weights[20968:20975] = '{32'h4288c101, 32'h425fee23, 32'hc1947cb5, 32'h42059c98, 32'h426d8848, 32'hc0f37420, 32'h40a61454, 32'h428273c5};
test_bias[2621:2621] = '{32'hc293761f};
test_output[2621:2621] = '{32'h4385676c};
test_input[20976:20983] = '{32'h426a1399, 32'h3f59fd7b, 32'h41858083, 32'hc1f296a0, 32'h426421ba, 32'hc2052659, 32'h41dca038, 32'hc2a51635};
test_weights[20976:20983] = '{32'h4267940c, 32'hc2bc7c1b, 32'h40d27d29, 32'h41b673ba, 32'hc2a6eebb, 32'hc171b48c, 32'hc2884fba, 32'hc2baf311};
test_bias[2622:2622] = '{32'h4290636a};
test_output[2622:2622] = '{32'h4588c5c0};
test_input[20984:20991] = '{32'hc29107bf, 32'h428b044c, 32'hc222c46e, 32'hc003b028, 32'hc29c8197, 32'h4292370c, 32'hc2b0635c, 32'hc23c5617};
test_weights[20984:20991] = '{32'hbf8742fe, 32'hc18f9b0d, 32'hc00d4336, 32'hc2587a8c, 32'hc289bf61, 32'hc1e868f0, 32'hc21537f5, 32'h426dac0d};
test_bias[2623:2623] = '{32'hc1da888c};
test_output[2623:2623] = '{32'h452c8e41};
test_input[20992:20999] = '{32'hc183ca91, 32'h40f31af9, 32'h4292fb0a, 32'h4049bd44, 32'hc226bec4, 32'h429c303e, 32'hc155358a, 32'hc2907762};
test_weights[20992:20999] = '{32'hc2541468, 32'hbfa6c7e8, 32'h42c0c272, 32'h42725cd2, 32'hc289f182, 32'h4292a3e0, 32'hc2bcceac, 32'h423b5368};
test_bias[2624:2624] = '{32'h42831714};
test_output[2624:2624] = '{32'h46655d3e};
test_input[21000:21007] = '{32'h41a8c94f, 32'h425187d7, 32'hc23e8702, 32'h42b5210b, 32'hc1e91a4d, 32'h41c7b68e, 32'h4231f87e, 32'h4199bbba};
test_weights[21000:21007] = '{32'hc2933cf8, 32'hc2261f53, 32'h3f5fea93, 32'h406f8296, 32'hc241a9ef, 32'h424c03d9, 32'h429fa15f, 32'hc287735a};
test_bias[2625:2625] = '{32'hc285d9fc};
test_output[2625:2625] = '{32'h44b36b4e};
test_input[21008:21015] = '{32'hc1d1d62e, 32'hc2c23ef8, 32'hc05b3866, 32'h41f7b197, 32'hc25832c4, 32'hc1ab9a78, 32'h425b6b71, 32'h41dbd0fa};
test_weights[21008:21015] = '{32'hc2852db6, 32'h4092fe54, 32'hc2855899, 32'hc2a9b709, 32'h427d3b9d, 32'h41887360, 32'h426e5f85, 32'hc21c07e8};
test_bias[2626:2626] = '{32'hc167c64a};
test_output[2626:2626] = '{32'hc528f73e};
test_input[21016:21023] = '{32'h4282cac0, 32'h429793db, 32'hc1909327, 32'hc1a8f55e, 32'h42902284, 32'h408b2dc0, 32'hc1bb6c2b, 32'hc207df67};
test_weights[21016:21023] = '{32'hc2b96061, 32'hc21a3d31, 32'h41ab6df9, 32'hc2402fb1, 32'h41de7090, 32'h41da59d7, 32'hc1d8bb2a, 32'h4280607a};
test_bias[2627:2627] = '{32'hc1e4e7ab};
test_output[2627:2627] = '{32'hc5f400ce};
test_input[21024:21031] = '{32'hc252d29e, 32'h42b6d9c3, 32'hc29aed42, 32'hc18267d4, 32'hc0a39d09, 32'hc27495ab, 32'hc28c1c40, 32'h41ee581e};
test_weights[21024:21031] = '{32'hc12d64cc, 32'h41c53332, 32'hc187ef3c, 32'h42c4805d, 32'h418021e9, 32'h427ba3d6, 32'hc204e625, 32'h4251524c};
test_bias[2628:2628] = '{32'hc2844715};
test_output[2628:2628] = '{32'h4517f690};
test_input[21032:21039] = '{32'hc0159f4c, 32'hc29171bd, 32'h42c6642d, 32'hc2809d98, 32'h4252f16e, 32'hc2b009b6, 32'hc1514d0e, 32'h407e4536};
test_weights[21032:21039] = '{32'h3fbe0c85, 32'hc28a7269, 32'hc2954a09, 32'h416f0bf6, 32'h4293c918, 32'h42aedc35, 32'hc2a7d29f, 32'hc0d64f27};
test_bias[2629:2629] = '{32'hc20ec6ca};
test_output[2629:2629] = '{32'hc5be8f8d};
test_input[21040:21047] = '{32'h429a767b, 32'hc1f6d5cd, 32'h426b3ef0, 32'h426b2c82, 32'hc2c116e2, 32'hc21419e1, 32'hc25d85b4, 32'h42069a91};
test_weights[21040:21047] = '{32'h42bc9661, 32'h429987b4, 32'h41ce75f3, 32'hc1d0ea05, 32'hc1f69ce7, 32'h421ae695, 32'hc18aa929, 32'h4283bbf6};
test_bias[2630:2630] = '{32'h411ea605};
test_output[2630:2630] = '{32'h461663d9};
test_input[21048:21055] = '{32'hc1c85a59, 32'hc29a82cf, 32'h422fd429, 32'h423f2ab8, 32'h41ddfe20, 32'hc2b28992, 32'hc22a4f85, 32'hc2c51c78};
test_weights[21048:21055] = '{32'hc2bc6b4e, 32'h42c42416, 32'hc26d8b14, 32'h420b467e, 32'hc2bc6f4e, 32'hc20d4f9e, 32'h402e9a0c, 32'h42c1b7fd};
test_bias[2631:2631] = '{32'hc2c55f93};
test_output[2631:2631] = '{32'hc6706484};
test_input[21056:21063] = '{32'h425a0af1, 32'hc1f4ea61, 32'hc28a7883, 32'hc2597494, 32'h42073a12, 32'h418316a0, 32'h410760e2, 32'hc1dd907f};
test_weights[21056:21063] = '{32'h41a2ba4d, 32'hc2843391, 32'hc2c52370, 32'h42b25d60, 32'h429c02bc, 32'h4053b7d6, 32'hc2931807, 32'hc18b77dd};
test_bias[2632:2632] = '{32'h420b34c9};
test_output[2632:2632] = '{32'h45f07a24};
test_input[21064:21071] = '{32'h428af183, 32'h41323070, 32'h4283460c, 32'h422e9524, 32'hc29c1960, 32'h3d940c5d, 32'hc2acb692, 32'hc211977d};
test_weights[21064:21071] = '{32'h421c7c12, 32'hc283cbc5, 32'h42b3c86f, 32'hc201a3b0, 32'hc2bf4a60, 32'h40b7469d, 32'h42bf7220, 32'hc239a6ba};
test_bias[2633:2633] = '{32'hc2afe36f};
test_output[2633:2633] = '{32'h45e33108};
test_input[21072:21079] = '{32'h42428f9c, 32'h42a506ea, 32'hc1e23793, 32'h40b8e1d5, 32'h41eabfd4, 32'h42b35828, 32'hc243d23c, 32'hc2182123};
test_weights[21072:21079] = '{32'hc1ae3e5f, 32'hc27dcbcb, 32'hc1de32ad, 32'hc257e87d, 32'h42551256, 32'hc17e9bed, 32'h42628618, 32'hc21d0964};
test_bias[2634:2634] = '{32'hc045c447};
test_output[2634:2634] = '{32'hc5d9bc1c};
test_input[21080:21087] = '{32'hc1817c0c, 32'hc26fb9b5, 32'hc284bcde, 32'h4180ebc0, 32'hc2aa743f, 32'hc22072a1, 32'hc27df7fd, 32'hc247a366};
test_weights[21080:21087] = '{32'hc12c46e4, 32'hbfef9a67, 32'hc1ab3a57, 32'h415737b5, 32'hc2adc4ec, 32'h428ef23a, 32'hc183bcc8, 32'h4293027f};
test_bias[2635:2635] = '{32'h3faf18fa};
test_output[2635:2635] = '{32'h457000dd};
test_input[21088:21095] = '{32'hc293cdb4, 32'hc2c3b474, 32'h409c6b1c, 32'h414e10e6, 32'hc2c3abc7, 32'h40f78af2, 32'h41e1a4e3, 32'hc295e54d};
test_weights[21088:21095] = '{32'hc23100f4, 32'hc28ebac4, 32'hc2983310, 32'hc2b5f6ef, 32'h42440433, 32'hc200cf0d, 32'hc205a8d9, 32'h4293618d};
test_bias[2636:2636] = '{32'h41d7192c};
test_output[2636:2636] = '{32'hc52d44e2};
test_input[21096:21103] = '{32'hc2b7f04c, 32'h4196fc39, 32'h41eb62b6, 32'h416a8715, 32'h4269821c, 32'h428666e5, 32'h42984084, 32'h41de5829};
test_weights[21096:21103] = '{32'hc10588e0, 32'h424421a7, 32'hc2072d93, 32'h42b689a0, 32'h4211ae6d, 32'h427ac210, 32'h3ec9590f, 32'hc28ee514};
test_bias[2637:2637] = '{32'hc21388d2};
test_output[2637:2637] = '{32'h45c77556};
test_input[21104:21111] = '{32'h42400e6e, 32'hc2a6e250, 32'hc2945de2, 32'hc2902dcb, 32'hc284123f, 32'h41472781, 32'h4278b1b8, 32'h424a9c81};
test_weights[21104:21111] = '{32'h42afd7cd, 32'hc219ea5a, 32'hc12d484b, 32'hc2a80c7f, 32'hc2c4ce5a, 32'hc20614fa, 32'hc1959516, 32'hc2698212};
test_bias[2638:2638] = '{32'hc19e82ef};
test_output[2638:2638] = '{32'h467daa02};
test_input[21112:21119] = '{32'h41888eb9, 32'h4232511f, 32'h42a29d9e, 32'hc1ba0559, 32'hc2848188, 32'h40288b7a, 32'h428c689f, 32'h42b5b22e};
test_weights[21112:21119] = '{32'hc1ca81f0, 32'h42922dac, 32'h41875099, 32'h4166daf7, 32'hc2766d53, 32'h41151d3b, 32'h40d16ba8, 32'h4289f70e};
test_bias[2639:2639] = '{32'hc28f4faf};
test_output[2639:2639] = '{32'h46648b4f};
test_input[21120:21127] = '{32'hc2ac7d71, 32'h41e87707, 32'h41b0de81, 32'h41f82810, 32'h429bae07, 32'h422a3342, 32'h4144cc28, 32'h42c62499};
test_weights[21120:21127] = '{32'h40c6e70d, 32'h41cd2005, 32'hc190b63c, 32'h42900321, 32'h41927d69, 32'hc20436e1, 32'hc24f5613, 32'hc2a67711};
test_bias[2640:2640] = '{32'h42a81fed};
test_output[2640:2640] = '{32'hc5d28f06};
test_input[21128:21135] = '{32'hc2947dca, 32'hc1336c4a, 32'h42b734f5, 32'h42a33c42, 32'h42044e8c, 32'h419c1400, 32'h4298dcab, 32'h4041af02};
test_weights[21128:21135] = '{32'h41c51d5f, 32'h41bfeefd, 32'h42122204, 32'h4232a172, 32'h428add52, 32'hc2c63e66, 32'h42512897, 32'h42b57f31};
test_bias[2641:2641] = '{32'h42889ee6};
test_output[2641:2641] = '{32'h4615ed06};
test_input[21136:21143] = '{32'hc1013a5f, 32'hc25188de, 32'h42a95329, 32'h41983747, 32'hc29fce07, 32'h3f94ffff, 32'h4283b240, 32'h428ffc7d};
test_weights[21136:21143] = '{32'hc2376bca, 32'hc251513e, 32'h3ffb48e0, 32'h427474ed, 32'h42b60500, 32'hc29457db, 32'h42b0a5fd, 32'hc0e8082a};
test_bias[2642:2642] = '{32'hc2953040};
test_output[2642:2642] = '{32'h450fdb7f};
test_input[21144:21151] = '{32'hc1c7dfb6, 32'h4204c200, 32'h42c6c076, 32'h42a40ca5, 32'h4183654a, 32'hc274b04d, 32'hc26ee9fa, 32'hc2826cf4};
test_weights[21144:21151] = '{32'hc28287c0, 32'hc2c15090, 32'hc1e6c07b, 32'hc2b7067f, 32'hc2492104, 32'hbefd199c, 32'h401464ae, 32'h40195938};
test_bias[2643:2643] = '{32'hc210cc99};
test_output[2643:2643] = '{32'hc64c52a9};
test_input[21152:21159] = '{32'h4231ff38, 32'hc24f9dd5, 32'h4237bc21, 32'h41d5f7ba, 32'hc265d15e, 32'hc15e18eb, 32'hc2498059, 32'h426e7378};
test_weights[21152:21159] = '{32'h4208e971, 32'h421cc2e4, 32'hc258c24d, 32'hc14fca0e, 32'h42928445, 32'h428b2ac1, 32'hc24a7221, 32'hc1fe3b20};
test_bias[2644:2644] = '{32'hc1b37ced};
test_output[2644:2644] = '{32'hc5f68dac};
test_input[21160:21167] = '{32'hc272164b, 32'hc2ab96b2, 32'h427ec929, 32'hc2912b82, 32'hc24e7ef4, 32'h42651e57, 32'hc1e003ed, 32'h40c7d9c5};
test_weights[21160:21167] = '{32'hc2bf8cc7, 32'hc1f3f6e0, 32'h4203b130, 32'h421d1b14, 32'hc2bd3c52, 32'h415c76db, 32'h429acf01, 32'h42647128};
test_bias[2645:2645] = '{32'hc285d958};
test_output[2645:2645] = '{32'h4632fc66};
test_input[21168:21175] = '{32'h428c6009, 32'h41802652, 32'hc29c91cc, 32'hbef4bcb1, 32'h42611898, 32'hc207c294, 32'hc2131848, 32'hc195ba88};
test_weights[21168:21175] = '{32'h420f02ca, 32'hc25d1f02, 32'hc26122ee, 32'h42576eb3, 32'h42ad6cad, 32'hc20452cb, 32'h42a16f7c, 32'hc28dd181};
test_bias[2646:2646] = '{32'hc24e5d18};
test_output[2646:2646] = '{32'h462127f9};
test_input[21176:21183] = '{32'hc2b924c4, 32'h42aa1fdb, 32'hc2909bd7, 32'h4244ea1d, 32'hc20b2ac3, 32'hc27525ba, 32'h3fb70f52, 32'hc2906d18};
test_weights[21176:21183] = '{32'h42961a47, 32'hc191f982, 32'hc2a206e9, 32'hc1a5fb09, 32'hc0801446, 32'hc2c7aa66, 32'h42013890, 32'h42aa2181};
test_bias[2647:2647] = '{32'hc2b5a2b7};
test_output[2647:2647] = '{32'hc5609425};
test_input[21184:21191] = '{32'hc2bad011, 32'h42bfb4bf, 32'hc2b23921, 32'hc2aa2acb, 32'hc29ea7ea, 32'hc25945b8, 32'hc24af057, 32'hc1e7242a};
test_weights[21184:21191] = '{32'hc1097170, 32'h42031b3e, 32'h4113845f, 32'h425f9171, 32'hc2987329, 32'hc1ef7ab4, 32'hc128dd30, 32'hc2bed89c};
test_bias[2648:2648] = '{32'hc2a5e516};
test_output[2648:2648] = '{32'h46108557};
test_input[21192:21199] = '{32'h42607fbf, 32'hc1fe4d9c, 32'h422e578b, 32'hc2483f34, 32'h41727311, 32'hc1a611cc, 32'hc1b439a6, 32'hc2894222};
test_weights[21192:21199] = '{32'hc21b0198, 32'h429b71f5, 32'hc286d664, 32'hc2757aa8, 32'hc0714bf9, 32'h428fe45d, 32'h421ef2b6, 32'h427f7866};
test_bias[2649:2649] = '{32'h4122a545};
test_output[2649:2649] = '{32'hc6310a72};
test_input[21200:21207] = '{32'hc2abcb52, 32'hc27a9d59, 32'h4212ab62, 32'h41cf2c14, 32'hc1d70d4c, 32'h42bc0d19, 32'hc211ea83, 32'hc1afe4ef};
test_weights[21200:21207] = '{32'h4253f41b, 32'h42b2e800, 32'hc27e1ad2, 32'h42681277, 32'hc2bfcc0f, 32'h3f366009, 32'h426c6584, 32'h41929308};
test_bias[2650:2650] = '{32'h4249ebe9};
test_output[2650:2650] = '{32'hc629795f};
test_input[21208:21215] = '{32'hc1754d4f, 32'hc01df5fe, 32'h415e950c, 32'h42a9f9ec, 32'hc1708adb, 32'hc2ab98dd, 32'hc1cc8273, 32'hc2a64466};
test_weights[21208:21215] = '{32'h42b2a9b2, 32'hc274e379, 32'h42aa02b8, 32'hc2662f60, 32'hc2942b5b, 32'h4030829d, 32'hc28ecdf0, 32'hc2afa3a0};
test_bias[2651:2651] = '{32'h3faadeeb};
test_output[2651:2651] = '{32'h459eaefb};
test_input[21216:21223] = '{32'h41aee26e, 32'hc0e57c94, 32'hc286a3c5, 32'hc2bdf17a, 32'h41cbe7a5, 32'h40e2c35f, 32'h42552b00, 32'h41ef2cdb};
test_weights[21216:21223] = '{32'h417f1cc8, 32'hc26024cf, 32'hc2b01b7d, 32'h40b21588, 32'hc2c363c6, 32'h428e7642, 32'h426ca25c, 32'h41ee12e2};
test_bias[2652:2652] = '{32'h416cfbab};
test_output[2652:2652] = '{32'h46007639};
test_input[21224:21231] = '{32'h4042b5de, 32'h40bf976c, 32'hc25d5e38, 32'h429c8086, 32'h42c5cb59, 32'h417bf472, 32'hc1a56da1, 32'hc2a51f1f};
test_weights[21224:21231] = '{32'h42a737ee, 32'hc075e344, 32'hc2862840, 32'hc1c328c1, 32'h41cdd0dc, 32'hc2af52a1, 32'hc2735856, 32'hc206a494};
test_bias[2653:2653] = '{32'hc2c53779};
test_output[2653:2653] = '{32'h45df0881};
test_input[21232:21239] = '{32'h42726288, 32'hc1ef1aa9, 32'h42a64aab, 32'h42a4741f, 32'h4231af18, 32'hc29e832a, 32'h42a84e03, 32'hc2503c8e};
test_weights[21232:21239] = '{32'hc1a2f2eb, 32'hc2376466, 32'h42025e83, 32'h428f3943, 32'hc194e763, 32'h4224e31a, 32'h40a32bf1, 32'h4277df86};
test_bias[2654:2654] = '{32'h4180a9f7};
test_output[2654:2654] = '{32'h44e874f1};
test_input[21240:21247] = '{32'h3f956a0d, 32'hc2844659, 32'h4244c93d, 32'hc1e32b25, 32'hc2b59cef, 32'h42c14dad, 32'h425bf241, 32'hc279fea7};
test_weights[21240:21247] = '{32'hc2927ae0, 32'h40f4fb2b, 32'hc242f4c8, 32'h422f4668, 32'h429a7207, 32'hc24c077d, 32'hc28b749f, 32'h4086e1d9};
test_bias[2655:2655] = '{32'h3e4a602e};
test_output[2655:2655] = '{32'hc69e62fa};
test_input[21248:21255] = '{32'h41437cc3, 32'hc15c9032, 32'h425a9de0, 32'h425907b5, 32'h42982dc3, 32'h426d12ed, 32'h425a96cc, 32'h425dd294};
test_weights[21248:21255] = '{32'hc27ddf3c, 32'hc28526eb, 32'hc27f7ea8, 32'hc2b7ca23, 32'h420f006a, 32'h41d84779, 32'hc28b294a, 32'hc293c362};
test_bias[2656:2656] = '{32'h41c8b76c};
test_output[2656:2656] = '{32'hc639ba2d};
test_input[21256:21263] = '{32'h41a5b7e2, 32'h414f45f4, 32'hc2998f6b, 32'h42913233, 32'h4236885f, 32'hc2b3b5fb, 32'h41e74dff, 32'hbfb5cbe2};
test_weights[21256:21263] = '{32'h42a97dee, 32'h42823cf7, 32'h41e4a75a, 32'hc2a9c53f, 32'h40c25cd8, 32'h42acd74a, 32'hc290b0f1, 32'hc1bdb06b};
test_bias[2657:2657] = '{32'h42455801};
test_output[2657:2657] = '{32'hc66e5b51};
test_input[21264:21271] = '{32'hc1aa1ded, 32'h42ba67b5, 32'hc297103d, 32'hc28678b1, 32'h42a1f293, 32'h42c352e4, 32'hc29d7f87, 32'h42829b33};
test_weights[21264:21271] = '{32'h42518b70, 32'h424500b4, 32'h42b897f8, 32'h4283a4d1, 32'h413efd13, 32'h4238663e, 32'h429f7176, 32'h42844b25};
test_bias[2658:2658] = '{32'hc291c708};
test_output[2658:2658] = '{32'hc58c191c};
test_input[21272:21279] = '{32'hc2a8f755, 32'h42afab8b, 32'hc27babdc, 32'h41592e89, 32'h428a7262, 32'hc2983246, 32'h4294c57e, 32'hc2bf72db};
test_weights[21272:21279] = '{32'h42bd9190, 32'hc2b24749, 32'hc15c1148, 32'hc11e2445, 32'h40943792, 32'hc143840e, 32'hc1cdb07e, 32'hc274d937};
test_bias[2659:2659] = '{32'h41e4c959};
test_output[2659:2659] = '{32'hc61a5fb0};
test_input[21280:21287] = '{32'h42afc756, 32'hc2a072a4, 32'h4259ee14, 32'hc2314fea, 32'h42c69238, 32'h42c7af41, 32'hc233462d, 32'h42bd211e};
test_weights[21280:21287] = '{32'hc1dff116, 32'h426a1c03, 32'hc2190466, 32'hc2115381, 32'hc2a74887, 32'hc2148854, 32'hc1b79c1f, 32'h42bcc141};
test_bias[2660:2660] = '{32'h4235ec4d};
test_output[2660:2660] = '{32'hc616a8d7};
test_input[21288:21295] = '{32'h419da194, 32'hc24887ed, 32'h42be9378, 32'hc06bab09, 32'h42797dd8, 32'hc1cf6d16, 32'hc1f21200, 32'h42509c63};
test_weights[21288:21295] = '{32'h4160c66c, 32'h422cc8d9, 32'h42a9e4c3, 32'h429520e1, 32'hc2ae104e, 32'h41b31cc6, 32'hc1c1d7d1, 32'h412d5043};
test_bias[2661:2661] = '{32'hc263dd58};
test_output[2661:2661] = '{32'h44916a0c};
test_input[21296:21303] = '{32'h428399d4, 32'h411cabaa, 32'h41838bac, 32'h41324eea, 32'hc2bea666, 32'h42b79145, 32'hc28b81f7, 32'hc142cb97};
test_weights[21296:21303] = '{32'hc2922592, 32'h4295e959, 32'hc2c6abbc, 32'hc22de8d6, 32'hc12055eb, 32'hc29430e5, 32'hc2ba2f35, 32'h420ba676};
test_bias[2662:2662] = '{32'hc2aaeab9};
test_output[2662:2662] = '{32'hc5bd3597};
test_input[21304:21311] = '{32'h419651f5, 32'hc1c9bf7c, 32'h40ad9716, 32'hc1184321, 32'h42b04974, 32'hc25a2a64, 32'h420d0267, 32'h428627dd};
test_weights[21304:21311] = '{32'h42996c91, 32'h42812216, 32'h406d080c, 32'h4091105a, 32'h421a36dd, 32'h418a8ad9, 32'hc1335188, 32'hc1cf67e7};
test_bias[2663:2663] = '{32'hc2938d14};
test_output[2663:2663] = '{32'h420f9cbd};
test_input[21312:21319] = '{32'hc244680e, 32'hc124b651, 32'h4225c977, 32'hc2276974, 32'h4205b39e, 32'hc196f1a9, 32'hc15817b8, 32'h408c226f};
test_weights[21312:21319] = '{32'h410c3a2b, 32'h4117c7b6, 32'hc1d5c6d5, 32'hc187c54d, 32'hc29a9300, 32'hc28b1cad, 32'hc2158f58, 32'hc29354c2};
test_bias[2664:2664] = '{32'hc25d436d};
test_output[2664:2664] = '{32'hc501522f};
test_input[21320:21327] = '{32'h42a6e7cc, 32'h429f4744, 32'h42b87a32, 32'hc2b411c6, 32'h429517d0, 32'hc2851294, 32'hc1c862e5, 32'h4291fbca};
test_weights[21320:21327] = '{32'hc2856697, 32'h42bf91b6, 32'h413fa80b, 32'hc1f06789, 32'hc275ef01, 32'hc0d5aea3, 32'hc29bf634, 32'hc1c6003b};
test_bias[2665:2665] = '{32'h4225921d};
test_output[2665:2665] = '{32'h44f02d14};
test_input[21328:21335] = '{32'hc24fd0b1, 32'hc26bba61, 32'hc26f8715, 32'h41a285b8, 32'hc26ab601, 32'h425f6dc3, 32'h42c784d1, 32'h420d1e3f};
test_weights[21328:21335] = '{32'h427c920a, 32'hc2bbe99f, 32'hc2863633, 32'hc29c9b18, 32'hc2077c76, 32'hc2b0e860, 32'hc26e5c66, 32'hc2920e23};
test_bias[2666:2666] = '{32'h426c6a52};
test_output[2666:2666] = '{32'hc5d25835};
test_input[21336:21343] = '{32'h4227ec85, 32'h428328f4, 32'h428cba74, 32'h40a7e167, 32'hc1591b13, 32'hc175fd4c, 32'hbf3b240b, 32'h4202a918};
test_weights[21336:21343] = '{32'h42083307, 32'hc23d1c9b, 32'h42a30be3, 32'h426ba62a, 32'h4215f75c, 32'hc2b65ee1, 32'hc292270b, 32'hc28c977d};
test_bias[2667:2667] = '{32'h423456a4};
test_output[2667:2667] = '{32'h453fdcf0};
test_input[21344:21351] = '{32'hc1fa5c38, 32'h3f0ea7fc, 32'hc23bcef2, 32'hc1885c1b, 32'h423f8228, 32'hc28d6434, 32'hc20ca481, 32'hc0bf3d54};
test_weights[21344:21351] = '{32'hc2adbd6f, 32'h40d9d199, 32'h3f5577aa, 32'h41a7f040, 32'hc1532ea1, 32'hc258a87a, 32'h4201bccd, 32'hc0ef1fd1};
test_bias[2668:2668] = '{32'h4292e9cf};
test_output[2668:2668] = '{32'h458ca33b};
test_input[21352:21359] = '{32'hc203973d, 32'h429824ce, 32'h42013652, 32'hc2b900da, 32'hc2a1d0ba, 32'h42b4950c, 32'hc20dab14, 32'hc29be95a};
test_weights[21352:21359] = '{32'hc1c6dbff, 32'hc2026662, 32'hc1bac972, 32'hc2af96e2, 32'hc2c6da65, 32'hc1c86ad0, 32'hc229917b, 32'hc2b0563b};
test_bias[2669:2669] = '{32'h4231f840};
test_output[2669:2669] = '{32'h469b8484};
test_input[21360:21367] = '{32'h419d916d, 32'hc2220cf2, 32'hc2286e5a, 32'h425719bb, 32'h42b0e314, 32'hc0ea9590, 32'h42b2a056, 32'h3fb8ceda};
test_weights[21360:21367] = '{32'h421fbd1d, 32'hc1a12e77, 32'h40a4e54e, 32'h4231709b, 32'hc0d59dae, 32'h424cf208, 32'hc20ef1ee, 32'hc2b5ed41};
test_bias[2670:2670] = '{32'hc1a70174};
test_output[2670:2670] = '{32'hc406aa5f};
test_input[21368:21375] = '{32'h40ae8164, 32'hc168dbd5, 32'h42c6e446, 32'h42bf78ae, 32'hc23971b8, 32'hc2a4353e, 32'hc2001f90, 32'h4276fdaa};
test_weights[21368:21375] = '{32'h42bb2183, 32'h422b968f, 32'h42a1e34e, 32'hc2c6c84e, 32'hc2c4ec1f, 32'hc2c2b1e1, 32'h42a749ef, 32'hc2bd4288};
test_bias[2671:2671] = '{32'h3f4b94ca};
test_output[2671:2671] = '{32'h45197f8a};
test_input[21376:21383] = '{32'hc07f3409, 32'hc1409570, 32'h4215096c, 32'hc18ae685, 32'hc20619f4, 32'hc1378cbb, 32'hc2584685, 32'h429d7da6};
test_weights[21376:21383] = '{32'hc2a9f6d2, 32'hc1bb1201, 32'hc2904f9c, 32'h42309a05, 32'h411d6667, 32'hc2b6c128, 32'h4198f068, 32'h421e117a};
test_bias[2672:2672] = '{32'h4243defe};
test_output[2672:2672] = '{32'h412ded14};
test_input[21384:21391] = '{32'hc214b3f5, 32'h42a7d278, 32'h42093b59, 32'hc1ed3d92, 32'hc27c1b6d, 32'h42af4b36, 32'h419e9168, 32'hc28d1ed4};
test_weights[21384:21391] = '{32'h4223816e, 32'h4199bf6f, 32'hc2347c5f, 32'h41fb1634, 32'hc2701986, 32'hc1da2338, 32'h42291a6d, 32'hc243c6d3};
test_bias[2673:2673] = '{32'hc1ec565b};
test_output[2673:2673] = '{32'h454c5780};
test_input[21392:21399] = '{32'h424d3089, 32'h429daf8a, 32'hc2b1d323, 32'hc0945b9c, 32'hc294dc49, 32'hc29ec049, 32'hc2a34b8f, 32'h410639c0};
test_weights[21392:21399] = '{32'hc21b165b, 32'hc1642a2e, 32'hc0e6895a, 32'h4287601b, 32'hc1c0676b, 32'h41e1693c, 32'hc29988d6, 32'hc141cde6};
test_bias[2674:2674] = '{32'hc1d27771};
test_output[2674:2674] = '{32'h4535b065};
test_input[21400:21407] = '{32'hc1bd7d5b, 32'h4264eec3, 32'hc2990166, 32'hc2b3aede, 32'h42a488eb, 32'h41987a89, 32'h429c9c66, 32'hc270a359};
test_weights[21400:21407] = '{32'h40a4cc55, 32'h408686da, 32'h425e7555, 32'hc2842bd0, 32'h41ca718e, 32'hc1355d63, 32'hc0c1d93d, 32'h41ce04be};
test_bias[2675:2675] = '{32'hc0b15889};
test_output[2675:2675] = '{32'h44ccb9c2};
test_input[21408:21415] = '{32'hc1b76e79, 32'hc28abd0c, 32'h41d7e4c7, 32'hc13614a3, 32'hc24c512d, 32'hc2711d99, 32'hc1a3156f, 32'hc2c56d46};
test_weights[21408:21415] = '{32'h42a10cf8, 32'h426a64ca, 32'hc2834f7a, 32'h423aceab, 32'h41aa75ee, 32'h42a6a151, 32'h41880936, 32'hc29d6b51};
test_bias[2676:2676] = '{32'h3f18e03f};
test_output[2676:2676] = '{32'hc5d7ab91};
test_input[21416:21423] = '{32'h42b5ad33, 32'h41c83a52, 32'hc2adc7a4, 32'h428039dd, 32'hc15c23b9, 32'h428f2f6b, 32'h42697d7d, 32'h4262ae72};
test_weights[21416:21423] = '{32'h41e191b4, 32'h41ac06ba, 32'hc2c37a16, 32'h405d5e21, 32'hc28398b4, 32'hc1a18600, 32'hc2994481, 32'h4255011b};
test_bias[2677:2677] = '{32'h422a3230};
test_output[2677:2677] = '{32'h461a1228};
test_input[21424:21431] = '{32'h4204648c, 32'hc2a46fd1, 32'h41ebab3d, 32'h4292cb4c, 32'h41ef477c, 32'h42ab5285, 32'hc0e017fc, 32'h429f4d4f};
test_weights[21424:21431] = '{32'h428cadc1, 32'hc21609bc, 32'hc281ab58, 32'h4291640e, 32'hc1058465, 32'hc2b6d7bb, 32'hc21a0103, 32'hc2194fb5};
test_bias[2678:2678] = '{32'hc229a2a0};
test_output[2678:2678] = '{32'hc5014b93};
test_input[21432:21439] = '{32'hc2411277, 32'hc2ad6fa6, 32'h40138676, 32'h425aeed3, 32'h42557ece, 32'hc214dbce, 32'hc2c0fc99, 32'hc249536b};
test_weights[21432:21439] = '{32'h42b06203, 32'h42916d78, 32'h41e4d50e, 32'h420dc772, 32'hc121383f, 32'hc258140a, 32'hc2434cb8, 32'h4265c752};
test_bias[2679:2679] = '{32'h428ff234};
test_output[2679:2679] = '{32'hc5a23ff3};
test_input[21440:21447] = '{32'h42983cb7, 32'hc19ee9d0, 32'hc29e9fb9, 32'hc287b1aa, 32'h42a783d0, 32'h42b7526d, 32'h42c04c15, 32'h4238b588};
test_weights[21440:21447] = '{32'hc1f7e39f, 32'h424dd6ab, 32'hc1f152ab, 32'hc24c9f7f, 32'h41861a52, 32'hc1ecbcd2, 32'hc2743dc2, 32'h42c3d42a};
test_bias[2680:2680] = '{32'h42030a5a};
test_output[2680:2680] = '{32'hc30eb47c};
test_input[21448:21455] = '{32'h4175ec87, 32'hbf222865, 32'h41e13b10, 32'hc063b5bc, 32'h42155b34, 32'h4285b193, 32'hc295d69c, 32'hc2597a83};
test_weights[21448:21455] = '{32'hbef9fa96, 32'h421f9e33, 32'h429f7848, 32'h4283c72f, 32'hc2ae0f84, 32'hc1882be9, 32'hc2bfa442, 32'h422d60a2};
test_bias[2681:2681] = '{32'hbf767aa1};
test_output[2681:2681] = '{32'h4516b684};
test_input[21456:21463] = '{32'h427e0d04, 32'hc1e60813, 32'h42b56bfa, 32'hc2987884, 32'hc2b1dfd4, 32'hc1aea42b, 32'hc239de1e, 32'hc272a065};
test_weights[21456:21463] = '{32'hc18f5eb4, 32'hc0d9ce2c, 32'hc0db7d05, 32'h41c09297, 32'h42bf94c8, 32'h421f7be6, 32'h4206235c, 32'h428b930e};
test_bias[2682:2682] = '{32'hc2886f33};
test_output[2682:2682] = '{32'hc691b220};
test_input[21464:21471] = '{32'hc2181153, 32'h4206ba28, 32'h429e192a, 32'hc2b2ac7e, 32'h426c9ace, 32'hc20f9b54, 32'hc11933dd, 32'h426cbca7};
test_weights[21464:21471] = '{32'h428a7caa, 32'hbe0cf976, 32'hc20322b4, 32'hc26022bd, 32'h41a3cc54, 32'hc1ae07a7, 32'hc2812573, 32'h4124a1a1};
test_bias[2683:2683] = '{32'h41f175f3};
test_output[2683:2683] = '{32'h453d2dad};
test_input[21472:21479] = '{32'hc2a514dd, 32'hc1c72c78, 32'hc1ade126, 32'h408f67db, 32'h426d1a25, 32'h40e78db3, 32'h42a9db22, 32'hc226e21c};
test_weights[21472:21479] = '{32'h4123c323, 32'h42722e5b, 32'h4240d62a, 32'h41cbef57, 32'hc118500b, 32'hc2a241fa, 32'h4107b150, 32'hc148301d};
test_bias[2684:2684] = '{32'hc29270e3};
test_output[2684:2684] = '{32'hc54c411b};
test_input[21480:21487] = '{32'hc20ab7c9, 32'h3f70496e, 32'hc26a7ec5, 32'h42b477c6, 32'hc2ad8399, 32'hc26cec08, 32'h423c0e7b, 32'h427261ad};
test_weights[21480:21487] = '{32'hc298520d, 32'hc2c1cf82, 32'hc1d36202, 32'hc299ada2, 32'h42abead0, 32'hc2244d01, 32'hc221d83b, 32'hc28e66ac};
test_bias[2685:2685] = '{32'h3e8731c1};
test_output[2685:2685] = '{32'hc65bed0e};
test_input[21488:21495] = '{32'h429c5864, 32'hc2214820, 32'h42379933, 32'h4244aabc, 32'h4298cd90, 32'h420bcebf, 32'hc23b8c92, 32'hc20b9e10};
test_weights[21488:21495] = '{32'hc1cbfb3f, 32'h429cf8f3, 32'h41d6db00, 32'hc29b3969, 32'h428a548b, 32'hbf5dab82, 32'h414eca70, 32'hc1f629ae};
test_bias[2686:2686] = '{32'hc2c4a35e};
test_output[2686:2686] = '{32'hc504544e};
test_input[21496:21503] = '{32'hc08e5f32, 32'h420933f9, 32'hc1b76eb8, 32'h42ba6766, 32'hc1cea063, 32'h425b59cc, 32'hc230e913, 32'h4286302b};
test_weights[21496:21503] = '{32'hc23603f3, 32'h4228d549, 32'hc28107c7, 32'h42728946, 32'hc0dc7de4, 32'hc267faa2, 32'hc1d2cd00, 32'h4297b1d7};
test_bias[2687:2687] = '{32'h3ffdd34e};
test_output[2687:2687] = '{32'h463c0ab2};
test_input[21504:21511] = '{32'hc18da93a, 32'hc2565706, 32'h428c29c9, 32'hc0c066a4, 32'h421e9acd, 32'hc1323213, 32'hc13a448d, 32'hc2a7027d};
test_weights[21504:21511] = '{32'h4034dd47, 32'h4155fac2, 32'h41f54a9e, 32'h41a994bd, 32'hc2a8df79, 32'hc293f9e8, 32'h42c35cc9, 32'h41e70f7f};
test_bias[2688:2688] = '{32'h40b585e8};
test_output[2688:2688] = '{32'hc5966529};
test_input[21512:21519] = '{32'hc29b60fd, 32'hc27bd23e, 32'h42951ab1, 32'hc292ec8f, 32'h41fafcd5, 32'hc1e48fbd, 32'h42062fd0, 32'hbfd1fe9b};
test_weights[21512:21519] = '{32'h4298eedf, 32'hc170696d, 32'h41065f5e, 32'h41d28df3, 32'hc2becc29, 32'hc1f12e68, 32'h429e4814, 32'h4262e296};
test_bias[2689:2689] = '{32'h414b41a6};
test_output[2689:2689] = '{32'hc5b71943};
test_input[21520:21527] = '{32'h40cdf194, 32'hc269ff6f, 32'hc259be9c, 32'hc29e80bf, 32'hc16011e8, 32'h4027a981, 32'hc230be00, 32'hc1b4dc1c};
test_weights[21520:21527] = '{32'hc2b1ded8, 32'h42816edf, 32'hc20e9648, 32'hc243bbcf, 32'h404e69bf, 32'hc2815ea5, 32'hc279095b, 32'hc0d34ed1};
test_bias[2690:2690] = '{32'h429401d8};
test_output[2690:2690] = '{32'h4583df1e};
test_input[21528:21535] = '{32'h42448917, 32'hc2a7b097, 32'h415aa94a, 32'hc20bf180, 32'h4214186e, 32'hc2bf3eff, 32'h425e9b4d, 32'h424304e0};
test_weights[21528:21535] = '{32'h42b78a7b, 32'h42451fce, 32'h420401a9, 32'h42aa67f8, 32'hc263bfaf, 32'h42bafd5f, 32'h41e34a0f, 32'hc276d438};
test_bias[2691:2691] = '{32'h42a334ba};
test_output[2691:2691] = '{32'hc6634b9e};
test_input[21536:21543] = '{32'h42a16fe5, 32'hc2c2b4c5, 32'hc202e97c, 32'hc2b766b2, 32'h41ccd13f, 32'hc2aa8cd4, 32'hc20003db, 32'hc21eef3d};
test_weights[21536:21543] = '{32'hc2866101, 32'h425bf172, 32'h40fb2b1b, 32'hc22fe148, 32'h426590e9, 32'h423964fd, 32'h42169098, 32'hc2596760};
test_bias[2692:2692] = '{32'hc2003510};
test_output[2692:2692] = '{32'hc605c5db};
test_input[21544:21551] = '{32'h42b1ceab, 32'hc218410b, 32'hc29d305d, 32'hc14a98b2, 32'h41a47416, 32'hc1853c88, 32'h42c2ffe8, 32'h429fc887};
test_weights[21544:21551] = '{32'hc217d992, 32'hc29299c0, 32'hc26ece06, 32'hc29c952a, 32'h42b07584, 32'hc1a97660, 32'hc23e97d8, 32'h42a87b65};
test_bias[2693:2693] = '{32'hc21b664c};
test_output[2693:2693] = '{32'h46117ac8};
test_input[21552:21559] = '{32'h4287fae1, 32'h41e5323a, 32'hc20119b8, 32'hc2c77744, 32'hc245ce05, 32'hc280075d, 32'hc266463c, 32'h4281d3f9};
test_weights[21552:21559] = '{32'h4250d855, 32'h428b178f, 32'h42193094, 32'h426db263, 32'h42ac6e0b, 32'hc29542e2, 32'hc2a03584, 32'h42765fb0};
test_bias[2694:2694] = '{32'hc28f668a};
test_output[2694:2694] = '{32'h45e83e45};
test_input[21560:21567] = '{32'hc2827735, 32'hc29a994a, 32'h42be9fef, 32'h428b00ca, 32'hc2bbb19a, 32'hc29d243f, 32'hc035a6b9, 32'h419ee73b};
test_weights[21560:21567] = '{32'h42c4735f, 32'h42b820fe, 32'hc2a333cb, 32'hc19c250d, 32'h417e73e0, 32'hc1777b7b, 32'hc2a64626, 32'h41953b59};
test_bias[2695:2695] = '{32'h42b21a48};
test_output[2695:2695] = '{32'hc6adbf9d};
test_input[21568:21575] = '{32'hc2278cc2, 32'h42160773, 32'hc19b9c35, 32'h42b3a49f, 32'hc2b9e56d, 32'h42a9113b, 32'h42727820, 32'hc17e2ebd};
test_weights[21568:21575] = '{32'h42408c2d, 32'h428cbb3b, 32'hc0de21fd, 32'h425c3071, 32'hc225e73e, 32'hc2a18293, 32'h42b3a9dc, 32'hc2055191};
test_bias[2696:2696] = '{32'h42483a2d};
test_output[2696:2696] = '{32'h4608cf58};
test_input[21576:21583] = '{32'h425a9a04, 32'hc223365e, 32'h418785e9, 32'hc2af1612, 32'h424f4228, 32'hc29e37ec, 32'hc259ca5c, 32'hc2ae6422};
test_weights[21576:21583] = '{32'h42868992, 32'h420ce698, 32'h41edfc54, 32'h42b59382, 32'h42527eef, 32'hc20f102e, 32'h41f9eaa6, 32'hc24bf50d};
test_bias[2697:2697] = '{32'h428bcb9d};
test_output[2697:2697] = '{32'h4545e271};
test_input[21584:21591] = '{32'h42a03439, 32'h425145bc, 32'hc279a291, 32'hc284bdcc, 32'hc20a1561, 32'hc25e4d38, 32'hc09e3015, 32'h4293522e};
test_weights[21584:21591] = '{32'h42a46355, 32'h423b4af4, 32'h42a68df0, 32'h42901589, 32'hc1f1564b, 32'h4200f069, 32'hc1848ce6, 32'hc1c6a570};
test_bias[2698:2698] = '{32'hc289a65b};
test_output[2698:2698] = '{32'hc55b7231};
test_input[21592:21599] = '{32'h408cb7e0, 32'hc2873dfc, 32'h422b8b30, 32'h41a895a1, 32'hc24a3e6b, 32'hc2b11d34, 32'h42b37694, 32'hc26f6bcd};
test_weights[21592:21599] = '{32'h420106b0, 32'hc2a750b4, 32'h42a5564d, 32'hc1c81926, 32'h42060957, 32'h4053edac, 32'h421546bf, 32'h42274da8};
test_bias[2699:2699] = '{32'h4284c0cc};
test_output[2699:2699] = '{32'h45f1e96b};
test_input[21600:21607] = '{32'hc225b384, 32'hc21a45ef, 32'h4121bd24, 32'h4285724e, 32'hc2222066, 32'hc21ab6cb, 32'hc23f454e, 32'h41bac4d3};
test_weights[21600:21607] = '{32'h42099454, 32'h42139a2c, 32'h413703e3, 32'h4223fa0e, 32'h42c1021a, 32'hc1d10b16, 32'hc272e6e9, 32'hc234a9b0};
test_bias[2700:2700] = '{32'hc2ae5a91};
test_output[2700:2700] = '{32'hc48df891};
test_input[21608:21615] = '{32'h41a0f236, 32'h41c23953, 32'hc2a2d270, 32'hc247ba46, 32'h41c12d51, 32'h42985411, 32'hc267fe28, 32'h42ad9c2c};
test_weights[21608:21615] = '{32'hc0689385, 32'h4215211c, 32'hc195b99a, 32'h42211994, 32'h4126b048, 32'h41c6646e, 32'h41cde777, 32'h42833cff};
test_bias[2701:2701] = '{32'h425ac134};
test_output[2701:2701] = '{32'h45d2b85f};
test_input[21616:21623] = '{32'h3f8442fa, 32'hc21b20cb, 32'h41083ec7, 32'h42aad7a7, 32'h42bb127e, 32'h41634ef3, 32'h41b36110, 32'h428e81a5};
test_weights[21616:21623] = '{32'h425f0560, 32'h42a063fa, 32'hc1a593a1, 32'h42af9fd4, 32'h42a284c7, 32'hc2b67347, 32'hc24e0aa8, 32'hbfa7a549};
test_bias[2702:2702] = '{32'h3cec5943};
test_output[2702:2702] = '{32'h4611c291};
test_input[21624:21631] = '{32'hc2bef596, 32'hc079ab14, 32'hc20fe3be, 32'hc1c8d974, 32'hc290ca7c, 32'hc25370f5, 32'h42948ce8, 32'h42bf4611};
test_weights[21624:21631] = '{32'h423a5625, 32'hc261564f, 32'hc28d1ef3, 32'hc2ac744d, 32'hc1bed95f, 32'hc2a4612d, 32'h4127c639, 32'h4250643d};
test_bias[2703:2703] = '{32'hc05d2c4b};
test_output[2703:2703] = '{32'h4640420a};
test_input[21632:21639] = '{32'h423bbe2b, 32'h42c0da41, 32'h42a866e9, 32'hc23473fe, 32'hc258430e, 32'hc25ec7f6, 32'hc272e5c7, 32'hc2280ca7};
test_weights[21632:21639] = '{32'hc2b7193e, 32'hc1154d42, 32'h42a23298, 32'hc1d3ac3b, 32'h41b9832c, 32'h42c391a1, 32'h420c98ce, 32'hc237b590};
test_bias[2704:2704] = '{32'h429184fb};
test_output[2704:2704] = '{32'hc57a6763};
test_input[21640:21647] = '{32'hc285c58a, 32'h429d6fec, 32'h41cb68b6, 32'hc2a1a054, 32'h42bbacc4, 32'h428d5d92, 32'h42504c10, 32'hc20167f1};
test_weights[21640:21647] = '{32'hc1ccc2f3, 32'hc0bb00c3, 32'hc29d16e0, 32'h3fc1cd04, 32'h4297dc73, 32'hc2ad3d27, 32'h41a313c0, 32'h40b31da2};
test_bias[2705:2705] = '{32'hc213f27a};
test_output[2705:2705] = '{32'h4474a440};
test_input[21648:21655] = '{32'hc28237c5, 32'hc2c3df07, 32'hc04df407, 32'hc2847d90, 32'hc1b29e3a, 32'h420759fd, 32'h4289584f, 32'h41cebf58};
test_weights[21648:21655] = '{32'h406a8c6b, 32'h4220d8b7, 32'h41fc8877, 32'hc2a9c419, 32'hc29c5980, 32'hc289516b, 32'h42be5392, 32'h3f1483f4};
test_bias[2706:2706] = '{32'hc26fcac7};
test_output[2706:2706] = '{32'h45e2c856};
test_input[21656:21663] = '{32'hc280278a, 32'hc12594e7, 32'h42af8599, 32'hc19f625a, 32'h42af442e, 32'h421210e9, 32'hc28cae95, 32'hc22a65a8};
test_weights[21656:21663] = '{32'h42bdafe3, 32'h4259f3fa, 32'h4261582e, 32'hc072bb36, 32'h410ca18e, 32'hc25ac80f, 32'hc1a71343, 32'h428d4b20};
test_bias[2707:2707] = '{32'hc216dec7};
test_output[2707:2707] = '{32'hc58a560a};
test_input[21664:21671] = '{32'h42910583, 32'hc1e8241f, 32'hbf2f46c8, 32'hc21ee169, 32'hc28e4539, 32'hc1dddf67, 32'hc111b02f, 32'hbfdd2ed7};
test_weights[21664:21671] = '{32'h41826c3b, 32'hc237765e, 32'hc292a43c, 32'hc2b9907c, 32'hc2a7a88a, 32'hc1b52b7c, 32'h41cf72cb, 32'hc21ecf58};
test_bias[2708:2708] = '{32'hc1f15625};
test_output[2708:2708] = '{32'h464588a9};
test_input[21672:21679] = '{32'hc06d6b3a, 32'hc24f2ac8, 32'h42a8bfe8, 32'hc1dac8d1, 32'h426ad851, 32'hc1b12645, 32'hc1498108, 32'h429175cd};
test_weights[21672:21679] = '{32'hc1db6644, 32'h41899ca0, 32'hc2a22955, 32'hc28d2e92, 32'hc210ee27, 32'h42b83923, 32'h4068951d, 32'hc230ac05};
test_bias[2709:2709] = '{32'hc2821827};
test_output[2709:2709] = '{32'hc64e17a3};
test_input[21680:21687] = '{32'hbfdde861, 32'h422d92cb, 32'hc26b6090, 32'hc18a382c, 32'h42861b47, 32'h4205717a, 32'h41e1d207, 32'hc166b4ce};
test_weights[21680:21687] = '{32'hc2ae1c18, 32'hc28c35f4, 32'hc2845d6e, 32'h41df8fc5, 32'hc24bfddc, 32'h42a1baf5, 32'h42438e56, 32'hc114956d};
test_bias[2710:2710] = '{32'h41022967};
test_output[2710:2710] = '{32'h44a5152b};
test_input[21688:21695] = '{32'hc29e0037, 32'h425142ca, 32'h425b790f, 32'hc279d3a7, 32'hc29a060f, 32'h42af3f9f, 32'hc291fc11, 32'h42013f75};
test_weights[21688:21695] = '{32'hc2be53cb, 32'h42a1ede8, 32'h41799fe0, 32'h4270c5aa, 32'hc29e53c0, 32'hc17b1b13, 32'hc2a9a415, 32'hc28c2f27};
test_bias[2711:2711] = '{32'hc0173663};
test_output[2711:2711] = '{32'h4688af47};
test_input[21696:21703] = '{32'hc2c13d86, 32'hc2ac6a05, 32'hc29e8b35, 32'hbfb99e39, 32'h420b34ac, 32'hc1acd5ee, 32'h418ed860, 32'h4138940e};
test_weights[21696:21703] = '{32'h4230af18, 32'hc2aed00c, 32'hc2c62c06, 32'hc2a78392, 32'hc283151d, 32'hc18e0865, 32'h41f88859, 32'h413dc19c};
test_bias[2712:2712] = '{32'h421157b5};
test_output[2712:2712] = '{32'h461d67bb};
test_input[21704:21711] = '{32'h423a1715, 32'h42b5a1e0, 32'hc2b86d2e, 32'hc1a424d5, 32'h420f60aa, 32'h429f985c, 32'h42174650, 32'hc2273aa1};
test_weights[21704:21711] = '{32'h40d3e0a4, 32'hc222fc95, 32'hc23b4e1f, 32'h42a89b6a, 32'hc22f1824, 32'hc1ebcba7, 32'h41ebecc1, 32'hc250e77c};
test_bias[2713:2713] = '{32'h40b15b65};
test_output[2713:2713] = '{32'hc4b19d59};
test_input[21712:21719] = '{32'hc195291c, 32'h40d20442, 32'hc0a8c585, 32'hc2a33107, 32'hc24559a9, 32'hc29f9e95, 32'h42a45d88, 32'hc0cf9a03};
test_weights[21712:21719] = '{32'h429ab746, 32'h3f563bc8, 32'hc23400a5, 32'h420a3a03, 32'h4141afd1, 32'hc2473875, 32'h42805a92, 32'hc27c96d3};
test_bias[2714:2714] = '{32'h4274176e};
test_output[2714:2714] = '{32'h459f7b52};
test_input[21720:21727] = '{32'hc2147401, 32'h42080df8, 32'h42c56238, 32'hc21fa168, 32'hc20d4279, 32'hc14783f4, 32'hc22869af, 32'hc2bdce6e};
test_weights[21720:21727] = '{32'hc20e4e71, 32'hc21383e5, 32'hc2508b36, 32'h40ac92ed, 32'hc1a4ac89, 32'h42831e16, 32'hc29b6eb7, 32'h42480013};
test_bias[2715:2715] = '{32'h4231b252};
test_output[2715:2715] = '{32'hc5d4eeb1};
test_input[21728:21735] = '{32'h429a5d55, 32'hc08cd844, 32'h41101ad4, 32'h42b51f32, 32'h42393de9, 32'h42833cab, 32'h426eb58a, 32'hc28279ed};
test_weights[21728:21735] = '{32'h4231cc34, 32'h4233eedc, 32'hc2be19bf, 32'h42431766, 32'h40d1c000, 32'h42b40be8, 32'h426dd482, 32'hc150dc5a};
test_bias[2716:2716] = '{32'h421c212c};
test_output[2716:2716] = '{32'h46884667};
test_input[21736:21743] = '{32'h40badf09, 32'hc18b63d7, 32'h421e46ae, 32'hc20ca676, 32'hc2397071, 32'h419637b0, 32'h4226dca7, 32'hc18165f8};
test_weights[21736:21743] = '{32'hc2b000a8, 32'h42252f9d, 32'hc1fb5246, 32'hc20f4cba, 32'hc26182f5, 32'hc19a21f7, 32'h42b44131, 32'hc25198e5};
test_bias[2717:2717] = '{32'h4185ce2a};
test_output[2717:2717] = '{32'h45b0d879};
test_input[21744:21751] = '{32'hc1e37aed, 32'hc281805a, 32'h423c7be5, 32'h42acdff8, 32'h42a69295, 32'h423fe796, 32'hc24c4395, 32'hc2b79368};
test_weights[21744:21751] = '{32'hc2adef52, 32'hc285dfa3, 32'hc1527450, 32'hc11a254a, 32'hc1b28a44, 32'h4115c3a0, 32'hc2aa47f2, 32'hc23878e0};
test_bias[2718:2718] = '{32'h42b50a00};
test_output[2718:2718] = '{32'h46452125};
test_input[21752:21759] = '{32'hc2a4d82e, 32'h428afd2e, 32'hc2b212c8, 32'hc1dc2344, 32'hc2c54e21, 32'hc1b82d49, 32'hc178ea47, 32'h42916682};
test_weights[21752:21759] = '{32'hc14ed144, 32'hc29202f7, 32'h42afb7ac, 32'h41b4cd15, 32'h41aa579a, 32'h40d66c04, 32'h4293bfbf, 32'h4285e9a1};
test_bias[2719:2719] = '{32'hc2bf3f5c};
test_output[2719:2719] = '{32'hc62d32a7};
test_input[21760:21767] = '{32'h42563208, 32'h42a2fa45, 32'hc29ece78, 32'hc2c5c654, 32'hc1935863, 32'h41d82be0, 32'hc2c507db, 32'h4222b4e5};
test_weights[21760:21767] = '{32'hc18d78d3, 32'hc2226733, 32'hc2583788, 32'h4253c382, 32'h42ab3dc0, 32'hc2c0a879, 32'hc2b14c53, 32'hc2be7b3f};
test_bias[2720:2720] = '{32'hc1be54e2};
test_output[2720:2720] = '{32'hc58df88a};
test_input[21768:21775] = '{32'hc2bcd8a1, 32'h42c74135, 32'h428f50e2, 32'h4232c59b, 32'hc2b3ebea, 32'h42990e7a, 32'h4138b3fc, 32'hc2187219};
test_weights[21768:21775] = '{32'hc2becad2, 32'hc29bb0a1, 32'h428d259f, 32'hc2a98dd8, 32'hc2877ee5, 32'hc223ba89, 32'hc22680dd, 32'hc2181e22};
test_bias[2721:2721] = '{32'hc29b7686};
test_output[2721:2721] = '{32'h45c72cd0};
test_input[21776:21783] = '{32'hc1d366ac, 32'hc291be58, 32'h427af324, 32'hc1bac63d, 32'hc2b3af04, 32'hc287d9b2, 32'hc2992740, 32'hc2bd9b01};
test_weights[21776:21783] = '{32'hc29c1321, 32'hc0e4d8b7, 32'hc267c952, 32'hc1b9517b, 32'hc0ae9fb1, 32'h41f11945, 32'hc21525a5, 32'h40adc923};
test_bias[2722:2722] = '{32'hc2212c72};
test_output[2722:2722] = '{32'h4368047e};
test_input[21784:21791] = '{32'h42802e3f, 32'hc2833c48, 32'hc25d1a8e, 32'h42341805, 32'h42bc75ae, 32'h42340458, 32'h42ae9ec0, 32'h425410c0};
test_weights[21784:21791] = '{32'hc22350a8, 32'hc2ac8ed9, 32'hc21c7439, 32'h428bedbf, 32'h4282653c, 32'hc17a8866, 32'hc25d8824, 32'hbed63495};
test_bias[2723:2723] = '{32'hc145a180};
test_output[2723:2723] = '{32'h460b768c};
test_input[21792:21799] = '{32'hc21451d5, 32'h4189cf04, 32'hc25ccfe7, 32'hc19c823d, 32'h42c4310c, 32'hc24970e9, 32'h41c18b55, 32'hc1fc3ba7};
test_weights[21792:21799] = '{32'hc22b5b64, 32'h3f27eff6, 32'h41cb16ed, 32'h4284e993, 32'hc2044e70, 32'h420589ac, 32'h42c4fc4c, 32'h3f86ce00};
test_bias[2724:2724] = '{32'h41867590};
test_output[2724:2724] = '{32'hc564d39a};
test_input[21800:21807] = '{32'h4209b23a, 32'h41cd5610, 32'h428a20c5, 32'h422fb06b, 32'hc26f3d90, 32'hc2076f00, 32'hc1b341cc, 32'hc22000a1};
test_weights[21800:21807] = '{32'hc1f1c351, 32'hc2733bdc, 32'h42148dec, 32'hc229ce24, 32'hc2a3ca96, 32'hc16d630f, 32'h42476edf, 32'h428de841};
test_bias[2725:2725] = '{32'h41b47302};
test_output[2725:2725] = '{32'hc3d87cb4};
test_input[21808:21815] = '{32'hc1df2756, 32'hbfe778b6, 32'h422682d3, 32'hc22aecc5, 32'h42b4d180, 32'h4270821e, 32'h42712018, 32'hc1abebd3};
test_weights[21808:21815] = '{32'hc296b1ea, 32'h41896257, 32'hc0854385, 32'hc28ee268, 32'h4264ef5e, 32'hc0c81ccd, 32'h41ab16a1, 32'hc2ac8690};
test_bias[2726:2726] = '{32'hc230c2c9};
test_output[2726:2726] = '{32'h4648bd99};
test_input[21816:21823] = '{32'hc10feef6, 32'h408ab8c0, 32'h428986d5, 32'h420d0d3b, 32'hc29945e2, 32'hc271793a, 32'h426827fb, 32'hc296098c};
test_weights[21816:21823] = '{32'h42993c9c, 32'h426f1585, 32'hc2375eef, 32'h40cc488d, 32'h4239ccac, 32'hc2ac7b36, 32'h40438f0a, 32'hc2126aec};
test_bias[2727:2727] = '{32'h429ce55d};
test_output[2727:2727] = '{32'h44a15e0d};
test_input[21824:21831] = '{32'h4212c2d6, 32'h425daf26, 32'hc192eac9, 32'h42a80bc2, 32'h429ceb5f, 32'h414f8a4c, 32'h42b4dca4, 32'hc2754d27};
test_weights[21824:21831] = '{32'hc12faac4, 32'h4295c832, 32'h42ab5391, 32'hc15566db, 32'hc1ccceaf, 32'h4286d583, 32'hc29a45ea, 32'hc24f3cff};
test_bias[2728:2728] = '{32'hc28277d9};
test_output[2728:2728] = '{32'hc5767d06};
test_input[21832:21839] = '{32'h421dddb6, 32'hc1632fc1, 32'h4246fcfb, 32'hc1830df2, 32'h42a377fa, 32'hc1c1a498, 32'hc21396e6, 32'hc25b8650};
test_weights[21832:21839] = '{32'h418e45f2, 32'hc259ec64, 32'h4293ad1a, 32'hc27ebea0, 32'h42bc166d, 32'h42bc6157, 32'hc2a0c024, 32'h41ce41d5};
test_bias[2729:2729] = '{32'h4253659d};
test_output[2729:2729] = '{32'h464e48db};
test_input[21840:21847] = '{32'h427341ce, 32'hc229a645, 32'h41d3974e, 32'h41e4d823, 32'hc10ae68a, 32'hc28b154f, 32'hc18ff6ea, 32'h42b1b841};
test_weights[21840:21847] = '{32'h428ceb69, 32'h429a55df, 32'h42b3f284, 32'hc2367a2e, 32'hc1946e04, 32'hbd8de70b, 32'h425b2d4c, 32'hc255f56f};
test_bias[2730:2730] = '{32'hc0c462d7};
test_output[2730:2730] = '{32'hc55a48e5};
test_input[21848:21855] = '{32'hc286abbb, 32'hc2bb034c, 32'hc214f7d9, 32'hc133bd03, 32'hc1612e9f, 32'hc21dea4c, 32'hc1d4e869, 32'h42435ff1};
test_weights[21848:21855] = '{32'hc24386f9, 32'h42a0790e, 32'hc238696f, 32'h42522d59, 32'h426c1e0a, 32'hc22c55e5, 32'h4235f5a7, 32'h40908fe1};
test_bias[2731:2731] = '{32'h41dcb569};
test_output[2731:2731] = '{32'hc5468b73};
test_input[21856:21863] = '{32'hc1f2da5a, 32'hc22de5b5, 32'hc119740a, 32'hc1b32f7a, 32'h4275c540, 32'h415e398e, 32'hc236ef66, 32'h42c29319};
test_weights[21856:21863] = '{32'h41dc395f, 32'hc289c2b1, 32'h4276df1b, 32'h4295e8e4, 32'h41c2aaf2, 32'hc2ab05fd, 32'hc0eb0798, 32'h400a08a9};
test_bias[2732:2732] = '{32'hc1bf2a6e};
test_output[2732:2732] = '{32'h443356ad};
test_input[21864:21871] = '{32'h426f7c24, 32'hc18cc70d, 32'hc180dfd7, 32'hc22b6dc1, 32'h42ab66da, 32'hc2c0cdfe, 32'h429eff03, 32'hc283d307};
test_weights[21864:21871] = '{32'h42662b88, 32'hc29b2b38, 32'h42b49aaf, 32'hc2612ccd, 32'hc2821645, 32'h428b76f9, 32'h41d49de4, 32'hc2b59d38};
test_bias[2733:2733] = '{32'h41730d4c};
test_output[2733:2733] = '{32'h44c61eab};
test_input[21872:21879] = '{32'hc2af83b6, 32'h41eaab42, 32'hc269fe28, 32'h4216e97d, 32'h41c28375, 32'hc2848f5b, 32'h424ff94a, 32'h41879cac};
test_weights[21872:21879] = '{32'h42750c19, 32'h4241d31c, 32'h426a9f64, 32'hc1c0acc3, 32'hc2a144ce, 32'hc11378a8, 32'h40cc361a, 32'hc2025ef9};
test_bias[2734:2734] = '{32'h41eed18f};
test_output[2734:2734] = '{32'hc619acb9};
test_input[21880:21887] = '{32'h42a0f617, 32'hc094aac1, 32'hc23a00ea, 32'hc2c25a1e, 32'hc1c1de7c, 32'hc2805170, 32'hc24bd864, 32'hc29b5778};
test_weights[21880:21887] = '{32'hc283a1a4, 32'hc2b2fed7, 32'hc1f57f2d, 32'hc1de74a4, 32'hc20eac97, 32'hc256c341, 32'h42659124, 32'h42b7dca2};
test_bias[2735:2735] = '{32'h423b3c6a};
test_output[2735:2735] = '{32'hc5c9e90d};
test_input[21888:21895] = '{32'hc1fff91a, 32'hc2a1f87a, 32'hc284081e, 32'hc1a013a4, 32'h428bd4c0, 32'h41346aec, 32'h41c44b9f, 32'h42a57459};
test_weights[21888:21895] = '{32'hc28f5eb8, 32'hc2b33259, 32'hc20fa9ee, 32'hc2c49af3, 32'h42219590, 32'h3eefb47c, 32'hc26ca9cd, 32'h42412266};
test_bias[2736:2736] = '{32'hc2c4e721};
test_output[2736:2736] = '{32'h4695b336};
test_input[21896:21903] = '{32'hc2a07bd6, 32'hc21e3314, 32'hc10bc6b4, 32'hc22c210b, 32'h423bd20e, 32'h40cde262, 32'hc199f49f, 32'hc240f5a9};
test_weights[21896:21903] = '{32'h40d201ea, 32'h421a1a1c, 32'h4292ff34, 32'h4229bdec, 32'hc2a4629d, 32'hc22f5c2f, 32'hc28ec816, 32'h4187c945};
test_bias[2737:2737] = '{32'hc205f12a};
test_output[2737:2737] = '{32'hc5fe524d};
test_input[21904:21911] = '{32'hc2157060, 32'hc234eae8, 32'hc28522aa, 32'h42c4b8d8, 32'h40af782a, 32'hc251ba99, 32'h41a58b29, 32'h42717182};
test_weights[21904:21911] = '{32'hc2325577, 32'hc1df071b, 32'hc2867973, 32'h422f451d, 32'h42893997, 32'hc15a19d4, 32'h4299d72b, 32'h4140f663};
test_bias[2738:2738] = '{32'h42696570};
test_output[2738:2738] = '{32'h466d351f};
test_input[21912:21919] = '{32'hc238729e, 32'hc231b936, 32'hc275e3b1, 32'hc0bdbb55, 32'h42448544, 32'h42b43312, 32'hc1072bd5, 32'h42bb42ce};
test_weights[21912:21919] = '{32'hc1ef779e, 32'hc265a163, 32'h4261788a, 32'hc1b74de0, 32'h41d95f41, 32'hc2566866, 32'hc295a64d, 32'h427721d4};
test_bias[2739:2739] = '{32'hc1977feb};
test_output[2739:2739] = '{32'h455b1254};
test_input[21920:21927] = '{32'h421a0f8a, 32'hc1e424d2, 32'h41177ea4, 32'hc27a347e, 32'hc2932c67, 32'h40e0dd9a, 32'hc2870c87, 32'h425dfa27};
test_weights[21920:21927] = '{32'hc10550e6, 32'hc28c4d18, 32'hc21d1248, 32'h416a75c6, 32'h42c6cd08, 32'hc206c6c7, 32'hc2c4583e, 32'h416001d4};
test_bias[2740:2740] = '{32'h42161b9f};
test_output[2740:2740] = '{32'h438db37c};
test_input[21928:21935] = '{32'hc1ef4ff0, 32'hc2c4115c, 32'h42be48fc, 32'h40c7d575, 32'hc201679f, 32'h41c557e4, 32'hc0c5fb66, 32'hc2c66605};
test_weights[21928:21935] = '{32'h4180152d, 32'h4199ea51, 32'h4282b2bb, 32'h429a4ec5, 32'hbe3d5d68, 32'h40a106c1, 32'hc231cc43, 32'h40e4d472};
test_bias[2741:2741] = '{32'h4286af17};
test_output[2741:2741] = '{32'h45800aaf};
test_input[21936:21943] = '{32'hc2a2158c, 32'h42892aaf, 32'h426594bc, 32'h41c3317e, 32'h415bf73f, 32'hc2c2fc5b, 32'h40deb0af, 32'hc2a58a72};
test_weights[21936:21943] = '{32'h41a6c712, 32'h428c821f, 32'h42936143, 32'h41feb64a, 32'h422042ce, 32'h410d90a0, 32'hc210944f, 32'hc21396a9};
test_bias[2742:2742] = '{32'h42863619};
test_output[2742:2742] = '{32'h4627135a};
test_input[21944:21951] = '{32'h41ed819a, 32'h427f7810, 32'hc23576bc, 32'h41131a7d, 32'hc28c7104, 32'h429647f2, 32'h42b44e2d, 32'hc18eea85};
test_weights[21944:21951] = '{32'h41c7b69a, 32'h426d2de0, 32'h42bb1227, 32'h4185a2a5, 32'hc2c100df, 32'h4249a673, 32'hc1ba50d3, 32'h4290eeaa};
test_bias[2743:2743] = '{32'hc26dfefb};
test_output[2743:2743] = '{32'h45ebe948};
test_input[21952:21959] = '{32'hc1b39ced, 32'h421f4469, 32'h4275ad7e, 32'hc294a09f, 32'hc202a1e1, 32'hc2363c1d, 32'h428043c2, 32'h4084708e};
test_weights[21952:21959] = '{32'h4276b085, 32'h42a1b70e, 32'hc24c0201, 32'h4100fa05, 32'hc1167146, 32'h409103ef, 32'hc21c689b, 32'h42b3b6f1};
test_bias[2744:2744] = '{32'h42490089};
test_output[2744:2744] = '{32'hc5729aa8};
test_input[21960:21967] = '{32'h42424f7b, 32'hc112740a, 32'hc29e3f24, 32'hc2b9394d, 32'h42a01ad7, 32'h42225020, 32'h42551fce, 32'hc1d851f4};
test_weights[21960:21967] = '{32'h42516abe, 32'hc1c037b3, 32'hc2ac827a, 32'hc2b0166a, 32'hc2ad8a71, 32'h42486a3b, 32'hc196518f, 32'hc2295d56};
test_bias[2745:2745] = '{32'h42ab869e};
test_output[2745:2745] = '{32'h464c0942};
test_input[21968:21975] = '{32'hc26da881, 32'hc213be11, 32'h42a8b80d, 32'h426df8b2, 32'h41cff870, 32'hc1279126, 32'hc2b317bc, 32'h42abf49f};
test_weights[21968:21975] = '{32'hc29813bf, 32'hc2a27d2a, 32'h3fe0f92e, 32'h41859925, 32'hc295506a, 32'hc255b8f1, 32'h41d24d39, 32'h42a7ed2e};
test_bias[2746:2746] = '{32'hc18e686d};
test_output[2746:2746] = '{32'h463d797c};
test_input[21976:21983] = '{32'hc2824faf, 32'h42c54e7c, 32'h41985891, 32'h41dc10d8, 32'h42a62e7a, 32'hc28f7dd6, 32'h42478c64, 32'hc28e6517};
test_weights[21976:21983] = '{32'h420c82ae, 32'hc2c3cb3e, 32'h42b480ed, 32'h427fc2d0, 32'hc2c6cded, 32'hc1d857d1, 32'hc21e5cab, 32'hc2984842};
test_bias[2747:2747] = '{32'hc2c7a28d};
test_output[2747:2747] = '{32'hc632c83f};
test_input[21984:21991] = '{32'hc2c26d21, 32'hc2b8ca94, 32'hc2928d4c, 32'h3f8bf91b, 32'hc2854714, 32'hc26cbc28, 32'hc10143c8, 32'h42a12939};
test_weights[21984:21991] = '{32'hc272aa8f, 32'hc26d7b37, 32'h41901920, 32'h4229d0ff, 32'hc10581ac, 32'h42c6f504, 32'hc22a69f2, 32'h416edc8e};
test_bias[2748:2748] = '{32'hc23ec0cc};
test_output[2748:2748] = '{32'h45c42dc1};
test_input[21992:21999] = '{32'hc28c1e46, 32'hc15eafb1, 32'h41a93b14, 32'hc2a39aa3, 32'h42879d4c, 32'hbff91e97, 32'h4212e17f, 32'h421240ac};
test_weights[21992:21999] = '{32'h41db85d3, 32'hc2a3a0f0, 32'hc20923af, 32'hc2a1ceaf, 32'hc0a09198, 32'hc2a3e308, 32'hbfcb8b26, 32'h4276a0e4};
test_bias[2749:2749] = '{32'hc1942458};
test_output[2749:2749] = '{32'h45de0e34};
test_input[22000:22007] = '{32'hbda325b8, 32'hc28b58ab, 32'hc291290a, 32'h426a491c, 32'h418a2249, 32'h41ed8f16, 32'h4203a89d, 32'hc1b33042};
test_weights[22000:22007] = '{32'h4147bc1e, 32'hc151f1a7, 32'h41503563, 32'h42afe1e9, 32'hc1b2515b, 32'h41ec83d7, 32'hc284bc2a, 32'h419e2c8f};
test_bias[2750:2750] = '{32'h42943123};
test_output[2750:2750] = '{32'h453f3630};
test_input[22008:22015] = '{32'h41fa7ab6, 32'hc16f049a, 32'h41a91c9a, 32'hc2a0e202, 32'hc2a4e9ab, 32'hc2be446c, 32'hc1d6272e, 32'hc273128d};
test_weights[22008:22015] = '{32'h4148d6ea, 32'h4285493d, 32'h41ca6906, 32'hc2b171ca, 32'h4228f255, 32'hc2b428bf, 32'h429cb040, 32'hc252faaf};
test_bias[2751:2751] = '{32'hc2882bb7};
test_output[2751:2751] = '{32'h464e304c};
test_input[22016:22023] = '{32'hc28aa857, 32'h4235ba98, 32'h42bb80c1, 32'hc29a6db7, 32'hc2c65dd5, 32'hc2b567df, 32'hc1675c61, 32'h4297a6d8};
test_weights[22016:22023] = '{32'hc2b2e3f1, 32'h41911973, 32'h4153a04c, 32'h425380fd, 32'hc2368348, 32'hc1fde9f1, 32'hc29898a1, 32'h41459bd7};
test_bias[2752:2752] = '{32'h428c74db};
test_output[2752:2752] = '{32'h46560319};
test_input[22024:22031] = '{32'hc1af9d12, 32'h42a0d9a2, 32'h4017b7f9, 32'h42bec2f6, 32'h42a69341, 32'h409ed23a, 32'hc2bfb8a6, 32'h42a0abd9};
test_weights[22024:22031] = '{32'hc1ae2bcc, 32'hc17ebec6, 32'h42c1102a, 32'h42702b6d, 32'hc2880aad, 32'h400dbe19, 32'hc1386f79, 32'hc2388436};
test_bias[2753:2753] = '{32'hc2a8dd94};
test_output[2753:2753] = '{32'hc547262a};
test_input[22032:22039] = '{32'h4196f039, 32'h42a5df95, 32'hc2201575, 32'hc1551412, 32'hc2ac90a1, 32'h4272e459, 32'h42af53d1, 32'h41accf21};
test_weights[22032:22039] = '{32'hc0e997be, 32'hc2c0b056, 32'hc2bab1a3, 32'hc23c2589, 32'h429cbf65, 32'hc283c391, 32'h421a7443, 32'hc2b1f1a9};
test_bias[2754:2754] = '{32'h42710eb5};
test_output[2754:2754] = '{32'hc64b35c0};
test_input[22040:22047] = '{32'hc21efbfb, 32'hc107f316, 32'h429f2855, 32'hc2c46bdf, 32'h42af7341, 32'hc2bf81cd, 32'h4258e7e3, 32'hc239c4dd};
test_weights[22040:22047] = '{32'hc230e928, 32'h424cd8e4, 32'h41c710bd, 32'hc2436575, 32'h421b0391, 32'hc2b16324, 32'h41acb436, 32'hc292eb74};
test_bias[2755:2755] = '{32'h42b606d0};
test_output[2755:2755] = '{32'h46c0b42d};
test_input[22048:22055] = '{32'h423fa136, 32'h42b4ba2c, 32'hc27555c6, 32'hc1aab983, 32'h42b50587, 32'hc2c2e24a, 32'hc14a33f9, 32'h427c6e51};
test_weights[22048:22055] = '{32'h429828e7, 32'hc29f8b42, 32'h4254cdd6, 32'hc29b2183, 32'hc2725c7c, 32'hc15d92bf, 32'hc185ce9f, 32'h3f8bbfdd};
test_bias[2756:2756] = '{32'hc21750b0};
test_output[2756:2756] = '{32'hc60d9e90};
test_input[22056:22063] = '{32'h421597e2, 32'h423519be, 32'h42be7819, 32'h426f1b33, 32'hc28e933d, 32'h4285e570, 32'h42b68853, 32'h42afaf26};
test_weights[22056:22063] = '{32'hc2b554a5, 32'hc21deb13, 32'hc2b5166b, 32'h42c2e6bd, 32'hc253d9d5, 32'h42be8e73, 32'h429dc675, 32'h4274298c};
test_bias[2757:2757] = '{32'h428f34c9};
test_output[2757:2757] = '{32'h46676f27};
test_input[22064:22071] = '{32'hc1e38751, 32'hc2061703, 32'hc23e8fb8, 32'hbfed99bb, 32'hc2aaadc3, 32'h42b62cea, 32'h4170d436, 32'hc271a8fd};
test_weights[22064:22071] = '{32'h428b9f36, 32'h425129fe, 32'hc2067dac, 32'hc286f25c, 32'h403df952, 32'h41132f5e, 32'hc1fec994, 32'hc292e0e8};
test_bias[2758:2758] = '{32'h3f7b4671};
test_output[2758:2758] = '{32'h451e3ab9};
test_input[22072:22079] = '{32'h428a26a6, 32'h42b33041, 32'h425319c6, 32'h41c3dbe9, 32'hc2921674, 32'hc1f97f0e, 32'h41b8caa7, 32'hc2bdcd2e};
test_weights[22072:22079] = '{32'hc1c8d037, 32'h42208a37, 32'hc246b1b1, 32'hc18ed2a9, 32'h42be025c, 32'h42138558, 32'h4208983c, 32'h42af0def};
test_bias[2759:2759] = '{32'hc1ab11fa};
test_output[2759:2759] = '{32'hc68372a7};
test_input[22080:22087] = '{32'hbf8457e1, 32'hc2a77312, 32'hc1ee92dc, 32'h401e7168, 32'h42b3bf50, 32'hc2653b44, 32'h428861b1, 32'h41d25cb5};
test_weights[22080:22087] = '{32'h42bb60cb, 32'h42ba8ebc, 32'hc219bd43, 32'h4256fc1b, 32'h4190a6b3, 32'hc24818c7, 32'h4241c0df, 32'hc1f94a5b};
test_bias[2760:2760] = '{32'hc26fe194};
test_output[2760:2760] = '{32'h439012c4};
test_input[22088:22095] = '{32'h4280cf0e, 32'h40258ef2, 32'h41cadfc6, 32'h4247068e, 32'h421cd275, 32'hc0bac1aa, 32'hc0fd293f, 32'h40bab630};
test_weights[22088:22095] = '{32'hc23dd419, 32'hc288371a, 32'h41e6bf57, 32'hbf8a221e, 32'hc2a7ca30, 32'h42b31abd, 32'hc1e4eae7, 32'hc289b2a4};
test_bias[2761:2761] = '{32'hc24a0aae};
test_output[2761:2761] = '{32'hc5ce0413};
test_input[22096:22103] = '{32'h41e6d3a0, 32'h420fc96f, 32'hc24d4123, 32'h4294dab4, 32'hc2075fce, 32'hc2742911, 32'hc261cad3, 32'hc121fe23};
test_weights[22096:22103] = '{32'h42736c73, 32'h429d3bf2, 32'h423d083a, 32'hc2a0269c, 32'h41d7d305, 32'hc2bf5d56, 32'h42046c54, 32'hc2b3a16d};
test_bias[2762:2762] = '{32'h42271456};
test_output[2762:2762] = '{32'h434eee4f};
test_input[22104:22111] = '{32'hc24a1162, 32'h40b0c17b, 32'hc2ade50d, 32'h40b9d7e7, 32'h4292d335, 32'hc21ec6eb, 32'hc15db219, 32'hc23518a3};
test_weights[22104:22111] = '{32'hc14fc860, 32'hc2313618, 32'hc1ceb287, 32'h3eb1fe77, 32'h4229c133, 32'h42c0ab0f, 32'h424373eb, 32'hbf80097f};
test_bias[2763:2763] = '{32'hc2a84249};
test_output[2763:2763] = '{32'h449a716f};
test_input[22112:22119] = '{32'hc1c11430, 32'h418d4fc7, 32'h4214c7e7, 32'hc1fb0752, 32'hc2965eb9, 32'h42549015, 32'h422edddf, 32'h42b7efc3};
test_weights[22112:22119] = '{32'hc2c2ecd7, 32'h406cb9a5, 32'hc14640da, 32'h4287c2c0, 32'hc2b428a5, 32'h3ffeefa8, 32'h4285353a, 32'h419e130e};
test_bias[2764:2764] = '{32'hc2a3745a};
test_output[2764:2764] = '{32'h46316182};
test_input[22120:22127] = '{32'h421ab4e9, 32'hc210128d, 32'h429b0791, 32'hc29050fc, 32'hc2950f4b, 32'hc28b786b, 32'hc1e42f56, 32'hc216afb0};
test_weights[22120:22127] = '{32'hc0a750fb, 32'h4061da72, 32'hc24be058, 32'h42a7f4fb, 32'hc0c6d4d6, 32'h426d87f6, 32'hc29d9f01, 32'hc2916ad9};
test_bias[2765:2765] = '{32'h3f83f961};
test_output[2765:2765] = '{32'hc60d1798};
test_input[22128:22135] = '{32'h428d973b, 32'h3fcddeb5, 32'h42af29c7, 32'h4207f55a, 32'h42b8840c, 32'hc25a1f87, 32'hc2221589, 32'hc261a01f};
test_weights[22128:22135] = '{32'h429ac80d, 32'h41af4d07, 32'h42479488, 32'hc2b690f0, 32'h42c57155, 32'hc2b519c4, 32'h427e82c0, 32'hc26c6aa5};
test_bias[2766:2766] = '{32'hc298042a};
test_output[2766:2766] = '{32'h46a80519};
test_input[22136:22143] = '{32'hc2938e9c, 32'hc2019247, 32'hc132e111, 32'h42672235, 32'hc249b177, 32'h418cb75e, 32'hc1e5342f, 32'hc192222d};
test_weights[22136:22143] = '{32'h4249c6a7, 32'hc286c314, 32'h4220daf3, 32'hc2239ed4, 32'h41a505a5, 32'hc24c8af9, 32'h427eeaba, 32'hc1e26273};
test_bias[2767:2767] = '{32'h4202ff7e};
test_output[2767:2767] = '{32'hc5ec803e};
test_input[22144:22151] = '{32'h417596e4, 32'h42c591e4, 32'h42b2ae25, 32'hc22d4a85, 32'hc2b7688e, 32'hc27b6c24, 32'h40b46d1a, 32'h41f5cc89};
test_weights[22144:22151] = '{32'hc1075d7d, 32'h42c27282, 32'h409af771, 32'h40a5dd6e, 32'h41ff38d7, 32'h42afc281, 32'hc26ffbb7, 32'hc1e76879};
test_bias[2768:2768] = '{32'h423e9f10};
test_output[2768:2768] = '{32'h4256f2ff};
test_input[22152:22159] = '{32'h42bc1cfe, 32'hc2afe076, 32'hc230a41d, 32'hc2495b97, 32'hc1275b2c, 32'h41b96138, 32'h429aebb5, 32'hc178fee3};
test_weights[22152:22159] = '{32'h42c6a163, 32'h41b1f2da, 32'h426974ba, 32'hc2014bef, 32'hc1819514, 32'hc27d09dd, 32'h42064dce, 32'hc222a78c};
test_bias[2769:2769] = '{32'h4258c1e6};
test_output[2769:2769] = '{32'h4603a96c};
test_input[22160:22167] = '{32'hc0e7eb7c, 32'hc1c4dbcc, 32'hc238e17b, 32'hc2876caa, 32'hc29b6364, 32'h422466e2, 32'h411b2d8c, 32'hc1a6e14c};
test_weights[22160:22167] = '{32'h42a50829, 32'h411357a3, 32'hc27342a4, 32'hc114a3a0, 32'hc1b80af3, 32'h4084bd5a, 32'h42abe661, 32'h42aa9d58};
test_bias[2770:2770] = '{32'hc24bdf57};
test_output[2770:2770] = '{32'h455f8463};
test_input[22168:22175] = '{32'hc2321cdc, 32'hc29a83cc, 32'hc25f8201, 32'h42a193ec, 32'h429485ea, 32'h424c4d4a, 32'h42beba66, 32'h42a39708};
test_weights[22168:22175] = '{32'hc24fda33, 32'hc2bcc960, 32'hc28d9a95, 32'h404936a4, 32'hc0fa5802, 32'h41917685, 32'hc2c76278, 32'hc15a9d2f};
test_bias[2771:2771] = '{32'h4194ca92};
test_output[2771:2771] = '{32'h455e644f};
test_input[22176:22183] = '{32'hc1c63667, 32'h421b328a, 32'hc2a470ce, 32'h42054175, 32'hc23e4e49, 32'h4189ae64, 32'hc2a28e70, 32'h40fa3b48};
test_weights[22176:22183] = '{32'hc25ffdbc, 32'hc1cd7589, 32'h411e0f62, 32'hc273feae, 32'h41ccee31, 32'hc2053c4d, 32'h4184cd98, 32'h41979666};
test_bias[2772:2772] = '{32'hc234af39};
test_output[2772:2772] = '{32'hc5ab9ccf};
test_input[22184:22191] = '{32'hc06a96c9, 32'h429f2788, 32'h4269517e, 32'h41c16c4a, 32'h4282218f, 32'hc2a1eb55, 32'h42af6adf, 32'hc12441f3};
test_weights[22184:22191] = '{32'hc2b53bcc, 32'h41e7ad90, 32'h42892893, 32'hc22f625c, 32'h412e555c, 32'h42a9c987, 32'hc239c48d, 32'hc22d06a7};
test_bias[2773:2773] = '{32'hc07ee352};
test_output[2773:2773] = '{32'hc583e401};
test_input[22192:22199] = '{32'hc2b46652, 32'h42b54399, 32'hc10fb5fd, 32'hc13c9db1, 32'hc202d5f5, 32'h425c8004, 32'h4121106c, 32'h425c7b55};
test_weights[22192:22199] = '{32'h4271572f, 32'hc27a834a, 32'hc2838232, 32'h42c6e35b, 32'hc1667840, 32'h419a86e5, 32'h42b374f3, 32'hc2bf2e17};
test_bias[2774:2774] = '{32'hc2be6ec3};
test_output[2774:2774] = '{32'hc664841c};
test_input[22200:22207] = '{32'h413208dc, 32'hc1fa3df3, 32'hc2bb225e, 32'h419f5416, 32'h41ecfcc8, 32'h4268771b, 32'h422f961c, 32'h422d8a99};
test_weights[22200:22207] = '{32'h3f0cec20, 32'hc210a0d6, 32'hc20c9576, 32'h429939e4, 32'hc2a61304, 32'hc27a9688, 32'hc25fda45, 32'hc204e23f};
test_bias[2775:2775] = '{32'h4249632a};
test_output[2775:2775] = '{32'hc579cbda};
test_input[22208:22215] = '{32'h4274ddc4, 32'h4218b6b2, 32'hc236bb79, 32'hc2b7ad7c, 32'h41df39b1, 32'h41a97d8c, 32'h4225e6b1, 32'h410c8405};
test_weights[22208:22215] = '{32'hbfa49e2a, 32'h42c473da, 32'h428c829a, 32'hc2b5ef5e, 32'h420dcd92, 32'hc25b4396, 32'hc2312681, 32'h420dde7c};
test_bias[2776:2776] = '{32'hc1819fe3};
test_output[2776:2776] = '{32'h45ddf46e};
test_input[22216:22223] = '{32'h41b85580, 32'h429324d8, 32'hc2ab7810, 32'hc188502d, 32'h419dc46a, 32'hc2ab4f49, 32'h4225081d, 32'h420d7314};
test_weights[22216:22223] = '{32'hc2b80c06, 32'hc22a3be8, 32'h42b7da44, 32'h40932b49, 32'hc2b84ef3, 32'h4267e8b2, 32'h4254c65f, 32'hc27758a5};
test_bias[2777:2777] = '{32'h4205d0ba};
test_output[2777:2777] = '{32'hc69be22a};
test_input[22224:22231] = '{32'hc28a2e10, 32'h4248017e, 32'hc2aec986, 32'hc13fc09f, 32'hc2b9bc8b, 32'hc17084ed, 32'hc085ad42, 32'hbfb2d348};
test_weights[22224:22231] = '{32'hc07eb9c3, 32'hc1f63914, 32'hc1bbb12a, 32'hc09ef7ef, 32'h42ab3355, 32'hc1fd5787, 32'hc238d884, 32'h41e04569};
test_bias[2778:2778] = '{32'hc0889144};
test_output[2778:2778] = '{32'hc5ca6f64};
test_input[22232:22239] = '{32'hc23cab81, 32'h40d86782, 32'h426309ee, 32'hc24b2caf, 32'h422160ad, 32'hc2afd623, 32'hc25a3dc2, 32'h41ba6bfb};
test_weights[22232:22239] = '{32'hc111b33f, 32'h42c70cd2, 32'h41f5c8f6, 32'h41ff8743, 32'h4277cfae, 32'hc26aaea7, 32'h423e784b, 32'hc2157135};
test_bias[2779:2779] = '{32'h420e3f29};
test_output[2779:2779] = '{32'h45aa44cf};
test_input[22240:22247] = '{32'h42c3a837, 32'hc1abfaef, 32'hc2064b1c, 32'h41d79679, 32'hc295f2dc, 32'h4284ac73, 32'h4079b0a8, 32'hc02ad91a};
test_weights[22240:22247] = '{32'h4229364e, 32'h42860f93, 32'hc0bddc1c, 32'hc1c5180b, 32'hc2921f60, 32'h411d1824, 32'hc258d64c, 32'h425e4107};
test_bias[2780:2780] = '{32'hc207b183};
test_output[2780:2780] = '{32'h45f90039};
test_input[22248:22255] = '{32'hc245485d, 32'hc2075190, 32'hc2c7a7e0, 32'hc27a1fa0, 32'h4263f2ce, 32'hc2bcace0, 32'hc18f869e, 32'h42b962ea};
test_weights[22248:22255] = '{32'hc2833c50, 32'hc2b44ec2, 32'hc1ac5347, 32'h418be722, 32'hc28ad672, 32'hc252d4cf, 32'h42be5660, 32'hc2942326};
test_bias[2781:2781] = '{32'h4284a8d6};
test_output[2781:2781] = '{32'hc3135c05};
test_input[22256:22263] = '{32'hc20886b5, 32'h419c261c, 32'hc168a00a, 32'h42095de6, 32'hc207c573, 32'h41171336, 32'h4289862e, 32'hc2a8530c};
test_weights[22256:22263] = '{32'h42408f96, 32'hc27e655a, 32'hc22d26ec, 32'h42321bff, 32'hc15aed24, 32'h42738420, 32'h40436f80, 32'h429fdfbe};
test_bias[2782:2782] = '{32'h422e10b8};
test_output[2782:2782] = '{32'hc5c086ea};
test_input[22264:22271] = '{32'hc2c11e95, 32'h4248cb9a, 32'hc23c5e0b, 32'hc2353c35, 32'hc1f7ad26, 32'h413d38c0, 32'hc26ea608, 32'hc25e1fe3};
test_weights[22264:22271] = '{32'h41c3d820, 32'hc2584ad0, 32'hc25cdc99, 32'h427532da, 32'hc1552e11, 32'h4293901e, 32'h42b12395, 32'h425d19a6};
test_bias[2783:2783] = '{32'h42acb6d4};
test_output[2783:2783] = '{32'hc63f3712};
test_input[22272:22279] = '{32'hc2876d83, 32'hc1961a3b, 32'h421c18e2, 32'h422edddb, 32'hc2a01ea9, 32'hc1718475, 32'hc0311ae6, 32'h4113b8ac};
test_weights[22272:22279] = '{32'h4249fb73, 32'hc25bf12c, 32'h42bfcc4e, 32'hc1788c1e, 32'h426de367, 32'h4259d95c, 32'h41f88c68, 32'hc25138ec};
test_bias[2784:2784] = '{32'h41ec50d5};
test_output[2784:2784] = '{32'hc5aa3873};
test_input[22280:22287] = '{32'h421cfc97, 32'hc1f66deb, 32'hc26d3228, 32'hc200ef33, 32'hbf101989, 32'h42acdd64, 32'h429092c4, 32'hc2bb4898};
test_weights[22280:22287] = '{32'hc24b4c07, 32'h40fa997c, 32'hc1a8dbe3, 32'h429f1cbc, 32'hc2b588ea, 32'hc2a027f3, 32'h41c9e937, 32'hc2ade5a8};
test_bias[2785:2785] = '{32'h4289a71c};
test_output[2785:2785] = '{32'hc3bfceab};
test_input[22288:22295] = '{32'h41dc4105, 32'hc18df56b, 32'hc2ac92a8, 32'h40dbcd81, 32'h425e24a1, 32'hc2c04c09, 32'hc2679c02, 32'hc2b984ef};
test_weights[22288:22295] = '{32'hc2613798, 32'hc19a75d7, 32'h421e6912, 32'hc1da950c, 32'hc2c52065, 32'hbfe38d1e, 32'h413b9ef1, 32'hc2422af6};
test_bias[2786:2786] = '{32'h42c030e9};
test_output[2786:2786] = '{32'hc5c19b35};
test_input[22296:22303] = '{32'h41a0fc6d, 32'hc2ab8e20, 32'h42c5e117, 32'hc2ae6c25, 32'h40b49185, 32'h422e4849, 32'h42652027, 32'h426491d3};
test_weights[22296:22303] = '{32'h401a51a2, 32'hc25939e6, 32'hc080ad19, 32'hc1bea4a5, 32'hc295680a, 32'h410de6cf, 32'hc26e307f, 32'h42c1ef1a};
test_bias[2787:2787] = '{32'h42c0506a};
test_output[2787:2787] = '{32'h46060901};
test_input[22304:22311] = '{32'h419ae6e3, 32'h42a786ed, 32'hc188537e, 32'h42bf767a, 32'h41e584d7, 32'h429b3a96, 32'h42227b20, 32'h416235c8};
test_weights[22304:22311] = '{32'h41358dc0, 32'h4216c4a6, 32'h405fdf72, 32'hc22881e1, 32'hc2aa6646, 32'h41d5c05a, 32'hc0eea92c, 32'h42820ca3};
test_bias[2788:2788] = '{32'h42ac5e85};
test_output[2788:2788] = '{32'hc3bfc9c6};
test_input[22312:22319] = '{32'hc1c6d69b, 32'hc20578b8, 32'h4277add5, 32'h41e9aff0, 32'hc1d2b815, 32'hc252897e, 32'hc246d116, 32'hc2c3ebca};
test_weights[22312:22319] = '{32'hc2854931, 32'hbefcb9fd, 32'h40b762d8, 32'hc28fd3d9, 32'hc0fcdac1, 32'hc1a8a9c4, 32'h418d647a, 32'h429848a3};
test_bias[2789:2789] = '{32'hc2b20adc};
test_output[2789:2789] = '{32'hc5e06c3d};
test_input[22320:22327] = '{32'hc1bec9a1, 32'hc2b8382b, 32'hc0be72bb, 32'h41dc0842, 32'h428add7b, 32'hc1e0271a, 32'hc2a7d8b8, 32'hc2ae1efb};
test_weights[22320:22327] = '{32'h418de07f, 32'h420c3a3e, 32'h421401c2, 32'hc2b2782d, 32'h42a11015, 32'h40f48c2f, 32'hc2b11360, 32'h41d2bd6b};
test_bias[2790:2790] = '{32'h4159d632};
test_output[2790:2790] = '{32'h45834b7f};
test_input[22328:22335] = '{32'hc132da82, 32'h424ea046, 32'h40e5a2e8, 32'h41707343, 32'h42afea8e, 32'h42c79b26, 32'h42083b02, 32'h3f701483};
test_weights[22328:22335] = '{32'hc2c7b459, 32'hc25c12f2, 32'h42560078, 32'hc229043a, 32'h4228e093, 32'h429c34b7, 32'hc0db6c4a, 32'h422b091e};
test_bias[2791:2791] = '{32'hc2234689};
test_output[2791:2791] = '{32'h461144f2};
test_input[22336:22343] = '{32'hc2aa048b, 32'hc214ac31, 32'h4173bf83, 32'h4231e426, 32'hc206f889, 32'h41a819e5, 32'h42ad4eb6, 32'hc2971df6};
test_weights[22336:22343] = '{32'h425c4101, 32'hc2bb4d18, 32'h42578bd1, 32'h426e62c0, 32'h41840ce4, 32'hc21b5759, 32'h42aa3ac8, 32'hc251f02d};
test_bias[2792:2792] = '{32'h42839724};
test_output[2792:2792] = '{32'h464044f7};
test_input[22344:22351] = '{32'h42a0a256, 32'hc2912237, 32'h42b988ed, 32'hc1da1dd8, 32'h402b205d, 32'h42b39b60, 32'h42bed26b, 32'h42ad941f};
test_weights[22344:22351] = '{32'hc2a1a118, 32'hc2c6b71d, 32'h4299ed3d, 32'h429e2801, 32'hc1d8c659, 32'hc241e62c, 32'hc170cb63, 32'hc09b3491};
test_bias[2793:2793] = '{32'hc273ebcb};
test_output[2793:2793] = '{32'hc42022e4};
test_input[22352:22359] = '{32'hc2959aba, 32'h41b8fc24, 32'hc26c8b32, 32'h41537ac4, 32'h4140b949, 32'h428f1c46, 32'hc1d615ef, 32'h418cbeb0};
test_weights[22352:22359] = '{32'h427793a1, 32'hc2b58495, 32'hc28c28ab, 32'hc2630862, 32'h42bf6f6f, 32'h42a8da1c, 32'hc2365d5d, 32'h412a20cb};
test_bias[2794:2794] = '{32'hc221b6ca};
test_output[2794:2794] = '{32'h45a35289};
test_input[22360:22367] = '{32'h42bda50e, 32'hc2213ea2, 32'h4117d037, 32'hc2b0926b, 32'h3f88e59e, 32'hc1f42693, 32'hc2a2626a, 32'h42bec1a0};
test_weights[22360:22367] = '{32'h42816ef5, 32'h426e78b0, 32'h426aba01, 32'h4242c33f, 32'h42a1f087, 32'hc24e48c7, 32'h428f4a7c, 32'hc24b6a30};
test_bias[2795:2795] = '{32'h42a5fdab};
test_output[2795:2795] = '{32'hc60b91f6};
test_input[22368:22375] = '{32'hc27a7b62, 32'h4247d4cb, 32'hc208c851, 32'hc2ac27cb, 32'hc2be186f, 32'h42b9d1a2, 32'hc2836bbc, 32'h42b3d221};
test_weights[22368:22375] = '{32'h41eb7dc2, 32'h42997641, 32'hc29b75a0, 32'h4294270e, 32'h42abcd67, 32'h4271fb86, 32'hc21fe032, 32'hc297d07b};
test_bias[2796:2796] = '{32'h42202663};
test_output[2796:2796] = '{32'hc603bb5e};
test_input[22376:22383] = '{32'h42b7a822, 32'h41c455d2, 32'hc180e139, 32'h428a6a71, 32'h42b89317, 32'h429871d1, 32'hc1828e14, 32'hc13ae6d5};
test_weights[22376:22383] = '{32'h41ff51ff, 32'h42539a9a, 32'hc2bf1daa, 32'hc28585cb, 32'hc2945a09, 32'hc2a3e8eb, 32'hc27fd4b2, 32'h41895309};
test_bias[2797:2797] = '{32'hc2acf8f0};
test_output[2797:2797] = '{32'hc62ece0b};
test_input[22384:22391] = '{32'hc2c0d43e, 32'h41e218e4, 32'hc21da2ad, 32'hc17081bb, 32'hc2c3a82b, 32'hc2905ed8, 32'hc28197de, 32'hc287ef83};
test_weights[22384:22391] = '{32'hc29ef6d3, 32'hc1db9d8b, 32'h422d1fba, 32'hc201805c, 32'hc290aef9, 32'h42c05363, 32'h4292cdc7, 32'hc2935bc5};
test_bias[2798:2798] = '{32'hc29b8fac};
test_output[2798:2798] = '{32'h45bace15};
test_input[22392:22399] = '{32'h42173865, 32'h419fc348, 32'h42868684, 32'h4227e9fc, 32'hc2457c13, 32'hc1dd3d3c, 32'hc22427d0, 32'hc2b2dff1};
test_weights[22392:22399] = '{32'h42a38060, 32'hc28cab66, 32'h42b8724c, 32'h42978456, 32'h41fbff64, 32'hc0f721b0, 32'hc2bb52db, 32'h42639db6};
test_bias[2799:2799] = '{32'hc2997e8a};
test_output[2799:2799] = '{32'h460355e8};
test_input[22400:22407] = '{32'h42bbaaab, 32'hc21106e4, 32'h42c48d15, 32'h41993363, 32'hc214e26c, 32'h42b91e27, 32'hc1a33aff, 32'hc238a47e};
test_weights[22400:22407] = '{32'hc29f6db2, 32'h429144d2, 32'hc21c8829, 32'hc25332e7, 32'hc2c5959c, 32'h42966fb2, 32'h4078155d, 32'hc107d9be};
test_bias[2800:2800] = '{32'h4182b634};
test_output[2800:2800] = '{32'hc57a1d39};
test_input[22408:22415] = '{32'h42696aa5, 32'hc2159c9a, 32'hc2b42ae1, 32'h426d13e3, 32'h40f46a06, 32'h410f7743, 32'hc23e46ed, 32'hc14e919b};
test_weights[22408:22415] = '{32'h42c4696b, 32'hc22efa5a, 32'h41437b62, 32'h42b74611, 32'h41e1a73f, 32'h4220fe64, 32'h426981d2, 32'hc11eb0a8};
test_bias[2801:2801] = '{32'hc290b6dc};
test_output[2801:2801] = '{32'h46154286};
test_input[22416:22423] = '{32'h42b9d6e9, 32'hc2716a17, 32'h41e54b89, 32'hc281d643, 32'hc2005d01, 32'h423689ab, 32'hc24b1d3a, 32'hc289dd19};
test_weights[22416:22423] = '{32'hc2a3b45f, 32'hc279c763, 32'hc20d99ac, 32'h4278de1c, 32'h42970e74, 32'h425a7694, 32'h42b4d921, 32'h42934705};
test_bias[2802:2802] = '{32'h424d1ffe};
test_output[2802:2802] = '{32'hc6900cbb};
test_input[22424:22431] = '{32'hc1df6336, 32'hc2c4f3ac, 32'h41afeff6, 32'hc2845d7f, 32'hc2a1fe5c, 32'hc294d9d8, 32'hc0af4422, 32'hc1fd8a73};
test_weights[22424:22431] = '{32'h429dce19, 32'hc2aa7a71, 32'h4290b231, 32'h40a5d2d3, 32'hc14e11bd, 32'hc2857d88, 32'hc2147029, 32'h42bc1d52};
test_bias[2803:2803] = '{32'hc29232b9};
test_output[2803:2803] = '{32'h46259b76};
test_input[22432:22439] = '{32'hc2ac8c74, 32'hc2bec470, 32'hc29e1fa5, 32'h3fa5056d, 32'h41abd9af, 32'h410fa104, 32'hc28427e2, 32'hc294fe6e};
test_weights[22432:22439] = '{32'hc200a4fa, 32'hc18e1d27, 32'hc2a55b4a, 32'h42234cee, 32'h42770703, 32'h42bec8d5, 32'h420b9566, 32'hc216ed4f};
test_bias[2804:2804] = '{32'hc2aa6ca2};
test_output[2804:2804] = '{32'h465574cc};
test_input[22440:22447] = '{32'h41d85df4, 32'hc2a6a43a, 32'h416a7e40, 32'hc1c7c461, 32'hbf88c1b8, 32'hc28074cd, 32'h423464d9, 32'hc1e96319};
test_weights[22440:22447] = '{32'hc2c0c354, 32'h41951a21, 32'hc211d937, 32'h425e4859, 32'hc23b2b49, 32'hc2ab24c5, 32'h4227b5cc, 32'hc2bd9fd5};
test_bias[2805:2805] = '{32'hc078af06};
test_output[2805:2805] = '{32'h4580ab5e};
test_input[22448:22455] = '{32'hc19f1eb5, 32'hc21af956, 32'hc25d8c47, 32'hc2a4cde0, 32'hbf365083, 32'hc2a04699, 32'h426a1551, 32'hc29eafb9};
test_weights[22448:22455] = '{32'hc1c02d95, 32'hc2c2e9d8, 32'h410337d1, 32'hc1d9673e, 32'h41d800d6, 32'h4147e007, 32'hc29c1cfb, 32'h4207935c};
test_bias[2806:2806] = '{32'hc2bf3d40};
test_output[2806:2806] = '{32'hc511e713};
test_input[22456:22463] = '{32'hc2a6dbb6, 32'hc1604c7c, 32'h411098b2, 32'h42acc312, 32'h418d0286, 32'h41de3f05, 32'h428876c9, 32'hc28512c7};
test_weights[22456:22463] = '{32'hc03993b1, 32'hc2bf7301, 32'hc295561d, 32'h41bb45e6, 32'h420da6e6, 32'hc1f8f32d, 32'hc0882b2b, 32'h429ea7f5};
test_bias[2807:2807] = '{32'h4286415a};
test_output[2807:2807] = '{32'hc52fa981};
test_input[22464:22471] = '{32'h41e21bc2, 32'hc1f7ca06, 32'hc29c6211, 32'h42866ef6, 32'hc1dbff0e, 32'hc2a1d1de, 32'hc2bbee64, 32'h4241d65b};
test_weights[22464:22471] = '{32'hc26f1b0c, 32'h42c1cda2, 32'h423ec3d4, 32'hc29b16a8, 32'h42a4eb11, 32'h41333f87, 32'h4294efcc, 32'hc2b43497};
test_bias[2808:2808] = '{32'hc18fd475};
test_output[2808:2808] = '{32'hc6dc37fd};
test_input[22472:22479] = '{32'h42581218, 32'hc23e759f, 32'h41b7227f, 32'hc1e09926, 32'hc1b09432, 32'hc2c106df, 32'h42954f94, 32'h418c0080};
test_weights[22472:22479] = '{32'h41eed368, 32'h41bbbe6a, 32'h42af8cd4, 32'hc2c64c59, 32'hc1852f5b, 32'h42bf6814, 32'h429cad6c, 32'h41d03f61};
test_bias[2809:2809] = '{32'h41fc9fb9};
test_output[2809:2809] = '{32'h452c272e};
test_input[22480:22487] = '{32'hc271eb95, 32'h42809d76, 32'h42ace435, 32'hc2c518f0, 32'h414ce01c, 32'hc294a592, 32'hc22c5f68, 32'hc1fcdbb3};
test_weights[22480:22487] = '{32'h425aacb9, 32'h4277a59d, 32'h42900589, 32'hc01ae7c8, 32'h41fc7f9f, 32'h42823fdf, 32'h41b65bde, 32'h418d2f16};
test_bias[2810:2810] = '{32'h420260f5};
test_output[2810:2810] = '{32'h44955d81};
test_input[22488:22495] = '{32'h42afeea7, 32'hc2792637, 32'h41546227, 32'h4239c488, 32'h422fbd9e, 32'h42b942d1, 32'h4260bafe, 32'h42a72b26};
test_weights[22488:22495] = '{32'hc22cd90e, 32'h42ae3c15, 32'hc28e19c3, 32'hc2c5819f, 32'hc22e7926, 32'hc2b653df, 32'hc2297420, 32'hc2b4fd25};
test_bias[2811:2811] = '{32'h4176f5a7};
test_output[2811:2811] = '{32'hc708e664};
test_input[22496:22503] = '{32'h420f154b, 32'h424ca788, 32'h419b48b2, 32'hc17ebabc, 32'h42670375, 32'hbee63815, 32'hc2b5d662, 32'h41dfcc36};
test_weights[22496:22503] = '{32'h41d55f9f, 32'hc14e3b3b, 32'hc1e1611b, 32'hc2c084a1, 32'h4245cc0f, 32'hc15eca19, 32'hc281af54, 32'hc2bd6423};
test_bias[2812:2812] = '{32'hbfcbdd0d};
test_output[2812:2812] = '{32'h45e6d8c6};
test_input[22504:22511] = '{32'hc296775c, 32'h42a15d53, 32'hc2ac43be, 32'hc26cd0be, 32'hc0f8ae84, 32'hc2756e46, 32'h421f5748, 32'h42a62a84};
test_weights[22504:22511] = '{32'h42bf4b9a, 32'h41c31130, 32'h3f7ca4b5, 32'hc21f3a59, 32'h42989b76, 32'hc25eaf49, 32'hc210f5df, 32'h4118f53e};
test_bias[2813:2813] = '{32'hc1a42bb5};
test_output[2813:2813] = '{32'hc448f6d0};
test_input[22512:22519] = '{32'h421f1343, 32'hc1c2a44b, 32'hc2193f7c, 32'hc0a77250, 32'hc2405226, 32'h427719b9, 32'hc295b7e6, 32'h41cd2854};
test_weights[22512:22519] = '{32'h426f4acb, 32'hc2ad47b3, 32'hc0905647, 32'h42bf0595, 32'hc21ff9d2, 32'h4285d59a, 32'hc2adeccf, 32'h40f4a2d4};
test_bias[2814:2814] = '{32'hc2ac9fbf};
test_output[2814:2814] = '{32'h46838903};
test_input[22520:22527] = '{32'hc16fdef1, 32'hc2b1c326, 32'hc22ef4d7, 32'h42854c42, 32'h420678d5, 32'h41514bbb, 32'hc21ef56a, 32'h4200af7a};
test_weights[22520:22527] = '{32'h42b02d07, 32'h42988d0a, 32'h40f227af, 32'hc1c06fdd, 32'hc18940f6, 32'hc20c992d, 32'h41b922e7, 32'hc29332bf};
test_bias[2815:2815] = '{32'h42b0efdd};
test_output[2815:2815] = '{32'hc65ef735};
test_input[22528:22535] = '{32'hc2943c26, 32'hc2532122, 32'h4221abd2, 32'hc1c65073, 32'hc26fbd18, 32'hc28a27c5, 32'hc2c3ea0e, 32'h4230c730};
test_weights[22528:22535] = '{32'hc2b8a844, 32'hc22ce1ea, 32'h42c03f76, 32'h429a8751, 32'h41ddc2ff, 32'hc25561c4, 32'hc229b6f4, 32'hc209e89e};
test_bias[2816:2816] = '{32'h42a68ed4};
test_output[2816:2816] = '{32'h4677665d};
test_input[22536:22543] = '{32'h42aebbc4, 32'h4189dab0, 32'h4060fd0a, 32'hc21228d1, 32'h42a00d36, 32'h42b6010c, 32'hc2ad33d9, 32'hc200cb34};
test_weights[22536:22543] = '{32'hc1fea8f4, 32'h4147958a, 32'h420a1a08, 32'hc018fa5a, 32'h426077a5, 32'hc2a02ee2, 32'hc24956bb, 32'hc1a357d9};
test_bias[2817:2817] = '{32'hc1205b15};
test_output[2817:2817] = '{32'hc314b07c};
test_input[22544:22551] = '{32'h427fcaec, 32'h421884ad, 32'hbeed7e6a, 32'hc1d37d76, 32'hc23ae6e7, 32'hc29e34cb, 32'h429e6d85, 32'hc124002e};
test_weights[22544:22551] = '{32'hc200a37a, 32'h42a96457, 32'h402d8716, 32'h427f6ccc, 32'hc068136a, 32'h419234ff, 32'hc28ade67, 32'h4142063c};
test_bias[2818:2818] = '{32'hc2bfd8d5};
test_output[2818:2818] = '{32'hc5eac91f};
test_input[22552:22559] = '{32'hc2a3d521, 32'h428baf1a, 32'hc1319797, 32'hc274f399, 32'hc277ec14, 32'h4293d210, 32'hc2b946e5, 32'hc2651248};
test_weights[22552:22559] = '{32'h42b90179, 32'hc2149601, 32'h425b22a6, 32'hc2a4b677, 32'h425b0989, 32'hc2949b5e, 32'hc1ac877f, 32'hc268c912};
test_bias[2819:2819] = '{32'hc2525583};
test_output[2819:2819] = '{32'hc6120177};
test_input[22560:22567] = '{32'h42148649, 32'hc294abc6, 32'h426e8ceb, 32'hc2af1cb5, 32'hc17ec3e1, 32'hc22593e3, 32'hc25b4806, 32'hc1387970};
test_weights[22560:22567] = '{32'h428e037e, 32'hc1ac8880, 32'h42855b15, 32'hc24f3ebe, 32'hc28cbdf9, 32'hc1bd6119, 32'h41c7c8ea, 32'hc24e1814};
test_bias[2820:2820] = '{32'h42984149};
test_output[2820:2820] = '{32'h465d28be};
test_input[22568:22575] = '{32'hc27c515c, 32'h42aa8128, 32'h42bd4d8c, 32'h42929b5c, 32'h427bd0ba, 32'hc11af88b, 32'hc1c2f44f, 32'hc2728419};
test_weights[22568:22575] = '{32'hc235a3f4, 32'h412745db, 32'hc23ee5a3, 32'hc21668bf, 32'hc222b8f3, 32'h4245a6ad, 32'h41af4f65, 32'hc2b4b5d1};
test_bias[2821:2821] = '{32'hc28faf70};
test_output[2821:2821] = '{32'hc4d2a4d2};
test_input[22576:22583] = '{32'h41d8aea7, 32'h428308bc, 32'hc2c335a9, 32'hc283252a, 32'h40f5739d, 32'hc2bfd65b, 32'hc1ce4afc, 32'h42aef23f};
test_weights[22576:22583] = '{32'h4289a897, 32'h415cd50d, 32'hc214263b, 32'hc271a356, 32'h4250630f, 32'hc1e5e133, 32'hc2ad1b7a, 32'h4245b7d4};
test_bias[2822:2822] = '{32'hc12f9e18};
test_output[2822:2822] = '{32'h469c9a90};
test_input[22584:22591] = '{32'h423e355c, 32'hc108d0e4, 32'h42b0639c, 32'hc281e0da, 32'hc0d364f4, 32'hc0fea50d, 32'hc1cbceea, 32'hc2a88064};
test_weights[22584:22591] = '{32'hc20c04db, 32'hc2993ab4, 32'hc1b343e2, 32'h41e7ab62, 32'hc27ed516, 32'h4292f17b, 32'hc2b94521, 32'hc28dbbe9};
test_bias[2823:2823] = '{32'h42127070};
test_output[2823:2823] = '{32'h45509229};
test_input[22592:22599] = '{32'hc21f5436, 32'h428fa3ac, 32'h4215a8ad, 32'hc2b00c7b, 32'h42a87a56, 32'hc23c7911, 32'hc247f11c, 32'h429eadad};
test_weights[22592:22599] = '{32'hc18f4610, 32'h4252d726, 32'h426b4de1, 32'hbff9ef15, 32'hc1cd5499, 32'h427115e2, 32'h42b0bbab, 32'hc2549c46};
test_bias[2824:2824] = '{32'h42aa56e1};
test_output[2824:2824] = '{32'hc5d0b8f0};
test_input[22600:22607] = '{32'h42b89bb9, 32'hc0d5b098, 32'h41e18d58, 32'hc2bc0660, 32'h428e48f7, 32'hc26ee90c, 32'h425e1419, 32'h429f0cec};
test_weights[22600:22607] = '{32'h429d3743, 32'h428ebdd1, 32'h42c1a8a1, 32'hc1a0247d, 32'hc15fb79d, 32'hc22b9c79, 32'hc2606dcf, 32'h41f932a3};
test_bias[2825:2825] = '{32'h4207b095};
test_output[2825:2825] = '{32'h46410be4};
test_input[22608:22615] = '{32'h42470eb2, 32'hc279ba85, 32'hc19cca50, 32'h42b77d92, 32'hc1f7bd5b, 32'h41f602f7, 32'h4284ca41, 32'hc2ba85c6};
test_weights[22608:22615] = '{32'hc1f4c827, 32'h42658316, 32'hc2c7fde4, 32'hc181039c, 32'hc2c0756c, 32'hc278e3f5, 32'h42168bac, 32'hc27bfc2f};
test_bias[2826:2826] = '{32'h41715c8f};
test_output[2826:2826] = '{32'h4596f790};
test_input[22616:22623] = '{32'hc25d0849, 32'h42a03ca6, 32'hc2bd31fd, 32'h426c9a22, 32'h420224cc, 32'h42232838, 32'h4265ccee, 32'hc20dde2f};
test_weights[22616:22623] = '{32'h424c67fe, 32'h4124fb92, 32'h422c1cbe, 32'h41a5ba63, 32'hc2c2b729, 32'hc29f4ce6, 32'h41d25741, 32'hc2ad6938};
test_bias[2827:2827] = '{32'hc2bcecef};
test_output[2827:2827] = '{32'hc5d37f2a};
test_input[22624:22631] = '{32'hc2c24288, 32'hc1c6934c, 32'h429608ec, 32'hc2a29dc8, 32'hc24a5782, 32'h42a5629c, 32'hc2796a23, 32'h41a85507};
test_weights[22624:22631] = '{32'h42a975ec, 32'hc1d119d6, 32'hc20cc4b6, 32'h4264fff6, 32'hc2b18313, 32'h4008bc27, 32'h42a20b47, 32'hc2c437f4};
test_bias[2828:2828] = '{32'h429e914e};
test_output[2828:2828] = '{32'hc686bd4a};
test_input[22632:22639] = '{32'hc2ab6759, 32'h422b6eeb, 32'h41788c86, 32'h41f18807, 32'hc1872b8e, 32'hc1aaaa80, 32'h41e11efe, 32'h41fc3e8a};
test_weights[22632:22639] = '{32'h4242e456, 32'hc1a3919e, 32'hc278c26a, 32'h42793361, 32'hc1f30b7a, 32'hc1b87737, 32'hc2555731, 32'hc249e784};
test_bias[2829:2829] = '{32'hc217b8b6};
test_output[2829:2829] = '{32'hc5c3b176};
test_input[22640:22647] = '{32'hc130c406, 32'hc2bd927f, 32'h4285e245, 32'h42c1b84f, 32'hc200537b, 32'hc292e39b, 32'h41ef33d2, 32'h42c39d39};
test_weights[22640:22647] = '{32'hc25b8d13, 32'hc2b67311, 32'hc2c10a2d, 32'hc119ed94, 32'h4134f38d, 32'hc23d853b, 32'h42701b48, 32'hc1042e3a};
test_bias[2830:2830] = '{32'h40d04fb9};
test_output[2830:2830] = '{32'h45ba93af};
test_input[22648:22655] = '{32'hc294bd9e, 32'hc15eec88, 32'hbf8252f3, 32'h422d1f52, 32'h420b6d2b, 32'hc22db1ad, 32'h42932ecd, 32'h41160c60};
test_weights[22648:22655] = '{32'h415442c3, 32'h4187b3f8, 32'hc2c0dca9, 32'h4247b82b, 32'hc1be6aa9, 32'h4285d479, 32'h4219b7ea, 32'h4217e728};
test_bias[2831:2831] = '{32'h41f6b7a7};
test_output[2831:2831] = '{32'h4400fc14};
test_input[22656:22663] = '{32'hc21414c3, 32'hc288af1d, 32'hc1bc12c2, 32'hc250269b, 32'h421f3728, 32'h423e8d75, 32'hc1a51f07, 32'h41940016};
test_weights[22656:22663] = '{32'hc2b06d0e, 32'hc21de02f, 32'hc1ee383d, 32'hc1f2a129, 32'h4189bbcf, 32'h4215b68d, 32'h424ecc00, 32'h42a120f2};
test_bias[2832:2832] = '{32'h41f96536};
test_output[2832:2832] = '{32'h462e70b5};
test_input[22664:22671] = '{32'h42c1b78e, 32'h41b052c2, 32'h4273db3a, 32'hc21287e2, 32'h4223c24b, 32'hc2a3c837, 32'h422d7e9e, 32'hc2334f76};
test_weights[22664:22671] = '{32'h41c1810f, 32'hc27815e5, 32'h4283f102, 32'h3f99dac9, 32'hc2c0b9d4, 32'h42b8a352, 32'h42a3c38f, 32'h422f8f06};
test_bias[2833:2833] = '{32'h4193bd3d};
test_output[2833:2833] = '{32'hc59aa807};
test_input[22672:22679] = '{32'h41874c61, 32'hc1137849, 32'h427c09e5, 32'hc00b67be, 32'h429d348d, 32'h4157e885, 32'hc2126469, 32'hc023d0b1};
test_weights[22672:22679] = '{32'hc2c2a1a4, 32'h40c63b7e, 32'h41825e7d, 32'h428fa2fe, 32'h41f6830e, 32'hc24fd98c, 32'hc277b451, 32'h425975bd};
test_bias[2834:2834] = '{32'h41e2553c};
test_output[2834:2834] = '{32'h453e3d46};
test_input[22680:22687] = '{32'h42b1b2bb, 32'hc199b27b, 32'hc0af7271, 32'hc1786473, 32'hc2ace0bf, 32'h42ac6902, 32'h4101b4ac, 32'h4268ab50};
test_weights[22680:22687] = '{32'hbdc4b4cd, 32'h428d3b6d, 32'hc0a3eab6, 32'hc2c63780, 32'hc285e26c, 32'hc0b3a4d6, 32'h4088551b, 32'h4252399c};
test_bias[2835:2835] = '{32'h42875724};
test_output[2835:2835] = '{32'h46075cd7};
test_input[22688:22695] = '{32'hc2615773, 32'h3e999aa4, 32'h42ac25fb, 32'h414a00af, 32'h42b254ef, 32'h42b76d97, 32'h40823799, 32'hc25fcd7f};
test_weights[22688:22695] = '{32'hc2c0c2c3, 32'hc21c7c75, 32'h42b98d20, 32'h4246c7bc, 32'hc220e972, 32'h428cb685, 32'h41eb1a53, 32'hc143a19e};
test_bias[2836:2836] = '{32'h42adf2a4};
test_output[2836:2836] = '{32'h468af68a};
test_input[22696:22703] = '{32'hc25308c6, 32'hc24ebdf2, 32'hc24f4638, 32'hbfa0949a, 32'hc234be76, 32'hc2343d50, 32'h429517c2, 32'h41566e9b};
test_weights[22696:22703] = '{32'h41d90c23, 32'h42acb21f, 32'h4207cac7, 32'hc2a0874a, 32'h42685fac, 32'hc21b80ca, 32'hc2bba87a, 32'hc25c45a0};
test_bias[2837:2837] = '{32'h415902ae};
test_output[2837:2837] = '{32'hc67c4476};
test_input[22704:22711] = '{32'hc29d2854, 32'hc2943cdd, 32'h4295259c, 32'h4297af54, 32'h421ad0df, 32'h42c63d3e, 32'h41b26baf, 32'h3f4a9aec};
test_weights[22704:22711] = '{32'hc2a98e92, 32'h410d1b26, 32'hc24d277f, 32'hc207f60d, 32'hc09c901d, 32'h4128cf82, 32'h42377f1a, 32'h4290a1dd};
test_bias[2838:2838] = '{32'hc2238bf9};
test_output[2838:2838] = '{32'h44bbaa57};
test_input[22712:22719] = '{32'hc13d336b, 32'h417501a5, 32'hc252f586, 32'h427ee010, 32'h42c03ce0, 32'h413ed0e1, 32'h428f6f29, 32'h422d40c3};
test_weights[22712:22719] = '{32'hc0c43abe, 32'h42161065, 32'h426e1e02, 32'hc150bd73, 32'hc1d5fc56, 32'hc2ab29b7, 32'hbf55c17f, 32'h40064c45};
test_bias[2839:2839] = '{32'h4242fe6b};
test_output[2839:2839] = '{32'hc5d59e13};
test_input[22720:22727] = '{32'h41872135, 32'hc26f7e50, 32'hc165c174, 32'h427f31c0, 32'hc2205356, 32'hc297a5a6, 32'hc217aa0d, 32'hc217f206};
test_weights[22720:22727] = '{32'hc08a972f, 32'hc2061396, 32'hc2bfe90b, 32'hc2bc908a, 32'h42b49a9f, 32'h42bad822, 32'hc105b9bd, 32'hc20e2739};
test_bias[2840:2840] = '{32'h40ea8c41};
test_output[2840:2840] = '{32'hc6375112};
test_input[22728:22735] = '{32'hc2c1bb7e, 32'h428655a0, 32'hc2c54873, 32'hc28011a4, 32'hc2970007, 32'h41c22b20, 32'hc208b778, 32'hc0ecf550};
test_weights[22728:22735] = '{32'hc28b8559, 32'h4270921a, 32'hc12961ea, 32'hc2a38bf7, 32'hc110a80e, 32'hc287a873, 32'hc1acfce1, 32'hc228ccf4};
test_bias[2841:2841] = '{32'h42c6d029};
test_output[2841:2841] = '{32'h4686e1cf};
test_input[22736:22743] = '{32'h421a6e7c, 32'hc286f17b, 32'h4286543e, 32'hc2c7b38e, 32'hc2b9698c, 32'h42b36aba, 32'hc2a33678, 32'hc038a67a};
test_weights[22736:22743] = '{32'hc2130ea2, 32'h426f69a2, 32'hc25cf96d, 32'h415fcc5f, 32'hc167ff2d, 32'hc25fc3f6, 32'h425293fb, 32'hc2576c2a};
test_bias[2842:2842] = '{32'hc201a070};
test_output[2842:2842] = '{32'hc68fd861};
test_input[22744:22751] = '{32'hc226dd93, 32'h423ce8b8, 32'hc1b5df02, 32'h429a7e7a, 32'h407f3271, 32'h428ee22f, 32'h42c180a7, 32'hc2a377c9};
test_weights[22744:22751] = '{32'hc0bc6e28, 32'hc0a7c6ea, 32'h421c5d64, 32'hbff867dd, 32'h41d2103d, 32'hc299531d, 32'h429a4a35, 32'hc2753ba8};
test_bias[2843:2843] = '{32'hc20c3744};
test_output[2843:2843] = '{32'h45bc5824};
test_input[22752:22759] = '{32'h42447335, 32'h42c290f1, 32'h41f701b1, 32'hc1610198, 32'hc1d141af, 32'h42b6ad34, 32'hc231ca02, 32'h420ba507};
test_weights[22752:22759] = '{32'h4195edf5, 32'h42bc4f57, 32'hc003b37e, 32'hc0a6877c, 32'h42739ad6, 32'hc0829547, 32'hc0c3f0c5, 32'hc2ad8404};
test_bias[2844:2844] = '{32'h4229796f};
test_output[2844:2844] = '{32'h45a90df3};
test_input[22760:22767] = '{32'h41912ddd, 32'hc1d9dcf6, 32'h4154471d, 32'h42709fe5, 32'hc2979b28, 32'hc2b7bdf9, 32'h42c21809, 32'hc1467d74};
test_weights[22760:22767] = '{32'hc2344d08, 32'hc245c31c, 32'h422fbd35, 32'h3bf47bb3, 32'hc273d36d, 32'hc0873cbc, 32'hc22fb6a6, 32'h4227233b};
test_bias[2845:2845] = '{32'h41a81533};
test_output[2845:2845] = '{32'h44aa07b3};
test_input[22768:22775] = '{32'h42a47c4b, 32'hc27526f6, 32'h425d1a0d, 32'hc2b99a65, 32'h41ca8ee0, 32'hc296a164, 32'h42134b01, 32'hc212a241};
test_weights[22768:22775] = '{32'h42aa1733, 32'hc299c83e, 32'h42143606, 32'h423039b8, 32'hc1d89e45, 32'h41eaa466, 32'hbdd0973c, 32'h41de895a};
test_bias[2846:2846] = '{32'h425b55f2};
test_output[2846:2846] = '{32'h45b559c5};
test_input[22776:22783] = '{32'hc2bf20a2, 32'h426a3dbc, 32'hc2adfb61, 32'hc169b4d7, 32'h425e2d3a, 32'h417cbd56, 32'hc29dbedf, 32'h4244eaa8};
test_weights[22776:22783] = '{32'hc2a91b97, 32'h41073ff5, 32'hc2b4f4d6, 32'hc2349a0c, 32'hc1277807, 32'h41c7b3da, 32'hc1b669ca, 32'h42190d4f};
test_bias[2847:2847] = '{32'h4296feaa};
test_output[2847:2847] = '{32'h46a1883b};
test_input[22784:22791] = '{32'hc2ba4534, 32'hc2249f1a, 32'h4126c9d8, 32'hc1eaa97a, 32'h429587d1, 32'h42341a1d, 32'h4121a009, 32'hc278a7ee};
test_weights[22784:22791] = '{32'hc16915a5, 32'hc1d03b63, 32'h41ce0402, 32'h42675cae, 32'h4224cee6, 32'hc12e6d33, 32'h42364178, 32'hc256c4a2};
test_bias[2848:2848] = '{32'hc204de94};
test_output[2848:2848] = '{32'h45e5d1c4};
test_input[22792:22799] = '{32'hc19a9fdf, 32'hc2a552bc, 32'hc285b1ae, 32'h421812ba, 32'h4207de71, 32'h41b3b1a5, 32'hc25660d8, 32'hc08875d8};
test_weights[22792:22799] = '{32'hc1318a78, 32'h4043872e, 32'h4234f89c, 32'hc2b648c3, 32'hc243eaeb, 32'hc2bde929, 32'h421c9e77, 32'hc13fe308};
test_bias[2849:2849] = '{32'h42b78467};
test_output[2849:2849] = '{32'hc63fde7e};
test_input[22800:22807] = '{32'hc2c2279f, 32'hc2939822, 32'h41cff44f, 32'hc29a9d28, 32'hc2a10aa4, 32'h42215459, 32'h425be0ba, 32'h428ea5dd};
test_weights[22800:22807] = '{32'hc238d09f, 32'h4092b8e5, 32'hc1f69641, 32'hc2606436, 32'h420082bc, 32'h42bc9f64, 32'h42a12535, 32'hc284bd9e};
test_bias[2850:2850] = '{32'h414eed63};
test_output[2850:2850] = '{32'h46067e17};
test_input[22808:22815] = '{32'h42bf2fb4, 32'h42694e15, 32'hc2741d64, 32'h41b83e28, 32'hc282ba20, 32'h42557652, 32'h42a0b3e7, 32'hc022aafc};
test_weights[22808:22815] = '{32'h42be9d97, 32'hc2009ec7, 32'h423aa71d, 32'hc211b746, 32'h42ba4421, 32'h423e1723, 32'hc2927e14, 32'hc25384e3};
test_bias[2851:2851] = '{32'h4295b9ea};
test_output[2851:2851] = '{32'hc5b178a7};
test_input[22816:22823] = '{32'h42c2cdd1, 32'h41ea159d, 32'hc28a7062, 32'hc23a717b, 32'hc2a8eda8, 32'hc1e4343d, 32'hc2c3cd1c, 32'h42a1a6b9};
test_weights[22816:22823] = '{32'h412200fc, 32'h41682f6b, 32'hc2384216, 32'h4286630e, 32'h4295eee3, 32'h42c1579d, 32'h40f585bf, 32'h420bdb7d};
test_bias[2852:2852] = '{32'hc281db3d};
test_output[2852:2852] = '{32'hc5af6182};
test_input[22824:22831] = '{32'hc2804893, 32'h42444f52, 32'h41c798b5, 32'hc2360913, 32'hc2af2686, 32'hc25bff9d, 32'hc2c471bb, 32'h428a9985};
test_weights[22824:22831] = '{32'hc24b471f, 32'h42943d90, 32'h42950ce8, 32'h423dee2d, 32'h42045eaa, 32'hc28785ff, 32'h41f62ffd, 32'hc1cb5c31};
test_bias[2853:2853] = '{32'hc2bbf36e};
test_output[2853:2853] = '{32'h451f25a7};
test_input[22832:22839] = '{32'h42bab402, 32'hc1688175, 32'h3f4133a6, 32'hc2a36a4c, 32'h4140a347, 32'h4298f9fd, 32'h42a684ab, 32'hbf13a4cd};
test_weights[22832:22839] = '{32'hc211b33e, 32'h4211ff59, 32'hc2915243, 32'h426a3a01, 32'hc23df2a8, 32'h42625a17, 32'h410fc086, 32'hc2c284b3};
test_bias[2854:2854] = '{32'h42682eb5};
test_output[2854:2854] = '{32'hc581baa4};
test_input[22840:22847] = '{32'hc255b582, 32'hc1d3b03a, 32'hc2360fe8, 32'hc22b81c3, 32'hc2af6f86, 32'h4250bd8f, 32'h425a4c50, 32'hc26744aa};
test_weights[22840:22847] = '{32'h4274bee9, 32'hc294e58d, 32'hc2a96ff6, 32'h42b75beb, 32'hc228d8d1, 32'h41890b14, 32'h419d9664, 32'h4243146e};
test_bias[2855:2855] = '{32'hc258b0e9};
test_output[2855:2855] = '{32'h44b1fb58};
test_input[22848:22855] = '{32'h42c56af2, 32'hc2b5a2f4, 32'h4280ed39, 32'hc1ce8f2f, 32'hc203fdde, 32'h42340920, 32'hc264da5f, 32'h428f0339};
test_weights[22848:22855] = '{32'h42a92961, 32'hc2bb0bb6, 32'hc213e13f, 32'h42027a7f, 32'h42092dfb, 32'hc2344ee0, 32'h40357ca8, 32'h427f8599};
test_bias[2856:2856] = '{32'h42c44316};
test_output[2856:2856] = '{32'h4669c0f2};
test_input[22856:22863] = '{32'h42605c92, 32'hc1cb2388, 32'hc184130b, 32'hc1f640b9, 32'h40d1525f, 32'hc1bec224, 32'h41d42f00, 32'hc287fc10};
test_weights[22856:22863] = '{32'hc1e8fd28, 32'h4285c82c, 32'hc238a560, 32'hc2aa3476, 32'hc2b45b09, 32'hc21df485, 32'h41fca9cb, 32'hc2aee023};
test_bias[2857:2857] = '{32'hc24bc829};
test_output[2857:2857] = '{32'h45dee93b};
test_input[22864:22871] = '{32'h415a8d59, 32'h42874f23, 32'hc2c4eeaf, 32'hc187ea23, 32'hc2117dde, 32'hc2024552, 32'h4287500f, 32'hc1e8f44f};
test_weights[22864:22871] = '{32'hc2629e5e, 32'hc2895554, 32'h42757c0a, 32'hc0439416, 32'hc1b67cab, 32'hc2392fc6, 32'h4192a09d, 32'hc2ac5c15};
test_bias[2858:2858] = '{32'h41bcfd98};
test_output[2858:2858] = '{32'hc5a59f62};
test_input[22872:22879] = '{32'hc2863ada, 32'hc2b90dc8, 32'hc2979ed6, 32'hc2057cfa, 32'h42a50b49, 32'hc1d09c1a, 32'h42718d9f, 32'hc1c85dee};
test_weights[22872:22879] = '{32'h42701d4e, 32'h404c3b1f, 32'h42994d1d, 32'h418afb61, 32'hc23e33dd, 32'hc265229a, 32'hc24f043e, 32'hc266a682};
test_bias[2859:2859] = '{32'hbfc8ee12};
test_output[2859:2859] = '{32'hc667aeb9};
test_input[22880:22887] = '{32'hc2a6e0f1, 32'h41d0b7e2, 32'hc17898ec, 32'h42afae2e, 32'hc2402907, 32'hc232a877, 32'hc013b58f, 32'hc1d4ce76};
test_weights[22880:22887] = '{32'h402bd30c, 32'h41d8b329, 32'h429962c9, 32'h41d20ba7, 32'h425ab003, 32'hc284e4a7, 32'h42bc9d96, 32'h42c194d8};
test_bias[2860:2860] = '{32'hc10f9a1e};
test_output[2860:2860] = '{32'hc457a5a2};
test_input[22888:22895] = '{32'hc24a55d2, 32'hc0ac1027, 32'h41ca0012, 32'h4146a394, 32'h41228a7c, 32'hc2ac812c, 32'h416369b1, 32'h4221cf22};
test_weights[22888:22895] = '{32'h425e341f, 32'hc2b627e5, 32'h428e621f, 32'hc278c114, 32'hc2458161, 32'h4285e9ce, 32'h42bb530d, 32'hc2a5e1b4};
test_bias[2861:2861] = '{32'h41e6dbd0};
test_output[2861:2861] = '{32'hc6157a25};
test_input[22896:22903] = '{32'hc28209f1, 32'hc299c764, 32'hc27887aa, 32'hc27a74cb, 32'h42c21d20, 32'h41841943, 32'hc2878870, 32'h4138b075};
test_weights[22896:22903] = '{32'hc286426e, 32'hc1e3ece3, 32'hc25be75f, 32'h42ab166e, 32'h426137b1, 32'hc2c502f7, 32'hc1e95ee5, 32'hc295ee63};
test_bias[2862:2862] = '{32'h40f27584};
test_output[2862:2862] = '{32'h461590a9};
test_input[22904:22911] = '{32'hc291781f, 32'h40bef8d7, 32'h41c67201, 32'h42730960, 32'hc2a9accf, 32'h42a3d258, 32'h428b8721, 32'hc1ebae5e};
test_weights[22904:22911] = '{32'hc2532f09, 32'h428a71c7, 32'h423746c9, 32'h424aafcf, 32'h41b36685, 32'hc2a7a011, 32'hc2bd4b8d, 32'h41cd9277};
test_bias[2863:2863] = '{32'hc24a6e06};
test_output[2863:2863] = '{32'hc5f0edc2};
test_input[22912:22919] = '{32'hc28cc1d9, 32'hc299284e, 32'hc2960a49, 32'hc0bce7f6, 32'h424a70e6, 32'h4289d9a5, 32'h429e3b35, 32'h426092ab};
test_weights[22912:22919] = '{32'hc29c6080, 32'h420892d0, 32'h427cdcd9, 32'hc1c0cde7, 32'h40bc6fc3, 32'h4261caff, 32'h428e5b74, 32'hc22d7cde};
test_bias[2864:2864] = '{32'hc2bae09e};
test_output[2864:2864] = '{32'h45ae5c72};
test_input[22920:22927] = '{32'h42445b19, 32'hc2a6df1b, 32'hc29721ac, 32'hc294d42e, 32'h42b23746, 32'h42bc10a2, 32'h4284bd28, 32'hc27ca63a};
test_weights[22920:22927] = '{32'h42a55457, 32'h41f4fc51, 32'h42184afd, 32'hc1320ff1, 32'hc1eeb21e, 32'h40d56b20, 32'h427ab56c, 32'h426ab2b7};
test_bias[2865:2865] = '{32'h42bf492a};
test_output[2865:2865] = '{32'hc4fd8440};
test_input[22928:22935] = '{32'hc2ae1ec6, 32'h40536c27, 32'hc2b95050, 32'h4190fb51, 32'hc2229400, 32'hc2147008, 32'hc281ac35, 32'h4210ed77};
test_weights[22928:22935] = '{32'hc29ecc3d, 32'hc29234d3, 32'hc2a38edb, 32'hc29b0da0, 32'hc2b327a7, 32'hc267f490, 32'hc2688c59, 32'h4161041f};
test_bias[2866:2866] = '{32'hc2bf2a68};
test_output[2866:2866] = '{32'h46b24700};
test_input[22936:22943] = '{32'hc239eb03, 32'h42bc4bca, 32'h4268aa25, 32'hc2a6b637, 32'h42c7bb31, 32'hc0ff6052, 32'hc2819962, 32'hc29477ad};
test_weights[22936:22943] = '{32'hc11524ed, 32'hc220044d, 32'hc29eb850, 32'hc2366ef5, 32'h42244f21, 32'hc23ee7d7, 32'h42553c53, 32'h42a9cde8};
test_bias[2867:2867] = '{32'h427b283a};
test_output[2867:2867] = '{32'hc6123a14};
test_input[22944:22951] = '{32'h42b5a48b, 32'h417d09d9, 32'hc2695548, 32'h423285d2, 32'h4208f426, 32'hc29fa1d7, 32'h42a8401a, 32'h419940a5};
test_weights[22944:22951] = '{32'hc1958f13, 32'h41a8c796, 32'h4279425a, 32'hc258e7a5, 32'hc277f737, 32'hc27284a6, 32'hc272b062, 32'h42a5318f};
test_bias[2868:2868] = '{32'hc291f868};
test_output[2868:2868] = '{32'hc601a5e5};
test_input[22952:22959] = '{32'hc22b3fd1, 32'h4297904d, 32'h41580140, 32'hbed149ee, 32'hc0451ef2, 32'h414c0a30, 32'hc278a3e4, 32'h42aa7330};
test_weights[22952:22959] = '{32'hc1240570, 32'hc0d8b16d, 32'hc1eaf4b5, 32'hc2c6b4fe, 32'hc20a8dff, 32'h406d20f8, 32'hc28f3650, 32'hc25d7f7c};
test_bias[2869:2869] = '{32'hc20e6d60};
test_output[2869:2869] = '{32'hc41105ef};
test_input[22960:22967] = '{32'h424a1644, 32'h42023e2a, 32'hc214b2fc, 32'hc2a1092b, 32'h42acccd2, 32'hc23dd3d2, 32'hc263bb3e, 32'hc2c529d8};
test_weights[22960:22967] = '{32'h41354364, 32'h42609bef, 32'h428b6ae0, 32'hc2b08452, 32'h4147ba23, 32'hc15cf80c, 32'h429321f4, 32'h42a78d4d};
test_bias[2870:2870] = '{32'hc1fc42cf};
test_output[2870:2870] = '{32'hc56f506e};
test_input[22968:22975] = '{32'hc2b8df16, 32'hc14220b3, 32'h42299b99, 32'hc2928616, 32'hc28c4d0a, 32'hc1ff0fd8, 32'hc28a9484, 32'h4207ea63};
test_weights[22968:22975] = '{32'h4105d956, 32'hc2ac45ac, 32'hc0fc5b0a, 32'hc264e69c, 32'hc2b61363, 32'hc1a5e1e6, 32'hc29d43b8, 32'h42c27f97};
test_bias[2871:2871] = '{32'h428a46a4};
test_output[2871:2871] = '{32'h469c3e95};
test_input[22976:22983] = '{32'hc29b1800, 32'h42ab1326, 32'h41de0bdb, 32'hc194f226, 32'hc1dafa9d, 32'h42a2add4, 32'h427b1609, 32'h4175305a};
test_weights[22976:22983] = '{32'hc222a309, 32'hc1edcfa3, 32'hc2059cd2, 32'hc22c80d5, 32'h4293b163, 32'h42b62795, 32'hc26b7165, 32'h4286a041};
test_bias[2872:2872] = '{32'hc227c121};
test_output[2872:2872] = '{32'h4545fb65};
test_input[22984:22991] = '{32'hc20ccecc, 32'hc20b8745, 32'h4265ed0c, 32'hc26089e6, 32'hc29f1189, 32'hc2b270c5, 32'hc15da013, 32'hc1a279d4};
test_weights[22984:22991] = '{32'h42159ed6, 32'h42acafa9, 32'h42502672, 32'h41a3fb17, 32'h42471aed, 32'h429bda70, 32'h424677d2, 32'h42aad9a8};
test_bias[2873:2873] = '{32'h422a6935};
test_output[2873:2873] = '{32'hc6768ca1};
test_input[22992:22999] = '{32'h41bfb249, 32'h41fe4afa, 32'h42215008, 32'h4268e519, 32'hc1bf273b, 32'hc29396a2, 32'h4275174f, 32'h422eb677};
test_weights[22992:22999] = '{32'hc24d50a2, 32'hc190e252, 32'hc1a7fe40, 32'h428c45a5, 32'h420376e5, 32'h423f423b, 32'h42850451, 32'hc1302ffc};
test_bias[2874:2874] = '{32'h426b065c};
test_output[2874:2874] = '{32'h444092fa};
test_input[23000:23007] = '{32'hc2b64fc7, 32'h42bdcb6a, 32'hc2098c66, 32'hc1e9b2bb, 32'hc184ea16, 32'h418420d9, 32'h426f4ce7, 32'hc29a266a};
test_weights[23000:23007] = '{32'hc25496ee, 32'hc25a239e, 32'h42747282, 32'hc29e1d65, 32'h40f79805, 32'h42a12f7a, 32'hc080404f, 32'h424e5f4f};
test_bias[2875:2875] = '{32'hc27afb4a};
test_output[2875:2875] = '{32'hc547f0d3};
test_input[23008:23015] = '{32'h41be8881, 32'hc23cd12d, 32'hc2a5abd3, 32'h424a7781, 32'hc2166fc9, 32'h42297651, 32'h411c3f8a, 32'h42702475};
test_weights[23008:23015] = '{32'hc294fca7, 32'h42a3f4f7, 32'h41885565, 32'h4290d336, 32'h4289269f, 32'hc2973f48, 32'h42336e69, 32'hc115d11a};
test_bias[2876:2876] = '{32'hc1360244};
test_output[2876:2876] = '{32'hc61172a0};
test_input[23016:23023] = '{32'hc2795004, 32'hc2714b70, 32'h418f0067, 32'hc28aecfe, 32'hc1958746, 32'h42b89499, 32'h422f18a2, 32'hc2c013cb};
test_weights[23016:23023] = '{32'h42b729e9, 32'h42678a67, 32'h42069ae2, 32'h41b149ab, 32'hc2960c23, 32'h3fec5902, 32'h4298f8f0, 32'hc2b51e86};
test_bias[2877:2877] = '{32'h42b6174c};
test_output[2877:2877] = '{32'h455f3400};
test_input[23024:23031] = '{32'hc13b5219, 32'hc1f22019, 32'h42979ef3, 32'hc102cafc, 32'hc210a1e2, 32'h41ede438, 32'hc2928f88, 32'hc1d2f9ff};
test_weights[23024:23031] = '{32'h4272266d, 32'hc14943f6, 32'hc220dd8a, 32'h4100d8c8, 32'h4236c781, 32'hc20dfb15, 32'hc2a9c0e4, 32'h40c6c9be};
test_bias[2878:2878] = '{32'hc2abfb40};
test_output[2878:2878] = '{32'hc334707f};
test_input[23032:23039] = '{32'hc2a1383c, 32'hc2982673, 32'hbda50024, 32'h429bc928, 32'hc2a60abc, 32'hc1c5f874, 32'h42b459bf, 32'hc2376c0f};
test_weights[23032:23039] = '{32'h410e965b, 32'hc24f8783, 32'h42acc182, 32'h42a015a6, 32'h42990070, 32'h425e7173, 32'hc2716e2b, 32'hc1b75d4d};
test_bias[2879:2879] = '{32'hc256d748};
test_output[2879:2879] = '{32'hc529c6dc};
test_input[23040:23047] = '{32'hc0a398c4, 32'h420e7b88, 32'h42ae3a1e, 32'h3decdc46, 32'h42afecc8, 32'h4287eb7e, 32'hc28686f2, 32'h41797239};
test_weights[23040:23047] = '{32'h4246e247, 32'hc2a7712f, 32'hc27c780e, 32'h41abe3df, 32'h4275f9f1, 32'h41f337be, 32'h429ce9f9, 32'hc2965d3d};
test_bias[2880:2880] = '{32'h40efac69};
test_output[2880:2880] = '{32'hc5f0971e};
test_input[23048:23055] = '{32'h4281fd7c, 32'hc2052928, 32'hc2b356e6, 32'hc1c4d5f0, 32'h42aebe8b, 32'hc22e38bb, 32'hc299948b, 32'h4133179f};
test_weights[23048:23055] = '{32'hc1f26d67, 32'hc2092e34, 32'hc2ae6ca4, 32'h418837f6, 32'hc204f533, 32'h4114a164, 32'hc27acbef, 32'h4143b57e};
test_bias[2881:2881] = '{32'h42acebcb};
test_output[2881:2881] = '{32'h4601bad3};
test_input[23056:23063] = '{32'hc2ac527d, 32'h42878bd3, 32'hc2364af6, 32'h41c53078, 32'hc11960ae, 32'h4235a80d, 32'h42bc89ad, 32'hc0005943};
test_weights[23056:23063] = '{32'hc2b9cfef, 32'hc1998147, 32'hc28c74f9, 32'hc2bd0d77, 32'h421cdb02, 32'h427279f1, 32'h41ccda71, 32'h424d905a};
test_bias[2882:2882] = '{32'h42559da7};
test_output[2882:2882] = '{32'h46407169};
test_input[23064:23071] = '{32'h4149bb45, 32'h42ae28dd, 32'h4063f9bf, 32'hc153bd3b, 32'h41f7847d, 32'h427308f1, 32'h425bec82, 32'h421f0a1a};
test_weights[23064:23071] = '{32'hc0ae07c6, 32'h424075ba, 32'h42287182, 32'h4054bec5, 32'h400609bf, 32'h42461c47, 32'h4281f0bc, 32'h40aac77f};
test_bias[2883:2883] = '{32'hc1a71d0f};
test_output[2883:2883] = '{32'h462ce2fc};
test_input[23072:23079] = '{32'h41830ab3, 32'hc202e5d5, 32'h3fa549f0, 32'hc2227d13, 32'h422c0dc4, 32'h42a7f3e5, 32'h4199b02b, 32'h42820a01};
test_weights[23072:23079] = '{32'hc14da4b1, 32'h41f8954d, 32'hc29ee06c, 32'hc0cc3485, 32'hc2c7c6e9, 32'h4295fdc0, 32'hc29cb05c, 32'h41f74f14};
test_bias[2884:2884] = '{32'hc2a9c468};
test_output[2884:2884] = '{32'h44a8d38c};
test_input[23080:23087] = '{32'h42b22646, 32'h426bb63b, 32'h428a9ccf, 32'hc2b3c783, 32'hc0c465d8, 32'hc22e0124, 32'hc20c40ee, 32'hc2b36969};
test_weights[23080:23087] = '{32'h412ae03b, 32'hc1a1a794, 32'hc217abe4, 32'hc253b3cb, 32'hc1aaae92, 32'hc259fe7a, 32'hc20b1fe3, 32'h411c8384};
test_bias[2885:2885] = '{32'h4210a90b};
test_output[2885:2885] = '{32'h45950fa0};
test_input[23088:23095] = '{32'h420d43d3, 32'h423ce981, 32'h42c72fcd, 32'h42b22f89, 32'hc2bbc207, 32'h428c37e5, 32'hc2c64fce, 32'h42c74269};
test_weights[23088:23095] = '{32'h423e611a, 32'hc2adf063, 32'h4286b03d, 32'hc288a88e, 32'hc145b958, 32'hc2534fba, 32'hc194681b, 32'hc2a7fabf};
test_bias[2886:2886] = '{32'hc265f603};
test_output[2886:2886] = '{32'hc62ae2a3};
test_input[23096:23103] = '{32'h422355ff, 32'h423b7a42, 32'h42711d7f, 32'hc2b9af2c, 32'hc2b2eb5b, 32'hc2103687, 32'hc2bdcdfd, 32'hc26f6e67};
test_weights[23096:23103] = '{32'h41f641a2, 32'h42bcf829, 32'hc1715395, 32'h420b2943, 32'h422edab4, 32'hc1a762d7, 32'hc2a60542, 32'h42612f0c};
test_bias[2887:2887] = '{32'h41592847};
test_output[2887:2887] = '{32'h4535fa52};
test_input[23104:23111] = '{32'h4153075f, 32'h417e5f23, 32'hc288d458, 32'h41f967ba, 32'hc252db72, 32'hc2929a91, 32'h42a3b968, 32'hc2c3622b};
test_weights[23104:23111] = '{32'hc2926fa2, 32'h429d5e03, 32'h4207d5ec, 32'h42787bd2, 32'h4216a606, 32'hc285558f, 32'hc18b2d86, 32'hc2a5f976};
test_bias[2888:2888] = '{32'hbf7ca30a};
test_output[2888:2888] = '{32'h46142869};
test_input[23112:23119] = '{32'hc2694a8d, 32'h42917baf, 32'hc201f058, 32'h426aacd5, 32'h42391100, 32'h42c517f9, 32'hc2b8a496, 32'h42b9d2a6};
test_weights[23112:23119] = '{32'h40ce9ee1, 32'h42380fe0, 32'h40e85c47, 32'hc2b0c39e, 32'hc2a9c7b4, 32'hc2c5ff74, 32'hc0961158, 32'h427a5e7e};
test_bias[2889:2889] = '{32'h422c6f14};
test_output[2889:2889] = '{32'hc619c9fe};
test_input[23120:23127] = '{32'h424c7703, 32'hc2a3a2c9, 32'hc28b7dca, 32'hc23bf831, 32'h4285b0e0, 32'h3f50a6b3, 32'hc21328e4, 32'hc232f923};
test_weights[23120:23127] = '{32'hc209f1e3, 32'hc2034323, 32'h429553f3, 32'h4293ef7b, 32'h42812b7a, 32'h4247a115, 32'h4138967a, 32'hc2a6976b};
test_bias[2890:2890] = '{32'h41f1050d};
test_output[2890:2890] = '{32'hc28d9e77};
test_input[23128:23135] = '{32'h42806c7c, 32'hc1134b77, 32'h42498a15, 32'h41c28fe9, 32'hc1709fe8, 32'h4219f2de, 32'h42af458a, 32'h4183148c};
test_weights[23128:23135] = '{32'h42a3a6a0, 32'hbd31838b, 32'h4201740a, 32'hc2b47b68, 32'hc2227b2e, 32'h42651a4f, 32'h419c3b1a, 32'h4210b93e};
test_bias[2891:2891] = '{32'hc23542af};
test_output[2891:2891] = '{32'h461892d4};
test_input[23136:23143] = '{32'h4120f4c9, 32'hc2154078, 32'h41d922ba, 32'h4240ec76, 32'hc283297a, 32'hc2c2ef4b, 32'h428f7fc6, 32'hc295c6a4};
test_weights[23136:23143] = '{32'h428428dc, 32'h422d2495, 32'hc2c36b8b, 32'h415e9def, 32'h42aa79ef, 32'hc185a409, 32'hc1905d49, 32'hc2438a26};
test_bias[2892:2892] = '{32'h42a9f9f3};
test_output[2892:2892] = '{32'hc58ad041};
test_input[23144:23151] = '{32'hc216d54b, 32'h41ef6f57, 32'hc20fea7f, 32'hc2a550f1, 32'hc2a9b5f6, 32'h425ece1c, 32'h429eb4a5, 32'hbff0ff7b};
test_weights[23144:23151] = '{32'hc254d6e1, 32'h42ac5f33, 32'hc0d0e7fb, 32'hc2a74552, 32'hc28c0e86, 32'hc1f4175d, 32'hc299151a, 32'hc2c266a7};
test_bias[2893:2893] = '{32'h42127d6c};
test_output[2893:2893] = '{32'h461e2a64};
test_input[23152:23159] = '{32'h42a3060b, 32'hc1b97ac9, 32'h41d0f2d7, 32'h42c21367, 32'h428e947c, 32'h41348780, 32'h41907315, 32'h4197469d};
test_weights[23152:23159] = '{32'hc214d63d, 32'h41d704d5, 32'h4298850c, 32'h41a4af80, 32'hc2900b20, 32'h41eaaf8a, 32'hc18d5991, 32'hc22fc811};
test_bias[2894:2894] = '{32'h42a6a77e};
test_output[2894:2894] = '{32'hc5ad06f5};
test_input[23160:23167] = '{32'h4283edce, 32'hc15608f4, 32'h424c6ba6, 32'hc2c77382, 32'hc2718445, 32'h3ffc11fc, 32'hc264cf19, 32'h3dc516c5};
test_weights[23160:23167] = '{32'hc1d26253, 32'hc2b08a05, 32'hc27afb67, 32'hc1079b5a, 32'hc2962430, 32'hc160db87, 32'hc2876bc0, 32'hc2bdc12e};
test_bias[2895:2895] = '{32'h41c88c5f};
test_output[2895:2895] = '{32'h45ab3693};
test_input[23168:23175] = '{32'hc27ce85c, 32'h424677c1, 32'h42a408d2, 32'h42c11a9d, 32'hc2884c24, 32'hc2382a30, 32'h4180317e, 32'h418ae1cf};
test_weights[23168:23175] = '{32'h4077d95c, 32'h4099b9cd, 32'h41536bdc, 32'hc2908b32, 32'hc1e6faa1, 32'h42ab5c9b, 32'hc291dd93, 32'h42595699};
test_bias[2896:2896] = '{32'h41001699};
test_output[2896:2896] = '{32'hc5fcfb10};
test_input[23176:23183] = '{32'hc2b4612a, 32'h428e8738, 32'h422dd1c7, 32'hc2b5c13d, 32'h425c7f8d, 32'h42bb07f5, 32'h42381382, 32'h40d930f5};
test_weights[23176:23183] = '{32'h423e47d4, 32'hc11ecdac, 32'hc2a51e3e, 32'h42951aa0, 32'h420a4f66, 32'hc1a71b8a, 32'hc26da988, 32'hc21d7987};
test_bias[2897:2897] = '{32'h42739823};
test_output[2897:2897] = '{32'hc68f586e};
test_input[23184:23191] = '{32'h423439b6, 32'hc20949d3, 32'h42237156, 32'h4190a344, 32'h425b5bcb, 32'hc2b22037, 32'h425f2770, 32'h428082f3};
test_weights[23184:23191] = '{32'h42189a7c, 32'h41b9dec5, 32'h420cde28, 32'hc2acb5ff, 32'h415f3ac5, 32'h3fbc6b5a, 32'hc210c890, 32'h42be802e};
test_bias[2898:2898] = '{32'hc28e61c6};
test_output[2898:2898] = '{32'h45aab8d5};
test_input[23192:23199] = '{32'h429bbb92, 32'hc1d45754, 32'hc23c61ad, 32'hc1e71974, 32'hc1dfc6da, 32'h4284b1d9, 32'h42b2c2f7, 32'h42c15134};
test_weights[23192:23199] = '{32'hc28c8711, 32'h42c4c682, 32'hbfc7aac4, 32'hc195eaba, 32'h41acfe8b, 32'h428c184e, 32'hc240a03e, 32'h4265f57f};
test_bias[2899:2899] = '{32'h41d6f0a3};
test_output[2899:2899] = '{32'hc5061c8a};
test_input[23200:23207] = '{32'h4200a4fd, 32'h420f38dd, 32'hc1c92331, 32'hc26f3ef6, 32'h4285d9ae, 32'hc2a55f11, 32'h426c89b4, 32'hc2b77ed9};
test_weights[23200:23207] = '{32'h4158aa1c, 32'hc249c19a, 32'h4205ac56, 32'h41869995, 32'h40039dfb, 32'h42955b68, 32'h4296ea21, 32'hc1b689c0};
test_bias[2900:2900] = '{32'h41923c60};
test_output[2900:2900] = '{32'hc5278656};
test_input[23208:23215] = '{32'h42b677a1, 32'hc2041a44, 32'hc03ab7a2, 32'h42914eec, 32'hc1f09dba, 32'hc2a1f515, 32'hc2be59af, 32'h4204e3f1};
test_weights[23208:23215] = '{32'hc222d49d, 32'h4214ac82, 32'h42966120, 32'h42c3291f, 32'hc21a43e8, 32'hc2585d71, 32'hc2962ec4, 32'hc215f58f};
test_bias[2901:2901] = '{32'h42277026};
test_output[2901:2901] = '{32'h465190d9};
test_input[23216:23223] = '{32'h40f4de41, 32'h42168424, 32'h42550cc7, 32'h4284c775, 32'h42bd80d7, 32'h40e12b23, 32'h42195bc7, 32'hc20bc7fc};
test_weights[23216:23223] = '{32'h42986d97, 32'hc277f652, 32'h42309ed3, 32'hc2c4c1ad, 32'h425eb53e, 32'hc2007d5f, 32'h3ff56b78, 32'hc2bf72c0};
test_bias[2902:2902] = '{32'hc263588c};
test_output[2902:2902] = '{32'h451b2500};
test_input[23224:23231] = '{32'hc28140d3, 32'h4214c181, 32'hc25a674d, 32'hc23b8663, 32'hc23acd68, 32'h427e78ce, 32'h421e9dc9, 32'hc2b52961};
test_weights[23224:23231] = '{32'hc0482e54, 32'h415d6e9e, 32'hc176f8a4, 32'hc1177f0a, 32'h42a38e17, 32'hc2047429, 32'h426c1d7e, 32'hc1dbc628};
test_bias[2903:2903] = '{32'hc1c778cb};
test_output[2903:2903] = '{32'h445c83f0};
test_input[23232:23239] = '{32'h4292315b, 32'h4282d3ca, 32'h411d85f7, 32'h4204229c, 32'h4187651d, 32'h42b43004, 32'hc25a7a2b, 32'hc1af0384};
test_weights[23232:23239] = '{32'hc2819e83, 32'hc2b3843b, 32'hc2129de8, 32'h41ee10cd, 32'hc023d582, 32'hc2c05211, 32'h423c4867, 32'hc21ed8bd};
test_bias[2904:2904] = '{32'hc2aa88fd};
test_output[2904:2904] = '{32'hc6a001b3};
test_input[23240:23247] = '{32'hc249263a, 32'hc2b66425, 32'hc18a2dc2, 32'hc2359d9e, 32'h40c7f3f9, 32'h4081403c, 32'h42a336e1, 32'hc112345c};
test_weights[23240:23247] = '{32'hc26c5343, 32'hc2c6b8b3, 32'hc2b31ced, 32'hc22e7141, 32'hc2bfdeb9, 32'h41e5279b, 32'hc25f223b, 32'h4132bbcf};
test_bias[2905:2905] = '{32'h41d80004};
test_output[2905:2905] = '{32'h46234057};
test_input[23248:23255] = '{32'hc2565305, 32'h42954772, 32'hc287254a, 32'hc25baf8d, 32'hc2487894, 32'h42be1f34, 32'hc21a4ec0, 32'h413c5810};
test_weights[23248:23255] = '{32'hc12ff1f4, 32'hc23db6a2, 32'hc2bba4b4, 32'hc28a3eab, 32'h40808c59, 32'hc1a0baff, 32'h414c4eda, 32'h40199d62};
test_bias[2906:2906] = '{32'h42914c0d};
test_output[2906:2906] = '{32'h459252d1};
test_input[23256:23263] = '{32'h4255703c, 32'hc15251c8, 32'h40af42c9, 32'hc27946cc, 32'h428f5fc0, 32'h42b53c02, 32'h42c33d6c, 32'hc29428b3};
test_weights[23256:23263] = '{32'h4266aa5c, 32'h4251b57f, 32'hc28fc20f, 32'h42b86f05, 32'hc09a43cf, 32'hc1f15c0e, 32'h41ec1275, 32'hc278dd1a};
test_bias[2907:2907] = '{32'hc1d03e6b};
test_output[2907:2907] = '{32'h441dda4b};
test_input[23264:23271] = '{32'h424e2645, 32'h4273debb, 32'hc2c2e170, 32'hc2afc2a5, 32'h4204bf48, 32'hc23a28b8, 32'hc257aeed, 32'h4048b77a};
test_weights[23264:23271] = '{32'h421ff4c1, 32'h42a52cfc, 32'h4237a180, 32'h423ca913, 32'h4166ac86, 32'h42790bdb, 32'hc10d23cd, 32'h41768352};
test_bias[2908:2908] = '{32'hc0e05d57};
test_output[2908:2908] = '{32'hc5560425};
test_input[23272:23279] = '{32'h420d4c21, 32'h429aa179, 32'h429dbd82, 32'h429e440d, 32'hc227b96a, 32'hc21dbe56, 32'hc2211850, 32'hbf8d1164};
test_weights[23272:23279] = '{32'hc119b094, 32'hc2412d15, 32'h4295d068, 32'hc0baec93, 32'h41537bec, 32'h40e75c76, 32'hc2b5195c, 32'hc2bff1dc};
test_bias[2909:2909] = '{32'h426273cf};
test_output[2909:2909] = '{32'h4587b25c};
test_input[23280:23287] = '{32'h429badf8, 32'h42be669f, 32'hc1918a48, 32'hc286f262, 32'h42529171, 32'hc188e2d1, 32'hc2bc3b9d, 32'h419adf60};
test_weights[23280:23287] = '{32'h4221836e, 32'hc221e3af, 32'hc28046eb, 32'hc2968237, 32'hc108d008, 32'h41baee18, 32'hc2916057, 32'h41815a84};
test_bias[2910:2910] = '{32'h40dc59ef};
test_output[2910:2910] = '{32'h463916b4};
test_input[23288:23295] = '{32'h414686cd, 32'hbf8b95b9, 32'h4230bcd6, 32'h42c4d11b, 32'h4223979b, 32'h425d49e8, 32'h425d8f6c, 32'hc236693b};
test_weights[23288:23295] = '{32'h428ef1fc, 32'h41b7a3e2, 32'hc254d84f, 32'hc203de7c, 32'h4260eb73, 32'h42b0b679, 32'h41a1d826, 32'h42c481fd};
test_bias[2911:2911] = '{32'hc226f2a7};
test_output[2911:2911] = '{32'hc46ce7e2};
test_input[23296:23303] = '{32'hc145a1b5, 32'h42829db3, 32'h42b55ff8, 32'h423fd205, 32'h4249f157, 32'hc1536dc4, 32'hc1eff1fb, 32'h421a13f5};
test_weights[23296:23303] = '{32'hc275e6ef, 32'h415d6d96, 32'hc2547c42, 32'hc0101637, 32'hc2a7f16a, 32'h41974ee9, 32'hc029e48a, 32'hc288db73};
test_bias[2912:2912] = '{32'h409fa396};
test_output[2912:2912] = '{32'hc620fb0a};
test_input[23304:23311] = '{32'hc176a6ea, 32'hc21f33b8, 32'h42659bc8, 32'h42179bf4, 32'hc167686a, 32'h42b96cf6, 32'h4283f851, 32'h42b3c1d8};
test_weights[23304:23311] = '{32'hc205a673, 32'h41485fd8, 32'hc22d6c74, 32'hc2b68ace, 32'hc13225ec, 32'h42746d4d, 32'hc2980811, 32'h42036a73};
test_bias[2913:2913] = '{32'h4199ccd2};
test_output[2913:2913] = '{32'hc5064dbe};
test_input[23312:23319] = '{32'hc2079f9a, 32'h429ce851, 32'h42baa3b3, 32'h4232aea4, 32'h4204d9df, 32'h42a50970, 32'hc247290d, 32'h429417cd};
test_weights[23312:23319] = '{32'h419b5ece, 32'hc1c2274a, 32'h41ff3262, 32'h426816d0, 32'hc1974723, 32'hc2488c16, 32'hc2805408, 32'hc2946750};
test_bias[2914:2914] = '{32'h41f6629f};
test_output[2914:2914] = '{32'hc57bbdb1};
test_input[23320:23327] = '{32'h42a848ab, 32'h4275785a, 32'hc06bd5ba, 32'h41301e0e, 32'hc170fb51, 32'h4289faf4, 32'h4297c314, 32'hc2307a02};
test_weights[23320:23327] = '{32'h428bc980, 32'hc1571618, 32'h429d2c0b, 32'h428554dc, 32'hc1bede9b, 32'hc1eb9dbd, 32'hc08fac81, 32'h4183a3f7};
test_bias[2915:2915] = '{32'hc2a10055};
test_output[2915:2915] = '{32'h45278855};
test_input[23328:23335] = '{32'hc2425d9b, 32'hc2a5379c, 32'h4185f39e, 32'h4110e322, 32'hc2c53774, 32'h4210c99b, 32'hc20123eb, 32'hc09fda94};
test_weights[23328:23335] = '{32'h42379e69, 32'hc29264b5, 32'h40b06aa2, 32'hc1a0f725, 32'h427b861c, 32'hc26fa7b2, 32'h4282e579, 32'h42ae6046};
test_bias[2916:2916] = '{32'h4232649c};
test_output[2916:2916] = '{32'hc5df5813};
test_input[23336:23343] = '{32'hc17e9906, 32'h41871b21, 32'h41c22e4a, 32'h41cc5c61, 32'h42905c03, 32'hc2a1a703, 32'hc234c9ae, 32'hc2659458};
test_weights[23336:23343] = '{32'hc23ea93f, 32'h4113a5ce, 32'hc0b5d235, 32'hc14a74eb, 32'h416c6f83, 32'hc2984935, 32'h42a81e9b, 32'hc29ca142};
test_bias[2917:2917] = '{32'hc2acb092};
test_output[2917:2917] = '{32'h46016da3};
test_input[23344:23351] = '{32'h42c77de9, 32'h420a1dcf, 32'hc2c441f0, 32'hc2a42251, 32'h42ab9282, 32'h4263d3b6, 32'hc29a7d8d, 32'hc158b31e};
test_weights[23344:23351] = '{32'hc2c04b2b, 32'h40a28abb, 32'h4293d689, 32'hc28aa687, 32'h42ab999d, 32'hc2863b83, 32'h41fc147a, 32'h423f3f1b};
test_bias[2918:2918] = '{32'h42b37b4b};
test_output[2918:2918] = '{32'hc62304cf};
test_input[23352:23359] = '{32'hc1f88e3b, 32'h41bc135c, 32'hc22da16c, 32'h421b582f, 32'h423ca8e2, 32'h42945932, 32'h42b26489, 32'hc14a7529};
test_weights[23352:23359] = '{32'h42bb336e, 32'hc1ff4509, 32'hc251724c, 32'hc2be0ecc, 32'hc2934570, 32'h4159411b, 32'h4224c8ce, 32'hc15f6dc8};
test_bias[2919:2919] = '{32'h4295eb9f};
test_output[2919:2919] = '{32'hc561f94c};
test_input[23360:23367] = '{32'hc0910ca8, 32'h419ab3f5, 32'hc2116cb0, 32'hc1ab093f, 32'h4226d2c1, 32'hc26c46b7, 32'h41ef1f2d, 32'hc1bf42b5};
test_weights[23360:23367] = '{32'h41b90218, 32'h41bbb8b6, 32'h42353734, 32'h42b5f283, 32'hc2699652, 32'hc2622093, 32'hc250a9c3, 32'h42892a72};
test_bias[2920:2920] = '{32'hc2c2ab8f};
test_output[2920:2920] = '{32'hc5b01c5b};
test_input[23368:23375] = '{32'h42b87076, 32'hc1fe8b08, 32'hc010b008, 32'h428f2d5b, 32'hc07343cb, 32'hc2280938, 32'h429dec69, 32'hc125c144};
test_weights[23368:23375] = '{32'hc2b61edf, 32'hc259a439, 32'hc1b4311c, 32'h4116b3f2, 32'h4236abb0, 32'hc278ccec, 32'hc20e1517, 32'hc2129505};
test_bias[2921:2921] = '{32'h42813d7f};
test_output[2921:2921] = '{32'hc5b731f9};
test_input[23376:23383] = '{32'hc2524799, 32'h4279acd8, 32'hc258f555, 32'hc22d0ed9, 32'hc29a77c9, 32'h42b277d9, 32'h4240392d, 32'h423127ac};
test_weights[23376:23383] = '{32'hc212f231, 32'h42045109, 32'hc2655af1, 32'h4218c4b2, 32'hc2028d60, 32'hc2b636e2, 32'hc29109a3, 32'h42679e0e};
test_bias[2922:2922] = '{32'hc2997791};
test_output[2922:2922] = '{32'hc4901371};
test_input[23384:23391] = '{32'h425cabf3, 32'h4283c03e, 32'hc134f25b, 32'h425c5de0, 32'hc2b86b9a, 32'h427d6a55, 32'hc19b8d64, 32'hc216c421};
test_weights[23384:23391] = '{32'hc14f1e43, 32'hc284be66, 32'h4198972a, 32'h40952821, 32'h428be433, 32'hc220c2f8, 32'hc265e2bb, 32'hc18e69f2};
test_bias[2923:2923] = '{32'h429b37c5};
test_output[2923:2923] = '{32'hc63e3ccd};
test_input[23392:23399] = '{32'h42725986, 32'hc29dbe18, 32'h3f82ffad, 32'h418e9112, 32'h41a0c6c0, 32'h428e12af, 32'hc2a9d9b5, 32'h42c2f214};
test_weights[23392:23399] = '{32'h423aced3, 32'hc2764d09, 32'h409e7616, 32'hc253bf2c, 32'hc13fc3b5, 32'hc0f3e55c, 32'hc216a080, 32'hc0769628};
test_bias[2924:2924] = '{32'hbfbd63eb};
test_output[2924:2924] = '{32'h460949c6};
test_input[23400:23407] = '{32'h41f9a947, 32'h42361377, 32'h42464700, 32'hc2c34a11, 32'h429f9a97, 32'h429f04dd, 32'h42654293, 32'hc288ce6c};
test_weights[23400:23407] = '{32'h4283eaa0, 32'h423acc78, 32'hc28bf6ff, 32'hc25a957f, 32'h4296cd23, 32'h424ebe2c, 32'h4011b2a6, 32'hc1b05d8c};
test_bias[2925:2925] = '{32'h42c241f9};
test_output[2925:2925] = '{32'h468bf284};
test_input[23408:23415] = '{32'h422be0c7, 32'hc25094e1, 32'h3e9a48d5, 32'h4196ec86, 32'hc2a3e0f5, 32'hc1f30b3f, 32'h4299e6ce, 32'h42335992};
test_weights[23408:23415] = '{32'hc262a080, 32'hc2b0407b, 32'hc2c32cef, 32'h40a08c5d, 32'hc20cc902, 32'hc2bbb2e7, 32'hc1bd2747, 32'hc23b04b6};
test_bias[2926:2926] = '{32'h428e6292};
test_output[2926:2926] = '{32'h4580a526};
test_input[23416:23423] = '{32'h428ed22e, 32'hc1d29bf9, 32'h428b9869, 32'h428ec142, 32'h418eeb0c, 32'hc22fc123, 32'hc261f000, 32'hc1c3742f};
test_weights[23416:23423] = '{32'hc26446a5, 32'hc0329125, 32'h41ad5caf, 32'h42216f60, 32'hc1d08fba, 32'hc2ad40d7, 32'h429269f4, 32'hc2137333};
test_bias[2927:2927] = '{32'hc195a941};
test_output[2927:2927] = '{32'h43ef5f03};
test_input[23424:23431] = '{32'h4200672a, 32'hc0e2bd0a, 32'h3eb7caa4, 32'hc2872518, 32'h42b46185, 32'hc129e3c8, 32'hc220f7ea, 32'h42a141e6};
test_weights[23424:23431] = '{32'hc265063e, 32'h4242fd83, 32'hc1ff3876, 32'hc2b82ddd, 32'hc22d86a0, 32'hc24573bd, 32'hc19f7b73, 32'hc2a691b3};
test_bias[2928:2928] = '{32'hc2098243};
test_output[2928:2928] = '{32'hc5a5de93};
test_input[23432:23439] = '{32'hc0f1dca8, 32'h41bf2faa, 32'h429b349e, 32'h4225cc97, 32'h42063331, 32'hc2c3accd, 32'h426012d9, 32'h403ac21f};
test_weights[23432:23439] = '{32'h428e0cea, 32'hc2c0573d, 32'h40de82eb, 32'h4205913d, 32'h4297e1e6, 32'hc23b72a7, 32'h42bce4fe, 32'hc27e7521};
test_bias[2929:2929] = '{32'h4055bc96};
test_output[2929:2929] = '{32'h463106f7};
test_input[23440:23447] = '{32'hc1811fe3, 32'h42af9ada, 32'hc2962cb1, 32'hc2b3d5e4, 32'hc297ac6c, 32'hc1e91e0b, 32'h42a09818, 32'hc2570f3c};
test_weights[23440:23447] = '{32'hc2a58974, 32'hc29097b9, 32'hc2c5372c, 32'h428d0175, 32'hc0bd86f9, 32'hc269ba60, 32'h42ac98b4, 32'hc2804d15};
test_bias[2930:2930] = '{32'h428b602f};
test_output[2930:2930] = '{32'h460733ca};
test_input[23448:23455] = '{32'h427dddc9, 32'h42889918, 32'hc273786d, 32'h41da6af4, 32'h42952cdb, 32'h42276257, 32'h41f567d9, 32'hc2804ea9};
test_weights[23448:23455] = '{32'hc257294b, 32'h427e4843, 32'hc21e40d4, 32'hc2312591, 32'hc0ca2734, 32'hc2b98257, 32'hbfc851c1, 32'h41cd3671};
test_bias[2931:2931] = '{32'hc2a7eaca};
test_output[2931:2931] = '{32'hc57a34b0};
test_input[23456:23463] = '{32'hc0b19933, 32'hc2b9be83, 32'h427ce575, 32'hc2c62ffb, 32'hc28f0a04, 32'hc281b5cc, 32'h41a1772a, 32'hc1d14b4b};
test_weights[23456:23463] = '{32'hc04e0012, 32'hc2570d14, 32'hc14db6cd, 32'h4299ac04, 32'hc1c8a79a, 32'hc2ba020e, 32'hc1bae61a, 32'h41b404e5};
test_bias[2932:2932] = '{32'hc1c34862};
test_output[2932:2932] = '{32'h454fd119};
test_input[23464:23471] = '{32'h416e5a1d, 32'h4216b0cc, 32'h41b9cd90, 32'h42c65316, 32'hc217dc51, 32'hc246197d, 32'h42a7858e, 32'h42a401b9};
test_weights[23464:23471] = '{32'h420a39d3, 32'h42af664e, 32'h42832544, 32'h42b45bf8, 32'hc11a6b7f, 32'hc24a9cd3, 32'h42445ee5, 32'hc2883d7c};
test_bias[2933:2933] = '{32'h42aea0ac};
test_output[2933:2933] = '{32'h4676714e};
test_input[23472:23479] = '{32'h4231ab09, 32'hc2bd8f56, 32'hc284efa0, 32'h42600f79, 32'hc1b8ff44, 32'h41802eb6, 32'hc079e80a, 32'hc2663e82};
test_weights[23472:23479] = '{32'hc207f6b8, 32'h423f2fd0, 32'h41db5faf, 32'h41c6799b, 32'h41d9c591, 32'h41db90bf, 32'hc08a02a3, 32'h42a4cc70};
test_bias[2934:2934] = '{32'hc1fcc2af};
test_output[2934:2934] = '{32'hc632718b};
test_input[23480:23487] = '{32'h3e7d6de5, 32'h42bba694, 32'hc24fb9e0, 32'hc2b93f48, 32'hc28f15f9, 32'h42b311b5, 32'hc27c6cc1, 32'hc256adcc};
test_weights[23480:23487] = '{32'hc21068bf, 32'hc298e509, 32'hc2632f98, 32'hc2bdf583, 32'hc2c13cd9, 32'hc105fbe4, 32'hc28bb3d2, 32'h41f349f9};
test_bias[2935:2935] = '{32'h41f92492};
test_output[2935:2935] = '{32'h46537b9c};
test_input[23488:23495] = '{32'h416b516b, 32'h42425afc, 32'hc28f1d10, 32'hc2aed31e, 32'hc2bc8dc7, 32'h41235f30, 32'h428d9d47, 32'hc2afc614};
test_weights[23488:23495] = '{32'hc280c7b2, 32'hc0caed87, 32'h4241d84f, 32'hc2b586f3, 32'hc27a90e7, 32'hc1242cae, 32'h42900cd3, 32'h4212fb2c};
test_bias[2936:2936] = '{32'h41f9ff47};
test_output[2936:2936] = '{32'h462a8652};
test_input[23496:23503] = '{32'h41a0fb9f, 32'h40f3d97c, 32'h424574b3, 32'h429ade75, 32'hc2935319, 32'hc2078e54, 32'h4223f6ad, 32'h41a37337};
test_weights[23496:23503] = '{32'h41b17b97, 32'hc1512f04, 32'hc2980798, 32'hc1e6bf4f, 32'h425cc7d8, 32'hc23eeb95, 32'h429d9a31, 32'h4290ac23};
test_bias[2937:2937] = '{32'h4195c4aa};
test_output[2937:2937] = '{32'hc5520925};
test_input[23504:23511] = '{32'hc128bae0, 32'h42a2833a, 32'hc202981a, 32'hc2c2ad36, 32'h4177e75a, 32'hc2062671, 32'hc2bf73fc, 32'hc0d74d7b};
test_weights[23504:23511] = '{32'h41e386c0, 32'hc28c6b2d, 32'h412aa267, 32'hc2b0d949, 32'h40c8a101, 32'hc244064b, 32'h4296fbfd, 32'h42a812b4};
test_bias[2938:2938] = '{32'h42b98fdb};
test_output[2938:2938] = '{32'hc5678886};
test_input[23512:23519] = '{32'hc29fd4b1, 32'hc280987f, 32'hc27fb4d9, 32'hc16ec2c0, 32'hc2ab4f3f, 32'hc2292eaa, 32'h42444b43, 32'h428f2c69};
test_weights[23512:23519] = '{32'hc291e13c, 32'hc2abf733, 32'h42c092d5, 32'hc24a8f87, 32'hc27a74e1, 32'hc1b116cf, 32'h42a3ae3b, 32'hc19310d2};
test_bias[2939:2939] = '{32'hc245d313};
test_output[2939:2939] = '{32'h4668f080};
test_input[23520:23527] = '{32'h42756b38, 32'hbf55e23f, 32'h42400146, 32'h4246e2e3, 32'hc2928247, 32'h42a00a77, 32'h42409245, 32'h4183258a};
test_weights[23520:23527] = '{32'hc20440c6, 32'h41dc79b6, 32'h4043214b, 32'h429648c8, 32'h423b2df2, 32'hc1b557a9, 32'hc10c2801, 32'h41f617fc};
test_bias[2940:2940] = '{32'h4286b230};
test_output[2940:2940] = '{32'hc54bcfb0};
test_input[23528:23535] = '{32'h41c2eb24, 32'h427b55f0, 32'hbf89ef3c, 32'hc1967fe0, 32'hc2322295, 32'h41598e46, 32'h41a66e77, 32'h4288052f};
test_weights[23528:23535] = '{32'hc29a22ee, 32'hc1b3cf2f, 32'hc2900903, 32'hc2b91793, 32'hc25ebef8, 32'h42a9aced, 32'hc2c3f920, 32'h4293b544};
test_bias[2941:2941] = '{32'hc2b195fb};
test_output[2941:2941] = '{32'h459e0cee};
test_input[23536:23543] = '{32'hc2b89e08, 32'h419512bc, 32'h42a621cb, 32'hc2bb3df0, 32'h425829ff, 32'hc2b379b5, 32'h42388e9e, 32'h42520177};
test_weights[23536:23543] = '{32'hc2bbd070, 32'hc2a6335d, 32'h42a316b0, 32'hc293b6ee, 32'hc0f51d23, 32'hc165f1d2, 32'hc239c928, 32'h4166cd3c};
test_bias[2942:2942] = '{32'h42ae8dd3};
test_output[2942:2942] = '{32'h469f42d8};
test_input[23544:23551] = '{32'h3f66b81a, 32'hc27d0094, 32'hc233dfaa, 32'hc22c7f6e, 32'h4162c223, 32'h4257f834, 32'h42acd8c1, 32'h42b33b54};
test_weights[23544:23551] = '{32'h42aed25d, 32'h4227035a, 32'h426c0663, 32'h4023ea96, 32'hc2272533, 32'hc216bdf3, 32'hc25a311f, 32'hc2977c7a};
test_bias[2943:2943] = '{32'hc20f67fd};
test_output[2943:2943] = '{32'hc698459c};
test_input[23552:23559] = '{32'hc17e6221, 32'hc1d73be4, 32'h4244e5cd, 32'hc271455b, 32'h42aa7cd5, 32'h40c058b4, 32'hc22157a7, 32'hc2734fc8};
test_weights[23552:23559] = '{32'h418f1be4, 32'h42494ecc, 32'hc1073ad3, 32'h4108661d, 32'h428f2672, 32'h41f21c9e, 32'h41ec65dd, 32'h40e29be7};
test_bias[2944:2944] = '{32'hc288beef};
test_output[2944:2944] = '{32'h44fcf19c};
test_input[23560:23567] = '{32'hc134c0b9, 32'hc0185213, 32'h42c79229, 32'h4127368b, 32'h42c56c04, 32'hc094d4c9, 32'h42993a37, 32'h41b74ca5};
test_weights[23560:23567] = '{32'h40aeeed5, 32'hc1922ddc, 32'h4175bf3c, 32'hc1d999a5, 32'hc2c5bc10, 32'hc209bd67, 32'hc19f38c5, 32'hc03eac80};
test_bias[2945:2945] = '{32'hc298738e};
test_output[2945:2945] = '{32'hc61cd964};
test_input[23568:23575] = '{32'hc2016086, 32'h40ad300b, 32'hc2951ad9, 32'hc2be794f, 32'hc29ee5bc, 32'hc29b117d, 32'hc1219168, 32'h4284c541};
test_weights[23568:23575] = '{32'hc2b5b6cb, 32'hc26ebe4c, 32'hc1389219, 32'hc27e4fa8, 32'hbfb57dd6, 32'h4231c16e, 32'hc2b4c52c, 32'hc2ab70b9};
test_bias[2946:2946] = '{32'hc1f3777a};
test_output[2946:2946] = '{32'h44adaf63};
test_input[23576:23583] = '{32'hc2828f4d, 32'h42ad2c06, 32'hc22b7c2a, 32'hc291160e, 32'hc281f723, 32'hc172f8e1, 32'hc12601d3, 32'h4296cece};
test_weights[23576:23583] = '{32'hc0d79c92, 32'h41fa0e9e, 32'hc2c31de7, 32'hc216857c, 32'hc25cbd43, 32'hc2407b48, 32'h4251e090, 32'hc246d393};
test_bias[2947:2947] = '{32'hc1f52bbb};
test_output[2947:2947] = '{32'h461d10f7};
test_input[23584:23591] = '{32'hc2c6daad, 32'h413762fd, 32'h42b935f2, 32'h42315681, 32'h3f8725d9, 32'hc24fe473, 32'h4261d7dc, 32'h41f6a685};
test_weights[23584:23591] = '{32'h413bcaaf, 32'hc2591fb1, 32'h42943848, 32'hc10de5dd, 32'hc1697b21, 32'hc287cb8a, 32'h42a13fe0, 32'h409bab1d};
test_bias[2948:2948] = '{32'h4299ddcd};
test_output[2948:2948] = '{32'h464ab4a2};
test_input[23592:23599] = '{32'h421572aa, 32'hc194958d, 32'h42b1da8e, 32'h422b5c92, 32'h40fae34b, 32'hc2c4ca7e, 32'h42c22667, 32'hc2b3909b};
test_weights[23592:23599] = '{32'h42527eaf, 32'h426f5500, 32'hc1f43d5c, 32'h42265f55, 32'hc2880b7d, 32'h4241d502, 32'h42ac57cf, 32'h429fbc48};
test_bias[2949:2949] = '{32'hc2a685d7};
test_output[2949:2949] = '{32'hc58563bf};
test_input[23600:23607] = '{32'h42b1f3e0, 32'hc1b95f58, 32'h4100d547, 32'h42c15702, 32'h42ab2461, 32'hc2990eb5, 32'h426786de, 32'hc286b20b};
test_weights[23600:23607] = '{32'h428874dc, 32'hc28e7bee, 32'hc0c8584a, 32'hc0e7cc99, 32'h4287649c, 32'h42a2a5dc, 32'hc22097f7, 32'hc10491fe};
test_bias[2950:2950] = '{32'h41b4b5da};
test_output[2950:2950] = '{32'h4595e689};
test_input[23608:23615] = '{32'hc24acc80, 32'h410a824b, 32'h4220502d, 32'hc1012d9c, 32'hc29a6c23, 32'h426f13ce, 32'h4282db80, 32'hc2c7f9cb};
test_weights[23608:23615] = '{32'hc0cffb46, 32'hc2a5d4b0, 32'hc2555ccd, 32'h420cf437, 32'h4265130d, 32'h4130bbda, 32'h40e69ff7, 32'h42b2b363};
test_bias[2951:2951] = '{32'hc2b0e5db};
test_output[2951:2951] = '{32'hc66c4bfe};
test_input[23616:23623] = '{32'hc27afef9, 32'h42ba72d6, 32'h421e6079, 32'hc2460f27, 32'hc05318bb, 32'hc2befad5, 32'h41d5b57a, 32'hc214022a};
test_weights[23616:23623] = '{32'h42a06e67, 32'hc2492a24, 32'hc25a9fd2, 32'hc1f244d6, 32'hc2b650b4, 32'hc1ac1cab, 32'h42c75545, 32'hc2864ef8};
test_bias[2952:2952] = '{32'hc2a4be85};
test_output[2952:2952] = '{32'hc5396699};
test_input[23624:23631] = '{32'hc184b959, 32'hc2b0eda3, 32'h42663751, 32'hc27dfc9a, 32'h421793c8, 32'hc1d7b23d, 32'h429f8ef1, 32'h42529af6};
test_weights[23624:23631] = '{32'hc23e9abb, 32'hc1cc03f9, 32'h42a40d95, 32'h42a121d6, 32'h42904f17, 32'hc21d6a50, 32'hc266f239, 32'hc0fc7804};
test_bias[2953:2953] = '{32'h4232d430};
test_output[2953:2953] = '{32'h44b7c8d3};
test_input[23632:23639] = '{32'hc10a92fa, 32'hc190e965, 32'h41a2d929, 32'hc1b4eeda, 32'h41d7fecc, 32'hc2427cf5, 32'hc1e4c17e, 32'h42a05d15};
test_weights[23632:23639] = '{32'h428b577b, 32'h42a5ecb4, 32'hc1c782db, 32'hc2a3b61b, 32'hc296d678, 32'h41caa808, 32'hc2815e31, 32'hc249f54e};
test_bias[2954:2954] = '{32'h4196ec89};
test_output[2954:2954] = '{32'hc5c2130a};
test_input[23640:23647] = '{32'h4233bc3d, 32'h41b962b0, 32'h429c1ce6, 32'hc20e5ba8, 32'h4270b53b, 32'h42674d58, 32'hc283cfef, 32'hc22a5645};
test_weights[23640:23647] = '{32'hc186f958, 32'h41e2a9c7, 32'hc2b78e31, 32'hc29ee36d, 32'h426821d3, 32'hc283d01a, 32'hc1492013, 32'hc191d99d};
test_bias[2955:2955] = '{32'hc2723d38};
test_output[2955:2955] = '{32'hc548c912};
test_input[23648:23655] = '{32'hc21ff503, 32'hc218e631, 32'hc179d6c3, 32'h42b5d9a5, 32'h42914d4d, 32'hc2b1d185, 32'h4281404c, 32'h423c72eb};
test_weights[23648:23655] = '{32'hc2c314a9, 32'h41ab0233, 32'h3ed85d22, 32'hc23524b4, 32'h40480fd2, 32'hc296c1b2, 32'h4193383d, 32'hc2a75871};
test_bias[2956:2956] = '{32'h4294caff};
test_output[2956:2956] = '{32'h45489d79};
test_input[23656:23663] = '{32'hc28b7ad3, 32'h40dd41ca, 32'hc2036559, 32'hc21f5dd7, 32'h4295f6b8, 32'h42627f0f, 32'hc0e3b932, 32'hc26f1381};
test_weights[23656:23663] = '{32'hc17566d7, 32'hc2777809, 32'h42b93153, 32'hc0047916, 32'h4291ad1d, 32'h4227d11e, 32'h429560db, 32'hc13ea1d4};
test_bias[2957:2957] = '{32'h4291dd7e};
test_output[2957:2957] = '{32'h45b46abd};
test_input[23664:23671] = '{32'hc2c5619d, 32'h426813a3, 32'hc14e26f6, 32'h4281ef7d, 32'h42c12f70, 32'h42a5fb4a, 32'h420f6d54, 32'hc1a83e18};
test_weights[23664:23671] = '{32'hc2114544, 32'hc17e1ec7, 32'hc22615e6, 32'hc2972c51, 32'h4280d87c, 32'hc247ca32, 32'hc21033e0, 32'hc2aa4f43};
test_bias[2958:2958] = '{32'h42612dd4};
test_output[2958:2958] = '{32'h4465c4c8};
test_input[23672:23679] = '{32'h405cab3c, 32'h423aec49, 32'hc1a7b434, 32'hc1962e46, 32'h429c469e, 32'hc23b6688, 32'h422d06c8, 32'h42444e10};
test_weights[23672:23679] = '{32'hc29edda8, 32'hc26743ac, 32'h4280d0b7, 32'h42a6131a, 32'hc21e0feb, 32'hc23ed398, 32'h42956622, 32'h414e3ba9};
test_bias[2959:2959] = '{32'h42909586};
test_output[2959:2959] = '{32'hc52f129a};
test_input[23680:23687] = '{32'hc1e7ced4, 32'hc2c7a57a, 32'hc201fac0, 32'hc27ff30d, 32'h41239c99, 32'h4291c902, 32'h40ec0b41, 32'hc27ecfa8};
test_weights[23680:23687] = '{32'h423a0024, 32'h41f6c943, 32'hc26cc923, 32'h42c38f6e, 32'h42b29e5b, 32'h42c2775f, 32'h428dc52b, 32'h4290c8dd};
test_bias[2960:2960] = '{32'hc2b4e3bb};
test_output[2960:2960] = '{32'hc59a51a4};
test_input[23688:23695] = '{32'h42b64df4, 32'h42c42316, 32'hc294b41c, 32'h429e62b6, 32'hc1805e11, 32'h428bd2b3, 32'h42562f3f, 32'h41747148};
test_weights[23688:23695] = '{32'hc21ec00f, 32'hc270d09a, 32'h42ad6c0c, 32'h413909cf, 32'h42a2210d, 32'h41c47d40, 32'hc0cf34df, 32'hc2aef8c1};
test_bias[2961:2961] = '{32'hc1ae7f6d};
test_output[2961:2961] = '{32'hc67f56e5};
test_input[23696:23703] = '{32'hc29d52e6, 32'h429a68f6, 32'hc1827f8a, 32'h3f1df348, 32'hc09991f1, 32'h416c5b45, 32'hc1fde995, 32'hc2a2a3ff};
test_weights[23696:23703] = '{32'h4293efb9, 32'hc23a901f, 32'h423ed799, 32'hc2265687, 32'hc1ee8fa2, 32'hc263a40c, 32'h40d82426, 32'h41f02504};
test_bias[2962:2962] = '{32'hc059b7a8};
test_output[2962:2962] = '{32'hc6542eff};
test_input[23704:23711] = '{32'hc21ad076, 32'hc2a4601e, 32'h41113e41, 32'hc1b19d2f, 32'h42acb80d, 32'hc29169d5, 32'hc23d5569, 32'h4071547f};
test_weights[23704:23711] = '{32'h411a4fe1, 32'hc24e4cc9, 32'hc2328af3, 32'h40d92545, 32'h4204c5cb, 32'h4242adb9, 32'hc2953926, 32'hc23c912f};
test_bias[2963:2963] = '{32'h42a00ff3};
test_output[2963:2963] = '{32'h45bdbc44};
test_input[23712:23719] = '{32'hc24654bf, 32'hc28f70b9, 32'hc2a3e0cb, 32'hc191490f, 32'hc212c223, 32'h4240cb9e, 32'h42aa8143, 32'hc1ec1cb5};
test_weights[23712:23719] = '{32'h427d94c4, 32'h42824bd4, 32'h41a09c81, 32'h4120b4e7, 32'h425c0f97, 32'hc1d33782, 32'hc2a05187, 32'h40dd05db};
test_bias[2964:2964] = '{32'h420f0afe};
test_output[2964:2964] = '{32'hc69bc032};
test_input[23720:23727] = '{32'hc29a1b64, 32'h4225b5eb, 32'hc1c63cb7, 32'h4212323a, 32'h42b3feb2, 32'h422d0bce, 32'hc2156511, 32'hc28c1c0a};
test_weights[23720:23727] = '{32'h4269c7e2, 32'hc24dbd0b, 32'hc2b6bf47, 32'hbee5fa2e, 32'h41cae588, 32'h41f50b1b, 32'hc21e8328, 32'hc1f94e17};
test_bias[2965:2965] = '{32'hbfea196e};
test_output[2965:2965] = '{32'h453428fa};
test_input[23728:23735] = '{32'hc1f01d2f, 32'hc1fce7c5, 32'h4276a5b1, 32'hc2b63f7c, 32'h41d39568, 32'h42baf252, 32'h4287d1d4, 32'hc2aa1ff1};
test_weights[23728:23735] = '{32'h420f56a2, 32'hc280a9d3, 32'h428d88cd, 32'hc220720b, 32'h42c75c1f, 32'h42677bc3, 32'hc2481cb3, 32'h429274ac};
test_bias[2966:2966] = '{32'h4256dc41};
test_output[2966:2966] = '{32'h45e8d01a};
test_input[23736:23743] = '{32'h42bacbf2, 32'hc2852879, 32'h418baa30, 32'hc2a3438b, 32'hc181ccb8, 32'h4224f4bd, 32'hc29c6501, 32'h4298abf3};
test_weights[23736:23743] = '{32'h42ad97a0, 32'hc19924b7, 32'h41e12706, 32'h40da4482, 32'h42c77a2a, 32'hc297ae2c, 32'hc2b0f975, 32'hc25748fc};
test_bias[2967:2967] = '{32'h42b28776};
test_output[2967:2967] = '{32'h45e9709f};
test_input[23744:23751] = '{32'hc2b28c5b, 32'hc2820a45, 32'h41fa3f6c, 32'h428ef226, 32'h4278b75d, 32'h42839ea2, 32'h422c5eeb, 32'h423b4b48};
test_weights[23744:23751] = '{32'hc2974530, 32'h423333ee, 32'hc2934ab3, 32'hc22b1dda, 32'hc2965b5c, 32'hc28d82fe, 32'h42a7ca9c, 32'h408efafe};
test_bias[2968:2968] = '{32'hc102c7d8};
test_output[2968:2968] = '{32'hc5dbe497};
test_input[23752:23759] = '{32'h42b9b3a9, 32'hc2b72031, 32'hc2aec7b7, 32'h417a8427, 32'h412993b7, 32'hc2c63aab, 32'hc27f245a, 32'h4261adaf};
test_weights[23752:23759] = '{32'hc2a50885, 32'hc05bc5f0, 32'hc08c2541, 32'hc26e193f, 32'h42c285a5, 32'hc262ad59, 32'h42aea630, 32'h41fa8f54};
test_bias[2969:2969] = '{32'h4289a97b};
test_output[2969:2969] = '{32'hc59bb93e};
test_input[23760:23767] = '{32'hc16d37cd, 32'h429f889a, 32'hc2740081, 32'hc2a35acd, 32'h4252957a, 32'h41a50d07, 32'h417f4927, 32'hc15eabac};
test_weights[23760:23767] = '{32'h426b8acd, 32'hc221164d, 32'hc21f3a34, 32'hc200ff3d, 32'hc2391335, 32'hc110c9a0, 32'h421d0fff, 32'h41b57d82};
test_bias[2970:2970] = '{32'h424bf44e};
test_output[2970:2970] = '{32'hc4a07d8f};
test_input[23768:23775] = '{32'h4290beb3, 32'hc23adfdc, 32'h426d9feb, 32'h4214f4cd, 32'h420636f5, 32'h3f6c1f44, 32'hc1426928, 32'h417abdef};
test_weights[23768:23775] = '{32'hc2c2a112, 32'hc2a86446, 32'hc2893c32, 32'hc1647fa1, 32'hc2a564e9, 32'h42bd08f2, 32'hc2a399c1, 32'hbf64bed6};
test_bias[2971:2971] = '{32'h42617592};
test_output[2971:2971] = '{32'hc6126351};
test_input[23776:23783] = '{32'hc2813bf6, 32'h42a03ef7, 32'h42b4975a, 32'hc2b4dbf6, 32'hc28ed9ea, 32'h42b0e3f6, 32'hc2234de3, 32'hc1a5c01e};
test_weights[23776:23783] = '{32'h4255fc41, 32'hc20ee6cc, 32'hc2985043, 32'h42aa9d89, 32'hc2719de5, 32'h3f766005, 32'hc1f8b120, 32'h41ad9e72};
test_bias[2972:2972] = '{32'hc08eb101};
test_output[2972:2972] = '{32'hc6753e6d};
test_input[23784:23791] = '{32'hc11c6196, 32'h416bdc42, 32'hc27069e3, 32'hc2a80d18, 32'hc1f35775, 32'hc2c77821, 32'hc2487822, 32'h4126f05f};
test_weights[23784:23791] = '{32'h429c41db, 32'hc27d6cad, 32'h42ba1a7e, 32'h42884de5, 32'h41e20507, 32'hc2687326, 32'h4236bee0, 32'hc2bdbf76};
test_bias[2973:2973] = '{32'hc222511d};
test_output[2973:2973] = '{32'hc632220b};
test_input[23792:23799] = '{32'hc25de07e, 32'hc21f9bdb, 32'h4277142f, 32'hc27ca97e, 32'h421b6e32, 32'h41585bf7, 32'h42ac5dde, 32'h4221410a};
test_weights[23792:23799] = '{32'hc2920130, 32'hc2b60522, 32'hc075f672, 32'h414ac933, 32'hc2a98903, 32'hc2abcee7, 32'h429b1683, 32'hc208b991};
test_bias[2974:2974] = '{32'hc2bcaa55};
test_output[2974:2974] = '{32'h45e730fc};
test_input[23800:23807] = '{32'h41423123, 32'h41c1ee59, 32'hc1d6bd6f, 32'hc179180f, 32'hc2575d3c, 32'h42ad7d1b, 32'h42077f75, 32'hc2905b01};
test_weights[23800:23807] = '{32'h40350ad7, 32'h427ef53f, 32'h42c49396, 32'h4287912d, 32'h426c2e21, 32'h428d364f, 32'hc18e7177, 32'hc2c4f9da};
test_bias[2975:2975] = '{32'hc298645f};
test_output[2975:2975] = '{32'h45e2e67d};
test_input[23808:23815] = '{32'hc21f685b, 32'h4118e1c7, 32'hc26b4f18, 32'h4197ac88, 32'h41cdf697, 32'hc291de24, 32'h419627b7, 32'h4163a983};
test_weights[23808:23815] = '{32'hc19de65a, 32'h4121e7b4, 32'hc23fd010, 32'hc228198c, 32'hc283fa30, 32'h421068f5, 32'h42794798, 32'h41d3a090};
test_bias[2976:2976] = '{32'hc24393a3};
test_output[2976:2976] = '{32'h429158ab};
test_input[23816:23823] = '{32'hc1d02783, 32'hc17ecd59, 32'hc14da5be, 32'h42844386, 32'hbf527bd2, 32'hc2a845ba, 32'h42afe8a7, 32'h4233f4d4};
test_weights[23816:23823] = '{32'hc10f15f2, 32'h42ba6b31, 32'hc28828be, 32'h425498a0, 32'h42935f68, 32'h42af1b1d, 32'h4299d342, 32'h4281f009};
test_bias[2977:2977] = '{32'h40e0dc10};
test_output[2977:2977] = '{32'h45a8ef94};
test_input[23824:23831] = '{32'hc1eb3dfb, 32'h40f3827f, 32'hc2b3f4b6, 32'hc2320965, 32'h42a6d4b9, 32'hc05861c9, 32'hc180c8c0, 32'hc28de026};
test_weights[23824:23831] = '{32'h41b51405, 32'hc1faf6c7, 32'hc2867be1, 32'h41ca36ce, 32'hc12f5f8f, 32'hc2a633ab, 32'h4278ea22, 32'h42bb0375};
test_bias[2978:2978] = '{32'h41887f8f};
test_output[2978:2978] = '{32'hc584320b};
test_input[23832:23839] = '{32'h4295c763, 32'hc1cb0927, 32'h4199fe7e, 32'hc28e395b, 32'h41a1ec3a, 32'hc2c4dafc, 32'h418fbbf2, 32'h429d3215};
test_weights[23832:23839] = '{32'hc2c7b4bb, 32'h41a89a2e, 32'hc2320d63, 32'hc193da05, 32'hc29e4e19, 32'hc22528a1, 32'h4216dfdb, 32'hc2a8fbc4};
test_bias[2979:2979] = '{32'hc1a7bdf9};
test_output[2979:2979] = '{32'hc62d1653};
test_input[23840:23847] = '{32'h4235945b, 32'h427fbe7d, 32'h41ffa48d, 32'h42c1f336, 32'h427a28f9, 32'h41bcc848, 32'h427d9f78, 32'hc2a3b260};
test_weights[23840:23847] = '{32'h422e66e3, 32'hc18999f8, 32'h4170bc4c, 32'h42bf3a29, 32'hc2b7300b, 32'h416158ad, 32'h4214e168, 32'h428a14d1};
test_bias[2980:2980] = '{32'h418f3878};
test_output[2980:2980] = '{32'h44f5712c};
test_input[23848:23855] = '{32'hc260b1a9, 32'hc2c3d1aa, 32'h427f77b9, 32'h42b330db, 32'h41ca4e21, 32'h42a9ddec, 32'h42b2ea9f, 32'h42370743};
test_weights[23848:23855] = '{32'h42c372c7, 32'h42530f74, 32'hc260d0c2, 32'h417bf509, 32'hc0c0c8d2, 32'hc1b4f3d7, 32'hc263e85f, 32'h42c588b6};
test_bias[2981:2981] = '{32'h42c5ca31};
test_output[2981:2981] = '{32'hc6706ae6};
test_input[23856:23863] = '{32'h4247629d, 32'h42be83a9, 32'h42903d7a, 32'hc24b2c8d, 32'hc2a8c059, 32'hc1d3c3fe, 32'hc22a4f25, 32'h4130ccec};
test_weights[23856:23863] = '{32'hc0d2b0e2, 32'h4149797c, 32'h425e58e6, 32'h420c7eb9, 32'h424df257, 32'hc2c2eca7, 32'h40e730d3, 32'h4290b226};
test_bias[2982:2982] = '{32'hbfe0ac17};
test_output[2982:2982] = '{32'h44e3bd7a};
test_input[23864:23871] = '{32'hc239f810, 32'hc2628d47, 32'h426bb891, 32'hc20b6886, 32'h42559fd1, 32'h41e244f6, 32'h42a9a2e3, 32'h42b8fb93};
test_weights[23864:23871] = '{32'h424b8a6e, 32'h41857952, 32'hc2457ced, 32'h427ed075, 32'hc2c06ca8, 32'hc0a852b2, 32'h42a44f14, 32'h4236eb8f};
test_bias[2983:2983] = '{32'h428b60ff};
test_output[2983:2983] = '{32'hc519c03c};
test_input[23872:23879] = '{32'hc198d983, 32'h41a8f549, 32'hc21ef42d, 32'hc27619d1, 32'hc2b342c5, 32'hc2c21500, 32'h42a333c9, 32'h422258c7};
test_weights[23872:23879] = '{32'hc2ab602a, 32'h3f5da534, 32'h40e37436, 32'hc1b43d27, 32'h42b68940, 32'h428a235b, 32'h4281ce57, 32'h41853d15};
test_bias[2984:2984] = '{32'h42b18c6c};
test_output[2984:2984] = '{32'hc5bd7703};
test_input[23880:23887] = '{32'h41f4ae57, 32'h41cd4b6d, 32'hc20567b0, 32'hc2c25684, 32'h407a76c0, 32'hc2933566, 32'h429bbf5c, 32'hc21c9cf6};
test_weights[23880:23887] = '{32'hc10a52ec, 32'h419b9b52, 32'hc2192ab2, 32'h42b6a8b3, 32'h41acf366, 32'hc2aee9c4, 32'hc21bfa11, 32'h41770791};
test_bias[2985:2985] = '{32'h4297e384};
test_output[2985:2985] = '{32'hc589afe2};
test_input[23888:23895] = '{32'hc00d30fb, 32'h429cb467, 32'hc2b8bf9a, 32'h420a873a, 32'hc2b1de25, 32'h428bd410, 32'hbc53159d, 32'h42c5f32b};
test_weights[23888:23895] = '{32'hc2a19e9d, 32'hc185b7a7, 32'h3ffca01e, 32'hc27bf547, 32'hc275b589, 32'h42b32b9b, 32'h42ac497b, 32'h428cbf1c};
test_bias[2986:2986] = '{32'hc0c736c7};
test_output[2986:2986] = '{32'h466d53dd};
test_input[23896:23903] = '{32'h427fc377, 32'h41fc83fe, 32'hc0476f1d, 32'hc1affbf3, 32'hc1ca13b3, 32'hc28cc253, 32'h42aebbbf, 32'h41b3a497};
test_weights[23896:23903] = '{32'h42c40644, 32'h422fb4f4, 32'h4295a2e9, 32'h4212aba8, 32'hc27a8261, 32'h41e7775c, 32'hc2974673, 32'h4204706f};
test_bias[2987:2987] = '{32'hc15b4e17};
test_output[2987:2987] = '{32'h438c7b28};
test_input[23904:23911] = '{32'hc0df5b66, 32'hc2ad49d0, 32'hc2092366, 32'hc26abf53, 32'h41f5677f, 32'h41b9896d, 32'h422c34fe, 32'h42afc60e};
test_weights[23904:23911] = '{32'h40c75eaf, 32'hc2b5f0cf, 32'hc2870836, 32'hc08d285b, 32'hc155fba4, 32'h42604b5c, 32'h4202e899, 32'h420708ae};
test_bias[2988:2988] = '{32'h42967e13};
test_output[2988:2988] = '{32'h4676262a};
test_input[23912:23919] = '{32'hc23b4c5c, 32'hc2673e55, 32'h426054d2, 32'hc1e337a1, 32'hc2bb8be3, 32'h4190ae25, 32'hc2969cf1, 32'h4295d0c4};
test_weights[23912:23919] = '{32'hc247f43d, 32'hc251d998, 32'hc1f84cca, 32'hc1ca4704, 32'hc18d1be0, 32'hc1a43eef, 32'h41f3f3ae, 32'hc0c98c1c};
test_bias[2989:2989] = '{32'hc28fc015};
test_output[2989:2989] = '{32'h452e9b9d};
test_input[23920:23927] = '{32'h428aeb8a, 32'h418c6655, 32'hc237838d, 32'h42398d2c, 32'hc2c37443, 32'hc29e22fd, 32'h42c7541d, 32'h42ba281c};
test_weights[23920:23927] = '{32'hc19e878a, 32'hc2699c97, 32'hc20f6f0f, 32'hc296958f, 32'h42916b97, 32'h42050e84, 32'hc2aa006d, 32'h42a8004e};
test_bias[2990:2990] = '{32'h41b803c9};
test_output[2990:2990] = '{32'hc6645ad9};
test_input[23928:23935] = '{32'hc09fcf16, 32'hc266e764, 32'h42bc9099, 32'hc19747ed, 32'h410cde6a, 32'h42320396, 32'h41eea6f2, 32'hc2c424da};
test_weights[23928:23935] = '{32'h4294173c, 32'h428c83cf, 32'h420545c2, 32'h42c349d4, 32'hc267b331, 32'h42aca5c6, 32'h42a53b6d, 32'h42177b3c};
test_bias[2991:2991] = '{32'h42410c62};
test_output[2991:2991] = '{32'hc47a05a1};
test_input[23936:23943] = '{32'h424813e6, 32'hc1af4870, 32'hc1c2d1b2, 32'h42c33da7, 32'h423dec89, 32'hc2bd5548, 32'hc2a0906e, 32'hc2840e39};
test_weights[23936:23943] = '{32'h42a4d523, 32'hc284474f, 32'h4229f68f, 32'hc2632d47, 32'h3fd24bfb, 32'h419a7f0e, 32'hc2229ddd, 32'hc2901f8d};
test_bias[2992:2992] = '{32'hc2659a22};
test_output[2992:2992] = '{32'h45a2b663};
test_input[23944:23951] = '{32'h42c02c6d, 32'hc2933936, 32'h4143d643, 32'hc2ab0485, 32'hc2ab4dc7, 32'h4233447a, 32'h429bb66f, 32'h422ed854};
test_weights[23944:23951] = '{32'h41c358f1, 32'hc15593a1, 32'h42b69e21, 32'hc2761c9b, 32'h42573caf, 32'h422c8834, 32'h4167a313, 32'hc20dafa1};
test_bias[2993:2993] = '{32'h4244dd9a};
test_output[2993:2993] = '{32'h45d01f9a};
test_input[23952:23959] = '{32'hc2a72864, 32'hc299fd35, 32'hc283000f, 32'h4184f72e, 32'h422a97e5, 32'hc276e561, 32'hc28347f5, 32'hc2b14c52};
test_weights[23952:23959] = '{32'hc26d8bb0, 32'hc1e19671, 32'h40bb0564, 32'hc29c1286, 32'h429f105f, 32'hc244acf0, 32'h4226d07b, 32'hc275bf45};
test_bias[2994:2994] = '{32'hc08cd0ab};
test_output[2994:2994] = '{32'h4663e81b};
test_input[23960:23967] = '{32'hc22ce55c, 32'hc2286d30, 32'hc1170d52, 32'hc1a88017, 32'h4198974c, 32'h422b7eaf, 32'h427b2198, 32'h426638df};
test_weights[23960:23967] = '{32'hc2014bdc, 32'hc2c3abed, 32'h4130fb16, 32'h424eb0aa, 32'h4108cf4b, 32'hc295ec5c, 32'hc275aadd, 32'hc289d0be};
test_bias[2995:2995] = '{32'h40b0756b};
test_output[2995:2995] = '{32'hc5cc7a52};
test_input[23968:23975] = '{32'h421ef1db, 32'h40897259, 32'hc22a9c72, 32'hc28650cb, 32'hc25354b2, 32'h42385e71, 32'hc0138a6c, 32'h40fc9b4b};
test_weights[23968:23975] = '{32'h4225fa50, 32'h42996962, 32'hc289794d, 32'h42c132fa, 32'h427bfbfa, 32'hc21f002b, 32'hc28c7b18, 32'h42329d7c};
test_bias[2996:2996] = '{32'hc2b0caef};
test_output[2996:2996] = '{32'hc5c53d91};
test_input[23976:23983] = '{32'h4165c52e, 32'hc24b9208, 32'hc276ca9a, 32'h41bbf464, 32'h4113f253, 32'hc289948a, 32'h4283a2f0, 32'hc2a226ad};
test_weights[23976:23983] = '{32'h40b1ddeb, 32'hc1d78fe6, 32'hc1cd4e5f, 32'hc28ae9d5, 32'h42a35d33, 32'hc2b3c290, 32'h427acb48, 32'hc1c1a672};
test_bias[2997:2997] = '{32'h42c3e4ec};
test_output[2997:2997] = '{32'h4662fffd};
test_input[23984:23991] = '{32'hbd1acad0, 32'hc1c98452, 32'hc260dae1, 32'h428dbdc0, 32'h428321bf, 32'hc2452c44, 32'hc2c3e7d7, 32'hc1cc52a0};
test_weights[23984:23991] = '{32'hc2ad557a, 32'hc28be923, 32'hc1cbd694, 32'h4265e278, 32'h4287764f, 32'hc2908678, 32'h41b2bab5, 32'hc2a2d966};
test_bias[2998:2998] = '{32'h40bf5141};
test_output[2998:2998] = '{32'h466d0b7d};
test_input[23992:23999] = '{32'h42b42455, 32'hc2a617c6, 32'hc10451b1, 32'h4242d20d, 32'hc0d1a0d7, 32'hc2909b2d, 32'hc2316ca6, 32'hc1bba77f};
test_weights[23992:23999] = '{32'h42123fc0, 32'h42bc5f50, 32'h41ed8cdf, 32'hc089a1ef, 32'h42b3e72e, 32'hc1e845c4, 32'hc205fec0, 32'h40959d11};
test_bias[2999:2999] = '{32'h41e0a353};
test_output[2999:2999] = '{32'hc5015667};
test_input[24000:24007] = '{32'h414b80ec, 32'hc2b82d64, 32'h405c2eb8, 32'hc2646491, 32'h42248f68, 32'hc1d3897f, 32'h4213deee, 32'hc12d35a9};
test_weights[24000:24007] = '{32'hc237eeee, 32'h4266155b, 32'h42aeeff9, 32'h41dfa104, 32'hc28149e9, 32'hc1b6cf4b, 32'h408c6cf3, 32'h41966438};
test_bias[3000:3000] = '{32'h425f891c};
test_output[3000:3000] = '{32'hc61006c8};
test_input[24008:24015] = '{32'hc096d6cb, 32'hc14eaa64, 32'h41a30d3a, 32'hc272bb26, 32'hc2ace11c, 32'h423a9c12, 32'hc1d7936b, 32'h4240318f};
test_weights[24008:24015] = '{32'hc1a05a3e, 32'h40f90d5b, 32'hc2305708, 32'hc24db398, 32'h4270e85e, 32'h4220bb08, 32'hc2a439e7, 32'h4271c255};
test_bias[3001:3001] = '{32'h423109f9};
test_output[3001:3001] = '{32'h457cdb03};
test_input[24016:24023] = '{32'hc23e97ab, 32'h4203fabb, 32'h42a92391, 32'h42aadf54, 32'h42ba03a7, 32'hc2b2378e, 32'hc024fdd3, 32'h4269bb50};
test_weights[24016:24023] = '{32'hc0f25715, 32'hc24e108a, 32'hc1c8e520, 32'h41d7ddf7, 32'hc260a019, 32'h41f3af5e, 32'hc2a05efa, 32'hc1a6a03f};
test_bias[3002:3002] = '{32'hc2924572};
test_output[3002:3002] = '{32'hc61f07ea};
test_input[24024:24031] = '{32'hc2a9c4c1, 32'h42086449, 32'h42c0dfea, 32'hc2b5cf4e, 32'hc287dd28, 32'h420947f6, 32'hc280ce09, 32'h42664567};
test_weights[24024:24031] = '{32'h411661f7, 32'hc1e1786f, 32'h411a37f3, 32'hc291cdac, 32'h4202dc83, 32'hc2580d85, 32'hc20d65a0, 32'h4292aace};
test_bias[3003:3003] = '{32'hc2b4bebe};
test_output[3003:3003] = '{32'h45fe0c14};
test_input[24032:24039] = '{32'hc2915cdb, 32'hc2441b2e, 32'h428467c4, 32'h42790ac0, 32'hc270ef40, 32'h424fda06, 32'hc28b11ce, 32'hc1929a67};
test_weights[24032:24039] = '{32'h4244f219, 32'hc2885305, 32'hc2a09a5f, 32'hbf526dd0, 32'h405ecb90, 32'h4157f616, 32'hc2bf7727, 32'hc17c71db};
test_bias[3004:3004] = '{32'hc014e2f7};
test_output[3004:3004] = '{32'h44e4e2ad};
test_input[24040:24047] = '{32'hc2a4494b, 32'hc24810c0, 32'h42859e14, 32'hc1166fec, 32'h412a1a5a, 32'hc241cf0a, 32'hc29a5813, 32'hc20b7183};
test_weights[24040:24047] = '{32'hc29fa766, 32'hc0ca8bdd, 32'h424f9170, 32'hc2980733, 32'hc224fc6e, 32'h422d1d20, 32'hc288579d, 32'hc23f4fa8};
test_bias[3005:3005] = '{32'hc281b5b1};
test_output[3005:3005] = '{32'h46705d29};
test_input[24048:24055] = '{32'h3fadafde, 32'hc19a2910, 32'hc21a65ed, 32'h426e0eb0, 32'h41bcaa8c, 32'hc1e17170, 32'h3ebaa8de, 32'h422ab090};
test_weights[24048:24055] = '{32'hc22182ef, 32'hc234a915, 32'h42630c3d, 32'h41555775, 32'hc14ae298, 32'hc1a887e4, 32'h41bc7262, 32'h41e164ae};
test_bias[3006:3006] = '{32'hc205cbe1};
test_output[3006:3006] = '{32'h445e8828};
test_input[24056:24063] = '{32'hc297f016, 32'h41e73d59, 32'hc13ebdb8, 32'h427da13a, 32'h421947a3, 32'hc2b13804, 32'h418b331e, 32'hc2b46d43};
test_weights[24056:24063] = '{32'hc25807a6, 32'hc2419fb7, 32'hc241ec34, 32'h428be51d, 32'hc29ce5d1, 32'h42469a7e, 32'hc297d001, 32'h4205d8ba};
test_bias[3007:3007] = '{32'hc2c389fa};
test_output[3007:3007] = '{32'hc580f06f};
test_input[24064:24071] = '{32'hc2b43069, 32'hc2891f22, 32'h42a5e869, 32'hc2c66195, 32'hc2b77105, 32'h3ec59852, 32'hc114deae, 32'h42a64318};
test_weights[24064:24071] = '{32'h4260a51a, 32'h42068804, 32'h423104af, 32'hc1a0478e, 32'h429a8450, 32'hc29954e2, 32'h41a31594, 32'h413d20c3};
test_bias[3008:3008] = '{32'h42bba442};
test_output[3008:3008] = '{32'hc5f802b3};
test_input[24072:24079] = '{32'h40e62e14, 32'h4289f461, 32'hc29524a6, 32'h429741b8, 32'h4235f342, 32'hc28c44b3, 32'h42511b25, 32'hc2a26c4f};
test_weights[24072:24079] = '{32'h4297e48a, 32'hc2608ed9, 32'h4234dcd0, 32'hc1a6c4ce, 32'hc2b88a75, 32'h41ac41ff, 32'h427313f3, 32'hc1991d81};
test_bias[3009:3009] = '{32'hc28a24f6};
test_output[3009:3009] = '{32'hc6119e88};
test_input[24080:24087] = '{32'hc2ada15d, 32'hc21a6662, 32'hc2c64a89, 32'h3f99e280, 32'h4295987c, 32'h41a1b112, 32'hc0418e1d, 32'hc11fa5cd};
test_weights[24080:24087] = '{32'h42a21a8d, 32'h42510062, 32'h42c124e7, 32'hbf066328, 32'h40d81a2b, 32'hc282f0eb, 32'h3e52933e, 32'h424735f0};
test_bias[3010:3010] = '{32'h42115970};
test_output[3010:3010] = '{32'hc69b8821};
test_input[24088:24095] = '{32'h428d2f9a, 32'hc29a8b37, 32'h4210b99b, 32'hc2543982, 32'h42c1cd52, 32'h42499fad, 32'h425bad56, 32'h41fc6c85};
test_weights[24088:24095] = '{32'hc29efe45, 32'hc2bf34b2, 32'h422bef94, 32'hc1ca8b40, 32'h425e2789, 32'hc20048e0, 32'hc28059c2, 32'hc264559b};
test_bias[3011:3011] = '{32'h42a4ceed};
test_output[3011:3011] = '{32'h4547bf63};
test_input[24096:24103] = '{32'hc2a82fdd, 32'hc2778240, 32'h410de7b6, 32'hc2a49f22, 32'hc2c77014, 32'h422ac7dc, 32'hc254fae5, 32'h42909f47};
test_weights[24096:24103] = '{32'h422893ba, 32'hc292cf8b, 32'hc26f9341, 32'h40a7df35, 32'h42af5d0d, 32'hc11f3b77, 32'hc1f46469, 32'hc246c8d4};
test_bias[3012:3012] = '{32'hc1962bc8};
test_output[3012:3012] = '{32'hc62dbc92};
test_input[24104:24111] = '{32'h42afad33, 32'h4250364a, 32'h421eec28, 32'hc23a5a41, 32'hc1459b0e, 32'hc29186ac, 32'h3f5f09b2, 32'hc270fab6};
test_weights[24104:24111] = '{32'h426657e2, 32'h4040ce28, 32'h42341127, 32'h40335f9a, 32'hc2820af4, 32'h4269c48d, 32'hc10da161, 32'h422e44db};
test_bias[3013:3013] = '{32'hc289a423};
test_output[3013:3013] = '{32'h44349a8c};
test_input[24112:24119] = '{32'hc1c2ae99, 32'hc18515a9, 32'hc28ff5fa, 32'h41e6ba63, 32'h42806f89, 32'h41f59fb0, 32'h4287f3bc, 32'hc2ae6df2};
test_weights[24112:24119] = '{32'hc18ddc6f, 32'h42136d32, 32'h42909471, 32'h40d78238, 32'h41dc1865, 32'h429bcc39, 32'hc2a3160b, 32'hc0146190};
test_bias[3014:3014] = '{32'h429b1d08};
test_output[3014:3014] = '{32'hc5c4bc7b};
test_input[24120:24127] = '{32'hc286a826, 32'hc1e71d59, 32'hc2bba87c, 32'h413945cb, 32'hbf705a1b, 32'hc2274a38, 32'h4166dd43, 32'hc20a9b33};
test_weights[24120:24127] = '{32'h4244d5d3, 32'h427746e4, 32'hc0f5a613, 32'h4228e08d, 32'h42105beb, 32'h4241823e, 32'hc2442bea, 32'hc2675ad9};
test_bias[3015:3015] = '{32'hc2a43ece};
test_output[3015:3015] = '{32'hc593e4d8};
test_input[24128:24135] = '{32'hc0bc8a5c, 32'hc2b26eba, 32'hc2c52475, 32'hc27bfbd9, 32'h4227e587, 32'hc2a354b2, 32'hc21ef99d, 32'hc02c4d25};
test_weights[24128:24135] = '{32'hc26b8c8e, 32'h4192cbf3, 32'h42a45f98, 32'hc2c6605c, 32'hc23b548c, 32'h42666979, 32'hc1695e4a, 32'hc23370d9};
test_bias[3016:3016] = '{32'h41e6caf1};
test_output[3016:3016] = '{32'hc60dee26};
test_input[24136:24143] = '{32'hc2c44707, 32'h42724ae8, 32'h40c6f41e, 32'h40473db8, 32'h41c816e5, 32'hc2c09967, 32'h429379a6, 32'h4209985e};
test_weights[24136:24143] = '{32'hc2b4868a, 32'h4271a20b, 32'h42bec609, 32'hc2b4043f, 32'h42931d92, 32'hc21b6469, 32'h42777828, 32'h42a37371};
test_bias[3017:3017] = '{32'hc2c6d942};
test_output[3017:3017] = '{32'h46c8a9aa};
test_input[24144:24151] = '{32'hc20ccd1a, 32'h4218bd98, 32'h42c4e050, 32'h3d566da0, 32'hc2a1078d, 32'hc25330f4, 32'h41a3fef5, 32'h42b2ab41};
test_weights[24144:24151] = '{32'h41de5d7a, 32'h41300a78, 32'h41454b49, 32'hc202acec, 32'h42461bc7, 32'hc1ae2e17, 32'hbfe072e0, 32'hc28fbf27};
test_bias[3018:3018] = '{32'hc09c6309};
test_output[3018:3018] = '{32'hc607178c};
test_input[24152:24159] = '{32'h42923c6f, 32'h425e490a, 32'h426b444b, 32'hc199a041, 32'hc09013c7, 32'hc1fb143c, 32'h42814595, 32'h42a3afa3};
test_weights[24152:24159] = '{32'hc25e5551, 32'hc10a072e, 32'h42786a69, 32'hc1ecb496, 32'hc0a91df5, 32'h411e4f32, 32'hc281b49b, 32'h410d391d};
test_bias[3019:3019] = '{32'hc19cff75};
test_output[3019:3019] = '{32'hc5801338};
test_input[24160:24167] = '{32'h42446157, 32'h41f7f442, 32'hc2a1987e, 32'hc106db08, 32'h427a52a1, 32'hc2518b28, 32'hc2b21574, 32'h429f6595};
test_weights[24160:24167] = '{32'hc1f331bf, 32'hc1496d1d, 32'h42765374, 32'hc2073309, 32'h41cab05c, 32'h428235b9, 32'h42977be8, 32'hc1926528};
test_bias[3020:3020] = '{32'h423ba716};
test_output[3020:3020] = '{32'hc681545a};
test_input[24168:24175] = '{32'hc13e03a8, 32'h420f8700, 32'hc1aa892e, 32'hc293c2c2, 32'h428b07ca, 32'h42894fa6, 32'h41db0346, 32'h419ffd7d};
test_weights[24168:24175] = '{32'h41d79760, 32'h42976bd4, 32'h429720ed, 32'hc26902c0, 32'hc17477da, 32'h4244e472, 32'h42afca6d, 32'hc292c51f};
test_bias[3021:3021] = '{32'h4193c803};
test_output[3021:3021] = '{32'h4602afd4};
test_input[24176:24183] = '{32'h4213ee4e, 32'h428c32ba, 32'h42a5525b, 32'hc28ad458, 32'hc2ba40d8, 32'h42aeb402, 32'hc2b96a17, 32'hc20b3a2e};
test_weights[24176:24183] = '{32'hc22f56f8, 32'hc27986cc, 32'h42a67e03, 32'h4107de33, 32'hc2612c32, 32'hc256463e, 32'h4265e934, 32'hc095a973};
test_bias[3022:3022] = '{32'h42b4d69f};
test_output[3022:3022] = '{32'hc583b4b5};
test_input[24184:24191] = '{32'h41da2027, 32'hc0841334, 32'h40c887f0, 32'hc1a7d0f6, 32'hc24e4314, 32'hc2c04fe3, 32'h419879bc, 32'h420801b6};
test_weights[24184:24191] = '{32'hc1d26037, 32'h41e074fd, 32'hc2a9c8d0, 32'hc27c594e, 32'h41eda48b, 32'hc2b0617d, 32'h41f355bb, 32'hc285e248};
test_bias[3023:3023] = '{32'h423543af};
test_output[3023:3023] = '{32'h45a43e1f};
test_input[24192:24199] = '{32'hc22bc694, 32'h42937c13, 32'h4260f6c7, 32'h42585d64, 32'hc0ca0faf, 32'hc1b815a5, 32'hc2bd8786, 32'h4295d4b1};
test_weights[24192:24199] = '{32'hc28c169a, 32'hc29197b8, 32'h3e582f75, 32'hc2583f23, 32'hc2b48285, 32'h41f52f2d, 32'h42b65b92, 32'h4262a2ce};
test_bias[3024:3024] = '{32'h42a9b133};
test_output[3024:3024] = '{32'hc617dbde};
test_input[24200:24207] = '{32'hbf88cad7, 32'hc2856a67, 32'h4255ee67, 32'h42472ea0, 32'hc0fafe65, 32'hc0b7b2f5, 32'hc280c6af, 32'h41f32c81};
test_weights[24200:24207] = '{32'hc2c16e56, 32'hc1d9e365, 32'h423d614d, 32'hc2359bde, 32'hc281dcbe, 32'hc29e2119, 32'hc2bbe60e, 32'h4238a9dc};
test_bias[3025:3025] = '{32'h413a1704};
test_output[3025:3025] = '{32'h4625eb5a};
test_input[24208:24215] = '{32'h4262bf52, 32'hbf2597bc, 32'hc21b8459, 32'hc2288816, 32'hc1533848, 32'h42b7e5fc, 32'hc2bdec0f, 32'hc1ed1ea9};
test_weights[24208:24215] = '{32'h427da715, 32'hc23daee2, 32'hc29edc6c, 32'h424923c2, 32'hc2c6df78, 32'hc1ea9812, 32'h408650c4, 32'hc1888e84};
test_bias[3026:3026] = '{32'h42790686};
test_output[3026:3026] = '{32'h45534df0};
test_input[24216:24223] = '{32'hc289deae, 32'h42866e8a, 32'hc26a3689, 32'h41acac30, 32'h42ac3df5, 32'h4270f747, 32'hc26ad010, 32'hc267b76c};
test_weights[24216:24223] = '{32'hc2c5837c, 32'hc1f21d82, 32'h429b9ab2, 32'h429e2aab, 32'h40eaa824, 32'hc261b3c8, 32'hc24326d8, 32'h41d863d5};
test_bias[3027:3027] = '{32'h41b5adb4};
test_output[3027:3027] = '{32'h43ee8b80};
test_input[24224:24231] = '{32'h42128d5d, 32'h4217e295, 32'h42b725e5, 32'hc28b8bb5, 32'hc170d68a, 32'h41a03df1, 32'hc2aa3167, 32'h4281897e};
test_weights[24224:24231] = '{32'h41f13834, 32'h41d8ff66, 32'hc2b5ac3c, 32'hc1c72183, 32'h4227334c, 32'hbf26a236, 32'h42a3b275, 32'h42a13556};
test_bias[3028:3028] = '{32'hc11131f8};
test_output[3028:3028] = '{32'hc5d5d44f};
test_input[24232:24239] = '{32'hc1434531, 32'h41b49a5d, 32'h42c145b8, 32'hc2afad9e, 32'hc1ec2ba9, 32'hc253f795, 32'hc2ba36f4, 32'hc2819e47};
test_weights[24232:24239] = '{32'h40a454e8, 32'hc194dcd5, 32'h427b9d1e, 32'hc181ba10, 32'hc2ae2c58, 32'hc1c47116, 32'h4274fb98, 32'h4106b95d};
test_bias[3029:3029] = '{32'h4294a5f3};
test_output[3029:3029] = '{32'h459375a8};
test_input[24240:24247] = '{32'h41d11bd6, 32'hc212419c, 32'hc06fab44, 32'hc21f43f7, 32'hc29af5b0, 32'h42624c8b, 32'h42351a8e, 32'h429e7348};
test_weights[24240:24247] = '{32'h41a4195f, 32'hc21bcd66, 32'hc109cae6, 32'hc0d7e5c5, 32'h4125f898, 32'h425cb61a, 32'h42a09cd3, 32'hc29d5cde};
test_bias[3030:3030] = '{32'h41116703};
test_output[3030:3030] = '{32'h44f8d5e8};
test_input[24248:24255] = '{32'h3fa47973, 32'h42b4a67c, 32'h3ff04f52, 32'hc2593e18, 32'h40818c90, 32'h422fdee0, 32'hc1e812d2, 32'h4126976e};
test_weights[24248:24255] = '{32'hc1af67fe, 32'hc1048a7d, 32'hc2c4bda7, 32'h4285f631, 32'h4120e584, 32'hc244510b, 32'h4263fcfe, 32'h42bafacc};
test_bias[3031:3031] = '{32'hc1804055};
test_output[3031:3031] = '{32'hc5e7a0d8};
test_input[24256:24263] = '{32'hc05d5a85, 32'hc2c60e90, 32'hc28ef6d3, 32'hc29dbb04, 32'hc29e710f, 32'h426bcd84, 32'hc16327d6, 32'h429df7d7};
test_weights[24256:24263] = '{32'h424592ba, 32'h4291866e, 32'h421b1630, 32'h420450bc, 32'h426db034, 32'h424d54a8, 32'h42b4fd0f, 32'h4298c749};
test_bias[3032:3032] = '{32'hc230b0d4};
test_output[3032:3032] = '{32'hc61815b3};
test_input[24264:24271] = '{32'h42863069, 32'hc284e898, 32'h42332503, 32'h425963ef, 32'hc2ae8474, 32'hc0ba955d, 32'hc22d83d5, 32'hbed5c36d};
test_weights[24264:24271] = '{32'hc124d0b1, 32'h425b2f4b, 32'h421c3967, 32'h4283a455, 32'h429c7217, 32'hc2ac476f, 32'hc1c70c65, 32'h42b7c700};
test_bias[3033:3033] = '{32'hc1f79e50};
test_output[3033:3033] = '{32'hc586fc92};
test_input[24272:24279] = '{32'h42af83be, 32'h413008c4, 32'h428c538e, 32'h42bfe442, 32'h428bc3f2, 32'h42b9bf47, 32'hc1a9d222, 32'hc2649886};
test_weights[24272:24279] = '{32'h4210a326, 32'h4278f751, 32'hc16eb783, 32'h428b1612, 32'hbf8112f0, 32'hc2864e6d, 32'h42800f69, 32'h4298088d};
test_bias[3034:3034] = '{32'hc1d815c7};
test_output[3034:3034] = '{32'hc51fa220};
test_input[24280:24287] = '{32'hc2397d79, 32'h421c6340, 32'h42a709d3, 32'h42147c0d, 32'hc2b8ebb3, 32'hc2946caa, 32'h420b0a65, 32'hc2788f16};
test_weights[24280:24287] = '{32'hc274929d, 32'h428e7d8c, 32'hc285f414, 32'hc2194cda, 32'h427c1100, 32'hc2945cca, 32'h42123579, 32'h41da8d7b};
test_bias[3035:3035] = '{32'hc2268981};
test_output[3035:3035] = '{32'hc5089bc3};
test_input[24288:24295] = '{32'hc2a8e60e, 32'h425947ad, 32'h4296104d, 32'hc2af5e13, 32'hc24270e3, 32'hc272f19c, 32'h41a9c116, 32'hc29cafa2};
test_weights[24288:24295] = '{32'hc234a4fd, 32'h425e4c32, 32'hc23cc4ee, 32'hc283db28, 32'h42a70628, 32'hc2ad7563, 32'h42bf1a24, 32'h42adecdb};
test_bias[3036:3036] = '{32'h413c3a98};
test_output[3036:3036] = '{32'h45ac1781};
test_input[24296:24303] = '{32'h4257946f, 32'h42a82b8d, 32'hc29f951f, 32'hc21ccc6b, 32'hc1e0a530, 32'hc2799ac2, 32'h40842f1a, 32'hc244d72e};
test_weights[24296:24303] = '{32'hc2469d00, 32'hc183b89a, 32'hc1a6f1b0, 32'h42b7eda9, 32'hc2c798c8, 32'hc2237b84, 32'hc231947f, 32'hc299706a};
test_bias[3037:3037] = '{32'hc265c584};
test_output[3037:3037] = '{32'h45346eaf};
test_input[24304:24311] = '{32'h423ecc55, 32'hc1cd648a, 32'hc2609cd7, 32'h42416c4a, 32'hc1c461c0, 32'hc2ba7bbd, 32'h41a4543c, 32'h413c363c};
test_weights[24304:24311] = '{32'h420d257f, 32'h429c487e, 32'h4222214a, 32'hc2b666c9, 32'hc166e5b4, 32'hc1ffbf05, 32'h40b64da3, 32'h428124fd};
test_bias[3038:3038] = '{32'h4220b471};
test_output[3038:3038] = '{32'hc52c55d8};
test_input[24312:24319] = '{32'h42c26bb6, 32'h4260ead9, 32'hc27f9ed6, 32'h42ba566e, 32'hc297a31f, 32'h41499f74, 32'hc2685b03, 32'hc2c43b82};
test_weights[24312:24319] = '{32'h3ec80adc, 32'h40e1b0d9, 32'h42aff52a, 32'h426d8f82, 32'h42a75d17, 32'h42b6125a, 32'h40b9c1b7, 32'h40c12506};
test_bias[3039:3039] = '{32'h4222e117};
test_output[3039:3039] = '{32'hc5b36499};
test_input[24320:24327] = '{32'hc2551515, 32'h42bcb625, 32'hc2bc0478, 32'h4296e3eb, 32'h4231dd06, 32'hc0eaa7b1, 32'hc18edc5b, 32'hc294140b};
test_weights[24320:24327] = '{32'hc24cb5cd, 32'h42990ee0, 32'h4281c7fc, 32'hc249f392, 32'h425e929a, 32'hc2938660, 32'h42922eb3, 32'hc22a5e09};
test_bias[3040:3040] = '{32'hc0595e76};
test_output[3040:3040] = '{32'h45990e8c};
test_input[24328:24335] = '{32'h4263fef7, 32'h428384a3, 32'hc25af664, 32'hc2b174cd, 32'h429faf3f, 32'h4047bd71, 32'h429e3309, 32'hc2a18032};
test_weights[24328:24335] = '{32'h42469f4b, 32'h40af90a7, 32'hc2be7745, 32'h4204893b, 32'hc12e704f, 32'h42a59238, 32'h4218bc55, 32'h42bc5169};
test_bias[3041:3041] = '{32'h41dba49a};
test_output[3041:3041] = '{32'h43944ca2};
test_input[24336:24343] = '{32'h411dbc18, 32'hc1fb2d3a, 32'hc03eb128, 32'hc2baf364, 32'hc187487c, 32'h423664c5, 32'hc26b7480, 32'h42b4ddf0};
test_weights[24336:24343] = '{32'hc226610a, 32'hc254895b, 32'h4291fd83, 32'hc24e816c, 32'hc2a0e321, 32'hc2c7d205, 32'h41b27091, 32'hc2c205a4};
test_bias[3042:3042] = '{32'h41d0f478};
test_output[3042:3042] = '{32'hc5e6e652};
test_input[24344:24351] = '{32'hc1e5b1c2, 32'hc2a701cc, 32'h422e8b42, 32'h42a680e3, 32'h42c1a1a3, 32'h41827099, 32'hc281880d, 32'h4170ed6a};
test_weights[24344:24351] = '{32'h42bb34ea, 32'hc2b57930, 32'h42c7be79, 32'hc210f701, 32'h4298e93d, 32'hc2277d8c, 32'h427b6574, 32'hc23396ce};
test_bias[3043:3043] = '{32'h41995e6e};
test_output[3043:3043] = '{32'h460078c3};
test_input[24352:24359] = '{32'h42619137, 32'hc2a5a23f, 32'hbee36641, 32'h4287cd3e, 32'hc26445fd, 32'hc05438fc, 32'hc18f3f4d, 32'hc137c15d};
test_weights[24352:24359] = '{32'h42c7572e, 32'h42578cf7, 32'h42685d1e, 32'hc1e95ae4, 32'h42865faf, 32'h429bd186, 32'h3f07254e, 32'hc2139c5f};
test_bias[3044:3044] = '{32'h41390bf1};
test_output[3044:3044] = '{32'hc58d1a77};
test_input[24360:24367] = '{32'h42a628c6, 32'h4234185d, 32'h42c440db, 32'h424c8a1f, 32'h4249163c, 32'h429445e9, 32'h42b469f9, 32'h4267bb2f};
test_weights[24360:24367] = '{32'h427c6ef2, 32'hc130afec, 32'h42af2d81, 32'hc1aeff63, 32'h4278c830, 32'h4205cb79, 32'hc01bd578, 32'hc276d3a8};
test_bias[3045:3045] = '{32'hc2b5a200};
test_output[3045:3045] = '{32'h4659dcd7};
test_input[24368:24375] = '{32'h4157de12, 32'hc2954f11, 32'h421d1dda, 32'hc29db0a6, 32'hc2638057, 32'h42702edb, 32'hc29cedbf, 32'hc232b88e};
test_weights[24368:24375] = '{32'hc2131598, 32'h42156a27, 32'h4045025f, 32'h416d5245, 32'hc21d2a13, 32'hc219a24e, 32'h4283c8c0, 32'hc273367d};
test_bias[3046:3046] = '{32'hc28c7bdb};
test_output[3046:3046] = '{32'hc5d884a2};
test_input[24376:24383] = '{32'hc2bf1ab7, 32'h426eb19f, 32'hc29074cf, 32'h417bbc3f, 32'h42a4cdc5, 32'hc1b1e509, 32'h419c5568, 32'h4112e724};
test_weights[24376:24383] = '{32'hc2b8240a, 32'h42187f6d, 32'h422c7be6, 32'h423406a1, 32'h42719380, 32'h41cdd89b, 32'hc2840817, 32'hc2ad32fa};
test_bias[3047:3047] = '{32'hc201776e};
test_output[3047:3047] = '{32'h462b23e9};
test_input[24384:24391] = '{32'hc1621db6, 32'h42a5d5bb, 32'h426e745a, 32'h423308fc, 32'hc1e18870, 32'hc2c4627d, 32'h42c6f33d, 32'hc2b8d319};
test_weights[24384:24391] = '{32'hc24d87eb, 32'h41c0b5ac, 32'h4228eddd, 32'h41d7b4a5, 32'h425dcc23, 32'h42990b8a, 32'h412e21b9, 32'hc28376f0};
test_bias[3048:3048] = '{32'h41e0796d};
test_output[3048:3048] = '{32'h458e5ff5};
test_input[24392:24399] = '{32'hc108146f, 32'h413392b0, 32'h428997a1, 32'hc2575b85, 32'hc29e3549, 32'h41ec2e3e, 32'hc22e7b9d, 32'h420983cc};
test_weights[24392:24399] = '{32'hc23c97ed, 32'h4280d678, 32'h423121e1, 32'h423ec2bf, 32'h42badd83, 32'h415a434b, 32'h41c5ce2e, 32'h418e1ddd};
test_bias[3049:3049] = '{32'hc223d216};
test_output[3049:3049] = '{32'hc5b8308f};
test_input[24400:24407] = '{32'h4292ce08, 32'h42b128d0, 32'hc272f9bc, 32'hc14f51a5, 32'hc07be280, 32'hc1529dea, 32'h42701c76, 32'hc2ac784d};
test_weights[24400:24407] = '{32'h420cd0f4, 32'h42776c5b, 32'h4108d1e0, 32'hc2814a02, 32'h425b80ad, 32'h41295e57, 32'hc1e8e2d3, 32'h420eab46};
test_bias[3050:3050] = '{32'hc114750c};
test_output[3050:3050] = '{32'h454799c2};
test_input[24408:24415] = '{32'h423a8542, 32'h3e6300b7, 32'hc115f207, 32'h42bd265d, 32'h41d44952, 32'hc1db455a, 32'h3e6a0509, 32'h4246b2c9};
test_weights[24408:24415] = '{32'h418cce6e, 32'hc115c333, 32'h42853758, 32'h42537e83, 32'hc1cfcbe1, 32'hc1ee27ad, 32'h42807956, 32'hc20371ea};
test_bias[3051:3051] = '{32'h4192f9a7};
test_output[3051:3051] = '{32'h4568a503};
test_input[24416:24423] = '{32'hc2af82c9, 32'h4244e0d7, 32'h42a8265c, 32'h42174ca5, 32'h413450f3, 32'h42238408, 32'hc2a885e8, 32'hc1fb6a00};
test_weights[24416:24423] = '{32'hc1ac77d0, 32'hc2520b1c, 32'h425d245c, 32'hc1a8c2ed, 32'hc2a2a6a8, 32'hc28eeaf0, 32'h42b464fb, 32'h41812265};
test_bias[3052:3052] = '{32'hc2801fa0};
test_output[3052:3052] = '{32'hc60a4eab};
test_input[24424:24431] = '{32'hc2a04360, 32'h42b20f86, 32'hc23f84d1, 32'h42665f44, 32'hc1f0f089, 32'h42b59d1f, 32'h420dc235, 32'hc1c2e205};
test_weights[24424:24431] = '{32'h415c2085, 32'h42c45e58, 32'hc1259a2b, 32'hc22b5184, 32'hc2b7b25f, 32'h427c9186, 32'hc25bb342, 32'hc25a045c};
test_bias[3053:3053] = '{32'hc2b2bc27};
test_output[3053:3053] = '{32'h46524e89};
test_input[24432:24439] = '{32'h42554745, 32'h42739310, 32'h4224c7da, 32'hc2610635, 32'hc2baab0c, 32'h424832b0, 32'h429866b0, 32'hc2c7bc66};
test_weights[24432:24439] = '{32'hc1fc8ef9, 32'hc2056ed6, 32'h42c58818, 32'hc1cae216, 32'hc0ebf0a2, 32'h420912a6, 32'hc1277dca, 32'h41fc2a42};
test_bias[3054:3054] = '{32'h4299e97a};
test_output[3054:3054] = '{32'h439db2f9};
test_input[24440:24447] = '{32'h424b7ae8, 32'h41ee19ac, 32'h418579f5, 32'h42510414, 32'hc24b1767, 32'h41d61cc1, 32'h42ab59f2, 32'hc20a5968};
test_weights[24440:24447] = '{32'hc29698cc, 32'h411e083a, 32'h41ef8786, 32'hc29e34c0, 32'hc05d8b75, 32'h42bcd48c, 32'h413fec36, 32'hc2479d94};
test_bias[3055:3055] = '{32'h42afeb87};
test_output[3055:3055] = '{32'hc4cb3f50};
test_input[24448:24455] = '{32'hc2755666, 32'hc29bebc5, 32'hc190a324, 32'hc20c2162, 32'h42bcae24, 32'h4191557a, 32'h42c77ecb, 32'h428d806f};
test_weights[24448:24455] = '{32'hc29ab7cc, 32'hc180bb91, 32'h424adeb2, 32'h3fe3c1e1, 32'hc2aea53a, 32'h41bf59d0, 32'hc027d91e, 32'h4210cf36};
test_bias[3056:3056] = '{32'h42a95d15};
test_output[3056:3056] = '{32'hc3c78c70};
test_input[24456:24463] = '{32'h41bf6af1, 32'hc1b810c7, 32'hc2c25a93, 32'hc2bfeb4e, 32'h418fdbb6, 32'hc22c2317, 32'hc234770f, 32'h3f295dd1};
test_weights[24456:24463] = '{32'h429cdb29, 32'hc2807456, 32'h41a9ef75, 32'h411daf8b, 32'h42612729, 32'hc0a458fa, 32'hc27efe81, 32'h41889655};
test_bias[3057:3057] = '{32'h41c59217};
test_output[3057:3057] = '{32'h458c4d64};
test_input[24464:24471] = '{32'hc29d1683, 32'hc0d4d25a, 32'hc2b77906, 32'h4258aa98, 32'hc2b27257, 32'h41b81b1f, 32'h41d91910, 32'hc181069d};
test_weights[24464:24471] = '{32'hc1af2284, 32'h42bfbfb7, 32'hc24f4871, 32'h40e2d79d, 32'hc174da9c, 32'h42a373c0, 32'h3f561f97, 32'hc2a0b266};
test_bias[3058:3058] = '{32'h42c054c0};
test_output[3058:3058] = '{32'h462a026f};
test_input[24472:24479] = '{32'h4298f457, 32'hc24213e9, 32'h42139c2d, 32'h420e0582, 32'h41ae97c5, 32'hc294e482, 32'h422ca6a8, 32'hc1ccee39};
test_weights[24472:24479] = '{32'h42806451, 32'hc2a2bfa5, 32'hc295cb0a, 32'h41e0001f, 32'hc2c0d88d, 32'hc2980988, 32'hc2820bab, 32'hc117b5c6};
test_bias[3059:3059] = '{32'hc2924a6c};
test_output[3059:3059] = '{32'h45fa3180};
test_input[24480:24487] = '{32'h41c6d2b7, 32'h429949da, 32'hc1aed25f, 32'h41d9fdd2, 32'hc201ac39, 32'h418f3f4a, 32'hc20a24a0, 32'h4245d2bf};
test_weights[24480:24487] = '{32'hc15ec815, 32'h3d5ec050, 32'h4288b5a4, 32'h427f1ffd, 32'hc24e1a00, 32'h42768e48, 32'h4215adc3, 32'h4133dd7f};
test_bias[3060:3060] = '{32'hbe4c01b5};
test_output[3060:3060] = '{32'h44f27b78};
test_input[24488:24495] = '{32'hc0cfea60, 32'hc29cc69b, 32'hc2099ad9, 32'hc1d1f2e4, 32'hc2989b2e, 32'h421be76c, 32'h42b1b575, 32'h42a622e9};
test_weights[24488:24495] = '{32'h4120347b, 32'hc21f4d6f, 32'h42907482, 32'hc2910c35, 32'h429bf614, 32'h4244bd40, 32'hc296f109, 32'hc28077ea};
test_bias[3061:3061] = '{32'h42a737eb};
test_output[3061:3061] = '{32'hc6532f94};
test_input[24496:24503] = '{32'hc29163f6, 32'h4231fe68, 32'hc28202b4, 32'hc2b69436, 32'hc251447a, 32'h410a7a4a, 32'h419744c5, 32'hc2790a67};
test_weights[24496:24503] = '{32'hc2c4ecc2, 32'hc27abccb, 32'h42721362, 32'h42ae993d, 32'hc2a12f1f, 32'h41c1dee0, 32'h4275e99f, 32'h414993b0};
test_bias[3062:3062] = '{32'hc29d7009};
test_output[3062:3062] = '{32'hc52f9be9};
test_input[24504:24511] = '{32'hc2820cfc, 32'h40e86baf, 32'hc1b6efab, 32'hc28369fe, 32'hc1557aa2, 32'hc0a5ceee, 32'h422b94bf, 32'h4278479a};
test_weights[24504:24511] = '{32'hc21ae613, 32'hc03be7f6, 32'h42b6ab28, 32'hc28cca1a, 32'hc076538b, 32'hc2c638da, 32'h42485c41, 32'hc2032dcf};
test_bias[3063:3063] = '{32'hc299f788};
test_output[3063:3063] = '{32'h45b014f7};
test_input[24512:24519] = '{32'h4128bf66, 32'hc298629b, 32'hc20d20cd, 32'h41cb5fee, 32'h42740ac0, 32'h4272d17b, 32'hc2b466c8, 32'hc1ff9cde};
test_weights[24512:24519] = '{32'hc2c59db4, 32'h41d269f2, 32'h4210fc15, 32'h42a20099, 32'hc205bb0e, 32'h42848553, 32'hc23fdfe9, 32'hc194e276};
test_bias[3064:3064] = '{32'h424c65ce};
test_output[3064:3064] = '{32'h45928afc};
test_input[24520:24527] = '{32'h42828601, 32'hc12c583a, 32'h42988d9b, 32'hc2b6d49e, 32'h4160a56d, 32'hc2743ce9, 32'h409dc11f, 32'h429b2190};
test_weights[24520:24527] = '{32'hc2a4b0c2, 32'h40f5495d, 32'h42c4fb4e, 32'h41aae2ea, 32'hc1d9f896, 32'h4262ffc5, 32'h4204c591, 32'h4294aeff};
test_bias[3065:3065] = '{32'hc2924e0a};
test_output[3065:3065] = '{32'h4504076f};
test_input[24528:24535] = '{32'hc29eb99b, 32'h4277c58d, 32'h41bb5503, 32'hc1f6ef0a, 32'hc1845dff, 32'hc23e6e5c, 32'h417adb1e, 32'h41bc0042};
test_weights[24528:24535] = '{32'h4239942e, 32'h424991dc, 32'h4286c53c, 32'h420ae538, 32'h42befd96, 32'hc224ffe9, 32'h426b2e50, 32'h40ad90a2};
test_bias[3066:3066] = '{32'h42acd561};
test_output[3066:3066] = '{32'h44b72102};
test_input[24536:24543] = '{32'hc279f032, 32'h42b2bee7, 32'hc103900a, 32'h4234cdc1, 32'hc2a53c49, 32'hbeb27e87, 32'hc29e5790, 32'h424717cd};
test_weights[24536:24543] = '{32'h429b1a2b, 32'hc27cb696, 32'h42a57722, 32'hc287566a, 32'h42a66e0c, 32'h42287710, 32'hc0435ed3, 32'hc2c7627e};
test_bias[3067:3067] = '{32'hc1a629e7};
test_output[3067:3067] = '{32'hc6ca0bec};
test_input[24544:24551] = '{32'h4193736c, 32'h42841ee1, 32'h4289f3c9, 32'hc1bdc593, 32'hc2b09b20, 32'h42a87879, 32'h429afdda, 32'hc2b1e0f7};
test_weights[24544:24551] = '{32'h42b91159, 32'h41af540f, 32'h42ac05ad, 32'hc19e019c, 32'h4204311e, 32'hc285cbcd, 32'h417f17e0, 32'hc2bbef6b};
test_bias[3068:3068] = '{32'hc1706a01};
test_output[3068:3068] = '{32'h46254c40};
test_input[24552:24559] = '{32'hc1e6ff03, 32'hc2436d24, 32'hc1b8a634, 32'h41d0d7f4, 32'hc2bc0142, 32'hc2091401, 32'h429ccb3d, 32'h42c370a7};
test_weights[24552:24559] = '{32'hc1dcf617, 32'hc2988787, 32'hc2b4d064, 32'hc2accaf3, 32'h425e50a3, 32'h42ad8de0, 32'hc29ca99d, 32'h4232ea43};
test_bias[3069:3069] = '{32'h40c6dc79};
test_output[3069:3069] = '{32'hc5af3ab5};
test_input[24560:24567] = '{32'hc1c9a3ed, 32'hc2a4d475, 32'h41db3e9a, 32'hc278dc27, 32'hc153cd99, 32'h4298d7cd, 32'hc29466ec, 32'hc21b1609};
test_weights[24560:24567] = '{32'h42847ecf, 32'h41cbd44e, 32'h42b60812, 32'hc178bce3, 32'h42963a75, 32'hc1bed8bb, 32'hc2463ac8, 32'h42ba103e};
test_bias[3070:3070] = '{32'hc186e90f};
test_output[3070:3070] = '{32'hc5400212};
test_input[24568:24575] = '{32'hc29a0a39, 32'hc2792be2, 32'hc273a1e7, 32'hc244e1de, 32'h42927a37, 32'hc2a88206, 32'hc1cd17ee, 32'hc23b0aef};
test_weights[24568:24575] = '{32'hc291059e, 32'h4242e9a8, 32'hc1be12dc, 32'hc2bffbca, 32'h406fe6c2, 32'h41bc9539, 32'h41c8f066, 32'hc2b3ba2f};
test_bias[3071:3071] = '{32'hc0b8ae03};
test_output[3071:3071] = '{32'h46250858};
test_input[24576:24583] = '{32'hc2048c23, 32'hc04a71e2, 32'h41d6bdd6, 32'hc0991803, 32'hc18120a7, 32'h4290d7f6, 32'hc2c2815e, 32'hc2680da4};
test_weights[24576:24583] = '{32'h4209a9e5, 32'h418236ec, 32'hc2bd7aad, 32'h42098318, 32'hc299d5da, 32'h4105747c, 32'h421e36b2, 32'hc130a855};
test_bias[3072:3072] = '{32'h423378d8};
test_output[3072:3072] = '{32'hc5a2f929};
test_input[24584:24591] = '{32'h4116a3f8, 32'hc204f875, 32'hc1202a10, 32'h428e97a8, 32'h4244f94c, 32'h4287a415, 32'hc2993017, 32'hc260de0f};
test_weights[24584:24591] = '{32'hc2be755f, 32'h42a14686, 32'h4287cb88, 32'hc2b28e0d, 32'hc2c4519b, 32'hc2861747, 32'h4238094e, 32'hc15c1cf2};
test_bias[3073:3073] = '{32'hc1f26803};
test_output[3073:3073] = '{32'hc6b1ff6d};
test_input[24592:24599] = '{32'h4234dbf2, 32'h420a4ad7, 32'hc2852767, 32'h426b0762, 32'h42933d72, 32'hc1341301, 32'hc10f98b6, 32'hc23118c1};
test_weights[24592:24599] = '{32'h42743db9, 32'hc215ae64, 32'hc27e8d8b, 32'h42b9a8ce, 32'h42042f1d, 32'hc28a4d62, 32'hc2ad199a, 32'hc22d172e};
test_bias[3074:3074] = '{32'hc13337c2};
test_output[3074:3074] = '{32'h468535c8};
test_input[24600:24607] = '{32'hc25ffae9, 32'hc1feccbd, 32'h42abc5f1, 32'hc19c30a3, 32'h42ad9f80, 32'hc2bb4311, 32'h41933c9e, 32'h4268a6db};
test_weights[24600:24607] = '{32'hc1b9894f, 32'hc25d770e, 32'hc229b238, 32'h42a7444c, 32'hc29679be, 32'h429066e6, 32'hc2986ad9, 32'hc2b4321c};
test_bias[3075:3075] = '{32'h42654aa4};
test_output[3075:3075] = '{32'hc6ac97a4};
test_input[24608:24615] = '{32'hc2c006d8, 32'hc277296d, 32'h42a1170e, 32'h429c812e, 32'h42a38672, 32'h4266ce7f, 32'h41d5911a, 32'h429fd0e7};
test_weights[24608:24615] = '{32'h42710f0d, 32'h41e7e35c, 32'hc2b86cea, 32'hc2afee7c, 32'hc20de340, 32'hc1ddfc69, 32'h4226712a, 32'hc21172d9};
test_bias[3076:3076] = '{32'h41e4b2d7};
test_output[3076:3076] = '{32'hc6dbf75f};
test_input[24616:24623] = '{32'hc2938763, 32'h428f9025, 32'h42686cc6, 32'h429fc7e9, 32'hc18b5de6, 32'hc2a8d31b, 32'hc2841133, 32'h41ca17cd};
test_weights[24616:24623] = '{32'hc247c4b0, 32'hc2b2859d, 32'hc193593e, 32'hc1da2621, 32'h424e1699, 32'h426d179b, 32'h42a9ad86, 32'h427fcc54};
test_bias[3077:3077] = '{32'h400e6ee0};
test_output[3077:3077] = '{32'hc677c622};
test_input[24624:24631] = '{32'h42177aae, 32'h41cc9d99, 32'h42660cec, 32'hc2984af8, 32'h428493ea, 32'hc26b9e1a, 32'hc104f822, 32'hc216eb54};
test_weights[24624:24631] = '{32'hc2bf4825, 32'h42c4814c, 32'hc28a07d9, 32'h426ad4de, 32'hc2bef232, 32'hc231e18a, 32'hc0eb8645, 32'hc22887dd};
test_bias[3078:3078] = '{32'hc1c75dfe};
test_output[3078:3078] = '{32'hc635bfd1};
test_input[24632:24639] = '{32'hc10ebb9e, 32'h41c39bac, 32'hc12f64d5, 32'hc17e2992, 32'h4186e6f5, 32'h42294c34, 32'h4188575c, 32'hc187e4a9};
test_weights[24632:24639] = '{32'hc16ddc30, 32'h41fdd19e, 32'hc2a19fa8, 32'h42bb00a5, 32'hc2a2eec7, 32'h42887053, 32'h429082c8, 32'hc261910f};
test_bias[3079:3079] = '{32'h41c5934c};
test_output[3079:3079] = '{32'h457c4989};
test_input[24640:24647] = '{32'h42b8f19c, 32'h417a4712, 32'hbfa27db7, 32'hc16b7676, 32'h41eda5b3, 32'h42812ec6, 32'h428e680a, 32'hc27e0eaf};
test_weights[24640:24647] = '{32'h42a1ddcd, 32'hc25247c0, 32'hc249c645, 32'hc1fbb9a2, 32'h405f5645, 32'hc2905aee, 32'hc061346b, 32'hc115c685};
test_bias[3080:3080] = '{32'h429e6bef};
test_output[3080:3080] = '{32'h453eda75};
test_input[24648:24655] = '{32'h42c1e615, 32'hc29ffc72, 32'hc2075179, 32'hc1e79d88, 32'h41dd4afb, 32'hc1442d65, 32'hbff5b054, 32'hc269594f};
test_weights[24648:24655] = '{32'hc2b0ee68, 32'h427b9b81, 32'hc18b1c7c, 32'hc1454b94, 32'h3fbcdec7, 32'h413642b4, 32'hc2a386df, 32'hc21d4e3c};
test_bias[3081:3081] = '{32'h42916c86};
test_output[3081:3081] = '{32'hc61ff895};
test_input[24656:24663] = '{32'hc293325b, 32'hc24ca670, 32'h41ccd6ac, 32'hc283351d, 32'hc2821ddb, 32'h4102dac5, 32'h42be3d55, 32'hc11573dc};
test_weights[24656:24663] = '{32'h42561068, 32'hc20a08db, 32'h42594bd1, 32'hc2c3d241, 32'hc202aa55, 32'h408f5196, 32'h41827367, 32'hc1a22e18};
test_bias[3082:3082] = '{32'h42b69d1b};
test_output[3082:3082] = '{32'h46168ac4};
test_input[24664:24671] = '{32'hc21cbbda, 32'h41caa9ae, 32'hc27e6a18, 32'hc2887478, 32'h42342af0, 32'hc28ef95d, 32'h40bea979, 32'hc2568464};
test_weights[24664:24671] = '{32'hc15f2730, 32'hc2c08eff, 32'hc24643e3, 32'h4138eda8, 32'h41aea3ed, 32'hc24899ba, 32'hc1890d4a, 32'h40f8d058};
test_bias[3083:3083] = '{32'h409238e7};
test_output[3083:3083] = '{32'h458d6abe};
test_input[24672:24679] = '{32'hc1f10206, 32'h429050b9, 32'h4222b3bf, 32'hc22f5002, 32'hc28ccc4b, 32'hc21b7cb4, 32'hc29ef7ce, 32'hc2a711b1};
test_weights[24672:24679] = '{32'h3faafd71, 32'h42c5b76d, 32'h4299f880, 32'h414dc38b, 32'h41f8af5a, 32'hc1ca8f42, 32'h42bb7393, 32'h41a48737};
test_bias[3084:3084] = '{32'h4296f91e};
test_output[3084:3084] = '{32'hc41edb9e};
test_input[24680:24687] = '{32'hc2c45210, 32'hc2bcccf4, 32'hc1a0d3c6, 32'h42b17016, 32'h41f2052e, 32'h42a86af4, 32'h42bf0626, 32'hc27b04c5};
test_weights[24680:24687] = '{32'hc10e494a, 32'hc1b10d78, 32'hc1885c87, 32'h42b657f4, 32'h41cc4376, 32'h42456077, 32'h41ed032f, 32'hc1b61e52};
test_bias[3085:3085] = '{32'hc1f0cb5d};
test_output[3085:3085] = '{32'h46a08aaa};
test_input[24688:24695] = '{32'hc2128a78, 32'hc2815a0e, 32'h414f57e6, 32'hc0d31b24, 32'hbedd325e, 32'hc2307988, 32'h408724cb, 32'h41cfa3c4};
test_weights[24688:24695] = '{32'hc29e69c7, 32'hc2435822, 32'hc02e8cb1, 32'h428df2b4, 32'h41088199, 32'hc1a8939d, 32'h4210e27e, 32'h41790d33};
test_bias[3086:3086] = '{32'h418949fe};
test_output[3086:3086] = '{32'h45dc86a4};
test_input[24696:24703] = '{32'hc2561376, 32'h427d52a3, 32'h429434c7, 32'h42bf0af2, 32'hc2608c10, 32'h4269a819, 32'hc1d17358, 32'h42648b66};
test_weights[24696:24703] = '{32'h4295e2c6, 32'hc23adfe3, 32'hc16f0358, 32'hc2be289c, 32'hc2664c3f, 32'hc216c91c, 32'h42b80de7, 32'h419b2c38};
test_bias[3087:3087] = '{32'h4292b8ae};
test_output[3087:3087] = '{32'hc68798d7};
test_input[24704:24711] = '{32'hc03286e6, 32'h424beaa2, 32'hc2b94ea7, 32'hc28b8d91, 32'h429af669, 32'hc21e59db, 32'h42aa3aab, 32'h408e3d15};
test_weights[24704:24711] = '{32'hc2bb8786, 32'h42841128, 32'h42ae30e4, 32'hc1965305, 32'hc2098b2b, 32'h409c267f, 32'h40971f90, 32'h4254e112};
test_bias[3088:3088] = '{32'h428c4122};
test_output[3088:3088] = '{32'hc5a4fbd5};
test_input[24712:24719] = '{32'hc28ddb2a, 32'hc2b1c2ec, 32'h42834cdd, 32'h41511542, 32'hc2826607, 32'h42852563, 32'hc22d64e9, 32'h4260fb44};
test_weights[24712:24719] = '{32'h42af3ea9, 32'h425c760b, 32'h426be809, 32'h4283e084, 32'h40d89e41, 32'hc1c3c1ae, 32'h410347cf, 32'h42b40faa};
test_bias[3089:3089] = '{32'hc1a9a729};
test_output[3089:3089] = '{32'hc56b387d};
test_input[24720:24727] = '{32'h426dba34, 32'hc0d9316f, 32'h4164d69c, 32'h408eb6a4, 32'hc20a2572, 32'hc1b98ab2, 32'hc0dec5e9, 32'h427a5d17};
test_weights[24720:24727] = '{32'hc22e5b99, 32'h4259e413, 32'h41850673, 32'h41a2bbeb, 32'h410925b8, 32'h4204b967, 32'hc2b51e2e, 32'h42440a2b};
test_bias[3090:3090] = '{32'h429d385e};
test_output[3090:3090] = '{32'h429e7fa5};
test_input[24728:24735] = '{32'h4040a90f, 32'h41bac7d0, 32'hc2a88b69, 32'h42c152a3, 32'hc19e6520, 32'hc2b3d938, 32'h421f0adf, 32'hc1e76d8b};
test_weights[24728:24735] = '{32'h4286bbf0, 32'h42ac6be9, 32'hc1978820, 32'h4153cdf7, 32'h41fb4852, 32'hc1940128, 32'h42a9c597, 32'hc0943a15};
test_bias[3091:3091] = '{32'h42b1df27};
test_output[3091:3091] = '{32'h46180ce9};
test_input[24736:24743] = '{32'hc2a75cd2, 32'h4262ce1a, 32'hc2a2fcc4, 32'h3f9eb4bd, 32'h42bb1494, 32'h41ea030d, 32'hc287f20c, 32'h3fbd58ba};
test_weights[24736:24743] = '{32'h42a3bf1e, 32'h41856eb2, 32'hc0bf1049, 32'h41df1820, 32'h4228bc81, 32'hc257afcf, 32'h4295292a, 32'hc1b2e97e};
test_bias[3092:3092] = '{32'hc1a1f6c4};
test_output[3092:3092] = '{32'hc5fe543a};
test_input[24744:24751] = '{32'hc2badb85, 32'hc2c48a84, 32'hc1ab1ca5, 32'hc23b8215, 32'h42362d7a, 32'hc1537c3c, 32'h427b5e7d, 32'h429762d4};
test_weights[24744:24751] = '{32'hc26cad4c, 32'h41a186f6, 32'hc207b178, 32'hc24e594e, 32'h42bc34cd, 32'h423e1c6f, 32'hc267c760, 32'hc2843b7a};
test_bias[3093:3093] = '{32'hc1b8b759};
test_output[3093:3093] = '{32'h44d18df6};
test_input[24752:24759] = '{32'hc19ac70f, 32'h4267b877, 32'h42702b70, 32'hc2c42b2c, 32'hc20709e5, 32'h4267d7a1, 32'h42bf8f5d, 32'h40c6d381};
test_weights[24752:24759] = '{32'h40ec9e7a, 32'h4280fbfd, 32'h42c23f2e, 32'hc2c69f76, 32'h42ad28b5, 32'hc2190349, 32'hc227dc69, 32'hc23c329a};
test_bias[3094:3094] = '{32'h42b9ce96};
test_output[3094:3094] = '{32'h461939de};
test_input[24760:24767] = '{32'hc234afae, 32'h428b7939, 32'h424bd6c1, 32'hc29a52f8, 32'h4280f51c, 32'hc2353016, 32'hc1af24c4, 32'h428f22c1};
test_weights[24760:24767] = '{32'h3fbc5fe5, 32'hc2454c28, 32'hc197eea7, 32'h42bb967c, 32'hc27d7240, 32'h42858287, 32'h40538490, 32'hc16286af};
test_bias[3095:3095] = '{32'h42a69d12};
test_output[3095:3095] = '{32'hc69addcd};
test_input[24768:24775] = '{32'hc2a08b27, 32'hc218d440, 32'h41b7f23d, 32'hc08eae33, 32'h42b401ae, 32'hc1c7fc94, 32'h428bc08d, 32'h420cfc42};
test_weights[24768:24775] = '{32'hc29efa5f, 32'hc1fea13e, 32'hc2b13a2e, 32'h425f080b, 32'hc22e294b, 32'h41dd15e4, 32'h42c1dca2, 32'h4247fc69};
test_bias[3096:3096] = '{32'h429e0d2e};
test_output[3096:3096] = '{32'h46118dc0};
test_input[24776:24783] = '{32'h426f94d5, 32'h4289788a, 32'h41844d99, 32'h4293d6ac, 32'hc2b425fd, 32'h427d7e7d, 32'hc1d79967, 32'h42b7ce82};
test_weights[24776:24783] = '{32'h42562269, 32'h42603d4f, 32'hc0c4241f, 32'h4262909d, 32'hc2a7c639, 32'hc29e5fee, 32'hc26645c7, 32'h4052f475};
test_bias[3097:3097] = '{32'hc1c77fd7};
test_output[3097:3097] = '{32'h4672616e};
test_input[24784:24791] = '{32'h4223c8ae, 32'h426c1b54, 32'hc293a720, 32'h420d10f8, 32'h42c4d48a, 32'hc2b0fe87, 32'h42c39c3c, 32'hc21034e1};
test_weights[24784:24791] = '{32'hc2a93fc5, 32'h41f46c16, 32'h429e3632, 32'hc2b42303, 32'h42b8d466, 32'hc2747750, 32'hc230b37d, 32'hc29753c3};
test_bias[3098:3098] = '{32'h42366da8};
test_output[3098:3098] = '{32'h450e6608};
test_input[24792:24799] = '{32'hc2a47ac6, 32'h42c7a310, 32'h415c36db, 32'hc28ed772, 32'hc25be0de, 32'h427f46a9, 32'h429c3d08, 32'h41872885};
test_weights[24792:24799] = '{32'h41abe5c9, 32'hc1f0de6c, 32'hc1b2cf55, 32'hc25b8527, 32'hc20e11f1, 32'h4296372c, 32'hc25a49b1, 32'hc1a61395};
test_bias[3099:3099] = '{32'hc19b6aba};
test_output[3099:3099] = '{32'h446df71d};
test_input[24800:24807] = '{32'hc11add55, 32'hc17f9ffb, 32'hc2b4191a, 32'hc219099d, 32'hc2bab362, 32'hc1339439, 32'h4158e116, 32'h40c92472};
test_weights[24800:24807] = '{32'h418c28be, 32'hc252cc5c, 32'h413251af, 32'h42950c00, 32'hc253cbde, 32'h420f2432, 32'hc185d8d4, 32'hbe80d99e};
test_bias[3100:3100] = '{32'hc286f29b};
test_output[3100:3100] = '{32'h4484dcd3};
test_input[24808:24815] = '{32'h42af6744, 32'h41d1c042, 32'h4296df45, 32'h41657ef0, 32'hc1a9ab7f, 32'hc2960caf, 32'hc21b4904, 32'h42a36d2a};
test_weights[24808:24815] = '{32'h3d8b2849, 32'h421ae426, 32'h42c089f9, 32'h4253131d, 32'h41b3095f, 32'hc2b89a3b, 32'hc290f564, 32'hc18902b5};
test_bias[3101:3101] = '{32'h420b1ae3};
test_output[3101:3101] = '{32'h46845739};
test_input[24816:24823] = '{32'hc285b182, 32'hc1c1b024, 32'hc23c1088, 32'hc2b90bd4, 32'hc217a23d, 32'hc13a9e78, 32'h42ba4924, 32'hc28b6fd5};
test_weights[24816:24823] = '{32'hc1e0f2ac, 32'h42a6a29a, 32'hc2c73666, 32'h4286899c, 32'h41b0bed9, 32'h40863890, 32'h425adbbd, 32'hc2aa5a1b};
test_bias[3102:3102] = '{32'hc137ecec};
test_output[3102:3102] = '{32'h46042923};
test_input[24824:24831] = '{32'h41443ef2, 32'h419d677e, 32'h41d1fb67, 32'h41cac028, 32'hc28abcef, 32'h42bf633d, 32'h4249f312, 32'h41dd4420};
test_weights[24824:24831] = '{32'hc27607ef, 32'hc2c2f55b, 32'hc2874915, 32'h42c28165, 32'h420edf28, 32'hc13538b1, 32'hc2755d16, 32'hc1c355e0};
test_bias[3103:3103] = '{32'hc283c224};
test_output[3103:3103] = '{32'hc6129b40};
test_input[24832:24839] = '{32'h4021946b, 32'h429f2421, 32'hc19ee5fe, 32'hc2b2a057, 32'hc270ab5d, 32'h42a29f20, 32'hc21a038d, 32'hc08d6c54};
test_weights[24832:24839] = '{32'hc26f35e6, 32'hc238b042, 32'h41887f88, 32'hc2aa5a43, 32'h428ec445, 32'hc2935e5c, 32'h4253c11c, 32'h4122146d};
test_bias[3104:3104] = '{32'hc2a1b396};
test_output[3104:3104] = '{32'hc60cbaaf};
test_input[24840:24847] = '{32'h4042c5e8, 32'hc159a0dd, 32'hc294e2c1, 32'hc270bcc7, 32'h420dfbac, 32'hc2989915, 32'h4238ec3d, 32'hc1a3650d};
test_weights[24840:24847] = '{32'h3f47748a, 32'hc1d78011, 32'h41d8a3a1, 32'hc01a0c54, 32'hc26d62d8, 32'h42188d52, 32'hc2c3755d, 32'h4292b223};
test_bias[3105:3105] = '{32'h424825b5};
test_output[3105:3105] = '{32'hc6431368};
test_input[24848:24855] = '{32'h428899d9, 32'h4262879b, 32'h429f1015, 32'h420f3289, 32'hc2be8424, 32'hc2bcdf22, 32'h4285808b, 32'h42b6e272};
test_weights[24848:24855] = '{32'h423f1688, 32'h428eb986, 32'hc2abe626, 32'h428fbb1c, 32'h42a1b142, 32'hc1eac5b4, 32'h42003706, 32'h4230f953};
test_bias[3106:3106] = '{32'hc206499f};
test_output[3106:3106] = '{32'h458539aa};
test_input[24856:24863] = '{32'h421170c5, 32'hc16c08f6, 32'h41dac3f6, 32'h415996bb, 32'hc212aaaa, 32'h426d51f6, 32'h4226fb99, 32'h4281c570};
test_weights[24856:24863] = '{32'hc288eeab, 32'h426c3898, 32'h422330d3, 32'hc23f9d58, 32'h4223411f, 32'h42b55711, 32'h4181bda5, 32'hc1edb047};
test_bias[3107:3107] = '{32'h428a93f6};
test_output[3107:3107] = '{32'hc3430195};
test_input[24864:24871] = '{32'hc2c43e60, 32'h428517e7, 32'h42018360, 32'h4120aa1a, 32'hc2878077, 32'hc25e508e, 32'h4221e88a, 32'hc283c3b3};
test_weights[24864:24871] = '{32'h41bf35c1, 32'h42a3c742, 32'hc2431b16, 32'h42ad3a7f, 32'h4298991c, 32'hc1bbb4cd, 32'h3e89b20e, 32'h415029a1};
test_bias[3108:3108] = '{32'hc238d84e};
test_output[3108:3108] = '{32'hc513b133};
test_input[24872:24879] = '{32'hc2a3f4e4, 32'h41cd7fd3, 32'hc21f73a0, 32'hc1c88683, 32'h41623ad5, 32'hc1ba5d9d, 32'hbf76b6d8, 32'hc1afc509};
test_weights[24872:24879] = '{32'hc1531087, 32'hc1d0f95f, 32'h42a9dd96, 32'hc0f69eab, 32'h42b04349, 32'hc2a6d55e, 32'hc1eba2dc, 32'h429ee363};
test_bias[3109:3109] = '{32'h41de067b};
test_output[3109:3109] = '{32'hc4a04150};
test_input[24880:24887] = '{32'hc234a4bd, 32'hc2a49af8, 32'h425f6d6b, 32'h429faf64, 32'h4289622a, 32'hc2714679, 32'h4227e339, 32'hc2ae8eda};
test_weights[24880:24887] = '{32'hc22d6443, 32'h420f0b8b, 32'hc2969eb1, 32'hc2026015, 32'h422a0061, 32'h42b376ec, 32'hc2b98ec0, 32'h428c3269};
test_bias[3110:3110] = '{32'h4123b458};
test_output[3110:3110] = '{32'hc69e835f};
test_input[24888:24895] = '{32'h42603c86, 32'h41f1e783, 32'hc2c10766, 32'hc2289d97, 32'h426a9217, 32'h4291afff, 32'hc2801b5c, 32'h40a942bc};
test_weights[24888:24895] = '{32'hc25a1357, 32'hc0dba709, 32'hc26f1d85, 32'h4295724a, 32'h42979f69, 32'h42851a28, 32'h41d8cf6d, 32'hc2bc65c2};
test_bias[3111:3111] = '{32'h41852499};
test_output[3111:3111] = '{32'h45c8ff01};
test_input[24896:24903] = '{32'h42b8749d, 32'h423e0ca4, 32'h4111ef38, 32'h42b3b806, 32'h4283cb54, 32'h422d1acb, 32'hc19f798e, 32'h42bb6ac3};
test_weights[24896:24903] = '{32'hc2b0c090, 32'hc298ba1c, 32'h41b494a9, 32'hc116ae8d, 32'h427ba644, 32'h42a7a13d, 32'hc277f4da, 32'hc27a5a14};
test_bias[3112:3112] = '{32'h423021b6};
test_output[3112:3112] = '{32'hc6103ea9};
test_input[24904:24911] = '{32'h4190c48c, 32'hbf8feb3b, 32'h40977676, 32'hc2b6147e, 32'hc0da32a9, 32'hc23a2a4b, 32'hc291e799, 32'h42902cdf};
test_weights[24904:24911] = '{32'hc29df896, 32'hc2b1ad20, 32'h4219458b, 32'h42ae827b, 32'h42bd894f, 32'hc224c809, 32'hc10b6240, 32'h426cef4a};
test_bias[3113:3113] = '{32'h4210b57a};
test_output[3113:3113] = '{32'hc533ef11};
test_input[24912:24919] = '{32'h3f68ddbd, 32'hc226c676, 32'hc2a2113a, 32'hc0185535, 32'hc255d0f5, 32'h42b11cfc, 32'hc26ca4f6, 32'h421cbdd7};
test_weights[24912:24919] = '{32'h428b7dfd, 32'hc18bb03c, 32'h4206f2d2, 32'h4249f10a, 32'hc2044174, 32'h42c37c06, 32'hc23a047d, 32'h42b562ef};
test_bias[3114:3114] = '{32'hc1c92ca8};
test_output[3114:3114] = '{32'h4664c21d};
test_input[24920:24927] = '{32'h4211c15c, 32'h41912d43, 32'hc24ac00c, 32'hc21d6dcf, 32'hc24eed37, 32'h4275d949, 32'h426eb743, 32'hc201fe6c};
test_weights[24920:24927] = '{32'hc234d358, 32'hc26f6647, 32'h429a7104, 32'h428698b2, 32'hc29a6cd9, 32'h42bbb321, 32'h41bc2821, 32'h42c5a969};
test_bias[3115:3115] = '{32'hc13d5c4b};
test_output[3115:3115] = '{32'hc4a935bd};
test_input[24928:24935] = '{32'hc2185478, 32'hbf21289f, 32'hc2a18f75, 32'hc15a064c, 32'h42ad7be5, 32'hc083090d, 32'hc29585d2, 32'h42a3f017};
test_weights[24928:24935] = '{32'hc223a4b2, 32'h4264584b, 32'hc24426d0, 32'h429fe84a, 32'hc21a3b25, 32'hc268d1c4, 32'h3fc5bdd0, 32'hc288ec9b};
test_bias[3116:3116] = '{32'hc2a11dec};
test_output[3116:3116] = '{32'hc58d41ab};
test_input[24936:24943] = '{32'hc240c8fb, 32'h427ddcd6, 32'hc2b27db6, 32'h41f8aed2, 32'h427c7932, 32'hc28a4ae0, 32'hc2609781, 32'hc2c316c1};
test_weights[24936:24943] = '{32'h4281205c, 32'h423a35ec, 32'hc29eca24, 32'hc2111b4d, 32'hc220bdd5, 32'h427ff9d1, 32'h4259cf32, 32'h41628263};
test_bias[3117:3117] = '{32'h41edab04};
test_output[3117:3117] = '{32'hc5ae09d3};
test_input[24944:24951] = '{32'h423d71fc, 32'hc2150202, 32'h4266b7cb, 32'h41ffef62, 32'h421f50c5, 32'h42af69d6, 32'h42707e83, 32'h427287e8};
test_weights[24944:24951] = '{32'h42201f6f, 32'h4140c380, 32'h4260705c, 32'h423c055d, 32'h418fe1bd, 32'hc0da9985, 32'hc2c7efcf, 32'h409a0e5d};
test_bias[3118:3118] = '{32'hc1ae1252};
test_output[3118:3118] = '{32'h440d0956};
test_input[24952:24959] = '{32'h421cb6ee, 32'h423d2ce7, 32'h42b5fec8, 32'hc21d8b12, 32'h4149591b, 32'h419a9212, 32'h4260b38f, 32'hc13cf3ab};
test_weights[24952:24959] = '{32'hc21c682a, 32'hc255fb93, 32'h41a65672, 32'hc29a44cb, 32'hc261abca, 32'h429c0bba, 32'hc23343ce, 32'h427f55fe};
test_bias[3119:3119] = '{32'h4284e4ee};
test_output[3119:3119] = '{32'hc4c06ba2};
test_input[24960:24967] = '{32'h408a058f, 32'hc154fb2d, 32'hc2a23178, 32'h4197cdb1, 32'h428fa0b6, 32'h40a3994a, 32'h422cdb2e, 32'hc28cd8b6};
test_weights[24960:24967] = '{32'h428f94f8, 32'h42a754e2, 32'h42887207, 32'hc050aabf, 32'hc2be2ffd, 32'hc22ee0df, 32'hc1a651d3, 32'h4218ab21};
test_bias[3120:3120] = '{32'h4109f17f};
test_output[3120:3120] = '{32'hc685098a};
test_input[24968:24975] = '{32'h41c25eba, 32'hc1cac759, 32'hc2020b28, 32'h4112155c, 32'hc2270d39, 32'h4234b21e, 32'hc0b0e7ff, 32'hc29834f4};
test_weights[24968:24975] = '{32'hc27de4a0, 32'h42bccd8d, 32'hc20fb797, 32'h4294f2be, 32'h4211fe00, 32'hc2615d98, 32'hc19291a4, 32'h4144eeff};
test_bias[3121:3121] = '{32'h4241f69b};
test_output[3121:3121] = '{32'hc5d8fa52};
test_input[24976:24983] = '{32'hc274eda7, 32'h415da8f0, 32'h417eeebf, 32'h42a16b8f, 32'h42577b5b, 32'h42ad0b26, 32'hc1c814e1, 32'hc160a588};
test_weights[24976:24983] = '{32'hc2b55fbd, 32'h42824872, 32'h4261d058, 32'hc23471d4, 32'h418e6745, 32'h421745df, 32'hc1e18254, 32'h41b9301a};
test_bias[3122:3122] = '{32'h428a37bf};
test_output[3122:3122] = '{32'h46032859};
test_input[24984:24991] = '{32'hc1873b59, 32'h4283fad7, 32'hc283fc0a, 32'h41b09c64, 32'h42441348, 32'hc1f0c486, 32'hc233034e, 32'hc294e95c};
test_weights[24984:24991] = '{32'hc28f8d47, 32'hc1fa2850, 32'hc2c65740, 32'hc2135827, 32'h41f82f18, 32'h4129cd13, 32'hc2b1a147, 32'hc2c1b2c4};
test_bias[3123:3123] = '{32'h4211e7da};
test_output[3123:3123] = '{32'h4687313c};
test_input[24992:24999] = '{32'h42c56c27, 32'hc1e21b50, 32'h4227e058, 32'h4107c4fa, 32'h42437e6c, 32'hc2bb580e, 32'h429854c5, 32'hc1ea1d3c};
test_weights[24992:24999] = '{32'h42c21991, 32'h42bc2d8d, 32'hc260a9bc, 32'hc2bed789, 32'h42945056, 32'hc28b03c2, 32'hc2442800, 32'h41aa1f51};
test_bias[3124:3124] = '{32'hc24118aa};
test_output[3124:3124] = '{32'h46142cf7};
test_input[25000:25007] = '{32'hc2c769b8, 32'hc215839d, 32'h429c116d, 32'hc2c32dd3, 32'h41cd451b, 32'hc0149dae, 32'hc1e9cfda, 32'hc1e855c9};
test_weights[25000:25007] = '{32'hc228b069, 32'hc20ee845, 32'h427e4037, 32'hc216b8d1, 32'hc2aa5692, 32'hc27eee27, 32'h4261da19, 32'hc193d98b};
test_bias[3125:3125] = '{32'hc28201eb};
test_output[3125:3125] = '{32'h462b46db};
test_input[25008:25015] = '{32'h41c43426, 32'hc230233b, 32'hc2a36399, 32'h426205da, 32'h40139305, 32'h428441f5, 32'h42bd3693, 32'h4297652c};
test_weights[25008:25015] = '{32'hc20453da, 32'hc24c8b3f, 32'hc23c74e4, 32'h42b9717d, 32'hc2b13392, 32'h421721dc, 32'h41329ec3, 32'h429aa738};
test_bias[3126:3126] = '{32'h41e57099};
test_output[3126:3126] = '{32'h469a6266};
test_input[25016:25023] = '{32'hc29e7c5e, 32'h42323243, 32'hc271cff1, 32'hc2b63739, 32'h423e8cd0, 32'hc223216e, 32'hc182b8df, 32'h42c0ad0f};
test_weights[25016:25023] = '{32'hc2794cbe, 32'h41a8532b, 32'hc2104e19, 32'h42971eed, 32'h4286d1d9, 32'hc22a5f8f, 32'hc2bcd045, 32'hc1e5138a};
test_bias[3127:3127] = '{32'h423fe508};
test_output[3127:3127] = '{32'h459ac9ee};
test_input[25024:25031] = '{32'h40e0161d, 32'h40efe4d3, 32'hc27ec964, 32'hc21f1ec8, 32'hc2392429, 32'h40df67c4, 32'h42acfc99, 32'h422b87d7};
test_weights[25024:25031] = '{32'h42a95e53, 32'h424fba3f, 32'h42ad937e, 32'h42764793, 32'hc2617f3d, 32'h42a03174, 32'hc2bb3488, 32'h3da49cdf};
test_bias[3128:3128] = '{32'hc1b85362};
test_output[3128:3128] = '{32'hc63a988e};
test_input[25032:25039] = '{32'hc1abec53, 32'h4228a089, 32'hc29d1581, 32'h42c14c33, 32'hc248ce6b, 32'h429866a7, 32'hc2371c55, 32'hc2381d5a};
test_weights[25032:25039] = '{32'h429aef8d, 32'hc2b51a3a, 32'h4281286f, 32'hc14d8bd5, 32'h42a0f4a3, 32'h410c4081, 32'hc1b33582, 32'h420d8b95};
test_bias[3129:3129] = '{32'h420a8085};
test_output[3129:3129] = '{32'hc675e322};
test_input[25040:25047] = '{32'h4085531d, 32'h428cc721, 32'h41fa94ac, 32'h4281441f, 32'hc189a209, 32'h3cedf37d, 32'hc253f614, 32'h41ce4c88};
test_weights[25040:25047] = '{32'h42438c2f, 32'h40eb740e, 32'hc2aed4a9, 32'h4291ce53, 32'h41d08cd9, 32'h428d2393, 32'h42ab7601, 32'h42b8718a};
test_bias[3130:3130] = '{32'h42c37a1a};
test_output[3130:3130] = '{32'h433608ac};
test_input[25048:25055] = '{32'h4259a391, 32'h420bb9c7, 32'hc1a30f53, 32'hc12ac16f, 32'h42c4ceb9, 32'hc2b673db, 32'hc2a80dff, 32'h424a9b24};
test_weights[25048:25055] = '{32'hc2242e10, 32'hc2802248, 32'hc25fe153, 32'h42a5cd4a, 32'h42af6a5e, 32'h4207ddc6, 32'hc220c727, 32'h4295d9cd};
test_bias[3131:3131] = '{32'h41230d9e};
test_output[3131:3131] = '{32'h4604ced8};
test_input[25056:25063] = '{32'hc28057ac, 32'hc2aad8af, 32'hc25888c1, 32'hc286628e, 32'hc209a851, 32'h423d803d, 32'hc280a187, 32'hc26ad808};
test_weights[25056:25063] = '{32'hc28ea05f, 32'h424f5630, 32'h426d5bbe, 32'h42070e8c, 32'h4243a5ff, 32'h41567f32, 32'h41add057, 32'h428db58c};
test_bias[3132:3132] = '{32'h411fe9b4};
test_output[3132:3132] = '{32'hc63a6018};
test_input[25064:25071] = '{32'h42b7b82a, 32'hc1a20d1c, 32'h427005a0, 32'h424195ce, 32'hc22d5ccc, 32'hc29733e9, 32'h419cee86, 32'h417490d6};
test_weights[25064:25071] = '{32'hc255e895, 32'hc260c2d9, 32'hc26b8286, 32'h42bcd15c, 32'h419c811e, 32'hc2be1b54, 32'hc0665fc0, 32'hc25f248d};
test_bias[3133:3133] = '{32'hc235568b};
test_output[3133:3133] = '{32'h45247885};
test_input[25072:25079] = '{32'h418f47eb, 32'hc2b186b0, 32'hc2ab3032, 32'hc264b706, 32'h41f24d84, 32'hc0daf215, 32'h427e7043, 32'hc2a1a6c9};
test_weights[25072:25079] = '{32'h418f6fd9, 32'h42a5d85a, 32'h428630f2, 32'hc2500210, 32'hc1cad966, 32'hc28580f2, 32'h429fc4a8, 32'h40aaa35f};
test_bias[3134:3134] = '{32'h4209cf1b};
test_output[3134:3134] = '{32'hc5a9daa8};
test_input[25080:25087] = '{32'hc2c139b3, 32'hc24dfc59, 32'hc10c4847, 32'h424eaa74, 32'hc2bb00fc, 32'hc2812603, 32'h41159ffc, 32'hc2863962};
test_weights[25080:25087] = '{32'h42287c97, 32'hc2c1dd40, 32'h42904919, 32'h42ae668d, 32'h4293e597, 32'hc1b86265, 32'hc2715790, 32'h429ef406};
test_bias[3135:3135] = '{32'h42abf0c5};
test_output[3135:3135] = '{32'hc5c9590c};
test_input[25088:25095] = '{32'h42ad552f, 32'h41dca32a, 32'hc1955842, 32'h42635f41, 32'h42b00f64, 32'h42191669, 32'h428058f5, 32'hc24089da};
test_weights[25088:25095] = '{32'h41cfddad, 32'hc2adca67, 32'h4289ebae, 32'h40b7ad23, 32'hc1e9f2b3, 32'h421bb824, 32'hc1fe6a59, 32'hc2859550};
test_bias[3136:3136] = '{32'h3fc2d2c4};
test_output[3136:3136] = '{32'hc47d9eec};
test_input[25096:25103] = '{32'hc2b3dd61, 32'hc28b7bad, 32'h423ce24e, 32'hc22fc9f7, 32'hc1c819f7, 32'hc2aca329, 32'h420b3a85, 32'hc1d80900};
test_weights[25096:25103] = '{32'hc18d7b2e, 32'hc19d1db3, 32'h428ccb02, 32'hc2aacafd, 32'h42af4135, 32'hc2ae6714, 32'hc2860f9e, 32'h41064565};
test_bias[3137:3137] = '{32'h410336b2};
test_output[3137:3137] = '{32'h46485426};
test_input[25104:25111] = '{32'h427d1210, 32'hc2139a26, 32'h41d7daaa, 32'hc10c9e9e, 32'h42854dc8, 32'h42b21d98, 32'hc0fbddc3, 32'hc201ed0e};
test_weights[25104:25111] = '{32'h416eb6d3, 32'h4276149d, 32'hc2620837, 32'h4159597e, 32'h417f7f2c, 32'h4287c52b, 32'hc1f4fc14, 32'hc26ab046};
test_bias[3138:3138] = '{32'h41f99a4d};
test_output[3138:3138] = '{32'h45c56dfd};
test_input[25112:25119] = '{32'hc2c72f5f, 32'h423467f0, 32'hc20728a2, 32'hc26859de, 32'h42837623, 32'hc17f8f10, 32'h42ab8b56, 32'hc25ad659};
test_weights[25112:25119] = '{32'h42254aef, 32'h42b0d17c, 32'hc29cb8e1, 32'h42c1ac82, 32'h42b2041d, 32'hc297ea8d, 32'h403275b7, 32'h42065e59};
test_bias[3139:3139] = '{32'h42824e16};
test_output[3139:3139] = '{32'h45178fad};
test_input[25120:25127] = '{32'hc25d409b, 32'hc26f7a01, 32'hc2a75675, 32'h4222b686, 32'h42204dc0, 32'h427523f7, 32'h4077e95e, 32'h419cf03b};
test_weights[25120:25127] = '{32'h41be89d7, 32'h42afd6d7, 32'hc1525fff, 32'hc289b7d6, 32'h41c36f7c, 32'hc2abb43d, 32'hc15d1e51, 32'hc21beed0};
test_bias[3140:3140] = '{32'h42563cc8};
test_output[3140:3140] = '{32'hc65044ae};
test_input[25128:25135] = '{32'h4264f224, 32'hc1f85021, 32'hc197c545, 32'h42090aa4, 32'h426dd190, 32'hc1ce3a7d, 32'hc2c181f9, 32'h41be127d};
test_weights[25128:25135] = '{32'h4049ca0f, 32'h42658ef2, 32'h426f531c, 32'hc21a9c41, 32'hc2a0487d, 32'hc2a833c1, 32'h40b59726, 32'hbf30d1f8};
test_bias[3141:3141] = '{32'h42a5335a};
test_output[3141:3141] = '{32'hc5df1ea8};
test_input[25136:25143] = '{32'hc2926711, 32'hc093febf, 32'hc2a3ce65, 32'hc239ccb8, 32'h428dbaa6, 32'hc2bb7f89, 32'hc2332bca, 32'h41cbf275};
test_weights[25136:25143] = '{32'h417c44a1, 32'h4118bf41, 32'h42493713, 32'hc19557f2, 32'hc1f1968c, 32'hc2903df2, 32'hc29120c5, 32'hc2058d85};
test_bias[3142:3142] = '{32'hc209d8bf};
test_output[3142:3142] = '{32'h451e6c3d};
test_input[25144:25151] = '{32'h429c3941, 32'h4292c58c, 32'h41c38c53, 32'hc146a083, 32'hc1d434fa, 32'hc21265ec, 32'h421880f7, 32'h429fc7bc};
test_weights[25144:25151] = '{32'h42918fdd, 32'hc24ecb37, 32'h41b05d66, 32'h428b7805, 32'hc1da0ad4, 32'hc2a6cdd1, 32'h42100062, 32'hc2ac1e4c};
test_bias[3143:3143] = '{32'hc136dfe8};
test_output[3143:3143] = '{32'hc32e6a96};
test_input[25152:25159] = '{32'h419ef7aa, 32'hc2b29f59, 32'h427905b7, 32'hc1351074, 32'hc1ebe274, 32'h424718de, 32'h429a66ae, 32'h4291e906};
test_weights[25152:25159] = '{32'h3edbd7e7, 32'h42b43089, 32'h41da3275, 32'hc252301e, 32'hc2a21840, 32'h4276ddd7, 32'hc1f7c121, 32'h42a56f81};
test_bias[3144:3144] = '{32'hc0d7b61e};
test_output[3144:3144] = '{32'h455196e1};
test_input[25160:25167] = '{32'hc25be6bf, 32'h42816e4e, 32'h415075e1, 32'h4284e832, 32'h42971404, 32'h3f9b40eb, 32'hc2447e6b, 32'h4267cc2a};
test_weights[25160:25167] = '{32'hc108dff2, 32'hc25898f4, 32'hc21a41f2, 32'hc2827591, 32'h41b13ebd, 32'h42bd472a, 32'h4263c43a, 32'h4130a0d2};
test_bias[3145:3145] = '{32'h41e1718a};
test_output[3145:3145] = '{32'hc6005036};
test_input[25168:25175] = '{32'hc292ba1e, 32'hc2bc1b8e, 32'h42ab5a66, 32'h4255a8ac, 32'h41fe20c1, 32'h412a3f13, 32'hc2140330, 32'h40586d2d};
test_weights[25168:25175] = '{32'hc289c674, 32'hc2a9c6c1, 32'hc230245d, 32'hc2a5f2cf, 32'hc298c23a, 32'hc21b5184, 32'hc290af34, 32'hc1e811b7};
test_bias[3146:3146] = '{32'hc1b3fc91};
test_output[3146:3146] = '{32'h458e2f35};
test_input[25176:25183] = '{32'h4183d904, 32'hc12f11db, 32'hc262a824, 32'hc114390f, 32'hc27dfc7a, 32'hc2c5b49a, 32'h42b56d3e, 32'h41e22b56};
test_weights[25176:25183] = '{32'h42b1b48b, 32'hc2a7217e, 32'hc2a62437, 32'hc03a4900, 32'h42991e8e, 32'h42207e68, 32'h424c4365, 32'h40bdb93b};
test_bias[3147:3147] = '{32'hc20f48ef};
test_output[3147:3147] = '{32'h453e965b};
test_input[25184:25191] = '{32'h41fce43b, 32'h4288531b, 32'h41534fc6, 32'h4268df26, 32'hc22fb536, 32'h4212544e, 32'h4237869f, 32'h42b8137d};
test_weights[25184:25191] = '{32'hc21db5aa, 32'hc2a6fd7c, 32'hc180eb54, 32'h428b5ae2, 32'h424b567f, 32'hc16f2188, 32'hc2a4149d, 32'h4279133d};
test_bias[3148:3148] = '{32'h40e88630};
test_output[3148:3148] = '{32'hc573b706};
test_input[25192:25199] = '{32'hc1cf02ef, 32'hc281f754, 32'hc22b4c77, 32'h429f3e3c, 32'hc29afb90, 32'hc21a7560, 32'h42b598ad, 32'h42212d38};
test_weights[25192:25199] = '{32'hc2b1e8c1, 32'hc2b84010, 32'h4215a71d, 32'h423d2873, 32'hc29f24b1, 32'hc218c605, 32'hc17aaacb, 32'h423f8341};
test_bias[3149:3149] = '{32'hc2bd4c66};
test_output[3149:3149] = '{32'h469090e5};
test_input[25200:25207] = '{32'h428d86d6, 32'h42235dd0, 32'h42a88f48, 32'hc1be70aa, 32'h40f9b64a, 32'h40fd1605, 32'hc1bcd925, 32'hc16b600d};
test_weights[25200:25207] = '{32'hc2a92c73, 32'hc29facf9, 32'h42957c66, 32'h40e2d8dc, 32'h427683b4, 32'h42b820ff, 32'h42911ef9, 32'h4244da71};
test_bias[3150:3150] = '{32'h41b31c25};
test_output[3150:3150] = '{32'hc5870970};
test_input[25208:25215] = '{32'hc2c79298, 32'hc2924a3d, 32'h42751ec0, 32'hc21e2d57, 32'hc1c06e3f, 32'hc213a684, 32'h42462e11, 32'hc21d6773};
test_weights[25208:25215] = '{32'hc2b55448, 32'hc2323b1e, 32'h41f5cddc, 32'hc2377002, 32'h42c0854c, 32'hc0546328, 32'hc29d031a, 32'h42513dec};
test_bias[3151:3151] = '{32'hc2511a69};
test_output[3151:3151] = '{32'h45f40ab4};
test_input[25216:25223] = '{32'h426bc59b, 32'h40b9fc7a, 32'h4295ca72, 32'h42847c8a, 32'hc28c1c76, 32'hc2c274c4, 32'h4231fa87, 32'hc2921cad};
test_weights[25216:25223] = '{32'h42693442, 32'hc0b098eb, 32'hc08eda4b, 32'hc1d8289b, 32'hc246ba01, 32'hc154deee, 32'hc25d7638, 32'hc194ed88};
test_bias[3152:3152] = '{32'hc1f152df};
test_output[3152:3152] = '{32'h4599c46f};
test_input[25224:25231] = '{32'hc1971369, 32'hc2354106, 32'hc2838f80, 32'h42a1d98f, 32'h42a8b8e5, 32'h426e1512, 32'hc2a7bece, 32'hc218d570};
test_weights[25224:25231] = '{32'hc167d08d, 32'h42605eda, 32'h41a6f2de, 32'h42319a63, 32'hc28bec74, 32'hc2b4e021, 32'h428b790b, 32'h424fe479};
test_bias[3153:3153] = '{32'h4244b4cd};
test_output[3153:3153] = '{32'hc6955cad};
test_input[25232:25239] = '{32'hc21f1889, 32'hc20ca47d, 32'hc298a7f5, 32'hc198e0a8, 32'h418e6963, 32'h42595f62, 32'hc29cc122, 32'hbfa97722};
test_weights[25232:25239] = '{32'h421a20fe, 32'h424a6871, 32'hc2041441, 32'hc24b4b49, 32'hc18d8312, 32'h410ce5b7, 32'h4195ab62, 32'hc2201f62};
test_bias[3154:3154] = '{32'h4277ae72};
test_output[3154:3154] = '{32'hc47bfe6b};
test_input[25240:25247] = '{32'hc08591b4, 32'h423cbadc, 32'h42ab1658, 32'h4121bfa5, 32'hbf8c4179, 32'h420f111d, 32'h42c4957c, 32'h4232ec00};
test_weights[25240:25247] = '{32'h4239d18b, 32'hc2959118, 32'hc1efd776, 32'h41be6f0a, 32'h42b755fa, 32'h41c69e92, 32'h40e336ad, 32'h428aa732};
test_bias[3155:3155] = '{32'hc1401236};
test_output[3155:3155] = '{32'hc4b7fbdf};
test_input[25248:25255] = '{32'h427bbc28, 32'h4291f277, 32'h41f244b5, 32'hc210784a, 32'hc2c14d7f, 32'h4283447e, 32'h40a02c5e, 32'hc202114a};
test_weights[25248:25255] = '{32'h42900a39, 32'hc2b919c1, 32'hc2864d88, 32'h42b8dae9, 32'h429b38cd, 32'hbfef72cf, 32'h42289105, 32'h418e538e};
test_bias[3156:3156] = '{32'hc2b1a1c0};
test_output[3156:3156] = '{32'hc674e5bf};
test_input[25256:25263] = '{32'h42b61f7c, 32'h41d85e59, 32'h427f0dad, 32'hc1f90238, 32'hc250f371, 32'hc2a30149, 32'hc0b53fa4, 32'hc2177cf9};
test_weights[25256:25263] = '{32'h42c15434, 32'h42b30ce3, 32'h410360c3, 32'h412b41fd, 32'h4179d21f, 32'h41a9a5b0, 32'hc2aaffd8, 32'hc26d9c5f};
test_bias[3157:3157] = '{32'h4276e15d};
test_output[3157:3157] = '{32'h46364768};
test_input[25264:25271] = '{32'hc20a53be, 32'h42aa020a, 32'hbf5f80d7, 32'hc20f603e, 32'h42743327, 32'h4180d2b6, 32'hc26caa75, 32'hc22d76ab};
test_weights[25264:25271] = '{32'hc16b2aa6, 32'h4233abde, 32'h4247ffb6, 32'hc2ba1a91, 32'h40bb285b, 32'hc299ac5c, 32'hc243c754, 32'h41d990b4};
test_bias[3158:3158] = '{32'h41ac5275};
test_output[3158:3158] = '{32'h46047002};
test_input[25272:25279] = '{32'h4294790b, 32'hc2669a38, 32'h428b5364, 32'hc26f96b9, 32'hc1889b9d, 32'h4288dd1e, 32'hc26aca26, 32'hc2815702};
test_weights[25272:25279] = '{32'hc2638812, 32'h41e97d41, 32'h4168b5b9, 32'hc2535294, 32'h42a953a8, 32'h40906266, 32'h42a0a6c8, 32'h4110d936};
test_bias[3159:3159] = '{32'hc1f2fd19};
test_output[3159:3159] = '{32'hc6000dd9};
test_input[25280:25287] = '{32'hc2989918, 32'h423995fd, 32'hc288607d, 32'h42b2304d, 32'hc1d2619f, 32'h42213252, 32'h42805619, 32'h4168c4a6};
test_weights[25280:25287] = '{32'hc2607c79, 32'hc2bf54a0, 32'hc2bd104f, 32'hc2c24ece, 32'h42534c32, 32'h4135a5c7, 32'h428fd156, 32'hc213ac31};
test_bias[3160:3160] = '{32'h416c627d};
test_output[3160:3160] = '{32'h44467a2f};
test_input[25288:25295] = '{32'hc2b22f95, 32'h4163c835, 32'h4201a4eb, 32'hc20e7de5, 32'h4282e60b, 32'hc272dfa7, 32'h410a9c9d, 32'hc181f526};
test_weights[25288:25295] = '{32'hc2313210, 32'hc1ac4191, 32'h42664ac6, 32'h423dcc76, 32'h423ef6d5, 32'h42b39ed8, 32'hc1d92c9c, 32'h41f93054};
test_bias[3161:3161] = '{32'h428eda73};
test_output[3161:3161] = '{32'h444c676f};
test_input[25296:25303] = '{32'h4269b3d5, 32'hc0e75ad6, 32'h4272e4d0, 32'h42855c20, 32'hc29a21b2, 32'hc12a7a91, 32'hc178617d, 32'h4280d3e5};
test_weights[25296:25303] = '{32'hc2061643, 32'hc19fb3d4, 32'h41059ccb, 32'hc249482e, 32'h402617f7, 32'hc2bc5052, 32'hc15a176c, 32'hc1e3861a};
test_bias[3162:3162] = '{32'hc20751a6};
test_output[3162:3162] = '{32'hc5ac4b7f};
test_input[25304:25311] = '{32'h42863bf8, 32'hc23728ae, 32'h42097ec4, 32'hc21aeedf, 32'h42a153c5, 32'hc28966e4, 32'hc1e9d92f, 32'h421e31f6};
test_weights[25304:25311] = '{32'h424fc493, 32'h41c5d7c0, 32'hc03f9501, 32'h428320fe, 32'h42c6ddca, 32'hc1d3df1a, 32'hc2a86206, 32'h4280f60f};
test_bias[3163:3163] = '{32'h3fb6a7a2};
test_output[3163:3163] = '{32'h46639033};
test_input[25312:25319] = '{32'hc24dd9d5, 32'h42256c28, 32'h416f75a4, 32'hc236f146, 32'h4148a65f, 32'h42a21d1a, 32'hc2bd0f4e, 32'hc205b3f2};
test_weights[25312:25319] = '{32'hc25a2966, 32'hc15745bd, 32'h424a6dd4, 32'h42a4a077, 32'hc27826e9, 32'h41e4e94d, 32'h40e6b902, 32'h42874ea9};
test_bias[3164:3164] = '{32'hc10e4cf1};
test_output[3164:3164] = '{32'hc50775a2};
test_input[25320:25327] = '{32'h41815b00, 32'hc29bfc41, 32'h41b6cacd, 32'h42a4dd21, 32'h41b5d540, 32'hc24a72ff, 32'hc2700139, 32'hbdf19d27};
test_weights[25320:25327] = '{32'h4202bd2f, 32'hbfb26d30, 32'h42039a15, 32'hc2117c72, 32'h42694b51, 32'hc23a65ed, 32'h42798d8d, 32'hc2aaa632};
test_bias[3165:3165] = '{32'hc1e681db};
test_output[3165:3165] = '{32'hc4d2e5c8};
test_input[25328:25335] = '{32'h42a9c404, 32'hc2599533, 32'hc2ac5778, 32'hc2473ba4, 32'hc2b75f61, 32'h4120a989, 32'h42b58578, 32'h4190f8f9};
test_weights[25328:25335] = '{32'hc276c330, 32'hc0061ed3, 32'h424bd9d9, 32'hc2990ea5, 32'h419f4e8a, 32'hc206dde9, 32'h41f2f927, 32'hc1066100};
test_bias[3166:3166] = '{32'h424e6987};
test_output[3166:3166] = '{32'hc5a2d4e9};
test_input[25336:25343] = '{32'hc251332a, 32'h41e388d3, 32'h41785c9e, 32'hc29f5c55, 32'h42c249d2, 32'h428578c1, 32'h42382db3, 32'hc0d48c42};
test_weights[25336:25343] = '{32'hc28fab8d, 32'h425593dd, 32'hc2b781ec, 32'h42b76fe3, 32'hc2a9a671, 32'hc29896f8, 32'hc2b52644, 32'h417e8751};
test_bias[3167:3167] = '{32'h41a04427};
test_output[3167:3167] = '{32'hc6a46995};
test_input[25344:25351] = '{32'hc21effdd, 32'h40a904d4, 32'h4183b6da, 32'h428cbfac, 32'h42b6a50d, 32'h42b846fc, 32'h429dae39, 32'h3e52574c};
test_weights[25344:25351] = '{32'h407b82d7, 32'h424737ff, 32'h42215cd3, 32'hc294960b, 32'hc287c66e, 32'hc17a01be, 32'hc06b28a1, 32'h42a93dd4};
test_bias[3168:3168] = '{32'h42b1379a};
test_output[3168:3168] = '{32'hc63fe168};
test_input[25352:25359] = '{32'h419085b0, 32'hc137f953, 32'h4247d014, 32'h427f1585, 32'h42948f31, 32'hc20bed91, 32'hc0ed8da4, 32'h42bd5a62};
test_weights[25352:25359] = '{32'h41501c19, 32'h423ef5f0, 32'hc284414d, 32'h42bdddc6, 32'hc29fb5dc, 32'hc0ea039c, 32'hc2a970a5, 32'h42367da7};
test_bias[3169:3169] = '{32'hc1bd2f76};
test_output[3169:3169] = '{32'h44d2b3bd};
test_input[25360:25367] = '{32'h41b07dc9, 32'h4292f300, 32'h42153c21, 32'h42b5e34e, 32'h41a51ad4, 32'h4221ebd2, 32'h429beed1, 32'h411cfd0b};
test_weights[25360:25367] = '{32'h42b138fd, 32'hc2b86bec, 32'hc251c3ed, 32'hc2aa6abd, 32'h42ad7315, 32'h42c03471, 32'h4289b313, 32'hc2544ce4};
test_bias[3170:3170] = '{32'h4125028f};
test_output[3170:3170] = '{32'hc57945d1};
test_input[25368:25375] = '{32'h42651d85, 32'h422ed6b6, 32'hc2b72155, 32'hc261d87e, 32'hc20ad55b, 32'h40630d3b, 32'hc2699e69, 32'h41cdcdbc};
test_weights[25368:25375] = '{32'h4204c20f, 32'hc2a42156, 32'h4202d78b, 32'h42be79f1, 32'h42a7d1bf, 32'h4180dcaa, 32'h40c085db, 32'hc0f27ab4};
test_bias[3171:3171] = '{32'hc2787d10};
test_output[3171:3171] = '{32'hc6534842};
test_input[25376:25383] = '{32'hc1a8c492, 32'h428b2982, 32'hc24a66e0, 32'h42705ba5, 32'h40c658df, 32'hc1fbee9e, 32'hc272b12f, 32'hc2c7930f};
test_weights[25376:25383] = '{32'h422ea622, 32'h42a3d4fb, 32'h429521d9, 32'h424fd78c, 32'hc1dca73c, 32'hc195cf3c, 32'hc2bc8e86, 32'h42248ddb};
test_bias[3172:3172] = '{32'h4138316e};
test_output[3172:3172] = '{32'h45c0e9cf};
test_input[25384:25391] = '{32'h4289973a, 32'h4293c3da, 32'h429f4cd1, 32'h426ff3e4, 32'h424829b9, 32'h42421cc7, 32'h429271b7, 32'h409c5f72};
test_weights[25384:25391] = '{32'h42c246bc, 32'hc181686b, 32'hc2555f8a, 32'h4231d450, 32'hc1f6a1ad, 32'hc13b1d14, 32'hc2088134, 32'h406963c8};
test_bias[3173:3173] = '{32'hc1a8217c};
test_output[3173:3173] = '{32'hc430a388};
test_input[25392:25399] = '{32'h42ab8457, 32'hc1f1380c, 32'h4274c69a, 32'h41d7a7b5, 32'h42b025ae, 32'h415ccb85, 32'hc2b1417d, 32'hc2af8b8b};
test_weights[25392:25399] = '{32'h4282faab, 32'h427806a7, 32'h41e06042, 32'hc2831d06, 32'h4188145c, 32'hc1260457, 32'h42a99c7c, 32'h42c00d8d};
test_bias[3174:3174] = '{32'h42b8ed6a};
test_output[3174:3174] = '{32'hc628c5ed};
test_input[25400:25407] = '{32'h42c166df, 32'h403cd4f1, 32'hc22834a3, 32'hc2ac202d, 32'hc1fe8e4d, 32'h42b6889a, 32'h42b8b3b5, 32'hc2bab1a0};
test_weights[25400:25407] = '{32'hbf17014e, 32'h413f7759, 32'hc29e2d62, 32'hc2905865, 32'h424713dd, 32'h413705d2, 32'h428a42a4, 32'h414a7b9f};
test_bias[3175:3175] = '{32'h41823609};
test_output[3175:3175] = '{32'h465dcbf4};
test_input[25408:25415] = '{32'h415ebd27, 32'h42ab99de, 32'h422f3b27, 32'hc26198c3, 32'hc2993087, 32'h4261425e, 32'hc2512e9e, 32'h4230f3cc};
test_weights[25408:25415] = '{32'h42a343fb, 32'hc2593d90, 32'h425646b9, 32'hc1e0c442, 32'hc17e76a2, 32'h428393bb, 32'hc2146065, 32'h42ab76c0};
test_bias[3176:3176] = '{32'h429758a7};
test_output[3176:3176] = '{32'h462e0c5a};
test_input[25416:25423] = '{32'h4212131a, 32'h4245099d, 32'h42a5f723, 32'hc220b434, 32'hc27d7c60, 32'hc20321d9, 32'h417e14b4, 32'hc0a9b7ec};
test_weights[25416:25423] = '{32'hc284edac, 32'hc2191b8e, 32'hc1c7e604, 32'h42adc816, 32'h4283225d, 32'h4233f001, 32'h42bf73ce, 32'h41766a43};
test_bias[3177:3177] = '{32'hc28a38ce};
test_output[3177:3177] = '{32'hc65ce655};
test_input[25424:25431] = '{32'hc28df51b, 32'hc2456b48, 32'h4237e121, 32'h4227c331, 32'hc1e5a7d5, 32'hc287ad9d, 32'h42757dc7, 32'h4119a996};
test_weights[25424:25431] = '{32'hc0ed78a8, 32'hc2364d5e, 32'h424742bd, 32'hc106ec94, 32'hc2b1fdcb, 32'h428ec40f, 32'h428a6408, 32'h42b3c7c6};
test_bias[3178:3178] = '{32'h42b1c8f9};
test_output[3178:3178] = '{32'h45ee3c90};
test_input[25432:25439] = '{32'hc1a7807e, 32'h41d645aa, 32'h41ac14d9, 32'hc2b2f9c7, 32'hc27d3f78, 32'hc299487c, 32'h42850010, 32'h424368fa};
test_weights[25432:25439] = '{32'hc2a43fa2, 32'h41a53842, 32'h4291874d, 32'hc0780ab6, 32'h42b1908d, 32'h4197bcbb, 32'hc2689284, 32'h409327e2};
test_bias[3179:3179] = '{32'h4283f89d};
test_output[3179:3179] = '{32'hc5ca0f21};
test_input[25440:25447] = '{32'hc22b21e6, 32'hc21c9d7e, 32'hc28ce0cc, 32'hc29def76, 32'h41c28ab2, 32'h418c3a41, 32'h41c43665, 32'h429f616d};
test_weights[25440:25447] = '{32'h4270e7f7, 32'h42b5ca26, 32'h4245c6a7, 32'h41ac7c73, 32'hc2874a59, 32'hc227eed6, 32'hc2c19e17, 32'hc1cec05a};
test_bias[3180:3180] = '{32'hc1d25141};
test_output[3180:3180] = '{32'hc68de406};
test_input[25448:25455] = '{32'hc184a13e, 32'hc2402920, 32'hc17a1e74, 32'h41f056e0, 32'hc2831877, 32'h4298d274, 32'h415cf410, 32'h3ff0d40a};
test_weights[25448:25455] = '{32'h42a5aa72, 32'hc28080c6, 32'h42a0b1eb, 32'hc1d0679f, 32'hc2c050d5, 32'hc1e9e695, 32'hc1c4d163, 32'h411c795c};
test_bias[3181:3181] = '{32'h42133258};
test_output[3181:3181] = '{32'h455830d4};
test_input[25456:25463] = '{32'hc2050637, 32'hc2347369, 32'hc205c648, 32'h41258533, 32'hc2766962, 32'h42a20428, 32'h42081711, 32'hc2839e4f};
test_weights[25456:25463] = '{32'hc298a123, 32'h4212c94c, 32'h41a98f73, 32'hc25f27dc, 32'hbf71cf01, 32'hc1f491c9, 32'hc1eab8aa, 32'h42156188};
test_bias[3182:3182] = '{32'h4226e5d4};
test_output[3182:3182] = '{32'hc5c2e028};
test_input[25464:25471] = '{32'h42163ad0, 32'hc2520fb3, 32'hc2911e53, 32'hc2986eed, 32'hc294abad, 32'hc1abe1f6, 32'h41f637a0, 32'h418657b2};
test_weights[25464:25471] = '{32'h42bd8db2, 32'hc141b095, 32'hc2494376, 32'h42bbc596, 32'h42a7d152, 32'hc2a9b63a, 32'hc2b4055c, 32'hc122f5d5};
test_bias[3183:3183] = '{32'h421fbaaf};
test_output[3183:3183] = '{32'hc5cf08b1};
test_input[25472:25479] = '{32'h42a3e23a, 32'hc218c29f, 32'hc285a439, 32'h42905ed4, 32'hc1dc50fa, 32'hc2abf444, 32'hc24ce34e, 32'h427289b5};
test_weights[25472:25479] = '{32'h41a36fad, 32'hc29d66e4, 32'h40ee98fe, 32'h41f79760, 32'hc2284809, 32'hc2920c16, 32'h41b84b03, 32'hc26f7cdd};
test_bias[3184:3184] = '{32'hc29629e2};
test_output[3184:3184] = '{32'h460c1c2a};
test_input[25480:25487] = '{32'h4282bcb0, 32'h42939ece, 32'hc1764098, 32'hc1c78d5b, 32'h40de9965, 32'h4233005a, 32'hc1671116, 32'hc1035bfa};
test_weights[25480:25487] = '{32'hc24fd373, 32'h41f9330e, 32'hc28064d6, 32'hc264f934, 32'h426c89f1, 32'hc2b6e088, 32'hc2c0ddb5, 32'h4213da0a};
test_bias[3185:3185] = '{32'h4255744c};
test_output[3185:3185] = '{32'hc49866eb};
test_input[25488:25495] = '{32'h42ae12f5, 32'hc27b8775, 32'hc212a9c8, 32'h4260ffb8, 32'h42073c10, 32'hc2bdbb04, 32'hc174feb5, 32'h4270366b};
test_weights[25488:25495] = '{32'hc2ab06cf, 32'h42c4a2ba, 32'hc2a71a93, 32'hc2c406d3, 32'hc2b7f048, 32'hbfb6fe3c, 32'h4261ef52, 32'h4230f5e6};
test_bias[3186:3186] = '{32'h42452c32};
test_output[3186:3186] = '{32'hc6866f24};
test_input[25496:25503] = '{32'h41a7184d, 32'h42541ebc, 32'hc299c600, 32'hc282c633, 32'hc23f3611, 32'h4279b38b, 32'h417c972a, 32'hc1320982};
test_weights[25496:25503] = '{32'hc0a04b39, 32'hc0ba252b, 32'h42a80145, 32'h4264078e, 32'hbf6d3d4a, 32'h41d145d0, 32'hc1c2beac, 32'hc2a807d1};
test_bias[3187:3187] = '{32'hc28196f7};
test_output[3187:3187] = '{32'hc603d113};
test_input[25504:25511] = '{32'hc1821bd0, 32'h421803e3, 32'hc2848f46, 32'hc262b97a, 32'hc26a53f2, 32'h426b93bc, 32'h4137dccc, 32'h42951517};
test_weights[25504:25511] = '{32'h401fb54a, 32'hc22c845f, 32'hbfe02445, 32'hc21c27da, 32'h4253ae32, 32'h41830992, 32'hc2678c88, 32'h42beaed2};
test_bias[3188:3188] = '{32'h4270ae34};
test_output[3188:3188] = '{32'h459cbc0b};
test_input[25512:25519] = '{32'h42008373, 32'h41fb9463, 32'hc2793dc2, 32'h419fb537, 32'h42b07324, 32'hc194f5d3, 32'hc0fdee1a, 32'h4280d374};
test_weights[25512:25519] = '{32'h424caaa7, 32'h41b64b70, 32'hc287faaa, 32'h422e11cf, 32'hc21c96ff, 32'hc226afb4, 32'hc1a992bd, 32'h42184580};
test_bias[3189:3189] = '{32'hc205b31a};
test_output[3189:3189] = '{32'h45e67582};
test_input[25520:25527] = '{32'h424837a4, 32'h422d012f, 32'hc193bac2, 32'h41fd98d1, 32'hc20ae9ae, 32'hc2684826, 32'hc2a92ab5, 32'hc2711ab3};
test_weights[25520:25527] = '{32'h42634316, 32'h429f0ca1, 32'h40e8ddd4, 32'hc28fe766, 32'h42501c8c, 32'h425cc3d1, 32'h4286dae8, 32'h42349dda};
test_bias[3190:3190] = '{32'h412878c1};
test_output[3190:3190] = '{32'hc6155856};
test_input[25528:25535] = '{32'h42bdc721, 32'h42a3c38e, 32'hc22e25c9, 32'hc2988820, 32'h42981169, 32'hc2b88f5e, 32'h428565f4, 32'h42121e2a};
test_weights[25528:25535] = '{32'h41dfa460, 32'h41edd87d, 32'h429d53bb, 32'hc2b136fd, 32'h41b42d38, 32'hc1128122, 32'h425d305a, 32'h41f9037d};
test_bias[3191:3191] = '{32'hc2879b9d};
test_output[3191:3191] = '{32'h4675dbb7};
test_input[25536:25543] = '{32'h40b35d2b, 32'hc284963c, 32'h4238035a, 32'h429a9e90, 32'hc2b1c6c1, 32'hc29554f0, 32'hc2c7f2d8, 32'hc203e414};
test_weights[25536:25543] = '{32'hc2a0510c, 32'hc288bcdf, 32'h425e40fb, 32'hc20de1ae, 32'hc15f088b, 32'h4280bfba, 32'hc2077f22, 32'hc1f6beed};
test_bias[3192:3192] = '{32'h417df267};
test_output[3192:3192] = '{32'h4594672c};
test_input[25544:25551] = '{32'h423d1564, 32'hc1e75813, 32'h42c3c796, 32'hc23938c8, 32'hc2813451, 32'hc10d6c4b, 32'hc176d9c3, 32'hc29dd7b1};
test_weights[25544:25551] = '{32'h42c1e915, 32'hc279a03d, 32'h42028df4, 32'h42ba52b9, 32'hc1abb797, 32'h4217934e, 32'h42c28582, 32'hc0ddd608};
test_bias[3193:3193] = '{32'h42165b83};
test_output[3193:3193] = '{32'h45a8e667};
test_input[25552:25559] = '{32'hc1bd4bf5, 32'hc2c55120, 32'h423bcb1e, 32'h423d62bc, 32'hc1d76eeb, 32'hc2c44242, 32'hc1b0c3e7, 32'hc1afb683};
test_weights[25552:25559] = '{32'hc2b008b7, 32'h42a6c227, 32'h4298d308, 32'h413ce236, 32'h421bc396, 32'hc12da431, 32'hc294b602, 32'h41b985f7};
test_bias[3194:3194] = '{32'h42227fb9};
test_output[3194:3194] = '{32'hc449a197};
test_input[25560:25567] = '{32'h41a47403, 32'h4156cd86, 32'hc25c2263, 32'h42804f03, 32'hc207200c, 32'h41d3faad, 32'h42ad9229, 32'h422812d8};
test_weights[25560:25567] = '{32'hc22128eb, 32'h422fd275, 32'hc282e7c9, 32'h408e4905, 32'hc13fc37f, 32'hc05e6f85, 32'h425d797b, 32'h41e631bd};
test_bias[3195:3195] = '{32'hc0947d35};
test_output[3195:3195] = '{32'h461bce7e};
test_input[25568:25575] = '{32'hc058c634, 32'hc0940363, 32'hc02bf4e5, 32'hc29a976a, 32'hc2a078c6, 32'hc1f483d5, 32'hbf4b3f18, 32'h42317afe};
test_weights[25568:25575] = '{32'hc29460ae, 32'hc1925920, 32'hc052fc80, 32'hc251c1c6, 32'h40d8a2a3, 32'hc283ee28, 32'hc119b587, 32'h42c2de45};
test_bias[3196:3196] = '{32'h42c6e68d};
test_output[3196:3196] = '{32'h4620f54c};
test_input[25576:25583] = '{32'hc2a3f045, 32'h42b53825, 32'h413232f8, 32'h426373fb, 32'h42bcbb64, 32'hc2823dad, 32'hc24d6d35, 32'hc2422031};
test_weights[25576:25583] = '{32'hc2211d57, 32'h41f86563, 32'hc2c1a8d3, 32'h427d093c, 32'h41ca2399, 32'h418e280d, 32'h40b47ec0, 32'hc210a269};
test_bias[3197:3197] = '{32'h429bb8dd};
test_output[3197:3197] = '{32'h46322fa3};
test_input[25584:25591] = '{32'hc161e351, 32'hc28695ce, 32'hc2986fe0, 32'h409c2cde, 32'h42a5b504, 32'hc2365eff, 32'hc154624c, 32'hc0928fae};
test_weights[25584:25591] = '{32'hc2565103, 32'hc1f02049, 32'h429845fb, 32'hc26369e9, 32'hc1bfd2a1, 32'hc2a7c94f, 32'hc2c08052, 32'h42259d45};
test_bias[3198:3198] = '{32'h4251a53f};
test_output[3198:3198] = '{32'hc3a2c570};
test_input[25592:25599] = '{32'h42a558f1, 32'hc1bcf100, 32'hc150328b, 32'hc2c0f73a, 32'hc287c50b, 32'hc20ca82d, 32'h4261cd96, 32'hc1c42244};
test_weights[25592:25599] = '{32'h42b0fc0d, 32'h40a7f445, 32'hc20f256d, 32'h428a8493, 32'h41a8f883, 32'hc2b52e8d, 32'h425d3d98, 32'hc226bd18};
test_bias[3199:3199] = '{32'h42573a06};
test_output[3199:3199] = '{32'h45d869b5};
test_input[25600:25607] = '{32'h3fbefece, 32'hc2afae48, 32'h42695ae1, 32'hc17c91f8, 32'hc2b032be, 32'h4240723c, 32'hc188a958, 32'hc29cbc39};
test_weights[25600:25607] = '{32'hc1e930d2, 32'h3f472ea3, 32'h41cb3ec8, 32'h42b5b7d4, 32'hc2c316a6, 32'h4238af87, 32'h42626195, 32'h42730e64};
test_bias[3200:3200] = '{32'hc0a2d9f4};
test_output[3200:3200] = '{32'h459cc924};
test_input[25608:25615] = '{32'hc27f44d9, 32'h4204a266, 32'h42b19375, 32'hc22a072a, 32'h4282f8d8, 32'hc18ad6fc, 32'h420e73b7, 32'h418c7657};
test_weights[25608:25615] = '{32'h41dc309a, 32'h41b32df9, 32'h42ac7ccb, 32'h4281d5b3, 32'hc249a2db, 32'hc078ecf1, 32'hc11f1d1e, 32'h40c70abf};
test_bias[3201:3201] = '{32'hc2024de6};
test_output[3201:3201] = '{32'h43ba84a1};
test_input[25616:25623] = '{32'hc151ba05, 32'hc268c6a7, 32'h429fd10b, 32'hc2178a31, 32'h422d3994, 32'h427e20e8, 32'hc1c22c6c, 32'h41d461c6};
test_weights[25616:25623] = '{32'h41ebb631, 32'hc28c49c6, 32'hc2b4f26c, 32'hc28ff1f3, 32'hc17a233b, 32'h4150a061, 32'hc2454df7, 32'hc16578a5};
test_bias[3202:3202] = '{32'hc2b25ac6};
test_output[3202:3202] = '{32'h428f0e17};
test_input[25624:25631] = '{32'h429c1c13, 32'h42311f20, 32'h429f99b9, 32'h40a70f68, 32'h41312d17, 32'h41bc9ac9, 32'h429cd3d0, 32'h40f0a523};
test_weights[25624:25631] = '{32'h4215a35f, 32'hc24fa372, 32'hc0ec6ab7, 32'hc0a243b1, 32'h4101a5a2, 32'hc2184cab, 32'h42b57c2b, 32'h4254b9b3};
test_bias[3203:3203] = '{32'hc16653e9};
test_output[3203:3203] = '{32'h45d153b3};
test_input[25632:25639] = '{32'h41f67e26, 32'hc230d8c7, 32'hc28e3154, 32'h42b7d54f, 32'hc124a427, 32'h4173159f, 32'h42b868c8, 32'hc1b57348};
test_weights[25632:25639] = '{32'hc26d4dd4, 32'hc1b47bf0, 32'h4288758a, 32'hc2c0361a, 32'h42bb1248, 32'h41f149a7, 32'hc12692cf, 32'h42811232};
test_bias[3204:3204] = '{32'hc2861465};
test_output[3204:3204] = '{32'hc688cc19};
test_input[25640:25647] = '{32'hc233b114, 32'h423654c1, 32'h424f1951, 32'hc225844c, 32'h421216ed, 32'hc2954cd6, 32'h41953571, 32'h42a39be2};
test_weights[25640:25647] = '{32'hc29b839b, 32'hc110d276, 32'h41ef81ba, 32'hc1a4012f, 32'h424e7531, 32'hc26377ed, 32'hc0c7bc8a, 32'h425373fe};
test_bias[3205:3205] = '{32'hc281024f};
test_output[3205:3205] = '{32'h46762254};
test_input[25648:25655] = '{32'h41f4924a, 32'hc2b2986c, 32'h4252afac, 32'h42bd2715, 32'h42a4bf44, 32'hc2a5cad1, 32'h412f8f4a, 32'hc2971a3b};
test_weights[25648:25655] = '{32'h42a6e4ff, 32'hc2493f29, 32'hc28b29b6, 32'hc2a18b18, 32'hc2762d2a, 32'hc2b15256, 32'h42270fc3, 32'h4281151e};
test_bias[3206:3206] = '{32'hc2224b92};
test_output[3206:3206] = '{32'hc5c93569};
test_input[25656:25663] = '{32'hc18cd357, 32'h428cc154, 32'h42a614e9, 32'hc1256a90, 32'hc146798e, 32'h41eca372, 32'h40838944, 32'h42459c8b};
test_weights[25656:25663] = '{32'h41f015f3, 32'h42a4b851, 32'h42aea153, 32'h41a3bc03, 32'hc1c245e8, 32'h408a36ed, 32'hc2053cd0, 32'h42b15e46};
test_bias[3207:3207] = '{32'hc2c5fff1};
test_output[3207:3207] = '{32'h4683e2ee};
test_input[25664:25671] = '{32'h41fe32d4, 32'h426e9d52, 32'h426e2f4e, 32'h42266338, 32'h42095a31, 32'hc28eeeb6, 32'h42ad44e0, 32'h42a6b9ec};
test_weights[25664:25671] = '{32'hc2c209c9, 32'hc2848007, 32'h424b041f, 32'hc28ea25a, 32'h4276bd07, 32'hc210ffa0, 32'hc21cdb74, 32'hc2875449};
test_bias[3208:3208] = '{32'h428c08c7};
test_output[3208:3208] = '{32'hc62f99d3};
test_input[25672:25679] = '{32'hc0fef4bf, 32'hc256ecbf, 32'h4205e973, 32'h41875694, 32'h42bd46a0, 32'hc20d6d06, 32'hc1af1b5f, 32'h41e8cb5c};
test_weights[25672:25679] = '{32'hc2c299c0, 32'h421f073d, 32'hc268f56b, 32'hc1b65ba1, 32'h419902ad, 32'hc2854ac6, 32'hc2c275b9, 32'hc23980b8};
test_bias[3209:3209] = '{32'hc083fb8f};
test_output[3209:3209] = '{32'h449b95e5};
test_input[25680:25687] = '{32'hc28dac84, 32'h42964e87, 32'h424ef1ee, 32'hc2a6fb34, 32'h4224d1b1, 32'h423af7f9, 32'hc22ecff2, 32'h41f3cfdd};
test_weights[25680:25687] = '{32'h41c9f860, 32'hc283bea2, 32'h42c15578, 32'h42bb33d2, 32'h417d15da, 32'hc1c094a7, 32'hbf0db102, 32'hc29fd4b2};
test_bias[3210:3210] = '{32'hc196bf29};
test_output[3210:3210] = '{32'hc642a0aa};
test_input[25688:25695] = '{32'h42485a54, 32'h417b08fa, 32'h422b09f6, 32'h41a51f0b, 32'h41b1179c, 32'h4266fa08, 32'hc1bc8532, 32'hc2a8a273};
test_weights[25688:25695] = '{32'hc0950c5c, 32'h41c1751f, 32'hc2866525, 32'h420efe1d, 32'hc2662063, 32'hc2c2cfda, 32'h4272308d, 32'h41d581d1};
test_bias[3211:3211] = '{32'hc19301a9};
test_output[3211:3211] = '{32'hc6449c25};
test_input[25696:25703] = '{32'h429d9ef4, 32'h41ce4b25, 32'h41204d11, 32'h426c3bb1, 32'h41cedeba, 32'hc21dfdf2, 32'hc2848f3c, 32'h42b67720};
test_weights[25696:25703] = '{32'h419f2aff, 32'hc112aa07, 32'hc2313c1f, 32'hc2631324, 32'h41740e4e, 32'h429d4d34, 32'h3f5ed859, 32'hc2bb6ee9};
test_bias[3212:3212] = '{32'hc26ce420};
test_output[3212:3212] = '{32'hc6584ff8};
test_input[25704:25711] = '{32'h42408ce5, 32'h41b05749, 32'hc2464d13, 32'h4187d207, 32'hbf261699, 32'h41b1bbd6, 32'hc2559413, 32'h429aefec};
test_weights[25704:25711] = '{32'h4236965e, 32'hc1d7e812, 32'h4239f77a, 32'h417b3139, 32'hc26ee9a6, 32'hc22ce17d, 32'h4199868f, 32'hc2be398e};
test_bias[3213:3213] = '{32'h42927824};
test_output[3213:3213] = '{32'hc61733f9};
test_input[25712:25719] = '{32'hc2bc049e, 32'hc2b5d42a, 32'h42a2eec9, 32'hc1d61787, 32'hc210753c, 32'h41a120af, 32'h41843813, 32'h429bd4d9};
test_weights[25712:25719] = '{32'hc29aad83, 32'hc108cc50, 32'hc0ea3ccf, 32'hc2262bfd, 32'hc2c4a87f, 32'h42337fe5, 32'h40e06e3b, 32'h42a26be2};
test_bias[3214:3214] = '{32'h42895fc0};
test_output[3214:3214] = '{32'h469894cf};
test_input[25720:25727] = '{32'h406a9544, 32'h42be0439, 32'hc248224a, 32'hc2bc0a6b, 32'h414e6ba3, 32'hc24dcac4, 32'h410e1b39, 32'hc279794e};
test_weights[25720:25727] = '{32'h42562d8c, 32'hc2132acd, 32'hc111d9f1, 32'h42a69265, 32'hc1b47aee, 32'hc2b2e0f3, 32'h428367ac, 32'h423722a7};
test_bias[3215:3215] = '{32'h4142caeb};
test_output[3215:3215] = '{32'hc606bc47};
test_input[25728:25735] = '{32'h429f9c35, 32'h4292c61b, 32'hc28d3c66, 32'hc26ccb41, 32'hc27f03e1, 32'hc27364de, 32'h4254d923, 32'h420b1446};
test_weights[25728:25735] = '{32'hc21af979, 32'h424deed8, 32'hc186c5b0, 32'hc2ae1672, 32'hc2177d85, 32'h42b7fd5b, 32'hc09df57c, 32'hc19f8a0e};
test_bias[3216:3216] = '{32'hc2620507};
test_output[3216:3216] = '{32'h45310ff4};
test_input[25736:25743] = '{32'h40f154de, 32'h425db871, 32'hbfa971d0, 32'hc221aed3, 32'hbf08598f, 32'h413d0d15, 32'h41e45259, 32'h422e6221};
test_weights[25736:25743] = '{32'h4239afce, 32'h42a657f3, 32'h42ba4eee, 32'hc228cf1e, 32'h4159e871, 32'hc242d896, 32'h409c81bc, 32'h428577e6};
test_bias[3217:3217] = '{32'h4258da0f};
test_output[3217:3217] = '{32'h460d9ca6};
test_input[25744:25751] = '{32'hc2aeb46e, 32'h4281cbfa, 32'h415f8381, 32'h428fc03a, 32'h41c48a18, 32'h41d893b2, 32'h42a55437, 32'hc0ad5ede};
test_weights[25744:25751] = '{32'hc2929147, 32'hc27a4f35, 32'hc2bcec02, 32'hc114f264, 32'hc22bd6dd, 32'h42313ea9, 32'hc281ecb8, 32'h41df15f5};
test_bias[3218:3218] = '{32'hc2a037a3};
test_output[3218:3218] = '{32'hc59f8b64};
test_input[25752:25759] = '{32'hc28ae37d, 32'hc2c7871b, 32'hc21c7fd1, 32'h4297a5c8, 32'hc0ac3617, 32'h42a43b27, 32'hc0ab0a9f, 32'hc2adc416};
test_weights[25752:25759] = '{32'hc25c7f25, 32'hc175e375, 32'hc2977a80, 32'hc11322c8, 32'h42ac3d08, 32'h41ed8b7e, 32'h4098432f, 32'h415ecdba};
test_bias[3219:3219] = '{32'h41782686};
test_output[3219:3219] = '{32'h4602f90c};
test_input[25760:25767] = '{32'hc2ad48a6, 32'hc2304f90, 32'h41c33e79, 32'hc1a4d7c1, 32'hc2802a74, 32'h42b217de, 32'h40eabd6b, 32'h41947ecd};
test_weights[25760:25767] = '{32'h422d0944, 32'h41bebfb3, 32'hc1bf5776, 32'h42b8602b, 32'h42391b9f, 32'hc2061528, 32'hc25f9372, 32'hc2622f5f};
test_bias[3220:3220] = '{32'h4261902b};
test_output[3220:3220] = '{32'hc664b001};
test_input[25768:25775] = '{32'hc28f65fc, 32'hc2a56128, 32'hc294c100, 32'hbfd01d10, 32'hc1255e68, 32'hc21e7ce5, 32'hc2852584, 32'h4286b7c7};
test_weights[25768:25775] = '{32'hc1cdbafa, 32'hc08adb90, 32'h4285a400, 32'h3e790aaf, 32'h422e214a, 32'hc2adb356, 32'hc235857a, 32'hc14d0c21};
test_bias[3221:3221] = '{32'hc1c4a8e4};
test_output[3221:3221] = '{32'h45134e9b};
test_input[25776:25783] = '{32'h42544d4c, 32'hc20f1963, 32'hc2427081, 32'h42390924, 32'h42bc7010, 32'hc194e35d, 32'h42b09b50, 32'h41cfea51};
test_weights[25776:25783] = '{32'hc06f3456, 32'h42c32fca, 32'hc2bcf671, 32'hc280910c, 32'hc2ab04e3, 32'hc2835a45, 32'hc18acfac, 32'hc209870e};
test_bias[3222:3222] = '{32'h42c670e7};
test_output[3222:3222] = '{32'hc62f7e30};
test_input[25784:25791] = '{32'hc1f0c745, 32'h428893b9, 32'hc28d1f00, 32'hc2adafdf, 32'hc235fee6, 32'hc2b83ec3, 32'hc28ddf98, 32'hc2ad574f};
test_weights[25784:25791] = '{32'h41a052b8, 32'h41da68be, 32'h409a8f6c, 32'h42216289, 32'hc2bde6bb, 32'h420b56fa, 32'hc25168eb, 32'hc1a5db27};
test_bias[3223:3223] = '{32'hc13319a4};
test_output[3223:3223] = '{32'h457bb045};
test_input[25792:25799] = '{32'h423211a3, 32'hc0d64a59, 32'h42aa036e, 32'h41b74b22, 32'hc290cf2d, 32'hc090bc2f, 32'h4161664d, 32'hc22e6644};
test_weights[25792:25799] = '{32'h42920bfa, 32'h4115377f, 32'hc2240ca9, 32'hc14ff435, 32'h41cb5718, 32'hc23a3107, 32'hc2a74cd7, 32'h40b7c2c7};
test_bias[3224:3224] = '{32'hc2a0bec8};
test_output[3224:3224] = '{32'hc5696be0};
test_input[25800:25807] = '{32'h40989925, 32'h41c92e00, 32'h4155d2ee, 32'hc285011b, 32'h4291ef80, 32'hc288bc00, 32'hc263a6b6, 32'h4036edb6};
test_weights[25800:25807] = '{32'h4269a0ba, 32'hc1bbbf64, 32'h42ad8221, 32'hc2a0864b, 32'hc295be4d, 32'h4249eeb7, 32'h42bfc8dd, 32'h42903093};
test_bias[3225:3225] = '{32'h42361291};
test_output[3225:3225] = '{32'hc5f7f965};
test_input[25808:25815] = '{32'hc2a5093f, 32'h41fb6585, 32'hc25d7e7d, 32'h425dcb2e, 32'hc201ebb2, 32'hc2b2fbeb, 32'h412b6215, 32'hc20066cb};
test_weights[25808:25815] = '{32'h40d1ab91, 32'hc21adc43, 32'h42586378, 32'hc2918857, 32'hc2a34532, 32'h4236e528, 32'h41109800, 32'h428d0237};
test_bias[3226:3226] = '{32'h4299f592};
test_output[3226:3226] = '{32'hc64075b9};
test_input[25816:25823] = '{32'hc21496a3, 32'h42b6ec22, 32'h4256bb91, 32'hc2b14fd2, 32'h419a90fc, 32'h4297bf78, 32'h41eaa6f4, 32'hc1832ae2};
test_weights[25816:25823] = '{32'h4284864c, 32'hc2c35cd3, 32'h41a32685, 32'hc269dff0, 32'hc2a017e7, 32'h42297acc, 32'hc1e333d5, 32'hc2c0f855};
test_bias[3227:3227] = '{32'h4272c839};
test_output[3227:3227] = '{32'hc524f42d};
test_input[25824:25831] = '{32'hc292a6d9, 32'hc225d87c, 32'hc1808c62, 32'h4218b6ff, 32'h42c72538, 32'hc2a2b00f, 32'h42972495, 32'hc23b255b};
test_weights[25824:25831] = '{32'h4123a2c4, 32'h426625d8, 32'hc29ec60b, 32'hc2849467, 32'h428a920f, 32'h42af8a19, 32'hc2213d6c, 32'h419475b9};
test_bias[3228:3228] = '{32'h42a03b8c};
test_output[3228:3228] = '{32'hc60446ea};
test_input[25832:25839] = '{32'h428f7cb6, 32'h420d94f0, 32'h41c13b74, 32'hc29d3dee, 32'hc2c247be, 32'h4037e51a, 32'h42867c8b, 32'hc025e564};
test_weights[25832:25839] = '{32'hc1653383, 32'hc0656e55, 32'h4275e07b, 32'h42ad2865, 32'h41b0a9bb, 32'hc271b062, 32'h41ba35a6, 32'h421cfc82};
test_bias[3229:3229] = '{32'h4232d82a};
test_output[3229:3229] = '{32'hc5e3bb45};
test_input[25840:25847] = '{32'hc2ac09ea, 32'h4234e4b0, 32'hc2884667, 32'h42aef078, 32'h42a84d83, 32'hc253f044, 32'hc1c6f7d0, 32'h4164b6e4};
test_weights[25840:25847] = '{32'h42bd095f, 32'h4280c34b, 32'hc25ceaf6, 32'h404ddc40, 32'h412ec0ed, 32'h429e21e4, 32'hc2b0c7c8, 32'hc1778f9a};
test_bias[3230:3230] = '{32'h427d72bb};
test_output[3230:3230] = '{32'hc5163f4b};
test_input[25848:25855] = '{32'h429d60ab, 32'hc2662e6e, 32'hc2b66d6b, 32'hc22e120a, 32'h4277592e, 32'h423ef910, 32'hc1c9cfbc, 32'hc29e7b31};
test_weights[25848:25855] = '{32'h41d1ed3f, 32'hc21cefaf, 32'h408577f1, 32'hc1f1952e, 32'hc2304046, 32'h4249cb1b, 32'hc02d365a, 32'h408e9175};
test_bias[3231:3231] = '{32'h42ab6393};
test_output[3231:3231] = '{32'h459428a0};
test_input[25856:25863] = '{32'hc22953f5, 32'hc1ff6e24, 32'hc22d99cb, 32'h42311d97, 32'hc268cecc, 32'hc2493c6b, 32'h42c7e9f8, 32'hc18d65b7};
test_weights[25856:25863] = '{32'hc2af7e20, 32'h42b52d61, 32'h42a1a8ad, 32'hc192d5a0, 32'hc2aace70, 32'hc27d5e2f, 32'h4294cee7, 32'hc2a12987};
test_bias[3232:3232] = '{32'hc281aee0};
test_output[3232:3232] = '{32'h46523d27};
test_input[25864:25871] = '{32'h423bd737, 32'h42899734, 32'hc2577641, 32'h41fcd0b1, 32'h42b67c64, 32'hc1d2613e, 32'hc1ba1455, 32'h429af869};
test_weights[25864:25871] = '{32'h42467167, 32'hc2c2957b, 32'hc25e177c, 32'hc2c233a0, 32'hc2be59cd, 32'h42a5fada, 32'h426556c4, 32'hc2ae8e9d};
test_bias[3233:3233] = '{32'hc264b08d};
test_output[3233:3233] = '{32'hc6b74ac3};
test_input[25872:25879] = '{32'h42b88ca4, 32'hc2aa0586, 32'hc1c432a0, 32'hc2036695, 32'hc2c016d3, 32'hc06b6a62, 32'hc283d625, 32'hc286dce7};
test_weights[25872:25879] = '{32'h42229b63, 32'hc219c3ec, 32'hc27329fb, 32'hc1b28e5f, 32'hc2847507, 32'hc2a28fc0, 32'h3f49f064, 32'hc2c26255};
test_bias[3234:3234] = '{32'hc21a4ca5};
test_output[3234:3234] = '{32'h46aebc7b};
test_input[25880:25887] = '{32'hc2a0799c, 32'h41eb534a, 32'hc297d0eb, 32'hc2856d55, 32'h429e5285, 32'h4244e3ae, 32'hc2997afa, 32'hc1de63d4};
test_weights[25880:25887] = '{32'h42a1c0c6, 32'hc2343326, 32'h427c5ef8, 32'hc2581921, 32'h425be555, 32'hc27c4156, 32'hc2b99d7a, 32'h41522389};
test_bias[3235:3235] = '{32'hc243070f};
test_output[3235:3235] = '{32'hc48276db};
test_input[25888:25895] = '{32'hc29e45d3, 32'h41a5b827, 32'hc2b8998e, 32'h41436708, 32'h428fa3ed, 32'hc2a2c9a5, 32'hc1a6f21c, 32'h40e3789f};
test_weights[25888:25895] = '{32'h422a1049, 32'hc1e31a37, 32'hc1bcd03a, 32'hc285d459, 32'h42762a0d, 32'hc2645732, 32'h428cb918, 32'hc2565c34};
test_bias[3236:3236] = '{32'h42207c00};
test_output[3236:3236] = '{32'h4591cdfb};
test_input[25896:25903] = '{32'hc24bc931, 32'hc2141521, 32'hc1317a78, 32'h42a91f90, 32'h424bb2fc, 32'hc298b3ed, 32'h42879a3e, 32'hc1a8ed89};
test_weights[25896:25903] = '{32'hc0730dc9, 32'h41f0a591, 32'h42c4ffcc, 32'hc2bce91e, 32'hc2362490, 32'hc212e7e0, 32'hc2174b69, 32'hc2124513};
test_bias[3237:3237] = '{32'hc1d6fec1};
test_output[3237:3237] = '{32'hc631180c};
test_input[25904:25911] = '{32'hc2997e9f, 32'hc15316be, 32'h410574ce, 32'h41187c4b, 32'h404b0538, 32'hc26b1013, 32'hc28f1716, 32'hc1a186ce};
test_weights[25904:25911] = '{32'h42b1f456, 32'hc2bfb105, 32'h41817559, 32'h428bb05c, 32'hc17314e4, 32'hc1a0570c, 32'hc1997854, 32'h426c86e2};
test_bias[3238:3238] = '{32'hc2643206};
test_output[3238:3238] = '{32'hc55b87db};
test_input[25912:25919] = '{32'hc1d942bf, 32'hc27b07ce, 32'hc28eeb54, 32'h3fd001fa, 32'hc2899620, 32'hc1e064cd, 32'hc1ae596c, 32'hc20fa028};
test_weights[25912:25919] = '{32'h42c188d7, 32'hc2c0b8e9, 32'h428cfb95, 32'h4293e78e, 32'hc210fd65, 32'hc155daf6, 32'h427ac7db, 32'hc2b808e9};
test_bias[3239:3239] = '{32'h411c442d};
test_output[3239:3239] = '{32'h454f63a3};
test_input[25920:25927] = '{32'h4282f291, 32'h421cbf29, 32'hc2aad6ed, 32'hc2303b21, 32'hc298ac11, 32'hc214db6e, 32'hc2225ffa, 32'h40c76e1c};
test_weights[25920:25927] = '{32'hc1982fdc, 32'hc2566098, 32'h3f73ae0c, 32'h4096ac82, 32'hc18e6f62, 32'h3b8037de, 32'hc2432b92, 32'h4204c759};
test_bias[3240:3240] = '{32'hc277a31c};
test_output[3240:3240] = '{32'hc315dd25};
test_input[25928:25935] = '{32'h42b27af6, 32'hc258fcaf, 32'h42ba0198, 32'h3f97578d, 32'hc2073a69, 32'h42bc12ca, 32'h42a1799a, 32'hbf18971e};
test_weights[25928:25935] = '{32'hc27ce3cf, 32'h42889f40, 32'hc1310be6, 32'h4299ed72, 32'h4246c98f, 32'h42c623e7, 32'h41e3af04, 32'hc06f2ce3};
test_bias[3241:3241] = '{32'hc20d44dc};
test_output[3241:3241] = '{32'hc3c0725b};
test_input[25936:25943] = '{32'hc11aeda9, 32'hc2ac10f8, 32'h427be6fc, 32'hc2c3e288, 32'h4195cf76, 32'hc24afc65, 32'hc13fa59e, 32'h40c2b62d};
test_weights[25936:25943] = '{32'h3ffddfe9, 32'h42bf22a6, 32'h42a8fb4d, 32'hc26e03f2, 32'h41c0fab4, 32'h428720da, 32'hc2c6903b, 32'h4236b0c0};
test_bias[3242:3242] = '{32'h4094e94a};
test_output[3242:3242] = '{32'h44af4e52};
test_input[25944:25951] = '{32'hc2a05d19, 32'hc08f4b87, 32'h42bd8b95, 32'hc1ab1546, 32'h428739e1, 32'h4242e205, 32'hc2c03a4a, 32'h41e7c75b};
test_weights[25944:25951] = '{32'h4296067f, 32'h41061a56, 32'h41583469, 32'h42b28db2, 32'hc1851c1b, 32'h4234206a, 32'hc26819fb, 32'hc27196e9};
test_bias[3243:3243] = '{32'h414824bd};
test_output[3243:3243] = '{32'hc4dd82aa};
test_input[25952:25959] = '{32'hc20ea1f5, 32'h42bb760f, 32'hc26915a7, 32'h424562c1, 32'h412b15c9, 32'hc2a8684c, 32'h42c53e3a, 32'h428ff238};
test_weights[25952:25959] = '{32'hc2917d83, 32'h42c3d0f0, 32'h4132b481, 32'hc2c52603, 32'h421b9355, 32'h42b2f05f, 32'hc2471d87, 32'h42299731};
test_bias[3244:3244] = '{32'hc1e9a502};
test_output[3244:3244] = '{32'hc52bcf09};
test_input[25960:25967] = '{32'h42a60d60, 32'h425697d9, 32'h42b15546, 32'h4285e118, 32'hc113371d, 32'h41cca958, 32'h428e5feb, 32'hc0758ecc};
test_weights[25960:25967] = '{32'hc1b785eb, 32'hc28b3684, 32'hc1676c49, 32'hc2a88e80, 32'hc292f50a, 32'h421881e3, 32'hc21c8ea7, 32'hc28f4b1a};
test_bias[3245:3245] = '{32'hc12d9d57};
test_output[3245:3245] = '{32'hc651e6a7};
test_input[25968:25975] = '{32'hbf1fe3ac, 32'hc2b75aa0, 32'hc2317d8a, 32'hc2935601, 32'h41f813e5, 32'hc245fe79, 32'h4260c7b0, 32'hc1b5dc5f};
test_weights[25968:25975] = '{32'h418bcc45, 32'h4200174c, 32'h41cd4f05, 32'hc17015f7, 32'h406dfece, 32'h42613c0e, 32'h4294d7ad, 32'hc2a3a141};
test_bias[3246:3246] = '{32'hc28216ca};
test_output[3246:3246] = '{32'h43a284ae};
test_input[25976:25983] = '{32'h429b02f5, 32'hc1cf0476, 32'h42011266, 32'h4276089f, 32'hc291e6ea, 32'h42683b1b, 32'hc24b0efd, 32'h427fbd41};
test_weights[25976:25983] = '{32'h419160f2, 32'hc2867e96, 32'hc1deead4, 32'hc29f5d92, 32'h41319a0a, 32'hc1bbca09, 32'hc2168530, 32'h42a6e315};
test_bias[3247:3247] = '{32'hc0f5005d};
test_output[3247:3247] = '{32'h4516d4f4};
test_input[25984:25991] = '{32'hc2b5f917, 32'hc204cfe9, 32'h4199ddeb, 32'hc282be8c, 32'hc28120c6, 32'h42b0ab06, 32'hc20d5f21, 32'hc29ab10b};
test_weights[25984:25991] = '{32'hc2be8f39, 32'h427eed63, 32'h42afcb76, 32'hc2a0cdcc, 32'h41ecfeb7, 32'h42b1734a, 32'hc0b63b9d, 32'h42ac43fb};
test_bias[3248:3248] = '{32'h428aa4e7};
test_output[3248:3248] = '{32'h464ba43d};
test_input[25992:25999] = '{32'h42813f3e, 32'h41bcec17, 32'hc1a6a398, 32'h428b5000, 32'hc25b45c6, 32'hc2ad0795, 32'h429505d6, 32'hc2c3aa01};
test_weights[25992:25999] = '{32'hc2ab062b, 32'h3f0eef40, 32'h42c75979, 32'hc2aadd31, 32'h415adb12, 32'hc1b441b6, 32'hc286352b, 32'h423e3876};
test_bias[3249:3249] = '{32'h4236c1cc};
test_output[3249:3249] = '{32'hc6ab7661};
test_input[26000:26007] = '{32'hc2b0ec1a, 32'h42be6c4b, 32'h428ed1c8, 32'h42b9f135, 32'hc167c960, 32'hc221f8ae, 32'h41fb4122, 32'hc18016bf};
test_weights[26000:26007] = '{32'hc20c1201, 32'h41e906d6, 32'hc0976fcb, 32'h4120061b, 32'h4255c6b3, 32'h420a1b75, 32'h42911e67, 32'h41e42a9b};
test_bias[3250:3250] = '{32'hc2198b79};
test_output[3250:3250] = '{32'h45bdd3ba};
test_input[26008:26015] = '{32'h42b9eb48, 32'h41af6851, 32'hc187de59, 32'hc1b6e03d, 32'h408cfab4, 32'hc253de33, 32'h3fd1ea1f, 32'h42b0b03d};
test_weights[26008:26015] = '{32'h425ca7fc, 32'h42657306, 32'hc21329e2, 32'hc2930cf4, 32'hc299d843, 32'hc23379cf, 32'hc20197f1, 32'hc21c80d4};
test_bias[3251:3251] = '{32'hc2754cd8};
test_output[3251:3251] = '{32'h45dfb037};
test_input[26016:26023] = '{32'h4292535c, 32'h424b9975, 32'hc1c37a38, 32'hc1544014, 32'hc2a63c35, 32'hc265e460, 32'hc25b68e7, 32'h420030b2};
test_weights[26016:26023] = '{32'h41aa318c, 32'h42996243, 32'hc130d42b, 32'h42b9ab0a, 32'hc21167a0, 32'hc27ca5cf, 32'h40b1c9c2, 32'h420c3d0a};
test_bias[3252:3252] = '{32'h429728a7};
test_output[3252:3252] = '{32'h463c323f};
test_input[26024:26031] = '{32'hc18ec19a, 32'hc1bf223f, 32'hc1f446e2, 32'hc25543ee, 32'h42b27c6c, 32'h42912a90, 32'hc23bc0e4, 32'hc270b302};
test_weights[26024:26031] = '{32'hc22db881, 32'hc28bf36b, 32'hc20a8862, 32'h4197f3f7, 32'hc2b72985, 32'h41ed1247, 32'h429d7e3a, 32'hc28e8a00};
test_bias[3253:3253] = '{32'h421fa433};
test_output[3253:3253] = '{32'hc53521a8};
test_input[26032:26039] = '{32'hc1088286, 32'hc13a4378, 32'hc2c7cf4c, 32'h41bc5586, 32'h428775d1, 32'h42c7bf5d, 32'h41cfa4c2, 32'h42628534};
test_weights[26032:26039] = '{32'hc29ff64c, 32'hc28dbbdb, 32'h42469005, 32'h4204c678, 32'h42ac5bbd, 32'hc1d86c12, 32'hc239c36b, 32'hc228fe7b};
test_bias[3254:3254] = '{32'hc20bcc4b};
test_output[3254:3254] = '{32'hc546055a};
test_input[26040:26047] = '{32'hc2c2f683, 32'h423de4a4, 32'h4248db88, 32'hc211533c, 32'h416e3051, 32'hc2adb30c, 32'hc2921b96, 32'h428a18ff};
test_weights[26040:26047] = '{32'h416fb2b0, 32'h41f9accc, 32'h420cd086, 32'hc232ccce, 32'hc200c4d2, 32'h42019ea3, 32'h42a5dee8, 32'h422cee07};
test_bias[3255:3255] = '{32'h42c7870c};
test_output[3255:3255] = '{32'hc5326774};
test_input[26048:26055] = '{32'h42b3bfd1, 32'hc2297bea, 32'hc1d0d523, 32'h41cf9586, 32'h419f5b7e, 32'h42967c31, 32'h4236d03f, 32'hc22b34a0};
test_weights[26048:26055] = '{32'hc2b689c4, 32'hc2aaa748, 32'h4159648b, 32'hbedb2b3d, 32'h40a51553, 32'h41f20e68, 32'h4019fad1, 32'hc1c0fc71};
test_bias[3256:3256] = '{32'hc265b224};
test_output[3256:3256] = '{32'hc4ba1838};
test_input[26056:26063] = '{32'h4296d498, 32'hc22630f0, 32'h408d34da, 32'hc29dfa61, 32'hc25c003a, 32'h4176c991, 32'h418a85ec, 32'hc214910f};
test_weights[26056:26063] = '{32'hc06cab2e, 32'h417f74ba, 32'h42368934, 32'h42365c3b, 32'hc1af8982, 32'h42c34b22, 32'hc2a01a2e, 32'hc257ecd4};
test_bias[3257:3257] = '{32'hc284030c};
test_output[3257:3257] = '{32'hc486866e};
test_input[26064:26071] = '{32'h4207ca9b, 32'hc24ea94e, 32'hc121bc0f, 32'h427f6ded, 32'h41691720, 32'hc2866eac, 32'h422b3041, 32'h40cda458};
test_weights[26064:26071] = '{32'hc26b9552, 32'h41d2d820, 32'hc24e5315, 32'hc26c09e1, 32'h421fd125, 32'h410c328f, 32'h41e0ccef, 32'h419b0c52};
test_bias[3258:3258] = '{32'h42ad3ea8};
test_output[3258:3258] = '{32'hc5a287eb};
test_input[26072:26079] = '{32'h425dab26, 32'hc29ab2f6, 32'h423d1d21, 32'hc280569a, 32'hc2adbebb, 32'h42be2e5a, 32'hc1d0ce6a, 32'h42b12e24};
test_weights[26072:26079] = '{32'h421d0bf4, 32'hc2a8ca5e, 32'h4215f8a4, 32'hc2090f98, 32'hc2889d2d, 32'h42b52f84, 32'hc230a075, 32'h4211eeae};
test_bias[3259:3259] = '{32'h42af5c13};
test_output[3259:3259] = '{32'h46f79fad};
test_input[26080:26087] = '{32'h42afdf08, 32'hc23643f4, 32'hc2bb6076, 32'h42a1fd40, 32'hc25a1d51, 32'hbfa167d5, 32'hc05975ce, 32'hc134ec66};
test_weights[26080:26087] = '{32'hc1d55073, 32'hc21e8e86, 32'hc2939fd5, 32'hc2c36840, 32'h42b10970, 32'h424c0f33, 32'hc1eda743, 32'h4131ccd2};
test_bias[3260:3260] = '{32'h41a7722d};
test_output[3260:3260] = '{32'hc5c8fc73};
test_input[26088:26095] = '{32'h41ddda92, 32'h419694a6, 32'hc26b4f4d, 32'h427e4ef7, 32'h42318186, 32'h42a39394, 32'h427ed5b2, 32'hc18beec3};
test_weights[26088:26095] = '{32'hc11a8e7d, 32'hc187fe46, 32'h4101aa52, 32'hc2b5c01f, 32'h42c6de0a, 32'hc213f118, 32'h411de580, 32'h420de95a};
test_bias[3261:3261] = '{32'h42845fb4};
test_output[3261:3261] = '{32'hc5a8226b};
test_input[26096:26103] = '{32'h4236f86e, 32'hc1933241, 32'hc1376116, 32'h42656368, 32'hc1f4fac7, 32'h420b0b91, 32'h41d0b4e2, 32'hc27655ee};
test_weights[26096:26103] = '{32'hc1447bef, 32'hc0e25d33, 32'hc2b6c270, 32'h423bb332, 32'hc2884ed3, 32'hc17b391d, 32'h429437d5, 32'h416fe5b0};
test_bias[3262:3262] = '{32'h413e901b};
test_output[3262:3262] = '{32'h45b76f65};
test_input[26104:26111] = '{32'hc2a34663, 32'h422ddc4d, 32'h4217c08a, 32'h41e35add, 32'h423fb2f9, 32'h428ea920, 32'h41f6ca79, 32'hc20b7847};
test_weights[26104:26111] = '{32'hc2988304, 32'h4150849b, 32'h4282c521, 32'h42755644, 32'h42c03740, 32'hc1bd34f4, 32'h409ff6a1, 32'h42621ee2};
test_bias[3263:3263] = '{32'hc2b44073};
test_output[3263:3263] = '{32'h463bed98};
test_input[26112:26119] = '{32'hc1cfdcb3, 32'hc2c00a30, 32'hc2b7d17d, 32'h427abd0b, 32'h4269e4e8, 32'h4268850e, 32'hc1121413, 32'h3fb918cf};
test_weights[26112:26119] = '{32'hc245748a, 32'hc25459b7, 32'hc061b369, 32'h417cf848, 32'h42bd51c9, 32'h42208e68, 32'hc27ade59, 32'h42c697fc};
test_bias[3264:3264] = '{32'hc2ac0a65};
test_output[3264:3264] = '{32'h467d074c};
test_input[26120:26127] = '{32'h42687bfc, 32'hc29b6ed9, 32'h4238654a, 32'h424ec85e, 32'hc122eb1b, 32'h4201c9b6, 32'hc2a08993, 32'hc0deda28};
test_weights[26120:26127] = '{32'hc28efadc, 32'hc23b433e, 32'hc2097204, 32'h41947ac1, 32'hc2c04991, 32'hc282cdc9, 32'h408a9779, 32'h41ba6ace};
test_bias[3265:3265] = '{32'h41855ba9};
test_output[3265:3265] = '{32'hc52d9a68};
test_input[26128:26135] = '{32'hc2be42c4, 32'hc22a0af2, 32'hc24f9894, 32'h4231f92a, 32'hc21a8abc, 32'hc09cbd97, 32'hc212ac80, 32'hc28d1890};
test_weights[26128:26135] = '{32'hc1bf798e, 32'h421206bd, 32'h419b3e32, 32'h421b5f02, 32'hc1b6d8c9, 32'hc2697a3c, 32'h428831e2, 32'hc2ba48fd};
test_bias[3266:3266] = '{32'h414ddad9};
test_output[3266:3266] = '{32'h45d16f29};
test_input[26136:26143] = '{32'hc13fd474, 32'h427c46d9, 32'hc18dd707, 32'hc0a02240, 32'hc24e2cd7, 32'h4269373a, 32'h422c82ab, 32'hc2b4b855};
test_weights[26136:26143] = '{32'hc16d4935, 32'hc29ca9fe, 32'h427cfcec, 32'hbef1dd84, 32'h4198f6f0, 32'hc1d49cab, 32'h42482956, 32'hc26ab32e};
test_bias[3267:3267] = '{32'h4258f3c9};
test_output[3267:3267] = '{32'hc461974a};
test_input[26144:26151] = '{32'hc1faba12, 32'h416b52af, 32'hc23defb1, 32'hc20c2c9e, 32'hbd968177, 32'h42166795, 32'h42899724, 32'hc279571d};
test_weights[26144:26151] = '{32'hc15ec435, 32'hc28edce9, 32'h4155490c, 32'hc03a27f5, 32'hc250dc60, 32'hc2744137, 32'hc25be21d, 32'hc203d742};
test_bias[3268:3268] = '{32'h42a55aad};
test_output[3268:3268] = '{32'hc59ecfe1};
test_input[26152:26159] = '{32'h40c1a5e8, 32'h41db3480, 32'hc050a166, 32'hc21eaacf, 32'hc26dca2a, 32'h42aac88e, 32'hc216ef4a, 32'hc2587d01};
test_weights[26152:26159] = '{32'h42b64bd4, 32'h42c29903, 32'h42c6e6a7, 32'hc1c12a84, 32'h4247af71, 32'hc280a3f0, 32'h42c0922f, 32'hc0eaac6e};
test_bias[3269:3269] = '{32'h42158885};
test_output[3269:3269] = '{32'hc5f3fe62};
test_input[26160:26167] = '{32'h4182433a, 32'hc2160e89, 32'h422096a0, 32'h42ae182a, 32'hc1aca794, 32'h4254d883, 32'hc291e397, 32'h42121e29};
test_weights[26160:26167] = '{32'hc0bbdc7d, 32'hc224554d, 32'hc28a911b, 32'hc2c055ae, 32'h4112bc08, 32'hc2c6d332, 32'h420ca693, 32'hc0ffe648};
test_bias[3270:3270] = '{32'hc2a5fafc};
test_output[3270:3270] = '{32'hc68dadb4};
test_input[26168:26175] = '{32'h41e17f4e, 32'h4255e3d6, 32'hc1be34c9, 32'hc00cbda6, 32'h3f633c2a, 32'hc2c3a6dd, 32'h429dbdcb, 32'hc28670d0};
test_weights[26168:26175] = '{32'hc1f7fdf5, 32'hc1cb058d, 32'hc21b8baf, 32'h42a095cc, 32'hc2598fda, 32'hc1845b10, 32'hc11b86b1, 32'h4259a6e9};
test_bias[3271:3271] = '{32'hc1ad7fa2};
test_output[3271:3271] = '{32'hc58834cf};
test_input[26176:26183] = '{32'hc27949dc, 32'hc18ca231, 32'hc2c03226, 32'hc29c8d78, 32'hc28c2261, 32'h4292d997, 32'hc2ba8b49, 32'hc2a61757};
test_weights[26176:26183] = '{32'hc2c62385, 32'h420ec7cf, 32'h422f99c2, 32'hc228e0ae, 32'h3f08ba9d, 32'h42b4e485, 32'h410947b7, 32'hc214f4d0};
test_bias[3272:3272] = '{32'hc1af9635};
test_output[3272:3272] = '{32'h46530acf};
test_input[26184:26191] = '{32'hc2a51c36, 32'hc2b4b7de, 32'hc25a0bc3, 32'h42b6578b, 32'h42b5c6da, 32'h42835450, 32'hc2487571, 32'h42821134};
test_weights[26184:26191] = '{32'h42976a47, 32'h42b941c8, 32'hc1356f61, 32'h425ac5c5, 32'h41f2f5b7, 32'hc26944b1, 32'hc1f5b8d7, 32'hc2756339};
test_bias[3273:3273] = '{32'hc2556cf2};
test_output[3273:3273] = '{32'hc644b04f};
test_input[26192:26199] = '{32'hc226b684, 32'h3f412cb8, 32'h41d5332c, 32'hc2ac4517, 32'hc2b504af, 32'h423c060f, 32'h42c0d7b1, 32'h424bfa34};
test_weights[26192:26199] = '{32'hc21b6f10, 32'hc1d97a15, 32'h4277b1f3, 32'hc2abaae2, 32'h4286e147, 32'hc1b46adb, 32'hc25cce85, 32'hc26545dd};
test_bias[3274:3274] = '{32'hc02089b4};
test_output[3274:3274] = '{32'hc5950baf};
test_input[26200:26207] = '{32'h422cc30f, 32'h429da0d2, 32'h42ab6233, 32'h4288dc90, 32'hc29ff55b, 32'hc17b32ff, 32'h42a858e8, 32'hc2aa51d7};
test_weights[26200:26207] = '{32'h42077816, 32'h41c10778, 32'hc2518450, 32'hc2a36e04, 32'h423df64d, 32'hc1adc68e, 32'h4004f138, 32'h41973266};
test_bias[3275:3275] = '{32'hc2201d05};
test_output[3275:3275] = '{32'hc635ff00};
test_input[26208:26215] = '{32'hc2749ec1, 32'h4240bb88, 32'h422d204c, 32'h42b517d0, 32'hc20e9544, 32'hc20d49d8, 32'hc28e5839, 32'hc2a96bd2};
test_weights[26208:26215] = '{32'h42879298, 32'h4216e47f, 32'hc2167454, 32'hc2116399, 32'h42989c3e, 32'h41efb081, 32'hc0d26107, 32'h429f9c1e};
test_bias[3276:3276] = '{32'hc2b3dc76};
test_output[3276:3276] = '{32'hc687ff12};
test_input[26216:26223] = '{32'h41f42742, 32'h423240a7, 32'h42af4762, 32'h4100c403, 32'h42121413, 32'hc2c515ea, 32'h412f279e, 32'hc07fc92c};
test_weights[26216:26223] = '{32'hc1d22f78, 32'hc28183aa, 32'h4291b761, 32'h42a81936, 32'h42c3d253, 32'hc12b8c7d, 32'hbdc03d12, 32'hc1fc70f4};
test_bias[3277:3277] = '{32'hc25affae};
test_output[3277:3277] = '{32'h45fc64d1};
test_input[26224:26231] = '{32'hc2a4d2f5, 32'hc198518f, 32'hc2ad406f, 32'hc2bc40ce, 32'h427eaece, 32'hc2b95276, 32'hc2b99921, 32'hc2a201c6};
test_weights[26224:26231] = '{32'hc1d010cf, 32'hc1ff969f, 32'h41a8cfc1, 32'h4244d448, 32'h41cfaf9b, 32'h429b6853, 32'hc28c7cf0, 32'hc29f4a8b};
test_bias[3278:3278] = '{32'hc2ae4999};
test_output[3278:3278] = '{32'h4562bdeb};
test_input[26232:26239] = '{32'hc2975c09, 32'h41ddf394, 32'h427e9426, 32'h42a5eab7, 32'hc0273636, 32'h42628d80, 32'h422bb5db, 32'h429c7b4a};
test_weights[26232:26239] = '{32'hc197662f, 32'h419d2e97, 32'hc27ddd80, 32'hc1f666a4, 32'hc20c9fb8, 32'hc26c24f4, 32'hc2982eff, 32'hc1a557c1};
test_bias[3279:3279] = '{32'hc28396f6};
test_output[3279:3279] = '{32'hc64848ed};
test_input[26240:26247] = '{32'h429623b7, 32'hc287c38d, 32'h4288d3a2, 32'hc2970efa, 32'h42c5b253, 32'h40d6f63c, 32'hc201c779, 32'hc2089bd5};
test_weights[26240:26247] = '{32'hc21676d2, 32'h42079459, 32'hc227e392, 32'hc255fdfb, 32'h42b483a7, 32'hc2a4b55d, 32'h42c082c7, 32'h41c4047a};
test_bias[3280:3280] = '{32'hc2b4c3d6};
test_output[3280:3280] = '{32'h43b57314};
test_input[26248:26255] = '{32'h424893cd, 32'hc23dbbd3, 32'h4052ded9, 32'h4254b4a2, 32'h42c44415, 32'h412fe92f, 32'h425200de, 32'h41b354b7};
test_weights[26248:26255] = '{32'hc26173c3, 32'h428f0147, 32'hc1638696, 32'hc25d57a8, 32'h4298ada8, 32'h42c0890b, 32'h42c617f3, 32'hc2802c11};
test_bias[3281:3281] = '{32'h428358d4};
test_output[3281:3281] = '{32'h45463a30};
test_input[26256:26263] = '{32'hc2c2c0f2, 32'hbfee4846, 32'h42a8f127, 32'hc2735920, 32'h429dcc0a, 32'h415b850a, 32'h415cd0f6, 32'hc0b64b1f};
test_weights[26256:26263] = '{32'hc24f37cd, 32'h41c86873, 32'hc2b0ec80, 32'h4291159a, 32'h426f658c, 32'h41269a65, 32'hc141c4fd, 32'hc2185a30};
test_bias[3282:3282] = '{32'h4244edc8};
test_output[3282:3282] = '{32'hc4f07b57};
test_input[26264:26271] = '{32'h42687a0a, 32'h421bea40, 32'h42b5faf0, 32'hc23e016b, 32'h42b12fcd, 32'hc2782cd5, 32'hc2c3593b, 32'h42c3ce84};
test_weights[26264:26271] = '{32'h420530ac, 32'h42b6ea9e, 32'h407141da, 32'hc14b5faa, 32'h42119522, 32'hc2a2e0fc, 32'hbecefadc, 32'hc2bd9bc0};
test_bias[3283:3283] = '{32'hc288d7d4};
test_output[3283:3283] = '{32'h45a92c98};
test_input[26272:26279] = '{32'hc25ca20b, 32'h417f318a, 32'hc1c70162, 32'hc2b20467, 32'h4154b4df, 32'hc2b55355, 32'hc19dd65b, 32'h40d37bb5};
test_weights[26272:26279] = '{32'h42bf6cbe, 32'h429d7d91, 32'h42009a20, 32'h3ed4c3fa, 32'h42beb590, 32'h420c81b8, 32'h424e128e, 32'hc1e77ca8};
test_bias[3284:3284] = '{32'hc0d9125b};
test_output[3284:3284] = '{32'hc5f9bccd};
test_input[26280:26287] = '{32'hc295ea13, 32'h428fc3d1, 32'hc205119d, 32'hc26dc9b3, 32'hc2386d6d, 32'hc26259be, 32'h42b5751c, 32'h426508ec};
test_weights[26280:26287] = '{32'h4280bffe, 32'h429aee1b, 32'h421708e6, 32'h42471d04, 32'hc2c63342, 32'h423084ff, 32'h42463abb, 32'hc288a7a4};
test_bias[3285:3285] = '{32'h41c0e3c0};
test_output[3285:3285] = '{32'hc4460ffe};
test_input[26288:26295] = '{32'h410462bc, 32'hc0ca97fe, 32'h4162e3bb, 32'h3f7ad119, 32'hc296d20b, 32'hc2960d20, 32'h42a1e740, 32'hc27bcd7f};
test_weights[26288:26295] = '{32'hc278de3a, 32'hc2951f08, 32'h428c9b6c, 32'hc264c21c, 32'hc267a6e9, 32'hc28a5b44, 32'hc1578c66, 32'h4293a3f5};
test_bias[3286:3286] = '{32'h42a1e48f};
test_output[3286:3286] = '{32'h4595f72f};
test_input[26296:26303] = '{32'hc124c681, 32'hc21d381e, 32'h4209ecda, 32'hc2c463c2, 32'h416a6be0, 32'h42b3e4d9, 32'hc28a50db, 32'hc0b895ad};
test_weights[26296:26303] = '{32'hc2bb9627, 32'h4288cebc, 32'h42b1bb7c, 32'h4294ce9e, 32'h41165a93, 32'h4298eb1a, 32'h4238fb47, 32'h41ae374c};
test_bias[3287:3287] = '{32'hc10da04d};
test_output[3287:3287] = '{32'hc50ea3e8};
test_input[26304:26311] = '{32'hc246cc3f, 32'hc2c02202, 32'hc05b9df5, 32'hc151e1d9, 32'hc251c764, 32'h42c124d5, 32'hc2be24d2, 32'h427b91e8};
test_weights[26304:26311] = '{32'h411b344c, 32'h428b17ba, 32'hc2ba5483, 32'h3fde23a8, 32'h42aa1289, 32'hc14467e8, 32'h428aeb44, 32'h42021eb5};
test_bias[3288:3288] = '{32'hc2ac5212};
test_output[3288:3288] = '{32'hc686069d};
test_input[26312:26319] = '{32'hc2c16de5, 32'h42835616, 32'hc28ce409, 32'hc200fb69, 32'hc1733efb, 32'hc1c0df11, 32'hc2c3901f, 32'hc2ab9c53};
test_weights[26312:26319] = '{32'hc283a8b4, 32'hc235acb3, 32'hc28b96e8, 32'hc19b7daa, 32'h41c3aedf, 32'hc200f52d, 32'h42862a67, 32'h41f9c3d7};
test_bias[3289:3289] = '{32'h4204a5c6};
test_output[3289:3289] = '{32'h42ff8986};
test_input[26320:26327] = '{32'h42b153da, 32'h429cfb47, 32'hc2b3d924, 32'hc2ba0140, 32'hc2b2ce8e, 32'h41a74678, 32'h421b525e, 32'h42c596a0};
test_weights[26320:26327] = '{32'hc2a86f47, 32'h427b5688, 32'hc27d6d92, 32'hc1ce67b0, 32'hc1b42c77, 32'hc2c7393d, 32'h429f994e, 32'hc18c239d};
test_bias[3290:3290] = '{32'hc26bc914};
test_output[3290:3290] = '{32'h45d48c2f};
test_input[26328:26335] = '{32'hc1682b3a, 32'h416759f1, 32'hc1dc7a1f, 32'h423605fb, 32'hc069d63d, 32'h42ac6225, 32'hc195c646, 32'h4083b651};
test_weights[26328:26335] = '{32'h42932a61, 32'h419fcba9, 32'hc2490c6b, 32'h424c8963, 32'h4229e10f, 32'h41e90040, 32'h41e085bd, 32'hc0e49a42};
test_bias[3291:3291] = '{32'h42a4eed4};
test_output[3291:3291] = '{32'h45968005};
test_input[26336:26343] = '{32'hc1cfac1e, 32'hc25fc1d6, 32'h41785d06, 32'h425ccb11, 32'h3f66d492, 32'hc20eb623, 32'hc200f6c3, 32'hc2c00230};
test_weights[26336:26343] = '{32'hc28afdc1, 32'hc25ccde7, 32'hc0da20f4, 32'h41e22eef, 32'h42810908, 32'hc1c23ced, 32'hc160a82b, 32'h428e3555};
test_bias[3292:3292] = '{32'hc1803102};
test_output[3292:3292] = '{32'h445c6326};
test_input[26344:26351] = '{32'h42ac89fb, 32'hc290485b, 32'hc1e4795e, 32'hc2866a9e, 32'h42aaa95e, 32'h41f00d91, 32'hc286b66d, 32'hc1ebeaf9};
test_weights[26344:26351] = '{32'hc25c984a, 32'hc2bf1274, 32'hc22cbacf, 32'h429b0c11, 32'h410cf0a5, 32'hbe4f4e26, 32'hc1a33e6e, 32'h4186b954};
test_bias[3293:3293] = '{32'h41f06710};
test_output[3293:3293] = '{32'hc33d1206};
test_input[26352:26359] = '{32'h4282cc21, 32'hc268c585, 32'h4217334a, 32'hc1e5304a, 32'h41037af0, 32'h42229804, 32'hc24db67c, 32'h427ee202};
test_weights[26352:26359] = '{32'hc212227c, 32'hc2bf8f8d, 32'h41e32a19, 32'hc2c41d57, 32'h41908d92, 32'hc17cc084, 32'hc26d9a35, 32'hc1add2b2};
test_bias[3294:3294] = '{32'hc18d7ae7};
test_output[3294:3294] = '{32'h46008842};
test_input[26360:26367] = '{32'h42727aae, 32'h4216a22d, 32'hc289c878, 32'h42550941, 32'h417ae50f, 32'h414ab323, 32'hc2b6d7b4, 32'hc030f527};
test_weights[26360:26367] = '{32'h419c8012, 32'hc2811e34, 32'hc26bcff3, 32'h4293a29c, 32'h42b00ff6, 32'hc222c580, 32'h4091dfc3, 32'h4291b484};
test_bias[3295:3295] = '{32'h42c5a6b9};
test_output[3295:3295] = '{32'h45dda84b};
test_input[26368:26375] = '{32'h42ae6981, 32'h428de4af, 32'hc291f3c7, 32'hc2a457bd, 32'h42bbb289, 32'hc22531f9, 32'h41bfe445, 32'hc2636eb1};
test_weights[26368:26375] = '{32'hc2584e98, 32'hc243f710, 32'h42ade3f5, 32'h42a228e0, 32'hc213521a, 32'hc26613b6, 32'hc292853f, 32'h403c4840};
test_bias[3296:3296] = '{32'hc20515b4};
test_output[3296:3296] = '{32'hc6bd5b7a};
test_input[26376:26383] = '{32'hc1528ee8, 32'hc282062c, 32'hc2916f27, 32'h426a5fe3, 32'hc2957035, 32'hc158e2bd, 32'h41f1c8aa, 32'hc1791e68};
test_weights[26376:26383] = '{32'hc2c63418, 32'hc26ee201, 32'hc29633ae, 32'h423deb02, 32'hc0801cfb, 32'hc2a86588, 32'hc2c4596f, 32'h428c1d22};
test_bias[3297:3297] = '{32'h4281f747};
test_output[3297:3297] = '{32'h4629f59d};
test_input[26384:26391] = '{32'hc09cc329, 32'hc2b0a32f, 32'h41f44dfa, 32'hc2a6e841, 32'hc127f8a2, 32'h40c8843c, 32'h4239f62e, 32'hc22bbd10};
test_weights[26384:26391] = '{32'hc2400ada, 32'hc1c20d03, 32'hc09807f0, 32'h422b91e7, 32'hc1f16577, 32'hc272d134, 32'hc1b21620, 32'h42b80dac};
test_bias[3298:3298] = '{32'hc240683b};
test_output[3298:3298] = '{32'hc5c96713};
test_input[26392:26399] = '{32'h4243bc59, 32'h4255803a, 32'hc29b06fa, 32'hc29e9f57, 32'h42a98efb, 32'h42964c2c, 32'h419f7971, 32'hc299afa5};
test_weights[26392:26399] = '{32'hc29701a1, 32'h4226f5c2, 32'hc2bafb5b, 32'h42a3d7ab, 32'h42253eb8, 32'h42c4638e, 32'hc22357a2, 32'h42a20d6c};
test_bias[3299:3299] = '{32'h4107ba3e};
test_output[3299:3299] = '{32'h4543c71b};
test_input[26400:26407] = '{32'hbfe7e03d, 32'h42b5c665, 32'h42050143, 32'hc261870b, 32'hc25d8aa5, 32'hc22a2455, 32'h421fd5aa, 32'hc23e5a23};
test_weights[26400:26407] = '{32'hc289b860, 32'h428f7e0a, 32'hc2a65f7f, 32'hc0acf25a, 32'h42545efc, 32'h41948d91, 32'hc210fb79, 32'hc1978174};
test_bias[3300:3300] = '{32'h425e1d8e};
test_output[3300:3300] = '{32'hc216f184};
test_input[26408:26415] = '{32'h428b2545, 32'hc2635c25, 32'h40cf9632, 32'hc235cf5f, 32'hc2b8de14, 32'h42550859, 32'h42c0464f, 32'hc2719445};
test_weights[26408:26415] = '{32'hc2454f05, 32'h42762739, 32'h41223a2b, 32'hc29ff6c4, 32'h42587648, 32'h4287a945, 32'h4146eee8, 32'hc1957469};
test_bias[3301:3301] = '{32'h42737868};
test_output[3301:3301] = '{32'hc50b99df};
test_input[26416:26423] = '{32'hc1ab48dd, 32'hc298a702, 32'hc2bf3ffe, 32'h417c993e, 32'h415b9640, 32'hc0e78ffc, 32'h421cdfad, 32'h41409c49};
test_weights[26416:26423] = '{32'h428a5682, 32'h421413f8, 32'hc270d1b3, 32'h422e522d, 32'h427710cb, 32'h427a9f6c, 32'h425fc688, 32'h42a10daa};
test_bias[3302:3302] = '{32'hc29a03ae};
test_output[3302:3302] = '{32'h45af9a79};
test_input[26424:26431] = '{32'hc1c0840b, 32'h42ad3385, 32'h4288fca3, 32'h42a50731, 32'hc2a768db, 32'hc2c3fe2b, 32'h428a12b7, 32'h42439911};
test_weights[26424:26431] = '{32'hc23818ee, 32'hc2b8628a, 32'hc26ee3b5, 32'h41d27ca4, 32'h4219c9cc, 32'hc200a7c3, 32'h4147b566, 32'hc1aa5207};
test_bias[3303:3303] = '{32'h42c6e7ae};
test_output[3303:3303] = '{32'hc60bb886};
test_input[26432:26439] = '{32'h42a899db, 32'h4275292a, 32'h4227a231, 32'h425a6f28, 32'hc272db9a, 32'h422e7acb, 32'h42c76ed0, 32'h420a41ec};
test_weights[26432:26439] = '{32'h4287fa7c, 32'h419fa1c5, 32'h40dc7684, 32'hc12bb26c, 32'hc25a5232, 32'hc225a920, 32'hc21e0d6e, 32'hc0192f66};
test_bias[3304:3304] = '{32'hc2bd64b0};
test_output[3304:3304] = '{32'h457cefaf};
test_input[26440:26447] = '{32'hc2b8e560, 32'h412a106f, 32'hc2a8f392, 32'h42b3cfdd, 32'hc1e24930, 32'hc25b47eb, 32'hc2a8eee2, 32'hc12a2520};
test_weights[26440:26447] = '{32'hc1537331, 32'h4016e4a5, 32'h40db70be, 32'h42bfa491, 32'hc28b05f4, 32'hc2bff9da, 32'h40bfb8e2, 32'hc1c0896e};
test_bias[3305:3305] = '{32'h42a8c09d};
test_output[3305:3305] = '{32'h467f63d4};
test_input[26448:26455] = '{32'hc16a433d, 32'h426e2ac6, 32'hc215a8f8, 32'hc26bc6a0, 32'h4249b833, 32'h41fad67a, 32'h4287c0dc, 32'hc261f214};
test_weights[26448:26455] = '{32'hc244a6ee, 32'hc1cbd372, 32'hc2858e56, 32'hc29043e7, 32'hc21d3e48, 32'hc2a42d39, 32'hc2911376, 32'hc2779751};
test_bias[3306:3306] = '{32'hc290809e};
test_output[3306:3306] = '{32'hc2cd73ab};
test_input[26456:26463] = '{32'hc224f14c, 32'hc24f1ef1, 32'h41dda805, 32'h42b039bc, 32'hc1119f3f, 32'hc2387233, 32'hc1a9c419, 32'hc2562dd1};
test_weights[26456:26463] = '{32'h4289878d, 32'h41264859, 32'hc2c6e093, 32'hc227e430, 32'h41c8787a, 32'h425d225f, 32'h424342c2, 32'h427e7555};
test_bias[3307:3307] = '{32'hc206e9fc};
test_output[3307:3307] = '{32'hc68570a1};
test_input[26464:26471] = '{32'h42c1dad0, 32'h4178176d, 32'hc1eec271, 32'hc1d9ba84, 32'hc2984136, 32'h40153b71, 32'hc28d3a1d, 32'hc1485849};
test_weights[26464:26471] = '{32'h41b0fddf, 32'h428df235, 32'h425fd52a, 32'hc2a881f1, 32'hc10feca6, 32'h423254ea, 32'h429e6297, 32'h42b6ce56};
test_bias[3308:3308] = '{32'h41c23702};
test_output[3308:3308] = '{32'hc5007a85};
test_input[26472:26479] = '{32'hc2c3a840, 32'hc1741c89, 32'h427b7e5f, 32'h4291a113, 32'hc20124f1, 32'hc21a18c2, 32'hc223d5ea, 32'hc2af3ab1};
test_weights[26472:26479] = '{32'hc29ad098, 32'h4291fc49, 32'hc2923b05, 32'hc143a862, 32'h429bdf65, 32'hc27e6979, 32'h42a71876, 32'h422f18ad};
test_bias[3309:3309] = '{32'h4199349c};
test_output[3309:3309] = '{32'hc5c5e460};
test_input[26480:26487] = '{32'hc2c040be, 32'h42ba3b24, 32'hc0d5f36b, 32'hc1fabafb, 32'h4229d704, 32'h428f75a2, 32'h42b57cb2, 32'hc199944f};
test_weights[26480:26487] = '{32'h429ac80b, 32'h42b43471, 32'hc24b4253, 32'hc27b0b0a, 32'hc18ffb3c, 32'h42635c20, 32'h4285cf10, 32'h4131c102};
test_bias[3310:3310] = '{32'h418d0feb};
test_output[3310:3310] = '{32'h4642774d};
test_input[26488:26495] = '{32'hc216098c, 32'h42328c9d, 32'hc290d148, 32'h4242a032, 32'h4121ab31, 32'h4292d1d5, 32'hc26046da, 32'h429cc2f3};
test_weights[26488:26495] = '{32'hc2c37be6, 32'h422dbb87, 32'h425af243, 32'h42869f28, 32'h42c7c388, 32'hc1f0bf72, 32'h42c412ae, 32'hc2a8636f};
test_bias[3311:3311] = '{32'h41a31c82};
test_output[3311:3311] = '{32'hc6029b91};
test_input[26496:26503] = '{32'h428ba791, 32'hc24a93ec, 32'h4290cf55, 32'h42313193, 32'hc29312d1, 32'hc2c7555f, 32'h421dec71, 32'hc0100787};
test_weights[26496:26503] = '{32'hc2865455, 32'h4237d0cb, 32'hc2bea928, 32'hc15e8abb, 32'hc2aebc3c, 32'hc2aab2b6, 32'h4251abab, 32'hc2b2b723};
test_bias[3312:3312] = '{32'h42996a99};
test_output[3312:3312] = '{32'h452b6b8e};
test_input[26504:26511] = '{32'h42a87097, 32'h429e9b2b, 32'hc1266bee, 32'hc1b15e66, 32'hc2be7cd9, 32'h424d7837, 32'hc2875e9b, 32'h428dc3b7};
test_weights[26504:26511] = '{32'hc12d373b, 32'h42b042a5, 32'h42980a60, 32'hc29d51cc, 32'h42b62990, 32'h41c4c5dc, 32'hc2b3ae19, 32'h4285fbd0};
test_bias[3313:3313] = '{32'hc1a095bc};
test_output[3313:3313] = '{32'h4622f12a};
test_input[26512:26519] = '{32'h4170e68d, 32'hc2892739, 32'hc25fdf31, 32'hc153476e, 32'h426c52f0, 32'h426dc77d, 32'hc23e1de6, 32'h3e63c709};
test_weights[26512:26519] = '{32'h42a620bb, 32'hc251486c, 32'h41ac7fc3, 32'hc2b9a29f, 32'hc0dff651, 32'h42483ccf, 32'hc2688814, 32'h41a2dede};
test_bias[3314:3314] = '{32'h424269bb};
test_output[3314:3314] = '{32'h461fef80};
test_input[26520:26527] = '{32'h41a24b99, 32'h42b35c3a, 32'hc23f8d00, 32'hc1f4ffe6, 32'h4232e607, 32'h3fd885f0, 32'hc20781bd, 32'hc2c0bb0b};
test_weights[26520:26527] = '{32'h4201efaf, 32'h428077f0, 32'h423cc5e1, 32'h427b0fc3, 32'hc28f857b, 32'h42a7fb67, 32'h427786f8, 32'h42955a54};
test_bias[3315:3315] = '{32'hc24ab31b};
test_output[3315:3315] = '{32'hc61ef50b};
test_input[26528:26535] = '{32'hc285918e, 32'hc2247614, 32'hc10c472b, 32'hc0f4d79d, 32'hc0f88856, 32'h42055495, 32'hc281ae3f, 32'h41c784f3};
test_weights[26528:26535] = '{32'h429c4996, 32'hc2075102, 32'hc2a66792, 32'h423bbaae, 32'h42683380, 32'h4192e86b, 32'h40fe430a, 32'hc245c62f};
test_bias[3316:3316] = '{32'hc08d0d46};
test_output[3316:3316] = '{32'hc59dc7e3};
test_input[26536:26543] = '{32'h416d89c0, 32'h42016dc3, 32'hc26f8eb4, 32'hc288d2cb, 32'hc2559d12, 32'hc25df2be, 32'hc1b2a0c1, 32'h4276dd27};
test_weights[26536:26543] = '{32'hc28ae487, 32'h42945a4a, 32'hc28cec77, 32'hc2c68031, 32'hc21846d7, 32'h42afd0ed, 32'h42a22840, 32'hc2c73127};
test_bias[3317:3317] = '{32'h40448fc1};
test_output[3317:3317] = '{32'h44c587a6};
test_input[26544:26551] = '{32'h41fd00c2, 32'hc2122489, 32'h40c11ebf, 32'hc2b4654a, 32'h42824fe6, 32'h42a4286a, 32'hc22def08, 32'hc2bcec20};
test_weights[26544:26551] = '{32'h4084b0b6, 32'h4235a2e6, 32'hc1fd2571, 32'h421276e3, 32'h414ae721, 32'hc21a8dcd, 32'h42699c08, 32'hc19ad2d0};
test_bias[3318:3318] = '{32'hc1af0ad3};
test_output[3318:3318] = '{32'hc5fd202e};
test_input[26552:26559] = '{32'hc08e3276, 32'hc1eeedd8, 32'hc025ff84, 32'hc0bae3ca, 32'hc1a2d891, 32'h428d7703, 32'hc06ba3d4, 32'hc267e315};
test_weights[26552:26559] = '{32'h41060fd8, 32'hc2a761a7, 32'h42bea4d6, 32'h428ddff6, 32'hc2997c91, 32'hc0bee519, 32'h4237a18a, 32'h42ba33cd};
test_bias[3319:3319] = '{32'hc17bb2e9};
test_output[3319:3319] = '{32'hc525107e};
test_input[26560:26567] = '{32'hc2828271, 32'h423c8007, 32'h42924ed7, 32'h41ab6fc9, 32'hc287f895, 32'h424f3c52, 32'h4292e58f, 32'h42a55c40};
test_weights[26560:26567] = '{32'hc2c78c4f, 32'hc234c6ae, 32'hc202c1fe, 32'h4290e868, 32'hc284ec2a, 32'hc2c2664a, 32'h418edcc0, 32'hc24b63c0};
test_bias[3320:3320] = '{32'hc2bf6bc2};
test_output[3320:3320] = '{32'h4212bf30};
test_input[26568:26575] = '{32'hc211372e, 32'h4212ee8c, 32'hc2817827, 32'h42b219ef, 32'hc1e16b6d, 32'hc0a14bd6, 32'hc128c073, 32'hbfef2721};
test_weights[26568:26575] = '{32'h40c18f63, 32'h3f281bab, 32'h42b36096, 32'hc2adc78c, 32'h421e2bea, 32'hc2b35c6d, 32'hc18ee58d, 32'hc2adc40e};
test_bias[3321:3321] = '{32'h41fa2a99};
test_output[3321:3321] = '{32'hc65b0cdc};
test_input[26576:26583] = '{32'h42adb707, 32'hc26512be, 32'h429bb8cc, 32'hc1142770, 32'hc2a7be3b, 32'hc28a4c7a, 32'hc27f32d9, 32'hc052eeb0};
test_weights[26576:26583] = '{32'h4087782b, 32'h4113141a, 32'h42b10886, 32'h42827e40, 32'h423a7d3f, 32'hc06f7d21, 32'hc202e964, 32'h422fd367};
test_bias[3322:3322] = '{32'h427530de};
test_output[3322:3322] = '{32'h458c1039};
test_input[26584:26591] = '{32'h4239e4aa, 32'hc22f727b, 32'h425f652c, 32'hc2ad7d51, 32'h41905a1f, 32'hc1fb54d3, 32'hc25a8daa, 32'hc1ff32a1};
test_weights[26584:26591] = '{32'hc1760732, 32'h4240193f, 32'h42a1fcbe, 32'hc212ff3c, 32'hc226721f, 32'hc2c06c83, 32'h42a81d83, 32'h429adae5};
test_bias[3323:3323] = '{32'h41650b62};
test_output[3323:3323] = '{32'h42e324d1};
test_input[26592:26599] = '{32'hc2531d3c, 32'hc27e8b91, 32'h42483e37, 32'hc2acf436, 32'h40546bb4, 32'hc2b8e4ec, 32'h42106e8f, 32'hc2b86795};
test_weights[26592:26599] = '{32'h421d7808, 32'hc2b85ce8, 32'hc1dfa7de, 32'h41859caa, 32'h42b12b55, 32'h42803689, 32'h4294a9b9, 32'hc29bea23};
test_bias[3324:3324] = '{32'hc1a7e373};
test_output[3324:3324] = '{32'h45a156fa};
test_input[26600:26607] = '{32'h417d3c27, 32'h4138500e, 32'h403dc996, 32'hc29c7513, 32'h42ae6b26, 32'h421b1aaa, 32'h429d1bcb, 32'h424f8531};
test_weights[26600:26607] = '{32'hc2a619c5, 32'hc12bf51e, 32'h4216bdbf, 32'h3f8ed388, 32'h422a701e, 32'h42129429, 32'h42455c08, 32'hc1ced75b};
test_bias[3325:3325] = '{32'hc1b05c36};
test_output[3325:3325] = '{32'h45c2dc3e};
test_input[26608:26615] = '{32'h4228d46e, 32'hc1ba8d24, 32'hc1f9c535, 32'hc2bb10fb, 32'h42239e42, 32'hc1e03638, 32'h42c51e1a, 32'hc22fc029};
test_weights[26608:26615] = '{32'h427841ae, 32'hc2758869, 32'hc28c8b14, 32'hc261f572, 32'hc0453b28, 32'h428c6b47, 32'h41d48a06, 32'h428e7c78};
test_bias[3326:3326] = '{32'h41b857c0};
test_output[3326:3326] = '{32'h460bc82e};
test_input[26616:26623] = '{32'h419de333, 32'hc01ecd9c, 32'h422ccdf8, 32'h429d0133, 32'h4132104a, 32'h4096c1b4, 32'hc25a34c1, 32'h420bbf7e};
test_weights[26616:26623] = '{32'hc25fd3bf, 32'hbec1c738, 32'hc206c580, 32'h3fdfe277, 32'h42ae25ae, 32'h42a135e5, 32'h423cc755, 32'h423b0973};
test_bias[3327:3327] = '{32'h3f471a30};
test_output[3327:3327] = '{32'hc4fba11d};
test_input[26624:26631] = '{32'h41d03e9a, 32'h41984c84, 32'h41c5bb29, 32'hc2c1cb25, 32'h41757bb2, 32'hc1d6e745, 32'hc1bbd075, 32'hc2823022};
test_weights[26624:26631] = '{32'hc2c72cb4, 32'hc1d4d124, 32'hc28be46e, 32'hc29bb9d9, 32'h4295cf52, 32'h41b29396, 32'hc123f649, 32'h420c5054};
test_bias[3328:3328] = '{32'hc229e7ab};
test_output[3328:3328] = '{32'h4493ad8d};
test_input[26632:26639] = '{32'hc2600f1a, 32'h4272e941, 32'hbee0c8ce, 32'h42316643, 32'h3fad4df9, 32'h4258e64a, 32'hc2428dcf, 32'h3eedd571};
test_weights[26632:26639] = '{32'h423944b5, 32'hc2276d5c, 32'hc24cab44, 32'hc2a48eb3, 32'h424fda86, 32'hc2789b6c, 32'h41b18657, 32'hc1d1b4d0};
test_bias[3329:3329] = '{32'h40a2056e};
test_output[3329:3329] = '{32'hc64d7495};
test_input[26640:26647] = '{32'h408b26c9, 32'hc14b0417, 32'hc1ef8dca, 32'hc1d4e4c2, 32'hc28e3081, 32'h41e0f17f, 32'h4193ca8a, 32'hc27daae9};
test_weights[26640:26647] = '{32'hc190d12e, 32'h41cfbc91, 32'hc261325e, 32'hc1bfdd60, 32'h41f9173a, 32'hc1cf06b3, 32'hc28b42a3, 32'h3fb24cd2};
test_bias[3330:3330] = '{32'h425ddb5c};
test_output[3330:3330] = '{32'hc51289ec};
test_input[26648:26655] = '{32'hc1b2c2af, 32'hc295cf44, 32'h41b15216, 32'hc1040dd3, 32'h405f217c, 32'h40afb03c, 32'hc29d4fd1, 32'h40f635d4};
test_weights[26648:26655] = '{32'hc25cd7da, 32'h42b2bb39, 32'hc186ec04, 32'hc20fc770, 32'h422778b4, 32'h42726266, 32'h41220ce1, 32'h40a0594a};
test_bias[3331:3331] = '{32'h427efce2};
test_output[3331:3331] = '{32'hc5b3c883};
test_input[26656:26663] = '{32'h42bd972e, 32'h42492eb0, 32'hc21e72bf, 32'h41b5ad6d, 32'hc270e298, 32'h425143ea, 32'h4162dbcc, 32'hc0b820eb};
test_weights[26656:26663] = '{32'hc23313cd, 32'h41c791d0, 32'h3f51b9a7, 32'h42b38d2f, 32'h42b36ce8, 32'h429b1134, 32'hc2aa7160, 32'h4282fceb};
test_bias[3332:3332] = '{32'hc216b64b};
test_output[3332:3332] = '{32'hc57701c1};
test_input[26664:26671] = '{32'h429b0afa, 32'hc2160e68, 32'h42a3df5b, 32'hc2a4d8a1, 32'h42bb8617, 32'hc2a86561, 32'h41486609, 32'h42bde85f};
test_weights[26664:26671] = '{32'hc286434a, 32'hc1ad0934, 32'h42815ccd, 32'h41eddddb, 32'h41a006e2, 32'h4229e952, 32'hc29be45f, 32'h41196dde};
test_bias[3333:3333] = '{32'h4258c180};
test_output[3333:3333] = '{32'hc54b838a};
test_input[26672:26679] = '{32'hc22c7b22, 32'h41f7affa, 32'h4218faf6, 32'hc12ede7f, 32'h4292affc, 32'hc2a2a447, 32'h4288e7b5, 32'hc2a8c642};
test_weights[26672:26679] = '{32'hc2a585e1, 32'hc2bfa499, 32'h4221f9ff, 32'hc2b420eb, 32'h40de1d02, 32'h42aff50e, 32'hc2010ba5, 32'hc2c76497};
test_bias[3334:3334] = '{32'hc134de76};
test_output[3334:3334] = '{32'h4527b086};
test_input[26680:26687] = '{32'hc192d1c5, 32'hc2bb9511, 32'h424a5e12, 32'h4250a84c, 32'hc159fe95, 32'hc2c1217c, 32'h40f4c4f5, 32'hc242d6e3};
test_weights[26680:26687] = '{32'h42867cfd, 32'hc2adaa19, 32'hc29fa71d, 32'h422aca64, 32'h42873af6, 32'hc0f1cf55, 32'hc17ec837, 32'hc2a59acd};
test_bias[3335:3335] = '{32'h4297b274};
test_output[3335:3335] = '{32'h460afa23};
test_input[26688:26695] = '{32'h41bd9088, 32'hc22c1807, 32'h426928b4, 32'hc188e910, 32'h4125c334, 32'h42bfae43, 32'hc01b1f0d, 32'h42211a23};
test_weights[26688:26695] = '{32'hc215b3eb, 32'h42841a54, 32'hbfdf0dc0, 32'hc2a67fdc, 32'h428683e6, 32'hc2a575fc, 32'h42520674, 32'hc27dbfea};
test_bias[3336:3336] = '{32'hc23b07cd};
test_output[3336:3336] = '{32'hc6413a36};
test_input[26696:26703] = '{32'h41331e64, 32'h41a3bca4, 32'hc260b557, 32'hc217465f, 32'hc1fcb10b, 32'hc036a357, 32'h4234c829, 32'h415ead47};
test_weights[26696:26703] = '{32'h4269518d, 32'h42a640f1, 32'hc228fafc, 32'hc294ba97, 32'hc1946697, 32'hc2a596fa, 32'hc2c49da2, 32'h42b8eebf};
test_bias[3337:3337] = '{32'h4149d1c9};
test_output[3337:3337] = '{32'h45a31488};
test_input[26704:26711] = '{32'hc2ab1c21, 32'h42c3c02b, 32'hc11d1fe8, 32'hc138f76c, 32'h422c47ee, 32'h42a58f45, 32'h42aa7adf, 32'h422f5633};
test_weights[26704:26711] = '{32'h42b65151, 32'h42435211, 32'h42a086e4, 32'h423484e9, 32'hc2a851d3, 32'hc2949437, 32'h40ad8168, 32'hc29b36af};
test_bias[3338:3338] = '{32'hc0935ef5};
test_output[3338:3338] = '{32'hc68530ee};
test_input[26712:26719] = '{32'hc2169738, 32'h4202740a, 32'h428abcc1, 32'h42a008c6, 32'h42a9a452, 32'hc283fe2b, 32'hc0aa0357, 32'hc12d6c94};
test_weights[26712:26719] = '{32'h41c05c95, 32'h419ce77c, 32'h41d5ceb8, 32'h4277ffa4, 32'h4222ebcd, 32'hc2bfefad, 32'h428fa1cb, 32'h428fdda9};
test_bias[3339:3339] = '{32'h424996aa};
test_output[3339:3339] = '{32'h466deb7d};
test_input[26720:26727] = '{32'hc27a3697, 32'hc11aa442, 32'hc225d042, 32'h429401a0, 32'hc16097c4, 32'h42a04444, 32'hc2175118, 32'h42c50f86};
test_weights[26720:26727] = '{32'h422cd6ae, 32'hc2a18cd5, 32'h42a86a3a, 32'h429a0ce0, 32'h423ebc45, 32'hc2c4943d, 32'hc2794784, 32'h42a43f66};
test_bias[3340:3340] = '{32'hc292a665};
test_output[3340:3340] = '{32'h450457a1};
test_input[26728:26735] = '{32'h41d715f3, 32'h41408bae, 32'hc25d46ee, 32'h41d9a6fa, 32'hc18d7d33, 32'hc29f9da7, 32'h420bc200, 32'hc284da1a};
test_weights[26728:26735] = '{32'h42ba3ca4, 32'h421b86db, 32'h42ac3e35, 32'hc29f1448, 32'hc14b1e88, 32'h40b7f9ba, 32'hc1c2e67d, 32'hc0d67d83};
test_bias[3341:3341] = '{32'h423a4ae4};
test_output[3341:3341] = '{32'hc58e3360};
test_input[26736:26743] = '{32'hc2253ea5, 32'hc23e350a, 32'hc29978de, 32'hc1dd2b67, 32'hc2ac197e, 32'hc20824f8, 32'hc200da62, 32'hc2be060e};
test_weights[26736:26743] = '{32'hc22acc3b, 32'hc2c0c46e, 32'hc2a19eec, 32'h420ab9e5, 32'h42a51531, 32'h42663e7b, 32'h421b8399, 32'hc288dc04};
test_bias[3342:3342] = '{32'h42a1304b};
test_output[3342:3342] = '{32'h45f58b85};
test_input[26744:26751] = '{32'hc20270ed, 32'h41a44c51, 32'hc189f49f, 32'hc25ef75b, 32'hc10e7eb4, 32'hc20208d4, 32'hc18c6fec, 32'h4203bedd};
test_weights[26744:26751] = '{32'h4239675e, 32'h4296746e, 32'h426b6fbe, 32'hc20be265, 32'hc24f03f7, 32'h42680adb, 32'h4299b55f, 32'hc2be3b5f};
test_bias[3343:3343] = '{32'h4240df4a};
test_output[3343:3343] = '{32'hc598d6b3};
test_input[26752:26759] = '{32'h428726f1, 32'hc29905f5, 32'hc2b94a5c, 32'hc2c09f46, 32'hc1eb3e9a, 32'hc232a1b5, 32'hc28eab30, 32'h4246d8b9};
test_weights[26752:26759] = '{32'h42c5b519, 32'hc26f4280, 32'hc15bdc60, 32'h42a14ca5, 32'hc1ec36fe, 32'h426a58ec, 32'hc2acc309, 32'h42a5ecee};
test_bias[3344:3344] = '{32'h42486159};
test_output[3344:3344] = '{32'h465099a8};
test_input[26760:26767] = '{32'hc29a53b7, 32'h41c01960, 32'h429d0b2a, 32'hc0cd85ba, 32'h4203e257, 32'hc22bcb90, 32'h42bbec46, 32'h42801554};
test_weights[26760:26767] = '{32'hc2162abf, 32'h4203bf4a, 32'h428a02f3, 32'h42ba1a13, 32'h4269c2a5, 32'hc2551e70, 32'hc2c2f1d0, 32'h41a2dc52};
test_bias[3345:3345] = '{32'h41caaede};
test_output[3345:3345] = '{32'h4598f10f};
test_input[26768:26775] = '{32'h41b2cf97, 32'hc2b9b855, 32'h42855dab, 32'h42179bf7, 32'h42b1f740, 32'h42121722, 32'hc2175c26, 32'hc1f5d933};
test_weights[26768:26775] = '{32'h42b37fe9, 32'h4292cb78, 32'hc2ac18eb, 32'h4267c1fb, 32'hc289e760, 32'hc2bfbfb7, 32'h420389c4, 32'hc167766f};
test_bias[3346:3346] = '{32'h4212cb26};
test_output[3346:3346] = '{32'hc6927f9a};
test_input[26776:26783] = '{32'hc1a9a72c, 32'h40d8ef3a, 32'h42b48389, 32'hc23c0d3b, 32'hc29de182, 32'h420dc460, 32'h41a6fe23, 32'h42745eb9};
test_weights[26776:26783] = '{32'h42a740c8, 32'hc29b198d, 32'h4006b62c, 32'h42b1062a, 32'hc219998e, 32'hc20d6537, 32'h429f9234, 32'hc2a0edfd};
test_bias[3347:3347] = '{32'hc2a3e0b9};
test_output[3347:3347] = '{32'hc5f4818f};
test_input[26784:26791] = '{32'hc223ed1f, 32'hc1fcf683, 32'h4283015f, 32'hc2953345, 32'h4201e56d, 32'hc1ade827, 32'h4075f1a7, 32'h42a2914a};
test_weights[26784:26791] = '{32'h42764019, 32'h41489204, 32'h40ae96a4, 32'hc24a6717, 32'h42575eae, 32'hc193c7f2, 32'hc06e5b9f, 32'hc1b5236f};
test_bias[3348:3348] = '{32'hc27672af};
test_output[3348:3348] = '{32'h44b4d1a1};
test_input[26792:26799] = '{32'hc28ecb55, 32'hc2b927ca, 32'h42478059, 32'h41fe32c9, 32'hc0b9150b, 32'hc20844a4, 32'h42ab1364, 32'h42c49069};
test_weights[26792:26799] = '{32'h40acd36d, 32'h422cbeaa, 32'hc16a8e76, 32'hc1d30b91, 32'h41807d61, 32'hc2706026, 32'hc29c56cb, 32'hc2c5cdb8};
test_bias[3349:3349] = '{32'hc26f1744};
test_output[3349:3349] = '{32'hc69fe283};
test_input[26800:26807] = '{32'hc294c41a, 32'h42c32b52, 32'hc0641fff, 32'hc2c04a3d, 32'hc236b0ae, 32'hc23dba33, 32'hc0947f51, 32'h41319a35};
test_weights[26800:26807] = '{32'hc1ff6ef1, 32'h41ef4a57, 32'hc18848c2, 32'hc1e6c2e8, 32'hc283654d, 32'hc29804ca, 32'h41c8d575, 32'h429b9650};
test_bias[3350:3350] = '{32'h424fb581};
test_output[3350:3350] = '{32'h4672b2da};
test_input[26808:26815] = '{32'h42af2289, 32'h42880e94, 32'hc1ea0fa7, 32'hc1815b12, 32'hc23f27dd, 32'h41f0ebdf, 32'hc21b9f25, 32'hc16e8d6e};
test_weights[26808:26815] = '{32'h41cb982a, 32'h4252e472, 32'hc1d5e172, 32'hc0b878cd, 32'h416d088e, 32'h4198c176, 32'hc2c46edf, 32'h426e1e8e};
test_bias[3351:3351] = '{32'h429ad514};
test_output[3351:3351] = '{32'h461582c2};
test_input[26816:26823] = '{32'hc1eba1cf, 32'h429eae42, 32'h41035f32, 32'hc1e4a766, 32'hc2ad01d3, 32'h42a12da5, 32'h40ff5137, 32'hc2c16172};
test_weights[26816:26823] = '{32'h42a96959, 32'hc1337692, 32'h42bbe4f9, 32'h403c2a24, 32'h415497a0, 32'hc2291728, 32'hc2c0c481, 32'h41357677};
test_bias[3352:3352] = '{32'hbe9752b5};
test_output[3352:3352] = '{32'hc60e7e01};
test_input[26824:26831] = '{32'hc28e3074, 32'h42082a3e, 32'hc2b2a8c9, 32'h41572fe1, 32'hc2753f63, 32'h42a0d8bf, 32'h42108f67, 32'hc281f735};
test_weights[26824:26831] = '{32'h42ada025, 32'hc243894f, 32'h42aa7083, 32'hc23e3f8f, 32'h41a288ac, 32'hc0ae3cfc, 32'h429ee645, 32'hc213055a};
test_bias[3353:3353] = '{32'hc2628782};
test_output[3353:3353] = '{32'hc64462f2};
test_input[26832:26839] = '{32'hc08481bd, 32'hc2935cc2, 32'h4262d9dc, 32'hc2bb780d, 32'h42086168, 32'h423f0374, 32'h4096365d, 32'h422d9e82};
test_weights[26832:26839] = '{32'h429485d2, 32'h420811ce, 32'hc2821e28, 32'hc290fd6b, 32'h42c68967, 32'hc1ef37b0, 32'h42a0dc4b, 32'hc23d6875};
test_bias[3354:3354] = '{32'hc28a8393};
test_output[3354:3354] = '{32'h43faa4e9};
test_input[26840:26847] = '{32'h41c72913, 32'h423037e7, 32'hc1709509, 32'hc2b9f382, 32'h42c5d77f, 32'hc2be705a, 32'h42926639, 32'h42b7cab6};
test_weights[26840:26847] = '{32'hc23763b4, 32'hc1c5b190, 32'hc2708fc1, 32'h420b136e, 32'h42ba06e3, 32'h4222b9a8, 32'hc06b4220, 32'hc2c26487};
test_bias[3355:3355] = '{32'h41cea29f};
test_output[3355:3355] = '{32'hc603591f};
test_input[26848:26855] = '{32'hc239ea1a, 32'h423f4766, 32'h41c398fb, 32'h4142f3d8, 32'hc24949b9, 32'h429240c5, 32'h420903cd, 32'hc212d0eb};
test_weights[26848:26855] = '{32'h42039d85, 32'h41f249e3, 32'h42a33dff, 32'hc2817351, 32'hc15fa163, 32'h42b17107, 32'h41aa1cdb, 32'h40c6d950};
test_bias[3356:3356] = '{32'hc283d690};
test_output[3356:3356] = '{32'h4608bde2};
test_input[26856:26863] = '{32'h4246f17d, 32'h41940ae8, 32'hc20fd82e, 32'hc23631f0, 32'hc24f13f5, 32'hc280ea3d, 32'h429c5870, 32'h42c01c4b};
test_weights[26856:26863] = '{32'h428c4cf3, 32'h420574bc, 32'hc21407bf, 32'h3fd3025b, 32'h4247ce8a, 32'hc22e49d8, 32'hc1c826b7, 32'hc25dee6f};
test_bias[3357:3357] = '{32'h42c271c9};
test_output[3357:3357] = '{32'hc4c868e3};
test_input[26864:26871] = '{32'h41c196a3, 32'h3fc378de, 32'hc2bfc721, 32'hc19182bf, 32'hc2b5c5f3, 32'hc2956a2f, 32'hc21f356c, 32'h423208f9};
test_weights[26864:26871] = '{32'hc2016beb, 32'h42b096c1, 32'hc23c7998, 32'hc2904319, 32'h42b48258, 32'h4279cf4a, 32'h42b53ee6, 32'hc2a6b1d4};
test_bias[3358:3358] = '{32'h420348ef};
test_output[3358:3358] = '{32'hc669e9a7};
test_input[26872:26879] = '{32'h425a1a57, 32'hc0d0da10, 32'hc27488ba, 32'hc29815dd, 32'hc28a9e63, 32'hc20cfbde, 32'hc1d5f8c2, 32'hc2bc7993};
test_weights[26872:26879] = '{32'h429f4726, 32'hc1f2cb97, 32'hc2a4cdbe, 32'h41626340, 32'h42472841, 32'hc24f482a, 32'hc276b7e9, 32'hc29de240};
test_bias[3359:3359] = '{32'h428bba87};
test_output[3359:3359] = '{32'h467a91e8};
test_input[26880:26887] = '{32'h41ad23e6, 32'h42bed2c0, 32'h41e61994, 32'hc2b41209, 32'hc11681d8, 32'h4276bd2c, 32'h42a7fa1d, 32'h41d1e7e5};
test_weights[26880:26887] = '{32'h42675bc6, 32'h42a52795, 32'hc2c53ac0, 32'h42a2bbff, 32'hc2c7465b, 32'hc1ccc09f, 32'hc29e4e70, 32'h405bcf66};
test_bias[3360:3360] = '{32'h41df5ad4};
test_output[3360:3360] = '{32'hc6002c74};
test_input[26888:26895] = '{32'hc288d1a8, 32'h4281ec0d, 32'hc16b5287, 32'h427d2100, 32'hc1c45648, 32'hc280ac40, 32'hc1f981d6, 32'h42700fd2};
test_weights[26888:26895] = '{32'hc2c4852a, 32'h41ad1d38, 32'h423377e4, 32'h4213e284, 32'h4270ea68, 32'h421e1314, 32'h4296e62d, 32'hc22ed795};
test_bias[3361:3361] = '{32'hc1f6eea3};
test_output[3361:3361] = '{32'h4442d9d7};
test_input[26896:26903] = '{32'hc1a5dc8e, 32'hc287061e, 32'hc2a2d8dc, 32'h421b6809, 32'h4298da28, 32'h428cbf32, 32'h4273ba52, 32'h41ef418b};
test_weights[26896:26903] = '{32'h42b7b49e, 32'h4289bd0e, 32'hc294db46, 32'h4281cd94, 32'h4213678d, 32'hc2adaa3b, 32'hc2a68c2e, 32'h427fc3af};
test_bias[3362:3362] = '{32'hc01ef91f};
test_output[3362:3362] = '{32'hc58a753f};
test_input[26904:26911] = '{32'h4297b51e, 32'hc207c0a6, 32'h41f12879, 32'h425b633a, 32'h41276b54, 32'h4248def0, 32'h428e473e, 32'hc2b49380};
test_weights[26904:26911] = '{32'h423160b8, 32'hc1e1e045, 32'hc2222ec9, 32'hc27152a2, 32'hc2bdd7d7, 32'hc176a2b9, 32'hc22fe7a6, 32'hc2754bc5};
test_bias[3363:3363] = '{32'hbf990ba6};
test_output[3363:3363] = '{32'h43d74d48};
test_input[26912:26919] = '{32'hc1a80fe5, 32'h41b5cfd4, 32'hc2135b4a, 32'hc261cb2d, 32'h429ee367, 32'h4007b195, 32'h41b91ecf, 32'hc2a91fb0};
test_weights[26912:26919] = '{32'h42ac3c38, 32'h4286cf36, 32'h42ac7e60, 32'hc2aff87c, 32'hc2c5f6e9, 32'h413229a4, 32'h429f2a8a, 32'h42aa63b4};
test_bias[3364:3364] = '{32'h428659ae};
test_output[3364:3364] = '{32'hc6359d5e};
test_input[26920:26927] = '{32'hc2991d24, 32'h41a32fa2, 32'h4298ce7e, 32'h41255f6f, 32'h42acb8b1, 32'hc297be91, 32'h409b4c58, 32'h42989b7f};
test_weights[26920:26927] = '{32'hc27ccea4, 32'h42903d92, 32'hc1e397bd, 32'hc12be4b8, 32'h429e076f, 32'h42bc112d, 32'hc15018d3, 32'h42c78e7c};
test_bias[3365:3365] = '{32'h42730558};
test_output[3365:3365] = '{32'h4630f54c};
test_input[26928:26935] = '{32'hc1ebfdcb, 32'h427e0d73, 32'h40846f66, 32'hc1d588b2, 32'hc29effca, 32'h41ad597e, 32'hc20f1aac, 32'h42bb861c};
test_weights[26928:26935] = '{32'h4161d5bd, 32'h42788adc, 32'h4279f9ae, 32'h41cbb77a, 32'hc20ce3fb, 32'h423e91bc, 32'h42294246, 32'hc1f60e28};
test_bias[3366:3366] = '{32'hc1a601d5};
test_output[3366:3366] = '{32'h451db1a3};
test_input[26936:26943] = '{32'hc1167d46, 32'h42c2d8f1, 32'h421738ff, 32'hc25ad644, 32'h4207cade, 32'hc2bda6ed, 32'hc250ecec, 32'h42918fdd};
test_weights[26936:26943] = '{32'hc2919aa1, 32'hc28c4fbd, 32'hc2a63eec, 32'h427eef03, 32'h4085dc1f, 32'hc128846e, 32'h423e7e7b, 32'hc2b8eb27};
test_bias[3367:3367] = '{32'h4291d325};
test_output[3367:3367] = '{32'hc6a25cf0};
test_input[26944:26951] = '{32'hc2590d43, 32'h42012f73, 32'h419b909a, 32'hc1d7e647, 32'hc1ab7388, 32'hc2b758c3, 32'hc20bef81, 32'hc1eb8c13};
test_weights[26944:26951] = '{32'h4217e8de, 32'h4296fc0b, 32'h41fc0ea5, 32'hc23b78cf, 32'hc206ab88, 32'hc21eb6bd, 32'h424319c7, 32'hc1bceedf};
test_bias[3368:3368] = '{32'h424cbcd5};
test_output[3368:3368] = '{32'h45b0b095};
test_input[26952:26959] = '{32'h4297e16e, 32'hc15dcac2, 32'hc235064f, 32'hc2b6ecf8, 32'h4218acbd, 32'hc1a3aa1a, 32'hc2bedbdb, 32'h42023e84};
test_weights[26952:26959] = '{32'h423dfb7b, 32'hc25f3cd8, 32'h4274c23c, 32'h421d5348, 32'hc29a833d, 32'h42526150, 32'hc294c5ad, 32'hc11020ef};
test_bias[3369:3369] = '{32'hc282c29a};
test_output[3369:3369] = '{32'h443643b2};
test_input[26960:26967] = '{32'h426a1d3c, 32'h42bf370e, 32'h427ce338, 32'h42a669f9, 32'h419501aa, 32'h41ab4484, 32'h42b8596f, 32'hc222160d};
test_weights[26960:26967] = '{32'hc17b0787, 32'h42a47a24, 32'h41bdc064, 32'h4263b40b, 32'hc264afb6, 32'hc28457e8, 32'hc2992d1a, 32'hc2391f43};
test_bias[3370:3370] = '{32'hc22d31a6};
test_output[3370:3370] = '{32'h45aafce0};
test_input[26968:26975] = '{32'hc1215b66, 32'hc2b105b7, 32'h41cffdb4, 32'hc28ad0fe, 32'h4250f51c, 32'h42bcd8e9, 32'h420e0aee, 32'hc2a72e13};
test_weights[26968:26975] = '{32'h42097dd7, 32'hc1ab9691, 32'hc2a851a4, 32'h41f7c94d, 32'h421ef4fc, 32'h42b5dba2, 32'h4289e824, 32'hc22c3f98};
test_bias[3371:3371] = '{32'h42b085a1};
test_output[3371:3371] = '{32'h465af08f};
test_input[26976:26983] = '{32'h425c16ea, 32'h4235f033, 32'h418dbf9d, 32'hc2a4b6bf, 32'h41f1fe16, 32'hc2b1f2d3, 32'h4203775d, 32'hc2a6d070};
test_weights[26976:26983] = '{32'h42b77201, 32'hc29dbd3f, 32'h4223e836, 32'h42c01e13, 32'hc26f8dd7, 32'hc2910a14, 32'hc2b16ac6, 32'hc2498069};
test_bias[3372:3372] = '{32'hc29b0878};
test_output[3372:3372] = '{32'h42f7a07c};
test_input[26984:26991] = '{32'hc2477519, 32'h420eaf19, 32'hc28be514, 32'h41eaae8e, 32'h42565f43, 32'h4081f6bf, 32'hc23e9c94, 32'h42ad157b};
test_weights[26984:26991] = '{32'h40ba777e, 32'hc2798b0a, 32'h429f4a6a, 32'h3fd6f95c, 32'h4214338f, 32'h41f95c5b, 32'h424c29de, 32'h4218cba4};
test_bias[3373:3373] = '{32'h425f48c9};
test_output[3373:3373] = '{32'hc59c2041};
test_input[26992:26999] = '{32'hc28ebb20, 32'h41bc6bd9, 32'hc2332188, 32'h42209625, 32'hc2658435, 32'hc1dfaa51, 32'hc28e1ed2, 32'hc2c1167a};
test_weights[26992:26999] = '{32'hc2a21599, 32'h420471c2, 32'h42a6a2fc, 32'hc0cf7f01, 32'hc2a511a7, 32'h421bc947, 32'hc2c1a79b, 32'hc18fa8f0};
test_bias[3374:3374] = '{32'h4286383d};
test_output[3374:3374] = '{32'h4668d0b0};
test_input[27000:27007] = '{32'h3f900569, 32'hc1ab7268, 32'h42907a6a, 32'h429a923a, 32'hc234518a, 32'hc22c1532, 32'hc28c1ff4, 32'h4259db85};
test_weights[27000:27007] = '{32'h41e6ab37, 32'h41943d26, 32'h40c58eb8, 32'h42512bb6, 32'h4219d648, 32'hc12843d5, 32'h423af9f3, 32'hc1e9bf2c};
test_bias[3375:3375] = '{32'hbffb412d};
test_output[3375:3375] = '{32'hc4fd5ae7};
test_input[27008:27015] = '{32'hc29c2428, 32'hc1d0a284, 32'hc2aac2e2, 32'hc24d999c, 32'hc29c1216, 32'h4117480e, 32'h42b7d7ca, 32'hc208fcf6};
test_weights[27008:27015] = '{32'h41ebb40e, 32'h4277d974, 32'h42b21996, 32'h42c4c299, 32'h41b1bcd7, 32'h427fcdcd, 32'hc1ac3823, 32'hc10d2c68};
test_bias[3376:3376] = '{32'hc28912ab};
test_output[3376:3376] = '{32'hc697f488};
test_input[27016:27023] = '{32'h41e478b3, 32'h41a2874b, 32'hc23ced81, 32'h42055e60, 32'hc122adac, 32'hc1070889, 32'h42a0cf9d, 32'hbfef95ca};
test_weights[27016:27023] = '{32'hc2ad06dc, 32'hc16144fb, 32'h415c51f8, 32'hc2043c1e, 32'h42870869, 32'hc287ea8d, 32'h42965e49, 32'hc2ae12fa};
test_bias[3377:3377] = '{32'hc21fad50};
test_output[3377:3377] = '{32'h44c13c42};
test_input[27024:27031] = '{32'h42b54bf2, 32'hc1f07baa, 32'hc23a9a67, 32'hc2b19e85, 32'hc1f97eca, 32'h4258b1fa, 32'h41a2f60f, 32'h413cc7ea};
test_weights[27024:27031] = '{32'h426ad51c, 32'h41f12f69, 32'hc230ccd2, 32'h41213bb8, 32'hc2c00728, 32'h4284e4e9, 32'h41c6593b, 32'hc267dddc};
test_bias[3378:3378] = '{32'h41e682c6};
test_output[3378:3378] = '{32'h463bea31};
test_input[27032:27039] = '{32'h411ad244, 32'h429ea9bc, 32'h421f8919, 32'hc1e8d02b, 32'h4297daab, 32'hc244521e, 32'h42aa6036, 32'hc1b350bd};
test_weights[27032:27039] = '{32'h42991e15, 32'hc081ce3c, 32'hc2c399b8, 32'hc1b2002e, 32'hc2b349ee, 32'hc2b74012, 32'hc2a33c38, 32'h4293c351};
test_bias[3379:3379] = '{32'hc2249a5f};
test_output[3379:3379] = '{32'hc6578659};
test_input[27040:27047] = '{32'hc21182cf, 32'hc201c75b, 32'h424cefc9, 32'hc2b788de, 32'hc20d1232, 32'hc1f1e9f2, 32'h42ad0433, 32'h425fe04d};
test_weights[27040:27047] = '{32'h42800cf3, 32'h4291ab64, 32'hc1cd6264, 32'h42a44f03, 32'h41b877e1, 32'h406ca4fb, 32'h4234f984, 32'hc2669fc6};
test_bias[3380:3380] = '{32'hc29943c2};
test_output[3380:3380] = '{32'hc6589525};
test_input[27048:27055] = '{32'hc2ba87cb, 32'h4241f9e0, 32'hc25f4e10, 32'h42ad823c, 32'hc1bd9229, 32'h42227d7d, 32'hc2ab8e8a, 32'hc1def48b};
test_weights[27048:27055] = '{32'h418c9273, 32'hc208044f, 32'hbf29732a, 32'h40adbb33, 32'h41491d16, 32'h4260b9d8, 32'h42c2405b, 32'h42927eaa};
test_bias[3381:3381] = '{32'h4203ea44};
test_output[3381:3381] = '{32'hc62dfc97};
test_input[27056:27063] = '{32'hc20732a1, 32'hc2acd154, 32'h425eba3e, 32'hc2c2549e, 32'h42bf5ddd, 32'hc2311250, 32'hc2087fb8, 32'h423f6123};
test_weights[27056:27063] = '{32'h425351c4, 32'h429658f4, 32'hc2593397, 32'h41ca467a, 32'hc2937d3e, 32'hc1ae91f7, 32'hc2b0a4ac, 32'h4033e40d};
test_bias[3382:3382] = '{32'hc2883f00};
test_output[3382:3382] = '{32'hc68306e5};
test_input[27064:27071] = '{32'h4289ec69, 32'hc294f5a4, 32'h42a098ae, 32'h42ae8d7d, 32'h429d9cc1, 32'h429bb901, 32'h40cfd2f4, 32'h428c1e81};
test_weights[27064:27071] = '{32'h42b24836, 32'hc2b64dd6, 32'hc25101b4, 32'h4231937f, 32'h42189a69, 32'h427fe717, 32'hc2bdb265, 32'h4180e1c3};
test_bias[3383:3383] = '{32'hc214ef91};
test_output[3383:3383] = '{32'h46a4acac};
test_input[27072:27079] = '{32'h42b96108, 32'h419ddb9a, 32'hc2698d63, 32'hc205d8a0, 32'h41e1f6ec, 32'hc152b33d, 32'hc2a04893, 32'hc25948fc};
test_weights[27072:27079] = '{32'h42b0be1a, 32'hc28c8b98, 32'hc2506abb, 32'hc0b2a667, 32'h42b1a1d7, 32'hc21b192a, 32'hbfcec142, 32'hc2675f4a};
test_bias[3384:3384] = '{32'h4256cf09};
test_output[3384:3384] = '{32'h467fe844};
test_input[27080:27087] = '{32'h4261bb10, 32'hc202d094, 32'hc29604eb, 32'h42aae8ce, 32'hc1491b05, 32'hbffacea0, 32'h41679c93, 32'h4276a9a1};
test_weights[27080:27087] = '{32'h426bfb6e, 32'hc26e7dfe, 32'hc207d6ba, 32'h4260da50, 32'h42ad06e5, 32'hc28387f4, 32'h4277c919, 32'h42a16613};
test_bias[3385:3385] = '{32'h412dd954};
test_output[3385:3385] = '{32'h4689272b};
test_input[27088:27095] = '{32'h420243c9, 32'h3c904b88, 32'h428e1ed1, 32'h41becfa5, 32'h420f987d, 32'hc2bb0422, 32'hc2a00b6e, 32'h42c2a849};
test_weights[27088:27095] = '{32'hc210f0dd, 32'h42326ed3, 32'hc21f6701, 32'hc251d881, 32'hc2566c7c, 32'h4202b77c, 32'hc28f943b, 32'h425bf102};
test_bias[3386:3386] = '{32'hc10ec346};
test_output[3386:3386] = '{32'h44534051};
test_input[27096:27103] = '{32'h42991143, 32'hc273c524, 32'hc28b94f3, 32'h42950285, 32'hc2afbb6d, 32'h41f85859, 32'hc2a4be4d, 32'hc1bed2cf};
test_weights[27096:27103] = '{32'h42947c04, 32'h42afb4d5, 32'hc08cb4f3, 32'hc267b3bf, 32'h42bd0a12, 32'h42803892, 32'hc1e51a63, 32'h408be1a8};
test_bias[3387:3387] = '{32'h4282b46d};
test_output[3387:3387] = '{32'hc5efdd5a};
test_input[27104:27111] = '{32'hc2129f41, 32'hc1c90973, 32'h4280648a, 32'hc2052075, 32'hc23941e2, 32'h4290ca15, 32'hc2ac7cf3, 32'h42c4e4dd};
test_weights[27104:27111] = '{32'h42b6e6b4, 32'hc297c21e, 32'h42b5a16d, 32'h42c48303, 32'hc2621400, 32'h42a9c6cd, 32'hc16c943c, 32'h42c48608};
test_bias[3388:3388] = '{32'hbe1e5da4};
test_output[3388:3388] = '{32'h46a2b49b};
test_input[27112:27119] = '{32'h40a0282a, 32'hc15ecd4f, 32'hc0cbf010, 32'hc2916482, 32'hc21c9999, 32'hc2920af4, 32'hc2b6124a, 32'h4184394c};
test_weights[27112:27119] = '{32'hc0faf2d5, 32'hc2c7cd48, 32'h425b62c1, 32'hc25d4e16, 32'hc2c74e91, 32'h429fa977, 32'h3dbe071e, 32'h424ff835};
test_bias[3389:3389] = '{32'h40d3a900};
test_output[3389:3389] = '{32'h45771eaf};
test_input[27120:27127] = '{32'hc240dabf, 32'hc26f20d3, 32'h42476a54, 32'hc2c29b82, 32'h4245e0a0, 32'h4273edf0, 32'h428d6648, 32'hc2604ec5};
test_weights[27120:27127] = '{32'h423b251b, 32'hc1bd10c5, 32'h424cbe40, 32'hc246cca0, 32'hc1cee13a, 32'h4293fe33, 32'h4243b333, 32'h4237a014};
test_bias[3390:3390] = '{32'h42b9a976};
test_output[3390:3390] = '{32'h46280e84};
test_input[27128:27135] = '{32'h42c5cd64, 32'h41e7e54c, 32'hc29124e7, 32'h421d73c6, 32'h4175870e, 32'hc1e157de, 32'hc0cbe69c, 32'hc190ede7};
test_weights[27128:27135] = '{32'hc2ae7fff, 32'h42b865ea, 32'hc143a612, 32'hc2a0155b, 32'h41de6351, 32'hc29dca33, 32'hc2c19332, 32'h4139b72f};
test_bias[3391:3391] = '{32'h42082a89};
test_output[3391:3391] = '{32'hc5a053a9};
test_input[27136:27143] = '{32'h424bc8e3, 32'hc1337555, 32'hc26aa5d4, 32'hc287a7d5, 32'hc1df31d5, 32'h41f471d7, 32'h42c0c549, 32'h4205bf6d};
test_weights[27136:27143] = '{32'hc20f29cb, 32'hc263b95b, 32'h42483bca, 32'hc27a30ef, 32'h4277fbb3, 32'h422506b8, 32'hc2852df9, 32'h42173e94};
test_bias[3392:3392] = '{32'hc1987831};
test_output[3392:3392] = '{32'hc5ac87cc};
test_input[27144:27151] = '{32'h428a8218, 32'h42925b55, 32'h42b10e9a, 32'h4244eb58, 32'h421dbeed, 32'h4286ef32, 32'hc24e953f, 32'h421ab86c};
test_weights[27144:27151] = '{32'h416e557f, 32'h4271966c, 32'hc2b67fdb, 32'hc28c37bb, 32'hc1d48f7c, 32'hc1e09bd8, 32'hc26df9b8, 32'hc2b0498c};
test_bias[3393:3393] = '{32'h403c5433};
test_output[3393:3393] = '{32'hc61228cf};
test_input[27152:27159] = '{32'hc18e4714, 32'h3ee05eaf, 32'hc19435e9, 32'h416c5aca, 32'hc265d91d, 32'h4058ca55, 32'hc1ae8dd9, 32'h413cf546};
test_weights[27152:27159] = '{32'h42c29162, 32'hc0b355dc, 32'h42780c8f, 32'hc2244afd, 32'hc29779e5, 32'hc2c40c7c, 32'hc2bf31b3, 32'hc0dbdcec};
test_bias[3394:3394] = '{32'hc215859f};
test_output[3394:3394] = '{32'h451c3220};
test_input[27160:27167] = '{32'h41938093, 32'hc1ad35ca, 32'hc2c28732, 32'h4245c278, 32'hc1d5ce0a, 32'h42b4a97d, 32'hc126a70d, 32'hc2531dfa};
test_weights[27160:27167] = '{32'h4111e9c1, 32'hc268b38e, 32'hc278a02d, 32'hc1bee3f7, 32'h40bcaacb, 32'hc2956e28, 32'hc1905025, 32'h42891e1a};
test_bias[3395:3395] = '{32'hc21a67a5};
test_output[3395:3395] = '{32'hc57f242a};
test_input[27168:27175] = '{32'hc217216a, 32'hc26f87f0, 32'h4288bbe6, 32'h4263aa99, 32'hc2ba4245, 32'hc1d43726, 32'h420e1be8, 32'hc2aa5d6d};
test_weights[27168:27175] = '{32'h41ca20e9, 32'h41e090b7, 32'h415468de, 32'hc240f247, 32'h41193732, 32'hc25098c0, 32'h42c4ae49, 32'hc19d6b33};
test_bias[3396:3396] = '{32'hc27c1650};
test_output[3396:3396] = '{32'h448ca158};
test_input[27176:27183] = '{32'hc1e324bc, 32'h4254f05c, 32'h4148c4ca, 32'h41924563, 32'h429629cb, 32'hc287a322, 32'h4282eda8, 32'hc29c6137};
test_weights[27176:27183] = '{32'hc1108b2c, 32'hc2b15c24, 32'hc13910fe, 32'hc13ce89b, 32'hc26da80c, 32'hc2178d11, 32'hc2c26435, 32'hc24f4958};
test_bias[3397:3397] = '{32'hc23bcf21};
test_output[3397:3397] = '{32'hc60dca90};
test_input[27184:27191] = '{32'h42b074f9, 32'hc10db2ee, 32'h42621141, 32'h41cef485, 32'hc224f769, 32'h428bf1f2, 32'hc2aaa45b, 32'h4183e5b0};
test_weights[27184:27191] = '{32'hc1572b98, 32'hc291fe6e, 32'hc21b00c6, 32'h41d858e7, 32'h421b4633, 32'h423a55b7, 32'hc2c51094, 32'h429b417d};
test_bias[3398:3398] = '{32'hc270f2f8};
test_output[3398:3398] = '{32'h46109a8f};
test_input[27192:27199] = '{32'hc0d1ca3b, 32'hc122fa46, 32'hc1d6872f, 32'hc281aaaf, 32'h410e6f74, 32'hc1b2e827, 32'hc245dc72, 32'hbfb1214d};
test_weights[27192:27199] = '{32'h41a9f55b, 32'h4264265e, 32'h4269631b, 32'h41ea7c3b, 32'hc028ec56, 32'h420e336a, 32'h429286fc, 32'h403c4bde};
test_bias[3399:3399] = '{32'hc28b356c};
test_output[3399:3399] = '{32'hc607f5a0};
test_input[27200:27207] = '{32'h42a7548d, 32'hc20ca432, 32'hc1056b5e, 32'hc0c3eae1, 32'h42998b4b, 32'h427524fb, 32'hc21d4bfe, 32'hc2231485};
test_weights[27200:27207] = '{32'hc251de7c, 32'hc283973b, 32'hc035d153, 32'hc005eb27, 32'hc22c9598, 32'h42bfa87c, 32'h427ba30a, 32'hc202c060};
test_bias[3400:3400] = '{32'hc275ef10};
test_output[3400:3400] = '{32'hc42a77a2};
test_input[27208:27215] = '{32'h42b1aefe, 32'hc0b31cba, 32'hc1a7341b, 32'h40cfd258, 32'hc2a75ec1, 32'h414b6828, 32'hc2636186, 32'hc12b3bdb};
test_weights[27208:27215] = '{32'hc0bafbf2, 32'h4284bdad, 32'h419d33a9, 32'h423add7d, 32'h424aaa92, 32'h4194d047, 32'h418be5aa, 32'h41769e5e};
test_bias[3401:3401] = '{32'h426db0ba};
test_output[3401:3401] = '{32'hc5bea891};
test_input[27216:27223] = '{32'hc1069dac, 32'hc295081b, 32'hc21810be, 32'hc2ac9a8e, 32'hc2b658f9, 32'h418e4834, 32'hc2a79ad2, 32'h424b8691};
test_weights[27216:27223] = '{32'h42889485, 32'hc2adff2e, 32'h42be178b, 32'h404a1d3c, 32'hc1e2c7f1, 32'h4074ebe3, 32'h40334265, 32'hc20385f1};
test_bias[3402:3402] = '{32'h41a39667};
test_output[3402:3402] = '{32'h452e3ade};
test_input[27224:27231] = '{32'h41860ca7, 32'h41b1f63d, 32'hc29953ac, 32'h426cbb83, 32'hc23eec68, 32'hc1fa18a7, 32'hc2708eb1, 32'hc291d45e};
test_weights[27224:27231] = '{32'h41b346ae, 32'hc0649ec2, 32'hc1888024, 32'hc26b7591, 32'h41f9fcfe, 32'hc2ad7bbd, 32'h42a00d80, 32'h4204a472};
test_bias[3403:3403] = '{32'hc217453c};
test_output[3403:3403] = '{32'hc5f7bf87};
test_input[27232:27239] = '{32'h4257e730, 32'hc2041db8, 32'hc2b435ea, 32'hc21ae38d, 32'h42bc92b1, 32'h420d21e7, 32'hc16e09ee, 32'h4263b870};
test_weights[27232:27239] = '{32'hc2bd60ac, 32'h4295f0d7, 32'hc25d426e, 32'hc2b6fe97, 32'h4272171a, 32'h41caddc4, 32'h41f75921, 32'h4245cc03};
test_bias[3404:3404] = '{32'h428984ea};
test_output[3404:3404] = '{32'h461bb490};
test_input[27240:27247] = '{32'h42af58ac, 32'hc28297e0, 32'h4233396d, 32'hc1c007e8, 32'h41a468c4, 32'h42a0fd83, 32'hc1ce1bcb, 32'h415182c0};
test_weights[27240:27247] = '{32'hc2c1a413, 32'hc28fb9ee, 32'hc201c2da, 32'h41240f24, 32'h4274fc51, 32'hc2c039e2, 32'h40ba2d9b, 32'hc2909cec};
test_bias[3405:3405] = '{32'h42a7b572};
test_output[3405:3405] = '{32'hc64aea5a};
test_input[27248:27255] = '{32'hbfb2222c, 32'h42814927, 32'h420a52a0, 32'h42550c42, 32'hc2641e03, 32'h42543719, 32'h41b7de9b, 32'h42c675e6};
test_weights[27248:27255] = '{32'hc2b45425, 32'hc216879c, 32'h42a29b5c, 32'hc0e49329, 32'hc2c0ad5c, 32'h4243420b, 32'h4198f962, 32'hc2676fee};
test_bias[3406:3406] = '{32'h42a09eaa};
test_output[3406:3406] = '{32'h453aa36a};
test_input[27256:27263] = '{32'h3f28212c, 32'hc2b3c6d8, 32'h41408b4b, 32'hc21becb3, 32'hc2bb4ca5, 32'hc2b1f2fb, 32'h4221395c, 32'h42a0b164};
test_weights[27256:27263] = '{32'h42723c91, 32'hc23469cb, 32'hc2448bf7, 32'hc295998f, 32'h429d8f45, 32'h42859351, 32'hc2418fc6, 32'hc2c5408d};
test_bias[3407:3407] = '{32'hc1e07bd2};
test_output[3407:3407] = '{32'hc68348b1};
test_input[27264:27271] = '{32'hc1473cbe, 32'h428f65c7, 32'hc2661f96, 32'hc2848c19, 32'h4285be05, 32'h42a5e1c3, 32'hc191adfa, 32'h425393a2};
test_weights[27264:27271] = '{32'h429f0588, 32'h42c6da38, 32'hc20c7718, 32'h41d38b32, 32'hc28882a7, 32'h42313545, 32'h41cad870, 32'h42c29144};
test_bias[3408:3408] = '{32'h4235b64a};
test_output[3408:3408] = '{32'h46201826};
test_input[27272:27279] = '{32'hc2986b6f, 32'h42a0fd9f, 32'h423f3d31, 32'h4155ec0d, 32'hc259d9c6, 32'h42a149cc, 32'h42c66cd0, 32'h41f970a7};
test_weights[27272:27279] = '{32'h421a5018, 32'h428561da, 32'hc2b2db61, 32'hc26015ca, 32'hc213cd7a, 32'hc287cb34, 32'hc28df5fd, 32'hc1e435c7};
test_bias[3409:3409] = '{32'h42b24775};
test_output[3409:3409] = '{32'hc659372b};
test_input[27280:27287] = '{32'hbf96413d, 32'hc2b13049, 32'h423a5181, 32'hc24947fc, 32'hc1cdc529, 32'h42a52d24, 32'hc1b2aa9c, 32'h422cf992};
test_weights[27280:27287] = '{32'hc1172e1a, 32'h4192b63e, 32'h42498d78, 32'h41911d8a, 32'h41da0aa2, 32'hc29e330a, 32'hc19531cd, 32'h424361d3};
test_bias[3410:3410] = '{32'hc20875e1};
test_output[3410:3410] = '{32'hc599b394};
test_input[27288:27295] = '{32'h42251c75, 32'hc2bbbc29, 32'h42aea069, 32'h42c12482, 32'h4273bcf5, 32'hc24c9336, 32'h42be04e4, 32'hc0add0fd};
test_weights[27288:27295] = '{32'hc1e1f5e7, 32'hc0afbdac, 32'hc1bc3ae4, 32'hc28f1528, 32'h417b2a54, 32'hc0020816, 32'h420bcb97, 32'hc2a5b753};
test_bias[3411:3411] = '{32'hc224c9cb};
test_output[3411:3411] = '{32'hc596be6f};
test_input[27296:27303] = '{32'hc1976b81, 32'h4296ecb4, 32'h424f220c, 32'hc108e6aa, 32'hc29229ce, 32'h41ec2092, 32'hc15b1661, 32'h42b7cf11};
test_weights[27296:27303] = '{32'h41909e03, 32'hc2a8d8dd, 32'h3fef503d, 32'hc1c8914d, 32'h42211b29, 32'h42a13686, 32'hc2a241d9, 32'h426c0aa8};
test_bias[3412:3412] = '{32'hc26249f3};
test_output[3412:3412] = '{32'hc3f424a4};
test_input[27304:27311] = '{32'h4251573d, 32'h428ee420, 32'hc2a6c306, 32'h4297f249, 32'h4249d939, 32'h42c29d12, 32'h41956e85, 32'hc227c62a};
test_weights[27304:27311] = '{32'hc297d53e, 32'hc22953bf, 32'h42bc8d40, 32'h411e743e, 32'h418712de, 32'h41cdc504, 32'h42a01374, 32'h42b93e4b};
test_bias[3413:3413] = '{32'h42be18e1};
test_output[3413:3413] = '{32'hc64bd787};
test_input[27312:27319] = '{32'hc00eceae, 32'hc28fdc83, 32'h422e2734, 32'h42260365, 32'hc25f2254, 32'h42b4aca2, 32'hc28ea42c, 32'h40c3d3a7};
test_weights[27312:27319] = '{32'hc1b5396b, 32'hc2825e6b, 32'hc1f6f53d, 32'h42a153de, 32'h41e7ad5b, 32'h4116cc04, 32'hc29c32bb, 32'hc2b570c3};
test_bias[3414:3414] = '{32'hc2515db0};
test_output[3414:3414] = '{32'h462af672};
test_input[27320:27327] = '{32'hc29e97a1, 32'h425592b8, 32'hc2b7a5e2, 32'hc29ccc57, 32'hc29e27ad, 32'hc27fb748, 32'h42be3d10, 32'h41f6952e};
test_weights[27320:27327] = '{32'h42a9dca9, 32'h4224aff6, 32'hc2ac2ec1, 32'hc2986eec, 32'h417bad61, 32'hc1fe12f7, 32'h41d3c231, 32'hc0658e51};
test_bias[3415:3415] = '{32'hc29f7cd1};
test_output[3415:3415] = '{32'h4642a878};
test_input[27328:27335] = '{32'h4207f74f, 32'hc05ebcda, 32'h42a7a9e2, 32'hc28ac7b2, 32'h426b0cd3, 32'h4225ca6f, 32'hc298ea10, 32'h4242d4ed};
test_weights[27328:27335] = '{32'h4298ca4f, 32'hc132c051, 32'hc279ff6e, 32'hc0a54f40, 32'hc289024c, 32'h42a84870, 32'h422f6676, 32'hc171ccbf};
test_bias[3416:3416] = '{32'h423a58bd};
test_output[3416:3416] = '{32'hc5d54bfd};
test_input[27336:27343] = '{32'h41f39639, 32'h42bb6f09, 32'hc25c25b8, 32'hc0e2900b, 32'hc13e00cf, 32'h41680eef, 32'h411e4ce4, 32'h421aa0a1};
test_weights[27336:27343] = '{32'h424e4862, 32'hc2986601, 32'h42997926, 32'hc192c1c7, 32'h42988103, 32'hc28b8062, 32'hc22b67f7, 32'h429d9ae0};
test_bias[3417:3417] = '{32'hc260dc63};
test_output[3417:3417] = '{32'hc60cddc1};
test_input[27344:27351] = '{32'h40df12ec, 32'h40166a9c, 32'h414c1505, 32'h429bf695, 32'hc27a229c, 32'h42c5ebd0, 32'hc2a890a6, 32'h3f9d5e8c};
test_weights[27344:27351] = '{32'h41689f24, 32'h428b9064, 32'h429e3895, 32'hc26cee12, 32'h42127dda, 32'h41c5837f, 32'h41bfbce9, 32'hc22f8e25};
test_bias[3418:3418] = '{32'hc2bb92cb};
test_output[3418:3418] = '{32'hc5a77a65};
test_input[27352:27359] = '{32'h41332c17, 32'h3dfdd04b, 32'h42c16f3a, 32'h42728c4d, 32'h426002fd, 32'hc2619354, 32'h4180aa00, 32'h41f4dd10};
test_weights[27352:27359] = '{32'hc1944903, 32'h42493946, 32'hc081e902, 32'h41b9ec7f, 32'h42b487d0, 32'h42a9769b, 32'h420a7609, 32'hc246182e};
test_bias[3419:3419] = '{32'hc2c1c79f};
test_output[3419:3419] = '{32'h42102b0e};
test_input[27360:27367] = '{32'hc1ae3b44, 32'hc2c7325f, 32'h402cbc96, 32'hc1bf2034, 32'h428cbc9d, 32'hc1857685, 32'h41643e2e, 32'hc148c4cd};
test_weights[27360:27367] = '{32'hc130afd5, 32'hc2b3eb1c, 32'h41039fe5, 32'h428a23a9, 32'h42bc4f8e, 32'h429992b9, 32'h418548e9, 32'h4270c806};
test_bias[3420:3420] = '{32'h4288fbe3};
test_output[3420:3420] = '{32'h4642cef6};
test_input[27368:27375] = '{32'hc24888ad, 32'h41a01d91, 32'h427799aa, 32'h42bd4ab9, 32'h42968a11, 32'hc2237dbf, 32'h401b7411, 32'hc2093a05};
test_weights[27368:27375] = '{32'h42c14ec2, 32'h42b67d93, 32'h424290b9, 32'hc2a76e11, 32'hc21cd1de, 32'hc2ad70aa, 32'hc1d50736, 32'hc25ece3f};
test_bias[3421:3421] = '{32'h42ab5253};
test_output[3421:3421] = '{32'hc5a8f256};
test_input[27376:27383] = '{32'h41d1c4b4, 32'hc229c7bf, 32'hc29a8aae, 32'h42ad078c, 32'h42ab9417, 32'hc2109cfa, 32'h42184dfd, 32'h429c6fb4};
test_weights[27376:27383] = '{32'h428e7e1e, 32'hc252ff3c, 32'hc2938634, 32'hc25c1216, 32'h40cd07eb, 32'h42a72845, 32'h41caa74e, 32'h42c11e6f};
test_bias[3422:3422] = '{32'h4291bb04};
test_output[3422:3422] = '{32'h462e7432};
test_input[27384:27391] = '{32'h41f769f0, 32'h4256206a, 32'hc295893e, 32'hc28bb4f8, 32'hc1715f12, 32'h42633746, 32'h41fe35b5, 32'h428971f0};
test_weights[27384:27391] = '{32'h4213c237, 32'hc277fa40, 32'h41965481, 32'h40e89a62, 32'h4289f3e5, 32'h423b5576, 32'hc1e9d735, 32'hc1d5ccef};
test_bias[3423:3423] = '{32'h42b9a171};
test_output[3423:3423] = '{32'hc5a0aea4};
test_input[27392:27399] = '{32'h427f76df, 32'h421c7f9f, 32'h4241eeec, 32'h42357b32, 32'h41908c1c, 32'hc2be3ad3, 32'hc1d80063, 32'hc2430a2c};
test_weights[27392:27399] = '{32'hc2a76d29, 32'hc2a81e94, 32'hc2a343ee, 32'hc29aca19, 32'h420e879c, 32'h416d777f, 32'h423732ac, 32'hc1dde712};
test_bias[3424:3424] = '{32'hc07b513c};
test_output[3424:3424] = '{32'hc682f0b6};
test_input[27400:27407] = '{32'h4200bee4, 32'hbdfd841f, 32'h414190ce, 32'hc2b70c87, 32'h41c412c9, 32'hc2ac9a3d, 32'hc202e59f, 32'hc27c86b6};
test_weights[27400:27407] = '{32'h423693c0, 32'hc2c6e698, 32'hc2b03036, 32'h42733918, 32'hc275b965, 32'h42061836, 32'hc1e6f49d, 32'hc27311bd};
test_bias[3425:3425] = '{32'h42079de4};
test_output[3425:3425] = '{32'hc593ea83};
test_input[27408:27415] = '{32'h42570c19, 32'hc29fd914, 32'hc298b4ca, 32'h429e64ad, 32'hc2b9e089, 32'h42be8ada, 32'h42a10dc9, 32'hc296b56d};
test_weights[27408:27415] = '{32'hc2aec9c0, 32'h41d2aa05, 32'hc12e0795, 32'h426f96ca, 32'hc2b185c6, 32'hc0f351a0, 32'hc0e37d60, 32'hc2c289a9};
test_bias[3426:3426] = '{32'hc282f547};
test_output[3426:3426] = '{32'h464aee9c};
test_input[27416:27423] = '{32'hc21d4225, 32'hbf98d35d, 32'hc217f265, 32'h414b88df, 32'h408468f9, 32'hc29488c9, 32'hc227e44b, 32'h4272e12f};
test_weights[27416:27423] = '{32'hc28b6a0c, 32'hc0a901b9, 32'hc2590ae2, 32'h40edd316, 32'hc2ab9c92, 32'h424b3a67, 32'h42525c28, 32'hc21dfdf1};
test_bias[3427:3427] = '{32'h42979c40};
test_output[3427:3427] = '{32'hc56ababb};
test_input[27424:27431] = '{32'hc2bd3388, 32'h422d30d2, 32'h40dcbdeb, 32'hc02f138c, 32'hc0dcf26d, 32'hc241f1c1, 32'hc2c15252, 32'hc298b1f8};
test_weights[27424:27431] = '{32'hc24cb0ec, 32'hc1bed0f5, 32'h4105bd4b, 32'hc2a992a2, 32'hc2bd0147, 32'hc1597464, 32'hc1ce172c, 32'h414360d0};
test_bias[3428:3428] = '{32'hc233055b};
test_output[3428:3428] = '{32'h45d852fc};
test_input[27432:27439] = '{32'h424bc1b9, 32'h42925348, 32'h429d3695, 32'h41655f5d, 32'h42b05775, 32'hc25a10a6, 32'h421cf441, 32'h41c718c3};
test_weights[27432:27439] = '{32'h410aa448, 32'h422eeca3, 32'hc240a447, 32'hc17c3bff, 32'h4276ef7d, 32'h424cf11d, 32'hc2abc6b7, 32'hc2bf1ed4};
test_bias[3429:3429] = '{32'h4261aea7};
test_output[3429:3429] = '{32'hc5554cec};
test_input[27440:27447] = '{32'hc19ffef7, 32'hc2c5da5c, 32'h41be52c4, 32'h41754529, 32'hc1887ff7, 32'h42b15e92, 32'hc2a44d4e, 32'h4195efb1};
test_weights[27440:27447] = '{32'hc153469f, 32'hc1f7be30, 32'hc1ac80f9, 32'hc2bd08fc, 32'h4259cb84, 32'hc18e65d8, 32'hc2b9367e, 32'hc1fe0fcc};
test_bias[3430:3430] = '{32'hc29160c4};
test_output[3430:3430] = '{32'h45b52fb7};
test_input[27448:27455] = '{32'hc254ffd6, 32'hbf5fb243, 32'h424b3012, 32'h421cb38c, 32'h429541d1, 32'h42894982, 32'h42b599e3, 32'hc202accf};
test_weights[27448:27455] = '{32'hc246e97d, 32'hc2a6be4c, 32'hc27c0797, 32'hc2aea568, 32'h4214ab15, 32'hc2b4fe31, 32'hc16abac2, 32'hc18660c1};
test_bias[3431:3431] = '{32'hc28173ea};
test_output[3431:3431] = '{32'hc5ffd7ea};
test_input[27456:27463] = '{32'h42894479, 32'h41b3a850, 32'hc280bfb9, 32'hc26fb67a, 32'hc28dca99, 32'hc2ad5f47, 32'h42131eb0, 32'h422b4d80};
test_weights[27456:27463] = '{32'hc17db4b1, 32'hc1f64d84, 32'hc2b7d56f, 32'h4252ccb3, 32'h425039ea, 32'h420b69dd, 32'hc2c61c17, 32'h4286a11d};
test_bias[3432:3432] = '{32'hc1f752df};
test_output[3432:3432] = '{32'hc5cbe07f};
test_input[27464:27471] = '{32'hc23a6897, 32'hc29562b5, 32'h42897144, 32'hc21f7e1e, 32'h41a2c159, 32'hc2a86397, 32'h42bf802d, 32'hc24d1382};
test_weights[27464:27471] = '{32'hc29a8745, 32'hc11fe0a8, 32'hc20cbded, 32'hc28a83ad, 32'hc0ad007d, 32'h41a3b564, 32'hc27cac9d, 32'h42a98be7};
test_bias[3433:3433] = '{32'hc2911c5c};
test_output[3433:3433] = '{32'hc5edcc96};
test_input[27472:27479] = '{32'h42807187, 32'h42a1d79e, 32'h41ba12f5, 32'h42a10f6d, 32'hc21ec519, 32'hc1ce1289, 32'hc28363c5, 32'hc27353ce};
test_weights[27472:27479] = '{32'hc2946214, 32'h429075bd, 32'hc1fecbb5, 32'hc1f0f785, 32'h427ec68b, 32'hbfebc8b6, 32'hc28e65c1, 32'hc2a6f0bb};
test_bias[3434:3434] = '{32'h3ff9ae42};
test_output[3434:3434] = '{32'h45a23070};
test_input[27480:27487] = '{32'hc20027c5, 32'h428b9679, 32'hc223576f, 32'h42953263, 32'h421ea8fe, 32'hc2a91fb1, 32'hc257b533, 32'h424f13f2};
test_weights[27480:27487] = '{32'h42a16a88, 32'hc2bd199c, 32'h41a498e4, 32'hc280ccb7, 32'h41b0f74f, 32'hc1de5c68, 32'h42b272ca, 32'hc25bf5cc};
test_bias[3435:3435] = '{32'h416942d8};
test_output[3435:3435] = '{32'hc6965a30};
test_input[27488:27495] = '{32'h3fafdb85, 32'hc1b79c63, 32'hc2aacdf2, 32'hc1dbc2de, 32'hc02af538, 32'h425a8717, 32'h4229b003, 32'hc2b27933};
test_weights[27488:27495] = '{32'hc240c67f, 32'hc2240ce0, 32'h4272c4d0, 32'hc2bc911d, 32'hc2c79e1c, 32'hc29c48f2, 32'hc1c8fc27, 32'h42af83db};
test_bias[3436:3436] = '{32'h4236ef91};
test_output[3436:3436] = '{32'hc663af86};
test_input[27496:27503] = '{32'hc28f650a, 32'hc1fee91e, 32'h427b6a00, 32'h42c7e144, 32'h4257a3fb, 32'h41904769, 32'hc2b9ac31, 32'hc299fc62};
test_weights[27496:27503] = '{32'h42a1b5b2, 32'h416aae9c, 32'h4289c49b, 32'h4229de00, 32'h4122b208, 32'h420c380f, 32'h42c6e8ea, 32'h424bb5b0};
test_bias[3437:3437] = '{32'hc20c7dc7};
test_output[3437:3437] = '{32'hc6178e1a};
test_input[27504:27511] = '{32'hc19cf5af, 32'hc2a486e6, 32'h42c1f1a7, 32'h4232bade, 32'hc145be48, 32'hc23990bd, 32'hc260b058, 32'h4213315e};
test_weights[27504:27511] = '{32'hc2be5d0d, 32'h42c3cdf1, 32'hc1882d78, 32'hc16b525c, 32'h413e6f91, 32'h421803bd, 32'hc2ab5dfc, 32'hc22c9ccc};
test_bias[3438:3438] = '{32'hc2b6e466};
test_output[3438:3438] = '{32'hc5e33560};
test_input[27512:27519] = '{32'h42209757, 32'hc2252d61, 32'h422f85b7, 32'hc209f735, 32'h42901f7e, 32'hc2c12b58, 32'hc29ec5f3, 32'hc2b18a06};
test_weights[27512:27519] = '{32'hc23eb5eb, 32'h42aac497, 32'hc19ba68a, 32'h421f60d6, 32'hc225f479, 32'h41f3b317, 32'h41060c3a, 32'h423f6fac};
test_bias[3439:3439] = '{32'h42468833};
test_output[3439:3439] = '{32'hc6903fd5};
test_input[27520:27527] = '{32'h41c7370d, 32'h412e6e03, 32'h427f9dd5, 32'h41a2cc46, 32'hc1b9e9b1, 32'hc1f55173, 32'hc2c62992, 32'h42a46fed};
test_weights[27520:27527] = '{32'hc2c3d184, 32'hc2303aa9, 32'h428d2153, 32'hc13a7f61, 32'hc10e8f6f, 32'hc11d67d2, 32'hc29864ae, 32'hc286800f};
test_bias[3440:3440] = '{32'hc18fe037};
test_output[3440:3440] = '{32'h45718f7c};
test_input[27528:27535] = '{32'h42a22751, 32'hc203f4ed, 32'h421eab4f, 32'hc288ddbe, 32'hc297b818, 32'h41d1ab0a, 32'h4141bc6d, 32'h4298e58c};
test_weights[27528:27535] = '{32'h42bfd027, 32'hc2bb685b, 32'h422489c7, 32'hc2766f15, 32'h3fa23219, 32'h428d988e, 32'hc10e52dd, 32'h42c06ca7};
test_bias[3441:3441] = '{32'h4290ef90};
test_output[3441:3441] = '{32'h46c98456};
test_input[27536:27543] = '{32'hc296c534, 32'hc22b18a6, 32'hc2b5dd97, 32'h422d9e3d, 32'hc1cbc815, 32'hc01fbbe7, 32'hc203b7d2, 32'h42a5e792};
test_weights[27536:27543] = '{32'h41bc4e69, 32'hc2033994, 32'hc10adaf2, 32'hc15f0977, 32'hc22e6d9e, 32'hc24b7544, 32'hc28b67e5, 32'hc2c692b9};
test_bias[3442:3442] = '{32'hc27b007c};
test_output[3442:3442] = '{32'hc59ac6d1};
test_input[27544:27551] = '{32'h42044110, 32'h42152a4b, 32'h415145d2, 32'h42c2f041, 32'hc2c13f23, 32'hc1a2c737, 32'h41b04e98, 32'h41aee0e4};
test_weights[27544:27551] = '{32'hc291e233, 32'h42a19090, 32'hbf6c7052, 32'h42c4c957, 32'hc14a995f, 32'hc240a991, 32'h4200010f, 32'h42a49f35};
test_bias[3443:3443] = '{32'hc226f6da};
test_output[3443:3443] = '{32'h4667f559};
test_input[27552:27559] = '{32'hc282f723, 32'h42ab7474, 32'hc02fa738, 32'h42935f30, 32'hc1801fd7, 32'hc104aee0, 32'h4285eee5, 32'h42b56b27};
test_weights[27552:27559] = '{32'h42834999, 32'hc1ab7d3e, 32'h429c9b72, 32'hc20a2268, 32'h4187b522, 32'h42c032ad, 32'hc0ed7865, 32'h418ce8c6};
test_bias[3444:3444] = '{32'hc29bff50};
test_output[3444:3444] = '{32'hc60bb64e};
test_input[27560:27567] = '{32'hc29d2024, 32'hc280c6c5, 32'h424d365b, 32'h40aa61d3, 32'hc1b38dca, 32'hc1f62f68, 32'hc20d3b6d, 32'hc00cb4f6};
test_weights[27560:27567] = '{32'hc271fb1f, 32'h41b7e267, 32'hc282a347, 32'h421eaa9d, 32'h42a13f85, 32'hc24a693a, 32'h427dff13, 32'h42bc87a3};
test_bias[3445:3445] = '{32'h424c94e9};
test_output[3445:3445] = '{32'hc51d5a69};
test_input[27568:27575] = '{32'h42b90809, 32'hc228ac56, 32'h4289f665, 32'hc27e8f3d, 32'h42752814, 32'h425de126, 32'h423246a0, 32'hc2af2ae2};
test_weights[27568:27575] = '{32'h42908175, 32'h42b6a584, 32'hc1bf30c4, 32'hc17a5dd6, 32'h42bf0e81, 32'h412e6dba, 32'hbf0bf156, 32'h4200b27f};
test_bias[3446:3446] = '{32'h42517f4a};
test_output[3446:3446] = '{32'h45b6d3c2};
test_input[27576:27583] = '{32'hc290d3f1, 32'hc1d9d640, 32'h4226a72e, 32'hc29f4dc7, 32'h3f602751, 32'hc25c1192, 32'hc2b6d1aa, 32'h421769fa};
test_weights[27576:27583] = '{32'hc2ac0a09, 32'hc2a7e18b, 32'h42838056, 32'hc280b6df, 32'h42aed2e5, 32'h4007e99c, 32'hc1beffe3, 32'hc12ed129};
test_bias[3447:3447] = '{32'hc1602b49};
test_output[3447:3447] = '{32'h468d5d7c};
test_input[27584:27591] = '{32'h42b88bf8, 32'h41f12f31, 32'hc27e80e6, 32'h42522888, 32'h41d8ed90, 32'hbf966247, 32'hc1684782, 32'hc216c4e6};
test_weights[27584:27591] = '{32'h411b19f0, 32'h417ab534, 32'h41fd9d96, 32'h42b46873, 32'h42381075, 32'hc1045095, 32'h4130e010, 32'hc1813e7a};
test_bias[3448:3448] = '{32'hc2c1631b};
test_output[3448:3448] = '{32'h45b212bc};
test_input[27592:27599] = '{32'hc18bc228, 32'h429b341b, 32'hc27387cb, 32'h41ca23ec, 32'h426fc0e7, 32'h4225433c, 32'hc28a58dd, 32'h419dcb2a};
test_weights[27592:27599] = '{32'h40d12684, 32'hc1cf17d1, 32'hc2b2a1b8, 32'hc2529959, 32'hc2ab3b5a, 32'h42a2ca75, 32'hc1ea13bb, 32'hc1e63272};
test_bias[3449:3449] = '{32'hc120733a};
test_output[3449:3449] = '{32'h44cfc1d0};
test_input[27600:27607] = '{32'hc1a1347d, 32'hc2a874db, 32'hc245fe24, 32'h42afd524, 32'h42901845, 32'h41c42530, 32'h4195fc97, 32'h42b163b5};
test_weights[27600:27607] = '{32'h418dc8ca, 32'h42339981, 32'h4291f082, 32'h4225b6e6, 32'hc262227a, 32'h40f84f6d, 32'h420f4ab1, 32'h42aa90c6};
test_bias[3450:3450] = '{32'hc1dee0bb};
test_output[3450:3450] = '{32'h435873df};
test_input[27608:27615] = '{32'h41775f1a, 32'hc216ab42, 32'hc1a290c9, 32'h41d94a5f, 32'hc2013253, 32'h4236f472, 32'h42023507, 32'h429a9f62};
test_weights[27608:27615] = '{32'hc20126c5, 32'hc2a8dadc, 32'h42be79fd, 32'hc2bb3835, 32'hc228f131, 32'h4294f297, 32'hc0a319f2, 32'hc2127a14};
test_bias[3451:3451] = '{32'hc21176da};
test_output[3451:3451] = '{32'hc26f1190};
test_input[27616:27623] = '{32'hc25da5cc, 32'hc242b81e, 32'h42564862, 32'hc2427411, 32'hc2893d4a, 32'hc2c7b9c6, 32'h425a2835, 32'hc2a925c1};
test_weights[27616:27623] = '{32'h418a6d12, 32'h42bb9b88, 32'hc2470686, 32'hc2939d19, 32'h419c1621, 32'hc2971500, 32'hc2c0c0a0, 32'h422c7a33};
test_bias[3452:3452] = '{32'hc205974d};
test_output[3452:3452] = '{32'hc5e53168};
test_input[27624:27631] = '{32'hc20f95b4, 32'hc28f58df, 32'h41b5ca8f, 32'hc22a4a01, 32'h419ce881, 32'h405cd878, 32'hc275d533, 32'hc29eb9ae};
test_weights[27624:27631] = '{32'hc22da992, 32'hc01e9b94, 32'h4051a064, 32'h4257ec4b, 32'h41ecb5e7, 32'hbf9c74fd, 32'h42b37120, 32'hc280353d};
test_bias[3453:3453] = '{32'h42160d0c};
test_output[3453:3453] = '{32'hc396480d};
test_input[27632:27639] = '{32'h42c70abd, 32'hc28f8100, 32'h426f7119, 32'h40df8a21, 32'hc1d347df, 32'h42a869c6, 32'h42123b0f, 32'h41e0aae8};
test_weights[27632:27639] = '{32'h418780e2, 32'h41aa403e, 32'hc236cb4e, 32'h42bb27d9, 32'h429465cd, 32'h425facbe, 32'hc1ca7d78, 32'h42418e94};
test_bias[3454:3454] = '{32'hc2a0bc00};
test_output[3454:3454] = '{32'h4493678b};
test_input[27640:27647] = '{32'hc1d49cc9, 32'hc2c79d50, 32'h4222e45d, 32'h42a1e709, 32'h42c43d6b, 32'h42a5c754, 32'h401d0bf6, 32'hc1755509};
test_weights[27640:27647] = '{32'hc2aa0d96, 32'hc2892b92, 32'h429b9811, 32'hc1c97f95, 32'h3ee7ef4b, 32'hc24b9620, 32'hc2b6feca, 32'hc1a48b5f};
test_bias[3455:3455] = '{32'h423d8c00};
test_output[3455:3455] = '{32'h45c1b0bc};
test_input[27648:27655] = '{32'hc1d3adb3, 32'h421e9b45, 32'h3ea04401, 32'h42b57cba, 32'h42bee4d9, 32'h423171e3, 32'h42a11a35, 32'hc1aaa6d7};
test_weights[27648:27655] = '{32'h42be596c, 32'h41c9fca2, 32'hc0ba8e29, 32'hc276bee4, 32'h41f3f4b5, 32'h42aaafd3, 32'hc243c7a1, 32'hc0168b85};
test_bias[3456:3456] = '{32'h4282d487};
test_output[3456:3456] = '{32'hc584b89b};
test_input[27656:27663] = '{32'hc289ac70, 32'h4268c1e0, 32'hc236002b, 32'hc284817d, 32'hc297a00c, 32'hc1dd3458, 32'hc20251a7, 32'h4148d962};
test_weights[27656:27663] = '{32'hc28b2b75, 32'hc1e9aafc, 32'hc2a477da, 32'h420d22c8, 32'h42abaf4f, 32'h41eadeb1, 32'hc22ee5c6, 32'h42bdda53};
test_bias[3457:3457] = '{32'hc212452c};
test_output[3457:3457] = '{32'hc375c3a8};
test_input[27664:27671] = '{32'h427d4fec, 32'h42bee59a, 32'hc13067cf, 32'h424d043d, 32'h42ae9ce0, 32'hc2331240, 32'hc19f09fe, 32'h420056d8};
test_weights[27664:27671] = '{32'h428b33ec, 32'h41a596b8, 32'h4298d94d, 32'h410cc72f, 32'hc1c91667, 32'h4224d607, 32'h425e4c08, 32'h423f3dac};
test_bias[3458:3458] = '{32'h428f9ec9};
test_output[3458:3458] = '{32'h4519558f};
test_input[27672:27679] = '{32'hc092af33, 32'hc2377746, 32'hc2bf6650, 32'hc2c3588c, 32'h42a6b699, 32'h42add0b2, 32'hc1dd5d9b, 32'hc24cb6b3};
test_weights[27672:27679] = '{32'h41fe5b07, 32'hc22deb5c, 32'h42a15c16, 32'h41b0f00a, 32'hc29debbf, 32'hc170e04c, 32'hc14e0b18, 32'h41494a0e};
test_bias[3459:3459] = '{32'h41b8d133};
test_output[3459:3459] = '{32'hc67cedc5};
test_input[27680:27687] = '{32'h423dfb76, 32'hc191cfa7, 32'h423484dd, 32'h42b48e01, 32'hc27f105c, 32'hc226e1a8, 32'h4298261d, 32'h4268b010};
test_weights[27680:27687] = '{32'hc2994999, 32'h42557c20, 32'hc2466a1c, 32'hc246a411, 32'hc2775471, 32'h428dbb64, 32'h41409a79, 32'h42bc6bba};
test_bias[3460:3460] = '{32'hc0b2e902};
test_output[3460:3460] = '{32'hc5775f86};
test_input[27688:27695] = '{32'hc16f645b, 32'h421fa0ad, 32'h42c7aca0, 32'h429e8c49, 32'hc28d5733, 32'h42c115af, 32'h420c9cb8, 32'hc16212b9};
test_weights[27688:27695] = '{32'hc1ce6003, 32'h3f368217, 32'h42bfbdfc, 32'hc1b0e606, 32'h420fb071, 32'h42ac291a, 32'h4266e376, 32'hc245ddae};
test_bias[3461:3461] = '{32'h41a2fdea};
test_output[3461:3461] = '{32'h4682e252};
test_input[27696:27703] = '{32'hc2af5c8c, 32'h41a33ea2, 32'hc17d1300, 32'h421ee68c, 32'h40f5bc40, 32'hc263643d, 32'h427d266f, 32'h4228d4a9};
test_weights[27696:27703] = '{32'h42744c0c, 32'hc240853c, 32'h428bdfbf, 32'h429c1ccf, 32'h417e76f0, 32'hc26866e6, 32'h41baeea0, 32'h42a5c382};
test_bias[3462:3462] = '{32'h428e9225};
test_output[3462:3462] = '{32'h45811662};
test_input[27704:27711] = '{32'h41b8a218, 32'hc2963636, 32'h425f5358, 32'h40d3f40a, 32'hc29616eb, 32'h42575c27, 32'h422aa088, 32'hc19a7c59};
test_weights[27704:27711] = '{32'h41a049c2, 32'h419c04b7, 32'h42c0a1d2, 32'hc28dacdd, 32'hc154d29e, 32'hc28e50fc, 32'hc028cbc9, 32'h41b4fc8d};
test_bias[3463:3463] = '{32'hc2bd3ac6};
test_output[3463:3463] = '{32'h43d67f50};
test_input[27712:27719] = '{32'h40960117, 32'hc295f2e1, 32'hc28728b3, 32'h424dbcb8, 32'hc25f1c8a, 32'h42407842, 32'h42321974, 32'hc17819db};
test_weights[27712:27719] = '{32'hc205b211, 32'h42771f27, 32'h41865def, 32'hc1185707, 32'h425a7a48, 32'hc23d31e3, 32'hc0865127, 32'hc2770349};
test_bias[3464:3464] = '{32'hc2003bc5};
test_output[3464:3464] = '{32'hc62bd4ef};
test_input[27720:27727] = '{32'hc2b46249, 32'h42089ea5, 32'h4243d7e6, 32'h42c35e67, 32'h42c052d8, 32'h41135621, 32'h4242d972, 32'hc285a1e6};
test_weights[27720:27727] = '{32'h42984cf7, 32'h42037bbb, 32'hc2abc15b, 32'h41bb6fb3, 32'h41a275c8, 32'hc298cb8e, 32'hc287f2d2, 32'hc1863d9e};
test_bias[3465:3465] = '{32'hc2b3a639};
test_output[3465:3465] = '{32'hc607cfac};
test_input[27728:27735] = '{32'h427309be, 32'h41b7648c, 32'h4183b143, 32'h42c28efc, 32'h41d76acb, 32'hc2c5e6ab, 32'h41c0d42c, 32'hc2b4bdee};
test_weights[27728:27735] = '{32'hc247869d, 32'h40075401, 32'h42477934, 32'h4275e162, 32'h41a6880f, 32'hc1c205af, 32'hc2b0ddb7, 32'h42087084};
test_bias[3466:3466] = '{32'hc1c90258};
test_output[3466:3466] = '{32'h44c0702d};
test_input[27736:27743] = '{32'h4212f6f4, 32'h41d2c586, 32'h4086acb9, 32'h41e3c2ef, 32'hbf7279e7, 32'hc1da37d2, 32'hc2991126, 32'h4284ceb0};
test_weights[27736:27743] = '{32'h41c6f759, 32'h42bdd3a6, 32'h42b113b6, 32'hc2b18c6a, 32'hc277dd6a, 32'hc2a34d5b, 32'h4280112e, 32'h42c14b77};
test_bias[3467:3467] = '{32'h415e1719};
test_output[3467:3467] = '{32'h459ea37e};
test_input[27744:27751] = '{32'h41b02823, 32'h42162a17, 32'hc1e5a825, 32'hc246ce18, 32'h42c170bd, 32'hc28a8ba2, 32'h4284f5d5, 32'hc27ef1ee};
test_weights[27744:27751] = '{32'h42331453, 32'hc0946995, 32'h403a2b92, 32'h4239ec78, 32'hc2bdfe28, 32'h42990f4e, 32'h427a4a73, 32'hc2b6c457};
test_bias[3468:3468] = '{32'hc27a99df};
test_output[3468:3468] = '{32'hc5c02eaf};
test_input[27752:27759] = '{32'hc1ac8304, 32'hc1b2e4c6, 32'hc20240b8, 32'h4166bbe6, 32'hc22f4994, 32'hc28dafa3, 32'h413aad4d, 32'hc2011530};
test_weights[27752:27759] = '{32'h42187418, 32'h42739290, 32'hc231c6cc, 32'h428abdfa, 32'h41d343f7, 32'h42608a11, 32'h42a3d5d2, 32'h41ba4573};
test_bias[3469:3469] = '{32'h4276ab19};
test_output[3469:3469] = '{32'hc58fdf2a};
test_input[27760:27767] = '{32'hc28bace3, 32'hc1f6ac68, 32'h4263af98, 32'h42b9cfcd, 32'h4296fa00, 32'hc2a691dc, 32'h42c304ef, 32'h42959892};
test_weights[27760:27767] = '{32'hc25d0010, 32'h4246124f, 32'hc2a4a79c, 32'h4255bc72, 32'hc2945355, 32'h42b4021f, 32'hc26e70d9, 32'hc20a4006};
test_bias[3470:3470] = '{32'hc0c37b46};
test_output[3470:3470] = '{32'hc69390ea};
test_input[27768:27775] = '{32'hc283dd0e, 32'hc123ff04, 32'h418a5d43, 32'h4253461c, 32'hc20a77cd, 32'hc1737c98, 32'hc28fdfcd, 32'hc2aad02c};
test_weights[27768:27775] = '{32'hc278176f, 32'h42817ccb, 32'h428d7d30, 32'hc285c4cf, 32'hc2c5f7a7, 32'hc2c21d7a, 32'hc0177660, 32'hc1e285d0};
test_bias[3471:3471] = '{32'hc24a2a8d};
test_output[3471:3471] = '{32'h4605b839};
test_input[27776:27783] = '{32'hc1b4dd33, 32'h3cec6017, 32'hc2937040, 32'hc26e8978, 32'h429f6414, 32'h4191833d, 32'hc2af8848, 32'hc2752619};
test_weights[27776:27783] = '{32'h41c766ed, 32'hc29736fd, 32'h415057d5, 32'h421b91c1, 32'hc241e3ef, 32'hc213a6f6, 32'h421d798f, 32'h41a9a62f};
test_bias[3472:3472] = '{32'h420975df};
test_output[3472:3472] = '{32'hc64cafc2};
test_input[27784:27791] = '{32'h42b4263c, 32'h4233641d, 32'h425e5aee, 32'hc1937a09, 32'hc05250db, 32'h425d9ec4, 32'hc2a64527, 32'h42674c7f};
test_weights[27784:27791] = '{32'hc2c55334, 32'hc27f032b, 32'hc1ccbb68, 32'h424431a6, 32'h3f6d78a7, 32'hc103267e, 32'h4102a86a, 32'h42a0e042};
test_bias[3473:3473] = '{32'h42a690df};
test_output[3473:3473] = '{32'hc623a9e0};
test_input[27792:27799] = '{32'hc08d0e1f, 32'hc2997122, 32'hc26f2374, 32'hc23ebc56, 32'hc2633276, 32'h428c7f66, 32'hc1758b12, 32'hc11f1e8f};
test_weights[27792:27799] = '{32'h42c272cb, 32'hc2b4d73c, 32'h425444e3, 32'hc21dbfb0, 32'h42791ce1, 32'h4296cf93, 32'h42a70ade, 32'hc258444d};
test_bias[3474:3474] = '{32'hc13c7e7b};
test_output[3474:3474] = '{32'h45c26372};
test_input[27800:27807] = '{32'h4242725f, 32'h411fb2b0, 32'hc27be735, 32'h409626bb, 32'hc2ad12fa, 32'hc29c9935, 32'h426e4e2b, 32'h40e503b0};
test_weights[27800:27807] = '{32'hc1003181, 32'hc2ada341, 32'hc2798ccd, 32'h42937367, 32'h42503c4d, 32'hc2212daf, 32'h42839499, 32'h42c18405};
test_bias[3475:3475] = '{32'h4244805d};
test_output[3475:3475] = '{32'h45c5cfa3};
test_input[27808:27815] = '{32'hc2c53102, 32'h414df8ad, 32'h41bb66fd, 32'hc2b2253c, 32'h41e348ac, 32'hc262ac52, 32'h421658d6, 32'h426b3ca9};
test_weights[27808:27815] = '{32'h42567272, 32'hc236feb2, 32'hc26e54a4, 32'hc24cd524, 32'hc2c5e19b, 32'hc1bfe446, 32'hc1920056, 32'h41ae8347};
test_bias[3476:3476] = '{32'hc1de567e};
test_output[3476:3476] = '{32'hc5607e19};
test_input[27816:27823] = '{32'h42b8557c, 32'hc209868d, 32'h41a0d286, 32'h410f4b49, 32'hc00c3e5a, 32'hc274b7dd, 32'h416410ca, 32'hc1ebea68};
test_weights[27816:27823] = '{32'hc2026e24, 32'h41f2902c, 32'hc2557f3c, 32'h41f3bd5e, 32'h40dca649, 32'hc21e4c55, 32'hc1f1888a, 32'hc2c47270};
test_bias[3477:3477] = '{32'h42286386};
test_output[3477:3477] = '{32'h4284dfc9};
test_input[27824:27831] = '{32'hc24ab115, 32'hc0947710, 32'hc2a1f01b, 32'hc014b74f, 32'hc20962c7, 32'h42c177f7, 32'hc189e763, 32'hc21ebc55};
test_weights[27824:27831] = '{32'h406908ef, 32'hc2bdcc07, 32'hc2bd9988, 32'h42b85989, 32'hc2b2b9bd, 32'hc263a02c, 32'hc2652e7c, 32'h42924385};
test_bias[3478:3478] = '{32'h4225661e};
test_output[3478:3478] = '{32'h45550c69};
test_input[27832:27839] = '{32'hc272ebde, 32'hbfc74648, 32'hc22ebe3a, 32'h425e483e, 32'h42aba94c, 32'h428733b4, 32'hc2b37aea, 32'hc14bf0b9};
test_weights[27832:27839] = '{32'hc218d974, 32'h423754f6, 32'hc250a6ea, 32'h422ec820, 32'h41c086fc, 32'hc2006dcf, 32'hc27d8078, 32'h427366b3};
test_bias[3479:3479] = '{32'h42a2b628};
test_output[3479:3479] = '{32'h463911b5};
test_input[27840:27847] = '{32'hc2c0fe87, 32'hc21ffa94, 32'h42911484, 32'hc2970201, 32'h42b0d446, 32'hc2c74e74, 32'hc2ac9a28, 32'hc1f79933};
test_weights[27840:27847] = '{32'hc2567130, 32'h414bbe3a, 32'h4268d43e, 32'hc2184e29, 32'h424336e4, 32'hc2c2b258, 32'hc21fe947, 32'hc2723144};
test_bias[3480:3480] = '{32'h42c59dc2};
test_output[3480:3480] = '{32'h46f3c051};
test_input[27848:27855] = '{32'h429ae68b, 32'hc205a071, 32'h42b4d998, 32'hc202da5e, 32'hc295b00d, 32'hc0e31d08, 32'h423c68f1, 32'hc12947ba};
test_weights[27848:27855] = '{32'h420d634e, 32'h4276d7fc, 32'hc2a92e4d, 32'hc1c5341e, 32'h42765bc5, 32'hc2c6b6a4, 32'hc22f24ec, 32'h42b4d52b};
test_bias[3481:3481] = '{32'hc263beeb};
test_output[3481:3481] = '{32'hc64d6c1f};
test_input[27856:27863] = '{32'h42c43cdc, 32'hc2a67c01, 32'hc295bcb7, 32'h425bdead, 32'h41a3bbfd, 32'hc2747721, 32'h42ab1bc8, 32'hbf5c4b1d};
test_weights[27856:27863] = '{32'hc21280f1, 32'h41272721, 32'hc188e5ab, 32'hc2b00d64, 32'hc23312b4, 32'h420beee0, 32'hc14bf03d, 32'hc206a0ba};
test_bias[3482:3482] = '{32'hc1908136};
test_output[3482:3482] = '{32'hc63dea91};
test_input[27864:27871] = '{32'h4280f5dd, 32'hc228cbce, 32'hc0abd95c, 32'h403a44af, 32'hc2924746, 32'hc25cbcf9, 32'hc1c55b7b, 32'hc26ce4fb};
test_weights[27864:27871] = '{32'hc2b0199b, 32'h419fa6b0, 32'h42208dda, 32'h41a5f472, 32'hc24d10d6, 32'h42b12115, 32'hc22d41cc, 32'h423b2c0c};
test_bias[3483:3483] = '{32'h424d9df7};
test_output[3483:3483] = '{32'hc613dfa6};
test_input[27872:27879] = '{32'hc142a002, 32'hbfb31f0a, 32'hc293dce0, 32'hc2c358b3, 32'hc1a95a69, 32'hc28e1937, 32'h42b0dbdf, 32'h422c54bc};
test_weights[27872:27879] = '{32'h428c20d1, 32'hc22a1dc5, 32'hc28222e2, 32'h420a2149, 32'hc2931880, 32'h4250ccb3, 32'h4240384e, 32'h42a2ad2d};
test_bias[3484:3484] = '{32'hc12b3bd9};
test_output[3484:3484] = '{32'h45c2e13e};
test_input[27880:27887] = '{32'hc175867d, 32'h41af6f3f, 32'h3f1d4ef0, 32'hc0252ae8, 32'hc238f791, 32'h42be09e5, 32'hc2790181, 32'hc29f86a9};
test_weights[27880:27887] = '{32'hc25c0ce9, 32'hc2bb3c6a, 32'hc14ff910, 32'hc21bd3f6, 32'h42bf8b4f, 32'h4284f80a, 32'hc1e22bcf, 32'hc197fcbf};
test_bias[3485:3485] = '{32'hc2a021cb};
test_output[3485:3485] = '{32'h4577fa2e};
test_input[27888:27895] = '{32'h41a1cc12, 32'hc25201ae, 32'hc29bb649, 32'hc2c47076, 32'h41a030fd, 32'hc1622808, 32'hc2a362e4, 32'hc298d33a};
test_weights[27888:27895] = '{32'hc27eb7fb, 32'hc2c5c096, 32'h427f2f29, 32'h420d191e, 32'h42947508, 32'hc24844a7, 32'h42c33b2f, 32'h427d65dd};
test_bias[3486:3486] = '{32'h42b48321};
test_output[3486:3486] = '{32'hc66b4cea};
test_input[27896:27903] = '{32'hc25dc909, 32'hc286f3f7, 32'hc2afa015, 32'h41407186, 32'hc18ec032, 32'h4269b172, 32'h428d13e3, 32'hc20c5444};
test_weights[27896:27903] = '{32'h4272e9db, 32'h41fc34c7, 32'h4277395b, 32'hc197cf63, 32'h40d35721, 32'h41fee6b2, 32'hc29d6b2d, 32'h42c0a51f};
test_bias[3487:3487] = '{32'hc28ff431};
test_output[3487:3487] = '{32'hc68fd32d};
test_input[27904:27911] = '{32'h42550e1f, 32'hc275b743, 32'h4279ef36, 32'hc2bb7bba, 32'h420e6293, 32'hc299baf3, 32'hc20baead, 32'hc1cf79b7};
test_weights[27904:27911] = '{32'hc118658e, 32'hc1957db4, 32'hc2aedaa8, 32'h42bdcc9f, 32'hc24833e7, 32'h4263256b, 32'hc2b75d47, 32'hc211ae81};
test_bias[3488:3488] = '{32'hc2340eb5};
test_output[3488:3488] = '{32'hc6764e99};
test_input[27912:27919] = '{32'hc28290b1, 32'h424e031f, 32'hc239389a, 32'hc224350c, 32'hc23ed59c, 32'hc20b6dd7, 32'h421197e3, 32'h42a4b145};
test_weights[27912:27919] = '{32'h42186a77, 32'hc28f6845, 32'hc1f5f336, 32'hc14672b9, 32'h42a9a4bb, 32'h42b20fc9, 32'hc28c1718, 32'h416736a4};
test_bias[3489:3489] = '{32'h42a8cb3c};
test_output[3489:3489] = '{32'hc64603e3};
test_input[27920:27927] = '{32'h42a0ebaf, 32'hc1e722a6, 32'hc16ae6ff, 32'h42106385, 32'hc22784a6, 32'hc1f515b9, 32'hc2530b03, 32'hc2a193bd};
test_weights[27920:27927] = '{32'hc0b1b9a6, 32'h417c75d3, 32'h41e00f97, 32'h423987a6, 32'h42082a08, 32'hc111a25a, 32'h428090a1, 32'h4282ec0f};
test_bias[3490:3490] = '{32'h42c0bf72};
test_output[3490:3490] = '{32'hc61268a2};
test_input[27928:27935] = '{32'h426e45df, 32'hc29882f1, 32'hc242e862, 32'hc231926a, 32'h4139bb10, 32'hc26899b0, 32'hc2c03266, 32'h41c4715a};
test_weights[27928:27935] = '{32'h42b15ef2, 32'hc26ea0cb, 32'h42c2137c, 32'hc2a9ad57, 32'h41cabfc3, 32'hc2887db9, 32'hc2aa894b, 32'h425d6f54};
test_bias[3491:3491] = '{32'hc2c38e44};
test_output[3491:3491] = '{32'h46b07891};
test_input[27936:27943] = '{32'hc0b7995e, 32'hc1391231, 32'h41c59e28, 32'h416708fd, 32'hc26eb84e, 32'hc1c15c6a, 32'hc1e68d17, 32'hc1b69dca};
test_weights[27936:27943] = '{32'hc2370403, 32'h42a291a5, 32'h4266953f, 32'hc2b82e24, 32'hc21fec33, 32'h4276337c, 32'hc2750490, 32'h40e659ab};
test_bias[3492:3492] = '{32'h40a7fa54};
test_output[3492:3492] = '{32'h44f02371};
test_input[27944:27951] = '{32'hbeb4249d, 32'hc18130c4, 32'hc1d6953f, 32'h4285994f, 32'h422d7bcf, 32'h42afdcd2, 32'hc2412fe7, 32'h419f0fb6};
test_weights[27944:27951] = '{32'h422ac270, 32'hc2a92b1c, 32'hc0c2aa98, 32'h420c8463, 32'hc18a9d92, 32'h417832f5, 32'h4225b703, 32'h4178edf5};
test_bias[3493:3493] = '{32'h4283bd82};
test_output[3493:3493] = '{32'h4531f944};
test_input[27952:27959] = '{32'h41c97ef9, 32'hc2376789, 32'hc237b483, 32'hc26b7c82, 32'hc289846e, 32'h42ab8f9a, 32'hc238696d, 32'hc2063692};
test_weights[27952:27959] = '{32'h42c19ae1, 32'h41858535, 32'h41e93801, 32'hc2451406, 32'hc1f10237, 32'h40b220cb, 32'h4200cfd1, 32'hc1555f3b};
test_bias[3494:3494] = '{32'hc1c93d99};
test_output[3494:3494] = '{32'h459389a1};
test_input[27960:27967] = '{32'hc20a2145, 32'hc1c75cb1, 32'hc2412620, 32'h415f4625, 32'hc12cdde0, 32'hc112ef79, 32'h42440df8, 32'hc2a42d5b};
test_weights[27960:27967] = '{32'h4074c8f4, 32'hc2c5f7f1, 32'h427ad750, 32'h414c0c1a, 32'h40d7cfb8, 32'hc294ebaa, 32'hc13247e3, 32'h41d77325};
test_bias[3495:3495] = '{32'hc220ed5a};
test_output[3495:3495] = '{32'hc528daef};
test_input[27968:27975] = '{32'hc29c1db2, 32'h41a5842e, 32'hc2a46f5c, 32'h4250d5c1, 32'hc1441047, 32'hc2748ae4, 32'h42c24cc9, 32'h428530cf};
test_weights[27968:27975] = '{32'h42b4bfcf, 32'hc19d55c7, 32'h42ad96d6, 32'hc28235b5, 32'hc285939c, 32'hc2c6f9cc, 32'hc2bf62c2, 32'h40bbe45d};
test_bias[3496:3496] = '{32'h41d6fc2d};
test_output[3496:3496] = '{32'hc69c0cdc};
test_input[27976:27983] = '{32'hc2a5edbf, 32'h4240ade4, 32'hc2003879, 32'hc2b958f3, 32'h4273ce5f, 32'hc2b804e0, 32'hc28a6051, 32'hc243f13a};
test_weights[27976:27983] = '{32'hc2237f2d, 32'hc01d13aa, 32'hc2874cc4, 32'h4114dd52, 32'h41f0bb85, 32'h41c5b771, 32'hc1f58f71, 32'h4290cfa8};
test_bias[3497:3497] = '{32'h411830fd};
test_output[3497:3497] = '{32'h452a5bb7};
test_input[27984:27991] = '{32'h42027883, 32'hc26c4e84, 32'hc10e31d9, 32'hc26760da, 32'h4214e726, 32'h41a07b35, 32'h423487f7, 32'hc1d09435};
test_weights[27984:27991] = '{32'hc28f1ff9, 32'h42492e8d, 32'h40ad085b, 32'hc2517573, 32'hc2b8bd3a, 32'hc20bc062, 32'h41ddd875, 32'h42087e20};
test_bias[3498:3498] = '{32'h4262a49d};
test_output[3498:3498] = '{32'hc5bceae9};
test_input[27992:27999] = '{32'hc2816beb, 32'hc2a3af6e, 32'hc2417c5a, 32'h4113d0b1, 32'hc03dc120, 32'h41384d65, 32'h42636cc2, 32'hc1c8d93d};
test_weights[27992:27999] = '{32'h42808a23, 32'hc1bd4024, 32'h42ad21a6, 32'hc2ad0fa0, 32'h41fa85a8, 32'h42b2f219, 32'h42772332, 32'h4284cabe};
test_bias[3499:3499] = '{32'h42814ef2};
test_output[3499:3499] = '{32'hc5884a02};
test_input[28000:28007] = '{32'hc146529c, 32'hc2b03f24, 32'h4092dcf0, 32'hc280c048, 32'h42c69ebb, 32'hc247a6b6, 32'h3e5a8e41, 32'hc24c16e0};
test_weights[28000:28007] = '{32'h42c5199d, 32'hc2819fcd, 32'hc259754f, 32'hc252e8eb, 32'hc1f581e5, 32'hc1cff0b5, 32'h419c17c8, 32'h4152c41a};
test_bias[3500:3500] = '{32'hc2a99deb};
test_output[3500:3500] = '{32'h45a05da6};
test_input[28008:28015] = '{32'hc2c76232, 32'h421e07b1, 32'hc2aac5cf, 32'h4206691a, 32'hc1c1c380, 32'hc2057589, 32'h41ade5ca, 32'hc23a00aa};
test_weights[28008:28015] = '{32'h4230fe3b, 32'h41e6dba9, 32'h417dd1b1, 32'hc2b2f05c, 32'h42c0f9c4, 32'h41048ffe, 32'hc29f1a9e, 32'h4286b2ce};
test_bias[3501:3501] = '{32'hc12c70bf};
test_output[3501:3501] = '{32'hc66c3518};
test_input[28016:28023] = '{32'h4252c197, 32'h42c33b37, 32'hc21a00f4, 32'h425a1306, 32'hc24dfd23, 32'h42860e11, 32'h42aa498a, 32'hc2b364aa};
test_weights[28016:28023] = '{32'h427ebf27, 32'h42c29efa, 32'hc263903d, 32'h40ec0d44, 32'h409c960c, 32'hc285f1bc, 32'hc21054f5, 32'h419f0a7a};
test_bias[3502:3502] = '{32'h4211b58f};
test_output[3502:3502] = '{32'h45b7f971};
test_input[28024:28031] = '{32'h4275072c, 32'h419b2b1d, 32'hc2b0df1d, 32'hc28b25a9, 32'h42569549, 32'hc296c744, 32'hc202fb2f, 32'hc17f288a};
test_weights[28024:28031] = '{32'h3f00c6de, 32'hc2c4b0cb, 32'hc2159ef1, 32'hc2a69021, 32'hc2a208b5, 32'hc292c963, 32'hc175cfcb, 32'h42857931};
test_bias[3503:3503] = '{32'h42ac53f2};
test_output[3503:3503] = '{32'h45f80a0f};
test_input[28032:28039] = '{32'hc297a251, 32'h4233885d, 32'h428a8d7e, 32'h421cf587, 32'h428649e6, 32'hc1bb518d, 32'hbe871700, 32'hc2c336b0};
test_weights[28032:28039] = '{32'hc1d4061a, 32'hc2a4d90b, 32'h42b9f728, 32'h4294a6bf, 32'h4159ef01, 32'hc2afe502, 32'hc296dbf5, 32'h4246dd13};
test_bias[3504:3504] = '{32'h42a1199a};
test_output[3504:3504] = '{32'h45b80d0f};
test_input[28040:28047] = '{32'h428643ca, 32'hc2935d43, 32'hc2929877, 32'h429d4214, 32'h410b6982, 32'h42a49bc8, 32'hc1db5b81, 32'hc18f0679};
test_weights[28040:28047] = '{32'h42a85bc8, 32'hc216bfbb, 32'h428ceb10, 32'hc253401c, 32'h426df363, 32'h42bd0b7e, 32'hc28613c6, 32'h42be1955};
test_bias[3505:3505] = '{32'hc2aba26e};
test_output[3505:3505] = '{32'h45e92f4e};
test_input[28048:28055] = '{32'h42966bde, 32'h41eff281, 32'hc286d2ca, 32'h4141c094, 32'h4234c9cb, 32'h42208a0c, 32'hc1cf2db7, 32'h42a6e8d4};
test_weights[28048:28055] = '{32'hc185ce3e, 32'hc20903c2, 32'hc295b9d1, 32'hc238c6f1, 32'h41890dee, 32'h421fd766, 32'h4215a8c6, 32'h4295e851};
test_bias[3506:3506] = '{32'h3fd522d9};
test_output[3506:3506] = '{32'h461a2ff1};
test_input[28056:28063] = '{32'hc2599277, 32'hc2512cbf, 32'hc190b4e3, 32'hc1f80cc8, 32'hbfa2f2d7, 32'h40ee8ccc, 32'h428a9968, 32'h42b11300};
test_weights[28056:28063] = '{32'h41e11895, 32'h42afc85c, 32'h427526d0, 32'hc2c43fa2, 32'h42771af8, 32'hc28dedd7, 32'h429f81fc, 32'h42856229};
test_bias[3507:3507] = '{32'hc2372cbf};
test_output[3507:3507] = '{32'h45cdcb34};
test_input[28064:28071] = '{32'h4232b001, 32'h415cef94, 32'hc2894a26, 32'h42696656, 32'hc254b291, 32'h421b953b, 32'h41b9ed8d, 32'h41d6d56b};
test_weights[28064:28071] = '{32'hc264c33b, 32'h4264f0cc, 32'h4287dd89, 32'hc28a4557, 32'h42bef73f, 32'h42497ed0, 32'h41d808ec, 32'h422531fd};
test_bias[3508:3508] = '{32'h42726b57};
test_output[3508:3508] = '{32'hc63819a9};
test_input[28072:28079] = '{32'h4283084f, 32'h419b2646, 32'h42b9a954, 32'hc2a5225e, 32'hc24a9ef9, 32'h429ea4d3, 32'hc260b331, 32'hc260a896};
test_weights[28072:28079] = '{32'hc2731cd7, 32'hc252eb4d, 32'hc2bc775f, 32'hc0d3e5bd, 32'h428da59b, 32'h41d60143, 32'h420cbf1a, 32'hc0514367};
test_bias[3509:3509] = '{32'h403bc01b};
test_output[3509:3509] = '{32'hc6809a8a};
test_input[28080:28087] = '{32'hc1cfcf2e, 32'hc1dce178, 32'h423dcd85, 32'hc0df5408, 32'h41b1e6f7, 32'h42343ff3, 32'hc19486f3, 32'h42c14695};
test_weights[28080:28087] = '{32'hc2c71207, 32'hc2684df2, 32'h4213dd82, 32'hc0aa8b31, 32'hc026c4ca, 32'h419505c5, 32'h42080792, 32'hc15702c5};
test_bias[3510:3510] = '{32'hc204e14e};
test_output[3510:3510] = '{32'h4595f44b};
test_input[28088:28095] = '{32'hc2844529, 32'h41a9dec7, 32'hc251d062, 32'h41931625, 32'hc25784b8, 32'h424b67a4, 32'hc1470de9, 32'hc29eef44};
test_weights[28088:28095] = '{32'h406f3de8, 32'hc267e071, 32'h4236a6b4, 32'h42a91b0a, 32'h4191cf78, 32'h424e6ebd, 32'hc24d9709, 32'hc2942c66};
test_bias[3511:3511] = '{32'h425564bb};
test_output[3511:3511] = '{32'h45b87eaa};
test_input[28096:28103] = '{32'h426408fd, 32'h42a42761, 32'h42826cd4, 32'h41847416, 32'h41b08247, 32'h42c6dc99, 32'hc272c2e4, 32'h42b1b551};
test_weights[28096:28103] = '{32'h41201f0f, 32'hc1cd3fa1, 32'h426ae42c, 32'hc2050dfb, 32'hc201094a, 32'h3e64a129, 32'h42bda115, 32'h4196bf34};
test_bias[3512:3512] = '{32'h41ac4547};
test_output[3512:3512] = '{32'hc53bc8ed};
test_input[28104:28111] = '{32'hc1884dee, 32'hc0b2f073, 32'hc1d984be, 32'h42b22d74, 32'hc2c11aca, 32'hc1a37df0, 32'hc1ded4c0, 32'hc1d69c02};
test_weights[28104:28111] = '{32'hc283da74, 32'hc27f352c, 32'h42899b94, 32'hc25d82f4, 32'hc0afe37d, 32'h4196c039, 32'hc2b3a3c0, 32'h42215443};
test_bias[3513:3513] = '{32'hc28e519e};
test_output[3513:3513] = '{32'hc56f5f84};
test_input[28112:28119] = '{32'hc09dd94a, 32'hc228108a, 32'h42510606, 32'h3f293c23, 32'h42a525b5, 32'hc262ecc6, 32'h41bffaeb, 32'h4286b462};
test_weights[28112:28119] = '{32'hc279cb10, 32'hc2b75eca, 32'h42976d42, 32'h42c4629a, 32'hc29d5936, 32'hc27a4408, 32'h421671cb, 32'hc1db0631};
test_bias[3514:3514] = '{32'hc2b4d19c};
test_output[3514:3514] = '{32'h45835768};
test_input[28120:28127] = '{32'hc2beb658, 32'hc2a0e992, 32'h41ac629c, 32'hc21cf4fe, 32'hc244a420, 32'hc1f0ac7a, 32'hc213b895, 32'hc28d9aee};
test_weights[28120:28127] = '{32'hc2a41ec9, 32'hc28cec30, 32'h42931275, 32'hc2845bfb, 32'h4133e12d, 32'hc2c3b235, 32'h40513269, 32'h42ab0cad};
test_bias[3515:3515] = '{32'hc1e829fa};
test_output[3515:3515] = '{32'h4658951f};
test_input[28128:28135] = '{32'h429e3d86, 32'h3f858d41, 32'hc2c23112, 32'hc2aad0a0, 32'h424dc8ac, 32'hc27856ae, 32'hc100c940, 32'hc225a61c};
test_weights[28128:28135] = '{32'h4284b2ad, 32'hc204d350, 32'h40603181, 32'hc10fde8a, 32'hc20d250e, 32'hc23dbcae, 32'h42c056e9, 32'hc2a473e5};
test_bias[3516:3516] = '{32'h42389007};
test_output[3516:3516] = '{32'h4613a64e};
test_input[28136:28143] = '{32'h42298bed, 32'hc1f85834, 32'hc2ad842b, 32'hc2044b5d, 32'hc1d702dd, 32'h41849a42, 32'h408c89a8, 32'hc263a369};
test_weights[28136:28143] = '{32'hc29d3650, 32'h42b4b2dd, 32'hc289cc33, 32'h4289e560, 32'hc2ac837f, 32'h40a932a9, 32'hc247ebd5, 32'hc26ceb68};
test_bias[3517:3517] = '{32'h42290422};
test_output[3517:3517] = '{32'h4545804e};
test_input[28144:28151] = '{32'hc2603b1f, 32'h42a69f8c, 32'hc29b4fda, 32'hc27359f5, 32'hc2c5531f, 32'hc262d260, 32'h4228d843, 32'h42b0fd07};
test_weights[28144:28151] = '{32'h41d1a744, 32'hc209f21d, 32'hc21bf3fb, 32'h415f444d, 32'hc292c09d, 32'h429ba707, 32'hc2b1271c, 32'hc29d3482};
test_bias[3518:3518] = '{32'h428457ba};
test_output[3518:3518] = '{32'hc61bb72e};
test_input[28152:28159] = '{32'hc29408b7, 32'hc1741033, 32'hc294c8de, 32'hc2ba9968, 32'hc2b8da41, 32'hc056882a, 32'hc198fb3e, 32'hc28ac478};
test_weights[28152:28159] = '{32'hc285eb2f, 32'hc26a6e11, 32'h429385e5, 32'hc1c6bee3, 32'h4080befe, 32'hc277c977, 32'h42bc436d, 32'h428ca669};
test_bias[3519:3519] = '{32'hc1260773};
test_output[3519:3519] = '{32'hc5826acf};
test_input[28160:28167] = '{32'hc10d8fae, 32'h42aeb122, 32'hc2b201b0, 32'hc26f9efd, 32'h41a686ec, 32'h4298f45e, 32'h41562fe1, 32'hc28d7208};
test_weights[28160:28167] = '{32'h42af9809, 32'h425444fe, 32'h40f04060, 32'hc0c226a6, 32'hc220101d, 32'h401eb169, 32'h3f003f68, 32'h42b5f6c0};
test_bias[3520:3520] = '{32'h427b675c};
test_output[3520:3520] = '{32'hc557e994};
test_input[28168:28175] = '{32'hc2c13f59, 32'h420d05d3, 32'hc0d09fc0, 32'hc26b2b7f, 32'h422e4de0, 32'h41fa4255, 32'h4172f0a9, 32'hc22b2105};
test_weights[28168:28175] = '{32'h42b867c8, 32'h42aabaf2, 32'hc05be7b0, 32'h41a38f94, 32'h4284b174, 32'hc16d778b, 32'h4229864f, 32'h4282c5c1};
test_bias[3521:3521] = '{32'hc2c477c2};
test_output[3521:3521] = '{32'hc5d7c1ea};
test_input[28176:28183] = '{32'h423b1ea4, 32'h40b29911, 32'h41c33b89, 32'h4182f552, 32'h42a03967, 32'hc2a2a02c, 32'h40ccff4b, 32'hc2b70791};
test_weights[28176:28183] = '{32'hc223a6aa, 32'h41367e7c, 32'hc2b306a5, 32'hbfbd20c3, 32'hc1832211, 32'hc2275062, 32'hc2ab22f3, 32'hc1098bf7};
test_bias[3522:3522] = '{32'h4241d2d3};
test_output[3522:3522] = '{32'hc4d27bb7};
test_input[28184:28191] = '{32'hc189bfda, 32'hc0c7a82f, 32'h42c58f48, 32'hc2962ae1, 32'hc1bbea70, 32'h427c29e6, 32'hc26b3a55, 32'hc227bfcc};
test_weights[28184:28191] = '{32'hc2aa21e9, 32'hc2182dbd, 32'h42296f36, 32'hc03dc48e, 32'hc0a4c3e0, 32'h428b04f3, 32'h4268e8a4, 32'h41e00498};
test_bias[3523:3523] = '{32'h422ecc8b};
test_output[3523:3523] = '{32'h45bd4807};
test_input[28192:28199] = '{32'h4232b2eb, 32'h41f54f14, 32'hc2a571e0, 32'hc1c4d8b7, 32'hc229e875, 32'h42071cff, 32'hc2401c70, 32'h42a15e47};
test_weights[28192:28199] = '{32'hc2943c7b, 32'hc28469da, 32'h41c33b92, 32'h424b7a94, 32'h42161c38, 32'hc282d409, 32'h4224984b, 32'h4287115f};
test_bias[3524:3524] = '{32'hc2940031};
test_output[3524:3524] = '{32'hc60ce337};
test_input[28200:28207] = '{32'h4221d2c4, 32'hc2a60f06, 32'h42429c7d, 32'h42435cd1, 32'hc2660bc4, 32'h42be0bc2, 32'h423f1808, 32'h4072ad69};
test_weights[28200:28207] = '{32'hc26127bd, 32'h40be46e1, 32'hc0a6f4db, 32'h4031f03e, 32'hc2c39a91, 32'hc20988a5, 32'hc1085135, 32'hc2b69124};
test_bias[3525:3525] = '{32'hc23ebb39};
test_output[3525:3525] = '{32'hc4a68921};
test_input[28208:28215] = '{32'h40205f57, 32'h41eac1c8, 32'h4119a177, 32'hc2c74576, 32'h42923aa6, 32'hc205512c, 32'hc2991085, 32'hc2b42fae};
test_weights[28208:28215] = '{32'hc28cd965, 32'h42b15aeb, 32'hc29b09e7, 32'h42aa39fc, 32'hc192e7d3, 32'hc2555c3f, 32'hc207fe53, 32'h42690ca5};
test_bias[3526:3526] = '{32'hc25c1d35};
test_output[3526:3526] = '{32'hc60da758};
test_input[28216:28223] = '{32'hc19d176c, 32'h42c1bf01, 32'h3f83f28f, 32'hc2a9618f, 32'hc21a2ed4, 32'h42455c1f, 32'h42457e59, 32'h42a0e85e};
test_weights[28216:28223] = '{32'h42419c9a, 32'hc173767d, 32'h424f56f1, 32'hc2adc954, 32'hc211fec5, 32'hc16d0d3c, 32'h4283c30a, 32'h425eda2f};
test_bias[3527:3527] = '{32'hc2bf3f1b};
test_output[3527:3527] = '{32'h464fdd21};
test_input[28224:28231] = '{32'hc23c711f, 32'h4133d80f, 32'h42c7548b, 32'hc27ab016, 32'hc2b5d06d, 32'hc12300bb, 32'h42b9c0f0, 32'hc239c7e9};
test_weights[28224:28231] = '{32'h3f8e5b30, 32'hc2a4b295, 32'h3e2a6830, 32'hc2c5487b, 32'h4121d2be, 32'hc2934ea6, 32'h42a70af8, 32'hc2b81e19};
test_bias[3528:3528] = '{32'hc2c4a504};
test_output[3528:3528] = '{32'h4684b445};
test_input[28232:28239] = '{32'h423228f2, 32'hc17bc453, 32'hc07ad883, 32'h42b7339d, 32'h42bfc6f5, 32'hc1fd8c26, 32'h42180c39, 32'h42aa915f};
test_weights[28232:28239] = '{32'h41bfd14a, 32'hc281ec74, 32'hc200497b, 32'hc25c9f37, 32'h4184388a, 32'h42891da8, 32'h42ae8580, 32'hc2ae037d};
test_bias[3529:3529] = '{32'hc1c9ee6b};
test_output[3529:3529] = '{32'hc5ec084e};
test_input[28240:28247] = '{32'hc1cf7cee, 32'h426ba14c, 32'h42c5f212, 32'h42841e23, 32'h400e7110, 32'hc28b2fd4, 32'h423c0847, 32'hc2ab60fb};
test_weights[28240:28247] = '{32'hc28c01bf, 32'hc25e52e1, 32'hc23bde1f, 32'hc190d0eb, 32'h428baaff, 32'h42936d17, 32'hc16db2a0, 32'h425d5b26};
test_bias[3530:3530] = '{32'h42b14e70};
test_output[3530:3530] = '{32'hc689b9ec};
test_input[28248:28255] = '{32'hc17e9dbc, 32'h42ab4e9f, 32'hc21dc386, 32'h42045a77, 32'hc114fd52, 32'h424a456f, 32'h426a4075, 32'hc20f8cb2};
test_weights[28248:28255] = '{32'hc1f5fe33, 32'h4288aac0, 32'h40be655c, 32'hc0841258, 32'hc2bc5fe1, 32'h42363f09, 32'h41b75679, 32'h41c4b070};
test_bias[3531:3531] = '{32'hc28d0b94};
test_output[3531:3531] = '{32'h46151567};
test_input[28256:28263] = '{32'hc06d89de, 32'hc2a832d3, 32'hc29970f1, 32'hc18a741f, 32'h4272609c, 32'h425580b9, 32'h4224a092, 32'hc2ab4daa};
test_weights[28256:28263] = '{32'hc1340ca3, 32'h4296ef18, 32'hc29a2feb, 32'h42b3e780, 32'hc265f39c, 32'hc0ee9349, 32'h427c9814, 32'hc1958dd4};
test_bias[3532:3532] = '{32'h42132079};
test_output[3532:3532] = '{32'hc4c6ef40};
test_input[28264:28271] = '{32'hc1cf5e4d, 32'hc23e7ae5, 32'h4139317a, 32'hc27174e9, 32'h42531e10, 32'hc0e9de76, 32'h4223ec24, 32'h418dd341};
test_weights[28264:28271] = '{32'h428fef56, 32'hc1f087b0, 32'hc2c7832f, 32'h428612c4, 32'hc27117dc, 32'hc23377b4, 32'h420c7e5e, 32'hc229a56e};
test_bias[3533:3533] = '{32'h4248dccf};
test_output[3533:3533] = '{32'hc5f2343c};
test_input[28272:28279] = '{32'hc294b936, 32'h42176adb, 32'h40ec1cd3, 32'h41ce3243, 32'h42012973, 32'h41cdfe93, 32'hc219ee3d, 32'h429ba561};
test_weights[28272:28279] = '{32'h424b8aac, 32'h426494e7, 32'hc1c9dae0, 32'h41e54926, 32'h41de8177, 32'hc230340d, 32'h42348127, 32'hc291dc79};
test_bias[3534:3534] = '{32'h4221192f};
test_output[3534:3534] = '{32'hc6079159};
test_input[28280:28287] = '{32'hc2b6dd25, 32'h427e05c0, 32'hc1226e9a, 32'hc20eb379, 32'h42b089b6, 32'hc284569d, 32'h42be46f8, 32'h42a6b34d};
test_weights[28280:28287] = '{32'hc2699d9f, 32'hc2b02ccb, 32'h42bc6f99, 32'h4290f087, 32'hc240ea1e, 32'h41f2fc0a, 32'hc2a60f62, 32'hc26f7dfb};
test_bias[3535:3535] = '{32'hc28af364};
test_output[3535:3535] = '{32'hc6b3dc21};
test_input[28288:28295] = '{32'hc165ccfa, 32'hc292c231, 32'hc17413e7, 32'hc00ff4a3, 32'h41697cbf, 32'hc186d7ce, 32'h40d4d473, 32'hc198ce1e};
test_weights[28288:28295] = '{32'h42a77e2a, 32'hc15bb851, 32'hc02fa0c2, 32'h42167750, 32'h4299d975, 32'h42bd65bf, 32'h4291a35f, 32'h4297984b};
test_bias[3536:3536] = '{32'h42b69306};
test_output[3536:3536] = '{32'hc4c5f5c9};
test_input[28296:28303] = '{32'h41c1a96e, 32'h42b6de2c, 32'h42822f6e, 32'hc2af10af, 32'h425f88ac, 32'hc2bce76b, 32'h425d63f9, 32'hc227873f};
test_weights[28296:28303] = '{32'hc26f1269, 32'hc0f6da75, 32'h416eff64, 32'h41ca64ed, 32'h4295d781, 32'hc280fe38, 32'h42ade9d7, 32'h42568fac};
test_bias[3537:3537] = '{32'hc1f5aa8e};
test_output[3537:3537] = '{32'h46132f6a};
test_input[28304:28311] = '{32'hc2887152, 32'hc25e6bc6, 32'hc22abdfd, 32'h4297eec4, 32'h41c7995b, 32'hc270e7ff, 32'hc1c45069, 32'hc21e1ab8};
test_weights[28304:28311] = '{32'h41cebd4a, 32'h42a5805c, 32'h3fd405be, 32'h41340c01, 32'hc1dfa6fc, 32'h41a28508, 32'hc2bc29b4, 32'h428aa22e};
test_bias[3538:3538] = '{32'hc2ad0121};
test_output[3538:3538] = '{32'hc5fa9714};
test_input[28312:28319] = '{32'hc2a4883a, 32'hc29ec470, 32'hc0e26319, 32'h42480f45, 32'h4229ef4c, 32'hc21e6e83, 32'h401fd4bf, 32'h41b22c93};
test_weights[28312:28319] = '{32'hc2abb396, 32'hc2997fbc, 32'hc25eda85, 32'h42c559b0, 32'hc28ca883, 32'hc2b53559, 32'h42bf83f0, 32'h40a365e4};
test_bias[3539:3539] = '{32'hc2a8c849};
test_output[3539:3539] = '{32'h469733d5};
test_input[28320:28327] = '{32'h42aaa581, 32'h42a1b317, 32'hc23e1dd6, 32'h4298d954, 32'hc2090f67, 32'hc277fa9f, 32'h41a29f00, 32'h41ff1188};
test_weights[28320:28327] = '{32'hc25110dc, 32'h42951e8b, 32'hc2a379eb, 32'h4228b00c, 32'h42788a61, 32'hc29a3c1e, 32'h421c8897, 32'hc2b6fa91};
test_bias[3540:3540] = '{32'hc235f956};
test_output[3540:3540] = '{32'h460f252f};
test_input[28328:28335] = '{32'h4051d0ea, 32'h4217b21b, 32'hc1f37fcc, 32'hc18d4781, 32'hc264d3ad, 32'hc298ba11, 32'hc2a42361, 32'hc20a0bb1};
test_weights[28328:28335] = '{32'hc27c5e94, 32'h41282d1d, 32'h428d511a, 32'h41f9f4de, 32'h4203a5e1, 32'h42066fd3, 32'hc258464e, 32'hc2a9ef22};
test_bias[3541:3541] = '{32'h427eb64c};
test_output[3541:3541] = '{32'h43ecb5eb};
test_input[28336:28343] = '{32'hc0f1e518, 32'h42755bf6, 32'h42266884, 32'h4289e513, 32'h42ab1a78, 32'hc2c00364, 32'hc2858580, 32'hc28871e5};
test_weights[28336:28343] = '{32'h42a14c92, 32'h4203213a, 32'hc2180318, 32'h42abe7ed, 32'h42b7b36c, 32'h427a8a3b, 32'h42b26a42, 32'h423e4778};
test_bias[3542:3542] = '{32'hc2be9c3a};
test_output[3542:3542] = '{32'hc4d524ef};
test_input[28344:28351] = '{32'hc2200d1e, 32'hc28811a0, 32'h4202f07d, 32'hc0c30482, 32'hc2c4f285, 32'hc279dae4, 32'h425587a5, 32'h40b6b9df};
test_weights[28344:28351] = '{32'hc279f446, 32'h40d0d360, 32'h421ede3d, 32'h4216bf6e, 32'h4167d130, 32'h428866d2, 32'h42a91238, 32'h42428ac3};
test_bias[3543:3543] = '{32'h42479596};
test_output[3543:3543] = '{32'h450e8540};
test_input[28352:28359] = '{32'h42253d5e, 32'hc12d222e, 32'h4295dfce, 32'h421fa689, 32'h42b72f59, 32'h4117e893, 32'hc1e3d681, 32'h42891e2a};
test_weights[28352:28359] = '{32'hc1a34332, 32'h41ded880, 32'h41d788a2, 32'h425c775b, 32'hc2b644aa, 32'hc2aa3aa6, 32'h40e183be, 32'h425746b2};
test_bias[3544:3544] = '{32'h42216433};
test_output[3544:3544] = '{32'hc51f791d};
test_input[28360:28367] = '{32'h422d13f3, 32'hc28a46ce, 32'h4299e154, 32'hc258f5ea, 32'h41eaa2ce, 32'h4204ad52, 32'hc2ab62b8, 32'hc2ab82f6};
test_weights[28360:28367] = '{32'h429af2ae, 32'h4291642f, 32'h42bc80f0, 32'h40c88f48, 32'h41f8b72c, 32'hc223ced2, 32'h4193503b, 32'hc2158bcd};
test_bias[3545:3545] = '{32'hc27129d3};
test_output[3545:3545] = '{32'h45c6bacb};
test_input[28368:28375] = '{32'h427b0243, 32'h429eedf5, 32'h42274f8d, 32'h425b9dd9, 32'hc1e37452, 32'h428fd44a, 32'h429673bc, 32'hc2afc31b};
test_weights[28368:28375] = '{32'h42609581, 32'h415d1312, 32'h420ce477, 32'h41d56c8f, 32'hc210307a, 32'hc1934292, 32'h428ddc12, 32'h42098839};
test_bias[3546:3546] = '{32'hc2c70ba6};
test_output[3546:3546] = '{32'h46140c32};
test_input[28376:28383] = '{32'hc2214851, 32'hc2952491, 32'hc297e5d2, 32'hc2074297, 32'h406b7099, 32'h40ce7e9b, 32'hc2b4e002, 32'h4208d644};
test_weights[28376:28383] = '{32'h42534fd2, 32'h41033b9e, 32'h429c1f89, 32'hc271a000, 32'hc2b0d9e5, 32'hc2945a31, 32'hc2949039, 32'h42673ea7};
test_bias[3547:3547] = '{32'h4151de47};
test_output[3547:3547] = '{32'h449f9e58};
test_input[28384:28391] = '{32'h40223880, 32'hc2a3838b, 32'h410377b0, 32'hc2473105, 32'h420d81f1, 32'hc29c2ad3, 32'hc288f01f, 32'hc2b745e3};
test_weights[28384:28391] = '{32'h4084d727, 32'h3e562780, 32'hc2bf7fa8, 32'h429f510b, 32'h41d01dd9, 32'hc26cade0, 32'hc2897af2, 32'hc2b8aa80};
test_bias[3548:3548] = '{32'hc218b022};
test_output[3548:3548] = '{32'h4659575f};
test_input[28392:28399] = '{32'h42151c41, 32'hc2a28d90, 32'hc29c4bee, 32'h42783a79, 32'h4290276d, 32'hc2c2696a, 32'hc2bf3294, 32'hc2c6da82};
test_weights[28392:28399] = '{32'hc220d37b, 32'hc1539157, 32'hc223014c, 32'h40129960, 32'hc263538d, 32'h4277e7e0, 32'h4274b92f, 32'h424fb519};
test_bias[3549:3549] = '{32'h42be4caf};
test_output[3549:3549] = '{32'hc68dad35};
test_input[28400:28407] = '{32'hc2bd904a, 32'hc279bb46, 32'h4287b80b, 32'hc296c226, 32'hc2892085, 32'hc2b298c1, 32'h40baa55d, 32'hc151d267};
test_weights[28400:28407] = '{32'hc250d3d2, 32'hc23417a6, 32'hc038aa94, 32'hc27a1288, 32'h424f3b1b, 32'h41bd3014, 32'hc2b6bcc4, 32'h428e3756};
test_bias[3550:3550] = '{32'h42acf4c8};
test_output[3550:3550] = '{32'h45a388d9};
test_input[28408:28415] = '{32'hc2433139, 32'h4066a22a, 32'h41a91961, 32'hc1f2b885, 32'hc0e26a07, 32'hc2c0de00, 32'h422f2cc2, 32'hc29818f2};
test_weights[28408:28415] = '{32'hc2c425ea, 32'hc24cf4ee, 32'h422326e8, 32'hc1b46493, 32'hc088b4cd, 32'hc22f7960, 32'hc2774844, 32'hc184c33e};
test_bias[3551:3551] = '{32'h422ce5e4};
test_output[3551:3551] = '{32'h460cb818};
test_input[28416:28423] = '{32'h3ee2100d, 32'h42bfd2a9, 32'hc1886508, 32'h41647b28, 32'hc245e99e, 32'hc2abbc3b, 32'h42467bbf, 32'hc2297211};
test_weights[28416:28423] = '{32'hc285820f, 32'h4299833c, 32'h42a0063b, 32'hc2a9e539, 32'h42a1795d, 32'hc20dd6a2, 32'h4259d594, 32'h4225199e};
test_bias[3552:3552] = '{32'h42c7b7af};
test_output[3552:3552] = '{32'h4597d744};
test_input[28424:28431] = '{32'h402f9dee, 32'h422f7d91, 32'h41a280cd, 32'h426f486c, 32'hc29da184, 32'h422a064c, 32'hc1308593, 32'h424d5d4b};
test_weights[28424:28431] = '{32'hc14089ba, 32'h4227729a, 32'hc27247f5, 32'h422724d2, 32'hc09e4dc5, 32'hc2041adc, 32'hc2505561, 32'h42b6eb2e};
test_bias[3553:3553] = '{32'hc20d5b7e};
test_output[3553:3553] = '{32'h45e3eee5};
test_input[28432:28439] = '{32'h4254686b, 32'h414a501c, 32'hc2937f86, 32'hc1ee5026, 32'h42963748, 32'h424c7b78, 32'h42c655e6, 32'hc1e38760};
test_weights[28432:28439] = '{32'h4221a755, 32'h40ec5808, 32'h42c18e30, 32'h4280672b, 32'h42a2d921, 32'h42311cd1, 32'hc2283d5e, 32'hc2217637};
test_bias[3554:3554] = '{32'hc1a83930};
test_output[3554:3554] = '{32'hc4b866ba};
test_input[28440:28447] = '{32'hc1c313a1, 32'h42903dad, 32'h42a1993e, 32'h42c0c8ac, 32'hc290598f, 32'hc277e87c, 32'hc216184d, 32'hc1f1c767};
test_weights[28440:28447] = '{32'hc2b6836f, 32'h41702031, 32'hc2c13baf, 32'hc23845ec, 32'hc227b4ee, 32'hc2c3a05a, 32'h4109a6c2, 32'h418801cc};
test_bias[3555:3555] = '{32'h42618ea5};
test_output[3555:3555] = '{32'hc41de303};
test_input[28448:28455] = '{32'h421ddba3, 32'hc21c5a9d, 32'hc24c3598, 32'h4220ef97, 32'hc298e791, 32'h4225829e, 32'h40bd1bf5, 32'hc1cdd633};
test_weights[28448:28455] = '{32'hc217f69e, 32'hc27f8a6c, 32'hc1b10990, 32'h4264aec0, 32'h42c49f11, 32'hc2967a4e, 32'h41d15603, 32'h42b5531a};
test_bias[3556:3556] = '{32'hc25435b5};
test_output[3556:3556] = '{32'hc603c223};
test_input[28456:28463] = '{32'hc261ea04, 32'h42c32ec3, 32'h41656853, 32'hc273b9f5, 32'hc1f9d9f7, 32'h42977779, 32'hc2a58edf, 32'h4102af62};
test_weights[28456:28463] = '{32'hc132db6f, 32'h41a248ef, 32'h42b3c9ae, 32'hc163a0ca, 32'h3eab8228, 32'hc2c707a9, 32'hc29097b2, 32'h427bf019};
test_bias[3557:3557] = '{32'hc1250f8d};
test_output[3557:3557] = '{32'h4567c7d2};
test_input[28464:28471] = '{32'hc28dcb61, 32'hc2a856ee, 32'h427be8c1, 32'h42b32444, 32'h429d060c, 32'h41ca89ef, 32'h41bc1028, 32'hc201d7ed};
test_weights[28464:28471] = '{32'hc293c2ec, 32'h413080ec, 32'h40869a5c, 32'hbf24bdd9, 32'h42bd5947, 32'hbfe9a30e, 32'h40bc072a, 32'hc2c33fe8};
test_bias[3558:3558] = '{32'h42ae8016};
test_output[3558:3558] = '{32'h466f0793};
test_input[28472:28479] = '{32'hc2245ed5, 32'hc2069c08, 32'hc1e2b635, 32'hc280d6cc, 32'hbf6626f4, 32'hc289342d, 32'h420e6639, 32'h4268e8bc};
test_weights[28472:28479] = '{32'hc25af1e2, 32'h42a1189d, 32'hc0cb7848, 32'h428cf3a0, 32'h423611c5, 32'hc2a0a1f0, 32'hc29f8e42, 32'hc295cf7d};
test_bias[3559:3559] = '{32'h40d6c9b5};
test_output[3559:3559] = '{32'hc5cc9963};
test_input[28480:28487] = '{32'hc2baa2b1, 32'hc2a6cf40, 32'h428db30e, 32'h42644f61, 32'hc2acf538, 32'hc10763c0, 32'h42185b0f, 32'h40f9c6e9};
test_weights[28480:28487] = '{32'hc2804020, 32'hc2420228, 32'hc2b0a5ee, 32'hbf3af209, 32'hc105852d, 32'h42b638d4, 32'hc2138d26, 32'hc2a55669};
test_bias[3560:3560] = '{32'h42c3e983};
test_output[3560:3560] = '{32'h44d808e9};
test_input[28488:28495] = '{32'hc20a2c52, 32'h42b71b46, 32'h410b2503, 32'hc2b117b0, 32'hc2b67cb3, 32'hc22ad646, 32'hc2b3b84d, 32'hc2b31bbb};
test_weights[28488:28495] = '{32'h42a0f837, 32'hc27395b7, 32'hc2235ea3, 32'hc252fd89, 32'hc198e553, 32'hc2b9ed09, 32'hc2986a89, 32'h42c550e0};
test_bias[3561:3561] = '{32'hc12ee02e};
test_output[3561:3561] = '{32'hc3a1f62a};
test_input[28496:28503] = '{32'h42bb1eb3, 32'h424da26c, 32'hc2abb9b9, 32'hc2a9d29f, 32'hc259e216, 32'h401f68d0, 32'h42b4b43c, 32'hc0f1aa6c};
test_weights[28496:28503] = '{32'h428f8eb2, 32'hc22bcb32, 32'h4240a101, 32'hc23508fc, 32'hc2804b95, 32'h42ade88f, 32'h42a69a7f, 32'h42bafdd0};
test_bias[3562:3562] = '{32'hc274167c};
test_output[3562:3562] = '{32'h46657795};
test_input[28504:28511] = '{32'hc26524a6, 32'hc2a22bbe, 32'hc28ce38e, 32'hc2a393de, 32'hc2a2961e, 32'h42b55774, 32'hc2bee6ee, 32'hc23842cb};
test_weights[28504:28511] = '{32'h419b03a3, 32'h416d2c7f, 32'hc1ca2aa3, 32'hc2909286, 32'h425ed8a6, 32'h41a64799, 32'hc282629f, 32'h407e2468};
test_bias[3563:3563] = '{32'h4295fbd8};
test_output[3563:3563] = '{32'h460a4b38};
test_input[28512:28519] = '{32'hc262940b, 32'h42646363, 32'hc1433467, 32'h41f17fff, 32'hc1ada516, 32'hc2c47640, 32'hc2b1fcac, 32'h42a6c5ea};
test_weights[28512:28519] = '{32'hc184aa5a, 32'h4284bfb2, 32'h426a89f3, 32'h4182422d, 32'h417e4014, 32'hc22315e2, 32'hc27150bf, 32'hc2566b16};
test_bias[3564:3564] = '{32'hc22e4190};
test_output[3564:3564] = '{32'h460cf331};
test_input[28520:28527] = '{32'hc07f56a1, 32'h424a3e08, 32'hc1f47400, 32'hc2bcc033, 32'hc24c35b5, 32'h428fc453, 32'hc2042ad2, 32'hc204454b};
test_weights[28520:28527] = '{32'h42882fa3, 32'h428ec2ab, 32'hc28b9cc9, 32'h42c56077, 32'hc25d99a0, 32'hc29f419d, 32'hc0a0a7fc, 32'hc2ae8b85};
test_bias[3565:3565] = '{32'hc11d46ee};
test_output[3565:3565] = '{32'hc56710a7};
test_input[28528:28535] = '{32'h4298a4be, 32'hc1d8c8eb, 32'hc2925ad7, 32'h427cdc86, 32'hc2afe48c, 32'hbf93fb01, 32'h423382e5, 32'h429939bd};
test_weights[28528:28535] = '{32'h413fd91b, 32'hc1b1fd4b, 32'hc297fb41, 32'hc22cbf21, 32'hc239e225, 32'hc2b67fcf, 32'hc2ade25b, 32'h42b8c0ea};
test_bias[3566:3566] = '{32'h42c78bab};
test_output[3566:3566] = '{32'h4638a1d5};
test_input[28536:28543] = '{32'h41f631bd, 32'hc22c7f90, 32'hbf320514, 32'h423cbc65, 32'h423c4900, 32'h40c453c8, 32'hc29067d0, 32'h42b201ee};
test_weights[28536:28543] = '{32'h42b76e83, 32'hc1b2b032, 32'h40eb6f60, 32'hc2a18526, 32'h42a03c3a, 32'h40446c81, 32'h425df8af, 32'hc2035f9e};
test_bias[3567:3567] = '{32'h4180e6a6};
test_output[3567:3567] = '{32'hc5451b6e};
test_input[28544:28551] = '{32'hc1e3aa33, 32'h4295eb12, 32'hc16571da, 32'h4273c4dd, 32'h4216690b, 32'hc26b85cc, 32'h41e394d6, 32'hc2c774a8};
test_weights[28544:28551] = '{32'hc26ab027, 32'h41702c43, 32'h426415f1, 32'h41ed2f24, 32'hc2a2cb0d, 32'hc20057bd, 32'h420acdf1, 32'h42ad7f6f};
test_bias[3568:3568] = '{32'hc2bb9025};
test_output[3568:3568] = '{32'hc5a0cb19};
test_input[28552:28559] = '{32'hc23bfff8, 32'h3fa3a8bc, 32'h4267c387, 32'hc13954e9, 32'h42aca2db, 32'h40c1c24b, 32'h42424897, 32'hc2a207ea};
test_weights[28552:28559] = '{32'hc144eb82, 32'h429113a0, 32'h42a02954, 32'hc2ad0eee, 32'h412c4edb, 32'hc2161818, 32'h420226b7, 32'hc23f6747};
test_bias[3569:3569] = '{32'hc20acfc0};
test_output[3569:3569] = '{32'h464258a6};
test_input[28560:28567] = '{32'hc26bdcb3, 32'h4299c4b9, 32'hc230e6de, 32'h4273c0cf, 32'h4283a9ea, 32'h42844248, 32'hc2657f2c, 32'h42bfa20b};
test_weights[28560:28567] = '{32'h4236a207, 32'hc20c1590, 32'h4291c162, 32'h41e14d3f, 32'hc294a472, 32'h41ea8a66, 32'h429b1fe6, 32'hc143c3a2};
test_bias[3570:3570] = '{32'hc2095d16};
test_output[3570:3570] = '{32'hc6723991};
test_input[28568:28575] = '{32'h42938877, 32'h428485ed, 32'hc223e151, 32'hc1f42e02, 32'h422ff308, 32'h41ca06e1, 32'hbf2405d1, 32'h4203d6f1};
test_weights[28568:28575] = '{32'h42798a45, 32'hc18c9cee, 32'h4264dda0, 32'h4297d022, 32'hc1b5afd6, 32'h428afa2f, 32'hc28fad52, 32'h42991226};
test_bias[3571:3571] = '{32'hc291cb4c};
test_output[3571:3571] = '{32'h44fd7a54};
test_input[28576:28583] = '{32'h4152f441, 32'h4293649f, 32'hc2831325, 32'h41f0c995, 32'h420deee1, 32'hc1f379dd, 32'h41525092, 32'h4289913d};
test_weights[28576:28583] = '{32'h41cbf103, 32'hc0f067d7, 32'hc29025ac, 32'hc2804dc7, 32'hc11fa577, 32'hc26737da, 32'hc2224fc6, 32'h418e942c};
test_bias[3572:3572] = '{32'h4276d277};
test_output[3572:3572] = '{32'h4593f413};
test_input[28584:28591] = '{32'hbfa686f3, 32'hc2018fa9, 32'h40731eb0, 32'h40cdaa54, 32'h429aba94, 32'h4238284a, 32'h4280863f, 32'h414ce1fb};
test_weights[28584:28591] = '{32'h4030aa1f, 32'hc1c84d67, 32'h4219e3a7, 32'hc282167f, 32'h41f8f8be, 32'hc2a75279, 32'hc095859e, 32'h42960f4b};
test_bias[3573:3573] = '{32'hc0ed64a2};
test_output[3573:3573] = '{32'hc37f6dba};
test_input[28592:28599] = '{32'h41318a28, 32'h41310564, 32'h42c72235, 32'h4022412f, 32'h42af0db0, 32'hc281c8ce, 32'h4262c4fc, 32'hc175a18c};
test_weights[28592:28599] = '{32'h429ffde9, 32'h4293be7f, 32'hc286978f, 32'h4278263f, 32'hc1a5f2de, 32'hc23ce73a, 32'h42aa2e64, 32'hc1dba8e5};
test_bias[3574:3574] = '{32'hc230fbdc};
test_output[3574:3574] = '{32'h44c980cd};
test_input[28600:28607] = '{32'hc2a32d07, 32'hc017b608, 32'hc1e75ab1, 32'h41309861, 32'h42b658e6, 32'h41be6bb4, 32'hc28446b4, 32'h4298c486};
test_weights[28600:28607] = '{32'hc24bdeb0, 32'h4202379e, 32'hc202e7bf, 32'h4202e23c, 32'hc2187f95, 32'h41e5ddd2, 32'h4263889c, 32'h41582dad};
test_bias[3575:3575] = '{32'h42c16d85};
test_output[3575:3575] = '{32'hc212d903};
test_input[28608:28615] = '{32'hc2ac4bb6, 32'h4254cfa9, 32'h42b318a8, 32'hc295190d, 32'h42467cdc, 32'h42957625, 32'h41891f52, 32'h42a567a9};
test_weights[28608:28615] = '{32'hbe08280f, 32'h428eb68d, 32'hc28aebc9, 32'hc259f610, 32'hc10d7b5d, 32'h428b8d82, 32'h42472630, 32'hc2098eda};
test_bias[3576:3576] = '{32'h42a6bfa0};
test_output[3576:3576] = '{32'h458d3209};
test_input[28616:28623] = '{32'h4238edc5, 32'h420ab555, 32'h42650164, 32'hc2b111a7, 32'h41905d25, 32'h423c0ddb, 32'h423ad8eb, 32'h405ac57e};
test_weights[28616:28623] = '{32'h42c0791a, 32'h428b5f46, 32'h40c68beb, 32'h427e56f6, 32'h42c51f56, 32'hc083fddf, 32'h42b961a9, 32'h41bd7cf6};
test_bias[3577:3577] = '{32'h427d8222};
test_output[3577:3577] = '{32'h45ef1218};
test_input[28624:28631] = '{32'h427f49e9, 32'hc1785af1, 32'h4290bfa3, 32'h42b2ca19, 32'h41edfded, 32'hc2c07471, 32'h4284b36b, 32'hc23fb2ec};
test_weights[28624:28631] = '{32'h42b3c29e, 32'hc2116e10, 32'h42c1cd03, 32'hc0d43903, 32'h41f548ea, 32'hc257376f, 32'h429ce102, 32'h41b7e3eb};
test_bias[3578:3578] = '{32'h42ba010a};
test_output[3578:3578] = '{32'h46b3bcbc};
test_input[28632:28639] = '{32'hc16268a4, 32'hc2bb77df, 32'h42b0bcfa, 32'hc2913473, 32'hc16f4e2a, 32'h42b78e0a, 32'h423405c3, 32'hc2173a2f};
test_weights[28632:28639] = '{32'h41b6ad36, 32'hc29913b1, 32'h428dacd4, 32'h42a6cc5c, 32'hc24ce874, 32'h428dc8f1, 32'h41a1f507, 32'hc1c0f10c};
test_bias[3579:3579] = '{32'h42a24bd5};
test_output[3579:3579] = '{32'h467da26c};
test_input[28640:28647] = '{32'h42c01dea, 32'h429e18b7, 32'hc2969412, 32'hc092495c, 32'hc1349b7f, 32'h42b50400, 32'h42bff66a, 32'h41d74d6f};
test_weights[28640:28647] = '{32'h428b223f, 32'hc20a9d5f, 32'hc28d8481, 32'h40b2fece, 32'h42acc222, 32'h40ccb956, 32'h41d83cb7, 32'h42a1a9a1};
test_bias[3580:3580] = '{32'hc1dce02c};
test_output[3580:3580] = '{32'h46545c5e};
test_input[28648:28655] = '{32'h4233c244, 32'h421ff05b, 32'hc2a5e34c, 32'hc2b6912e, 32'h426e404b, 32'hc23ec9df, 32'hc20c196c, 32'h3fcc2839};
test_weights[28648:28655] = '{32'h42c5b9c3, 32'hc21f4c9c, 32'h4191d3e8, 32'hc171b2f4, 32'h410718fd, 32'h42421980, 32'hc2129b95, 32'h4275491f};
test_bias[3581:3581] = '{32'hc23801ee};
test_output[3581:3581] = '{32'h450c1720};
test_input[28656:28663] = '{32'hc23ea7d1, 32'h4115ab9c, 32'hc1732c7d, 32'h4195a54f, 32'h4286d06b, 32'hc2941879, 32'h41d34406, 32'hc1ce83d6};
test_weights[28656:28663] = '{32'h40a47e25, 32'hc22cd003, 32'h4284cca2, 32'h42589815, 32'h4267a2f2, 32'hc2be2b8c, 32'h41afca54, 32'h4287293c};
test_bias[3582:3582] = '{32'hc105ee58};
test_output[3582:3582] = '{32'h460e990d};
test_input[28664:28671] = '{32'h429b854e, 32'h42c3980c, 32'h42b64892, 32'hc28c765c, 32'h41b56b32, 32'hc125523e, 32'h428b6e52, 32'hc1c8a0be};
test_weights[28664:28671] = '{32'hc0f2add8, 32'hc25bfda0, 32'h426a45b8, 32'hc1c414bb, 32'hc214f6a1, 32'hc214e1f5, 32'h42afd5d7, 32'hc16dc3a3};
test_bias[3583:3583] = '{32'h4286b51c};
test_output[3583:3583] = '{32'h45e102e5};
test_input[28672:28679] = '{32'h422eabd6, 32'hc2587142, 32'h428fecc5, 32'h42639735, 32'h420771cf, 32'hc28eca66, 32'hc2c58637, 32'hc1d56d48};
test_weights[28672:28679] = '{32'hc2b4aece, 32'h40ab9968, 32'hc1e9669b, 32'h429b9456, 32'hc27710bf, 32'h415acd7e, 32'hc13cfba6, 32'h42a5231c};
test_bias[3584:3584] = '{32'hc2988c62};
test_output[3584:3584] = '{32'hc5be4809};
test_input[28680:28687] = '{32'h421bd161, 32'hc28e5f4a, 32'h42b39088, 32'h4242d602, 32'hc155ee69, 32'hc2595627, 32'hc231d50e, 32'hc259ca82};
test_weights[28680:28687] = '{32'h42c0d8e3, 32'h429999b4, 32'hc2a54c7f, 32'hc1619128, 32'h416b8b4a, 32'hc1992003, 32'hc1f17636, 32'h418e3992};
test_bias[3585:3585] = '{32'hc1f5b9ee};
test_output[3585:3585] = '{32'hc606df36};
test_input[28688:28695] = '{32'hc28e425f, 32'h420b90a0, 32'hc24219b4, 32'h42097510, 32'h4253fec1, 32'hc2ad2692, 32'hc19bbd24, 32'h41d32683};
test_weights[28688:28695] = '{32'h4292215f, 32'h429ddab5, 32'hc1e9691a, 32'hc214f41c, 32'hc2a69cee, 32'hc2970eed, 32'hc2778605, 32'hc29aa75f};
test_bias[3586:3586] = '{32'hc0b0cbbd};
test_output[3586:3586] = '{32'hc48023e6};
test_input[28696:28703] = '{32'h413058be, 32'h423ed202, 32'h428014de, 32'h4260d424, 32'hc22e06a3, 32'hc1f9a64a, 32'hc2b0d2df, 32'hc25794b4};
test_weights[28696:28703] = '{32'hc2ba5984, 32'h421696e6, 32'h41f11880, 32'h421d7255, 32'hc1e05028, 32'h426cf50b, 32'hc142f8ca, 32'hc1f2676b};
test_bias[3587:3587] = '{32'hc1a161ca};
test_output[3587:3587] = '{32'h45d9e764};
test_input[28704:28711] = '{32'hc2c53ed0, 32'hc2bc8b54, 32'h41d3ca74, 32'h4220a846, 32'hc13585d1, 32'h4104792b, 32'hc19caa11, 32'hc1ef1cb9};
test_weights[28704:28711] = '{32'h4146fba1, 32'h42222aa4, 32'hc1f59733, 32'hc2c4db67, 32'h416550c0, 32'hc0e8bcb1, 32'hc21daaa7, 32'h429d3591};
test_bias[3588:3588] = '{32'hc2897932};
test_output[3588:3588] = '{32'hc6368e44};
test_input[28712:28719] = '{32'h4246649e, 32'hc2b4f0af, 32'hc064e186, 32'h425d2cff, 32'hc280a1bd, 32'h42ab1aa6, 32'hc18c1ba6, 32'hc2a7cca6};
test_weights[28712:28719] = '{32'h417e6581, 32'hc1f97bb4, 32'hc2167c37, 32'hc2155a8c, 32'hc1ec0c57, 32'h4214bc2d, 32'h4188dae0, 32'h429707fd};
test_bias[3589:3589] = '{32'hc28f169b};
test_output[3589:3589] = '{32'h424f7f3b};
test_input[28720:28727] = '{32'h41fcf915, 32'h42b300c5, 32'h42903320, 32'h41fdfe4e, 32'hc167e8cc, 32'hc01b2e18, 32'hc23a8e48, 32'h42c718d9};
test_weights[28720:28727] = '{32'hc1c645e9, 32'h417a1566, 32'h3ee52c63, 32'hc241d9b8, 32'hc2441807, 32'hc28f4145, 32'h423cd568, 32'hc29259d7};
test_bias[3590:3590] = '{32'h426eafed};
test_output[3590:3590] = '{32'hc613660e};
test_input[28728:28735] = '{32'hc1905ffd, 32'hc273ce3c, 32'hc22855a8, 32'hc2198ed1, 32'h429101c6, 32'hc2526f49, 32'h41e9f2dd, 32'hc2b09a4e};
test_weights[28728:28735] = '{32'h42adb5bd, 32'h42af9cc6, 32'h3f67aef6, 32'h41b9138b, 32'h42146d7a, 32'h42a23d22, 32'h429f4b08, 32'h425c53a6};
test_bias[3591:3591] = '{32'h42b09991};
test_output[3591:3591] = '{32'hc639747e};
test_input[28736:28743] = '{32'hc2870aab, 32'h42abee72, 32'hc239ffeb, 32'hc261a018, 32'h429dcca9, 32'hc163216d, 32'hc28a887e, 32'h42919068};
test_weights[28736:28743] = '{32'hbfd27bfd, 32'hc20f7b37, 32'hc1e29814, 32'hc1e53dd5, 32'h41d4a86f, 32'h4219d58d, 32'h42836f04, 32'h42c527ef};
test_bias[3592:3592] = '{32'h42a25927};
test_output[3592:3592] = '{32'h4583c0e7};
test_input[28744:28751] = '{32'hc28e9a38, 32'h4243e1f2, 32'h4289af61, 32'hc2bf54a4, 32'hc2bc8050, 32'hc1f749e7, 32'hc2c587d6, 32'hc2582607};
test_weights[28744:28751] = '{32'h4284e071, 32'hc28aa03a, 32'hbfc7acd9, 32'hc25882ea, 32'hc29aa899, 32'h42560851, 32'h429cdfed, 32'h401d0c57};
test_bias[3593:3593] = '{32'hc201bd41};
test_output[3593:3593] = '{32'hc5a6d209};
test_input[28752:28759] = '{32'h42a75531, 32'hc2ac9669, 32'h40d54953, 32'h42473906, 32'h420e8f72, 32'h42c182bd, 32'h41eeb4d6, 32'h42b77b84};
test_weights[28752:28759] = '{32'h42be8ff7, 32'hc28bdfbb, 32'h42a7656f, 32'hc13cfc11, 32'h428a6727, 32'hc272cd99, 32'hc20ed2e9, 32'h41b10810};
test_bias[3594:3594] = '{32'h41faa3d2};
test_output[3594:3594] = '{32'h4634b74a};
test_input[28760:28767] = '{32'h4233c326, 32'hc1b6fc45, 32'h429e3226, 32'h428847cd, 32'h4274e2c1, 32'h420b6ef4, 32'h421b4371, 32'h41dc411b};
test_weights[28760:28767] = '{32'h3f840725, 32'hc20f10a4, 32'h42b43da8, 32'h42c3b53d, 32'hc20e8b87, 32'h421c4a96, 32'h4254ec79, 32'hc20a5b89};
test_bias[3595:3595] = '{32'hc299c8ae};
test_output[3595:3595] = '{32'h46687792};
test_input[28768:28775] = '{32'h427d825c, 32'h41520612, 32'hc2781b41, 32'h4270f4f4, 32'hc2a8d533, 32'h42a5c471, 32'h4261dedd, 32'h427f0cd0};
test_weights[28768:28775] = '{32'h4292a3fd, 32'hc0da8e53, 32'h42ac51ee, 32'h42333a71, 32'h4277a4c8, 32'hc092b872, 32'h42145332, 32'hc2b31ccf};
test_bias[3596:3596] = '{32'h4292c011};
test_output[3596:3596] = '{32'hc5e22a25};
test_input[28776:28783] = '{32'h420044bc, 32'h422c3b50, 32'hc07b57ed, 32'h41695520, 32'h41562cc3, 32'hc2c794b8, 32'hc1b2ec33, 32'hc1a45295};
test_weights[28776:28783] = '{32'hc1ef2a9f, 32'hc28d207d, 32'hc1970ce5, 32'hc2724ca8, 32'h42926bf3, 32'h425116bf, 32'hc21cd275, 32'hc1497a15};
test_bias[3597:3597] = '{32'h4233e168};
test_output[3597:3597] = '{32'hc5f5b035};
test_input[28784:28791] = '{32'h42c2c5e2, 32'hc276e0b9, 32'h42a86051, 32'hc2974736, 32'hc1713c06, 32'hc214a02d, 32'h42a855f1, 32'hc2aec0ee};
test_weights[28784:28791] = '{32'hc21ec0e7, 32'hc1c74922, 32'hc2aa17a9, 32'hc0d8f86a, 32'h4217ec97, 32'hc248fab1, 32'h42a27ee6, 32'hc2410f63};
test_bias[3598:3598] = '{32'hc2a35485};
test_output[3598:3598] = '{32'h454dda5c};
test_input[28792:28799] = '{32'h42ace45c, 32'h42548476, 32'hc2985314, 32'h42bf2274, 32'hc26edcab, 32'hc2b7e525, 32'h42364f74, 32'hc2b09186};
test_weights[28792:28799] = '{32'hc2ba3ed3, 32'hc263e94c, 32'h41b81f5f, 32'h425009b9, 32'h42c16157, 32'hc2b8184f, 32'hc17e66eb, 32'h4266ada2};
test_bias[3599:3599] = '{32'h40f6d8cd};
test_output[3599:3599] = '{32'hc62b89ae};
test_input[28800:28807] = '{32'hc1c93ea7, 32'hc28c4894, 32'hc2c2d48f, 32'hc296651c, 32'h42a017e2, 32'hc14e876a, 32'hc219ad1e, 32'h42352a14};
test_weights[28800:28807] = '{32'hc2999090, 32'hc2bee45a, 32'h42b0b556, 32'hc2c15961, 32'hc211ee86, 32'hc2c70459, 32'hc2ae41ff, 32'hc209c557};
test_bias[3600:3600] = '{32'h42b65f6f};
test_output[3600:3600] = '{32'h45eb5d6b};
test_input[28808:28815] = '{32'h42555a80, 32'hc13f0edb, 32'h42c5e4ae, 32'h42b29c86, 32'hc00c8a1b, 32'hc0a978a7, 32'h4198f3b1, 32'h42c6dabf};
test_weights[28808:28815] = '{32'hc26880e3, 32'h420306f7, 32'hc196dd34, 32'h41f38949, 32'h423f4e72, 32'h429955fa, 32'hc199249c, 32'h4227c9e6};
test_bias[3601:3601] = '{32'h419b6227};
test_output[3601:3601] = '{32'h44289230};
test_input[28816:28823] = '{32'h42a6fcc4, 32'h42b6f569, 32'hc224a70f, 32'hc219d4e1, 32'hc2867779, 32'hc0319e8e, 32'hc1229b4d, 32'h4261574e};
test_weights[28816:28823] = '{32'hc0cd9cfe, 32'h4298ffc0, 32'hc2151315, 32'h428e2fee, 32'h42550913, 32'hc2b48001, 32'h429b12f8, 32'h42ab0386};
test_bias[3602:3602] = '{32'hc2c00475};
test_output[3602:3602] = '{32'h45b742ee};
test_input[28824:28831] = '{32'h42830eb5, 32'h429f1afa, 32'h3fbbdd2f, 32'h429ff469, 32'hc2a6007a, 32'hc29457ac, 32'hc2a84c7b, 32'h421fd3f8};
test_weights[28824:28831] = '{32'hc1f12e87, 32'h4203f485, 32'h4221a501, 32'hc0878eff, 32'hc2a379a9, 32'h41a2f6ec, 32'hc2be46b7, 32'hbfa19ba3};
test_bias[3603:3603] = '{32'h41f47040};
test_output[3603:3603] = '{32'h4654f27e};
test_input[28832:28839] = '{32'h42b908d7, 32'h424deb48, 32'h418f4599, 32'hc2879adc, 32'h4211ca0a, 32'hc2098ec5, 32'h4283893e, 32'h42bdaa84};
test_weights[28832:28839] = '{32'h42680837, 32'hc2979394, 32'h41a1fd2f, 32'hc2067bd3, 32'hc21fdf54, 32'hc2897df8, 32'hc1864ade, 32'h425b1f3d};
test_bias[3604:3604] = '{32'hc2c4b755};
test_output[3604:3604] = '{32'h460cbdb6};
test_input[28840:28847] = '{32'hc1cf8bf0, 32'hc250bb90, 32'hc29ca94c, 32'hc292503e, 32'hc24d95f1, 32'hc2b7f1fd, 32'h4294f550, 32'h4298137e};
test_weights[28840:28847] = '{32'hc1a22819, 32'h42a34c54, 32'hc1e33bd7, 32'hc099f9af, 32'h3f9592ac, 32'h41848977, 32'h42550ced, 32'h425a87dd};
test_bias[3605:3605] = '{32'h41431238};
test_output[3605:3605] = '{32'h45a87ce7};
test_input[28848:28855] = '{32'h428f3b50, 32'hc2b964f3, 32'h4274cf2f, 32'h4263caf6, 32'h422314fe, 32'h42477d5c, 32'h429e6092, 32'h42055ab7};
test_weights[28848:28855] = '{32'h42c351c5, 32'h4147b879, 32'h4229e18f, 32'hc1abb0e1, 32'h4199cd5a, 32'h42353d91, 32'h408d70f3, 32'hc224773d};
test_bias[3606:3606] = '{32'h4252d1fe};
test_output[3606:3606] = '{32'h461125f2};
test_input[28856:28863] = '{32'hc2762b72, 32'h40184c8e, 32'hc226eb48, 32'h42b00d35, 32'hc13b60af, 32'hc0ed33ce, 32'h42b95877, 32'hc295b25f};
test_weights[28856:28863] = '{32'hc1d62599, 32'hc2c56708, 32'h42018ae0, 32'hc2a00d55, 32'hc2ac13ad, 32'hc27aebb5, 32'h428324f9, 32'hc2422372};
test_bias[3607:3607] = '{32'hc1f0c68b};
test_output[3607:3607] = '{32'h458245ad};
test_input[28864:28871] = '{32'hc2c2fdf7, 32'hc17952b2, 32'h424417b6, 32'hc237ab38, 32'hc2a1f693, 32'h4077ee8d, 32'h4083d461, 32'h429f4cf9};
test_weights[28864:28871] = '{32'hc2c78a54, 32'hbfcb5fce, 32'h422dbc21, 32'hc28f88e5, 32'h42c55d90, 32'h42be00f1, 32'hbeda6a8a, 32'hc131dd64};
test_bias[3608:3608] = '{32'hc22b5d5d};
test_output[3608:3608] = '{32'h45cef8a3};
test_input[28872:28879] = '{32'hc2b75c5c, 32'h4247d52f, 32'h424c2dff, 32'h4252791a, 32'h4221c906, 32'h4193751f, 32'hc2664e95, 32'h424db7fd};
test_weights[28872:28879] = '{32'h42c065c8, 32'h3fa6437b, 32'h428a7dce, 32'hc237019f, 32'hc2442b20, 32'hc2b6920b, 32'hc220a0b4, 32'h41bee957};
test_bias[3609:3609] = '{32'h4284e064};
test_output[3609:3609] = '{32'hc5f03d6f};
test_input[28880:28887] = '{32'h427acf98, 32'hc2281200, 32'hc146fa2b, 32'h42ba232c, 32'hc2257661, 32'h429bf3f4, 32'h42945cc1, 32'h42b016eb};
test_weights[28880:28887] = '{32'h42b42f7a, 32'h41313d41, 32'hc1e993a0, 32'hc287d33a, 32'hc2507182, 32'h429937c8, 32'hc2914e42, 32'hc0f1cf01};
test_bias[3610:3610] = '{32'h41ade44e};
test_output[3610:3610] = '{32'h44a54d79};
test_input[28888:28895] = '{32'h42ad56ac, 32'hc242ade9, 32'hc27cb4fe, 32'hc2131895, 32'hc2acc977, 32'h425f6f97, 32'hc280563c, 32'h42c28fab};
test_weights[28888:28895] = '{32'h3d0d732c, 32'hc2bf12f3, 32'hc285438b, 32'hc143d000, 32'hc2852783, 32'hc20a2b5d, 32'h4244d10e, 32'hc2b64eb4};
test_bias[3611:3611] = '{32'hc285dee5};
test_output[3611:3611] = '{32'h44825ead};
test_input[28896:28903] = '{32'hc290734b, 32'hc2b02e3b, 32'hc2817e2a, 32'hc1e47abf, 32'h4180897b, 32'hc2bd9f32, 32'hc1cb8d3f, 32'hc2a48c1d};
test_weights[28896:28903] = '{32'hc29a37f6, 32'h4225ab62, 32'h41f66e22, 32'h41b568af, 32'h423b0308, 32'h4208ba57, 32'hc13b28ff, 32'h4293cea3};
test_bias[3612:3612] = '{32'h42aecb62};
test_output[3612:3612] = '{32'hc60b28e8};
test_input[28904:28911] = '{32'hbf905bfd, 32'hc2373074, 32'hc22d2f83, 32'hc2643054, 32'hc2a0b36f, 32'hc2c07740, 32'hc1fdce41, 32'h414f124d};
test_weights[28904:28911] = '{32'hc283ca9d, 32'h4200d135, 32'h42bcceb6, 32'h42abee09, 32'hc201cb81, 32'h42c668f4, 32'h428633f7, 32'h41682f5a};
test_bias[3613:3613] = '{32'hc23f616e};
test_output[3613:3613] = '{32'hc696f0b1};
test_input[28912:28919] = '{32'hc197190f, 32'h4262f3db, 32'h42ad112e, 32'h42010142, 32'h42bacfad, 32'h41c5d8f3, 32'hc05a7960, 32'hc0f288af};
test_weights[28912:28919] = '{32'hc119ee33, 32'h4276dbfd, 32'h41ce870e, 32'hc2c6ed56, 32'hc2b91f15, 32'h41942624, 32'h4287a3a1, 32'hc2412c44};
test_bias[3614:3614] = '{32'hc2718edf};
test_output[3614:3614] = '{32'hc5a8e15d};
test_input[28920:28927] = '{32'hc293e9b3, 32'hc26d5845, 32'h409b397b, 32'h420bf0cd, 32'hc0a07d13, 32'h426c8048, 32'hc14c343a, 32'hc2b4e93e};
test_weights[28920:28927] = '{32'h41bbe5c8, 32'h411e2a20, 32'hc1ed5e73, 32'h421a1f74, 32'h42829f09, 32'h4133e98e, 32'hc290c37c, 32'hc29289d2};
test_bias[3615:3615] = '{32'h41a73e78};
test_output[3615:3615] = '{32'h45d4309d};
test_input[28928:28935] = '{32'hc24676eb, 32'hc1d3e439, 32'hc13201ae, 32'h422c9506, 32'hc2acc8aa, 32'h42910790, 32'hc1feb3c6, 32'hc29d5768};
test_weights[28928:28935] = '{32'h421cc27e, 32'hc0e056c0, 32'h42a8f7a4, 32'hc29ebdb7, 32'h41104efd, 32'h41df9a35, 32'hc25b501f, 32'h42a968e1};
test_bias[3616:3616] = '{32'hc2a7f43d};
test_output[3616:3616] = '{32'hc61a56d6};
test_input[28936:28943] = '{32'hc1dcb73d, 32'h41162e42, 32'h42b971c5, 32'h4095cb6c, 32'hc1da3d62, 32'hc22aab8c, 32'hc2a6dd07, 32'hc2900f97};
test_weights[28936:28943] = '{32'h427f09ba, 32'h42525b2d, 32'hc05906fb, 32'h3fef9698, 32'h41ed5ffe, 32'hc1c88d14, 32'hc2b9b8fc, 32'h424fe04e};
test_bias[3617:3617] = '{32'h4286e9dd};
test_output[3617:3617] = '{32'h452c8b81};
test_input[28944:28951] = '{32'hbf9d470b, 32'h42afdf22, 32'h3f9c3b19, 32'hc2ab2834, 32'h4234ef56, 32'h4206b13a, 32'hc183e8bf, 32'hc297b7a4};
test_weights[28944:28951] = '{32'hc15b1e59, 32'hc2456691, 32'hc28a981b, 32'hc2a7358a, 32'hc20e87a2, 32'hc29522f6, 32'hc27a8b0e, 32'hc27a488a};
test_bias[3618:3618] = '{32'hc267f608};
test_output[3618:3618] = '{32'h4587cfa2};
test_input[28952:28959] = '{32'h42b6002b, 32'h41c4f6f7, 32'h41b27ef5, 32'hc235e6ac, 32'h414b4e35, 32'h4219acf6, 32'h427dc162, 32'h4267e7a0};
test_weights[28952:28959] = '{32'h42b8f81b, 32'hc297273a, 32'hc0d4e231, 32'hc22c7ad1, 32'h42ad8f00, 32'h41b4f131, 32'h424baf31, 32'h428b0ddc};
test_bias[3619:3619] = '{32'h41e8eba2};
test_output[3619:3619] = '{32'h4689bbbd};
test_input[28960:28967] = '{32'h4286c7d0, 32'hc2754e2f, 32'hc2afb958, 32'h4098aba6, 32'hc2844267, 32'h4230c23b, 32'h4103dd49, 32'hc2a5994e};
test_weights[28960:28967] = '{32'hc21b4b6a, 32'hc1b7c08f, 32'h42b8787b, 32'h421055ca, 32'hc29696f1, 32'h41f78bd4, 32'h42b95a53, 32'hc2a18116};
test_bias[3620:3620] = '{32'hc28e6a3f};
test_output[3620:3620] = '{32'h458f4edd};
test_input[28968:28975] = '{32'h42a6b8e9, 32'h4237c339, 32'h417d81ca, 32'h41ecd092, 32'h4203973b, 32'h41c1e4cd, 32'hc23c4545, 32'h42c2ffd9};
test_weights[28968:28975] = '{32'h41f1f4a9, 32'hc2013440, 32'hc0aa455b, 32'hc23a36b0, 32'h42b84b16, 32'hc1a6db59, 32'hc117cfa4, 32'h41888b64};
test_bias[3621:3621] = '{32'h4252375a};
test_output[3621:3621] = '{32'h458540b0};
test_input[28976:28983] = '{32'hc26a4cab, 32'hc2b499d6, 32'hc2a806c4, 32'hc17df75d, 32'h41bd831d, 32'h42ba6572, 32'h41b2ea6d, 32'hc23d3187};
test_weights[28976:28983] = '{32'h427bd289, 32'hc222545a, 32'hc239bf56, 32'h4283126f, 32'hc190302f, 32'h429a3c4a, 32'h42b8d852, 32'hc2653b00};
test_bias[3622:3622] = '{32'hc2950ddf};
test_output[3622:3622] = '{32'h465f7556};
test_input[28984:28991] = '{32'h4216f3fa, 32'hc1191e99, 32'h42bd8c89, 32'hc27f5319, 32'h40e4c287, 32'hc09671e6, 32'h42ad3bf6, 32'hc22d3c5e};
test_weights[28984:28991] = '{32'hc2aae3ef, 32'h42a8eddc, 32'hc2bd33aa, 32'hc275e671, 32'h42a61894, 32'hc2ae7464, 32'hc2c39502, 32'hc22f816a};
test_bias[3623:3623] = '{32'hc28cb89f};
test_output[3623:3623] = '{32'hc665dd4a};
test_input[28992:28999] = '{32'hc2aa7fac, 32'h4282ece2, 32'hc11eb2e6, 32'h427455b8, 32'h42639859, 32'h429e5b9e, 32'h42506712, 32'h429fe9a3};
test_weights[28992:28999] = '{32'hc2268d22, 32'hc28e170d, 32'hc1343385, 32'hc234dc49, 32'h4299ce3e, 32'hc29ed311, 32'h422e1beb, 32'hc2b2fb4f};
test_bias[3624:3624] = '{32'hc2161da0};
test_output[3624:3624] = '{32'hc6257257};
test_input[29000:29007] = '{32'hc1444375, 32'h42a9cd1b, 32'h426e957e, 32'hc1affa20, 32'h40a9e56c, 32'hc1a1b168, 32'h421a6416, 32'h414a62ba};
test_weights[29000:29007] = '{32'hbf0688be, 32'h41491a3b, 32'hc26d5984, 32'hc2c3cc2f, 32'hc221984a, 32'h42a1efbd, 32'hc1dff1d7, 32'hc18c8df6};
test_bias[3625:3625] = '{32'h4209a14b};
test_output[3625:3625] = '{32'hc55677a5};
test_input[29008:29015] = '{32'hc1e37794, 32'hc1c8288c, 32'h42849deb, 32'hc2b388f6, 32'h42a81907, 32'hc0e5b3a4, 32'h422a2062, 32'hc24a2efb};
test_weights[29008:29015] = '{32'hc2151d36, 32'hc189ce65, 32'hc10a79f8, 32'h4124e330, 32'hc1b7a4d9, 32'hc2b62a50, 32'hc25ce01b, 32'h423e41fa};
test_bias[3626:3626] = '{32'hc2862090};
test_output[3626:3626] = '{32'hc5bebb4e};
test_input[29016:29023] = '{32'hc2bee4f3, 32'hc2333327, 32'hc2c324c6, 32'h411132fe, 32'hc173273d, 32'h4209b2ef, 32'h402d1a43, 32'h42c3c195};
test_weights[29016:29023] = '{32'hc1a7c636, 32'h4295b9e9, 32'hc294ce63, 32'h4285d2fe, 32'h422e5f2b, 32'hc1884cd9, 32'hc20db0e0, 32'hc1d9805b};
test_bias[3627:3627] = '{32'h42adb204};
test_output[3627:3627] = '{32'h45223aae};
test_input[29024:29031] = '{32'h40c7d644, 32'hc2925375, 32'h406fa88d, 32'h42422cf7, 32'hc2a91235, 32'hbfe82787, 32'h42a3d660, 32'h427ead31};
test_weights[29024:29031] = '{32'hc2a8e8cb, 32'h42a14c17, 32'hc2af5c30, 32'h420c9f82, 32'hc1ae9c15, 32'hc2241814, 32'hc21c9599, 32'h42c220ab};
test_bias[3628:3628] = '{32'h421e4063};
test_output[3628:3628] = '{32'hc2ead1dc};
test_input[29032:29039] = '{32'hc25b4cef, 32'hc1992a46, 32'hc224e0d8, 32'hc10cff0a, 32'h42862c09, 32'hc26cc7fd, 32'h42930ed1, 32'h40a593ca};
test_weights[29032:29039] = '{32'h42c2d7c1, 32'h41bf4505, 32'h42bcaf1c, 32'h423f0613, 32'h41f704eb, 32'hc03967ef, 32'hc2a6c523, 32'hc1d0d1d1};
test_bias[3629:3629] = '{32'hc2a324a6};
test_output[3629:3629] = '{32'hc65e1586};
test_input[29040:29047] = '{32'hc2962bd9, 32'h42b3221c, 32'hc2a5fff4, 32'h4079735c, 32'hc281b35e, 32'hc2ae8190, 32'h42030065, 32'h4293de6b};
test_weights[29040:29047] = '{32'h42674a1a, 32'hc1ffb615, 32'h41534693, 32'hc2bd2c71, 32'h41ce03fc, 32'hc22948b4, 32'hc25f2ec5, 32'h42039b8d};
test_bias[3630:3630] = '{32'h427ace7d};
test_output[3630:3630] = '{32'hc5bad4f3};
test_input[29048:29055] = '{32'hc1fe1453, 32'h428e5156, 32'h41b3692f, 32'hc25ec1e5, 32'hc2997eea, 32'h42c1e2cb, 32'hc27d708a, 32'h41f681ef};
test_weights[29048:29055] = '{32'h424cb595, 32'hc0f4c8e8, 32'h4107ef6d, 32'h429c3d3c, 32'h42a5f92b, 32'h41cf50f5, 32'hc2a13981, 32'h4244fad3};
test_bias[3631:3631] = '{32'h410b4659};
test_output[3631:3631] = '{32'hc55e0bc1};
test_input[29056:29063] = '{32'hc2ab96c2, 32'hc2bbc390, 32'h4234b32f, 32'hc0708647, 32'h421cb7e5, 32'h42a73d61, 32'hc2272786, 32'hc2848426};
test_weights[29056:29063] = '{32'hc2a5471a, 32'hc02a4ffb, 32'hc29d153c, 32'hc21eb3b1, 32'hc23f7ff4, 32'hc1a10227, 32'hc2530893, 32'hc1cfc1a9};
test_bias[3632:3632] = '{32'hc2bd3b45};
test_output[3632:3632] = '{32'h4583a73c};
test_input[29064:29071] = '{32'h4292b384, 32'h42babab6, 32'h42aad100, 32'h415bfa59, 32'h41a9d320, 32'hc2c482fc, 32'h415b60db, 32'hc1b4079e};
test_weights[29064:29071] = '{32'h409a2c55, 32'hc2bf0e59, 32'hc291d91d, 32'h42b37a0f, 32'h41bb76f4, 32'hc1020c34, 32'hc290675b, 32'hc2649b31};
test_bias[3633:3633] = '{32'hc2c69dd7};
test_output[3633:3633] = '{32'hc63c8cb2};
test_input[29072:29079] = '{32'hc208f562, 32'hc2ab9018, 32'hc180894d, 32'h429bc456, 32'h42a3fccd, 32'hc1bd76b4, 32'hc2166bc9, 32'hc296f285};
test_weights[29072:29079] = '{32'h41fa94af, 32'h42c22eb6, 32'hc22597b8, 32'h4234ae37, 32'hc2b88ddb, 32'hc2640d51, 32'hc14f4330, 32'h4195dca4};
test_bias[3634:3634] = '{32'hc276b28e};
test_output[3634:3634] = '{32'hc64218e2};
test_input[29080:29087] = '{32'h410d2a88, 32'hc2a44c51, 32'hc05c0a43, 32'hc11d8f61, 32'h42a8a071, 32'h42c33435, 32'h40f1ca5d, 32'h4277a5fe};
test_weights[29080:29087] = '{32'hc298992c, 32'h42beb336, 32'hc2056718, 32'hc296b2f2, 32'h41bfca54, 32'h4242fb9d, 32'hc2174222, 32'hc26d19b1};
test_bias[3635:3635] = '{32'h41e21361};
test_output[3635:3635] = '{32'hc595edfa};
test_input[29088:29095] = '{32'hc1e7f7ef, 32'h42b47775, 32'hc0c751fd, 32'hc2c00c06, 32'h4286cdad, 32'h41f5c77e, 32'hc2a9002d, 32'hc28379f7};
test_weights[29088:29095] = '{32'hc2a0f1a1, 32'hc29ec098, 32'hc2c09cf4, 32'h4226cc1f, 32'hc29ad274, 32'hc1c28483, 32'hc28d0310, 32'h4299e477};
test_bias[3636:3636] = '{32'hc293ea6e};
test_output[3636:3636] = '{32'hc650f183};
test_input[29096:29103] = '{32'h41252672, 32'h40fcd7f4, 32'h42bdb032, 32'h40a152c9, 32'h40afb5cb, 32'hc1de7599, 32'h4288565d, 32'hc28bf636};
test_weights[29096:29103] = '{32'hc0ccefc4, 32'h41f923e0, 32'h42aee1ce, 32'hc2462ecc, 32'hc1064a9d, 32'hc0c4eacb, 32'h429c6fce, 32'h42711188};
test_bias[3637:3637] = '{32'h422c4b03};
test_output[3637:3637] = '{32'h46148839};
test_input[29104:29111] = '{32'hc2195a4c, 32'h423057ea, 32'hc1e6142f, 32'h421f8a06, 32'hc25848a4, 32'h42aa2eb4, 32'h41b96597, 32'hc2761538};
test_weights[29104:29111] = '{32'h40cb7413, 32'h41b13f04, 32'hc29390b1, 32'hc2aeaa6b, 32'hc24c9b3d, 32'h419f7291, 32'h42b3ba87, 32'hc2892e2b};
test_bias[3638:3638] = '{32'h40e11fac};
test_output[3638:3638] = '{32'h461e7b42};
test_input[29112:29119] = '{32'h4137d686, 32'hc1574ae3, 32'hc23b351d, 32'hc00ab024, 32'h424765d9, 32'h410a2f76, 32'hc2c59fb2, 32'hc2c15824};
test_weights[29112:29119] = '{32'hc1564074, 32'hc2028c1b, 32'hc17beae7, 32'h42b00cfc, 32'hc1bf46e3, 32'hc254bfd2, 32'h4195ccb5, 32'hc1813e3c};
test_bias[3639:3639] = '{32'hc2a5a4b5};
test_output[3639:3639] = '{32'hc494e328};
test_input[29120:29127] = '{32'hc0ca0df5, 32'h425c7f07, 32'hc2b756af, 32'hc2010ae7, 32'hc0bc82e6, 32'hc2af3fc9, 32'h422af962, 32'h40912b09};
test_weights[29120:29127] = '{32'h4025ca2d, 32'h422ca611, 32'hc1890adf, 32'hc2badf31, 32'hc19eed33, 32'h425474b5, 32'hc2bd10cd, 32'h42650ecd};
test_bias[3640:3640] = '{32'h419c11f3};
test_output[3640:3640] = '{32'hc4a8dc9f};
test_input[29128:29135] = '{32'hc29831ff, 32'hc2103f41, 32'hc08158d9, 32'hc29554db, 32'h41bd0e7e, 32'h41b6531b, 32'h4140df0f, 32'hc2955a8c};
test_weights[29128:29135] = '{32'h42572ee8, 32'hc2883dd2, 32'h426affaf, 32'h429a9acb, 32'hc18d04e4, 32'h42602b65, 32'hc2ab5184, 32'hc2605c78};
test_bias[3641:3641] = '{32'h42baa4b8};
test_output[3641:3641] = '{32'hc55d06d6};
test_input[29136:29143] = '{32'h4177a58e, 32'h42b6883f, 32'h42a07ee2, 32'h42c20bf9, 32'h42b35081, 32'h4293a898, 32'hc1dc68f3, 32'hc26dfc40};
test_weights[29136:29143] = '{32'h42525343, 32'hc2520806, 32'h422327c2, 32'h41928568, 32'h42bd9364, 32'h423ff3ce, 32'hc1a6fd4d, 32'h42a14e4a};
test_bias[3642:3642] = '{32'h42baf6c5};
test_output[3642:3642] = '{32'h460c5cfa};
test_input[29144:29151] = '{32'hc0b8c6ef, 32'h416d250f, 32'hc27c84c7, 32'hc1c22b04, 32'h424efffd, 32'h3f8c382c, 32'h42c55381, 32'hc2068a17};
test_weights[29144:29151] = '{32'hc265f869, 32'h42651037, 32'h40afa62f, 32'h42bef713, 32'h4239533a, 32'hc194eb3e, 32'h41442a2f, 32'hc283bbf9};
test_bias[3643:3643] = '{32'h42948115};
test_output[3643:3643] = '{32'h45894abb};
test_input[29152:29159] = '{32'h41f5d4c5, 32'h41faaafb, 32'hc23bbd1a, 32'h4205d769, 32'hc2c3ecc0, 32'hc2244187, 32'hc08e53f6, 32'hc2608933};
test_weights[29152:29159] = '{32'hc285de0e, 32'hc24d2f7b, 32'hc24d5128, 32'h4290705f, 32'hc07c6da7, 32'hc2b8a589, 32'h42b1c5b8, 32'h42711efc};
test_bias[3644:3644] = '{32'hc27c879d};
test_output[3644:3644] = '{32'h44bb1a30};
test_input[29160:29167] = '{32'h3e87f77c, 32'h429658fb, 32'h413b3396, 32'h429cff2a, 32'hc1d61b75, 32'hc220325e, 32'hc246fa56, 32'hc2bb509b};
test_weights[29160:29167] = '{32'h42c28aa9, 32'hc258373b, 32'h42b3e759, 32'hc297dfc7, 32'hc19f573e, 32'h42a81ee2, 32'h420bf93d, 32'h4293bc92};
test_bias[3645:3645] = '{32'hc28e8217};
test_output[3645:3645] = '{32'hc6a03bc3};
test_input[29168:29175] = '{32'hbfae0ea7, 32'hc143a68b, 32'hc2aa07f0, 32'hc145d927, 32'h421e7d31, 32'h3f8a8f17, 32'h417cbf11, 32'h42c01f36};
test_weights[29168:29175] = '{32'h41972ded, 32'h411c6fb2, 32'hc21033e1, 32'hc28d470d, 32'h429f2fe2, 32'hc22d28b4, 32'h42861ec8, 32'hc2c4bf52};
test_bias[3646:3646] = '{32'hc25c260c};
test_output[3646:3646] = '{32'hc4c13588};
test_input[29176:29183] = '{32'hc28f9403, 32'hc255f2df, 32'h42c49824, 32'hc0cc4fcc, 32'hc23487dc, 32'h42ab7f9f, 32'hc19389ca, 32'hc2921176};
test_weights[29176:29183] = '{32'h423b6bfa, 32'hc2a8e174, 32'hc28378ca, 32'hc20febf3, 32'hc0965a10, 32'h42a9a220, 32'h423e14c4, 32'hc11b1ce0};
test_bias[3647:3647] = '{32'h41359725};
test_output[3647:3647] = '{32'h450c8dba};
test_input[29184:29191] = '{32'h42bc1c02, 32'hc1dd4056, 32'h42460a04, 32'hc29481e7, 32'h42299172, 32'hc2598c38, 32'hc1e11572, 32'hc1557a82};
test_weights[29184:29191] = '{32'hc2750c57, 32'hc2489428, 32'hc22178b3, 32'hc24532af, 32'hc22a3ee9, 32'hc262b7c6, 32'hc2581d72, 32'h42a3ea55};
test_bias[3648:3648] = '{32'h41868bce};
test_output[3648:3648] = '{32'hc477d3cf};
test_input[29192:29199] = '{32'hc28c51b1, 32'hc2b78ad7, 32'hc2c7e445, 32'hc02c4d56, 32'hc2490a49, 32'hc29117f4, 32'hc2758f21, 32'h429d9ffb};
test_weights[29192:29199] = '{32'h41fa7157, 32'h422e7d23, 32'h41a4ef54, 32'h425aebdb, 32'hc2a317be, 32'h41fb642b, 32'hc2a27759, 32'hc236dda6};
test_bias[3649:3649] = '{32'h41453653};
test_output[3649:3649] = '{32'hc5a24458};
test_input[29200:29207] = '{32'h41ba63b3, 32'h4263e549, 32'hc2251e21, 32'h4184a160, 32'h422c09ff, 32'h403c2a0f, 32'hc2c5c9c6, 32'hc26023d1};
test_weights[29200:29207] = '{32'h41c525be, 32'hc2bfd1cd, 32'h42c3de51, 32'h424dff9b, 32'hc1de0fb3, 32'hc2ae6b92, 32'hc255408d, 32'hc19908e7};
test_bias[3650:3650] = '{32'h424986f6};
test_output[3650:3650] = '{32'hc543ead5};
test_input[29208:29215] = '{32'h42955674, 32'hc2980d6c, 32'hc28fd6b7, 32'h41115f24, 32'hbf82b1fb, 32'h428c3842, 32'hc29fb042, 32'h41bf82ae};
test_weights[29208:29215] = '{32'h429f5c2b, 32'hc21b8d89, 32'hc28d9957, 32'h4292a2c2, 32'hc2a135ca, 32'h4203144d, 32'hc2c2832b, 32'hc20d35a2};
test_bias[3651:3651] = '{32'h412513dd};
test_output[3651:3651] = '{32'h46bb4cff};
test_input[29216:29223] = '{32'h42494500, 32'hc1c054bf, 32'hc2b819a0, 32'hc161c4ab, 32'hc280be0b, 32'h42a9b0f6, 32'hbfa6e3e7, 32'h42c15e01};
test_weights[29216:29223] = '{32'h42c69640, 32'h420fdb88, 32'hc1bc7af3, 32'h4105654e, 32'h4154cefd, 32'hc191de3a, 32'h42c2fb58, 32'h41c963aa};
test_bias[3652:3652] = '{32'hc2313318};
test_output[3652:3652] = '{32'h45bccf06};
test_input[29224:29231] = '{32'hc15323ad, 32'hc1b53fcf, 32'h4281b6b6, 32'h4194c86e, 32'hc17678b1, 32'hc2b66803, 32'h4272ea19, 32'h41d53b45};
test_weights[29224:29231] = '{32'hc2b5178e, 32'hbb957a47, 32'h42a1ba79, 32'hc2a2ac24, 32'hc28d1939, 32'h4207b812, 32'h41be2283, 32'h41de5a89};
test_bias[3653:3653] = '{32'h3f8c37cb};
test_output[3653:3653] = '{32'h459f8341};
test_input[29232:29239] = '{32'h4244fadf, 32'h429f3d2c, 32'h427cf30b, 32'h4212f221, 32'hc24cd9b4, 32'hc2078198, 32'h4296c22d, 32'hc11976f3};
test_weights[29232:29239] = '{32'h42543906, 32'h427a86ee, 32'hc1bcb787, 32'h40554df7, 32'h42b96de1, 32'hc2b0c8f9, 32'h41f76652, 32'hc2934344};
test_bias[3654:3654] = '{32'hc2937728};
test_output[3654:3654] = '{32'h45e8801b};
test_input[29240:29247] = '{32'h41204f7d, 32'hc14c14e8, 32'h4221bc6d, 32'h418b7803, 32'h42a9bcd5, 32'hc29b606b, 32'hc1d8b8cd, 32'hc2302515};
test_weights[29240:29247] = '{32'h42b328b2, 32'h425a2aa8, 32'hc25c4931, 32'hc1cb31df, 32'h42791b72, 32'h41e32845, 32'hc2aef03d, 32'h42c64ec4};
test_bias[3655:3655] = '{32'h4287f49e};
test_output[3655:3655] = '{32'hc4a4a383};
test_input[29248:29255] = '{32'h42545116, 32'hc2b3ef96, 32'hc1b5e258, 32'hc20a8efd, 32'hc1caae9f, 32'h429ce0db, 32'hc2918328, 32'h428a1e7b};
test_weights[29248:29255] = '{32'h413018e9, 32'h42aad787, 32'hc2b6741f, 32'hc228c9fa, 32'h4237f9b5, 32'h42aeb08c, 32'hc24d8e46, 32'h41e81eaf};
test_bias[3656:3656] = '{32'h422e148c};
test_output[3656:3656] = '{32'h45f717b6};
test_input[29256:29263] = '{32'h41bdaf6e, 32'hc183ef57, 32'h425f4d6b, 32'hc2271d7b, 32'hc2b72459, 32'h42146539, 32'h42700506, 32'hc26a0103};
test_weights[29256:29263] = '{32'hc1dc0d8a, 32'h42aa3d5e, 32'h41f6e7bb, 32'h40826b2b, 32'h42be68a7, 32'hc28a588a, 32'h42c16a03, 32'h412e1dc8};
test_bias[3657:3657] = '{32'hbf4158ea};
test_output[3657:3657] = '{32'hc5ceefdb};
test_input[29264:29271] = '{32'hc2692c74, 32'hc0222cd9, 32'hc2767e17, 32'h429db2be, 32'h428b67dc, 32'hc16c36a3, 32'h426f6432, 32'h42930855};
test_weights[29264:29271] = '{32'h4197987c, 32'h40c8f8b8, 32'hc1e8ed35, 32'h4261069d, 32'h41e72ee8, 32'h40f5cd3d, 32'h41c9e2fd, 32'hbe846999};
test_bias[3658:3658] = '{32'hc2931f2b};
test_output[3658:3658] = '{32'h4603b027};
test_input[29272:29279] = '{32'hc26d983a, 32'hc24c6788, 32'h4249ac00, 32'hc29b3690, 32'hc2738418, 32'hc269f7fd, 32'h42a5ffe2, 32'h41cb6558};
test_weights[29272:29279] = '{32'hc21782a9, 32'hc1f2cb8d, 32'h41ede0fc, 32'h41181303, 32'hc217faa6, 32'h408834a4, 32'h41ea2a3b, 32'hc2c68878};
test_bias[3659:3659] = '{32'h42bb59cd};
test_output[3659:3659] = '{32'h45cf0e15};
test_input[29280:29287] = '{32'h41787120, 32'hc122643d, 32'h4290e551, 32'h428dfa9c, 32'hc285c63d, 32'hc17a5dbd, 32'hc212b871, 32'hc282ff63};
test_weights[29280:29287] = '{32'hc2bc1017, 32'h3fdd342a, 32'hc19f2e08, 32'h42a51184, 32'h40b3b93c, 32'hbe8b55a6, 32'h42229c8d, 32'h42c0e610};
test_bias[3660:3660] = '{32'hc2bfd70c};
test_output[3660:3660] = '{32'hc5a6bf19};
test_input[29288:29295] = '{32'hc29b7370, 32'h4246eea0, 32'hc23d590d, 32'h4174ff56, 32'hc1df7e00, 32'hc1a21af5, 32'hc16d854a, 32'h3fd834d3};
test_weights[29288:29295] = '{32'h421ecd26, 32'hc20c4a38, 32'h40b3056b, 32'h41e9dc3a, 32'hc2590b3b, 32'h42a8cf38, 32'hc28a7615, 32'h41b21ba1};
test_bias[3661:3661] = '{32'hc282f55a};
test_output[3661:3661] = '{32'hc5701c73};
test_input[29296:29303] = '{32'hc29420c1, 32'hc1972858, 32'h42b87327, 32'hc28219fc, 32'hc24153e5, 32'hc1f2f974, 32'hc26ad825, 32'h42691468};
test_weights[29296:29303] = '{32'h42967dce, 32'h413b0a28, 32'hc257ad49, 32'hc2a91e43, 32'h408a12d9, 32'h4215837b, 32'hc264cc03, 32'h3e554f07};
test_bias[3662:3662] = '{32'hc1a49501};
test_output[3662:3662] = '{32'hc54bbef5};
test_input[29304:29311] = '{32'hc28b1189, 32'h42212180, 32'h42c56794, 32'h422995ec, 32'h4233ee8a, 32'h41e1850d, 32'h421db3b0, 32'h41f846e9};
test_weights[29304:29311] = '{32'hc2812306, 32'hc28e5964, 32'h429a3c21, 32'h4282254d, 32'hc2904b08, 32'hc254c57b, 32'hc2074cee, 32'h41fd9493};
test_bias[3663:3663] = '{32'hc29f2bd8};
test_output[3663:3663] = '{32'h45d516a0};
test_input[29312:29319] = '{32'hc2892f76, 32'h408f0dbd, 32'hc299945c, 32'hc2ad8717, 32'h428eac0a, 32'hc2745081, 32'h42233b8a, 32'hc2408d06};
test_weights[29312:29319] = '{32'hc1c4687b, 32'hc2a11638, 32'hc2bc5318, 32'hc2713d5e, 32'hc2b5b954, 32'hc2c3f3c0, 32'h3ff3a3ba, 32'hc2b1f03a};
test_bias[3664:3664] = '{32'hc257eed3};
test_output[3664:3664] = '{32'h468978b7};
test_input[29320:29327] = '{32'h42687659, 32'h41cb4344, 32'hc1d2f28c, 32'hc21e1cd5, 32'h4283cc11, 32'hc2c7d680, 32'h41025ee2, 32'hc284635d};
test_weights[29320:29327] = '{32'h41daaa71, 32'hc2ae4dab, 32'h42c67527, 32'hc2497fb6, 32'h429312b7, 32'h429757e5, 32'h423fddde, 32'hc24fc02b};
test_bias[3665:3665] = '{32'hc1014035};
test_output[3665:3665] = '{32'hc3117ddb};
test_input[29328:29335] = '{32'hc2a9a05e, 32'h425b96b4, 32'h42c40f7f, 32'hc294d988, 32'hc0c27d65, 32'hc21fa431, 32'h4297ed1f, 32'h3feb4be7};
test_weights[29328:29335] = '{32'h428fe41e, 32'hc28bfcea, 32'h421e1201, 32'h429756a9, 32'h42a2be24, 32'h42a6d012, 32'h42935eb5, 32'h42a5e1ad};
test_bias[3666:3666] = '{32'hc24cc35c};
test_output[3666:3666] = '{32'hc6198b84};
test_input[29336:29343] = '{32'hc2c5eb0a, 32'h42a4e793, 32'hc176a861, 32'h42463d06, 32'hc28e0d72, 32'h427bb040, 32'hc2acff4c, 32'h3fffa598};
test_weights[29336:29343] = '{32'h41c5a17d, 32'h42bafaf6, 32'h41e6c95b, 32'h410e1b88, 32'h42a17fd2, 32'hc27047c7, 32'h41efcc67, 32'hc215dd63};
test_bias[3667:3667] = '{32'hc2aa0320};
test_output[3667:3667] = '{32'hc5db038d};
test_input[29344:29351] = '{32'h42ae093a, 32'h4281d1aa, 32'hc2279bd6, 32'hc2168935, 32'hc1e68a94, 32'hc2c4466e, 32'h42bab5f8, 32'h42293caf};
test_weights[29344:29351] = '{32'h427334fd, 32'h42a2db80, 32'hc2b406be, 32'hc24db9e1, 32'hc292d12e, 32'hc1e0ff98, 32'hc2a64043, 32'h40bbb740};
test_bias[3668:3668] = '{32'hc245a644};
test_output[3668:3668] = '{32'h4654772a};
test_input[29352:29359] = '{32'h42c02361, 32'hc28bb0e7, 32'hc1ad8e9a, 32'h4273781a, 32'h4209ee7b, 32'h4290e417, 32'hc2147a05, 32'hc2ad11d0};
test_weights[29352:29359] = '{32'h42c73e1e, 32'h42a665a2, 32'hc222fd33, 32'hc2a2d531, 32'h3fe19ccc, 32'h4253cba7, 32'h4246b323, 32'hc2aba366};
test_bias[3669:3669] = '{32'h411c1e52};
test_output[3669:3669] = '{32'h460f6324};
test_input[29360:29367] = '{32'hc20b024b, 32'hc2724be3, 32'hc2386758, 32'hc2b103fb, 32'hc271fa03, 32'hc113e002, 32'hc28315be, 32'h40b6b06e};
test_weights[29360:29367] = '{32'hc2a3448c, 32'hc107cf50, 32'h41cb98b5, 32'hc22b27ce, 32'hc1c78ec0, 32'h428a7710, 32'h41b6867b, 32'h4184a3cb};
test_bias[3670:3670] = '{32'h42a86133};
test_output[3670:3670] = '{32'h45ac6cf3};
test_input[29368:29375] = '{32'h429d5710, 32'h3fd97142, 32'h424284ad, 32'hc29600f7, 32'hc19ae3f0, 32'h429f399c, 32'h42b9301c, 32'hc284ad1a};
test_weights[29368:29375] = '{32'hc28c8732, 32'h42bff597, 32'h4209aa88, 32'hc2c14c9c, 32'h42b4e152, 32'h42af2e3b, 32'hc283edf2, 32'hc2a26276};
test_bias[3671:3671] = '{32'h423a07e1};
test_output[3671:3671] = '{32'h45fd472b};
test_input[29376:29383] = '{32'h41a2c8be, 32'hc21c27ea, 32'h42c79949, 32'hc2b7b1de, 32'h42782827, 32'h41a36d5b, 32'h40aefceb, 32'hc1f1241a};
test_weights[29376:29383] = '{32'hc29c4bce, 32'hc1ce4149, 32'h4281b6ce, 32'hc2504c3c, 32'hc17533bc, 32'hc2a41ccc, 32'h429a02eb, 32'hc28cb837};
test_bias[3672:3672] = '{32'h429b96f0};
test_output[3672:3672] = '{32'h4626a279};
test_input[29384:29391] = '{32'hc07f0821, 32'h412ae73a, 32'hc1e24f24, 32'h42629146, 32'h41942996, 32'hc0660075, 32'hc25ad1f0, 32'hc2852188};
test_weights[29384:29391] = '{32'hc0c7c261, 32'h41b1b381, 32'h418daa30, 32'hc2b90d4b, 32'hc28b6fc4, 32'hc29ab7ed, 32'h40a31d38, 32'h42909fef};
test_bias[3673:3673] = '{32'h42abcc42};
test_output[3673:3673] = '{32'hc633ad2c};
test_input[29392:29399] = '{32'hc26bf9e4, 32'hc208fb04, 32'hc2ab32d5, 32'hc125ef29, 32'hc2342526, 32'h427be5a0, 32'h42a40c56, 32'hc251ced1};
test_weights[29392:29399] = '{32'hc2afc363, 32'h427442aa, 32'hc2bab655, 32'h410a1083, 32'h41fc6bb3, 32'h4296ce0e, 32'h4281f023, 32'hc19e6662};
test_bias[3674:3674] = '{32'h426fe942};
test_output[3674:3674] = '{32'h46a21bf9};
test_input[29400:29407] = '{32'h41c2537f, 32'hc18e7027, 32'h42a01bb3, 32'h41fe5004, 32'hc00fbb54, 32'hc00fb735, 32'h4235e1a7, 32'hc2884f0e};
test_weights[29400:29407] = '{32'h429c68eb, 32'hc2b1dd3c, 32'hc1c6f8be, 32'hc1f7b8b1, 32'h42ae5f98, 32'hc2aeedbd, 32'hc27cc1f0, 32'hc1165dbb};
test_bias[3675:3675] = '{32'h41d0b772};
test_output[3675:3675] = '{32'hc4d44c7d};
test_input[29408:29415] = '{32'h42773d17, 32'h409c9f13, 32'hc211c1ca, 32'hc296a337, 32'hc23df8a5, 32'h419119ab, 32'h421d8b02, 32'h42991677};
test_weights[29408:29415] = '{32'h40762b35, 32'hc1fed55e, 32'h4283e51b, 32'h40f2dc0c, 32'hc2244340, 32'h41b541fe, 32'h42aef8cb, 32'h4168cad3};
test_bias[3676:3676] = '{32'h422a823e};
test_output[3676:3676] = '{32'h457e6696};
test_input[29416:29423] = '{32'hc1708ea0, 32'h4145c45e, 32'hc217e7c7, 32'hc2a37949, 32'hc27e86f5, 32'h40de8ee5, 32'hbf836ce0, 32'h42a89bbb};
test_weights[29416:29423] = '{32'hc261c701, 32'h4273ec89, 32'h4141fc8c, 32'h41514c14, 32'h41b26047, 32'h42b7203c, 32'hc20718a0, 32'h4274ad9d};
test_bias[3677:3677] = '{32'hc2b1dc9c};
test_output[3677:3677] = '{32'h45894ad8};
test_input[29424:29431] = '{32'hc2b6162a, 32'h423eaee0, 32'h42c48038, 32'h42b73337, 32'h428b3a29, 32'h4242145d, 32'hc28350b2, 32'hbe007a15};
test_weights[29424:29431] = '{32'hc27a19ab, 32'hc1e778b0, 32'hbf4b95e0, 32'hc29fb2f5, 32'h41d02dac, 32'h429d49cc, 32'hc147399e, 32'h427f9b25};
test_bias[3678:3678] = '{32'hc2a639f4};
test_output[3678:3678] = '{32'h454ca8d2};
test_input[29432:29439] = '{32'hc2149da6, 32'h41ee9c14, 32'h41ace447, 32'h41b85ccf, 32'hc0806e1d, 32'hc0b99711, 32'hc13dfa98, 32'hc12ddaee};
test_weights[29432:29439] = '{32'hc27d6b1a, 32'h3fd85b0a, 32'hc163d271, 32'hc2b8a2ca, 32'hc1d087e5, 32'hc24341c3, 32'h429cf7df, 32'h3f9bc52a};
test_bias[3679:3679] = '{32'h4274f076};
test_output[3679:3679] = '{32'hc403c5df};
test_input[29440:29447] = '{32'hc2c21d36, 32'hc1af4325, 32'h42bdfee6, 32'h414293b0, 32'hc1cafb57, 32'hc2428bea, 32'hc26c4643, 32'h428868fb};
test_weights[29440:29447] = '{32'hc255f3e4, 32'h41ac74df, 32'h42b92253, 32'hc2148f58, 32'hc11c50c2, 32'h42b7aea7, 32'h40c38d4f, 32'hc1ce48dd};
test_bias[3680:3680] = '{32'h40ac4605};
test_output[3680:3680] = '{32'h45d23f29};
test_input[29448:29455] = '{32'hc28b1cdb, 32'hc21d1555, 32'h420cdd3c, 32'hc28284da, 32'hc132ab7e, 32'h42c3248c, 32'h4250c21e, 32'hc2c5ba09};
test_weights[29448:29455] = '{32'h4007c059, 32'h4215ce5e, 32'hc28b44de, 32'hc239834d, 32'hc10b04f1, 32'h422c6510, 32'hc279543e, 32'h42198a87};
test_bias[3681:3681] = '{32'hc1d2c0b7};
test_output[3681:3681] = '{32'hc56e808d};
test_input[29456:29463] = '{32'hc2934c90, 32'hc2a2d783, 32'hc2ad8ef8, 32'hc2afdd03, 32'h412b0e29, 32'h424f0ccb, 32'h42302d4f, 32'hc296360f};
test_weights[29456:29463] = '{32'hc24800fb, 32'hc22b10cc, 32'hc20b4d09, 32'h420354f3, 32'hc2359d6d, 32'hc274efb6, 32'h421d9234, 32'hbe22e826};
test_bias[3682:3682] = '{32'h4278520e};
test_output[3682:3682] = '{32'h45aa6d89};
test_input[29464:29471] = '{32'hc2a9aa81, 32'h3fb7fcba, 32'h426be3a2, 32'hc1d0e4e3, 32'h4233969c, 32'hc1dc4d65, 32'h42547cf8, 32'hc10b8e36};
test_weights[29464:29471] = '{32'h4257e829, 32'hc18021f2, 32'hc1cc422f, 32'hc1f2eff3, 32'hc2373b99, 32'h4239a322, 32'h422e16d2, 32'hc2bc3b85};
test_bias[3683:3683] = '{32'hc1f0ed4e};
test_output[3683:3683] = '{32'hc5ad5565};
test_input[29472:29479] = '{32'hbd5354e9, 32'h422d258b, 32'h40cbdf18, 32'hc2b86900, 32'hc070196b, 32'hc20c5bee, 32'h428a67bf, 32'h41897f02};
test_weights[29472:29479] = '{32'h4236f88f, 32'h42c42054, 32'h42251a28, 32'h4292b6bd, 32'hc22686d1, 32'hc2925c3d, 32'hc22bbda3, 32'h42c5ae59};
test_bias[3684:3684] = '{32'hc2c69f45};
test_output[3684:3684] = '{32'hc46289fb};
test_input[29480:29487] = '{32'hc281e46d, 32'h41a76d68, 32'h411beac0, 32'hc2c25f37, 32'hc2870dd6, 32'hc15aaa9e, 32'h419d3496, 32'hc2806998};
test_weights[29480:29487] = '{32'hc2b62146, 32'hc27e70ac, 32'hc21895e9, 32'h42a9a3ef, 32'h42538be9, 32'hc26da2a7, 32'h42787770, 32'hc204d82e};
test_bias[3685:3685] = '{32'h42ada810};
test_output[3685:3685] = '{32'hc5517884};
test_input[29488:29495] = '{32'hc2894491, 32'h4233fddb, 32'hc1adf001, 32'h4110fd35, 32'hc2270a07, 32'hc2bde86f, 32'h42a4dbdd, 32'h428a7715};
test_weights[29488:29495] = '{32'h414c4518, 32'hc1105951, 32'h4291871a, 32'hc2bb0c57, 32'hc16166fc, 32'h4275b72b, 32'hc28cd76d, 32'h4195889c};
test_bias[3686:3686] = '{32'h42b1041f};
test_output[3686:3686] = '{32'hc6510a19};
test_input[29496:29503] = '{32'hc116cce2, 32'h42b15127, 32'h41d234d4, 32'hc281eaac, 32'hc18e6ebe, 32'hc286dab2, 32'hc28a2451, 32'hc269252c};
test_weights[29496:29503] = '{32'hc2027dfe, 32'h421f0136, 32'hc1cd5a4f, 32'hc29f899c, 32'h423905b1, 32'hc2048a22, 32'hc13776bd, 32'hc29fd166};
test_bias[3687:3687] = '{32'h422aa4ab};
test_output[3687:3687] = '{32'h466e275b};
test_input[29504:29511] = '{32'hc29d3338, 32'h42b5d2ba, 32'h408b8cd7, 32'h429fd91c, 32'h42b2df8c, 32'h41df264a, 32'hc2828dee, 32'hc2bcec80};
test_weights[29504:29511] = '{32'h423c4c60, 32'hc2859f3b, 32'hc2929125, 32'hc24e24ad, 32'hc2b3ab3c, 32'hc0078e93, 32'hc2b54e5a, 32'h40ce2656};
test_bias[3688:3688] = '{32'h421da7da};
test_output[3688:3688] = '{32'hc6847b39};
test_input[29512:29519] = '{32'hc121202f, 32'h4209a440, 32'h40927234, 32'h41ba0e0d, 32'h4279f2f2, 32'hc2867626, 32'h420b5401, 32'hc2a3e193};
test_weights[29512:29519] = '{32'hc2ad3c85, 32'h425f43cb, 32'hc23d8d16, 32'hc1e1da68, 32'hc1e195c1, 32'h4286ef2c, 32'hc28e8f9a, 32'hc2870839};
test_bias[3689:3689] = '{32'h424956fa};
test_output[3689:3689] = '{32'hc49fd368};
test_input[29520:29527] = '{32'h42bdc623, 32'hc21861ba, 32'h4034daa8, 32'h42b49486, 32'h4237764e, 32'hc04d0f85, 32'h427c064e, 32'h4235a8d0};
test_weights[29520:29527] = '{32'hc28872d8, 32'hc28e3240, 32'hc0a5145d, 32'hc08dc6ea, 32'hc298cceb, 32'h41e6761e, 32'hc29f4d5c, 32'h428ebe14};
test_bias[3690:3690] = '{32'h429314d9};
test_output[3690:3690] = '{32'hc6141f26};
test_input[29528:29535] = '{32'h42c7b91c, 32'h42b00b99, 32'hc2c64447, 32'h4223adbb, 32'hc263a809, 32'h41a9c0b6, 32'h41a3704d, 32'hc2b6f5e4};
test_weights[29528:29535] = '{32'h4232c0da, 32'hc297c442, 32'h42ad709c, 32'hc1cc068f, 32'hc28fc7a8, 32'hc22596a1, 32'hc1220427, 32'hc2884f94};
test_bias[3691:3691] = '{32'hc2205801};
test_output[3691:3691] = '{32'hc52602a8};
test_input[29536:29543] = '{32'h421709a8, 32'hc2a62ef2, 32'h426076c2, 32'hc281b92f, 32'hc2ab4f0b, 32'hc27ee53c, 32'hc28588ad, 32'hc28b4494};
test_weights[29536:29543] = '{32'hc24c84cd, 32'hc0732eed, 32'h422f4b94, 32'hc2a0a0c7, 32'h41c9245b, 32'h3e5ad177, 32'hc27f0c92, 32'hc0358bf9};
test_bias[3692:3692] = '{32'h41f4b49c};
test_output[3692:3692] = '{32'h4602cef8};
test_input[29544:29551] = '{32'hc2c67b88, 32'h42177bb0, 32'h422055ef, 32'hc23bd7c5, 32'hc21fce8c, 32'hc1a76e85, 32'hc28f7175, 32'h41869fde};
test_weights[29544:29551] = '{32'h42a480a4, 32'hc286e675, 32'h42181a5a, 32'hc2496cc2, 32'h415f0bae, 32'hc2709de1, 32'hc2a79455, 32'hc1e43948};
test_bias[3693:3693] = '{32'hc2b64bdf};
test_output[3693:3693] = '{32'hc42bf256};
test_input[29552:29559] = '{32'hc224618a, 32'hc2325ec2, 32'h4248e43f, 32'hbffbbba7, 32'h42638364, 32'hc1ef4d3a, 32'hc26b5c5e, 32'hc2b4d55e};
test_weights[29552:29559] = '{32'hc27c8ce7, 32'h42530877, 32'h41eabae8, 32'h4280cafa, 32'h41f2f57a, 32'hc2c46846, 32'hc288f318, 32'hc101056a};
test_bias[3694:3694] = '{32'hc2969bee};
test_output[3694:3694] = '{32'h462ae321};
test_input[29560:29567] = '{32'hc26981ab, 32'hc0fca8c7, 32'h423b0ade, 32'h42250f59, 32'hc2549179, 32'hc10e870b, 32'h429e468f, 32'hc2797905};
test_weights[29560:29567] = '{32'hc29dc132, 32'h42bf3a9a, 32'hc2c40ec4, 32'hc2a904e9, 32'hc2a875a7, 32'h41feab07, 32'h4285cc3d, 32'hc29d8296};
test_bias[3695:3695] = '{32'h429a7714};
test_output[3695:3695] = '{32'h46203953};
test_input[29568:29575] = '{32'h4225b448, 32'h425ce665, 32'hc25d0121, 32'h4266059f, 32'hc24727cf, 32'hc18c12fe, 32'h418b2bf8, 32'hc045bcba};
test_weights[29568:29575] = '{32'h42c7068f, 32'hc190bd6f, 32'hc24a33b6, 32'hc1b86a0c, 32'hc2983ec9, 32'h423fd79e, 32'h41f6b747, 32'h42c61a13};
test_bias[3696:3696] = '{32'h41efd3b5};
test_output[3696:3696] = '{32'h45f3cb0e};
test_input[29576:29583] = '{32'h426bb035, 32'hc2593184, 32'h425fb5a3, 32'h42c2c3a2, 32'h42acba9a, 32'h41fa58a6, 32'hc18ed1f3, 32'h42448274};
test_weights[29576:29583] = '{32'h4260c699, 32'hc2ad24ed, 32'hc23e1e2c, 32'hc254514e, 32'hc2c7ad05, 32'h40ebc221, 32'hc28302bd, 32'hc28f72f3};
test_bias[3697:3697] = '{32'h42946da5};
test_output[3697:3697] = '{32'hc623dd1f};
test_input[29584:29591] = '{32'h42457e86, 32'h42105961, 32'h41d0a5f4, 32'hc1a126e3, 32'h42631a8d, 32'h42881c6f, 32'hc2745374, 32'hc2bdc8ff};
test_weights[29584:29591] = '{32'h42963090, 32'hc1fba8a8, 32'h42acb287, 32'hc123c16c, 32'h4216e6d6, 32'h42acec00, 32'h41ac7db9, 32'h41bf55cf};
test_bias[3698:3698] = '{32'hc2091e19};
test_output[3698:3698] = '{32'h46136fc8};
test_input[29592:29599] = '{32'hc1b7e54c, 32'hc2919289, 32'hc22bed40, 32'h42871ad5, 32'hc1c700ad, 32'hc1fd6b18, 32'h424ca3a6, 32'h428f31a6};
test_weights[29592:29599] = '{32'h4208158f, 32'h4292cdd7, 32'hc253cd83, 32'h424be8e2, 32'h401803cb, 32'hc2a7dd2a, 32'h428316cb, 32'hc1b9be04};
test_bias[3699:3699] = '{32'h42c6fac7};
test_output[3699:3699] = '{32'h45790ed6};
test_input[29600:29607] = '{32'h429e101c, 32'hc2509318, 32'hc1b5db4d, 32'h409d5307, 32'hc2a21750, 32'h42587959, 32'h4218a5c1, 32'hc1adf0f8};
test_weights[29600:29607] = '{32'h428fb479, 32'hc1650404, 32'hc2b89eed, 32'h42596c19, 32'hc1d51679, 32'h425feda7, 32'h41b17d23, 32'hc294c243};
test_bias[3700:3700] = '{32'h4241a978};
test_output[3700:3700] = '{32'h4680d691};
test_input[29608:29615] = '{32'hc121e2b4, 32'h41239106, 32'h42415715, 32'hc1a5f76f, 32'hc22ac73f, 32'h4258cf88, 32'hc1164ffa, 32'hc1d09664};
test_weights[29608:29615] = '{32'h4179f149, 32'h4259fef8, 32'hc2b02fc7, 32'h41942af4, 32'hc28caeb7, 32'hc29b04a6, 32'hc16cd60a, 32'h419d9d05};
test_bias[3701:3701] = '{32'h418ba26c};
test_output[3701:3701] = '{32'hc5b532a1};
test_input[29616:29623] = '{32'h418087fc, 32'h42a1bd99, 32'h41be79b9, 32'h3ea59491, 32'hc0fd81c0, 32'h421ac72a, 32'hc22602a3, 32'h42c0f700};
test_weights[29616:29623] = '{32'h3f4e9925, 32'hc03df17c, 32'hc24b7cd2, 32'h411c3f18, 32'hc29a92f5, 32'hc10f0a0b, 32'hc2b87f43, 32'h42014915};
test_bias[3702:3702] = '{32'hc1e3bd9c};
test_output[3702:3702] = '{32'h45b3ae10};
test_input[29624:29631] = '{32'hc1e26306, 32'hc28d3e24, 32'hc2c424b8, 32'hc1d9264b, 32'hc2ae9cc3, 32'h42bb490a, 32'h4240acbe, 32'hc25fb7b9};
test_weights[29624:29631] = '{32'h42002a03, 32'hc2952f71, 32'hc2aa933e, 32'h42994e4d, 32'hc2a96833, 32'h4189b8c1, 32'h40c24576, 32'hc2c3b1e6};
test_bias[3703:3703] = '{32'h423e0612};
test_output[3703:3703] = '{32'h46c6f0fb};
test_input[29632:29639] = '{32'h42af45fe, 32'hc275b023, 32'hc220868a, 32'h418a8930, 32'h41e7e87e, 32'hc18a0e68, 32'hc1a5a448, 32'h42540624};
test_weights[29632:29639] = '{32'h4161869a, 32'h4207d75d, 32'hc2af178d, 32'h4253cd64, 32'h41c1d334, 32'hc29f4b1b, 32'hc146402f, 32'hc209bdac};
test_bias[3704:3704] = '{32'hc1f42831};
test_output[3704:3704] = '{32'h457d9356};
test_input[29640:29647] = '{32'h42a5df77, 32'hc28e4b1c, 32'hc09ea38e, 32'hc2501007, 32'h41f681e0, 32'h428f9311, 32'h42b1ffa8, 32'h4259a1fc};
test_weights[29640:29647] = '{32'hc25a4cb3, 32'h41d983f1, 32'h42b01d40, 32'h410f4bb0, 32'hc2a85b9c, 32'h426414fb, 32'h42b59343, 32'hbf8f2d54};
test_bias[3705:3705] = '{32'hc28fb4d5};
test_output[3705:3705] = '{32'h45023c03};
test_input[29648:29655] = '{32'hc2401dd1, 32'hc2a4409d, 32'hc29a6ba0, 32'hc1729e59, 32'h4159c2af, 32'h41f2317d, 32'h41c69174, 32'h4207b201};
test_weights[29648:29655] = '{32'h42a5d309, 32'hc2620be3, 32'h4268c7f0, 32'h42c64a92, 32'h42582f83, 32'h4294d0e7, 32'h4282446e, 32'h416c162c};
test_bias[3706:3706] = '{32'h424381cd};
test_output[3706:3706] = '{32'hc337758b};
test_input[29656:29663] = '{32'hc24ac823, 32'hc23d1712, 32'hc22f47e3, 32'hc2c2129b, 32'h41ca1d00, 32'hc2c52e47, 32'hc0a3e09a, 32'h41840d56};
test_weights[29656:29663] = '{32'h429c0e7f, 32'hc27fe595, 32'h42541f87, 32'h4291529a, 32'hc031f68e, 32'h4224219d, 32'h422ee21e, 32'h41e02033};
test_bias[3707:3707] = '{32'h42b45f09};
test_output[3707:3707] = '{32'hc65c3424};
test_input[29664:29671] = '{32'hc0fe8273, 32'hc1ce5642, 32'h3fb76340, 32'h4267a871, 32'hc1a98fc6, 32'hc2777f51, 32'h42954293, 32'h42c10ad6};
test_weights[29664:29671] = '{32'hc2a3e347, 32'hc1b59c96, 32'h424ef803, 32'h420cc4d1, 32'hc21bf765, 32'hc16362e8, 32'hc1a39960, 32'h424fc26b};
test_bias[3708:3708] = '{32'hc23e7da0};
test_output[3708:3708] = '{32'h4604bb2b};
test_input[29672:29679] = '{32'hc1cea9d9, 32'hc26b7fd9, 32'h408a923d, 32'h3fc06830, 32'hc2745e50, 32'h4294f02f, 32'h423b2b60, 32'h4248515c};
test_weights[29672:29679] = '{32'hbf030cac, 32'h4169d3ef, 32'h40958db3, 32'h427f5a44, 32'hc1cd8da8, 32'h41780ada, 32'h419e21c0, 32'hc211fad0};
test_bias[3709:3709] = '{32'h41e1f3b6};
test_output[3709:3709] = '{32'h448bd6ab};
test_input[29680:29687] = '{32'hc2c5a03b, 32'hc2883cf3, 32'h422501d0, 32'hc288e6ac, 32'hc14f8d6e, 32'hc228bb6a, 32'hc27adfe1, 32'hc2822095};
test_weights[29680:29687] = '{32'hc1705bd5, 32'h42bd77bc, 32'h423406b7, 32'h4271bfbf, 32'hc0a4dfe0, 32'hc17633da, 32'hc1b4b712, 32'hc22c8118};
test_bias[3710:3710] = '{32'hc2b3edf8};
test_output[3710:3710] = '{32'hc516072b};
test_input[29688:29695] = '{32'h4214bedd, 32'hc18bdbe0, 32'hc2240244, 32'h42a4af9f, 32'h429ad7cd, 32'hc2bc36ed, 32'h4214e75b, 32'h4140c5f3};
test_weights[29688:29695] = '{32'hc251eade, 32'hc2412f19, 32'h41a5b40a, 32'hc27fbcc2, 32'h41b395d4, 32'h41bc7ca3, 32'h3fbe7f31, 32'h41a3f807};
test_bias[3711:3711] = '{32'h42151ade};
test_output[3711:3711] = '{32'hc5e60557};
test_input[29696:29703] = '{32'hc2a7a1b7, 32'hc29a470d, 32'h406f7a31, 32'hc2999480, 32'hc2826294, 32'h4286f002, 32'h423852e9, 32'h42ad5487};
test_weights[29696:29703] = '{32'hc2a2ebc9, 32'hc2a559a2, 32'hc1a9cf6f, 32'h42a29318, 32'h41f43e67, 32'hc18635d2, 32'hc244e0ae, 32'hc2a756da};
test_bias[3712:3712] = '{32'hc26a9994};
test_output[3712:3712] = '{32'hc5b5c458};
test_input[29704:29711] = '{32'hc289fcde, 32'hc28783ac, 32'hc28bb7bc, 32'h420db74c, 32'h42b32590, 32'h4251292c, 32'hc21f7400, 32'hc2a2f2ac};
test_weights[29704:29711] = '{32'h422963a7, 32'h427b3611, 32'h42333981, 32'h414fcdd3, 32'h42c49093, 32'hc1eda192, 32'h41eea454, 32'hc10aa281};
test_bias[3713:3713] = '{32'h4219ef9d};
test_output[3713:3713] = '{32'hc53e1737};
test_input[29712:29719] = '{32'hc21de864, 32'h416c58b8, 32'h4254db4c, 32'h427363ab, 32'h41d63ae0, 32'hc0f28288, 32'h424eadf4, 32'hc2c61566};
test_weights[29712:29719] = '{32'hc2950480, 32'hc28142ea, 32'h42b74a41, 32'hc28dfa84, 32'hc2b1f398, 32'hc116e57d, 32'h42395bf2, 32'h413669e5};
test_bias[3714:3714] = '{32'hc237b08d};
test_output[3714:3714] = '{32'h44b58297};
test_input[29720:29727] = '{32'h423412db, 32'hc2bd9424, 32'h42a6b4aa, 32'hc25340a5, 32'h426d2d4b, 32'h423d84c3, 32'hc22be71e, 32'h42c7d955};
test_weights[29720:29727] = '{32'hc1bd5bbd, 32'h429f3ca6, 32'hc2943e45, 32'hc10781c0, 32'h4241b2d2, 32'h423cf2e0, 32'hc2b32c30, 32'h4057d16c};
test_bias[3715:3715] = '{32'hc2a6f578};
test_output[3715:3715] = '{32'hc5a05500};
test_input[29728:29735] = '{32'h4146ccb9, 32'h42a6758c, 32'hc263ccc7, 32'hc2c49104, 32'hc238842c, 32'hc22c427b, 32'h42b9db2f, 32'h42be7212};
test_weights[29728:29735] = '{32'hc1ed0afa, 32'hc2981d89, 32'h41de5508, 32'h4196597c, 32'h42056670, 32'h41256e9a, 32'hc2596e9d, 32'h42819429};
test_bias[3716:3716] = '{32'hc1346e54};
test_output[3716:3716] = '{32'hc62bf49c};
test_input[29736:29743] = '{32'h42a5f111, 32'hc143f783, 32'hc23d8b33, 32'h421d9449, 32'hc2884572, 32'hc116260b, 32'h42aa895d, 32'hc2310005};
test_weights[29736:29743] = '{32'h4200f23e, 32'h42346493, 32'h42a8cdf0, 32'hc277e66a, 32'hc032c31d, 32'hc17bf9fb, 32'hc202dfd9, 32'h3f47ba3e};
test_bias[3717:3717] = '{32'hc23f852e};
test_output[3717:3717] = '{32'hc5d62661};
test_input[29744:29751] = '{32'hc0bf3115, 32'hc28ab197, 32'hc296b603, 32'hc2948309, 32'h41b98415, 32'hc26a6587, 32'hc2ad9127, 32'h422c9fd0};
test_weights[29744:29751] = '{32'h41b5fb91, 32'hc1f31882, 32'h42606d36, 32'h425879ff, 32'hc1cb499b, 32'h41efe0b9, 32'h42c23a9d, 32'hbf3884bf};
test_bias[3718:3718] = '{32'h42513639};
test_output[3718:3718] = '{32'hc68508bc};
test_input[29752:29759] = '{32'h41f3632a, 32'hc1e3a3ca, 32'h40d1b7d4, 32'h42ae0949, 32'hc16de415, 32'hc288e987, 32'h42b35d2c, 32'h4299e4b7};
test_weights[29752:29759] = '{32'h429c58f8, 32'hc2aea6cf, 32'hc23da9ca, 32'h423b5062, 32'h42a1d22f, 32'hc280d147, 32'h42b0c0f3, 32'hc297bc9c};
test_bias[3719:3719] = '{32'h41f66796};
test_output[3719:3719] = '{32'h465a0143};
test_input[29760:29767] = '{32'hbf79a5cb, 32'hc202dcfb, 32'h428801bc, 32'h424d8d73, 32'h41f18369, 32'h427aa721, 32'h42524ce2, 32'hc29053d5};
test_weights[29760:29767] = '{32'h404d3f59, 32'hc163544d, 32'hc2b01e23, 32'hbfd0512a, 32'hc1ab31b9, 32'hc217a5a0, 32'hc2262ff5, 32'hc245087e};
test_bias[3720:3720] = '{32'hc18d8f26};
test_output[3720:3720] = '{32'hc5e37a54};
test_input[29768:29775] = '{32'h42b2a7d4, 32'hc21f241f, 32'hbfc47d49, 32'hc0f2d72c, 32'hc2a81d13, 32'hc244208e, 32'h42bb18ca, 32'hc280a3d5};
test_weights[29768:29775] = '{32'h42a93bf7, 32'h41c637bb, 32'hc2ae19a9, 32'h41801483, 32'h42b42e8f, 32'h42be229f, 32'h42b3767a, 32'hc2ad39fe};
test_bias[3721:3721] = '{32'h41b78d3b};
test_output[3721:3721] = '{32'h46024c4a};
test_input[29776:29783] = '{32'h413da615, 32'hc1d122e0, 32'hc2764203, 32'h41990c44, 32'hc2804b46, 32'hc2acf254, 32'hbfb7b3b6, 32'hc27f5d5f};
test_weights[29776:29783] = '{32'hc2ac92dd, 32'h42b9fdbf, 32'h42ba50fc, 32'h426424f3, 32'h4107a5ac, 32'h418442ac, 32'h42a03b77, 32'h417cb738};
test_bias[3722:3722] = '{32'hc0fb4b1a};
test_output[3722:3722] = '{32'hc62f0a51};
test_input[29784:29791] = '{32'h41553dda, 32'h4246aa5d, 32'h42289cb4, 32'hc2b7e149, 32'h42b1a0fb, 32'hc20da7bc, 32'hc192ac1f, 32'h425fa692};
test_weights[29784:29791] = '{32'h412f64bc, 32'h41d125b1, 32'hc284aa59, 32'hc18e5b50, 32'hc21a24f7, 32'h4295161e, 32'h422fa850, 32'hc2798eec};
test_bias[3723:3723] = '{32'hc2994f98};
test_output[3723:3723] = '{32'hc61e9074};
test_input[29792:29799] = '{32'hc29624a4, 32'h42ad661b, 32'hc222103e, 32'h40b670cb, 32'hc2a38a5a, 32'h429e07ca, 32'h42874bd1, 32'hc14851f7};
test_weights[29792:29799] = '{32'h41d4d450, 32'hc2a6e167, 32'hc1d1900f, 32'h4202ac94, 32'h423913d8, 32'h429ae09e, 32'hc2991416, 32'hc2bfce80};
test_bias[3724:3724] = '{32'h423afef6};
test_output[3724:3724] = '{32'hc615aadb};
test_input[29800:29807] = '{32'hc2943169, 32'hc2020800, 32'hc23b05fe, 32'hc2a1d7db, 32'h424b6b65, 32'hc21cfd22, 32'hc2810a6c, 32'hc2be9f79};
test_weights[29800:29807] = '{32'hc2b9f506, 32'h423c2fa6, 32'hc2b8fd8d, 32'h42281303, 32'h42b9761f, 32'hc21c8b3a, 32'hc1ce3d99, 32'hc1ec29fe};
test_bias[3725:3725] = '{32'h4112a1fb};
test_output[3725:3725] = '{32'h4684fcd9};
test_input[29808:29815] = '{32'hbff02318, 32'hc1ae966b, 32'h4293a84a, 32'h42a3e715, 32'hc2338337, 32'h42a7b5df, 32'h41e23665, 32'hc2409fde};
test_weights[29808:29815] = '{32'h42a42955, 32'h427c2d8f, 32'hc16ca009, 32'h41ffd146, 32'h41ea9d1c, 32'h40f1ed51, 32'hc2c056c9, 32'h42903aa3};
test_bias[3726:3726] = '{32'hc28e9c5a};
test_output[3726:3726] = '{32'hc5d91586};
test_input[29816:29823] = '{32'h425cefe1, 32'hc285d4a8, 32'hbfeac73c, 32'h423acdc2, 32'h41020903, 32'hc21c776c, 32'h420956e0, 32'hc2a99505};
test_weights[29816:29823] = '{32'h428d0fd7, 32'h42b3de18, 32'hc2b71755, 32'hc2a60e64, 32'h425a475f, 32'h4104fa6d, 32'h4299db77, 32'hc2216687};
test_bias[3727:3727] = '{32'hc0dd8ced};
test_output[3727:3727] = '{32'h43ab2a5c};
test_input[29824:29831] = '{32'h42bd026b, 32'h4164540a, 32'hc2aae61f, 32'h42844aac, 32'h411b0154, 32'hc2592c3c, 32'hc20c6acf, 32'hc2b55681};
test_weights[29824:29831] = '{32'h4207fed4, 32'hc2c14c98, 32'hc2a8d315, 32'hc23a9d77, 32'h41e8f01b, 32'hc1d80a64, 32'h42bd7232, 32'h42192d7e};
test_bias[3728:3728] = '{32'h429799d6};
test_output[3728:3728] = '{32'h4476e75f};
test_input[29832:29839] = '{32'hc296e1cf, 32'h4280151f, 32'hc241255c, 32'h428a5a5e, 32'hc2c36a81, 32'hc29ae818, 32'h42bef860, 32'h41a2840f};
test_weights[29832:29839] = '{32'h428dfa91, 32'h4229ab97, 32'hc1c0115c, 32'h42a9ce8d, 32'h4262190a, 32'hc22decde, 32'hc26726f1, 32'h427f4c27};
test_bias[3729:3729] = '{32'hc2b3e536};
test_output[3729:3729] = '{32'hc5018d66};
test_input[29840:29847] = '{32'hc1365d57, 32'h426a582c, 32'hc265758f, 32'h424fe056, 32'hc2b41321, 32'hc2916e52, 32'hc2b55224, 32'h42c24e41};
test_weights[29840:29847] = '{32'h42abb3f7, 32'h41690c06, 32'hc291c0ed, 32'h42788cb6, 32'hc1a6cafe, 32'hc2c64b58, 32'hc0364348, 32'h42759190};
test_bias[3730:3730] = '{32'h422ca7a7};
test_output[3730:3730] = '{32'h46b0da37};
test_input[29848:29855] = '{32'hc19b0ed7, 32'h42183824, 32'hc1d5e89c, 32'h418265de, 32'h424d1cb0, 32'hc29f5853, 32'h426a74d4, 32'h40c8ac02};
test_weights[29848:29855] = '{32'hc1a48492, 32'h427cdf2c, 32'hc1e0ac70, 32'h42b094b2, 32'hbfd2197e, 32'h423576d5, 32'h4203c0a2, 32'h42b8b11d};
test_bias[3731:3731] = '{32'hc2aa0e08};
test_output[3731:3731] = '{32'h456887f6};
test_input[29856:29863] = '{32'hc152560b, 32'h41d6a777, 32'h413cddec, 32'h42b3896e, 32'hc090d470, 32'h41a790f6, 32'hc2ab1f17, 32'hc2bdb973};
test_weights[29856:29863] = '{32'h41526a70, 32'h410e9be1, 32'hc2b9a72c, 32'h42575181, 32'h4286996b, 32'hc2bc713b, 32'hc054c9b8, 32'hc0c92462};
test_bias[3732:3732] = '{32'hc29c3145};
test_output[3732:3732] = '{32'h451173fb};
test_input[29864:29871] = '{32'hc2b4b5ca, 32'hbd345096, 32'h42ba2263, 32'h42932d78, 32'hc292d104, 32'hc2c2c48a, 32'h42bc8568, 32'hc20197b1};
test_weights[29864:29871] = '{32'hc204fa66, 32'h42bf3ec5, 32'h423c7681, 32'h42a35fe1, 32'hc231237c, 32'h422fc78b, 32'hc29114b6, 32'h422c81f0};
test_bias[3733:3733] = '{32'h427cbe15};
test_output[3733:3733] = '{32'h45831b16};
test_input[29872:29879] = '{32'hc19902df, 32'h41b783e0, 32'hc16c2278, 32'h41fe5bee, 32'hc02161a6, 32'h40d84e34, 32'h42823396, 32'hc1f2fb45};
test_weights[29872:29879] = '{32'h4262cd4e, 32'hc2774a1e, 32'h425a253e, 32'h42c7caad, 32'h4218edeb, 32'hc29af226, 32'h40f376a7, 32'h40ad362e};
test_bias[3734:3734] = '{32'hc2609124};
test_output[3734:3734] = '{32'hc3ee5592};
test_input[29880:29887] = '{32'h405644c6, 32'hc14c2389, 32'h42a6f003, 32'h42bb1a45, 32'h429d583a, 32'h428e42e4, 32'hc247de1b, 32'hc2a9abfe};
test_weights[29880:29887] = '{32'h4176784c, 32'hc1b14c12, 32'hc2a8a6cf, 32'hc1cab0d2, 32'h4283a924, 32'h42c676af, 32'hc10f7fcd, 32'hc23abddd};
test_bias[3735:3735] = '{32'h42bf6d50};
test_output[3735:3735] = '{32'h45ef9b52};
test_input[29888:29895] = '{32'h42829193, 32'h428f4dc4, 32'hc1574780, 32'hc22dea4f, 32'h42069c2b, 32'h417399e3, 32'hc21b96fd, 32'hc2052d60};
test_weights[29888:29895] = '{32'h42c684ca, 32'h420a660d, 32'h401970d0, 32'h42a5b82c, 32'h420e6ba6, 32'hc2a067e7, 32'h429ef061, 32'h40c0feb3};
test_bias[3736:3736] = '{32'hc2bbd5b2};
test_output[3736:3736] = '{32'h44ef7134};
test_input[29896:29903] = '{32'h42bf04f6, 32'hc22d91f1, 32'hc1cd5042, 32'hc16eab1f, 32'h42c2df6c, 32'h41d43ae8, 32'h4289c103, 32'h41d8c505};
test_weights[29896:29903] = '{32'hc1920efd, 32'h426388d7, 32'hc29f6af5, 32'h42239493, 32'h42ac2230, 32'h428f0b3b, 32'h40de3625, 32'h4263e4bb};
test_bias[3737:3737] = '{32'h425e51eb};
test_output[3737:3737] = '{32'h4615c27a};
test_input[29904:29911] = '{32'hc0e10fac, 32'h41d63a70, 32'hc288b72a, 32'h4213bc7e, 32'h402094bb, 32'h42c2868b, 32'h42a27833, 32'h41f63910};
test_weights[29904:29911] = '{32'h42aafd2b, 32'h4208713c, 32'hc1f51bcf, 32'hc2b0df2f, 32'hc1c637b9, 32'h42927a38, 32'h4292dc97, 32'h4052faef};
test_bias[3738:3738] = '{32'h42b3a7ea};
test_output[3738:3738] = '{32'h46411785};
test_input[29912:29919] = '{32'h42a77ce4, 32'hc182cde1, 32'h421f9222, 32'hc2784b82, 32'h4275bb5c, 32'h42b38a7d, 32'h425113d4, 32'hc2930e6c};
test_weights[29912:29919] = '{32'h42b11fe7, 32'h41ac5899, 32'h42319a68, 32'hc2a30c7c, 32'hbfb3e932, 32'hc2149edb, 32'h42138802, 32'h42a63a15};
test_bias[3739:3739] = '{32'h420b9257};
test_output[3739:3739] = '{32'h45c5af03};
test_input[29920:29927] = '{32'h41e532be, 32'h41a06d75, 32'hc2900dc8, 32'hc23cc3a4, 32'h4209263b, 32'h42beefa1, 32'hc28b1e64, 32'h425882c0};
test_weights[29920:29927] = '{32'h410bb9f2, 32'hc28430d6, 32'h42bcdccf, 32'h41f417ee, 32'h4285ef8e, 32'h4235cc9f, 32'h40c16467, 32'hc2b4c1c6};
test_bias[3740:3740] = '{32'h41bf7f4e};
test_output[3740:3740] = '{32'hc5f90fde};
test_input[29928:29935] = '{32'hc255498a, 32'hc2b39ac6, 32'hc1eb0310, 32'hc189a669, 32'hc16f1048, 32'h41d87186, 32'hc2745b80, 32'h42216770};
test_weights[29928:29935] = '{32'h42b09bab, 32'hc2b90b5e, 32'hc23cbd49, 32'h419825c0, 32'hc19f07a5, 32'hc1274664, 32'h425509e1, 32'hc1b48693};
test_bias[3741:3741] = '{32'h42855a1b};
test_output[3741:3741] = '{32'h440ff04e};
test_input[29936:29943] = '{32'h4273e806, 32'h42ba5c76, 32'h42a39dc1, 32'h41cb07b5, 32'h40e12964, 32'h416f4703, 32'hc25d0628, 32'h421cf009};
test_weights[29936:29943] = '{32'hc2686167, 32'h4234d9af, 32'hc1b66527, 32'h429181a0, 32'h423b55ce, 32'h4273c80f, 32'h429a0441, 32'h4185a6bf};
test_bias[3742:3742] = '{32'hc1a43f0e};
test_output[3742:3742] = '{32'hc4d7f231};
test_input[29944:29951] = '{32'hc27c9714, 32'h4171c12d, 32'hc246daa2, 32'h423ac847, 32'hc0c35b8b, 32'hc1422dd9, 32'hc1ecb8e0, 32'h419e754f};
test_weights[29944:29951] = '{32'hc1f6052f, 32'h4279e08f, 32'h41f41fcf, 32'h42a735ce, 32'h4256f728, 32'h42860fe5, 32'h42422e2f, 32'h427d80c5};
test_bias[3743:3743] = '{32'hc1b9424a};
test_output[3743:3743] = '{32'h45756e20};
test_input[29952:29959] = '{32'hc1cf5202, 32'h42b53d7d, 32'hc0a70bf8, 32'hc263062d, 32'h42952fc1, 32'h4295b38a, 32'hc2ab3256, 32'h425548a2};
test_weights[29952:29959] = '{32'h42a85034, 32'hc1e3a1d6, 32'hc250039f, 32'hc02b6a99, 32'h42959de3, 32'hc2356ebe, 32'hc2a160d9, 32'h4268345e};
test_bias[3744:3744] = '{32'h3ea52650};
test_output[3744:3744] = '{32'h45f55d7f};
test_input[29960:29967] = '{32'h4286a75e, 32'h42401b12, 32'hc08e2f05, 32'h4292063f, 32'h41d91df1, 32'h401be46c, 32'hc2bf08fe, 32'hc1b809c2};
test_weights[29960:29967] = '{32'h4295aba9, 32'hc1bf09c6, 32'hc0a2f0fc, 32'hc2abc5ed, 32'hc1e92861, 32'hc2abb251, 32'hbdbfd1c6, 32'hc27c6e91};
test_bias[3745:3745] = '{32'h42041b57};
test_output[3745:3745] = '{32'hc4e8dd0a};
test_input[29968:29975] = '{32'h420cc978, 32'hc126b253, 32'h418bbba2, 32'hc28d55ba, 32'h429ef4ec, 32'h4238028a, 32'h42be9815, 32'h41d64d8b};
test_weights[29968:29975] = '{32'hc291af98, 32'hc28792be, 32'hc15eb849, 32'hc0fb5254, 32'hc2005f21, 32'hc25c85de, 32'h41bb5358, 32'hc246511e};
test_bias[3746:3746] = '{32'h429448e6};
test_output[3746:3746] = '{32'hc5b0b8cb};
test_input[29976:29983] = '{32'h42a7bf77, 32'h41bd9d68, 32'hc14693a6, 32'h42110b79, 32'h41d95b74, 32'h42900c24, 32'h42042870, 32'hc1fc5c18};
test_weights[29976:29983] = '{32'h425418c7, 32'hc2b51712, 32'h42898cec, 32'hc282e1db, 32'hc2ae3201, 32'h42395e00, 32'h42c51d03, 32'hc274e725};
test_bias[3747:3747] = '{32'h41e4f516};
test_output[3747:3747] = '{32'h45a4720d};
test_input[29984:29991] = '{32'hc1e28b58, 32'h41be7ab0, 32'h4124cd7c, 32'hc2b00762, 32'h42ae338e, 32'h4283dcf1, 32'hc27d941d, 32'hc27892c2};
test_weights[29984:29991] = '{32'h41da4d45, 32'hc2bf49c7, 32'hc20c1c70, 32'h420d2466, 32'hc204a89d, 32'hc02b4b9a, 32'hc1cfcc39, 32'hc240531e};
test_bias[3748:3748] = '{32'h42b054f6};
test_output[3748:3748] = '{32'hc597d696};
test_input[29992:29999] = '{32'hc2049c71, 32'hbf9d5634, 32'hc1d6c741, 32'hc29c1bde, 32'h419d005f, 32'hc08fcb74, 32'hc19b63cd, 32'h4284288b};
test_weights[29992:29999] = '{32'hc2b7bc61, 32'hc2a374c9, 32'h427ac1a0, 32'hc2734204, 32'h41d47c30, 32'h42a64180, 32'hc149e176, 32'h42a43287};
test_bias[3749:3749] = '{32'hc23d8267};
test_output[3749:3749] = '{32'h463b317f};
test_input[30000:30007] = '{32'hc28f9c75, 32'hc18b671e, 32'h42b75fac, 32'h42695ce9, 32'h4283433a, 32'hc276cdd8, 32'h42bfef4b, 32'hc2c536ad};
test_weights[30000:30007] = '{32'hc0ace299, 32'hc1a4763c, 32'h41c11a26, 32'h41786219, 32'h428e9e57, 32'hc0f8fd5c, 32'hc2b49c6f, 32'h4284b63e};
test_bias[3750:3750] = '{32'hc20c6c33};
test_output[3750:3750] = '{32'hc5c25bb9};
test_input[30008:30015] = '{32'h40bb54b6, 32'h4296ba90, 32'hc17b94cd, 32'h423156cf, 32'hc18cf93d, 32'hc21ed63c, 32'hc2c03ba1, 32'hc246ee71};
test_weights[30008:30015] = '{32'hc2c0e03b, 32'h4246f0c7, 32'h4266e06a, 32'hc1451da6, 32'h410fd2d9, 32'hc2adb67d, 32'hc1a008e9, 32'h413a8e53};
test_bias[3751:3751] = '{32'h4252993a};
test_output[3751:3751] = '{32'h45c88087};
test_input[30016:30023] = '{32'hc2bf4366, 32'hc295735f, 32'h4244a699, 32'hc179a02a, 32'h42a0373e, 32'h42b455d4, 32'h4292e57a, 32'h4206cd92};
test_weights[30016:30023] = '{32'hc13a3957, 32'hc2100eb8, 32'hc2c395fb, 32'h42bd6d4a, 32'hc1905e35, 32'hc22c8d95, 32'hc2a0dfdc, 32'h4202af02};
test_bias[3752:3752] = '{32'h420081df};
test_output[3752:3752] = '{32'hc644bd41};
test_input[30024:30031] = '{32'h426f777a, 32'h4249d79b, 32'h42b2e10f, 32'h42bb50bf, 32'hc26cea9b, 32'hc2bf1ceb, 32'hc2623a7c, 32'hc2a28968};
test_weights[30024:30031] = '{32'hc2b55acc, 32'h4150f642, 32'h41535c15, 32'hc088251a, 32'h42ac6548, 32'h42641690, 32'hc121c702, 32'hc10a9492};
test_bias[3753:3753] = '{32'h421c39cc};
test_output[3753:3753] = '{32'hc64ea7ce};
test_input[30032:30039] = '{32'h4211144b, 32'h41d8603a, 32'h42b030a2, 32'hc1f0edcc, 32'hc1f79900, 32'h42180b6b, 32'hc2c0fbeb, 32'hc20baaf8};
test_weights[30032:30039] = '{32'h422974f9, 32'h4206a81d, 32'h42afaab2, 32'hc2015cad, 32'h42bc4f32, 32'hc23ef7b1, 32'hc25e3964, 32'h40b9a704};
test_bias[3754:3754] = '{32'hc2b7a0ad};
test_output[3754:3754] = '{32'h4633a102};
test_input[30040:30047] = '{32'hc144a2d1, 32'h424db363, 32'h40fadd2c, 32'h422a1d9e, 32'hc1f0987e, 32'hc2a9c754, 32'hc264872f, 32'hc2931db3};
test_weights[30040:30047] = '{32'hc1d07fe0, 32'hc28c63b0, 32'hc098f59d, 32'hc2b3d900, 32'h41f469d8, 32'h41af0125, 32'h42c707fc, 32'h423cbd21};
test_bias[3755:3755] = '{32'hc19b1e2c};
test_output[3755:3755] = '{32'hc6953dbb};
test_input[30048:30055] = '{32'hc18657f5, 32'h42b30634, 32'hc1a56d55, 32'h415b8be5, 32'h41724138, 32'hc28acc61, 32'h4208fd11, 32'h419ca4a9};
test_weights[30048:30055] = '{32'h41b904ba, 32'h42adec87, 32'h420b094e, 32'h429406b6, 32'hc1f57774, 32'h4194a92d, 32'hc2a7d5b4, 32'hc29fb758};
test_bias[3756:3756] = '{32'hc1c275b9};
test_output[3756:3756] = '{32'h44b89065};
test_input[30056:30063] = '{32'hc28e07df, 32'hc1b0a10e, 32'hc2248a41, 32'hc2720e87, 32'h41a04b1b, 32'hc27b5955, 32'hc2af5aeb, 32'hc20ad457};
test_weights[30056:30063] = '{32'hc291acd4, 32'h41950aff, 32'h42abc077, 32'h414eee74, 32'hc0a93d4b, 32'h41d06531, 32'h42bcf42d, 32'h42357b76};
test_bias[3757:3757] = '{32'hc29d57b0};
test_output[3757:3757] = '{32'hc62f866f};
test_input[30064:30071] = '{32'hc1a4dd77, 32'h40d3de91, 32'h42c3a17f, 32'hc2132e33, 32'hc15ee5d5, 32'hc27a22d1, 32'h4270acd0, 32'h429f24ed};
test_weights[30064:30071] = '{32'h42468fd6, 32'h41a7c37d, 32'hc2b36c99, 32'h424b1d66, 32'hc2016b5f, 32'hc29096ee, 32'hc24aad26, 32'h42393cfa};
test_bias[3758:3758] = '{32'h42186eb6};
test_output[3758:3758] = '{32'hc5b7ce78};
test_input[30072:30079] = '{32'h42b6d619, 32'hc1a372c2, 32'hc253a999, 32'hc1010d88, 32'hc288ab6b, 32'hc28a1c5c, 32'h42c15f9c, 32'hc20fa13f};
test_weights[30072:30079] = '{32'hc20bd198, 32'hbffcec42, 32'hc255daf0, 32'h423819d2, 32'h41d53bd1, 32'hc213ac62, 32'h4207d6e4, 32'hc2941098};
test_bias[3759:3759] = '{32'hc23a7166};
test_output[3759:3759] = '{32'h45b92f23};
test_input[30080:30087] = '{32'h4107a870, 32'hc2a3a5fc, 32'h42a2fa90, 32'hc2638216, 32'hc14db7e4, 32'h42c17d75, 32'h42a2abdd, 32'hc276143a};
test_weights[30080:30087] = '{32'hc270d4c7, 32'hc20d4145, 32'h42bc6d4b, 32'hc2a0094f, 32'h4151ca75, 32'h42838b79, 32'h429039c6, 32'hc23cef2d};
test_bias[3760:3760] = '{32'hc28e4f3a};
test_output[3760:3760] = '{32'h46e67c62};
test_input[30088:30095] = '{32'h4292fe22, 32'hc231d8be, 32'hc1057f92, 32'h42b623c6, 32'h421d36c3, 32'h42074317, 32'hc0aa16b1, 32'h42b7e7d2};
test_weights[30088:30095] = '{32'hc2c45689, 32'hc0bba141, 32'hc2819c18, 32'hc23301c4, 32'h426a9859, 32'hc28a1f79, 32'hc0f5b6ea, 32'h42a54816};
test_bias[3761:3761] = '{32'h42a368b1};
test_output[3761:3761] = '{32'hc52eddf0};
test_input[30096:30103] = '{32'h428639fc, 32'h4293c969, 32'hc1bf6125, 32'h427adc22, 32'h42c774c6, 32'h418f18e5, 32'h42b74771, 32'hc1bd6594};
test_weights[30096:30103] = '{32'hc280d5aa, 32'h429a2f72, 32'h42413614, 32'hc1c2c4ae, 32'hc13a9ed2, 32'hc1bd27e2, 32'hc28f1e21, 32'h42be886e};
test_bias[3762:3762] = '{32'hc22d7c9c};
test_output[3762:3762] = '{32'hc6379e19};
test_input[30104:30111] = '{32'hc244f9e4, 32'hc2147462, 32'h4281e8c4, 32'hc2c3d2e8, 32'h40b1c636, 32'h41e04e50, 32'h41256430, 32'hc2b61d60};
test_weights[30104:30111] = '{32'hc24560a9, 32'h40d7f2b1, 32'h42abc0f4, 32'h423a509b, 32'hc2836277, 32'h420a5344, 32'hc28166d8, 32'h418347e3};
test_bias[3763:3763] = '{32'h42910357};
test_output[3763:3763] = '{32'h44d5e107};
test_input[30112:30119] = '{32'h413e3905, 32'hc05abe04, 32'h42872a6d, 32'hc15c7452, 32'hc27b4553, 32'h42b4a22a, 32'hc2bd8084, 32'h420ace32};
test_weights[30112:30119] = '{32'hc23aca4c, 32'h427c7a76, 32'hc0820426, 32'hc2c727fb, 32'h41b92f77, 32'h422e87ef, 32'hc1867e85, 32'h40d7a191};
test_bias[3764:3764] = '{32'hc2c62ada};
test_output[3764:3764] = '{32'h458de6d7};
test_input[30120:30127] = '{32'h41ad9d05, 32'h42c335c2, 32'hc1bccddc, 32'h4157c88b, 32'h42c42553, 32'h420bc5d2, 32'hc2556f2b, 32'hc296e305};
test_weights[30120:30127] = '{32'hc1fe8f60, 32'h42afd490, 32'h42926114, 32'h427a104d, 32'h42a9fb01, 32'h42ad4142, 32'h42b8e187, 32'h425f9579};
test_bias[3765:3765] = '{32'hc19137ac};
test_output[3765:3765] = '{32'h460fc37b};
test_input[30128:30135] = '{32'h42887732, 32'hc2b2d89e, 32'h428914ef, 32'hc2ad04c6, 32'h429b9350, 32'hc1e598eb, 32'hc28050c7, 32'h42ad154d};
test_weights[30128:30135] = '{32'hc269efad, 32'hc290afca, 32'hc1258aaa, 32'h42844e35, 32'h3f904f23, 32'hc2b83308, 32'h42bbbcd9, 32'hc02e9631};
test_bias[3766:3766] = '{32'hc25d000d};
test_output[3766:3766] = '{32'hc5eb8146};
test_input[30136:30143] = '{32'hc2711701, 32'hc1f930e5, 32'hc24b7910, 32'hc10c94ff, 32'h42b98af1, 32'h42a86b5f, 32'h425e070d, 32'h40a15cbc};
test_weights[30136:30143] = '{32'h407d90c9, 32'h40b57296, 32'hc22626eb, 32'hc20f0dff, 32'h40ff8849, 32'hc251d6cb, 32'hc22a4da5, 32'h40c28b92};
test_bias[3767:3767] = '{32'hc221d087};
test_output[3767:3767] = '{32'hc57c6134};
test_input[30144:30151] = '{32'h429ae05f, 32'hc254cd0b, 32'hc2835b61, 32'h429cc6dc, 32'hc1948aa1, 32'hc25dd384, 32'h42871540, 32'h40f24632};
test_weights[30144:30151] = '{32'hc27f2d57, 32'h41d795cc, 32'h42085d87, 32'hc1cda42b, 32'hc0a6b493, 32'hc2814379, 32'h428837ba, 32'h42b30bb0};
test_bias[3768:3768] = '{32'hc232eaf3};
test_output[3768:3768] = '{32'hc4d6334f};
test_input[30152:30159] = '{32'hc234f0f1, 32'h42896790, 32'hc26cb888, 32'hc1a1fdce, 32'h42a925bd, 32'hc18db7b8, 32'h4217e9fa, 32'h41ba3287};
test_weights[30152:30159] = '{32'hc1a144de, 32'h41fe9896, 32'hc219a484, 32'hc1c34f42, 32'h42663624, 32'h426d9de1, 32'hc29d1772, 32'h420d4125};
test_bias[3769:3769] = '{32'hc1c3c41b};
test_output[3769:3769] = '{32'h45ea3a96};
test_input[30160:30167] = '{32'hc23d9db2, 32'h424c5f2d, 32'h426aa39c, 32'h42033fa7, 32'h4230e7c6, 32'h421899be, 32'hc173b96c, 32'hc2bf60a5};
test_weights[30160:30167] = '{32'h4241197d, 32'h41910fa6, 32'h42ab88be, 32'hc2355a2d, 32'hc23870b1, 32'hc13b57f7, 32'h42b6f203, 32'h427ff41a};
test_bias[3770:3770] = '{32'h420d2e98};
test_output[3770:3770] = '{32'hc5f34c8c};
test_input[30168:30175] = '{32'h421adab8, 32'h42a9a5b3, 32'hc1fbb7e5, 32'h423ed8e9, 32'hc29a920f, 32'hc26af744, 32'h4283eef7, 32'hc10abe89};
test_weights[30168:30175] = '{32'h429900f5, 32'hbfe545b4, 32'hc2c40d68, 32'hc2a55b0f, 32'hc282ad4b, 32'h418e72f9, 32'h41ee4855, 32'h40605221};
test_bias[3771:3771] = '{32'hc2bd126e};
test_output[3771:3771] = '{32'h45f38855};
test_input[30176:30183] = '{32'hc1fbbf63, 32'hc2a7de20, 32'h40ea7284, 32'h419e6060, 32'hc0a44bcb, 32'h42440b7c, 32'hc1f6ec41, 32'h41268ece};
test_weights[30176:30183] = '{32'hc2a39c42, 32'h4212c0e0, 32'h429a20f1, 32'h42a6dd4f, 32'hc2c7d487, 32'h4264485d, 32'hc1c319fb, 32'h421d4880};
test_bias[3772:3772] = '{32'hc292cd99};
test_output[3772:3772] = '{32'h45beefb0};
test_input[30184:30191] = '{32'h428a8c00, 32'h41f2af18, 32'hc2b9a23a, 32'hc2265492, 32'hc29a490c, 32'hc2814de4, 32'hc29191ab, 32'h3e06ecfa};
test_weights[30184:30191] = '{32'h42a05a06, 32'h42b6c15d, 32'h41fa1e11, 32'h42a9c7b8, 32'hc20d66c4, 32'hc1967d94, 32'hc09ee731, 32'h4206159d};
test_bias[3773:3773] = '{32'h419a1864};
test_output[3773:3773] = '{32'h45c2742f};
test_input[30192:30199] = '{32'hc102dbf9, 32'h42ae9dce, 32'h4279d07c, 32'hc1705f5c, 32'hc1f710df, 32'h421ffebe, 32'hc29ca21c, 32'hc1be085c};
test_weights[30192:30199] = '{32'h427f66e2, 32'h42a4e319, 32'h424c15fe, 32'hc2709106, 32'hc297aceb, 32'h41330cdc, 32'h424279b0, 32'h42459b0b};
test_bias[3774:3774] = '{32'hc252a60b};
test_output[3774:3774] = '{32'h460526cd};
test_input[30200:30207] = '{32'h41d8744f, 32'hc2a4af85, 32'h415fbaca, 32'hc0e8425e, 32'hc1c08a97, 32'hc2bcc5c2, 32'h42b0be12, 32'h429d6e5e};
test_weights[30200:30207] = '{32'hc15ad655, 32'h42391dbf, 32'h42abfe35, 32'hc2c6a98f, 32'h4297514e, 32'h41508da9, 32'h40243fc5, 32'h42b8762c};
test_bias[3775:3775] = '{32'h423f110f};
test_output[3775:3775] = '{32'h450b1fcc};
test_input[30208:30215] = '{32'hc130eed3, 32'h429c111a, 32'h41e2eb4c, 32'hbdea4bec, 32'hc2663bb1, 32'hc26f0ed2, 32'h41ba5960, 32'h42bfab84};
test_weights[30208:30215] = '{32'h4250115e, 32'h42456615, 32'hc288edae, 32'h426aee30, 32'hc2b3e880, 32'h420cce85, 32'hbfc51051, 32'h411b7e49};
test_bias[3776:3776] = '{32'hc2aad281};
test_output[3776:3776] = '{32'h45a2d710};
test_input[30216:30223] = '{32'hc2399beb, 32'h4251a4bb, 32'hc2894a79, 32'h421ac15f, 32'h428b7ea6, 32'hc2685fee, 32'hc221bd05, 32'h413973ff};
test_weights[30216:30223] = '{32'h42923c0e, 32'hc1395412, 32'h41f592ca, 32'h42828f8c, 32'hc097b28f, 32'h4196247d, 32'h4022add0, 32'h421767d6};
test_bias[3777:3777] = '{32'hc24c13bf};
test_output[3777:3777] = '{32'hc5936b9e};
test_input[30224:30231] = '{32'hc296b9c2, 32'hc2b290d7, 32'h40c992f8, 32'hc2b7ca57, 32'h42bc1c07, 32'hc1ad1a47, 32'h428a065d, 32'hc15673e6};
test_weights[30224:30231] = '{32'h42b90a98, 32'h423c0839, 32'h42bcde95, 32'h41cf0be4, 32'hc2b9ecac, 32'h41f8950f, 32'h41b3cf5c, 32'h42c5f479};
test_bias[3778:3778] = '{32'hc29ad15b};
test_output[3778:3778] = '{32'hc6ad9bbe};
test_input[30232:30239] = '{32'h4238c8fc, 32'h41f7ae8c, 32'hc29fcdc4, 32'h42325f39, 32'h42c172e6, 32'h41dd0b76, 32'h4258fcc2, 32'hc2029dce};
test_weights[30232:30239] = '{32'hc1d178e0, 32'h413fe12d, 32'hc206fe68, 32'hc149e938, 32'hc27823e7, 32'hc124272d, 32'hc1ace539, 32'hc2b5f434};
test_bias[3779:3779] = '{32'h3f108a4b};
test_output[3779:3779] = '{32'hc5475506};
test_input[30240:30247] = '{32'hc291b156, 32'hbf9e2ca7, 32'hbdc95957, 32'hc28a8649, 32'hc281233d, 32'h42b703e3, 32'hc1bd573e, 32'hc296bb15};
test_weights[30240:30247] = '{32'h4201e7c8, 32'h423ed995, 32'h422b82af, 32'h421cfee7, 32'hc12a55b9, 32'h42384fda, 32'hc2019a75, 32'hc1e10da6};
test_bias[3780:3780] = '{32'h42adf01e};
test_output[3780:3780] = '{32'h452aa6c7};
test_input[30248:30255] = '{32'h41f53bb0, 32'h42c0c37c, 32'h428298d4, 32'hc23d8030, 32'h4298b465, 32'h40651b33, 32'h429980b0, 32'hc2208bae};
test_weights[30248:30255] = '{32'hc2bf7340, 32'h429f5c19, 32'hc2a87b73, 32'h4129847b, 32'h42549539, 32'h42b84c08, 32'h423cf914, 32'h42287222};
test_bias[3781:3781] = '{32'hc219753c};
test_output[3781:3781] = '{32'h459d1d41};
test_input[30256:30263] = '{32'h420b464f, 32'hc16ce55f, 32'h41d9ea08, 32'hc2b4ff20, 32'h4126d8d5, 32'hc2468c29, 32'h42972716, 32'h42a4ed20};
test_weights[30256:30263] = '{32'h42946631, 32'hc20f47e1, 32'h423bde14, 32'hc1d769ee, 32'hc22b2e22, 32'h428499a6, 32'h41be769e, 32'h420b23a1};
test_bias[3782:3782] = '{32'h420b2cb6};
test_output[3782:3782] = '{32'h45f39b6d};
test_input[30264:30271] = '{32'hc2a24898, 32'h4299cd2e, 32'hc2535d52, 32'h42813499, 32'h4092798d, 32'h42afc188, 32'h425ddf36, 32'hc2bd4291};
test_weights[30264:30271] = '{32'h41bd83d6, 32'hc2a00cc9, 32'h419f09ea, 32'h42893435, 32'h42156961, 32'hc291559c, 32'h4251da52, 32'hc23c8da1};
test_bias[3783:3783] = '{32'hc2674f0a};
test_output[3783:3783] = '{32'hc560cbfa};
test_input[30272:30279] = '{32'hc23a97a2, 32'hc2c5bf97, 32'hc0bebdf7, 32'h428985e2, 32'h4287fcc2, 32'h429aea7e, 32'hc15cd989, 32'h4026e95b};
test_weights[30272:30279] = '{32'h42b205cd, 32'h420b7f26, 32'h4203b60a, 32'hc285d95b, 32'h41d70073, 32'hc2b18b28, 32'hc2970986, 32'hc2c15f6a};
test_bias[3784:3784] = '{32'hc2c6c1a4};
test_output[3784:3784] = '{32'hc682e8b3};
test_input[30280:30287] = '{32'h4209f932, 32'h4256cd91, 32'hc262b375, 32'hc2ad5bcf, 32'hc241e10e, 32'hc29ae9ef, 32'h40ee2108, 32'hc0569a83};
test_weights[30280:30287] = '{32'h419611ba, 32'hc27f9285, 32'hc2a88d18, 32'h417f2c6a, 32'h4182180a, 32'h42b903ef, 32'h402fecd2, 32'hc1b438d2};
test_bias[3785:3785] = '{32'h42b11e9e};
test_output[3785:3785] = '{32'hc5dfb8ee};
test_input[30288:30295] = '{32'hc2989fe3, 32'h4245b4dc, 32'hc1a1226a, 32'h42a62473, 32'h42a8d776, 32'hc2a7cc33, 32'h42b8a20c, 32'hc2c5051e};
test_weights[30288:30295] = '{32'hc2a28114, 32'h42345e7d, 32'hc14392a2, 32'h40f0d483, 32'h4169954a, 32'hc25dc5c6, 32'hc1bb4f91, 32'h4218b8d3};
test_bias[3786:3786] = '{32'h42c6a1fb};
test_output[3786:3786] = '{32'h461245b0};
test_input[30296:30303] = '{32'h41065648, 32'hc2aab323, 32'hc2a37d1c, 32'h421317c5, 32'hc243c27f, 32'hc142513d, 32'h4222810c, 32'hc2692f0a};
test_weights[30296:30303] = '{32'h42a40943, 32'hc252cefd, 32'hc2b67d2d, 32'hc2aa2016, 32'hc1aa48d0, 32'h3fa6bde0, 32'h4115fbdb, 32'h3fbe4ced};
test_bias[3787:3787] = '{32'h41bd0e3f};
test_output[3787:3787] = '{32'h4629b481};
test_input[30304:30311] = '{32'hc12bcb0c, 32'h42a54750, 32'hc09c9532, 32'h4228fbc8, 32'h42aaa4c6, 32'hc2aab597, 32'hc27d89c7, 32'h410ed107};
test_weights[30304:30311] = '{32'hc0b4b346, 32'h41a3a83a, 32'h42c09a8c, 32'hc2a4951a, 32'hc28673e5, 32'hc27f669b, 32'h41996fa2, 32'hc2b731ae};
test_bias[3788:3788] = '{32'hc2927c32};
test_output[3788:3788] = '{32'hc58f67dd};
test_input[30312:30319] = '{32'h42043147, 32'hc2be2f69, 32'hc22510c2, 32'h42096b1c, 32'hc23aacdb, 32'hc1dafd62, 32'hbfa66646, 32'h4287a10e};
test_weights[30312:30319] = '{32'hc136c406, 32'hc091bb59, 32'h415087f7, 32'h42879722, 32'hc21a76e7, 32'hc016ff7a, 32'hc2ab9635, 32'hc1716212};
test_bias[3789:3789] = '{32'h4245ffd7};
test_output[3789:3789] = '{32'h45323815};
test_input[30320:30327] = '{32'h4231f8d4, 32'h42860e6e, 32'h4256cd16, 32'h40a11846, 32'h42992ae2, 32'hc24d5ef6, 32'h421ead4d, 32'hc18bd6be};
test_weights[30320:30327] = '{32'h424c084b, 32'h41fb92f6, 32'hc270d39f, 32'hc2a998d1, 32'h412944e1, 32'h422329fa, 32'h41c72355, 32'hc1114d8a};
test_bias[3790:3790] = '{32'hc29e2950};
test_output[3790:3790] = '{32'h43fa2852};
test_input[30328:30335] = '{32'h4224e3e6, 32'h42519f3a, 32'hc149b551, 32'hc20ac273, 32'hc0e0cdc1, 32'h4221bf56, 32'h420d58af, 32'h419a9c3a};
test_weights[30328:30335] = '{32'hc2807080, 32'h42a987ea, 32'hc1115cac, 32'h42ae9f5a, 32'hc1a56dbf, 32'h40c61f91, 32'hc2886e31, 32'h42924ad6};
test_bias[3791:3791] = '{32'hc2c0a3b4};
test_output[3791:3791] = '{32'hc4e31e71};
test_input[30336:30343] = '{32'h42839190, 32'h429f2f7e, 32'h42294b40, 32'hc24d3151, 32'hc161e446, 32'hc1b3151b, 32'hc1cf5821, 32'h4017eaac};
test_weights[30336:30343] = '{32'hc28fcc91, 32'hc2388aea, 32'h42847028, 32'hc1f87bed, 32'hc21b4c58, 32'h4258e84f, 32'h414123a6, 32'h419db82e};
test_bias[3792:3792] = '{32'h4155b1ac};
test_output[3792:3792] = '{32'hc599e356};
test_input[30344:30351] = '{32'h41603ff7, 32'hc2977a01, 32'h42a1a637, 32'hc27083d7, 32'h429430b0, 32'hc2539a3f, 32'h4286f785, 32'hc1f6bb8e};
test_weights[30344:30351] = '{32'hc1decd94, 32'hc29e5b3a, 32'hc22521c0, 32'h426d844a, 32'hc2c7c3b0, 32'h426e69ea, 32'h42655913, 32'hc233274d};
test_bias[3793:3793] = '{32'h40eed516};
test_output[3793:3793] = '{32'hc5ce22aa};
test_input[30352:30359] = '{32'hc1d84cae, 32'hc2010a17, 32'h424ceda9, 32'h42ab0af9, 32'h42ba1a49, 32'hc29fc727, 32'h40a00db7, 32'hc2380a5b};
test_weights[30352:30359] = '{32'h40e5b7d0, 32'hc2188131, 32'h42b07b0b, 32'h41aebba1, 32'h4264e9da, 32'hc2812f72, 32'hc067277d, 32'h4242081b};
test_bias[3794:3794] = '{32'hc218fac8};
test_output[3794:3794] = '{32'h46741711};
test_input[30360:30367] = '{32'hc2a3f6d9, 32'h41d9e3f5, 32'h420197c5, 32'h4202471d, 32'h40d9ee73, 32'h4287a8a4, 32'h423d7372, 32'h428a4194};
test_weights[30360:30367] = '{32'hc2bac266, 32'hc26dc4f6, 32'hc0a57b47, 32'hc12b9a71, 32'hc1ac7adb, 32'h4265a331, 32'hc28c1df0, 32'hc2329ea8};
test_bias[3795:3795] = '{32'hc2b8bc6a};
test_output[3795:3795] = '{32'h452d1641};
test_input[30368:30375] = '{32'hc24f283f, 32'hc283dee5, 32'h426eaeeb, 32'h42a79877, 32'h42c604f0, 32'h42a9549a, 32'h42a5276f, 32'hc2bc06c2};
test_weights[30368:30375] = '{32'h4284bfb1, 32'h4175691d, 32'h40008546, 32'hc244495e, 32'hc1cedaf7, 32'hc29b7fe9, 32'hc28b1818, 32'h419f75bd};
test_bias[3796:3796] = '{32'h4209f202};
test_output[3796:3796] = '{32'hc6c49c95};
test_input[30376:30383] = '{32'h41dc3069, 32'h4239cdff, 32'hc2bb32bb, 32'h42b168fe, 32'h3fec6b9d, 32'hc29f8629, 32'hc288008b, 32'h41c29b75};
test_weights[30376:30383] = '{32'hc244b776, 32'hc283c6a3, 32'hc26c6023, 32'h40a38508, 32'hc1e86869, 32'hc211b00e, 32'hc28d71c6, 32'hc29042be};
test_bias[3797:3797] = '{32'h3fbe82af};
test_output[3797:3797] = '{32'h45e9adc1};
test_input[30384:30391] = '{32'hc28d19f2, 32'hc1dd095e, 32'h423ee670, 32'h4285eced, 32'hc26f58d7, 32'h42459c4f, 32'h426110c3, 32'hc159b7e5};
test_weights[30384:30391] = '{32'hc28b2f78, 32'hc2be4d11, 32'h41daf987, 32'h4288c207, 32'hc12e0b7a, 32'h429c0d01, 32'h4267bac0, 32'hc2c1d71f};
test_bias[3798:3798] = '{32'h41bf308e};
test_output[3798:3798] = '{32'h46b007bf};
test_input[30392:30399] = '{32'hc246e8f9, 32'h42889aeb, 32'hc21b5cf6, 32'hc211ce1a, 32'hc2b74d6a, 32'hc246cbb3, 32'h428adfa0, 32'hc179109b};
test_weights[30392:30399] = '{32'h4212d756, 32'h42826281, 32'h427a3bfe, 32'h41f3b272, 32'h42131452, 32'hc17a48fa, 32'hc1f36087, 32'hc2156af8};
test_bias[3799:3799] = '{32'hc243ec03};
test_output[3799:3799] = '{32'hc59eeb2a};
test_input[30400:30407] = '{32'hc20099e3, 32'hc26fbf32, 32'hc1f1611e, 32'hc1f41c84, 32'hc1441cfa, 32'hc2bdeb47, 32'h42acbf80, 32'h4294b723};
test_weights[30400:30407] = '{32'h425870a1, 32'h42084edc, 32'hc2846b48, 32'hc2861732, 32'h422c876d, 32'hc20d5a2e, 32'h42492240, 32'hc1deed18};
test_bias[3800:3800] = '{32'hc2c13c1c};
test_output[3800:3800] = '{32'h45a4778f};
test_input[30408:30415] = '{32'h4284859e, 32'h4262b60f, 32'hc147a244, 32'hc212de14, 32'hc24910d0, 32'h42b676ca, 32'h420c8713, 32'hc22eb1ff};
test_weights[30408:30415] = '{32'h42608217, 32'h42c5275c, 32'hc1977f6e, 32'h3d8fced8, 32'hc2a1e4a9, 32'h41395b3b, 32'hc1819901, 32'h42503e49};
test_bias[3801:3801] = '{32'hc29f39a9};
test_output[3801:3801] = '{32'h46377ce0};
test_input[30416:30423] = '{32'hbfc6cc1d, 32'h3fccca13, 32'hc2a79e62, 32'h42b06ac2, 32'hc29fe915, 32'h42b75112, 32'hc1932e86, 32'hc1c38f4f};
test_weights[30416:30423] = '{32'h421ccd8c, 32'hc1eb3c2a, 32'hc294143e, 32'h41063365, 32'hc2abaae0, 32'h42b99479, 32'h427418cd, 32'h4219aa8d};
test_bias[3802:3802] = '{32'hc25e01f9};
test_output[3802:3802] = '{32'h469cef54};
test_input[30424:30431] = '{32'hc297eedb, 32'hc2bd4ca1, 32'h4263e5eb, 32'hc1d60b28, 32'hc040c172, 32'h4262df5d, 32'hc20d4092, 32'hc2a7ae81};
test_weights[30424:30431] = '{32'h424bad61, 32'h42c7ea36, 32'hc2730b0f, 32'h42c7548c, 32'h414bc9ba, 32'hc06f07fc, 32'h42a60a23, 32'hc2817f14};
test_bias[3803:3803] = '{32'h3e845b1d};
test_output[3803:3803] = '{32'hc6867529};
test_input[30432:30439] = '{32'hc224c8bc, 32'h42ad83c3, 32'h4172fa9b, 32'hc27bbab1, 32'hc2ae8f16, 32'hc150ac12, 32'h42c5f736, 32'h41a88054};
test_weights[30432:30439] = '{32'h422d1eeb, 32'hc23672fd, 32'h429e75ff, 32'hc098fa74, 32'hc2c6784a, 32'h41d917b2, 32'h420cebfa, 32'hc18483a8};
test_bias[3804:3804] = '{32'hc2c31ca2};
test_output[3804:3804] = '{32'h45de3f47};
test_input[30440:30447] = '{32'h42b3177c, 32'h42a81116, 32'hc26872d1, 32'hc1dbb0fe, 32'hc25ba13b, 32'hc2ad4113, 32'h40d40968, 32'hc1db6bab};
test_weights[30440:30447] = '{32'h42beb9a8, 32'hc28b4aa6, 32'hc20f0c8b, 32'h40f1b91a, 32'h4126ee8a, 32'h426321db, 32'hc1dea8ef, 32'h42641000};
test_bias[3805:3805] = '{32'h422960b3};
test_output[3805:3805] = '{32'hc525027a};
test_input[30448:30455] = '{32'h4298782d, 32'hc2342120, 32'h41a69893, 32'hc1c47bb5, 32'hc2bdf812, 32'hc216d4ff, 32'h42a86a84, 32'hc22334c5};
test_weights[30448:30455] = '{32'hc29853df, 32'hc20d0bf1, 32'hc2887f39, 32'h42c5ddeb, 32'h429be608, 32'h4230a612, 32'h408588ac, 32'hc1b6ceb4};
test_bias[3806:3806] = '{32'h429f3854};
test_output[3806:3806] = '{32'hc6767d87};
test_input[30456:30463] = '{32'hc2133a68, 32'hc1c61a7e, 32'h41807865, 32'h42a08175, 32'hc2c5bad8, 32'hc0860b68, 32'hc1a74e40, 32'h426333dc};
test_weights[30456:30463] = '{32'hc2942d47, 32'hc2b7a637, 32'hc2b51e58, 32'h42c4e62e, 32'h42c225d7, 32'hc286e2ac, 32'h427b1cc4, 32'h423d6372};
test_bias[3807:3807] = '{32'hc25831d0};
test_output[3807:3807] = '{32'h4557f1f1};
test_input[30464:30471] = '{32'hc2537099, 32'hc18c0f98, 32'h41fb948f, 32'hc1dca79f, 32'hc269d1a3, 32'hc0216245, 32'h4242e835, 32'h40326ad6};
test_weights[30464:30471] = '{32'h428ecf5a, 32'hc1c8ee91, 32'h4267d7c3, 32'hc23055c0, 32'h41c81429, 32'h3f384629, 32'h42c21312, 32'hc2817b9a};
test_bias[3808:3808] = '{32'hc28eb39f};
test_output[3808:3808] = '{32'h4529c9d9};
test_input[30472:30479] = '{32'h42a5c11d, 32'h41095bda, 32'h41fd8e38, 32'h42ac5efb, 32'h422acf87, 32'hc0807549, 32'hc01caae0, 32'hc28d609b};
test_weights[30472:30479] = '{32'hc2b672a4, 32'hc270fcab, 32'h424f4f30, 32'h4284aeae, 32'h41ceb0d3, 32'hbea6835f, 32'h42a700e1, 32'h42985c23};
test_bias[3809:3809] = '{32'h42a756fe};
test_output[3809:3809] = '{32'hc59ff429};
test_input[30480:30487] = '{32'h41b133d2, 32'h426c694c, 32'h4183d79e, 32'h428bf173, 32'hc2983ea7, 32'h40755002, 32'hc209fc14, 32'h42b4991f};
test_weights[30480:30487] = '{32'h42544e99, 32'hc206891c, 32'hc24ce2df, 32'hc18b321c, 32'h41862205, 32'hc2155f7b, 32'h413a8790, 32'h42669325};
test_bias[3810:3810] = '{32'hc22fb2f7};
test_output[3810:3810] = '{32'h43e8ea51};
test_input[30488:30495] = '{32'hc20e72d4, 32'h429d0273, 32'h41d0b76e, 32'hc118adcf, 32'h42a39ae8, 32'hc23e0997, 32'h4244fdfa, 32'h42afc2a7};
test_weights[30488:30495] = '{32'hc02da48c, 32'hc2c2a990, 32'h42bddf66, 32'h41ca09db, 32'h42ba8265, 32'h41bd8354, 32'h4244abf7, 32'hc2c310e6};
test_bias[3811:3811] = '{32'hc0d61f58};
test_output[3811:3811] = '{32'hc59b0fa6};
test_input[30496:30503] = '{32'hc282c58c, 32'h42adc5be, 32'h42be230a, 32'hc0ac9f2d, 32'hc26356bd, 32'hc1f4e8ce, 32'h40e5c933, 32'hc1f3c8d9};
test_weights[30496:30503] = '{32'hc2b8e96d, 32'hc290b9b9, 32'h4270e8ec, 32'hc2c76ed4, 32'h4289a76b, 32'hc1f6b425, 32'hc2705382, 32'h412b6f1e};
test_bias[3812:3812] = '{32'hc261c60f};
test_output[3812:3812] = '{32'h450bf8ae};
test_input[30504:30511] = '{32'hc1d1ed9f, 32'h42729a38, 32'h42c37383, 32'h42befeb8, 32'h426da4af, 32'hc2543674, 32'hc0609bc1, 32'h4103a719};
test_weights[30504:30511] = '{32'h42aeb69f, 32'h42a000e9, 32'hc20ce151, 32'h41a1bdbe, 32'hc235528e, 32'hc18d8a91, 32'h42954b1a, 32'h428966ea};
test_bias[3813:3813] = '{32'hc091159f};
test_output[3813:3813] = '{32'hc3cb83da};
test_input[30512:30519] = '{32'hc25fc81a, 32'hc2015ba2, 32'h422c06a3, 32'h42b2fe9c, 32'h428919a7, 32'h422451e3, 32'h42bdfcb8, 32'h41785547};
test_weights[30512:30519] = '{32'h4163066b, 32'h42adbadd, 32'hc296025e, 32'h425ec4ae, 32'hc2c479f9, 32'hc22a776c, 32'hc26f1010, 32'h4254920a};
test_bias[3814:3814] = '{32'hc0b47747};
test_output[3814:3814] = '{32'hc66d4df3};
test_input[30520:30527] = '{32'h420e306a, 32'h42935fda, 32'hc2be7da3, 32'hc2b5b774, 32'h425c4a9c, 32'h42b87c8e, 32'h428337ff, 32'hc19fb58a};
test_weights[30520:30527] = '{32'h4262bdf0, 32'hc1c11f1d, 32'hc2675ea7, 32'h3fc989ce, 32'h42b50970, 32'hc29fdfcd, 32'h427e4752, 32'hc25dc7d6};
test_bias[3815:3815] = '{32'hc29dd03d};
test_output[3815:3815] = '{32'h46037235};
test_input[30528:30535] = '{32'h420db7b6, 32'hc00bb273, 32'h423c95e3, 32'h428931fb, 32'hc19cd9d1, 32'h4196f6c0, 32'hc290d86e, 32'hc2c3cfd3};
test_weights[30528:30535] = '{32'hc134ce2b, 32'h4278327e, 32'h42c232c3, 32'hc2b9b728, 32'h41542811, 32'hc215b2dd, 32'hc2163730, 32'hc2bc8886};
test_bias[3816:3816] = '{32'hc27ed278};
test_output[3816:3816] = '{32'h46063d74};
test_input[30536:30543] = '{32'hc2918902, 32'h3f38080e, 32'h421c3ef9, 32'hc25360e9, 32'hc205ace1, 32'hc2b5486d, 32'hc28323d9, 32'h418b2ab8};
test_weights[30536:30543] = '{32'hc20ad81b, 32'h42aa79f6, 32'hc2208a75, 32'hc16744d5, 32'h41ea1820, 32'h42844954, 32'h41b8c420, 32'hc2ac0872};
test_bias[3817:3817] = '{32'h40b55d86};
test_output[3817:3817] = '{32'hc6000c3d};
test_input[30544:30551] = '{32'h4105fc7a, 32'h426e54ad, 32'hc0c466a2, 32'hc10bac06, 32'hc23737d2, 32'h426658e2, 32'h428abbc6, 32'hc2323c47};
test_weights[30544:30551] = '{32'hc15e8c7e, 32'h42b21f5a, 32'h424ea9de, 32'hc1302289, 32'hc2861e28, 32'hc2680351, 32'h42634939, 32'h42a8cf65};
test_bias[3818:3818] = '{32'h42845675};
test_output[3818:3818] = '{32'h459a98d5};
test_input[30552:30559] = '{32'hc1be82e2, 32'h41f695ef, 32'hc2422f2c, 32'h41c9e5e8, 32'h428c4e37, 32'h425fc7b5, 32'h4143afa0, 32'h4272ab52};
test_weights[30552:30559] = '{32'hc29aadb4, 32'h4270f764, 32'hc286512e, 32'h41b82494, 32'h424cc435, 32'hc28769c2, 32'h42893a97, 32'h42c030fe};
test_bias[3819:3819] = '{32'hc27baf62};
test_output[3819:3819] = '{32'h4659f52d};
test_input[30560:30567] = '{32'hc20b2008, 32'h41a545c7, 32'hc2060da9, 32'h41dfe7a6, 32'hc2a2d1b6, 32'hc22cce9f, 32'hc1e7bf1b, 32'h412f293d};
test_weights[30560:30567] = '{32'hc2939136, 32'hc1b004aa, 32'h42a05c87, 32'h41a20540, 32'h42123eaf, 32'h425fc61c, 32'hc249badc, 32'hc2511384};
test_bias[3820:3820] = '{32'hc23b30f0};
test_output[3820:3820] = '{32'hc58e7f51};
test_input[30568:30575] = '{32'hc201e9d7, 32'hc189535d, 32'h42266ef3, 32'h42c59254, 32'h42868666, 32'hc26fee92, 32'hc289c29e, 32'h42679441};
test_weights[30568:30575] = '{32'h4274aa16, 32'h422105a6, 32'hc28a1552, 32'h41272691, 32'h4191848d, 32'hc203f4d2, 32'hc27e2ff8, 32'h42091adb};
test_bias[3821:3821] = '{32'hc213df6e};
test_output[3821:3821] = '{32'h459c844f};
test_input[30576:30583] = '{32'h42c3b52e, 32'hc18f7814, 32'hc2883647, 32'h42c5e2a3, 32'hc26e6d0e, 32'h42638d66, 32'hc24cb8c1, 32'h42428c51};
test_weights[30576:30583] = '{32'hc1204571, 32'hc0b13392, 32'h42a901cf, 32'h42927068, 32'h42a4b404, 32'h422f0472, 32'h426a6e90, 32'h42918823};
test_bias[3822:3822] = '{32'h41bfa418};
test_output[3822:3822] = '{32'hc49bf4d1};
test_input[30584:30591] = '{32'hc1d60ae1, 32'h41328137, 32'hc2b48eb2, 32'h4297020c, 32'h420b2301, 32'h41d3fad2, 32'hc206470b, 32'hc1900d53};
test_weights[30584:30591] = '{32'h426db904, 32'hc1dd8b57, 32'hc2bc1e81, 32'h427c80c4, 32'h425be396, 32'hc2b535b7, 32'hc26774a6, 32'hc2c25f97};
test_bias[3823:3823] = '{32'hc286089a};
test_output[3823:3823] = '{32'h46627e4b};
test_input[30592:30599] = '{32'hc2b94d03, 32'h4285d073, 32'hc24c5993, 32'h4207d389, 32'hc29fba13, 32'hc2907f9f, 32'h42c31e57, 32'h425dbb7f};
test_weights[30592:30599] = '{32'hc2adee0f, 32'hc2982a7d, 32'h4259b473, 32'h41c019f2, 32'h42c0b9f5, 32'h4285a451, 32'hc2550e46, 32'hc29c8c86};
test_bias[3824:3824] = '{32'hc2b5920b};
test_output[3824:3824] = '{32'hc6a53830};
test_input[30600:30607] = '{32'hc07c0a6b, 32'h4199552b, 32'hc23d9cf5, 32'h41c5d44d, 32'hc2996d59, 32'h42acd337, 32'h414342dd, 32'h428785f7};
test_weights[30600:30607] = '{32'hc2907527, 32'hc137c5f9, 32'hc1d1d339, 32'h428ffccd, 32'hc180eb90, 32'h4189e301, 32'hc1f7c4f9, 32'hc2671ef9};
test_bias[3825:3825] = '{32'hc118a02a};
test_output[3825:3825] = '{32'h44bcd823};
test_input[30608:30615] = '{32'hc1724396, 32'hc260571c, 32'hc0dfaef3, 32'h42c1ef9e, 32'hc13c9ddb, 32'hc1d351e6, 32'hc25673f6, 32'hc2780935};
test_weights[30608:30615] = '{32'hc284a558, 32'h4266e704, 32'hc26fae43, 32'hc28a4a42, 32'hc283fc08, 32'hc21960fd, 32'hc18d8bcd, 32'h427d5d14};
test_bias[3826:3826] = '{32'h4231d250};
test_output[3826:3826] = '{32'hc616fc9b};
test_input[30616:30623] = '{32'h42c3dd7c, 32'h41ff4ef4, 32'h42477ab4, 32'hc2634e49, 32'hc294b2c2, 32'h41281f53, 32'h429c9038, 32'h42c05721};
test_weights[30616:30623] = '{32'hc12d0234, 32'h42b3fe70, 32'hc1cc5c49, 32'hc20fb716, 32'hc29dab74, 32'hc1727586, 32'h4298c138, 32'hc1d95852};
test_bias[3827:3827] = '{32'h4262b44d};
test_output[3827:3827] = '{32'h4636e78d};
test_input[30624:30631] = '{32'hc10ba5ee, 32'h42be2e83, 32'hc2336dea, 32'h42bd6a81, 32'hc20ca202, 32'h42a97d60, 32'hc205ea02, 32'h4278522f};
test_weights[30624:30631] = '{32'hc27bf825, 32'hc1c3e498, 32'hc29662d4, 32'hc24e1499, 32'h41fd0c47, 32'hc2a3036b, 32'h41cf38c3, 32'h4159812a};
test_bias[3828:3828] = '{32'h4245767c};
test_output[3828:3828] = '{32'hc630394c};
test_input[30632:30639] = '{32'h4280054a, 32'h426cc15b, 32'h41dee4d7, 32'hc2278baa, 32'hc1f37ca5, 32'h41a64577, 32'h424cc1da, 32'hc2c4dd79};
test_weights[30632:30639] = '{32'hc22695e6, 32'h4261b7f4, 32'hc1a60c1a, 32'hc28985e9, 32'hc08678e0, 32'h41964959, 32'hc19fbf0a, 32'h42285214};
test_bias[3829:3829] = '{32'hc2696955};
test_output[3829:3829] = '{32'hc4d804bf};
test_input[30640:30647] = '{32'h42849412, 32'hc15ef035, 32'h41bee143, 32'h427696df, 32'hc299484c, 32'h41f0b02a, 32'hc1f36427, 32'h429339cc};
test_weights[30640:30647] = '{32'hc1ebe16b, 32'h42275bed, 32'h3fb912c9, 32'hc216679d, 32'h41973c99, 32'hc27f7ea8, 32'h428fb484, 32'h416517af};
test_bias[3830:3830] = '{32'h3ff78e4a};
test_output[3830:3830] = '{32'hc611a6d0};
test_input[30648:30655] = '{32'hc29767f3, 32'h41f3aaea, 32'h40e635c6, 32'h425de6e7, 32'h427dc36c, 32'hc285e1b2, 32'h423ca96a, 32'hc2af380c};
test_weights[30648:30655] = '{32'h424c4f8d, 32'h413d0fa7, 32'hc22cf573, 32'h425a7cd6, 32'h403b96f2, 32'hc1519201, 32'hc234a0f4, 32'h4218bbd2};
test_bias[3831:3831] = '{32'h42604a9b};
test_output[3831:3831] = '{32'hc5a0bfdf};
test_input[30656:30663] = '{32'h429dedd6, 32'h4243672f, 32'hc283a660, 32'h42ba404d, 32'hc05bd39b, 32'hc215f853, 32'h42b731b2, 32'hc19d08c6};
test_weights[30656:30663] = '{32'hc2acfad9, 32'h42ba0622, 32'hc236d426, 32'h4255d39d, 32'h40f27434, 32'hc1ab7756, 32'hc29a9048, 32'h42ab8d75};
test_bias[3832:3832] = '{32'hbecd4412};
test_output[3832:3832] = '{32'hc50ec6d3};
test_input[30664:30671] = '{32'h42c1919d, 32'h42a30fd5, 32'hc2bd0682, 32'h4285ecd1, 32'h42b890ac, 32'h41a2f87b, 32'h4286ac89, 32'hc1399b6d};
test_weights[30664:30671] = '{32'hc2b9a06a, 32'hc27afe54, 32'hc187daa8, 32'h4078b8d8, 32'h41d40ce8, 32'hc2a4501d, 32'h41dea52c, 32'hc1eba18a};
test_bias[3833:3833] = '{32'h4185b0ef};
test_output[3833:3833] = '{32'hc61032ec};
test_input[30672:30679] = '{32'hc024dd05, 32'hc2909bea, 32'h42163a94, 32'h415416e4, 32'h420c6803, 32'h42c5b12e, 32'hc1774083, 32'hc299af26};
test_weights[30672:30679] = '{32'h42c67326, 32'h42431ce9, 32'h4200f2eb, 32'hc286cd28, 32'hc1c94770, 32'h4196f798, 32'hc292c090, 32'h425347e2};
test_bias[3834:3834] = '{32'h416e8192};
test_output[3834:3834] = '{32'hc5a88840};
test_input[30680:30687] = '{32'hc20886b8, 32'h420fd8d1, 32'hc202315b, 32'h4177fcb6, 32'hc186e8ee, 32'hc2933c17, 32'h428a46a5, 32'h42a5f626};
test_weights[30680:30687] = '{32'hc222a146, 32'h42238b7e, 32'hc2a54cdd, 32'hc2a690a9, 32'h42afaadd, 32'h42c4bf39, 32'h42bf4fc4, 32'hc26377e4};
test_bias[3835:3835] = '{32'h4295d4e8};
test_output[3835:3835] = '{32'hc51c05de};
test_input[30688:30695] = '{32'hc2c6660a, 32'hc18c211e, 32'h4226e4bc, 32'h4082af7c, 32'h42861945, 32'hc22a77ac, 32'h424f1030, 32'h4201eba4};
test_weights[30688:30695] = '{32'h421cb0d6, 32'h42555a0e, 32'hc16d2bb2, 32'hc0e72721, 32'h4210431d, 32'hc107dde1, 32'h40f2e4e3, 32'hc2bdcacf};
test_bias[3836:3836] = '{32'h41d5e670};
test_output[3836:3836] = '{32'hc5a73557};
test_input[30696:30703] = '{32'h422fef4a, 32'hc262f61e, 32'hc289f413, 32'hc2617885, 32'h4268be83, 32'hc29bd07c, 32'hc04a8edb, 32'hc13c669b};
test_weights[30696:30703] = '{32'h4049efb5, 32'h42b6a1b5, 32'h411fe5a6, 32'h4204480f, 32'h4291f522, 32'hc234705d, 32'hc280577c, 32'h419fa937};
test_bias[3837:3837] = '{32'h42bde50c};
test_output[3837:3837] = '{32'h4363d3a7};
test_input[30704:30711] = '{32'hc1a106db, 32'hc28ebe1f, 32'h4289d21e, 32'h4111cee1, 32'hbeca13fe, 32'hc2029ff6, 32'h4232e59c, 32'h42630644};
test_weights[30704:30711] = '{32'h42267f50, 32'hc2a39183, 32'hc2a6d8b4, 32'h420ca30e, 32'hc2a849de, 32'h429294f1, 32'h428b1c74, 32'h41efde00};
test_bias[3838:3838] = '{32'h42958962};
test_output[3838:3838] = '{32'h45032089};
test_input[30712:30719] = '{32'h426b093b, 32'h4196e711, 32'hc24fa3a3, 32'hc0b97c3e, 32'hc210b026, 32'hc186b665, 32'h421f654b, 32'hc2977953};
test_weights[30712:30719] = '{32'hc24cc06d, 32'h4286edff, 32'h42ac18a6, 32'h4286f9d0, 32'hc207b529, 32'h42c68be7, 32'hc28f157a, 32'h40dd3107};
test_bias[3839:3839] = '{32'h41031f54};
test_output[3839:3839] = '{32'hc6228f03};
test_input[30720:30727] = '{32'hc2bb10c5, 32'hc2a31feb, 32'hc2331571, 32'hc275e02d, 32'hc188def1, 32'h3ffea558, 32'hc29ecb07, 32'hc220d630};
test_weights[30720:30727] = '{32'hc2964cda, 32'hbf5c6df1, 32'hc2b660bf, 32'h4148c291, 32'h42106b7f, 32'h428706e9, 32'h4199759f, 32'h4252e043};
test_bias[3840:3840] = '{32'h4292cfc0};
test_output[3840:3840] = '{32'h45c6ae0d};
test_input[30728:30735] = '{32'hc1021a5e, 32'hc1bf6174, 32'hc2833d02, 32'h416ab44e, 32'h42ab7d25, 32'h41a4c98c, 32'h428a222d, 32'hc2b1a832};
test_weights[30728:30735] = '{32'hc25767cb, 32'hc2bf8017, 32'h422e2317, 32'hc281fba0, 32'hc0eb5f23, 32'hc21f9259, 32'h423711ba, 32'h42c2c99f};
test_bias[3841:3841] = '{32'h42bdaae6};
test_output[3841:3841] = '{32'hc5f7cbe5};
test_input[30736:30743] = '{32'hc277b3dc, 32'h423e3983, 32'hc2945531, 32'h42bbb3ac, 32'hc1e9b3e7, 32'hc21d8361, 32'h419474bc, 32'hc252192b};
test_weights[30736:30743] = '{32'hc230d36d, 32'hc260fd79, 32'h414827ed, 32'h42bcde83, 32'hc2569e38, 32'hc13c5e2f, 32'h42608157, 32'h42389ea0};
test_bias[3842:3842] = '{32'h3fd76545};
test_output[3842:3842] = '{32'h46071e16};
test_input[30744:30751] = '{32'h41268b93, 32'hc21f6f51, 32'h41059575, 32'h42ade440, 32'h42b06765, 32'h42a9cfd9, 32'hc2989ef4, 32'h42adbee9};
test_weights[30744:30751] = '{32'h4217d3cc, 32'hc2b257fb, 32'hc1e09b6b, 32'h420fbb5c, 32'h423e29fc, 32'h42b23044, 32'hc1ad3bb2, 32'hc13b0b9b};
test_bias[3843:3843] = '{32'hc0c1e1a5};
test_output[3843:3843] = '{32'h469637ab};
test_input[30752:30759] = '{32'h427f559b, 32'h42a408db, 32'hc13a4833, 32'h41b0760b, 32'h426fd965, 32'h4217f408, 32'h40c8f659, 32'hc269ed04};
test_weights[30752:30759] = '{32'hc109781d, 32'h4240389f, 32'hc28bfcd3, 32'h424490b3, 32'hc25e328b, 32'hc2af5959, 32'hc27d96f6, 32'h4143dcc3};
test_bias[3844:3844] = '{32'h42907276};
test_output[3844:3844] = '{32'hc516b839};
test_input[30760:30767] = '{32'hc28a2a9e, 32'h4282ef1b, 32'h421c6866, 32'h423c585c, 32'h42c28eb6, 32'h427a7c94, 32'hc26ab552, 32'hc2c618f4};
test_weights[30760:30767] = '{32'h41e0ff36, 32'hc26f4211, 32'h42af2fdb, 32'hc1d829e5, 32'h42994a59, 32'h42a22c9a, 32'hc29a0c5a, 32'hc2b02643};
test_bias[3845:3845] = '{32'hc2b74bb7};
test_output[3845:3845] = '{32'h46abb6a3};
test_input[30768:30775] = '{32'hc2099e9b, 32'h429d25c5, 32'h429e2314, 32'hc0eb1a42, 32'h4176aba1, 32'h429ecea1, 32'hc2c6ef5e, 32'hc2c202f5};
test_weights[30768:30775] = '{32'h41e6451a, 32'h417bb552, 32'h40dd2777, 32'hc036233b, 32'hc2944a1f, 32'h4253c38d, 32'h3fe48f8f, 32'h418e0203};
test_bias[3846:3846] = '{32'hc25afb72};
test_output[3846:3846] = '{32'h44efef26};
test_input[30776:30783] = '{32'h424afe1b, 32'hc2abeb6e, 32'h40c07b78, 32'hc21e8207, 32'hc2995536, 32'h41bbada7, 32'h42879cf7, 32'hc26eaec9};
test_weights[30776:30783] = '{32'hc14f4303, 32'h4161dfd9, 32'hc1d77430, 32'hc2a60e41, 32'hc22fe340, 32'hc26716d2, 32'h429cb815, 32'hc27f7d32};
test_bias[3847:3847] = '{32'hc2a6490a};
test_output[3847:3847] = '{32'h46406a32};
test_input[30784:30791] = '{32'h4282a7ff, 32'h41aadb50, 32'hc28cd0a7, 32'hc1ea110c, 32'h4299ffc8, 32'h424a5b6e, 32'h4297db93, 32'hc0a7b8fc};
test_weights[30784:30791] = '{32'h422ab94a, 32'hc263d2c3, 32'hc212aea6, 32'hc2bf48ba, 32'hc2278959, 32'h40aa6e5a, 32'h41fd38ea, 32'h4251ce63};
test_bias[3848:3848] = '{32'hc2c26edd};
test_output[3848:3848] = '{32'h45bc5d5b};
test_input[30792:30799] = '{32'h421acae1, 32'hc182db83, 32'hc14e0932, 32'hc1e0d0e9, 32'h42178444, 32'hc20cb6fd, 32'h41836197, 32'h427c5bbb};
test_weights[30792:30799] = '{32'h428712c9, 32'h42b629a8, 32'h42921512, 32'h4249b91d, 32'hc1047745, 32'hc2b607e1, 32'h429d628b, 32'h41e47570};
test_bias[3849:3849] = '{32'h42b3f0ca};
test_output[3849:3849] = '{32'h459730e3};
test_input[30800:30807] = '{32'h424a27b6, 32'hc07767da, 32'hc2bbbe9e, 32'h41a8e8d1, 32'hc265e90d, 32'hc2903add, 32'hc2405a4a, 32'hc2a228cd};
test_weights[30800:30807] = '{32'h3f264cd6, 32'h418875a3, 32'hc2416cea, 32'h40a5df68, 32'hc246cf2e, 32'h4144118a, 32'h41e2fb52, 32'h428f5780};
test_bias[3850:3850] = '{32'h428f798f};
test_output[3850:3850] = '{32'hc400bfeb};
test_input[30808:30815] = '{32'hc22afe3c, 32'h42624762, 32'h423ab677, 32'hc25cb08e, 32'hc28ec88d, 32'h4256b50d, 32'hc1bf8d3e, 32'hc26d078f};
test_weights[30808:30815] = '{32'h42852ee8, 32'hc2be3eee, 32'hc22e18cd, 32'h41a54d66, 32'hc2af0153, 32'h41c94c7d, 32'h4279db58, 32'hc1897b5d};
test_bias[3851:3851] = '{32'h42b2ff67};
test_output[3851:3851] = '{32'hc582ecc8};
test_input[30816:30823] = '{32'hc0e535ec, 32'h3f0bd4df, 32'hc29ebd84, 32'hc226d70c, 32'h417ce099, 32'hc24e4215, 32'h4059691e, 32'h3eb70b82};
test_weights[30816:30823] = '{32'hc1e8bb93, 32'h429549d2, 32'hc1bbb9b6, 32'h42b94458, 32'h42801cef, 32'h42969d92, 32'hc29d1a1f, 32'hc28795af};
test_bias[3852:3852] = '{32'h423678af};
test_output[3852:3852] = '{32'hc5982315};
test_input[30824:30831] = '{32'hc2ac8ad1, 32'hc2bce222, 32'h3fdd7ede, 32'hc1175569, 32'h4138f9ef, 32'hc2c21f38, 32'hc2baa7e0, 32'hc25840c8};
test_weights[30824:30831] = '{32'h42bd1a44, 32'hc2a48be0, 32'h425415e0, 32'h42b43161, 32'h424f2205, 32'hc123b64f, 32'h428cc731, 32'hbf6dcbcd};
test_bias[3853:3853] = '{32'h4238f348};
test_output[3853:3853] = '{32'hc5bc639d};
test_input[30832:30839] = '{32'hc1eafe05, 32'h4295259f, 32'hc1d0d4ea, 32'hc15fe1f7, 32'hc15d6bd1, 32'hc25f5ae4, 32'hc1a96b0c, 32'h426d59e8};
test_weights[30832:30839] = '{32'hc2a1a1cd, 32'h41caadc4, 32'hc2910369, 32'h42371b8d, 32'h4173887a, 32'hc18b66c1, 32'hc2a89cca, 32'h427d5bb7};
test_bias[3854:3854] = '{32'h429fed1d};
test_output[3854:3854] = '{32'h4639f601};
test_input[30840:30847] = '{32'h428a24cf, 32'h42736bf8, 32'hc0114446, 32'hc1826b78, 32'h41f92edf, 32'hc107895c, 32'h42ac9b36, 32'h41beac43};
test_weights[30840:30847] = '{32'hc2a152a0, 32'h42bccb7d, 32'hc25563c8, 32'hc29fe40b, 32'h42737932, 32'hbf25db7d, 32'hc1d1e2c1, 32'h41df6400};
test_bias[3855:3855] = '{32'h4230c8b6};
test_output[3855:3855] = '{32'h44f30f4f};
test_input[30848:30855] = '{32'hc1f08fff, 32'h41926b3e, 32'h41dc9e61, 32'hc2337408, 32'h40a8702e, 32'hc1ccbf33, 32'hc1b12f6a, 32'h409bd8d3};
test_weights[30848:30855] = '{32'hc286b644, 32'hc26f66c9, 32'h42a90556, 32'hc23ecc19, 32'hc0441b60, 32'h41bb6bfb, 32'hc25fec29, 32'h40af10f0};
test_bias[3856:3856] = '{32'h422ae55f};
test_output[3856:3856] = '{32'h45be705e};
test_input[30856:30863] = '{32'h41f875da, 32'h422756e1, 32'h42984637, 32'h428d0820, 32'h4284e922, 32'hc25bf884, 32'h414d6ac5, 32'h42c2dec7};
test_weights[30856:30863] = '{32'hc28c8731, 32'h419939c0, 32'h42928b8f, 32'hc18d7040, 32'h41a7a6f4, 32'hc204dab0, 32'h416d19c7, 32'hc105108b};
test_bias[3857:3857] = '{32'h429575ff};
test_output[3857:3857] = '{32'h45afc77a};
test_input[30864:30871] = '{32'h4193205c, 32'hc17fb9b1, 32'h425e42c2, 32'hc1ce23dc, 32'hc28d3539, 32'hc26454c7, 32'hc1a6c422, 32'h41bcb96d};
test_weights[30864:30871] = '{32'hc242f662, 32'hc139542a, 32'h42ab84be, 32'hc286ddb9, 32'hc1f398e7, 32'hbfb45002, 32'h427a1685, 32'h4247a10e};
test_bias[3858:3858] = '{32'hc28a8b83};
test_output[3858:3858] = '{32'h45f494b7};
test_input[30872:30879] = '{32'hc2816439, 32'h40ef7b4e, 32'h412c8bf6, 32'h4182aa40, 32'h4298680a, 32'hc2a1053d, 32'hc2c441c1, 32'h427d4770};
test_weights[30872:30879] = '{32'h40b4228c, 32'h4021190b, 32'hc29b9a5d, 32'hc1909e43, 32'hc13fc50c, 32'hc233501a, 32'h422171f7, 32'hc2648c92};
test_bias[3859:3859] = '{32'hc1d458e8};
test_output[3859:3859] = '{32'hc5c7a729};
test_input[30880:30887] = '{32'hc2b8d6ae, 32'hc19cb034, 32'hc2173799, 32'hc2bca350, 32'h40608333, 32'hc2c01513, 32'h42061568, 32'hc1de5b1f};
test_weights[30880:30887] = '{32'h42a61d84, 32'h426cd2c6, 32'h4289b5b9, 32'h42867f42, 32'hc13f879f, 32'h4289fe98, 32'h428221b1, 32'hc28971e3};
test_bias[3860:3860] = '{32'hc29c4ff4};
test_output[3860:3860] = '{32'hc69faa3d};
test_input[30888:30895] = '{32'h41a2f8af, 32'h42aab83e, 32'h42069965, 32'hc2c177e0, 32'hc2488c42, 32'h41560b87, 32'h4299c40c, 32'hc05c3dc1};
test_weights[30888:30895] = '{32'hc278da2d, 32'hc091e8b2, 32'h42679833, 32'hc20a4af3, 32'h42436da0, 32'hc16d5889, 32'hc21a7911, 32'hc22b0fa3};
test_bias[3861:3861] = '{32'h4212f961};
test_output[3861:3861] = '{32'hc4e0a1e4};
test_input[30896:30903] = '{32'hc1421501, 32'hc2c5277d, 32'h42119324, 32'hc276b357, 32'hc1077aed, 32'hc2816900, 32'h4281aa36, 32'h420baad2};
test_weights[30896:30903] = '{32'hc1f9bbc8, 32'hbf6cc3b5, 32'h4230e826, 32'hc2be92c7, 32'hc24359a0, 32'hc2c4efd6, 32'hc292a884, 32'hc282b448};
test_bias[3862:3862] = '{32'hc204b413};
test_output[3862:3862] = '{32'h45efbff5};
test_input[30904:30911] = '{32'hc1a68a0b, 32'h415f00d3, 32'hbfcda5d7, 32'hc1ca057e, 32'hc29c07b1, 32'hc2a0b18e, 32'h426795f0, 32'h4161d0f3};
test_weights[30904:30911] = '{32'h4102e9d3, 32'hc059116f, 32'h41e0146f, 32'h425d9901, 32'h41a2e75a, 32'hc2b6548b, 32'hc087a10a, 32'hc283d9b9};
test_bias[3863:3863] = '{32'hc225fe43};
test_output[3863:3863] = '{32'h453294bf};
test_input[30912:30919] = '{32'hc2455866, 32'hc2bced9e, 32'h41a0ce5f, 32'h42c0f452, 32'h42a72027, 32'h420d53ce, 32'hc1ba3701, 32'h42ae2097};
test_weights[30912:30919] = '{32'hc26115f0, 32'hc20c4cae, 32'h427b5e5d, 32'h3fe16614, 32'h416c8ab1, 32'hc2b3bcb3, 32'hc022a6c5, 32'h42ada4c7};
test_bias[3864:3864] = '{32'hc276cc7d};
test_output[3864:3864] = '{32'h464d4cff};
test_input[30920:30927] = '{32'h42827f51, 32'hc29e99a3, 32'hc2b2f88c, 32'h42c5dded, 32'hc29f7b4a, 32'hc20a7551, 32'hc25ec806, 32'h42af28ce};
test_weights[30920:30927] = '{32'hc2872ce4, 32'hc1b1d0e5, 32'hbfc9a07e, 32'hc1d63f08, 32'hc1bd1800, 32'h429839ae, 32'hc206d963, 32'h42b71bcb};
test_bias[3865:3865] = '{32'hc0d52ece};
test_output[3865:3865] = '{32'h4578f7f2};
test_input[30928:30935] = '{32'h4291fcb2, 32'h415c293e, 32'h426282c3, 32'hc299317b, 32'hc047b77e, 32'h41fce0b3, 32'h41eb3318, 32'hc2b858ac};
test_weights[30928:30935] = '{32'hc18d7be0, 32'hc2b621c7, 32'h41bcdf57, 32'hc25f1fda, 32'h42c723ab, 32'hc28e309a, 32'hc14361a9, 32'hc291e993};
test_bias[3866:3866] = '{32'hc12d4377};
test_output[3866:3866] = '{32'h45d672a3};
test_input[30936:30943] = '{32'hc2b6f434, 32'h42691fb2, 32'hc2b7a81e, 32'hc0f7f413, 32'h42aa2440, 32'hc2a14992, 32'hc28173cf, 32'h4265cc2c};
test_weights[30936:30943] = '{32'hc1307a80, 32'h41042619, 32'hc1df5bde, 32'hc2af9303, 32'hc1bd1f0c, 32'hc21f263a, 32'hc1bd1053, 32'hc1b39cb7};
test_bias[3867:3867] = '{32'h4230ef5a};
test_output[3867:3867] = '{32'h45c23fe9};
test_input[30944:30951] = '{32'hc26ba645, 32'h425387ae, 32'h4196a1d9, 32'hc1355c23, 32'hc2a26f4e, 32'hc2a3aeef, 32'hc28b77e1, 32'h3fbfab84};
test_weights[30944:30951] = '{32'h420327ba, 32'hc28a69bd, 32'h4292b5bb, 32'h42b2e1f1, 32'h401c2b6d, 32'hc28ad432, 32'hc22e464c, 32'hc2086506};
test_bias[3868:3868] = '{32'h42923d67};
test_output[3868:3868] = '{32'h454f6ffd};
test_input[30952:30959] = '{32'h4136816f, 32'hc2c4044d, 32'h402ccb06, 32'hc253bf71, 32'h42924b8f, 32'h42adcd24, 32'hc0a45e11, 32'h41242492};
test_weights[30952:30959] = '{32'hc24a6de8, 32'h414d304f, 32'hc1868e4a, 32'hc111d318, 32'h429f827c, 32'hc2af5686, 32'hc2961c1b, 32'hc268f0d3};
test_bias[3869:3869] = '{32'hc2b8ef96};
test_output[3869:3869] = '{32'hc559e163};
test_input[30960:30967] = '{32'h41a44304, 32'hc218f5ca, 32'h41ef39c5, 32'h3f78e87e, 32'h428bab52, 32'hc284dc97, 32'hc29e5551, 32'hc298ef2d};
test_weights[30960:30967] = '{32'h423130cd, 32'hc248fd58, 32'h428852c3, 32'h411073de, 32'hc1604a8e, 32'h42b0280f, 32'h429952a4, 32'h4225a4f7};
test_bias[3870:3870] = '{32'hc2365006};
test_output[3870:3870] = '{32'hc62f84dc};
test_input[30968:30975] = '{32'hc224571e, 32'hc2af0262, 32'hc1775bd1, 32'hc2b831c0, 32'hc1fc1acd, 32'h4233f097, 32'hc2a7c4bc, 32'h4248a155};
test_weights[30968:30975] = '{32'h416e240b, 32'h4236f849, 32'h42287a60, 32'hc2bfec2d, 32'hc2b57989, 32'hc251d48a, 32'h42adaa95, 32'h42c03664};
test_bias[3871:3871] = '{32'h4199d9f7};
test_output[3871:3871] = '{32'h44cb7902};
test_input[30976:30983] = '{32'hc278e8fa, 32'h41a47ba5, 32'h4297068c, 32'h41b2f21b, 32'h42121b2a, 32'hc2668ed5, 32'hc1f3913e, 32'h4267cb37};
test_weights[30976:30983] = '{32'hc2370fa1, 32'hc25c21d6, 32'h42ad5910, 32'hc1bb7c09, 32'hc05304a3, 32'hc2a7ac92, 32'h417e7bf7, 32'h423e6389};
test_bias[3872:3872] = '{32'hc1bdfd46};
test_output[3872:3872] = '{32'h4665acdb};
test_input[30984:30991] = '{32'h42c65b9b, 32'h4284c945, 32'hc1adf270, 32'h4255bead, 32'hc1ca5fd5, 32'h42c1bdb6, 32'h422f17cc, 32'hc29dc051};
test_weights[30984:30991] = '{32'hbf99614c, 32'h41a866aa, 32'h4237db53, 32'h428cca64, 32'h4276c559, 32'hc213e393, 32'hc2b65d57, 32'hc2ad1717};
test_bias[3873:3873] = '{32'h4208716a};
test_output[3873:3873] = '{32'h44dcfca8};
test_input[30992:30999] = '{32'h42963ee1, 32'h4146d949, 32'hc1dd2589, 32'h412148bb, 32'h428c3c90, 32'h4186e8f2, 32'h4208af36, 32'h42a86f19};
test_weights[30992:30999] = '{32'h41753e46, 32'h4214b3ee, 32'hc2a5474f, 32'hc2b67de6, 32'h428b8bae, 32'hc2c3b2e4, 32'hc1b6418e, 32'h42581c12};
test_bias[3874:3874] = '{32'hc2b44ef9};
test_output[3874:3874] = '{32'h461ab703};
test_input[31000:31007] = '{32'hc1d1a447, 32'h4127e977, 32'hc1ea6d18, 32'h4113daaa, 32'hc28a803c, 32'h42c68cd0, 32'h41021d30, 32'hc27b7f35};
test_weights[31000:31007] = '{32'hc2a90e9e, 32'hc29e7f91, 32'h4230169b, 32'h41ec5496, 32'h40dede23, 32'h423f81f1, 32'hc203f786, 32'hc20a2bf6};
test_bias[3875:3875] = '{32'hc103fe28};
test_output[3875:3875] = '{32'h45cc2335};
test_input[31008:31015] = '{32'hc1512d9a, 32'h3f5ae8bb, 32'h4271a4f0, 32'h429fd1c8, 32'h424d6f73, 32'h42b77c65, 32'hc25f06d9, 32'h42c43db8};
test_weights[31008:31015] = '{32'hc2c6d81b, 32'hc2329e17, 32'h42add7d2, 32'hc2650780, 32'hc28a693f, 32'hc2546173, 32'hc2a60704, 32'h42249a7a};
test_bias[3876:3876] = '{32'h40477328};
test_output[3876:3876] = '{32'h450853be};
test_input[31016:31023] = '{32'hc2b25232, 32'hc2c11a2c, 32'h42a83d89, 32'hc2810977, 32'hc2b0a74d, 32'hc2b916d4, 32'hc281e82e, 32'h428e66c4};
test_weights[31016:31023] = '{32'h4227ab69, 32'hc0fec470, 32'h429528bf, 32'hc2062501, 32'h4272e3bc, 32'h3f592cff, 32'hc2c52649, 32'h4265991d};
test_bias[3877:3877] = '{32'h41d75334};
test_output[3877:3877] = '{32'h4624bd44};
test_input[31024:31031] = '{32'h41aea1bf, 32'hc0b36017, 32'h42ac5cb4, 32'hc2390979, 32'hc24f0aa0, 32'h429c9751, 32'hc2940f26, 32'h4191971f};
test_weights[31024:31031] = '{32'h428c7b04, 32'hc20e1c2e, 32'h42b16387, 32'h40e09893, 32'h42532674, 32'hc2982c4e, 32'hc0fb8dbd, 32'hc219f210};
test_bias[3878:3878] = '{32'hc17ba94a};
test_output[3878:3878] = '{32'h4363cc3e};
test_input[31032:31039] = '{32'h42b0c698, 32'hc2a0398c, 32'h423776c1, 32'hc1a7b96c, 32'h4286de32, 32'h42a4726e, 32'hc2a46c97, 32'h42b35e2d};
test_weights[31032:31039] = '{32'h429525b8, 32'hc1b0e703, 32'h42883f54, 32'h421d1132, 32'hc266d771, 32'h42a1797f, 32'hc2c1fce4, 32'h429f37f9};
test_bias[3879:3879] = '{32'hc1704a07};
test_output[3879:3879] = '{32'h46debba4};
test_input[31040:31047] = '{32'h42828b09, 32'h41f1ef11, 32'h40dccd95, 32'h41b0e865, 32'hc247441a, 32'hbf558fea, 32'hc157d16f, 32'h42a4898d};
test_weights[31040:31047] = '{32'hc21648c2, 32'h426e1799, 32'h42691c69, 32'h42ad229f, 32'hc2b546e7, 32'h429ee01e, 32'hc1da2e24, 32'h42281fbe};
test_bias[3880:3880] = '{32'h41bf0a9f};
test_output[3880:3880] = '{32'h461bab31};
test_input[31048:31055] = '{32'hc27d74f4, 32'hc28ff1cd, 32'h428104b8, 32'hc2c56eec, 32'h41ae59fc, 32'h4298226b, 32'h420399dd, 32'h424a928e};
test_weights[31048:31055] = '{32'h412952e7, 32'hc22252b6, 32'hc29b3cbd, 32'hc080a3f9, 32'hc25b87b6, 32'hc2c133c4, 32'h41be17c3, 32'h41c749b5};
test_bias[3881:3881] = '{32'h40de59d6};
test_output[3881:3881] = '{32'hc60a589d};
test_input[31056:31063] = '{32'h40c66191, 32'hc21f58dd, 32'hc150efa6, 32'h4230fc75, 32'h41ad5266, 32'hc2c6c0ed, 32'hc2a171ea, 32'h415edaa2};
test_weights[31056:31063] = '{32'h42a4bae1, 32'hc1e2b469, 32'h42258b0b, 32'h41d01978, 32'hc2c02bb9, 32'h4244d360, 32'hc2aed817, 32'h41351621};
test_bias[3882:3882] = '{32'h41817323};
test_output[3882:3882] = '{32'h451cd17e};
test_input[31064:31071] = '{32'hc295a3c2, 32'hc27c4869, 32'hc18e46ab, 32'h429e8034, 32'h42a26d1d, 32'h42932bfb, 32'h41fbf856, 32'h4297f1b1};
test_weights[31064:31071] = '{32'h42384636, 32'hc28d38f3, 32'h4236bfe9, 32'hc2ac32dc, 32'hc24c9ec4, 32'hc1b1d8ca, 32'hc206b517, 32'hc28dac36};
test_bias[3883:3883] = '{32'hc2149921};
test_output[3883:3883] = '{32'hc693a615};
test_input[31072:31079] = '{32'h4085b2f4, 32'h42c6cf3b, 32'hc2045c44, 32'hc1f4a147, 32'hc2745ea4, 32'hc23a3404, 32'h40e79def, 32'hc2061786};
test_weights[31072:31079] = '{32'hc29bf972, 32'h42968aa4, 32'hc2292a51, 32'h41bd7d62, 32'hc283ba94, 32'hc1b8f99e, 32'h4154f627, 32'h41c6faa0};
test_bias[3884:3884] = '{32'h4229552c};
test_output[3884:3884] = '{32'h463f3266};
test_input[31080:31087] = '{32'h42c6e298, 32'hc289f573, 32'h4290fd0c, 32'hc28a3ad5, 32'h42014df5, 32'h42c25493, 32'h42159c9f, 32'h42ac5e12};
test_weights[31080:31087] = '{32'hc2687c4d, 32'h41fcacce, 32'h42b78ad5, 32'hc1ed8449, 32'h415c56cf, 32'hc1d88dea, 32'hc28cf700, 32'h4280f732};
test_bias[3885:3885] = '{32'h413c8c27};
test_output[3885:3885] = '{32'h44bacaea};
test_input[31088:31095] = '{32'hc1364db5, 32'hc26cc1eb, 32'hc18e2911, 32'hc25a2388, 32'hc221adb7, 32'hc2429420, 32'h42748efe, 32'hc202e2e1};
test_weights[31088:31095] = '{32'hc284c380, 32'h424565ca, 32'h4296bd26, 32'h4193e620, 32'h42084e0b, 32'hc294514b, 32'h42bd0db6, 32'hc18c8794};
test_bias[3886:3886] = '{32'hc2b019a9};
test_output[3886:3886] = '{32'h4579006f};
test_input[31096:31103] = '{32'h413fd0d9, 32'hc2a4684d, 32'h414875ca, 32'h41ddd596, 32'h4263c513, 32'h3ff97046, 32'hc1e8f0ef, 32'h42a01f56};
test_weights[31096:31103] = '{32'hc22a85d8, 32'hc168253b, 32'h4237498c, 32'hc1b3f302, 32'hc217a143, 32'h4184242c, 32'h418818dc, 32'h423b2b47};
test_bias[3887:3887] = '{32'hc28bee10};
test_output[3887:3887] = '{32'h44d2d19e};
test_input[31104:31111] = '{32'hc1b6ec13, 32'hc27c7072, 32'h4118ed16, 32'h42bde1be, 32'hc2b39328, 32'hc0fffde8, 32'h426b12e2, 32'hc2b83a30};
test_weights[31104:31111] = '{32'hc256e491, 32'h415c4fb6, 32'hc15506a3, 32'h42123daf, 32'h4211b5d7, 32'h426edc78, 32'h41208106, 32'h42bea832};
test_bias[3888:3888] = '{32'hc1262bf3};
test_output[3888:3888] = '{32'hc600dc8c};
test_input[31112:31119] = '{32'hc1ca458c, 32'hc2527b74, 32'hc1fb1ea3, 32'h42b4aa37, 32'hc070c21a, 32'h4235e9fc, 32'hc28a5a99, 32'h41aeaa37};
test_weights[31112:31119] = '{32'hc1eb4f96, 32'hc27a4d3d, 32'hc2bc0410, 32'hc2078363, 32'hc11075c3, 32'h41b36b2d, 32'hc2940b69, 32'h42654d91};
test_bias[3889:3889] = '{32'hc13607d9};
test_output[3889:3889] = '{32'h46313755};
test_input[31120:31127] = '{32'hc2bc19ee, 32'h42c10158, 32'h4280bf15, 32'h410890b8, 32'hc1fac0e2, 32'h4188c992, 32'h422d982c, 32'h42373766};
test_weights[31120:31127] = '{32'hc28f96b5, 32'hc224ea17, 32'h41f09c63, 32'hc2a44e72, 32'h4256a43e, 32'hc2136e4e, 32'hc29057b5, 32'h4224ad6b};
test_bias[3890:3890] = '{32'h41ac1a45};
test_output[3890:3890] = '{32'h43ebbf9b};
test_input[31128:31135] = '{32'h4281b6d7, 32'hc11ef885, 32'h429b6912, 32'h4251ce39, 32'h4152a421, 32'hc09774d8, 32'h41a938d7, 32'hc19a1894};
test_weights[31128:31135] = '{32'hc28caea6, 32'h42a8ada3, 32'h42afb6ef, 32'h3f90e296, 32'h3d5e75ec, 32'h4248c7b6, 32'hc2c02d5a, 32'hc2a3e1f1};
test_bias[3891:3891] = '{32'hc0a740f2};
test_output[3891:3891] = '{32'h44457ede};
test_input[31136:31143] = '{32'h421b604a, 32'hc22fcb55, 32'hc28eb37e, 32'h42477ee1, 32'h41ea04fa, 32'h4246aed9, 32'h42a94698, 32'hc26120d1};
test_weights[31136:31143] = '{32'h419e6336, 32'hc29e8dbc, 32'h41fdd3f9, 32'h42992193, 32'hc1e6d19b, 32'h4204dc17, 32'hc193f6b4, 32'hc2857f0e};
test_bias[3892:3892] = '{32'hc06bc80b};
test_output[3892:3892] = '{32'h46098574};
test_input[31144:31151] = '{32'hc20df2f3, 32'h416d988d, 32'hc29797f9, 32'h4253c3aa, 32'h42b81986, 32'h40c7036a, 32'h40980d9f, 32'hc06d6534};
test_weights[31144:31151] = '{32'h429ee771, 32'h425aabc9, 32'h42a826b8, 32'hbf8a5a40, 32'hc26a69d0, 32'h42a4c081, 32'hc2a28a73, 32'hc2a49d69};
test_bias[3893:3893] = '{32'h4226be07};
test_output[3893:3893] = '{32'hc650bbad};
test_input[31152:31159] = '{32'h425e916b, 32'hbf09b29b, 32'hc2b37aa5, 32'h40c23c08, 32'hc151de06, 32'h428ca2a6, 32'h41e32d86, 32'hc2900f8c};
test_weights[31152:31159] = '{32'h4222c1b0, 32'hc26643bb, 32'h41e5a419, 32'hc22edb36, 32'h4219ba76, 32'h424a9bfc, 32'h41bec0a6, 32'h42039ece};
test_bias[3894:3894] = '{32'hc2186962};
test_output[3894:3894] = '{32'h44430a0f};
test_input[31160:31167] = '{32'hc2a07ba5, 32'h4196063b, 32'hc2c4b4ed, 32'h42befe01, 32'hc2bd3c66, 32'hc2952caa, 32'hc28e5a83, 32'hc16a9095};
test_weights[31160:31167] = '{32'h4281a4c6, 32'hc2a039fc, 32'hc2527488, 32'hc0600b9a, 32'hc2c58ef9, 32'h420a0bbe, 32'h42c16b06, 32'hc20f1461};
test_bias[3895:3895] = '{32'h426f76a1};
test_output[3895:3895] = '{32'hc4adca61};
test_input[31168:31175] = '{32'hc2127774, 32'h42b4e113, 32'hc29040fc, 32'hc268e15d, 32'h418148c3, 32'hc2b66f9c, 32'h428aa8f2, 32'h3f90e132};
test_weights[31168:31175] = '{32'hc1bedbb6, 32'h420c105e, 32'hc292b057, 32'h41e1cc1d, 32'hc2b668d1, 32'hc1a464ea, 32'hc1f7cf67, 32'hc2941782};
test_bias[3896:3896] = '{32'hc1044061};
test_output[3896:3896] = '{32'h45b6c140};
test_input[31176:31183] = '{32'hc24c8f59, 32'hc2a239e3, 32'hc1ca0433, 32'h4194099e, 32'h419368bd, 32'h42aceb85, 32'hc22c4bd8, 32'h4126898f};
test_weights[31176:31183] = '{32'hc238b6f8, 32'hc1244653, 32'hc2bcfac4, 32'hc1f8b586, 32'h42a6ea70, 32'hc271a932, 32'hc2570a47, 32'h4266b0cd};
test_bias[3897:3897] = '{32'hc2385594};
test_output[3897:3897] = '{32'h4582eaa5};
test_input[31184:31191] = '{32'hc2c4c6e9, 32'h42586199, 32'h41ae3b23, 32'h426def1a, 32'h4267133a, 32'h428b3001, 32'hc2118df9, 32'h40df8194};
test_weights[31184:31191] = '{32'h42b1a7b4, 32'h40bc64cf, 32'hc227f94f, 32'h41e196c6, 32'hc2a2c29c, 32'hc2b7eb0c, 32'h41842394, 32'h41df9abb};
test_bias[3898:3898] = '{32'hc232e10f};
test_output[3898:3898] = '{32'hc69613cd};
test_input[31192:31199] = '{32'hc14b2f78, 32'h429d9b42, 32'h42979d8c, 32'hc1f22714, 32'h41cbbd9c, 32'h422cd608, 32'h42bcf955, 32'h4210eeae};
test_weights[31192:31199] = '{32'hc222a9ba, 32'h42a9fab4, 32'h427cba8d, 32'h42746dbf, 32'h3f5f9e63, 32'h42c17976, 32'hc0c8fe86, 32'hc283f678};
test_bias[3899:3899] = '{32'hc1ec9d47};
test_output[3899:3899] = '{32'h46313944};
test_input[31200:31207] = '{32'hc2aa7d4e, 32'hc1c0dd66, 32'h427bd75f, 32'h402111da, 32'hc0b659b7, 32'h42bea1ff, 32'hc19b400d, 32'h4299592a};
test_weights[31200:31207] = '{32'hc23da5f9, 32'h41ac9857, 32'h41e658cb, 32'hc2c64b5f, 32'h42add3a2, 32'h42a14337, 32'h42850b05, 32'h42563c73};
test_bias[3900:3900] = '{32'h40175e9b};
test_output[3900:3900] = '{32'h466bd43f};
test_input[31208:31215] = '{32'hc25049e3, 32'h4290f401, 32'h422f312b, 32'h40afc150, 32'h423379eb, 32'hc2881009, 32'h41fac913, 32'hc29be42f};
test_weights[31208:31215] = '{32'h4271d3ac, 32'h424ccf4b, 32'h428dd32e, 32'h3f7be024, 32'h42c27090, 32'hc0627ad0, 32'hc2a2ca2a, 32'hc1547e13};
test_bias[3901:3901] = '{32'hc289a64d};
test_output[3901:3901] = '{32'h45d11e38};
test_input[31216:31223] = '{32'h42a5bc02, 32'h42a97437, 32'h42af76f4, 32'hc2c4810d, 32'h41f1ca76, 32'h424749a4, 32'hc28f5b2e, 32'hc23fbe39};
test_weights[31216:31223] = '{32'h412a63f3, 32'h417f7909, 32'h42b675a6, 32'hbc24b301, 32'h42c168f4, 32'hc1141441, 32'hbfe208c5, 32'h42267e89};
test_bias[3902:3902] = '{32'h40c7807d};
test_output[3902:3902] = '{32'h46295d77};
test_input[31224:31231] = '{32'hc2a968c0, 32'hc1e00c18, 32'hc2395996, 32'hc2bebd82, 32'hc19d437c, 32'h4298c254, 32'hc0fd0a3f, 32'hc2851970};
test_weights[31224:31231] = '{32'h4274b1e4, 32'hc1d0f24a, 32'hc265daec, 32'hc2619752, 32'hc1b057b2, 32'h420e9624, 32'hc25b3c2a, 32'h41d50e8f};
test_bias[3903:3903] = '{32'h409539e2};
test_output[3903:3903] = '{32'h45a926db};
test_input[31232:31239] = '{32'h41c9f295, 32'h423733a8, 32'hc1ac9e5d, 32'h4236eaa3, 32'h412ae393, 32'h4146eba1, 32'hc2074866, 32'h428f7671};
test_weights[31232:31239] = '{32'hc15e8299, 32'hc0c0327e, 32'h420e7281, 32'hc2525ee3, 32'hc09a456d, 32'h42900888, 32'hc2c5cc74, 32'hc28280ff};
test_bias[3904:3904] = '{32'h426d8811};
test_output[3904:3904] = '{32'hc58440bb};
test_input[31240:31247] = '{32'h408178d6, 32'h42965e70, 32'h4286951d, 32'h412f9ca1, 32'h427efa24, 32'h41c901b4, 32'h4299d106, 32'h428131d5};
test_weights[31240:31247] = '{32'hc2a098c7, 32'hc2181912, 32'hc29dbef6, 32'hc2b6421b, 32'h421a74bb, 32'h427c3718, 32'hc1ef0468, 32'hc2935485};
test_bias[3905:3905] = '{32'hc2c61871};
test_output[3905:3905] = '{32'hc644e47b};
test_input[31248:31255] = '{32'hc281152d, 32'hc2a2a509, 32'hc121c05f, 32'hc0b27f93, 32'h429f6f12, 32'hc29be1f1, 32'h41927a6d, 32'h41a30cda};
test_weights[31248:31255] = '{32'h42b29928, 32'hc1bafa89, 32'h414f71c0, 32'h42c4c6ce, 32'h41df3273, 32'h428eb7b5, 32'h411ffb4d, 32'hc28baf61};
test_bias[3906:3906] = '{32'h40788ce9};
test_output[3906:3906] = '{32'hc60e73b5};
test_input[31256:31263] = '{32'h41610104, 32'h425e1510, 32'hc1b6fe5c, 32'hc25b37ec, 32'h42739156, 32'h42894199, 32'hc218796e, 32'h42a88d04};
test_weights[31256:31263] = '{32'h42ba5bf9, 32'h41f134d8, 32'h40e6436a, 32'hc2b36677, 32'h42c3667c, 32'hc109f27a, 32'h4101ffba, 32'hc262b488};
test_bias[3907:3907] = '{32'hc29271b9};
test_output[3907:3907] = '{32'h45f7eec1};
test_input[31264:31271] = '{32'hc0d1a5eb, 32'h426daa31, 32'hc2a89768, 32'hc1a26730, 32'hc28ef9e9, 32'h42c6d01f, 32'hc2921e05, 32'hc1f7dd45};
test_weights[31264:31271] = '{32'h42398359, 32'hc2a1a3e9, 32'h42b931e3, 32'hc1a5d00f, 32'hc2b54944, 32'h419ec80b, 32'hc2bdedb4, 32'h42bbeb0e};
test_bias[3908:3908] = '{32'h425ec761};
test_output[3908:3908] = '{32'h4232e56b};
test_input[31272:31279] = '{32'h422f0fc5, 32'hc212218a, 32'hc2551ed8, 32'hc2b90c8a, 32'h411bb43a, 32'hc288cbeb, 32'hc273ecfe, 32'h41a182a8};
test_weights[31272:31279] = '{32'hc22ac4fe, 32'hc28452e8, 32'hc2a76f2b, 32'h42694ffa, 32'hc2904640, 32'h429f661a, 32'h42513ff0, 32'hc2685549};
test_bias[3909:3909] = '{32'hc216716d};
test_output[3909:3909] = '{32'hc62af54f};
test_input[31280:31287] = '{32'h4283cbf9, 32'h4291be66, 32'h425a0632, 32'hc10af9eb, 32'h4199ce67, 32'hc2531b3d, 32'h425db3d4, 32'hc285805c};
test_weights[31280:31287] = '{32'h42968b17, 32'h42a4d344, 32'hc2c27770, 32'h42006157, 32'h4274dbc1, 32'h4214a391, 32'hc295f4c1, 32'h42994155};
test_bias[3910:3910] = '{32'hc1e60920};
test_output[3910:3910] = '{32'hc592c341};
test_input[31288:31295] = '{32'h4280d6eb, 32'hc22bdf1d, 32'h4283a7da, 32'hc1b1d466, 32'hc2ba226e, 32'h41a7ddd3, 32'hc1934873, 32'h429f48a9};
test_weights[31288:31295] = '{32'hc298088a, 32'h42c03dfe, 32'hc0d457ba, 32'hc22e045d, 32'h41e6b778, 32'hc2adbd0b, 32'hc23c7260, 32'hc098e548};
test_bias[3911:3911] = '{32'hc299b183};
test_output[3911:3911] = '{32'hc644c6e3};
test_input[31296:31303] = '{32'hc2ba1a00, 32'hc12edd4e, 32'hc1aa5b07, 32'hc27ce664, 32'hc265df1f, 32'hbfdb9471, 32'hc2131b1e, 32'h42c2d476};
test_weights[31296:31303] = '{32'hc1c1a009, 32'h42a1a403, 32'hc136c6e8, 32'hc2c2902d, 32'h41e75209, 32'h42b88d48, 32'hc14988b1, 32'h40deb3da};
test_bias[3912:3912] = '{32'h41ee48a0};
test_output[3912:3912] = '{32'h45de4dab};
test_input[31304:31311] = '{32'h4092d30f, 32'h3efeab87, 32'hc24ec13c, 32'hc2a01f93, 32'hc28df9d3, 32'hc28a355c, 32'hc285be14, 32'h42909561};
test_weights[31304:31311] = '{32'hc272b6a9, 32'hc18ca31b, 32'hc1b37863, 32'hc2909150, 32'h41868bfd, 32'h429b0a2c, 32'h421a198d, 32'h41cea24f};
test_bias[3913:3913] = '{32'hc242494a};
test_output[3913:3913] = '{32'hc42233b4};
test_input[31312:31319] = '{32'hc299ed27, 32'h41f4eaec, 32'hc2a3a572, 32'h418a25f5, 32'hc2019921, 32'h400b3f68, 32'hc24b45e6, 32'h41491f1b};
test_weights[31312:31319] = '{32'hc2afc13c, 32'h42c79115, 32'hc1d8ca93, 32'h429b9d68, 32'hc178aa9b, 32'hc2226643, 32'h411c6fb0, 32'h42be3dfd};
test_bias[3914:3914] = '{32'hc1e51f91};
test_output[3914:3914] = '{32'h466201f2};
test_input[31320:31327] = '{32'h42beab84, 32'hc016d8a3, 32'h422630e8, 32'h4197e3ee, 32'h41f34b6c, 32'h41b5de9f, 32'h42b2ca9d, 32'h41dc6d35};
test_weights[31320:31327] = '{32'h428903a9, 32'hc2814a8a, 32'h42468016, 32'hc2a4fe70, 32'hc13ca5f9, 32'hc12113c2, 32'hc2261654, 32'h42490018};
test_bias[3915:3915] = '{32'hc160ac7c};
test_output[3915:3915] = '{32'h4584d199};
test_input[31328:31335] = '{32'h427c192b, 32'hc1d252f9, 32'h42bc9f04, 32'h41a1e828, 32'h423833ab, 32'h4207e2c4, 32'h42a8ebdf, 32'h4280353d};
test_weights[31328:31335] = '{32'h4180e1c8, 32'hc1fe0bbc, 32'h421e5a47, 32'h42216b94, 32'hc1f20e0a, 32'h42052b9a, 32'h429c29b2, 32'hc248da7a};
test_bias[3916:3916] = '{32'hc2396468};
test_output[3916:3916] = '{32'h4613ef0b};
test_input[31336:31343] = '{32'hc23935b1, 32'hc21c3ae5, 32'h4287a780, 32'hc1c9b2fc, 32'hc19431ad, 32'h4235dad8, 32'hc17a1f05, 32'h42c036ea};
test_weights[31336:31343] = '{32'hc2599e1f, 32'hc2ab1781, 32'h42094043, 32'hc2bd2b87, 32'hc29f0a20, 32'h3f20af0f, 32'hc2a8f132, 32'h42846645};
test_bias[3917:3917] = '{32'h42bdb0d0};
test_output[3917:3917] = '{32'h469b170b};
test_input[31344:31351] = '{32'h410bf9f1, 32'h42b1d131, 32'h40ad9248, 32'hc2985d22, 32'h42b651ab, 32'hc1f6fd13, 32'hc14551c2, 32'hc20d2758};
test_weights[31344:31351] = '{32'h42c306d1, 32'hc21ee537, 32'hc29062ed, 32'h41aaebf1, 32'hc2374acb, 32'h424ceb56, 32'h41a4360b, 32'h42be99c6};
test_bias[3918:3918] = '{32'h415426e6};
test_output[3918:3918] = '{32'hc65bae9b};
test_input[31352:31359] = '{32'hc24b22b3, 32'h41b446c2, 32'hc2a6f921, 32'hc2a04d79, 32'h42a3d001, 32'hc1bce7af, 32'h419f731d, 32'hc2aa9425};
test_weights[31352:31359] = '{32'hc2208eb5, 32'hc0bcc3a0, 32'hc1143678, 32'h423f25bf, 32'hc2a2b731, 32'hc2c67ef8, 32'h42184b7d, 32'hc1807206};
test_bias[3919:3919] = '{32'hc29845a8};
test_output[3919:3919] = '{32'hc555b5ff};
test_input[31360:31367] = '{32'h412fdb68, 32'hc2aefa4c, 32'h42c2f48c, 32'hc203935f, 32'hc29b2059, 32'hc1a5c3b3, 32'hc241245e, 32'h427b4c9a};
test_weights[31360:31367] = '{32'hc1eba25c, 32'hc15a81e1, 32'h42b034cc, 32'h4191299f, 32'h42833515, 32'hc2013bb4, 32'hc0361cac, 32'h40e2e785};
test_bias[3920:3920] = '{32'hc242d9f5};
test_output[3920:3920] = '{32'h459b8bb6};
test_input[31368:31375] = '{32'hc2a60cc3, 32'hc13a476b, 32'hc191b500, 32'h40505a42, 32'h41050fb9, 32'hbfd836a5, 32'hc1c0c9f6, 32'hc2b96ae7};
test_weights[31368:31375] = '{32'h4289418e, 32'hc1a2258b, 32'hc2bf561c, 32'hc2c3590d, 32'h425cbd59, 32'hc2347188, 32'h427d79ba, 32'hc1476115};
test_bias[3921:3921] = '{32'h42b5058f};
test_output[3921:3921] = '{32'hc56c7982};
test_input[31376:31383] = '{32'h429b538c, 32'h419df966, 32'hc205020d, 32'h42b226a7, 32'hc2127b07, 32'h42af0ed9, 32'h42b26e83, 32'h41db4750};
test_weights[31376:31383] = '{32'h3f97c435, 32'hc2882c56, 32'hc1286333, 32'h42c1f3d2, 32'h42327913, 32'h42ba15c8, 32'h41796329, 32'hc1a30788};
test_bias[3922:3922] = '{32'h42c0668e};
test_output[3922:3922] = '{32'h466d17ca};
test_input[31384:31391] = '{32'h42c556a0, 32'h42305f9d, 32'hc245c0be, 32'h41ae02eb, 32'hc29cbe8c, 32'hc1e9ebab, 32'h4291d68a, 32'h42241d95};
test_weights[31384:31391] = '{32'h423b9fb0, 32'hc150c832, 32'h42ab65e4, 32'h402327b4, 32'hc2abeee1, 32'h42aede68, 32'h424acc7f, 32'hc2609f3d};
test_bias[3923:3923] = '{32'hc149b5b2};
test_output[3923:3923] = '{32'h45a9c4e6};
test_input[31392:31399] = '{32'h4232d6e5, 32'h40658284, 32'h414749ad, 32'h42915a0a, 32'hc189b4f4, 32'hc2bd1728, 32'h42ae4832, 32'h42acb832};
test_weights[31392:31399] = '{32'hc284805f, 32'hc2846a8d, 32'hc2717db4, 32'hc1fd6a79, 32'hc280f65a, 32'h42a8402c, 32'hc21b6b2c, 32'hc2b727cf};
test_bias[3924:3924] = '{32'hc0951a47};
test_output[3924:3924] = '{32'hc6be98e6};
test_input[31400:31407] = '{32'hc27deb05, 32'h41df9570, 32'h42668807, 32'hc28d4e2c, 32'hc2b4513f, 32'h42be6624, 32'hc2b2f95b, 32'h40ca53ef};
test_weights[31400:31407] = '{32'h41dffb6e, 32'h425e8b18, 32'hc2a1bcf3, 32'hc15f10cb, 32'hc17e4537, 32'h428dc4e2, 32'hc1211493, 32'hbc057a57};
test_bias[3925:3925] = '{32'hc29c90a0};
test_output[3925:3925] = '{32'h459f8bba};
test_input[31408:31415] = '{32'h42b70f85, 32'h42b1f872, 32'hc244e745, 32'h42b45e80, 32'hc28466e8, 32'hc1c021b8, 32'h41a40f68, 32'hc2c212f8};
test_weights[31408:31415] = '{32'hc28a5c61, 32'hc2b8de29, 32'hc006eced, 32'h4280e931, 32'h42b01148, 32'hc1a78225, 32'h42827706, 32'hc2aa6ffc};
test_bias[3926:3926] = '{32'h42910626};
test_output[3926:3926] = '{32'hc585f0d7};
test_input[31416:31423] = '{32'hc2bf8699, 32'hc27e8614, 32'hc1c9e6fe, 32'h42a502ff, 32'hc1b32b2f, 32'hc2b7b845, 32'hc289520c, 32'h41667238};
test_weights[31416:31423] = '{32'hc112f500, 32'hc28e2b7c, 32'hc294950d, 32'h42aa098d, 32'h422bdd80, 32'hc26409d9, 32'h419b83c6, 32'h413e86a2};
test_bias[3927:3927] = '{32'hc299ddfb};
test_output[3927:3927] = '{32'h46875d75};
test_input[31424:31431] = '{32'hc2b340a6, 32'hc0c18042, 32'h41afc429, 32'hc2ac70a7, 32'h421f876f, 32'h42c40802, 32'h42acf2e4, 32'h424256a4};
test_weights[31424:31431] = '{32'h42aa3c72, 32'hc2330a02, 32'hc2b0aa4b, 32'h420e3149, 32'hc2276152, 32'hc1ea19b8, 32'h428376e1, 32'hc23e2cad};
test_bias[3928:3928] = '{32'hc294349e};
test_output[3928:3928] = '{32'hc6548306};
test_input[31432:31439] = '{32'hc284bdb3, 32'h41f77644, 32'h422b5801, 32'h425b8e10, 32'hc2a7ecad, 32'hc23253b6, 32'hc08df36e, 32'h42c28dec};
test_weights[31432:31439] = '{32'h42aa8639, 32'h412885ef, 32'h41d6a597, 32'h4293c597, 32'h428b9bc0, 32'hc252bad7, 32'hc2079925, 32'h428e872d};
test_bias[3929:3929] = '{32'h424fef99};
test_output[3929:3929] = '{32'h455a6399};
test_input[31440:31447] = '{32'h42293e11, 32'hc29047ce, 32'h419c96bb, 32'h428172c4, 32'h41052e7c, 32'h42aeaebe, 32'h42b3e783, 32'hc2b0fba8};
test_weights[31440:31447] = '{32'h428488a7, 32'h429f9289, 32'hc2c5061b, 32'hc07b4e9f, 32'h4249dfc7, 32'hc285b907, 32'h4203f7b7, 32'h4200a06a};
test_bias[3930:3930] = '{32'hc29881a4};
test_output[3930:3930] = '{32'hc62430d1};
test_input[31448:31455] = '{32'hc14de2e6, 32'h42040cc4, 32'h42b5cd57, 32'hc24b0a64, 32'hc24773a1, 32'hc289b856, 32'h4139feeb, 32'h42970b01};
test_weights[31448:31455] = '{32'hc291553b, 32'h42395287, 32'h40061180, 32'h42adf95f, 32'hc264b5fe, 32'hc2507706, 32'h4269b0c5, 32'hc2c2ee09};
test_bias[3931:3931] = '{32'hc17a838a};
test_output[3931:3931] = '{32'hc4fc3de2};
test_input[31456:31463] = '{32'hc29193b2, 32'hc1ee78cb, 32'hbf75c00b, 32'h419a0b16, 32'h42859132, 32'hc0e0c144, 32'h41ae25f4, 32'hc225e9ee};
test_weights[31456:31463] = '{32'h428fa2e1, 32'h4290ed59, 32'hc1ecf344, 32'h42b7fced, 32'hc28f50b4, 32'hc27161fb, 32'hc0c7aae7, 32'h41ffdeb3};
test_bias[3932:3932] = '{32'hc24865ba};
test_output[3932:3932] = '{32'hc6331836};
test_input[31464:31471] = '{32'hc2636f92, 32'hc11b5e20, 32'h426470a3, 32'hc2b9409a, 32'h42a6e227, 32'hc127f9aa, 32'hc2bb9b5f, 32'hc2b9ddba};
test_weights[31464:31471] = '{32'hc2109ad8, 32'hc1d8f4de, 32'hc20d20d9, 32'hc2157652, 32'h42003844, 32'h42bba81d, 32'hc23e6380, 32'h429000b2};
test_bias[3933:3933] = '{32'h41f6a5fc};
test_output[3933:3933] = '{32'h454bae70};
test_input[31472:31479] = '{32'h4216482c, 32'h4205ba10, 32'h4286ce53, 32'hc2a8d7a0, 32'h42a364e4, 32'h41cd0817, 32'hc0e6b6f0, 32'h4204c7f1};
test_weights[31472:31479] = '{32'hc144612b, 32'h4290adf5, 32'h42b23d6d, 32'h4243e7db, 32'hc2af3f58, 32'h42ad8f7c, 32'h42196789, 32'h3e60105a};
test_bias[3934:3934] = '{32'hc280c5b3};
test_output[3934:3934] = '{32'hc4b3d0c0};
test_input[31480:31487] = '{32'h42b11b8f, 32'h41fb8a52, 32'h42974f7e, 32'hc2642635, 32'hc139cca1, 32'hc139c512, 32'hc190dd2c, 32'hc1cf6d7b};
test_weights[31480:31487] = '{32'h424ec6af, 32'h425a4c60, 32'h42bacd50, 32'h428f9f6f, 32'h41d3d6be, 32'h41d323ec, 32'h42786c4a, 32'h418702a3};
test_bias[3935:3935] = '{32'h41296557};
test_output[3935:3935] = '{32'h45ddd3e4};
test_input[31488:31495] = '{32'h419b588f, 32'hc217f08d, 32'hc2beb1ab, 32'h4273b0e7, 32'h42a84755, 32'h4261ec44, 32'h4264f2e2, 32'h40edc9c2};
test_weights[31488:31495] = '{32'h40dc7e5b, 32'hc288d811, 32'h42663d10, 32'hc20cffb9, 32'h42bbee5a, 32'hc2158dc9, 32'hc2b24268, 32'hc28ad87e};
test_bias[3936:3936] = '{32'hc2ad506d};
test_output[3936:3936] = '{32'hc5966387};
test_input[31496:31503] = '{32'h415ab8ae, 32'hc2b3e62b, 32'h42a074ac, 32'hc219f1ac, 32'h429061c8, 32'h4299297f, 32'h42b65cae, 32'h42420451};
test_weights[31496:31503] = '{32'hc25fd692, 32'h425d17f8, 32'h42194db5, 32'hc20dc1d6, 32'hc295e215, 32'h42739a40, 32'h41d33d73, 32'h42c65d1b};
test_bias[3937:3937] = '{32'hc1bb61de};
test_output[3937:3937] = '{32'h45a0f4e2};
test_input[31504:31511] = '{32'h41b2cee8, 32'hc2390fda, 32'hc12469ac, 32'hc21cfe9b, 32'hc09f541c, 32'h42c1a46f, 32'h42b5fd4d, 32'h429d3782};
test_weights[31504:31511] = '{32'hc2aaed7e, 32'h4209ca33, 32'h40cecdb0, 32'h42b1e3fc, 32'h429e52a7, 32'h41ce3423, 32'h426a773f, 32'hc1ba6e1e};
test_bias[3938:3938] = '{32'h42ba7b94};
test_output[3938:3938] = '{32'hc4aa9678};
test_input[31512:31519] = '{32'hc27eda50, 32'h42ac1695, 32'hc2c533bb, 32'hc29f8de8, 32'h42bbe9d8, 32'h41c9174b, 32'hc1c43a26, 32'hc0fd44c3};
test_weights[31512:31519] = '{32'h41b42d32, 32'h41f38f8b, 32'h42a1e95a, 32'hc1fd96dd, 32'h42a0a167, 32'h41282760, 32'hc2bb0e02, 32'h4283ae1f};
test_bias[3939:3939] = '{32'h42697e89};
test_output[3939:3939] = '{32'h45a7e6d3};
test_input[31520:31527] = '{32'hc1c10761, 32'h41cf7102, 32'h4256d568, 32'h403f05d9, 32'hc2b693ce, 32'h40b0c475, 32'hc272414c, 32'h42934176};
test_weights[31520:31527] = '{32'h429f868c, 32'h41575ad9, 32'h42bcb037, 32'hc291db98, 32'h4218ffed, 32'h42a83412, 32'h42b51a1f, 32'hc21fdc1a};
test_bias[3940:3940] = '{32'h42760ea4};
test_output[3940:3940] = '{32'hc5fdb3eb};
test_input[31528:31535] = '{32'hc2715c74, 32'hc28b4f15, 32'hc2533988, 32'h408d5d8d, 32'h428a4aef, 32'h427d40f9, 32'h41ef3e4d, 32'h41ee3ca0};
test_weights[31528:31535] = '{32'h41015245, 32'hc2c00403, 32'hc1281cf3, 32'hc2ab72e1, 32'h42c1dd20, 32'h3dccdfc7, 32'h41ad2e9e, 32'h41752bfb};
test_bias[3941:3941] = '{32'hc2bebf46};
test_output[3941:3941] = '{32'h465c33d3};
test_input[31536:31543] = '{32'h42288566, 32'h421996ca, 32'h4283d571, 32'h429c8488, 32'hc242798d, 32'hc202693f, 32'hc1b52426, 32'h42c4e27f};
test_weights[31536:31543] = '{32'hbebb9f33, 32'h42a35798, 32'hc2248ec2, 32'hc227edee, 32'h41a2f232, 32'h41bda1a3, 32'h425233a3, 32'hc2b23ed3};
test_bias[3942:3942] = '{32'h3eb27ed3};
test_output[3942:3942] = '{32'hc6642b5c};
test_input[31544:31551] = '{32'hc19842c0, 32'h41045f83, 32'h42ac5427, 32'hc279d348, 32'hc213813d, 32'h42361ab0, 32'h426254dd, 32'hc1b1cf5f};
test_weights[31544:31551] = '{32'hc1e16fdf, 32'h42698466, 32'h4211b8a7, 32'hc1389710, 32'hbfb3d725, 32'h426ebaf8, 32'hc14b6cbe, 32'hc21bf856};
test_bias[3943:3943] = '{32'h415b321a};
test_output[3943:3943] = '{32'h45f40606};
test_input[31552:31559] = '{32'hc2923dc3, 32'h42942a28, 32'h419739a3, 32'hc2110f0b, 32'hc2c19675, 32'hc2a6d6ee, 32'hc2c639b9, 32'hc22424cd};
test_weights[31552:31559] = '{32'hbf77704e, 32'hc26d1b9a, 32'hc290004a, 32'hc2b0396e, 32'h42521ef6, 32'h421199b5, 32'hc20d5bfc, 32'hc2a8aea7};
test_bias[3944:3944] = '{32'h42b91c16};
test_output[3944:3944] = '{32'hc55df456};
test_input[31560:31567] = '{32'hc09b1d9d, 32'h42183951, 32'hc2471ec1, 32'hc233c151, 32'h415c8223, 32'h42769e9a, 32'h428438d5, 32'hc258d861};
test_weights[31560:31567] = '{32'hc0ee63c4, 32'hc2993617, 32'h41f54b29, 32'hc1d107f6, 32'h426d043c, 32'hc0f27a75, 32'hc11181cb, 32'hc29f2ca3};
test_bias[3945:3945] = '{32'h422a8a76};
test_output[3945:3945] = '{32'h445a82d0};
test_input[31568:31575] = '{32'hc20f69c2, 32'h41fb38d7, 32'hc2bc9781, 32'h42b291b9, 32'hc2c07b0f, 32'h41dec205, 32'hc2b6745d, 32'hc1a3e965};
test_weights[31568:31575] = '{32'h42187d7e, 32'h42a4e393, 32'h413f0d9c, 32'h42321779, 32'h429ed52a, 32'hc2b4c975, 32'h42126b46, 32'hc08c13fc};
test_bias[3946:3946] = '{32'h42955468};
test_output[3946:3946] = '{32'hc610be86};
test_input[31576:31583] = '{32'h429c233f, 32'h4204b7ea, 32'hc20fd329, 32'hc0b2e90c, 32'hc16e90c1, 32'hc1fe81d7, 32'hc26bb171, 32'hc1c83100};
test_weights[31576:31583] = '{32'hc2b4db53, 32'h42266a77, 32'h4105e32b, 32'h403c59ae, 32'hc202b14e, 32'h42b1356f, 32'h41ee3f52, 32'hc2ba276a};
test_bias[3947:3947] = '{32'hc150c5f3};
test_output[3947:3947] = '{32'hc5f2b725};
test_input[31584:31591] = '{32'h42061ab1, 32'h41c130b0, 32'h428b3088, 32'h42b38d6a, 32'hc2461f9e, 32'hc28e2b92, 32'hc272134e, 32'hc26abef8};
test_weights[31584:31591] = '{32'hc29a1288, 32'hc25a69b3, 32'hc2a5597a, 32'h40b26d20, 32'hbe2036d5, 32'hc24b4b64, 32'hc23dfb89, 32'h4192e840};
test_bias[3948:3948] = '{32'h42148209};
test_output[3948:3948] = '{32'hc567419f};
test_input[31592:31599] = '{32'h41d9ee55, 32'h42bdab97, 32'h42aa566f, 32'hc222cbcf, 32'h42a6ef63, 32'h3f5a402c, 32'h42343f00, 32'h42ad8b15};
test_weights[31592:31599] = '{32'h41fc578e, 32'h423332c2, 32'hc2bd460a, 32'hc20abbe0, 32'h41b9f6db, 32'hc2b86e17, 32'hc273b3ba, 32'h428c0415};
test_bias[3949:3949] = '{32'h41e85e09};
test_output[3949:3949] = '{32'h4565f4ee};
test_input[31600:31607] = '{32'h420fd6be, 32'h42958211, 32'h425bd959, 32'hc0766b67, 32'hc12ddb10, 32'hc252a464, 32'hc2820f91, 32'hc2b36a1e};
test_weights[31600:31607] = '{32'hc0a0ef98, 32'h3fb8ec0b, 32'h41a0559b, 32'h426d686b, 32'h42026481, 32'h415008db, 32'h41844d8d, 32'hc1f09804};
test_bias[3950:3950] = '{32'h40046ec8};
test_output[3950:3950] = '{32'h44ad378f};
test_input[31608:31615] = '{32'hc0800d7a, 32'h420fc78f, 32'h428ad173, 32'h428ddbd3, 32'h4122569a, 32'h41f69117, 32'hc200461c, 32'hc14cdd2e};
test_weights[31608:31615] = '{32'h42226e2b, 32'h42a7c58e, 32'hc26a24d1, 32'h424a7e76, 32'hc2c3777f, 32'h42b00f77, 32'h428f3c23, 32'hc2661571};
test_bias[3951:3951] = '{32'hc20d92a5};
test_output[3951:3951] = '{32'h451ca869};
test_input[31616:31623] = '{32'hc28c906d, 32'hc02bc1ba, 32'h42c23288, 32'hc1d7e368, 32'h428b1a01, 32'hc2b59733, 32'h41e3e6d9, 32'hc1a6508e};
test_weights[31616:31623] = '{32'h428dfd67, 32'h3fe7f639, 32'hc2a87b45, 32'h42bbde9e, 32'h42329077, 32'h41a3e7cc, 32'hc236a5a8, 32'hc269022a};
test_bias[3952:3952] = '{32'hc29af5e3};
test_output[3952:3952] = '{32'hc6649f30};
test_input[31624:31631] = '{32'h42309b03, 32'hc1a72d5c, 32'hc2c07f04, 32'hc2284718, 32'hc29a1019, 32'hc1905bc2, 32'hc22c3763, 32'hc2bac446};
test_weights[31624:31631] = '{32'hc27b4f54, 32'h41d93fc8, 32'hc191d035, 32'h4258bf53, 32'h41623e90, 32'hc07a27c5, 32'h426c73fc, 32'hc2c0bfeb};
test_bias[3953:3953] = '{32'hc28cc91f};
test_output[3953:3953] = '{32'h44bb5cb4};
test_input[31632:31639] = '{32'h4117fca9, 32'hc2b1071a, 32'hbf1d81b7, 32'hc1e5da39, 32'h41080681, 32'hc20840bf, 32'h42b4c235, 32'hc00ce597};
test_weights[31632:31639] = '{32'h41bdeba3, 32'h424ea98a, 32'h42b5e167, 32'h425ac51d, 32'h413b9a07, 32'hc2073cd0, 32'h4089dd59, 32'hc2396856};
test_bias[3954:3954] = '{32'h428f8294};
test_output[3954:3954] = '{32'hc582038c};
test_input[31640:31647] = '{32'h40be1f50, 32'h4253dabf, 32'hc2021e41, 32'hc2052b9d, 32'hc2100dcd, 32'h424ae2b5, 32'hc198f374, 32'hc0fca7ee};
test_weights[31640:31647] = '{32'hc2a2e9d6, 32'h41f84fb3, 32'h42966a70, 32'hc200876b, 32'h4023f71c, 32'h415d4434, 32'h42a86143, 32'h41b12f12};
test_bias[3955:3955] = '{32'h42496778};
test_output[3955:3955] = '{32'hc4a7b69d};
test_input[31648:31655] = '{32'h4136e377, 32'h41f63fc7, 32'hc26d7f8f, 32'hc12ddffc, 32'h42ac615c, 32'hc1dd3e2e, 32'h42abc752, 32'h42aa4602};
test_weights[31648:31655] = '{32'hc2a750a3, 32'hc2a2401d, 32'h4296670d, 32'hc2be206d, 32'h42bcc299, 32'hc112ed1c, 32'hc23d146f, 32'h428fb736};
test_bias[3956:3956] = '{32'h426d7969};
test_output[3956:3956] = '{32'h456245df};
test_input[31656:31663] = '{32'hc27e9502, 32'h42150b66, 32'hc236d1ef, 32'h42a41ddc, 32'h4222b2b8, 32'hc28fb5fe, 32'h42880047, 32'hc2b712ec};
test_weights[31656:31663] = '{32'hc20f114a, 32'hbf0ed9a1, 32'h4285bae4, 32'h4221adb1, 32'hc2520d81, 32'hc1e183f0, 32'h42a208dc, 32'hc29f062c};
test_bias[3957:3957] = '{32'hc2223a4c};
test_output[3957:3957] = '{32'h466cc384};
test_input[31664:31671] = '{32'hc2849695, 32'h42538872, 32'h427e0f25, 32'h429b0e14, 32'h41e820b1, 32'h41387f4d, 32'hc28201d1, 32'hc12a9a28};
test_weights[31664:31671] = '{32'hc012280c, 32'h41b02d83, 32'hc01be29b, 32'h42b45bb3, 32'h41242b52, 32'hc2c532e7, 32'hc28a0bfa, 32'hc2b09b52};
test_bias[3958:3958] = '{32'h42504a22};
test_output[3958:3958] = '{32'h4647e739};
test_input[31672:31679] = '{32'hc2bdcc35, 32'hc230f9c3, 32'h42b5e607, 32'h421cb40b, 32'h412ceec6, 32'hbf7e6dc0, 32'h428df257, 32'h4261d352};
test_weights[31672:31679] = '{32'h42baec8b, 32'hc2b111b1, 32'h41c15063, 32'hc18c66a7, 32'h42565625, 32'h4262e7b6, 32'hc2a36958, 32'h42a38b6e};
test_bias[3959:3959] = '{32'hc28f9375};
test_output[3959:3959] = '{32'hc5826c1b};
test_input[31680:31687] = '{32'h42c76314, 32'h4259d31e, 32'hc2b7d268, 32'h422b749d, 32'h42285da9, 32'h42808c0f, 32'h428bf685, 32'h40821ed7};
test_weights[31680:31687] = '{32'hc192949d, 32'h40f12164, 32'h423c2d5e, 32'hc2929485, 32'h4253f595, 32'h41b786ed, 32'h41f07188, 32'h42a676c6};
test_bias[3960:3960] = '{32'h42af3d5c};
test_output[3960:3960] = '{32'hc525761b};
test_input[31688:31695] = '{32'h42485de0, 32'hc2141faf, 32'hc23b41c8, 32'h429f0351, 32'hc051d866, 32'hc2b563e9, 32'h42181176, 32'hc28fee2d};
test_weights[31688:31695] = '{32'h421d1ee1, 32'h426e2c90, 32'h42b8f9b4, 32'hc1fa4d5a, 32'h4180d6c9, 32'h4273a928, 32'hc2b44869, 32'h3efbb51c};
test_bias[3961:3961] = '{32'hc2921c41};
test_output[3961:3961] = '{32'hc67c9e1d};
test_input[31696:31703] = '{32'h42c24a85, 32'hc218ae94, 32'h41105e30, 32'h41d77d14, 32'h41e9de3c, 32'h4293996d, 32'h4290215d, 32'h42a4164b};
test_weights[31696:31703] = '{32'h420e0a0d, 32'hc2c62c81, 32'h41d9678b, 32'h4287302b, 32'hc276bc7f, 32'hc156285f, 32'h42bc8d8f, 32'h424aab66};
test_bias[3962:3962] = '{32'hc241abca};
test_output[3962:3962] = '{32'h46880287};
test_input[31704:31711] = '{32'h41218df1, 32'hc210544f, 32'hc2b2b25f, 32'h426060ce, 32'hc297eeda, 32'hc2b4de33, 32'h42025aca, 32'hc2acc37f};
test_weights[31704:31711] = '{32'hc2b0563c, 32'h425e7331, 32'hc246f937, 32'hc20e163b, 32'h4108f206, 32'hc2bd85ae, 32'h41ca4dd2, 32'hc28f4d69};
test_bias[3963:3963] = '{32'h42b56fbe};
test_output[3963:3963] = '{32'h4663ca8d};
test_input[31712:31719] = '{32'h428043d8, 32'hc1bc21d5, 32'h428a54e8, 32'hc1ba52ef, 32'hc27fe053, 32'h420be4fb, 32'hc29c7603, 32'hc2b963a9};
test_weights[31712:31719] = '{32'h4129b403, 32'h429e4d16, 32'hc2c6bd28, 32'hc2c5e25f, 32'hc2a00cd8, 32'hc20aec13, 32'h41f9fd5f, 32'hbf11e646};
test_bias[3964:3964] = '{32'h4232bd99};
test_output[3964:3964] = '{32'hc5830263};
test_input[31720:31727] = '{32'h41c6af9e, 32'hc237b225, 32'h428e7887, 32'h429e8d24, 32'h42b69d7b, 32'hc2b4b4c0, 32'hc13e0e59, 32'h4248d9b4};
test_weights[31720:31727] = '{32'hc2b2dc12, 32'h423b6185, 32'hc1ea995f, 32'h41ee794d, 32'hc157fc0f, 32'h41c8b998, 32'h4253da1e, 32'h40f48f5f};
test_bias[3965:3965] = '{32'hc1f72e6a};
test_output[3965:3965] = '{32'hc5f61060};
test_input[31728:31735] = '{32'hbf0b118a, 32'h412cfda6, 32'h42a23a47, 32'h42b7e01a, 32'h429e26ee, 32'hc18e8e2d, 32'hc2b9aa83, 32'hc297efb9};
test_weights[31728:31735] = '{32'hc1fab95e, 32'hc1243771, 32'hc228a69e, 32'hc2810070, 32'h4296db5e, 32'h42420ed2, 32'h422ace39, 32'hc1d6de0d};
test_bias[3966:3966] = '{32'h429bef6c};
test_output[3966:3966] = '{32'hc5c16d27};
test_input[31736:31743] = '{32'hc26652ba, 32'hc25bbe52, 32'hc26ea21b, 32'h40f271a3, 32'h41f88440, 32'hbfab553c, 32'hc2795cbe, 32'hc1d815d8};
test_weights[31736:31743] = '{32'hc2b9553a, 32'h42894dcb, 32'hc2a9f5dc, 32'hc2adab0e, 32'h4246196d, 32'hc1464900, 32'hc2999cc7, 32'h42b9359e};
test_bias[3967:3967] = '{32'hc2a9c9e3};
test_output[3967:3967] = '{32'h461814ec};
test_input[31744:31751] = '{32'hc2b1664a, 32'hc17d9ce0, 32'hc201ef9f, 32'hc290280e, 32'hc096b09a, 32'hc20349a6, 32'h42548596, 32'h41491524};
test_weights[31744:31751] = '{32'hc2a866c1, 32'h41531d89, 32'hc29287ab, 32'h42a181b4, 32'hc296a932, 32'h42c2697e, 32'h406ac798, 32'hc288e155};
test_bias[3968:3968] = '{32'h413f546a};
test_output[3968:3968] = '{32'h43a4e60d};
test_input[31752:31759] = '{32'h421855e6, 32'h428c3460, 32'h42c549fb, 32'h41688735, 32'hc2abfbd6, 32'h4234b58d, 32'hc11f4e87, 32'hc29e557d};
test_weights[31752:31759] = '{32'hc091900b, 32'h42045854, 32'h42601b7a, 32'hc1d22410, 32'hc20a78e7, 32'h420772ee, 32'hc1fe632f, 32'hc27a2e5f};
test_bias[3969:3969] = '{32'h4177c4ef};
test_output[3969:3969] = '{32'h468572ee};
test_input[31760:31767] = '{32'h4256646f, 32'hc2b2515d, 32'hc29fbd92, 32'h420ea05b, 32'hc242e9eb, 32'hc21fcd38, 32'h40f9e4fd, 32'hbff7da9d};
test_weights[31760:31767] = '{32'hc29cd281, 32'h42b8aefd, 32'h423f9f98, 32'h42a67ac3, 32'hc025c859, 32'h42b6a555, 32'hbf414be4, 32'hc0fd0dee};
test_bias[3970:3970] = '{32'h407c0488};
test_output[3970:3970] = '{32'hc6834597};
test_input[31768:31775] = '{32'h42b5217d, 32'h42b96703, 32'h4298f2c7, 32'hc23803e6, 32'h4169d240, 32'hc2935473, 32'hc2098006, 32'h42900ef1};
test_weights[31768:31775] = '{32'h4103a282, 32'h42a779f2, 32'hc2c52332, 32'hc2a3073b, 32'hc226d9a7, 32'hc2223f7e, 32'hc21b0649, 32'hc2a6dc1e};
test_bias[3971:3971] = '{32'h4203f672};
test_output[3971:3971] = '{32'h45195fc9};
test_input[31776:31783] = '{32'h429b42c4, 32'h4084d86c, 32'hc18fe0e9, 32'h421627cf, 32'hc1733101, 32'hc2358680, 32'h422186e8, 32'h429e4a00};
test_weights[31776:31783] = '{32'h4297c879, 32'h42b9934d, 32'h415353cf, 32'h422c50a5, 32'h41dd6cf8, 32'h4291505d, 32'h42472cf2, 32'hc1f57d4c};
test_bias[3972:3972] = '{32'hc23cda4c};
test_output[3972:3972] = '{32'h45591386};
test_input[31784:31791] = '{32'hc15a68ab, 32'hc2a3edb7, 32'hc2614dbe, 32'h42b01af2, 32'h4195db7a, 32'h42636f30, 32'hc246ef28, 32'hc1bd2780};
test_weights[31784:31791] = '{32'hc28c5f90, 32'h420d4fe9, 32'h429bc2a8, 32'hbfe3ff8c, 32'hc257a368, 32'hc18116be, 32'h41b7c8d2, 32'h40c80dfe};
test_bias[3973:3973] = '{32'h4283a12e};
test_output[3973:3973] = '{32'hc61683ae};
test_input[31792:31799] = '{32'hc0c5d9ed, 32'hc1ed9e75, 32'h4200351c, 32'hc1d9d67e, 32'h4281bab5, 32'hc26c264b, 32'hc125496e, 32'h40e15636};
test_weights[31792:31799] = '{32'hc2790d0b, 32'h41197278, 32'h3fa44b15, 32'hbf25a84d, 32'hc232de15, 32'h424dd6ef, 32'hc108f496, 32'h4064905c};
test_bias[3974:3974] = '{32'h42826ec8};
test_output[3974:3974] = '{32'hc5af079b};
test_input[31800:31807] = '{32'h423c8031, 32'h41d0048d, 32'hc18f0bb9, 32'hc0853a08, 32'h428151ac, 32'h428e2221, 32'h4284c5ea, 32'h41a196e2};
test_weights[31800:31807] = '{32'hc2b10ef2, 32'hc25de0fa, 32'h42bc592a, 32'hc28d6a96, 32'h42ad7b46, 32'hc2b88520, 32'h42084070, 32'h408e4049};
test_bias[3975:3975] = '{32'hc2322715};
test_output[3975:3975] = '{32'hc5b069dd};
test_input[31808:31815] = '{32'h428ff527, 32'hc158c38e, 32'hc2be5b98, 32'hc28a354e, 32'h42c1e2cb, 32'h42a12e18, 32'hc24735d6, 32'hc251f7d0};
test_weights[31808:31815] = '{32'h42875107, 32'hc17bb026, 32'h42c04537, 32'h429fbc4a, 32'hc291c9a4, 32'hc2372afb, 32'hc191e9ac, 32'h42be0533};
test_bias[3976:3976] = '{32'hc279cc37};
test_output[3976:3976] = '{32'hc6bf48e4};
test_input[31816:31823] = '{32'h4222e12c, 32'h40a9fd58, 32'h42c66fd2, 32'h41e8c757, 32'hc1cc87c1, 32'hc1c3e87a, 32'h410aee9d, 32'hc1f9331a};
test_weights[31816:31823] = '{32'hc2a00c20, 32'h4290f5cd, 32'hc2c31cd0, 32'h402f731b, 32'hc2820444, 32'hc256c5b1, 32'hc27dec70, 32'hc2c7d73c};
test_bias[3977:3977] = '{32'hc16c61a6};
test_output[3977:3977] = '{32'hc5d92ddd};
test_input[31824:31831] = '{32'h4234ce3c, 32'h42110cfa, 32'h425ff490, 32'hc1eb1bb3, 32'hc2b0c77b, 32'h42586fdf, 32'h41e52cfc, 32'h42a2ca7c};
test_weights[31824:31831] = '{32'hc130eab8, 32'hc2c10d99, 32'h42a9321e, 32'hc198b089, 32'h412af98c, 32'hc280b696, 32'hc283b502, 32'hc256f8dc};
test_bias[3978:3978] = '{32'h425e673d};
test_output[3978:3978] = '{32'hc611db47};
test_input[31832:31839] = '{32'h42557b53, 32'hc21aa035, 32'hc29a524e, 32'h40fdb05c, 32'h4233581c, 32'hc2c6a075, 32'h423d7fb9, 32'h42b89f58};
test_weights[31832:31839] = '{32'h426f9f0d, 32'h41d3e9c8, 32'hc232fb5c, 32'hc2324e34, 32'hc2b08578, 32'h4267964a, 32'hc21c2567, 32'hc15463d7};
test_bias[3979:3979] = '{32'h3f642251};
test_output[3979:3979] = '{32'hc5eaa4e8};
test_input[31840:31847] = '{32'h415fad6d, 32'hc28425b3, 32'h429cb706, 32'h4107de20, 32'h414691c9, 32'hc2617c52, 32'h424693d6, 32'h41d78179};
test_weights[31840:31847] = '{32'hc270a56c, 32'hc2bc368c, 32'h42561b8f, 32'h427c0b31, 32'h420dfa7a, 32'hc2674e1c, 32'h426a8fe6, 32'hc2bd83d9};
test_bias[3980:3980] = '{32'h413f428a};
test_output[3980:3980] = '{32'h465d8402};
test_input[31848:31855] = '{32'hc1fa1f1f, 32'h42af2fd7, 32'hc25a3f91, 32'h4265c62c, 32'hc2b2a942, 32'h426ec4cc, 32'hc0d095a5, 32'hc2c64c40};
test_weights[31848:31855] = '{32'hc25177e7, 32'hc270bc76, 32'h42b08bb4, 32'h41abb516, 32'hc2bf3d15, 32'h42b535d3, 32'hc2a73d91, 32'hc2aa1c07};
test_bias[3981:3981] = '{32'hc2bd7d55};
test_output[3981:3981] = '{32'h4673feae};
test_input[31856:31863] = '{32'h424ef609, 32'hc0d161cd, 32'hc23a990f, 32'hc2169d01, 32'hc29b7851, 32'h4279cd0a, 32'hc1cc7366, 32'h426da386};
test_weights[31856:31863] = '{32'hc19f35e2, 32'hc28aaf51, 32'hc26edc67, 32'hc1aab5eb, 32'hc28c746e, 32'h422c1f41, 32'hc12689a2, 32'hc281c70d};
test_bias[3982:3982] = '{32'hc2b1c066};
test_output[3982:3982] = '{32'h45e9cd79};
test_input[31864:31871] = '{32'h41c4e490, 32'h418fd223, 32'hc1ce1fb9, 32'hc1f217d9, 32'hc1e43f30, 32'hc18b58a5, 32'h42a2db84, 32'h41f06458};
test_weights[31864:31871] = '{32'hc290a127, 32'hc28f18ff, 32'hc232578f, 32'h42c7d985, 32'h41fafb65, 32'h422f046e, 32'h42358935, 32'h42910d42};
test_bias[3983:3983] = '{32'h4283dad1};
test_output[3983:3983] = '{32'hc4246502};
test_input[31872:31879] = '{32'h420c2bca, 32'h423d279c, 32'hc23dd01c, 32'h42bebfc6, 32'hc025329f, 32'h429ae9db, 32'h421c426c, 32'hc2a93aa5};
test_weights[31872:31879] = '{32'hc0c76200, 32'h429c6ad3, 32'hc268b2de, 32'h4216e895, 32'hc1913f74, 32'hc0a9027d, 32'h427acd7f, 32'hc205b0ba};
test_bias[3984:3984] = '{32'hc27a261d};
test_output[3984:3984] = '{32'h46658df8};
test_input[31880:31887] = '{32'h412fa2d3, 32'hc29e5385, 32'h42c52cc8, 32'h41f8bd83, 32'hc2219520, 32'h42a7c535, 32'hc2c2b0c5, 32'h41014a55};
test_weights[31880:31887] = '{32'hc178793d, 32'hc24c55e3, 32'hc1f4cf73, 32'hc247ab09, 32'h40e0f1b8, 32'h419044e7, 32'h417bcfe7, 32'h42643489};
test_bias[3985:3985] = '{32'hc26dc6e5};
test_output[3985:3985] = '{32'hc4154972};
test_input[31888:31895] = '{32'hc27f05ee, 32'h42244225, 32'h421ad67b, 32'hc21b0653, 32'h42c6a05d, 32'hc1bee964, 32'h42b499c0, 32'h425edf6b};
test_weights[31888:31895] = '{32'h41aceb82, 32'h4268dca8, 32'hc292d4c3, 32'h42a39355, 32'hc218f648, 32'hc28b4740, 32'h428f3e09, 32'h421a3a63};
test_bias[3986:3986] = '{32'hc2212235};
test_output[3986:3986] = '{32'h44b40c85};
test_input[31896:31903] = '{32'hc2c48e64, 32'hc2c501ee, 32'h429f8835, 32'hc17e27f1, 32'h41e8ae0c, 32'h42763faa, 32'hc2954ba6, 32'h42927547};
test_weights[31896:31903] = '{32'h42843260, 32'h42053c63, 32'h414a1a97, 32'hc22c9a66, 32'h426ba561, 32'h41a825ba, 32'hc24386dd, 32'h42272278};
test_bias[3987:3987] = '{32'h41dc0732};
test_output[3987:3987] = '{32'h44cf6fb0};
test_input[31904:31911] = '{32'hc2462fad, 32'h429f4787, 32'h4159c7a0, 32'hc2bb1bda, 32'h4149df05, 32'h42b23cfb, 32'hc275fc1c, 32'hc208d200};
test_weights[31904:31911] = '{32'hc291e118, 32'h40ffe332, 32'hc2ae9468, 32'hc28bb8f7, 32'h422e61df, 32'hc286888d, 32'h42b47655, 32'h425d9b96};
test_bias[3988:3988] = '{32'hc2c5e5f6};
test_output[3988:3988] = '{32'hc553d1a2};
test_input[31912:31919] = '{32'h427c19c2, 32'h429ce03e, 32'hc28f6d88, 32'hc2998931, 32'hc265676b, 32'h418a76c7, 32'hc2805260, 32'h41f9ca7f};
test_weights[31912:31919] = '{32'hc2693076, 32'hc2c2eef5, 32'hc16db629, 32'h420aacdf, 32'h429d2a2e, 32'h41650afa, 32'h4184ca92, 32'hc22621bc};
test_bias[3989:3989] = '{32'hc1d7b067};
test_output[3989:3989] = '{32'hc698d62b};
test_input[31920:31927] = '{32'h41f6b637, 32'h42bb959d, 32'h42ac4cdb, 32'hc0505615, 32'h424c8422, 32'hc2890c1c, 32'hc0525f09, 32'hc284c043};
test_weights[31920:31927] = '{32'h41859a5e, 32'h41f5b85c, 32'hc2b1fbf1, 32'hc22b3d18, 32'h42b44a40, 32'hc24e7029, 32'h428866f7, 32'hc1735887};
test_bias[3990:3990] = '{32'hc2953021};
test_output[3990:3990] = '{32'h4593a62b};
test_input[31928:31935] = '{32'h41965194, 32'hc213213b, 32'hc11dfd64, 32'hc29cb6e6, 32'hc0a66cf1, 32'h4230f0cb, 32'hc2a919de, 32'hc284ed62};
test_weights[31928:31935] = '{32'h42a6838a, 32'hc270b930, 32'hc11edb8a, 32'h41d012e8, 32'hc2a91df0, 32'h428e3d5e, 32'h428be410, 32'hc298a5e5};
test_bias[3991:3991] = '{32'hc18c6222};
test_output[3991:3991] = '{32'h458ea8a2};
test_input[31936:31943] = '{32'h41e378cd, 32'h42a691aa, 32'h41d336ff, 32'hc2674e60, 32'hc26d2c7b, 32'hc23aeff4, 32'h41985b92, 32'h42a26b76};
test_weights[31936:31943] = '{32'h4283febc, 32'hc24fa92f, 32'hc2483611, 32'hc2b485e5, 32'h4276d7af, 32'h42a862ae, 32'hc21c4039, 32'h425ca929};
test_bias[3992:3992] = '{32'hc29ad603};
test_output[3992:3992] = '{32'hc51b4426};
test_input[31944:31951] = '{32'h420f955a, 32'hc29bb26c, 32'h42a3369b, 32'h42b37142, 32'h421f7cf9, 32'hc121d962, 32'hc2b30597, 32'h4256f629};
test_weights[31944:31951] = '{32'hc2b7fed7, 32'h41869891, 32'hc28ea5ff, 32'h42754fe6, 32'h4206c29a, 32'hc2a8a398, 32'h417c1d85, 32'hc2245ff4};
test_bias[3993:3993] = '{32'h4243ca90};
test_output[3993:3993] = '{32'hc5c4fedf};
test_input[31952:31959] = '{32'hc2b1c55a, 32'hc2931403, 32'hc29cf149, 32'h42672e1e, 32'h4223f5fb, 32'h415caa4c, 32'h421bdf90, 32'hc244f1f5};
test_weights[31952:31959] = '{32'h42412a15, 32'h42aee5da, 32'hc28396c7, 32'h428bf75b, 32'hc2a9428b, 32'h428d7bcd, 32'h420ec5cf, 32'h4285d84c};
test_bias[3994:3994] = '{32'h42643d87};
test_output[3994:3994] = '{32'hc5b70060};
test_input[31960:31967] = '{32'hc1d763c3, 32'hc2ae0308, 32'h4280ff96, 32'hc2bce85a, 32'h42a5b8c3, 32'h41b2afd0, 32'h4263c889, 32'h4285c33f};
test_weights[31960:31967] = '{32'h42c57888, 32'h4214e166, 32'h4295eadf, 32'h42897e23, 32'h425ef4d2, 32'h4181d485, 32'h41eebbfb, 32'h42085aad};
test_bias[3995:3995] = '{32'h4222971e};
test_output[3995:3995] = '{32'h44b4b669};
test_input[31968:31975] = '{32'h41697528, 32'hc29bd8d5, 32'hc20f3ac3, 32'h42b7ca0e, 32'h426abfb3, 32'h41847626, 32'hc21e841c, 32'h425ff605};
test_weights[31968:31975] = '{32'hc2b14776, 32'hc2242008, 32'h42a7056d, 32'hc1718fba, 32'h424c6848, 32'hc28f2f15, 32'h428461a8, 32'h42ba825c};
test_bias[3996:3996] = '{32'hc2886b31};
test_output[3996:3996] = '{32'h44e9bec6};
test_input[31976:31983] = '{32'h42169c1b, 32'hc263cd07, 32'hc21be780, 32'hc1c0a1f7, 32'hbf263c2f, 32'hc20ad184, 32'hc2aa76a2, 32'hc2662271};
test_weights[31976:31983] = '{32'hc256b810, 32'h41f4fdf5, 32'h42682b58, 32'hc2a78cae, 32'h41baa857, 32'h42aab5ba, 32'hc10f0514, 32'hc0b05ea9};
test_bias[3997:3997] = '{32'hc2c2452a};
test_output[3997:3997] = '{32'hc5bbae55};
test_input[31984:31991] = '{32'h4216b857, 32'hc2bc6df3, 32'hc2ad73da, 32'h42840869, 32'h42a7b845, 32'hc222a6a8, 32'h428f8e01, 32'hc256c278};
test_weights[31984:31991] = '{32'h410d7318, 32'h42077079, 32'h4282b8e3, 32'h426310fa, 32'h428a41cf, 32'hc19b6ff6, 32'h4236edac, 32'h429a7607};
test_bias[3998:3998] = '{32'hc2215767};
test_output[3998:3998] = '{32'h446238eb};
test_input[31992:31999] = '{32'hc1b0afc9, 32'h42608e90, 32'hc03612c5, 32'h4283d7b8, 32'hc26d644e, 32'h42840be7, 32'h4269ce75, 32'hc24d7922};
test_weights[31992:31999] = '{32'h40fa5571, 32'hc26564be, 32'h408b02d7, 32'hc1652d3e, 32'h3f9464f5, 32'hc2b3345f, 32'hc2bb8385, 32'h415603f2};
test_bias[3999:3999] = '{32'h42b863bb};
test_output[3999:3999] = '{32'hc6803148};
test_input[32000:32007] = '{32'h428690ed, 32'h41fb9609, 32'hc2b9e8e1, 32'hc1953418, 32'hc2bf385c, 32'h42b0dd03, 32'h41f0673b, 32'h4290af12};
test_weights[32000:32007] = '{32'hc20aa28d, 32'hc2983c5a, 32'hc1ec4861, 32'h42c6b3fe, 32'h4212ddfb, 32'hc18a6391, 32'hc295845b, 32'hc2aadeba};
test_bias[4000:4000] = '{32'hc2403d5a};
test_output[4000:4000] = '{32'hc6878926};
test_input[32008:32015] = '{32'hc27ca76a, 32'h41d9d06e, 32'hc237396c, 32'h41d2012f, 32'hc20790cb, 32'hc1eebca2, 32'hbf2c3432, 32'hc2c7a699};
test_weights[32008:32015] = '{32'h421482cc, 32'h3f9b77f6, 32'h425152c3, 32'h40ebcc29, 32'h41d97d7d, 32'h41ed7b92, 32'h40d82a1d, 32'hc235ba48};
test_bias[4001:4001] = '{32'hc1ac6a6b};
test_output[4001:4001] = '{32'hc4e2b8d7};
test_input[32016:32023] = '{32'hc2389bad, 32'hbfbe454a, 32'h42227ebe, 32'hc04275a3, 32'hc29146f7, 32'h42b5ea73, 32'hc19dd7c6, 32'hc1b7c1c4};
test_weights[32016:32023] = '{32'h42c2c584, 32'h416c67d5, 32'h4211dd7f, 32'hc28874ec, 32'hc14cb67f, 32'h426c39f4, 32'hc2c48ee6, 32'h42b5e2e4};
test_bias[4002:4002] = '{32'h427059b0};
test_output[4002:4002] = '{32'h4553779b};
test_input[32024:32031] = '{32'hc1b54082, 32'hc28a9276, 32'hc20dfbc4, 32'hc211a94b, 32'hc22c03f3, 32'h4206720b, 32'h428d24d6, 32'h41ad5ef3};
test_weights[32024:32031] = '{32'hc1304414, 32'h42236888, 32'h42a52797, 32'h4269097b, 32'h42baf8b9, 32'hc2a4ca95, 32'h4216dc73, 32'h3f8bd1f4};
test_bias[4003:4003] = '{32'h42b75003};
test_output[4003:4003] = '{32'hc635f91b};
test_input[32032:32039] = '{32'h423d94e8, 32'h42ab9f0f, 32'hc2accc42, 32'hc18745d5, 32'hbfad4161, 32'hc249fddb, 32'h41eb4f9e, 32'h406ab9ed};
test_weights[32032:32039] = '{32'h41fbcfc6, 32'h42af1fe8, 32'hc19c27a2, 32'h42a88dc0, 32'hc297b8a9, 32'h429cf859, 32'hc1c6cb3c, 32'h424a63b1};
test_bias[4004:4004] = '{32'h41bf0aa5};
test_output[4004:4004] = '{32'h4598a752};
test_input[32040:32047] = '{32'h419237ae, 32'h42ab67de, 32'hc2b9d768, 32'hbfe81132, 32'hc20eec3c, 32'h40bce454, 32'h42a94113, 32'h426cca6a};
test_weights[32040:32047] = '{32'h3fff4f65, 32'h42c0c1fb, 32'hc268eb59, 32'h40ba6b1f, 32'hc10220cd, 32'hc2c0f19a, 32'hc294e793, 32'h415d8656};
test_bias[4005:4005] = '{32'hc2488c79};
test_output[4005:4005] = '{32'h45f67430};
test_input[32048:32055] = '{32'h42a4e7de, 32'hc2c30609, 32'h428c631f, 32'h4183d77a, 32'hc1b94cd7, 32'h4237474c, 32'hc2bf8816, 32'hc29753d8};
test_weights[32048:32055] = '{32'hc20315f9, 32'h42088e2e, 32'h420e66c3, 32'hc2ab98c7, 32'h401a55ed, 32'hc0c34965, 32'h42a5e379, 32'hc2c0ea28};
test_bias[4006:4006] = '{32'hc213ad88};
test_output[4006:4006] = '{32'hc5ba5b32};
test_input[32056:32063] = '{32'hc0ea4f4d, 32'h427a5241, 32'hc292c5e4, 32'h42aaf2d3, 32'h42ad6cd8, 32'h42958742, 32'hc257f354, 32'h4210d6d6};
test_weights[32056:32063] = '{32'h429ee005, 32'h41b9804f, 32'h4127d784, 32'h42ba0ce2, 32'hc1d1e446, 32'h42006f72, 32'h42a62938, 32'h41767e7e};
test_bias[4007:4007] = '{32'hc1dbdfc1};
test_output[4007:4007] = '{32'h4583ebac};
test_input[32064:32071] = '{32'h427f83ae, 32'hc20e8f23, 32'hc1ac3c7f, 32'hc182c7a2, 32'hc2aa3917, 32'h41995053, 32'hc1b70df0, 32'h42a3a735};
test_weights[32064:32071] = '{32'h4282e0cb, 32'hc2be0a0b, 32'hc2b0f8d0, 32'h42022a6d, 32'h420ad4bb, 32'hc1d48fa9, 32'hc2bb5679, 32'hc23c1e9e};
test_bias[4008:4008] = '{32'hc2a07168};
test_output[4008:4008] = '{32'h4566b4be};
test_input[32072:32079] = '{32'h4296710b, 32'h42a78bef, 32'hc292ed70, 32'h4223bac3, 32'h41b6133c, 32'hc25ef76f, 32'h4111e335, 32'hc1a1d6a4};
test_weights[32072:32079] = '{32'hc26d90a4, 32'h4271b212, 32'h410f7927, 32'h41e29be2, 32'h4247b496, 32'h429e20d1, 32'hc2967061, 32'hc2b0ca0a};
test_bias[4009:4009] = '{32'hc1eee46c};
test_output[4009:4009] = '{32'hc489e708};
test_input[32080:32087] = '{32'h41f09ca2, 32'hbfb91840, 32'h4282c136, 32'hc12528ed, 32'h429cab38, 32'h42953b3c, 32'h427e7bd7, 32'h41f65b93};
test_weights[32080:32087] = '{32'hc2a1ece4, 32'hc1f0c153, 32'hc232471f, 32'h41db0fca, 32'h4238ac82, 32'h41dad8a1, 32'hc22f6cf3, 32'hc2b02984};
test_bias[4010:4010] = '{32'hc2b15fac};
test_output[4010:4010] = '{32'hc5ac8ccd};
test_input[32088:32095] = '{32'hc25794c8, 32'h4228e637, 32'hc0d632a1, 32'hc0e6d597, 32'h422cc0ba, 32'hc1c98076, 32'hc2200bb0, 32'hc25f75ac};
test_weights[32088:32095] = '{32'hc172ed53, 32'h42c38012, 32'hc28ec269, 32'hc238d394, 32'hc200680f, 32'hc271c984, 32'h403b6c69, 32'hc159972b};
test_bias[4011:4011] = '{32'h419e88a8};
test_output[4011:4011] = '{32'h45ccdadd};
test_input[32096:32103] = '{32'h4298b6da, 32'h4245dab8, 32'h42ab75c1, 32'hc29d7e24, 32'hc2c36bc6, 32'hc255f3f9, 32'h41489711, 32'h423ae086};
test_weights[32096:32103] = '{32'hc2bf9c7b, 32'hc277de6a, 32'h42114dc7, 32'h42a9d40c, 32'h424d5465, 32'h41869954, 32'h4224ffff, 32'hc2b51b36};
test_bias[4012:4012] = '{32'hc2b4d588};
test_output[4012:4012] = '{32'hc6b8f108};
test_input[32104:32111] = '{32'hc2b6fecd, 32'h429427ac, 32'hc21ee820, 32'hc0ecbe79, 32'h4107b684, 32'h4230543c, 32'hc2027461, 32'h429b0dd5};
test_weights[32104:32111] = '{32'hc257bee8, 32'h428e4baf, 32'h41a71342, 32'hc10612ef, 32'hc2af2f48, 32'hc2165127, 32'hc2b39d69, 32'h423faf66};
test_bias[4013:4013] = '{32'hc2acbcb4};
test_output[4013:4013] = '{32'h46547045};
test_input[32112:32119] = '{32'hc282039d, 32'h428e894d, 32'h419d7df6, 32'h423ef248, 32'h426043a1, 32'hc27f5aac, 32'h426aa96f, 32'h42398844};
test_weights[32112:32119] = '{32'hc0c1f336, 32'h40ee3614, 32'h423a2c21, 32'h42bd3bdc, 32'hc24a6940, 32'h42423aab, 32'h42b75daf, 32'hc2a07142};
test_bias[4014:4014] = '{32'h42b3a249};
test_output[4014:4014] = '{32'h450781a5};
test_input[32120:32127] = '{32'hbff0eb6a, 32'hc250dfeb, 32'h42b9d35f, 32'hc25fae9f, 32'hc2700cf8, 32'h42991795, 32'h40e0f8e2, 32'hc2be1ea9};
test_weights[32120:32127] = '{32'hc246a553, 32'hc23f8949, 32'h4035dd76, 32'hc29762b6, 32'hc1e4979a, 32'hc1fbab55, 32'h4291f957, 32'h429aa92d};
test_bias[4015:4015] = '{32'h427caaa9};
test_output[4015:4015] = '{32'hc3bc9ec9};
test_input[32128:32135] = '{32'h422e6845, 32'h4079a714, 32'hc2397003, 32'hc11a18e3, 32'h404fd744, 32'h4285236d, 32'h428aacb0, 32'hc2329241};
test_weights[32128:32135] = '{32'hc2431858, 32'h4295e1f2, 32'h42c68d09, 32'h41e6f7ee, 32'h429844bb, 32'hc2b26d6c, 32'h42a976fb, 32'h41c5464c};
test_bias[4016:4016] = '{32'hc297ade9};
test_output[4016:4016] = '{32'hc5f0df6c};
test_input[32136:32143] = '{32'hc2109e81, 32'h41e7dd56, 32'hc208c842, 32'h41d0f1c6, 32'h42ab1496, 32'hc12ad87d, 32'hc2156da1, 32'hc2a77ace};
test_weights[32136:32143] = '{32'hc2866376, 32'h428669b3, 32'hc29d26fe, 32'h41b46048, 32'h420e61b7, 32'hc27336d7, 32'h42a76bb4, 32'hc27e218b};
test_bias[4017:4017] = '{32'hc282ab03};
test_output[4017:4017] = '{32'h46528b91};
test_input[32144:32151] = '{32'hc28d6886, 32'h42bcde36, 32'hc2a0c231, 32'hc2254e7e, 32'h409e7da2, 32'hc29c7b1d, 32'hc2ab956f, 32'hc1592775};
test_weights[32144:32151] = '{32'h42aa33aa, 32'hc294e678, 32'hc137d90e, 32'h41efe6ba, 32'h42b8835d, 32'hc1c082df, 32'hc243330a, 32'h4272288d};
test_bias[4018:4018] = '{32'hc2bcdf81};
test_output[4018:4018] = '{32'hc5f2487a};
test_input[32152:32159] = '{32'h4204203e, 32'h427f046f, 32'h4283997f, 32'hc0bf0de2, 32'h41bdbd18, 32'h42a26c26, 32'h3fd4efe7, 32'h40c8c5b2};
test_weights[32152:32159] = '{32'h422b0ed7, 32'hc1ab8064, 32'h42234648, 32'hc22c241d, 32'h42959bfe, 32'hc27c39b4, 32'hc12a3085, 32'h41a631cf};
test_bias[4019:4019] = '{32'h412442dd};
test_output[4019:4019] = '{32'hc36b2d75};
test_input[32160:32167] = '{32'h428cb6c9, 32'hc2078b05, 32'hc22a4cfe, 32'h4287f643, 32'h4241479b, 32'h42933d61, 32'hc282983a, 32'h4128431b};
test_weights[32160:32167] = '{32'h40dcb07a, 32'hc259d0b6, 32'h4118f610, 32'h42a69c68, 32'h42992e7d, 32'h42bba6dd, 32'hc2b274d4, 32'h4296d6b9};
test_bias[4020:4020] = '{32'h4203f1e9};
test_output[4020:4020] = '{32'h46c21eca};
test_input[32168:32175] = '{32'h42c1ed0a, 32'h42a9f910, 32'hc2067e2d, 32'h4293e432, 32'h41e8d634, 32'hc2b33e10, 32'hc1bd4894, 32'hc24844b2};
test_weights[32168:32175] = '{32'hc2a3b65e, 32'h424a035a, 32'hc2623e84, 32'h421772fe, 32'hc1378cd6, 32'hc22781da, 32'hc2ab2e01, 32'h429e50ff};
test_bias[4021:4021] = '{32'hc202de94};
test_output[4021:4021] = '{32'h451c8ea6};
test_input[32176:32183] = '{32'hc29fee5c, 32'hbf0a6fcd, 32'hc2a11972, 32'h42c5499b, 32'hc182b91d, 32'h410005ee, 32'hc28e7bf6, 32'h40cd7fbd};
test_weights[32176:32183] = '{32'h42902ddd, 32'hc2abdd74, 32'h42c7f729, 32'h42bff959, 32'h4290a382, 32'hbc4776a2, 32'h421afb3e, 32'hc1c770c4};
test_bias[4022:4022] = '{32'hc1e49b90};
test_output[4022:4022] = '{32'hc603c847};
test_input[32184:32191] = '{32'hc2842502, 32'hc2153c50, 32'hc298df29, 32'hc2c249cb, 32'h429e8f36, 32'hc12ffab2, 32'h42a5ad7b, 32'hc252a405};
test_weights[32184:32191] = '{32'hc0f68809, 32'h424d0cbf, 32'h42b7a77d, 32'hc2411444, 32'hc28e234e, 32'h4280ddd6, 32'hc241683b, 32'h429c0b91};
test_bias[4023:4023] = '{32'h4186dc92};
test_output[4023:4023] = '{32'hc68dfb08};
test_input[32192:32199] = '{32'hc22e8032, 32'h418e367c, 32'hc2b76763, 32'hc2112f1a, 32'hc1540b06, 32'hbf3aac40, 32'h41df67c0, 32'h4274d9e8};
test_weights[32192:32199] = '{32'h41642f8b, 32'hc17064c2, 32'hc209a2db, 32'hc0a12c7c, 32'h420e7701, 32'h42c1187c, 32'hc028e313, 32'hc1afb714};
test_bias[4024:4024] = '{32'hc22f190d};
test_output[4024:4024] = '{32'h43de46e6};
test_input[32200:32207] = '{32'hc2c3107f, 32'h425a0d85, 32'h41a74b99, 32'hc22ee9a9, 32'h410911ee, 32'h4015f1fa, 32'hc262262a, 32'h420cd01f};
test_weights[32200:32207] = '{32'hc158c176, 32'hc22b2187, 32'h41a6e426, 32'h42b6e923, 32'hc1a2df35, 32'h428922b3, 32'h42a92b3b, 32'hc2b0b817};
test_bias[4025:4025] = '{32'h4224198a};
test_output[4025:4025] = '{32'hc6425d42};
test_input[32208:32215] = '{32'h3ff4f0f7, 32'hc205cd6c, 32'hc2bd4a1d, 32'hc2b1392a, 32'hc23ad1e2, 32'hc2037646, 32'hc234c257, 32'h4190bd93};
test_weights[32208:32215] = '{32'h42bda920, 32'hc2babec0, 32'h41bb363f, 32'h42a08dde, 32'hc2a8d1e3, 32'h4279eb8b, 32'hc1119a9b, 32'hc20ffc7b};
test_bias[4026:4026] = '{32'h42bfa935};
test_output[4026:4026] = '{32'hc585b605};
test_input[32216:32223] = '{32'h42a7d6b7, 32'h42ab0226, 32'hc238d6bf, 32'hc2a827f3, 32'h428d522f, 32'h4226038a, 32'hc243b215, 32'hc2c2bc76};
test_weights[32216:32223] = '{32'hc11d7f26, 32'h421f35d5, 32'h4232f8f1, 32'h422f7637, 32'h42c3dbb8, 32'hc29de90a, 32'hc0f9ea6a, 32'h41f0214a};
test_bias[4027:4027] = '{32'hc24fa767};
test_output[4027:4027] = '{32'hc505019f};
test_input[32224:32231] = '{32'h42b96a2c, 32'h428d18b9, 32'hc2879494, 32'h42a42b58, 32'hc28ae33c, 32'h429200f8, 32'h40f6b79a, 32'h42ae49d1};
test_weights[32224:32231] = '{32'hc2baf2ba, 32'h421d6445, 32'h42a4a66c, 32'hc2574c81, 32'h423617db, 32'hc18fdbce, 32'h41b887a1, 32'h414ceb90};
test_bias[4028:4028] = '{32'hc2bba5b4};
test_output[4028:4028] = '{32'hc695b586};
test_input[32232:32239] = '{32'hc28d3087, 32'h41f3548d, 32'h42c1c70c, 32'hc1534337, 32'h42679544, 32'hc0b4a994, 32'h42af4509, 32'hc2b5ab3c};
test_weights[32232:32239] = '{32'hc2a68199, 32'h42c181fa, 32'hc1dbb0db, 32'hc15faa09, 32'hc28365e6, 32'h42c540b8, 32'hc28eefd8, 32'h41419e4f};
test_bias[4029:4029] = '{32'h413a779d};
test_output[4029:4029] = '{32'hc5a7b962};
test_input[32240:32247] = '{32'hc236ee40, 32'hbf885edc, 32'h419420c1, 32'hc240f759, 32'hc2b4a256, 32'hc0cf2fd3, 32'hc20705a4, 32'hc2b43cdc};
test_weights[32240:32247] = '{32'h42948322, 32'h42802e7c, 32'h42238aae, 32'hc2a7367b, 32'h41fc8bd3, 32'h424fac43, 32'h41fcfba4, 32'h4227c709};
test_bias[4030:4030] = '{32'h42394368};
test_output[4030:4030] = '{32'hc5d0324d};
test_input[32248:32255] = '{32'h42836964, 32'h41fc5df0, 32'h428cb33c, 32'hc0da044d, 32'hc2adbbbc, 32'h4299faaf, 32'h3f28f605, 32'h40b426d3};
test_weights[32248:32255] = '{32'h42a17b7a, 32'hc2026a88, 32'hc0b6d9b4, 32'h42b87239, 32'hc256f8b1, 32'hc22fe205, 32'hc211c3cc, 32'hc2215d55};
test_bias[4031:4031] = '{32'hc198d1a2};
test_output[4031:4031] = '{32'h45851a01};
test_input[32256:32263] = '{32'h41e51291, 32'h40925907, 32'hc28d54ca, 32'hc242b07c, 32'h42c4a84b, 32'hc2027ce4, 32'h42783453, 32'hc2a86990};
test_weights[32256:32263] = '{32'h4236b3ad, 32'hc23e5667, 32'h41a78d8f, 32'hc1eaf399, 32'h4280ef74, 32'hc26303a8, 32'h429c52f1, 32'h42af7bff};
test_bias[4032:4032] = '{32'hc2a69f43};
test_output[4032:4032] = '{32'h45ce8345};
test_input[32264:32271] = '{32'h41bc4eab, 32'h42bfc8e3, 32'hc28d6a35, 32'hbd38d31a, 32'h4255a4a2, 32'h4292d223, 32'hc203522c, 32'h427a4cca};
test_weights[32264:32271] = '{32'hc2aed539, 32'hc209330d, 32'h41fbabed, 32'hc1c069c7, 32'h41ce69c9, 32'h4254825c, 32'hc2c3049a, 32'hc02a28c3};
test_bias[4033:4033] = '{32'h41e5c4e7};
test_output[4033:4033] = '{32'h4440ef9d};
test_input[32272:32279] = '{32'h41c06a94, 32'hc21093f8, 32'hc18d45d0, 32'hc2b98d88, 32'hc2904ae9, 32'hc23ee12f, 32'hc1b395d9, 32'hc25addf1};
test_weights[32272:32279] = '{32'h42352748, 32'h42c60415, 32'h428f2132, 32'h4231a6df, 32'h41183763, 32'hc23735a7, 32'h422776c8, 32'hc2ac8d42};
test_bias[4034:4034] = '{32'h4289789f};
test_output[4034:4034] = '{32'hc51dc95a};
test_input[32280:32287] = '{32'hc1907855, 32'hc2659464, 32'h41426c8c, 32'h419183f3, 32'hc2b9b862, 32'hc2891632, 32'h42a0542d, 32'hc17a4667};
test_weights[32280:32287] = '{32'h3fdaab58, 32'h429ae498, 32'hc25d4645, 32'hc1d798ef, 32'hc2005ce3, 32'hc27572e8, 32'h42616fc4, 32'h41670752};
test_bias[4035:4035] = '{32'hc238457b};
test_output[4035:4035] = '{32'h45b50d96};
test_input[32288:32295] = '{32'h42872e02, 32'hc2894b91, 32'h428b66eb, 32'h42307a2b, 32'hc158e8d2, 32'h419ff676, 32'h420214c3, 32'hc2c0fb1b};
test_weights[32288:32295] = '{32'hc1f2e85b, 32'hc15b6ddb, 32'hc2af06dd, 32'h4252b103, 32'h426eeec6, 32'hc1eabb1f, 32'hc09dd218, 32'h412a9a98};
test_bias[4036:4036] = '{32'h419112c9};
test_output[4036:4036] = '{32'hc5e8f23a};
test_input[32296:32303] = '{32'hc292fa23, 32'h41c63b35, 32'hc29b055e, 32'hc2a1e7d4, 32'h41ff94df, 32'hc24577a7, 32'hc2ba8c60, 32'hc27ca4fa};
test_weights[32296:32303] = '{32'hc26bb208, 32'hc1d27fa3, 32'hc26f18bf, 32'hc299a3b9, 32'hc2518e3e, 32'hc0a38467, 32'h42c4839b, 32'hc2b654ba};
test_bias[4037:4037] = '{32'h41409c58};
test_output[4037:4037] = '{32'h4617c800};
test_input[32304:32311] = '{32'h42afcabe, 32'h42c0bba9, 32'hc28ed6ea, 32'hc1a619e7, 32'h41ff204f, 32'h422e2041, 32'h401c3676, 32'h42862de9};
test_weights[32304:32311] = '{32'hc1e0bb8c, 32'h4269af50, 32'h42483963, 32'h428f9e78, 32'h41b31a28, 32'h42ab4704, 32'hc1b41cb0, 32'h423e54ae};
test_bias[4038:4038] = '{32'hc2393d37};
test_output[4038:4038] = '{32'h45afde0a};
test_input[32312:32319] = '{32'hc2854317, 32'hc20a8cb5, 32'h41ebed42, 32'hc0ee5d47, 32'hc23e9f00, 32'h41a39619, 32'hc2548a82, 32'h42292a09};
test_weights[32312:32319] = '{32'hc1e319ee, 32'h426935c3, 32'h41f6bb32, 32'h41e61551, 32'h41f1044d, 32'hc2c39d3e, 32'hc18657e5, 32'h42b28c60};
test_bias[4039:4039] = '{32'hc13d499b};
test_output[4039:4039] = '{32'h44df73ca};
test_input[32320:32327] = '{32'hc2a6564b, 32'h420a72bc, 32'hc29b7587, 32'h421b3310, 32'hc28166da, 32'hc236dd1a, 32'h428ef3ff, 32'h41a09cff};
test_weights[32320:32327] = '{32'hc2390a82, 32'hc1ad126f, 32'hc29948e4, 32'hc2a9df7c, 32'hc2836005, 32'hc189456f, 32'hc26d3065, 32'h42aae42e};
test_bias[4040:4040] = '{32'h424eb63b};
test_output[4040:4040] = '{32'h46020ed3};
test_input[32328:32335] = '{32'hc2bca9cb, 32'hc276b92c, 32'hc292704e, 32'h4211b550, 32'hc20302a9, 32'h42b169db, 32'h42980503, 32'h415649e2};
test_weights[32328:32335] = '{32'hbf104efe, 32'h40d391d5, 32'hc2035d48, 32'hc222e983, 32'hc28ddfc3, 32'h41ea2325, 32'hc231cb41, 32'h414f9d36};
test_bias[4041:4041] = '{32'hc1fedc66};
test_output[4041:4041] = '{32'h450c9585};
test_input[32336:32343] = '{32'h42bb4ca2, 32'h42a3189b, 32'h42970040, 32'hc2161c2d, 32'h41cf981c, 32'h40eca75f, 32'hc18d464e, 32'h423cedef};
test_weights[32336:32343] = '{32'h42293238, 32'hc269f6db, 32'h40b52352, 32'h421012b6, 32'h4241aac2, 32'h424cc436, 32'hc2a22b7d, 32'h40c90818};
test_bias[4042:4042] = '{32'h423ddd80};
test_output[4042:4042] = '{32'h44d1c6f3};
test_input[32344:32351] = '{32'h42c3717e, 32'hc179a041, 32'h42973fde, 32'h423810cc, 32'hc18e2fc6, 32'h429b979f, 32'h42bc16ab, 32'hc1a2feb5};
test_weights[32344:32351] = '{32'h42735112, 32'h42a34455, 32'hc19875f4, 32'h41a625c0, 32'h42bba863, 32'hc230010c, 32'h4271ab22, 32'hc2b70111};
test_bias[4043:4043] = '{32'hbf4058ea};
test_output[4043:4043] = '{32'h45cf7ec5};
test_input[32352:32359] = '{32'h4164831e, 32'hc2112870, 32'h42314884, 32'hc29e0713, 32'hc25db93a, 32'hc1f65d08, 32'h4234985f, 32'hc294688f};
test_weights[32352:32359] = '{32'h427f97aa, 32'hc2a03415, 32'hc1e9f12a, 32'hc16e2915, 32'hc24364e0, 32'h417ed9c3, 32'h42ba077e, 32'hc2733f24};
test_bias[4044:4044] = '{32'hc2b82310};
test_output[4044:4044] = '{32'h46632279};
test_input[32360:32367] = '{32'hbfc263a0, 32'h42852ab1, 32'hc2023461, 32'hc09259de, 32'hc2a2de52, 32'hc120046f, 32'hc296302f, 32'hc2800b11};
test_weights[32360:32367] = '{32'hc281538b, 32'h41a7fd82, 32'h42be364b, 32'hc2a88067, 32'hc29a8d67, 32'hc25b4dff, 32'hc222daba, 32'h4259dc0a};
test_bias[4045:4045] = '{32'h40177b61};
test_output[4045:4045] = '{32'h45a27f51};
test_input[32368:32375] = '{32'hc23f230c, 32'hc1f9edee, 32'hc27b381f, 32'h428f2482, 32'hc2c7e9ea, 32'h425fe996, 32'hc1cabbc6, 32'hc2b30580};
test_weights[32368:32375] = '{32'h40e4e77d, 32'hc296a31d, 32'hc2a9ff48, 32'h41d76a4d, 32'hc1fb82b2, 32'h42600f08, 32'hc054bab1, 32'h407b7c73};
test_bias[4046:4046] = '{32'hc2296885};
test_output[4046:4046] = '{32'h466e340f};
test_input[32376:32383] = '{32'h42a54b76, 32'h41895f35, 32'hc18a779f, 32'h429d98ed, 32'h41e12209, 32'h4228aa19, 32'h421b2897, 32'h421fd4e7};
test_weights[32376:32383] = '{32'h411fc860, 32'hc29239b8, 32'h41b1f756, 32'hc28f3295, 32'hc293b691, 32'h421151fb, 32'hc28a8e69, 32'h4276e99c};
test_bias[4047:4047] = '{32'hc18d912b};
test_output[4047:4047] = '{32'hc5e2502b};
test_input[32384:32391] = '{32'hc21f6a0b, 32'h42be027e, 32'hc1e37b5a, 32'h42747a13, 32'h41f670a7, 32'h4222df57, 32'h429159e6, 32'h42a79abf};
test_weights[32384:32391] = '{32'hc25d05c0, 32'h41dd018f, 32'hc22bdb60, 32'h4175d610, 32'hc2732e01, 32'h41bd402e, 32'h41ff52cf, 32'hc03d6fb0};
test_bias[4048:4048] = '{32'hc29efb91};
test_output[4048:4048] = '{32'h45fc2f09};
test_input[32392:32399] = '{32'h423a691b, 32'h424378b0, 32'hc2ba5131, 32'h41a3f3c8, 32'hc184143d, 32'h4268801b, 32'h4134ddf9, 32'h412137d4};
test_weights[32392:32399] = '{32'hc24aba8b, 32'hc2c68b9a, 32'hc0ee5089, 32'hc221ddc3, 32'hc21280bf, 32'hc29a9c0f, 32'hc2c0e568, 32'h422de9b5};
test_bias[4049:4049] = '{32'h42bd1079};
test_output[4049:4049] = '{32'hc6384c0c};
test_input[32400:32407] = '{32'h426a5552, 32'h4184c239, 32'hc24f588d, 32'hc22e8b89, 32'hc2a16ef1, 32'h421e5b90, 32'h41dd4d55, 32'h4203fd2a};
test_weights[32400:32407] = '{32'hc291beb0, 32'hc1171b83, 32'hc27f7706, 32'h42136bec, 32'hc1bcb40b, 32'hc046cd33, 32'hc1fbfba9, 32'hc1fd104a};
test_bias[4050:4050] = '{32'h4244c2ae};
test_output[4050:4050] = '{32'hc52f86e7};
test_input[32408:32415] = '{32'h425fb76f, 32'hc1a6ae28, 32'hc1782f7c, 32'hc2afba60, 32'h424fe536, 32'hc2ab4035, 32'h42b39776, 32'h42977f6e};
test_weights[32408:32415] = '{32'hc22f9825, 32'h42677e11, 32'h4200a62c, 32'h40c34078, 32'hc2c01ba1, 32'hc0e9cb5f, 32'hc10f3f52, 32'h403585af};
test_bias[4051:4051] = '{32'hc221715c};
test_output[4051:4051] = '{32'hc61770a4};
test_input[32416:32423] = '{32'h41d4e6c9, 32'hc2b638b8, 32'hc2542ac0, 32'h41b39b29, 32'h42368a4b, 32'h42aed2a1, 32'h40318ed1, 32'hc028c549};
test_weights[32416:32423] = '{32'h42b6bda9, 32'hc26729c8, 32'hc1516f5c, 32'hc26ea3dd, 32'h419f2ccc, 32'h4245f0d0, 32'h41256be5, 32'h427d5bb5};
test_bias[4052:4052] = '{32'h3f9d12ad};
test_output[4052:4052] = '{32'h463dd13c};
test_input[32424:32431] = '{32'hc25469f1, 32'hc27a53f2, 32'h4294cb10, 32'hc224cec8, 32'hc2aa5e53, 32'hc26e9635, 32'h428eaa6e, 32'h421fad22};
test_weights[32424:32431] = '{32'h41202cd2, 32'hc250b70f, 32'hc0a4ac9b, 32'h4258af40, 32'h4243d657, 32'h428636b5, 32'hc21b09e9, 32'h42c3f984};
test_bias[4053:4053] = '{32'h42ad64f8};
test_output[4053:4053] = '{32'hc5d52680};
test_input[32432:32439] = '{32'h42c02401, 32'h40214140, 32'hc24866b7, 32'hc15ea858, 32'h42af69f3, 32'hc2780761, 32'hc2ad7036, 32'hc2437a0c};
test_weights[32432:32439] = '{32'h4272a47c, 32'hc22fb1b0, 32'h42c4776d, 32'hc2657b05, 32'h424eff33, 32'hc242661c, 32'h426233aa, 32'h4207cadd};
test_bias[4054:4054] = '{32'hc2b346f2};
test_output[4054:4054] = '{32'h451bd80c};
test_input[32440:32447] = '{32'hc198101b, 32'hc2a5c346, 32'h4220a9a8, 32'hc1a2e6f4, 32'hc2b8d1ae, 32'hbf97184c, 32'hc2c59a85, 32'h41e36e95};
test_weights[32440:32447] = '{32'h42c7836b, 32'h421a63d7, 32'hc13271ae, 32'h420df45c, 32'h4250798e, 32'hc115f1dc, 32'hc1ebe163, 32'h4229ee1b};
test_bias[4055:4055] = '{32'h4241f785};
test_output[4055:4055] = '{32'hc5d7aca4};
test_input[32448:32455] = '{32'hc2408c29, 32'h4225545f, 32'hc29919a8, 32'h42953969, 32'h4251f25a, 32'h4288a689, 32'hc2300864, 32'h428b073c};
test_weights[32448:32455] = '{32'hc2c0debf, 32'h4289c4b3, 32'hc25d5d29, 32'h42959f36, 32'hc20c41eb, 32'hc20f3a29, 32'hc24bad71, 32'h41d83723};
test_bias[4056:4056] = '{32'hc223209f};
test_output[4056:4056] = '{32'h468596a1};
test_input[32456:32463] = '{32'h40f785c9, 32'hc1c1805b, 32'h420b6292, 32'hc28e785c, 32'hc238cc23, 32'h42802d0f, 32'h406011a4, 32'h40cfbd0c};
test_weights[32456:32463] = '{32'h41a0d19b, 32'h4200f8f9, 32'h41947281, 32'hc14afc82, 32'hc2aba529, 32'h419e9624, 32'h41c919f1, 32'hc28a7ce0};
test_bias[4057:4057] = '{32'hc1c8f7ee};
test_output[4057:4057] = '{32'h45b47595};
test_input[32464:32471] = '{32'h42c6dff1, 32'h42a88602, 32'hc26e7ede, 32'h420afb5f, 32'h42c1a4af, 32'h42979161, 32'hc2b1d321, 32'hc244fef7};
test_weights[32464:32471] = '{32'hc2b6ec1b, 32'hbdd07cb4, 32'hc2b80bc8, 32'h42004355, 32'hc279f286, 32'h4270505b, 32'hc12ddcea, 32'h42a4cf83};
test_bias[4058:4058] = '{32'h41c9af39};
test_output[4058:4058] = '{32'hc5dcd36b};
test_input[32472:32479] = '{32'hc2a2370a, 32'h420c0bae, 32'h4207c346, 32'h41b7a79b, 32'h42c659dd, 32'hc2732181, 32'hc184bc37, 32'hc2ba3980};
test_weights[32472:32479] = '{32'h42b2e32c, 32'hc29b9c10, 32'h3f826aeb, 32'h42410dc5, 32'hc26b7e32, 32'h42154c0b, 32'h4246f5e1, 32'hc289929e};
test_bias[4059:4059] = '{32'hc2567860};
test_output[4059:4059] = '{32'hc6326633};
test_input[32480:32487] = '{32'h418994b2, 32'hc246de78, 32'h429791fa, 32'hc1017bb9, 32'h42b6045c, 32'h42a23ba6, 32'hc222fb57, 32'h4112ea64};
test_weights[32480:32487] = '{32'hc18a9981, 32'h42bfe714, 32'h41171665, 32'hc27878cb, 32'hc2a2dc9c, 32'h42926c2f, 32'hc116ae5d, 32'h42a051f9};
test_bias[4060:4060] = '{32'hc202ec05};
test_output[4060:4060] = '{32'hc5845a1d};
test_input[32488:32495] = '{32'hc1f8d16a, 32'h4197b493, 32'hc2b17858, 32'hc26b71e0, 32'hc15a00fe, 32'hc243c8d6, 32'hc2bc8ba7, 32'hc2b0deae};
test_weights[32488:32495] = '{32'h4232b286, 32'hc2bd1b37, 32'h429f65ea, 32'h424a3955, 32'hc03a77af, 32'h419e2167, 32'hc264aabf, 32'hc2a7dcf6};
test_bias[4061:4061] = '{32'hc2b65863};
test_output[4061:4061] = '{32'hc4b3b31f};
test_input[32496:32503] = '{32'hc1d07731, 32'h4288b553, 32'hc1c9f009, 32'h425174b6, 32'hc2953288, 32'h42a05e87, 32'hc1b209c8, 32'h42c5b563};
test_weights[32496:32503] = '{32'h40d09867, 32'hc1c5854c, 32'hc2b4063f, 32'hc246393b, 32'hc23ce8f2, 32'h41a2cb75, 32'hc1f1e474, 32'hc2ad33eb};
test_bias[4062:4062] = '{32'h428d0774};
test_output[4062:4062] = '{32'hc597586c};
test_input[32504:32511] = '{32'hc259b12e, 32'h425c838c, 32'h419b66ed, 32'hbfb407ae, 32'hc2a6ed7d, 32'h429e7cba, 32'h427b4ca4, 32'h41e945b5};
test_weights[32504:32511] = '{32'hc2945782, 32'hc16bb603, 32'hc1c91675, 32'hc2ae44ae, 32'hc1e31fdb, 32'h42b1d0b7, 32'hc2462541, 32'h41ce7517};
test_bias[4063:4063] = '{32'h424593bd};
test_output[4063:4063] = '{32'h461bade7};
test_input[32512:32519] = '{32'hc2b26df9, 32'hc2784d0e, 32'hc2510fb2, 32'hc249d5e3, 32'h40e49042, 32'hc2c7b34b, 32'hc0d02a92, 32'hc0e4d17c};
test_weights[32512:32519] = '{32'hc0d708f2, 32'hc244cd40, 32'hc249f2d6, 32'hc29783b2, 32'hc2b847f2, 32'h42a780f9, 32'hc1343991, 32'hc18e9e33};
test_bias[4064:4064] = '{32'hc221962e};
test_output[4064:4064] = '{32'h449cd278};
test_input[32520:32527] = '{32'hc24bf427, 32'h429c8ce1, 32'hc24f2c0e, 32'hc25db769, 32'h42387c85, 32'hc2501d85, 32'h4256a032, 32'hc2161906};
test_weights[32520:32527] = '{32'hc2765658, 32'h429075cf, 32'h4290899f, 32'hc1bfdf87, 32'hc2b889b7, 32'hc28b4c81, 32'h42b2c184, 32'hc2531795};
test_bias[4065:4065] = '{32'hc2880d3e};
test_output[4065:4065] = '{32'h4642a1cd};
test_input[32528:32535] = '{32'h41f7a5ba, 32'h40d6e51a, 32'h40ccd99f, 32'hc29cef0b, 32'h425a5232, 32'hc2799546, 32'hc1e9aae3, 32'h4201895d};
test_weights[32528:32535] = '{32'h42630858, 32'hc291fad5, 32'h415bba7d, 32'h4245972b, 32'hc2c4c9b1, 32'hc1972a33, 32'h426e9feb, 32'hc28b3a47};
test_bias[4066:4066] = '{32'hc13af126};
test_output[4066:4066] = '{32'hc62784df};
test_input[32536:32543] = '{32'h429f4e41, 32'h421366b3, 32'h42719eb2, 32'hc299a433, 32'hc2b7a70d, 32'h4030dca2, 32'hc26bb504, 32'h41ad74c6};
test_weights[32536:32543] = '{32'h420c5a9d, 32'h420ed5e9, 32'hc1a2c7b1, 32'h41b5dfc0, 32'h40ed6d8f, 32'h41f9f97f, 32'h42a885a4, 32'hc2802ec2};
test_bias[4067:4067] = '{32'h4008a88d};
test_output[4067:4067] = '{32'hc5b5a3b1};
test_input[32544:32551] = '{32'h42411dab, 32'h42c619c5, 32'hc2b41311, 32'hc1bb07a9, 32'h41dc26dd, 32'hc254f7fb, 32'h42196da7, 32'h4263b6ed};
test_weights[32544:32551] = '{32'h42c79073, 32'h428549c1, 32'hc17fce71, 32'h42a989e8, 32'hc23519a0, 32'hc28a2096, 32'h407c1f5a, 32'h42af8060};
test_bias[4068:4068] = '{32'hc111bead};
test_output[4068:4068] = '{32'h469019cd};
test_input[32552:32559] = '{32'h421346b1, 32'h418f6f1a, 32'h4279b649, 32'hc2311bf0, 32'hc2b6d2c6, 32'hc2a4cff2, 32'h42869e86, 32'h410d4462};
test_weights[32552:32559] = '{32'hc2a09293, 32'hc28896ab, 32'hc283b899, 32'h428c10af, 32'hbfe88e51, 32'hc24a9933, 32'h41061949, 32'hc203b6c8};
test_bias[4069:4069] = '{32'h416e9b2d};
test_output[4069:4069] = '{32'hc5d36584};
test_input[32560:32567] = '{32'h4188b51c, 32'h4143fc56, 32'h422428df, 32'hc2b70ce8, 32'hc0a5dc5f, 32'h428640cd, 32'hc2646b64, 32'hc2586fb5};
test_weights[32560:32567] = '{32'hc280ed68, 32'h42c129d9, 32'h41a9240e, 32'hbf4a0c37, 32'h423696eb, 32'h42985dc6, 32'h4228d65c, 32'h42b355b0};
test_bias[4070:4070] = '{32'h4220b239};
test_output[4070:4070] = '{32'hc4a569c1};
test_input[32568:32575] = '{32'h41f423a1, 32'hc26f196f, 32'h41a2d8bc, 32'hc245aa1f, 32'h42b9e927, 32'hc2519c11, 32'hc0f1f765, 32'hc280ec2e};
test_weights[32568:32575] = '{32'h42a47c34, 32'hc28604d6, 32'h42965214, 32'h421c1c73, 32'h42c1f7cd, 32'h42bc1c61, 32'hc2349fbb, 32'h42654736};
test_bias[4071:4071] = '{32'hc2a2e569};
test_output[4071:4071] = '{32'h45d381b5};
test_input[32576:32583] = '{32'h425da012, 32'h41e0ae45, 32'h42985657, 32'h429588e2, 32'hc109ddff, 32'hc2907bc7, 32'h423ea909, 32'h420c57f4};
test_weights[32576:32583] = '{32'hc13ceee1, 32'h42049b54, 32'h4202c589, 32'h42552346, 32'h4017386c, 32'hc2956970, 32'hc157ce9b, 32'hc28c8b2b};
test_bias[4072:4072] = '{32'h40aced43};
test_output[4072:4072] = '{32'h460d019d};
test_input[32584:32591] = '{32'h42a19a8b, 32'hc1cc07d3, 32'hc294d6c9, 32'hc2bc11bf, 32'h424e82a5, 32'hbeda0b77, 32'hc28d81d8, 32'hc2aabad6};
test_weights[32584:32591] = '{32'h41fad55d, 32'h4256de2f, 32'h41b8864f, 32'hc2a6ca3a, 32'hc2161465, 32'h4219e2cd, 32'hc295fd67, 32'hc1f2d52c};
test_bias[4073:4073] = '{32'hc26ef1d3};
test_output[4073:4073] = '{32'h464dd484};
test_input[32592:32599] = '{32'hc22aacc5, 32'h41beaeab, 32'hc1d5437a, 32'h42bcf4ab, 32'hc22f9ed6, 32'h41ffdac9, 32'hc1ec9f63, 32'hc2aa7494};
test_weights[32592:32599] = '{32'hc0dabc2e, 32'h42857b2b, 32'h41e7b58b, 32'h42a9d8df, 32'hc2a15eab, 32'hc26f63b7, 32'hc27a75de, 32'h41a005fc};
test_bias[4074:4074] = '{32'h421e74dc};
test_output[4074:4074] = '{32'h462b1409};
test_input[32600:32607] = '{32'h4211bf1e, 32'h42b68708, 32'h426e72f2, 32'hc2731488, 32'hc2a2880f, 32'hc231ec77, 32'hc23b88ee, 32'h425b9cb2};
test_weights[32600:32607] = '{32'hc2c0d7cd, 32'hc2bb4cdf, 32'hc16963f4, 32'hc25f4d81, 32'h4089f454, 32'hc291cdc8, 32'hc0b76065, 32'hc25ae882};
test_bias[4075:4075] = '{32'h426bf3a2};
test_output[4075:4075] = '{32'hc611a727};
test_input[32608:32615] = '{32'hc1b6a7c3, 32'h425414bc, 32'hc2958297, 32'hc2344270, 32'hc100e28a, 32'h4257be3c, 32'h428abfb1, 32'hc2539456};
test_weights[32608:32615] = '{32'hc25d0c64, 32'h42417bf2, 32'hc22e6c2c, 32'h42013a34, 32'h42bf4adb, 32'h4240489e, 32'h41c8a3e5, 32'h41073cfa};
test_bias[4076:4076] = '{32'h412d49e0};
test_output[4076:4076] = '{32'h4608d0a3};
test_input[32616:32623] = '{32'hc28ecab2, 32'hc2564656, 32'h4286c819, 32'hc10df660, 32'h420e1c11, 32'h42426296, 32'hc29b4ad3, 32'h42252fb8};
test_weights[32616:32623] = '{32'h42b33dba, 32'hc116f674, 32'hc299a17b, 32'hc2887828, 32'hc2b53980, 32'hc2bef6db, 32'hc2b5275c, 32'hc20b0937};
test_bias[4077:4077] = '{32'hc1b9c6a3};
test_output[4077:4077] = '{32'hc647355e};
test_input[32624:32631] = '{32'hc222eb5d, 32'hc2aff671, 32'hc2bad7a6, 32'hc0edb219, 32'hc2811440, 32'hc21fc3b1, 32'h41e63acb, 32'hc1b0430a};
test_weights[32624:32631] = '{32'hc1186ae8, 32'hc2bcb627, 32'hc01fed1d, 32'hc2904d8a, 32'hc2813a7e, 32'h4299adf2, 32'h40ca800a, 32'hc1e30a6b};
test_bias[4078:4078] = '{32'h4161f188};
test_output[4078:4078] = '{32'h4631d644};
test_input[32632:32639] = '{32'hc2a9598b, 32'h40f621a9, 32'h421612cf, 32'h42aed9fb, 32'hc2ba66e4, 32'h42c04cc0, 32'h42bef056, 32'h410f2b40};
test_weights[32632:32639] = '{32'hc1a628ee, 32'h421d6897, 32'h4296ddb3, 32'hc2c58157, 32'h4264e968, 32'hc26383e9, 32'hc296ffc5, 32'hbf99722e};
test_bias[4079:4079] = '{32'h42363e3a};
test_output[4079:4079] = '{32'hc6a9ab5a};
test_input[32640:32647] = '{32'hc28c1b39, 32'hc2993c25, 32'h42bc5da0, 32'hc0b6d181, 32'h41d1ecb4, 32'hc22224c4, 32'h40a35bbc, 32'h426bf5fd};
test_weights[32640:32647] = '{32'h42c46a9b, 32'hc2a98a32, 32'h429e8165, 32'hc22364b3, 32'h417dffbf, 32'h407bdb64, 32'hc1bde8f0, 32'hc2304e99};
test_bias[4080:4080] = '{32'hc15bb45c};
test_output[4080:4080] = '{32'h459715af};
test_input[32648:32655] = '{32'hc202e4f3, 32'hc2bbb48c, 32'h42bad5ac, 32'hc21a688c, 32'h41fb7300, 32'hc23fa0fd, 32'h4236970d, 32'h40daf225};
test_weights[32648:32655] = '{32'h42a00851, 32'hc28a0e01, 32'h41a41054, 32'h41fa2837, 32'hc259e641, 32'hc29bad2d, 32'hc26cc556, 32'hc2708021};
test_bias[4081:4081] = '{32'h42202cc5};
test_output[4081:4081] = '{32'h455b82d3};
test_input[32656:32663] = '{32'h41a41114, 32'h418d4828, 32'hc2955294, 32'hc28f566a, 32'hc2192554, 32'hc27236c0, 32'hc241e450, 32'h4154ef01};
test_weights[32656:32663] = '{32'hc1abf2ed, 32'h41bca92e, 32'hc0c9df88, 32'hc25120d6, 32'h42b651c6, 32'hc23da68d, 32'h427b41b0, 32'hc1a329cb};
test_bias[4082:4082] = '{32'h41d97a29};
test_output[4082:4082] = '{32'h438eba88};
test_input[32664:32671] = '{32'hc27fabbf, 32'h426a8ff3, 32'hc1ada47e, 32'h42b10824, 32'h424128d7, 32'h42afa96a, 32'h42b853b2, 32'hc1edf96b};
test_weights[32664:32671] = '{32'hc2c29c17, 32'hc2b455cb, 32'h42452a31, 32'hc2610131, 32'hc29d13ac, 32'h4284f1cf, 32'hc252615c, 32'h423b9fe4};
test_bias[4083:4083] = '{32'h42afb8a6};
test_output[4083:4083] = '{32'hc610283d};
test_input[32672:32679] = '{32'hc28ca16c, 32'h41649229, 32'hc21f10f7, 32'hc19e1478, 32'hc182d8d1, 32'hc146bc1b, 32'hc2552504, 32'h408d545d};
test_weights[32672:32679] = '{32'h4112d809, 32'hc29d69f8, 32'h423b12be, 32'h4238d012, 32'h4249ab40, 32'hc050274c, 32'h424d5529, 32'h423d84ed};
test_bias[4084:4084] = '{32'h42798da0};
test_output[4084:4084] = '{32'hc5f37373};
test_input[32680:32687] = '{32'hc2170118, 32'hc282bfcb, 32'h41d1855c, 32'hc248e002, 32'h42672df2, 32'h422fe3aa, 32'h410ef712, 32'hc2a776df};
test_weights[32680:32687] = '{32'h428c253e, 32'h42a514f7, 32'h42329706, 32'h4209f3bc, 32'h426f0fb4, 32'h41b4a461, 32'h429115f6, 32'h414cc797};
test_bias[4085:4085] = '{32'h426aa511};
test_output[4085:4085] = '{32'hc58d4e64};
test_input[32688:32695] = '{32'hc2b84930, 32'h40ce0e5a, 32'hc2899382, 32'h41bb6ead, 32'hc2aca81e, 32'h4164280a, 32'hc0683760, 32'h42a687fd};
test_weights[32688:32695] = '{32'hc216c0f2, 32'hc21ff8ec, 32'hc1ae9d90, 32'h429c5052, 32'h41e51f8b, 32'h420edf56, 32'h40edc8d4, 32'h3ecf8357};
test_bias[4086:4086] = '{32'h41488dd4};
test_output[4086:4086] = '{32'h458fdf8f};
test_input[32696:32703] = '{32'h4256525c, 32'h41c0845c, 32'h42b3f6d7, 32'h4188896c, 32'h419e974b, 32'h42b7e6cc, 32'hc21a5982, 32'h42a00a80};
test_weights[32696:32703] = '{32'hc2154c22, 32'hc287b9a4, 32'h424ce692, 32'hc2496e36, 32'hc0e0d812, 32'h42b9534b, 32'hc0e3a298, 32'hc2854a18};
test_bias[4087:4087] = '{32'h42a328e4};
test_output[4087:4087] = '{32'h455c131b};
test_input[32704:32711] = '{32'h4238c8ca, 32'hc2862db6, 32'hc28c232f, 32'hc22f6381, 32'hc266e46a, 32'hc1cc4c87, 32'hc23500d8, 32'h41649cb3};
test_weights[32704:32711] = '{32'h41ecd551, 32'hc1f2d593, 32'h429a9847, 32'h428de9d9, 32'hc2b6226c, 32'h429bffb9, 32'hc2aed186, 32'hc2844cac};
test_bias[4088:4088] = '{32'hc26964e1};
test_output[4088:4088] = '{32'h4488a87b};
test_input[32712:32719] = '{32'hc271d785, 32'h41c513f9, 32'h42b8b4fc, 32'hc22c6da7, 32'h419d663e, 32'h41dd1eca, 32'hc2b8aacf, 32'hc2831a54};
test_weights[32712:32719] = '{32'hc0d929d1, 32'h41c456ef, 32'h418bcb93, 32'hc26f7f7b, 32'h428afca7, 32'hc2ba3b08, 32'h41138875, 32'h42191b9d};
test_bias[4089:4089] = '{32'h41d7d3ab};
test_output[4089:4089] = '{32'h4427724c};
test_input[32720:32727] = '{32'h427fef22, 32'h429332a5, 32'hc23ffa8b, 32'h429497c3, 32'hc27188d2, 32'h428e2a4c, 32'h40b92b64, 32'h4245d7ed};
test_weights[32720:32727] = '{32'hc291d9a6, 32'hc2902ec9, 32'hc12488ba, 32'hc0c89d63, 32'h41d4d90e, 32'hc1c7e44c, 32'hc2886c1f, 32'h423a7533};
test_bias[4090:4090] = '{32'h40d4634c};
test_output[4090:4090] = '{32'hc63244ee};
test_input[32728:32735] = '{32'hc235b3ed, 32'hc1bc50b2, 32'h420f977c, 32'hc2980ef0, 32'h423c66c3, 32'hc27f7087, 32'h429a61ec, 32'h42a50ac8};
test_weights[32728:32735] = '{32'h4225d7c2, 32'hc1db1e0a, 32'hc209a19c, 32'h42569a60, 32'h42bd4553, 32'hc2392986, 32'h41b311ba, 32'hc0d7a538};
test_bias[4091:4091] = '{32'h41382f05};
test_output[4091:4091] = '{32'h44ff7ba1};
test_input[32736:32743] = '{32'hc2174c80, 32'h41e77e56, 32'h4237d462, 32'hc2220c26, 32'hc0899a00, 32'h42ae2c8a, 32'h429cc686, 32'h4292846b};
test_weights[32736:32743] = '{32'h41144572, 32'h42199634, 32'h42a54484, 32'hc29564f5, 32'hc2a1e386, 32'h42bf5819, 32'h429862ab, 32'hc2b55cec};
test_bias[4092:4092] = '{32'hc2c6f6d4};
test_output[4092:4092] = '{32'h4672183d};
test_input[32744:32751] = '{32'h42a3f69f, 32'hc2c75077, 32'h3fa95c16, 32'hc28d2364, 32'hc24dbd7b, 32'hc228efd6, 32'hc171a7a3, 32'hc278f9f0};
test_weights[32744:32751] = '{32'hc212c231, 32'hc1ef72a3, 32'h42a73050, 32'hc2983c3d, 32'hc2bade6c, 32'hc289fd9d, 32'hc2528273, 32'h42a14445};
test_bias[4093:4093] = '{32'hc2c5b1da};
test_output[4093:4093] = '{32'h460a57c7};
test_input[32752:32759] = '{32'hc272e994, 32'hc29b00b8, 32'h404af34e, 32'hc1a2511f, 32'hc2b1ab4e, 32'hc2b3e5e2, 32'hc224b628, 32'h429aa664};
test_weights[32752:32759] = '{32'hc2581993, 32'hc1e0c77f, 32'hc13035a2, 32'hc28af0d6, 32'h42543be6, 32'h42b8a91f, 32'h42b407c9, 32'h41f36c5c};
test_bias[4094:4094] = '{32'h4185b863};
test_output[4094:4094] = '{32'hc5eb140b};
test_input[32760:32767] = '{32'h423d3c31, 32'h4248af24, 32'h42c3819e, 32'hc25357be, 32'hc21810c2, 32'hc19d1b6e, 32'hc2b16ee4, 32'h42490ccf};
test_weights[32760:32767] = '{32'h419a3e62, 32'h414731f8, 32'h4287ee96, 32'h425dbe89, 32'h40ed3e7e, 32'h4212f184, 32'h427828f5, 32'hc1b7499a};
test_bias[4095:4095] = '{32'hc1de90fe};
test_output[4095:4095] = '{32'hc518300d};
test_input[32768:32775] = '{32'h420c4fbf, 32'h42b8d9eb, 32'hc2981856, 32'h42917b00, 32'h42274bb8, 32'hc1c8b21d, 32'hc21ad288, 32'hc28e93af};
test_weights[32768:32775] = '{32'hc2a1f185, 32'hc1de76ea, 32'hc1dfb654, 32'hc1869aa4, 32'hc1e17490, 32'h423cfeb1, 32'h42b42b24, 32'h426cd88b};
test_bias[4096:4096] = '{32'h427d58ad};
test_output[4096:4096] = '{32'hc662d146};
test_input[32776:32783] = '{32'hc28c413a, 32'hc219500b, 32'h428a398c, 32'hc2772c98, 32'hc28bdc46, 32'h4208a1f3, 32'h4289b3fe, 32'h428e5616};
test_weights[32776:32783] = '{32'hc288a3ad, 32'hc2bace64, 32'h412cd12e, 32'h429bd7bc, 32'hc1c8671e, 32'hbdc986f9, 32'h40c08233, 32'hc15b4c20};
test_bias[4097:4097] = '{32'h4217b373};
test_output[4097:4097] = '{32'h45acbce0};
test_input[32784:32791] = '{32'hc2c04807, 32'h42c37465, 32'hc2a6a0bb, 32'hc1638cb3, 32'h409cf6ad, 32'hc205271f, 32'h41f19a9a, 32'h4198142b};
test_weights[32784:32791] = '{32'hbef4aa5c, 32'h428fe31f, 32'h4137a548, 32'h3f887154, 32'h4228b82b, 32'h429bd488, 32'h41f553be, 32'h4194c343};
test_bias[4098:4098] = '{32'h428e1c02};
test_output[4098:4098] = '{32'h459e6a53};
test_input[32792:32799] = '{32'h42c1e3c0, 32'h424a4dda, 32'hc2743fb9, 32'hc21cf67f, 32'hc2969d1d, 32'h42b19276, 32'hc1720fa9, 32'h42844c72};
test_weights[32792:32799] = '{32'h41a051b1, 32'hc1b51b8b, 32'hbf3e74b5, 32'h42381387, 32'hc26e9f76, 32'hc1d16749, 32'h420aa27d, 32'h423ec664};
test_bias[4099:4099] = '{32'hc24d643b};
test_output[4099:4099] = '{32'h456c9184};
test_input[32800:32807] = '{32'h41aeee53, 32'hc2a9c1f4, 32'hc148ff7c, 32'h420381cc, 32'h415fb8cb, 32'h42b1cdeb, 32'h42a0e8b8, 32'h424d45e9};
test_weights[32800:32807] = '{32'hc113b076, 32'hc2a87bd1, 32'h423df102, 32'hc0e224f3, 32'h40588de6, 32'h41de4b9f, 32'h427b4f4a, 32'hc2816d17};
test_bias[4100:4100] = '{32'h41ab75ae};
test_output[4100:4100] = '{32'h462261f6};
test_input[32808:32815] = '{32'h41dbe253, 32'h427702c2, 32'hc287c623, 32'h42901a3c, 32'hc297bba3, 32'hc297b4ad, 32'h408bb33e, 32'hc1d734ff};
test_weights[32808:32815] = '{32'h42762442, 32'hc2bd5614, 32'hc1ec544c, 32'hc20ee644, 32'h4284e4c4, 32'hbfb7c71d, 32'hc27e973c, 32'h4245231b};
test_bias[4101:4101] = '{32'hc122550e};
test_output[4101:4101] = '{32'hc63014df};
test_input[32816:32823] = '{32'h42a0617f, 32'h4207a6f2, 32'hc1eda710, 32'h411b53c1, 32'h4236c275, 32'h414fdd96, 32'h42898611, 32'hc1f994b2};
test_weights[32816:32823] = '{32'h423c7aba, 32'hc2b39969, 32'h41b42897, 32'hc2912372, 32'hc12a1e02, 32'h41edd67f, 32'hc270556d, 32'h429bfd90};
test_bias[4102:4102] = '{32'hc2766bb6};
test_output[4102:4102] = '{32'hc5e63161};
test_input[32824:32831] = '{32'h4212f882, 32'h42bf6ed7, 32'hc2813ab5, 32'h42927a3d, 32'hc2a0b575, 32'hc283392e, 32'h4112aea8, 32'hc28c747d};
test_weights[32824:32831] = '{32'h42b02407, 32'hc2ab6197, 32'hc2825a10, 32'h42ad3e9f, 32'h42515409, 32'h4273c461, 32'h41a555c5, 32'hc2a17893};
test_bias[4103:4103] = '{32'hc297290a};
test_output[4103:4103] = '{32'h45461805};
test_input[32832:32839] = '{32'h421d2587, 32'h42c3d80c, 32'h42110d94, 32'h4111f11d, 32'h420d59a2, 32'h425b4d2a, 32'hc25457bc, 32'hc24f9971};
test_weights[32832:32839] = '{32'hc0b77ef4, 32'hc2805653, 32'h423a1f76, 32'h42a754d2, 32'h4226fe91, 32'hc28a1640, 32'h42b9c7d5, 32'hc217009a};
test_bias[4104:4104] = '{32'h42777fd4};
test_output[4104:4104] = '{32'hc610f96a};
test_input[32840:32847] = '{32'h42b0f2c9, 32'h4218fcce, 32'h40bcec0d, 32'h41adbd20, 32'h40ef851a, 32'hc138fce0, 32'h4242cd57, 32'h41e58a52};
test_weights[32840:32847] = '{32'h42914441, 32'hc266bef9, 32'hc2b4da9b, 32'h42c14074, 32'hc28c75db, 32'h4249148e, 32'hc2a34446, 32'hc1bb25f7};
test_bias[4105:4105] = '{32'hc10054d5};
test_output[4105:4105] = '{32'h41b5d41d};
test_input[32848:32855] = '{32'h42076f68, 32'h42aa8671, 32'hc299682c, 32'hc2212498, 32'hc1e860eb, 32'hc2825d8a, 32'hc1d8c0b9, 32'hc2c63a09};
test_weights[32848:32855] = '{32'h4295d585, 32'h42bfe9ab, 32'h42ae1e03, 32'hc2b5556e, 32'hc027a03c, 32'hc2243d65, 32'h42b4abd7, 32'h3ebd42c1};
test_bias[4106:4106] = '{32'h421e2740};
test_output[4106:4106] = '{32'h45fa0651};
test_input[32856:32863] = '{32'hc25ce6d5, 32'hc048ae50, 32'hc23b8973, 32'h42c1242f, 32'hc2a86741, 32'hc1740207, 32'hc2ade7ab, 32'hc0a03bba};
test_weights[32856:32863] = '{32'h42624cee, 32'h42c655ce, 32'h42a56d65, 32'h3fc1c599, 32'h3f89a341, 32'hbf15d6e0, 32'hc1978026, 32'hc2a78295};
test_bias[4107:4107] = '{32'hc288d33b};
test_output[4107:4107] = '{32'hc5a418af};
test_input[32864:32871] = '{32'hc22743b4, 32'h42911e41, 32'h42c30330, 32'hc2a4997e, 32'h4218807c, 32'h4284b8fc, 32'hc276bdd2, 32'hc2551012};
test_weights[32864:32871] = '{32'hc2be0831, 32'h40bb85ea, 32'hc226fda2, 32'hc17b8954, 32'hbfa25101, 32'hc2346fe7, 32'h41370d35, 32'hc2b18c6f};
test_bias[4108:4108] = '{32'hc2c65d83};
test_output[4108:4108] = '{32'h451c7709};
test_input[32872:32879] = '{32'h426e9ea5, 32'h424be2c4, 32'h4258e107, 32'hc1048308, 32'hc1e3f987, 32'hc2c46073, 32'h428b57fa, 32'hc2b629b3};
test_weights[32872:32879] = '{32'hc2a341df, 32'h423cc523, 32'h413f8c44, 32'hc18062c3, 32'h42465206, 32'hc2bdb421, 32'h42a5bc0d, 32'h42b432c8};
test_bias[4109:4109] = '{32'h41fbc087};
test_output[4109:4109] = '{32'h456e906e};
test_input[32880:32887] = '{32'h428b84c2, 32'h4210a03f, 32'hc23d1ea5, 32'hc249bc62, 32'h428a170f, 32'hc28943c4, 32'hc0345f98, 32'h4085b336};
test_weights[32880:32887] = '{32'hc1d9055c, 32'h4238364d, 32'h428cc14e, 32'hc2056dbc, 32'h42987ed5, 32'h424abca2, 32'hc0b2667c, 32'h425ba358};
test_bias[4110:4110] = '{32'h427db9a3};
test_output[4110:4110] = '{32'h435e1d02};
test_input[32888:32895] = '{32'h42a4db82, 32'hc22aeeba, 32'hc25eefa5, 32'h42bced8e, 32'hc2637c3a, 32'hc1a05308, 32'hc2aeb161, 32'hc284efca};
test_weights[32888:32895] = '{32'h423c3195, 32'hbf292dcf, 32'hc160e293, 32'h427e95c1, 32'hc242abf9, 32'hc22fa121, 32'hc248745e, 32'hc2b22b6f};
test_bias[4111:4111] = '{32'hc23fa90c};
test_output[4111:4111] = '{32'h46c030d1};
test_input[32896:32903] = '{32'h4180e0b3, 32'hc225311c, 32'h41ab1859, 32'h41d41588, 32'hc21c2fde, 32'hc03a41c7, 32'hc2c223b0, 32'hc1cf6264};
test_weights[32896:32903] = '{32'hc13b32d6, 32'h424d45f1, 32'hc22d944a, 32'hc260d11f, 32'h4117fecd, 32'h42c28866, 32'hc28c4a59, 32'hc2934693};
test_bias[4112:4112] = '{32'h423d748b};
test_output[4112:4112] = '{32'h45539588};
test_input[32904:32911] = '{32'hc261ee46, 32'hc1afd255, 32'hc2bbca01, 32'hc291f5e8, 32'hc2b1562f, 32'h42c0b1a7, 32'hc288e034, 32'hc29d3bd1};
test_weights[32904:32911] = '{32'hc2837699, 32'hc1fcd335, 32'hc28a715f, 32'h4291e870, 32'hc203e337, 32'hc1c6da63, 32'h428bdcb2, 32'h42c60c38};
test_bias[4113:4113] = '{32'hc2bf9067};
test_output[4113:4113] = '{32'hc5ccdb0d};
test_input[32912:32919] = '{32'h40832da4, 32'hc240d02d, 32'h3f9b30dd, 32'hc2a73e1e, 32'hc2b23f39, 32'hc2a64fea, 32'h4250587f, 32'hc2c6e818};
test_weights[32912:32919] = '{32'hc0807ea0, 32'h422c4fb1, 32'hc262f025, 32'h42c1d162, 32'hc23d96b4, 32'h427ebe72, 32'hc252a159, 32'h42529391};
test_bias[4114:4114] = '{32'h42ac47f8};
test_output[4114:4114] = '{32'hc6963a9c};
test_input[32920:32927] = '{32'hc2c0f806, 32'hc253f488, 32'h42575045, 32'hc28cda80, 32'h415f21bd, 32'hc1323629, 32'hc2b1b894, 32'hc256d883};
test_weights[32920:32927] = '{32'hc2840c25, 32'h41ae736a, 32'hc25e573e, 32'h42a00e35, 32'h42a54025, 32'hc2311b40, 32'h423d78e5, 32'hc25dc904};
test_bias[4115:4115] = '{32'h42bfe38c};
test_output[4115:4115] = '{32'hc53570f6};
test_input[32928:32935] = '{32'hc2a4a1ef, 32'hc14b52e5, 32'h42874c00, 32'h429cdab5, 32'hc12ffd45, 32'h421ccc45, 32'hc241cfa8, 32'hc2ae243c};
test_weights[32928:32935] = '{32'h42770176, 32'hc2705cd4, 32'h42b126d5, 32'h424c14b7, 32'hc29bdfd1, 32'h4283b5c6, 32'hc1f64897, 32'h42b3e2bf};
test_bias[4116:4116] = '{32'hc215201f};
test_output[4116:4116] = '{32'h452af900};
test_input[32936:32943] = '{32'h42b3a08b, 32'hc2bcde2d, 32'hc2932b87, 32'hc1e9b8af, 32'hc21879cc, 32'h426ad01d, 32'h42312eea, 32'h42471b11};
test_weights[32936:32943] = '{32'h429f3b41, 32'hc1e0c07d, 32'h4254bb21, 32'hc1c9eed4, 32'h4280a931, 32'h42af5c66, 32'hc23569be, 32'hc298e3dc};
test_bias[4117:4117] = '{32'hc1c1ead6};
test_output[4117:4117] = '{32'h4559c240};
test_input[32944:32951] = '{32'hc2900886, 32'h424507d1, 32'h4228cbf4, 32'hc0d18740, 32'h429192ec, 32'h42b14ce1, 32'hc2808f05, 32'hc1920f15};
test_weights[32944:32951] = '{32'h42b0be52, 32'h42baed4b, 32'hc0b7be02, 32'h426f9bf3, 32'h40a60667, 32'hc1a7a0e8, 32'h40de652f, 32'h4296d47a};
test_bias[4118:4118] = '{32'hc29c4b33};
test_output[4118:4118] = '{32'hc5b4850f};
test_input[32952:32959] = '{32'hc1ed661e, 32'h41af5bab, 32'h42c159b6, 32'hc1551e18, 32'hc20a58e3, 32'h41664c1b, 32'hc2484590, 32'h41c5420a};
test_weights[32952:32959] = '{32'h4250366c, 32'hc2c4d9f6, 32'hc284eab9, 32'h40e42215, 32'hc19d7eb1, 32'hc25d65a2, 32'h423edcac, 32'hc2c6dc60};
test_bias[4119:4119] = '{32'h4175aebb};
test_output[4119:4119] = '{32'hc66cec5e};
test_input[32960:32967] = '{32'h4294b135, 32'h42b111d0, 32'h4296a08d, 32'hc0b01fe9, 32'hc28c6b0c, 32'h425625fc, 32'hc2bc1a87, 32'h425cc3af};
test_weights[32960:32967] = '{32'hc2b2542e, 32'h42a47ebd, 32'h4214099f, 32'hc2350af7, 32'hc2a54563, 32'hc27ba90e, 32'hc14d0484, 32'h41ac58f1};
test_bias[4120:4120] = '{32'hc28943a7};
test_output[4120:4120] = '{32'h46040099};
test_input[32968:32975] = '{32'h41d2785f, 32'h4263b83f, 32'hc138c55c, 32'hc2a59b43, 32'hc273ec12, 32'hc2bb557f, 32'h41c8049e, 32'hc0746a20};
test_weights[32968:32975] = '{32'h416cef6d, 32'hc2336c97, 32'hc1664b8a, 32'hc265777f, 32'hc2094b28, 32'h418ed3df, 32'h420d84e9, 32'h423468d6};
test_bias[4121:4121] = '{32'h429ba1fd};
test_output[4121:4121] = '{32'h4577b3bd};
test_input[32976:32983] = '{32'hc15723eb, 32'hc2c0d968, 32'h42b26181, 32'h40688070, 32'hc29816d1, 32'hc18ed0b4, 32'h427015fd, 32'hc191da31};
test_weights[32976:32983] = '{32'h428cf739, 32'h41ef5efb, 32'hc259d766, 32'hc1acd52a, 32'hc0540834, 32'h4213e7ea, 32'h41e84a31, 32'h42887454};
test_bias[4122:4122] = '{32'h421d205a};
test_output[4122:4122] = '{32'hc606fac1};
test_input[32984:32991] = '{32'hc2bdefbe, 32'hc2bb79bc, 32'hc171eead, 32'h429085a3, 32'hc2a4d28f, 32'h41a7f3ca, 32'hc2aacf05, 32'hbf1c448e};
test_weights[32984:32991] = '{32'hc2c39912, 32'hc2822b74, 32'hc112ec7a, 32'h429328e9, 32'h41822463, 32'hc185d83f, 32'h41f06a17, 32'h42703b4d};
test_bias[4123:4123] = '{32'hc2552cf0};
test_output[4123:4123] = '{32'h4680e03c};
test_input[32992:32999] = '{32'hc12b85e5, 32'h4242eb6a, 32'hc26d1485, 32'h4295e3cf, 32'hc2a508f9, 32'h423efb8d, 32'hc1484bb7, 32'h42bef6ef};
test_weights[32992:32999] = '{32'h42c6fbc1, 32'hc1af94d2, 32'h421b4331, 32'h4139cdc9, 32'hc09cc1ea, 32'h419dcf5b, 32'h429e79fc, 32'h41d30193};
test_bias[4124:4124] = '{32'hbfde8219};
test_output[4124:4124] = '{32'hc42de3b7};
test_input[33000:33007] = '{32'h4253ac8e, 32'h4263de1f, 32'hc29387d0, 32'hc23085f8, 32'hc2bcb029, 32'h4043ac0a, 32'h41a6bff5, 32'hc2be888e};
test_weights[33000:33007] = '{32'h42aaf63d, 32'hc1bea487, 32'h42c0f7c9, 32'hc227afbe, 32'h41a64019, 32'hc23c0879, 32'h42b6d22b, 32'h42bc4086};
test_bias[4125:4125] = '{32'h41c43193};
test_output[4125:4125] = '{32'hc62faab4};
test_input[33008:33015] = '{32'h42a76902, 32'hc11b984f, 32'hc1ba5c11, 32'hc20ea2a9, 32'hc19ee258, 32'h40970bad, 32'hc15d1f84, 32'hc2c16589};
test_weights[33008:33015] = '{32'hc2b04a80, 32'hc22d849d, 32'h429d4009, 32'hc25ce35d, 32'h410a1699, 32'hc1c0c5b6, 32'h42a84353, 32'hc2865a1c};
test_bias[4126:4126] = '{32'hc24b3336};
test_output[4126:4126] = '{32'hc4e3b4a2};
test_input[33016:33023] = '{32'h4294a8a6, 32'hc1436bca, 32'hc1f82955, 32'hc1eb2cbb, 32'h418bdc11, 32'h427962f3, 32'hc1ba60db, 32'h428040dc};
test_weights[33016:33023] = '{32'h4264f366, 32'hc26bd9c2, 32'hc207f1c5, 32'h427c0506, 32'hc2ba7598, 32'h420c8a77, 32'hc0d61568, 32'hc26234bb};
test_bias[4127:4127] = '{32'h411ce016};
test_output[4127:4127] = '{32'h449f9320};
test_input[33024:33031] = '{32'hc2024baa, 32'hc23ee2d7, 32'h42bcba4c, 32'h42a84921, 32'h42bb649c, 32'h42a1d7b8, 32'hc2a398a2, 32'h42a74239};
test_weights[33024:33031] = '{32'hc290743b, 32'hc282ad3e, 32'h41117e87, 32'hc1cacc77, 32'h4123b76b, 32'h42b1df7c, 32'hc22d2643, 32'hc206b12d};
test_bias[4128:4128] = '{32'hc29bc6f4};
test_output[4128:4128] = '{32'h464b1941};
test_input[33032:33039] = '{32'h40785564, 32'h42be7a12, 32'hc29aaf32, 32'hc212157a, 32'hc2b7a606, 32'hc2c762a2, 32'hc2a40696, 32'h42a6dc57};
test_weights[33032:33039] = '{32'hc27b9552, 32'h413c7a3f, 32'h4129c8d0, 32'h409b7ac9, 32'hc2a96b1e, 32'hc2a81cf5, 32'hc29f43ab, 32'h42af3d28};
test_bias[4129:4129] = '{32'hc29a1cb9};
test_output[4129:4129] = '{32'h46e8d394};
test_input[33040:33047] = '{32'hc0abac36, 32'hc13c3c6d, 32'h42b8d0b8, 32'hc29466be, 32'hc279612f, 32'h42369f7b, 32'hc18304fe, 32'hc2a197d8};
test_weights[33040:33047] = '{32'h42801259, 32'h41e72aa8, 32'hc186a17f, 32'h425b358d, 32'hc28f7dff, 32'hc248055d, 32'h42a76ef1, 32'h42246680};
test_bias[4130:4130] = '{32'hc295d4bc};
test_output[4130:4130] = '{32'hc60ac6e4};
test_input[33048:33055] = '{32'hc29f6654, 32'h41b2e34b, 32'h42c1bec0, 32'hc014b40d, 32'hc1fc2067, 32'hc29609fb, 32'h426f3630, 32'h421384ed};
test_weights[33048:33055] = '{32'hc28275bf, 32'h4228c20d, 32'h42aa6327, 32'hc2966baa, 32'hc26c4ac4, 32'h42b29823, 32'h41fdb2f2, 32'h42c40f9c};
test_bias[4131:4131] = '{32'h420f535c};
test_output[4131:4131] = '{32'h466ec119};
test_input[33056:33063] = '{32'h424496b6, 32'h41330252, 32'hc1f1ade6, 32'h42c0fcee, 32'hc288fa57, 32'h41cc3c53, 32'hc1dd87b7, 32'h420ee3c6};
test_weights[33056:33063] = '{32'h41f7f065, 32'hc21413d8, 32'hc0c9026d, 32'h42a3f28e, 32'h428b0735, 32'hc2035ac2, 32'hc099ae2a, 32'h42b26c9a};
test_bias[4132:4132] = '{32'hc2947aca};
test_output[4132:4132] = '{32'h45d6389c};
test_input[33064:33071] = '{32'hc2a32340, 32'h424db317, 32'h4194dbf1, 32'h413314cf, 32'hc2c12b73, 32'h42c4ea7c, 32'h41c425c9, 32'hc1e369d2};
test_weights[33064:33071] = '{32'hc18544b6, 32'hc2bcf850, 32'h4292d7f7, 32'hc1c452a9, 32'h42c41c15, 32'hc2a8220a, 32'h4295479d, 32'hc261bf7c};
test_bias[4133:4133] = '{32'hc2ab1b23};
test_output[4133:4133] = '{32'hc6834eb6};
test_input[33072:33079] = '{32'h42068bf3, 32'hc165a711, 32'hc1911841, 32'h417bd9c8, 32'hc299f17e, 32'h41a950ea, 32'hc1f7eab4, 32'h42240448};
test_weights[33072:33079] = '{32'hc23e5d19, 32'hc284fa47, 32'h426e9b2b, 32'hc2857726, 32'hc2492345, 32'h42c6ce8c, 32'h42325552, 32'h423b29d9};
test_bias[4134:4134] = '{32'h413fe6c1};
test_output[4134:4134] = '{32'h456a085c};
test_input[33080:33087] = '{32'h405d9431, 32'h429e647a, 32'h429fd0ca, 32'hc127a7e8, 32'h42b19719, 32'hc2a082a9, 32'h4280fe6c, 32'h42a139c7};
test_weights[33080:33087] = '{32'hc21af81e, 32'h4054c954, 32'h429914de, 32'h42808d8e, 32'hc2a2dced, 32'h412d4f1c, 32'h416971fd, 32'hc26d11b1};
test_bias[4135:4135] = '{32'hc21c5242};
test_output[4135:4135] = '{32'hc5c81f5d};
test_input[33088:33095] = '{32'h42a68ded, 32'hc1e0cc3f, 32'h4208914c, 32'h42a61c2e, 32'h42c79624, 32'h42717685, 32'h41d7d838, 32'hc1a5c12c};
test_weights[33088:33095] = '{32'h42c1a8cc, 32'hc28404b8, 32'hc2a763a9, 32'h411758ed, 32'hc200bb3b, 32'h42bb40a3, 32'hc0b34e68, 32'h42b38f68};
test_bias[4136:4136] = '{32'h42a8da1a};
test_output[4136:4136] = '{32'h46029fc0};
test_input[33096:33103] = '{32'h42698f08, 32'h42ba78ee, 32'h427904c5, 32'hc18df2a1, 32'hc28a1865, 32'h424c6ac6, 32'hc250c1d1, 32'hc22cf971};
test_weights[33096:33103] = '{32'hc2314d5a, 32'h42bc0b87, 32'h4219af87, 32'hbfb5d803, 32'h42ac7422, 32'h42271427, 32'h4262214c, 32'hc1e919e0};
test_bias[4137:4137] = '{32'h4265f7b9};
test_output[4137:4137] = '{32'h454473bb};
test_input[33104:33111] = '{32'hbea129c8, 32'hc28eb1ae, 32'hc295c904, 32'hc0bfa7e7, 32'h42b32d7c, 32'h427642be, 32'hc19e2393, 32'h4213794a};
test_weights[33104:33111] = '{32'hc2c5399b, 32'h428abaea, 32'h415b3552, 32'h423a19e1, 32'h4206a536, 32'h419ca413, 32'hc2762445, 32'h42076811};
test_bias[4138:4138] = '{32'h42b1341a};
test_output[4138:4138] = '{32'h4409e104};
test_input[33112:33119] = '{32'h42adfbfa, 32'h41d16041, 32'h42bc9caf, 32'h42038171, 32'hc28e56ea, 32'h42b006d3, 32'hc23a9aae, 32'h41cca94f};
test_weights[33112:33119] = '{32'hc2c77eb1, 32'h42b2e987, 32'h4284767b, 32'hc25e1634, 32'h42c60753, 32'hc28b2917, 32'hc2730f2b, 32'hc1923293};
test_bias[4139:4139] = '{32'hc10813eb};
test_output[4139:4139] = '{32'hc646ddb2};
test_input[33120:33127] = '{32'hc2741da7, 32'hc23bd727, 32'hc2c4b56e, 32'h42a2ce44, 32'hc2a4d735, 32'h42a1e661, 32'h41d1eb1b, 32'hc177cf59};
test_weights[33120:33127] = '{32'h42c515e2, 32'h4297da82, 32'h40b01537, 32'hc2076e04, 32'h42a1d16a, 32'hc154d304, 32'hc1c46cea, 32'h429aa815};
test_bias[4140:4140] = '{32'h419bd65e};
test_output[4140:4140] = '{32'hc6af591a};
test_input[33128:33135] = '{32'h41eba40d, 32'hc1882bcd, 32'h41b94128, 32'h42849aaf, 32'hc24d7a5c, 32'hc2a918fb, 32'hc29c95a4, 32'hc1c118f5};
test_weights[33128:33135] = '{32'hc2a2a634, 32'hc268b329, 32'hc10efaba, 32'h426e2b71, 32'hc19faddc, 32'h41375df6, 32'h428f443c, 32'hc02f2514};
test_bias[4141:4141] = '{32'hc29e144e};
test_output[4141:4141] = '{32'hc549d4de};
test_input[33136:33143] = '{32'h42c34742, 32'hc1c77571, 32'hc0faa1e8, 32'hc257199c, 32'h424df7a0, 32'hc28181b2, 32'hc2a62c05, 32'hc2ab8cbc};
test_weights[33136:33143] = '{32'hc2277e12, 32'h4240a104, 32'h3f4194f7, 32'hc1e72528, 32'h426c540e, 32'h42bc2618, 32'h425d821d, 32'h423e6e87};
test_bias[4142:4142] = '{32'hc2bf72fd};
test_output[4142:4142] = '{32'hc6734c37};
test_input[33144:33151] = '{32'hc0073466, 32'hc254b4e1, 32'hc1fe9f61, 32'hc2699edd, 32'hc298152c, 32'h41eb3157, 32'h41ba68c2, 32'h421417fe};
test_weights[33144:33151] = '{32'hc2418a9d, 32'hc113fa0b, 32'h41f18678, 32'h41408b5e, 32'hc21465a9, 32'hc220a600, 32'hc2c0b5b8, 32'h41dcd115};
test_bias[4143:4143] = '{32'h423d1b32};
test_output[4143:4143] = '{32'hc41756e7};
test_input[33152:33159] = '{32'h42c68fd4, 32'h40edd810, 32'hc2006b27, 32'hc15189d5, 32'hc1223681, 32'hbf93dea3, 32'h42b0a8b3, 32'h4235b913};
test_weights[33152:33159] = '{32'h41b01184, 32'h42852271, 32'hc08c776e, 32'hc1d89f3c, 32'hc28a20c3, 32'h42bde71a, 32'hc2ac4fbb, 32'hc2829fa1};
test_bias[4144:4144] = '{32'hc231826c};
test_output[4144:4144] = '{32'hc5d63e53};
test_input[33160:33167] = '{32'h425b8068, 32'h41d399c1, 32'hc2c43c3c, 32'h421ebb67, 32'h4107b6a1, 32'h42bfa6fa, 32'h42ad0830, 32'hc285fcb9};
test_weights[33160:33167] = '{32'h4298c0b1, 32'h42598d67, 32'h4226e93b, 32'h41cb52b8, 32'h424ddaa2, 32'hc23bcde8, 32'hc23bf3fa, 32'h42528609};
test_bias[4145:4145] = '{32'hc25f0bcb};
test_output[4145:4145] = '{32'hc60f35e3};
test_input[33168:33175] = '{32'h41652eb5, 32'hc2ab07b4, 32'hc21351d7, 32'h41abe401, 32'h4256b006, 32'hc20bb488, 32'h414ccdbe, 32'h41785d5e};
test_weights[33168:33175] = '{32'h413f6a6a, 32'hc27f0295, 32'hc284419b, 32'h420a798c, 32'h42b5b8c8, 32'h422cb932, 32'hc24f0d08, 32'hc21a152e};
test_bias[4146:4146] = '{32'hc20662f4};
test_output[4146:4146] = '{32'h4629f395};
test_input[33176:33183] = '{32'h42ad6229, 32'h426d24af, 32'h3ffcdafe, 32'hc110f8d2, 32'hc2320fec, 32'hc2b72bc2, 32'h4203f6cc, 32'h4290ce12};
test_weights[33176:33183] = '{32'hc20d6357, 32'h4292ff70, 32'h42821d63, 32'hc1e619c6, 32'h42a55a48, 32'hc1b12f08, 32'h42a7c05d, 32'hc1b07128};
test_bias[4147:4147] = '{32'hc2aa99ed};
test_output[4147:4147] = '{32'h448b6a19};
test_input[33184:33191] = '{32'hc1dec844, 32'hc17760f1, 32'hc19e0ab9, 32'hc149808b, 32'h426b1697, 32'h42530226, 32'hc2aaddc6, 32'h428552f7};
test_weights[33184:33191] = '{32'h42ad46c4, 32'hc2c29dd4, 32'h4265455c, 32'h42bea99e, 32'hc20246ff, 32'hc235a3bc, 32'h428fb570, 32'hc2818d70};
test_bias[4148:4148] = '{32'h42634aef};
test_output[4148:4148] = '{32'hc68c3d8b};
test_input[33192:33199] = '{32'hc2a93fc5, 32'hc2a7ed85, 32'hc2b05b46, 32'h4282aa14, 32'hc2c4d5c9, 32'hc2608570, 32'h42c43c53, 32'h41756b15};
test_weights[33192:33199] = '{32'hc2bd1b33, 32'hc278cbda, 32'hc2abeece, 32'h420a42df, 32'hc259ee8f, 32'h41b25344, 32'h42356fed, 32'hc19d207a};
test_bias[4149:4149] = '{32'h42980a9c};
test_output[4149:4149] = '{32'h46f54d9a};
test_input[33200:33207] = '{32'h3f906209, 32'hc22864fa, 32'hc2516867, 32'h42b1d255, 32'hc2bbed26, 32'h4131c882, 32'hc2c18a93, 32'hc243a6ca};
test_weights[33200:33207] = '{32'hc2bdb5b5, 32'h427a1e53, 32'h42612666, 32'hc26a9231, 32'hc2c24618, 32'h41ab24e7, 32'h4224a5d0, 32'hc2a9e767};
test_bias[4150:4150] = '{32'h417a12b8};
test_output[4150:4150] = '{32'hc4a87113};
test_input[33208:33215] = '{32'hc1e887a0, 32'h4298c84e, 32'hc28065b5, 32'h4223e8af, 32'hc051ed9d, 32'h42bf6f50, 32'hc266479e, 32'hc239cac3};
test_weights[33208:33215] = '{32'h3fd2e2f9, 32'h427995d0, 32'hc221fb92, 32'hc29dbf4a, 32'h42bbff48, 32'h42ab011b, 32'h41d8dcc9, 32'h42bcbca8};
test_bias[4151:4151] = '{32'hc1a5e18c};
test_output[4151:4151] = '{32'h45bb6c61};
test_input[33216:33223] = '{32'h42c57e7e, 32'h4293b889, 32'h4231d87d, 32'hc2258755, 32'hc1944275, 32'h42c4e192, 32'h418b931f, 32'h4217fe7c};
test_weights[33216:33223] = '{32'hc2b1ea20, 32'h428757fd, 32'hc16b7ecd, 32'h42235934, 32'hc2bcc118, 32'hc298b863, 32'h421ab0ba, 32'hc2224ef7};
test_bias[4152:4152] = '{32'h426de517};
test_output[4152:4152] = '{32'hc64687a0};
test_input[33224:33231] = '{32'h41659c67, 32'hc280fc32, 32'h4193ce84, 32'h42bbe114, 32'h4281a87e, 32'hc2c3fe56, 32'hc2c341b2, 32'hc262d4bc};
test_weights[33224:33231] = '{32'hc1ae657e, 32'h42bb8927, 32'h42979990, 32'h425236c6, 32'h429ef623, 32'hc2920d22, 32'hc20bf932, 32'h42bbd846};
test_bias[4153:4153] = '{32'h42b2b707};
test_output[4153:4153] = '{32'h462386a5};
test_input[33232:33239] = '{32'h4299a17a, 32'hc2847605, 32'hc24eebbb, 32'h40f50c12, 32'h4270b3ac, 32'h421daef6, 32'hc2a98fbf, 32'h427e8948};
test_weights[33232:33239] = '{32'h41903cb1, 32'hc11f9aac, 32'hc2803f59, 32'hc257144d, 32'hbd2250c7, 32'hc285afd1, 32'hc1c4258b, 32'hc274e25e};
test_bias[4154:4154] = '{32'h42b88ac3};
test_output[4154:4154] = '{32'h44133326};
test_input[33240:33247] = '{32'hc2c48f18, 32'hc1e06e10, 32'hc2282371, 32'h41d1e82d, 32'hc293f1ab, 32'hc26c2a1d, 32'h42bc0390, 32'h4172f7eb};
test_weights[33240:33247] = '{32'hc20b3d2d, 32'h419d8a01, 32'hc274c16f, 32'hc19172c0, 32'h41cea3dc, 32'h42a827d3, 32'hc2ab05a3, 32'hc14fa8bb};
test_bias[4155:4155] = '{32'hc180879e};
test_output[4155:4155] = '{32'hc61ecb85};
test_input[33248:33255] = '{32'h42126afc, 32'h4265daee, 32'h4296f863, 32'hc26a3e98, 32'h427818ad, 32'hc2ba6e3a, 32'hc294ce7a, 32'h4285e043};
test_weights[33248:33255] = '{32'h427641c9, 32'hc2767dd6, 32'hc2b8eb19, 32'h424ed1ad, 32'hc2183f25, 32'hc17d4db0, 32'hc28ded6e, 32'h42296240};
test_bias[4156:4156] = '{32'hc08a54da};
test_output[4156:4156] = '{32'hc57e594a};
test_input[33256:33263] = '{32'hc2c45c1f, 32'h41c7bc26, 32'hc1aa2cfe, 32'h4243cbe5, 32'h4205785f, 32'hc107246b, 32'hc2aa3936, 32'hc151eeac};
test_weights[33256:33263] = '{32'hc21e8c76, 32'hc26d13c9, 32'hc2601ed6, 32'hc165c8e2, 32'hc1d01aaa, 32'hc2745727, 32'hc2bee0d8, 32'hc26b7cf7};
test_bias[4157:4157] = '{32'h42c30241};
test_output[4157:4157] = '{32'h4634565e};
test_input[33264:33271] = '{32'h42137351, 32'h42b74ad6, 32'hc2557e7c, 32'h41c9517c, 32'hc1616fc5, 32'hc2a3455b, 32'hc0452aa0, 32'h42323a8a};
test_weights[33264:33271] = '{32'hc204d31e, 32'hc2874ed3, 32'hc18c8463, 32'h424ac7b2, 32'hc2907657, 32'h4216fc86, 32'h4175a796, 32'hc2608560};
test_bias[4158:4158] = '{32'hc18f9647};
test_output[4158:4158] = '{32'hc619c447};
test_input[33272:33279] = '{32'h4287c16b, 32'hc1f0133b, 32'h4205336f, 32'hc1e06507, 32'hc241fdd6, 32'hc2764d6b, 32'hc21efd8a, 32'hc121012d};
test_weights[33272:33279] = '{32'h42027469, 32'hc2b4a44a, 32'hc107ed1e, 32'h42b92889, 32'hc2a8e837, 32'hc157d262, 32'h421741c8, 32'h41623e64};
test_bias[4159:4159] = '{32'h42a6c0c3};
test_output[4159:4159] = '{32'h45a90802};
test_input[33280:33287] = '{32'h4273de67, 32'h429c8cd4, 32'h41e45eba, 32'hc1da6e9f, 32'h41eadc93, 32'h420d7fc2, 32'h41c27559, 32'hc23a314e};
test_weights[33280:33287] = '{32'h42573ac0, 32'h4208add6, 32'h41afd9fe, 32'h425c1519, 32'hc1f84171, 32'hc164cf69, 32'hbfb4f138, 32'hc1c9bb39};
test_bias[4160:4160] = '{32'hc2ba14c0};
test_output[4160:4160] = '{32'h45932e5f};
test_input[33288:33295] = '{32'h42a24e07, 32'h425d5ea4, 32'h429445ae, 32'hc29ff39e, 32'hc05eb9d2, 32'h41d85bae, 32'h42c2fd42, 32'hc2bef817};
test_weights[33288:33295] = '{32'h42b3649e, 32'hc21e01b3, 32'hc2648b85, 32'hc280bd7f, 32'hc1d98ce7, 32'hc291ff52, 32'h41809d20, 32'hc23d353e};
test_bias[4161:4161] = '{32'hc1b90986};
test_output[4161:4161] = '{32'h461f29c6};
test_input[33296:33303] = '{32'hc2884199, 32'h41c57625, 32'hc113889b, 32'hc29e1f39, 32'h4282442c, 32'h4123a6f3, 32'hc2929947, 32'hc229427e};
test_weights[33296:33303] = '{32'h42666b00, 32'h416e966e, 32'h420339a3, 32'hc15541f2, 32'h42c22753, 32'hc26a2bb4, 32'h429dbe63, 32'hc2acab16};
test_bias[4162:4162] = '{32'h4220dd9c};
test_output[4162:4162] = '{32'h444fca1f};
test_input[33304:33311] = '{32'h41d84fb4, 32'hc1d088b6, 32'hc133b815, 32'h42bb3976, 32'hc08147f4, 32'hc20ca4d2, 32'h426adf6e, 32'hc27f4eed};
test_weights[33304:33311] = '{32'hc2b53934, 32'hc2205f2a, 32'h41e3594e, 32'h42b20128, 32'hc2094551, 32'h4265e895, 32'h42661a98, 32'hc24ed16e};
test_bias[4163:4163] = '{32'h42068476};
test_output[4163:4163] = '{32'h4632b354};
test_input[33312:33319] = '{32'hc24ca11b, 32'h42959a0d, 32'h420a7047, 32'h42c28f41, 32'hc2b4eafb, 32'hc299f64f, 32'h421c2f56, 32'h42994652};
test_weights[33312:33319] = '{32'h42a11cd7, 32'h41ab04d9, 32'hc2bf04a6, 32'hc299b12e, 32'h417d99b5, 32'hc1b185e8, 32'hc27b2e06, 32'h421f3d16};
test_bias[4164:4164] = '{32'h42b0f4d4};
test_output[4164:4164] = '{32'hc640d4a7};
test_input[33320:33327] = '{32'h41f4edb7, 32'h40269073, 32'hc2525d0f, 32'h4204be51, 32'hc2c5b1c4, 32'h42bd5559, 32'hc28b585b, 32'hc2b9bf69};
test_weights[33320:33327] = '{32'hbf0a79fc, 32'h40cc2316, 32'h41fe277b, 32'hc209827f, 32'hc29a2e1a, 32'h42a8ef3b, 32'hc139f801, 32'hc2292258};
test_bias[4165:4165] = '{32'h4251c02a};
test_output[4165:4165] = '{32'h46897425};
test_input[33328:33335] = '{32'h422cada3, 32'h4249b455, 32'h419833b4, 32'hc1b6bfe6, 32'hc28bbd70, 32'hc2430628, 32'h4200a400, 32'hc247e55b};
test_weights[33328:33335] = '{32'h423efa9c, 32'hc25a5a19, 32'hc1356545, 32'hc25f2ba0, 32'hc2945552, 32'h41c5b2b5, 32'hc2796ce0, 32'h41f3582d};
test_bias[4166:4166] = '{32'hc25f5cc6};
test_output[4166:4166] = '{32'h443ec58d};
test_input[33336:33343] = '{32'h40c7932f, 32'hc2c1a029, 32'h42a265ea, 32'h42bcfecc, 32'hc1cee00b, 32'hc2a498e7, 32'h41ea69b2, 32'h41408ffd};
test_weights[33336:33343] = '{32'h42b6d2a5, 32'h422101f1, 32'h424b3f01, 32'hc22c3c3e, 32'h42602e90, 32'h41694080, 32'hc26c4dfa, 32'h42b7216e};
test_bias[4167:4167] = '{32'hc2bd2050};
test_output[4167:4167] = '{32'hc5cf947e};
test_input[33344:33351] = '{32'h426d948a, 32'hc2a2f924, 32'hc2a5b177, 32'h40b9091a, 32'h41b71450, 32'h41a69235, 32'hc17bc9ac, 32'hbfad467a};
test_weights[33344:33351] = '{32'h40fe1a53, 32'h4200cd53, 32'h4293017b, 32'hc2149322, 32'h4240dee0, 32'hc2b89869, 32'hc2b2f60d, 32'hc2380ff9};
test_bias[4168:4168] = '{32'h42127e00};
test_output[4168:4168] = '{32'hc5f2be37};
test_input[33352:33359] = '{32'hc28f7a1f, 32'h4174e644, 32'h421704d1, 32'h4120814d, 32'hc28bfe96, 32'hc10dc353, 32'h41fa7534, 32'h421ced5e};
test_weights[33352:33359] = '{32'hc074088d, 32'h41a1080b, 32'hc290ac7e, 32'hc197b6bb, 32'hc2b4b6ee, 32'hc2be88e4, 32'h420bff85, 32'hc27be556};
test_bias[4169:4169] = '{32'hc1f26dd9};
test_output[4169:4169] = '{32'h4556009e};
test_input[33360:33367] = '{32'hc233f734, 32'h42a04822, 32'h42af1c69, 32'h4272108f, 32'hc231c0ee, 32'hc158f0da, 32'h41a64d6c, 32'hc2a61e08};
test_weights[33360:33367] = '{32'hc10c8ba2, 32'hc189d4bd, 32'hc1f3c984, 32'hc2aa46fa, 32'hc2b75e41, 32'hc2b46885, 32'h42925271, 32'hc27bab3d};
test_bias[4170:4170] = '{32'hc2650bec};
test_output[4170:4170] = '{32'h4546cdd6};
test_input[33368:33375] = '{32'hc1747e27, 32'hc2b1dd88, 32'h427da05e, 32'h41e83c74, 32'h42c3b230, 32'h41ffeff2, 32'hc280873c, 32'hc11caa08};
test_weights[33368:33375] = '{32'h4192e916, 32'hc1ea94e7, 32'hc2c057b6, 32'h42b2273a, 32'h42c78868, 32'h41bdb9b4, 32'h42b4ae94, 32'hc1b1d6fe};
test_bias[4171:4171] = '{32'hc282d995};
test_output[4171:4171] = '{32'h456624e9};
test_input[33376:33383] = '{32'hc2c30b9e, 32'hc2ab5782, 32'h41f9e529, 32'hbf8b6182, 32'hc2b2f517, 32'hc263866b, 32'hc2218151, 32'hc212594a};
test_weights[33376:33383] = '{32'h42befec7, 32'hbef2c828, 32'h42413549, 32'hc20be943, 32'hc262296e, 32'hc1a01046, 32'h419a0f80, 32'hc296fa72};
test_bias[4172:4172] = '{32'hc2a30ef0};
test_output[4172:4172] = '{32'h43bb37ad};
test_input[33384:33391] = '{32'hc29f49bb, 32'hc2142d2e, 32'h42416685, 32'h4091f890, 32'h4215b614, 32'hc2b5e601, 32'h42898b22, 32'h41759ad7};
test_weights[33384:33391] = '{32'hc259dde0, 32'hc2aa6ed1, 32'hc269e40b, 32'h427fb924, 32'hc264fdd4, 32'hc29829ed, 32'hc2936312, 32'hc2073dc8};
test_bias[4173:4173] = '{32'hc1c69944};
test_output[4173:4173] = '{32'h4580e1fd};
test_input[33392:33399] = '{32'hc1827092, 32'hc276e6ad, 32'hc18ce544, 32'h428743f8, 32'h429320e2, 32'hc29b5b95, 32'hc29381eb, 32'h41d8a821};
test_weights[33392:33399] = '{32'hc28986ca, 32'hc12f637b, 32'hc296ee26, 32'h428902de, 32'h3fb36dee, 32'h41a42421, 32'hc081b0af, 32'hc249c660};
test_bias[4174:4174] = '{32'hc29cc7fc};
test_output[4174:4174] = '{32'h45a01ec2};
test_input[33400:33407] = '{32'hc23c04c7, 32'hc0a43632, 32'h41dde231, 32'h41a7871d, 32'h4247aeaf, 32'hc2a17552, 32'hc2691e1b, 32'h415b4042};
test_weights[33400:33407] = '{32'h418b3981, 32'hc29a90d7, 32'hc17d9109, 32'h418ab62c, 32'h41a992e6, 32'hc1be3637, 32'h426acecd, 32'h420f4f8a};
test_bias[4175:4175] = '{32'hc268efce};
test_output[4175:4175] = '{32'hc3fe5758};
test_input[33408:33415] = '{32'h428fa784, 32'hc185de90, 32'hc0cbfa5a, 32'hc2064689, 32'h412e0757, 32'hc17580ae, 32'hc2afd063, 32'hc21f6834};
test_weights[33408:33415] = '{32'hc23edf8a, 32'h420c74df, 32'h42a83e05, 32'h42583160, 32'h42ae4df4, 32'hc2a9cce1, 32'h40b656c0, 32'h419072cb};
test_bias[4176:4176] = '{32'hc2756dc5};
test_output[4176:4176] = '{32'hc5a8a664};
test_input[33416:33423] = '{32'hc2a4e18e, 32'h426d60f8, 32'hc2a810c0, 32'h4210dc2b, 32'hc22ae015, 32'h4212e80c, 32'h42af04ff, 32'h41c758e7};
test_weights[33416:33423] = '{32'h42939087, 32'hc283e8c2, 32'hc1f93edb, 32'h420dedce, 32'hc201956e, 32'hc298b06f, 32'h3ebd3f14, 32'hc25fa760};
test_bias[4177:4177] = '{32'h42965963};
test_output[4177:4177] = '{32'hc6097d58};
test_input[33424:33431] = '{32'hc2304faa, 32'hc1cd6b92, 32'h429cd001, 32'h4228a5eb, 32'hc23af4ac, 32'h42bf96ca, 32'hc147d69d, 32'h42a1109d};
test_weights[33424:33431] = '{32'hc23ec678, 32'h41896487, 32'hc22ff4b9, 32'h410c058d, 32'hc21cb9e9, 32'hc1542bce, 32'h4286ce8a, 32'hc1cad8eb};
test_bias[4178:4178] = '{32'h42a92351};
test_output[4178:4178] = '{32'hc56490ce};
test_input[33432:33439] = '{32'hc002f829, 32'hc2a40594, 32'hc0dda532, 32'hc1cc49ee, 32'h42864a9b, 32'h425aa994, 32'hc157a7ca, 32'h428f3331};
test_weights[33432:33439] = '{32'h42764ca9, 32'hc12618de, 32'h409c3d58, 32'hc293d4ec, 32'h4122240e, 32'h423c7bb6, 32'h42a5a194, 32'hc2809f0f};
test_bias[4179:4179] = '{32'h42854cf7};
test_output[4179:4179] = '{32'h43352b57};
test_input[33440:33447] = '{32'hc2a722d1, 32'h42a6eb70, 32'h425be4c0, 32'hc1bbd443, 32'h427f04a6, 32'h428e9ad1, 32'h42629943, 32'h4257f1b7};
test_weights[33440:33447] = '{32'hc2224351, 32'hc1622c81, 32'h42247a16, 32'hc1d4371c, 32'h42936a7b, 32'h418bafa5, 32'h41036ccd, 32'hc2341406};
test_bias[4180:4180] = '{32'h421ee78b};
test_output[4180:4180] = '{32'h460e6156};
test_input[33448:33455] = '{32'hc2876b68, 32'hc277a74b, 32'hc2c57406, 32'hc272803b, 32'h42a75a66, 32'hc2650247, 32'h429fc664, 32'hc2b50ec6};
test_weights[33448:33455] = '{32'hc0ae317c, 32'h42103f3e, 32'h4292f766, 32'hc094b1a9, 32'hc0e434e0, 32'hc26f9886, 32'hc2a2abcc, 32'hc22ad9ed};
test_bias[4181:4181] = '{32'hc1f2058e};
test_output[4181:4181] = '{32'hc6076704};
test_input[33456:33463] = '{32'hc1e2aab3, 32'hc25cac55, 32'h404dd1c7, 32'hc0cde38a, 32'hc252bce9, 32'h42910ec3, 32'hc1c3eeda, 32'h42b5cfed};
test_weights[33456:33463] = '{32'h4282d760, 32'hc2b67ea9, 32'h42829caf, 32'hc24004aa, 32'h4226eb9f, 32'h419379cf, 32'hc162a0c7, 32'hc070ebd9};
test_bias[4182:4182] = '{32'h426af7b9};
test_output[4182:4182] = '{32'h4535533b};
test_input[33464:33471] = '{32'h4239294e, 32'h427d23a1, 32'hc2a08f7b, 32'h426b822c, 32'h42561a56, 32'h414f1175, 32'hc15b9c2f, 32'h425d1e0e};
test_weights[33464:33471] = '{32'h42c17b39, 32'h4220a836, 32'h4291c48d, 32'hc28951d3, 32'h4290a11d, 32'hc28a9ab0, 32'hc2ae8041, 32'h428347ee};
test_bias[4183:4183] = '{32'hc216ea99};
test_output[4183:4183] = '{32'h4598c430};
test_input[33472:33479] = '{32'hc236177c, 32'h42b46af0, 32'hc2801c8a, 32'hc1da9ed5, 32'hc2313f68, 32'h41dcbb4a, 32'h40ae80c7, 32'hc1e1e2bf};
test_weights[33472:33479] = '{32'h40772241, 32'hc1624f62, 32'h424e03c1, 32'hc205ecad, 32'h429ec4d8, 32'h42c4344d, 32'hc296b205, 32'h42c7bf18};
test_bias[4184:4184] = '{32'h4149e1fd};
test_output[4184:4184] = '{32'hc5f5c854};
test_input[33480:33487] = '{32'h42a6e9c0, 32'hc2759448, 32'h4153b8c0, 32'hc22dd7e5, 32'h42b7ddcc, 32'h4276cd1e, 32'h4280c62a, 32'hc194697b};
test_weights[33480:33487] = '{32'h4238cd17, 32'h41937984, 32'hc287f845, 32'hc2175e25, 32'h42708478, 32'h429d79cb, 32'h3f6cb066, 32'hc247580f};
test_bias[4185:4185] = '{32'hc20a0d8e};
test_output[4185:4185] = '{32'h46675237};
test_input[33488:33495] = '{32'h42811e13, 32'hc23c7f39, 32'h404abd0d, 32'h42a0be3b, 32'hc1d6f1d3, 32'hc20b8bfd, 32'hc2c69c5a, 32'h41325bd8};
test_weights[33488:33495] = '{32'h4256937c, 32'hc2766ddc, 32'h4281e863, 32'h41dedf17, 32'hc1941b07, 32'h42a69b17, 32'hc190dedf, 32'hc2024c23};
test_bias[4186:4186] = '{32'hc2b48d34};
test_output[4186:4186] = '{32'h45f21af6};
test_input[33496:33503] = '{32'hc29c27f0, 32'h42a69cb9, 32'hc22d80ea, 32'hc06eb0c7, 32'hc2c6b2a6, 32'h42a821af, 32'h4122d8a2, 32'hc2226951};
test_weights[33496:33503] = '{32'hc1dbed21, 32'hc2b125ac, 32'h3fb6a54c, 32'hc2a22728, 32'h41956934, 32'hc2b4da74, 32'h41ca5b80, 32'h4264ce32};
test_bias[4187:4187] = '{32'hc2b8a9e5};
test_output[4187:4187] = '{32'hc681bcff};
test_input[33504:33511] = '{32'hc2807e59, 32'h42550968, 32'h42a4b7ba, 32'hc1ebd47f, 32'hc27b784b, 32'hc24901b4, 32'hc2b8a123, 32'h427ae9d5};
test_weights[33504:33511] = '{32'h40333a41, 32'h429d4820, 32'h429a2b9f, 32'h40bbc7af, 32'h42b70f09, 32'hc1cad41e, 32'hc2b7386d, 32'h429622d8};
test_bias[4188:4188] = '{32'hc2bc254a};
test_output[4188:4188] = '{32'h4692af73};
test_input[33512:33519] = '{32'h429c3904, 32'hc27edeb9, 32'hc2b4a10a, 32'hc24b6338, 32'h41af61a4, 32'hc28f20cc, 32'hc14e9fc9, 32'hc2439034};
test_weights[33512:33519] = '{32'h4281ec0f, 32'hc1fb8ac0, 32'h4249de81, 32'hc1b28849, 32'hc155c314, 32'hc29fa067, 32'h4171ee90, 32'hc272d241};
test_bias[4189:4189] = '{32'h40ae129e};
test_output[4189:4189] = '{32'h46392db1};
test_input[33520:33527] = '{32'hc214b5ca, 32'hc044951e, 32'h4299056c, 32'h42ac1211, 32'h41d6651a, 32'hc13db7f4, 32'h42bcab9f, 32'hc1972412};
test_weights[33520:33527] = '{32'h425be751, 32'h42557a96, 32'hc2985541, 32'hc1df7d87, 32'h41c98066, 32'h429556a5, 32'hc1a3d5b2, 32'hc2306b82};
test_bias[4190:4190] = '{32'hc2898dc0};
test_output[4190:4190] = '{32'hc638a2a4};
test_input[33528:33535] = '{32'hc253afc7, 32'hc28ac724, 32'h429319c0, 32'hc20e0c16, 32'h421ebccd, 32'hc261a4f8, 32'h41975d7e, 32'hc0beabb2};
test_weights[33528:33535] = '{32'h42ad6bdc, 32'hc2bd3450, 32'hc1b01d39, 32'h4197fc7b, 32'hc2bb5224, 32'h41861a2f, 32'hc15168b3, 32'hc290e851};
test_bias[4191:4191] = '{32'hc2bc9882};
test_output[4191:4191] = '{32'hc598d83b};
test_input[33536:33543] = '{32'hc27fc9c6, 32'h41afc11c, 32'hc00ef67c, 32'h4154e430, 32'hc237ebc6, 32'hc21e6b12, 32'h429c7c01, 32'h41c2bcf6};
test_weights[33536:33543] = '{32'h4228dc25, 32'h426c594b, 32'hc0d742cd, 32'h42314359, 32'h415e2072, 32'h41429826, 32'hc13c34a1, 32'h42b1af54};
test_bias[4192:4192] = '{32'hc25900e2};
test_output[4192:4192] = '{32'hc4362ee5};
test_input[33544:33551] = '{32'h41781561, 32'h4093ae08, 32'h423ed707, 32'h4292437d, 32'hc27e9088, 32'h40760074, 32'hc2413adb, 32'hc217dc1c};
test_weights[33544:33551] = '{32'h425b28cc, 32'hc28163f7, 32'hc262770d, 32'h41005bb0, 32'h429f5b4b, 32'hc1f4db96, 32'hc111b330, 32'h4239e71a};
test_bias[4193:4193] = '{32'h42b6c865};
test_output[4193:4193] = '{32'hc5f9890b};
test_input[33552:33559] = '{32'h422ce57e, 32'hc2aee50e, 32'hc24e9122, 32'hc1433900, 32'hc2ad2f49, 32'hc26c2d5c, 32'h4288f478, 32'h4266f1ab};
test_weights[33552:33559] = '{32'h42b522af, 32'h420d73eb, 32'h423cdaa8, 32'hc1a79a3f, 32'h421ae5b4, 32'hc22f70b2, 32'hc270ee22, 32'hc22a7ecb};
test_bias[4194:4194] = '{32'hc12e0c6e};
test_output[4194:4194] = '{32'hc60840cb};
test_input[33560:33567] = '{32'h41ef3dee, 32'h41e03fec, 32'hc2a8921f, 32'h4256b80a, 32'h4280affb, 32'h42c52794, 32'hc1e88d64, 32'h40977009};
test_weights[33560:33567] = '{32'h41e2fdd1, 32'h418d1595, 32'hc1d530b2, 32'h427605c6, 32'hc1fb3d7c, 32'hc0f91d96, 32'hc29348f5, 32'hc0a31a11};
test_bias[4195:4195] = '{32'hc2174877};
test_output[4195:4195] = '{32'h45c129da};
test_input[33568:33575] = '{32'h4126f2e8, 32'hc22d41e3, 32'h41eb4d53, 32'hc2a2ccee, 32'h428fd987, 32'hc28c4446, 32'h41afe50d, 32'h4217cb93};
test_weights[33568:33575] = '{32'h42bab5d9, 32'h420bc96d, 32'hc1baeafc, 32'h41d5b83a, 32'hc182b3b1, 32'hc2c70fbb, 32'hc2bb54dd, 32'h424b1677};
test_bias[4196:4196] = '{32'hc1cb713c};
test_output[4196:4196] = '{32'h450c5cce};
test_input[33576:33583] = '{32'h42a46963, 32'hc2119e5f, 32'h42adfc65, 32'hc06a0025, 32'h42963e76, 32'h419ff808, 32'h42b65dcc, 32'hc2a2539d};
test_weights[33576:33583] = '{32'h428c8d8f, 32'h41d8f93a, 32'h42aa9bb5, 32'h416469db, 32'hc2a908ca, 32'hc1db05c1, 32'hc2bd5578, 32'h42a33913};
test_bias[4197:4197] = '{32'hc1961b72};
test_output[4197:4197] = '{32'hc61c730a};
test_input[33584:33591] = '{32'hc294e1db, 32'hc2710fd9, 32'h4146e290, 32'hc24d0ca4, 32'h425982df, 32'hc2303c03, 32'h42c40b96, 32'h42a9ee2c};
test_weights[33584:33591] = '{32'hc25fb900, 32'hc2ac3502, 32'hc0c43864, 32'hc29a6c2d, 32'hc1b4ed3f, 32'hc1e2e841, 32'h426e4ca7, 32'hc19bab8e};
test_bias[4198:4198] = '{32'hc1d28267};
test_output[4198:4198] = '{32'h46880ca7};
test_input[33592:33599] = '{32'h42c5f702, 32'hc23cdf48, 32'hc24f12ee, 32'h4285413a, 32'hc2703048, 32'hc2156e36, 32'hc2a80d89, 32'hc166ec52};
test_weights[33592:33599] = '{32'hc038e6cf, 32'hc1c8d902, 32'hc23e3efa, 32'h4220b3ae, 32'hc2c6d06b, 32'hc25873cc, 32'h4241eec2, 32'h4163d78b};
test_bias[4199:4199] = '{32'h41d0cd9c};
test_output[4199:4199] = '{32'h4618bf44};
test_input[33600:33607] = '{32'h424da8fd, 32'hbf61544c, 32'hbe46482a, 32'hc281b876, 32'h42207d0c, 32'h42661e79, 32'hc1c60382, 32'hc1d21c7a};
test_weights[33600:33607] = '{32'hc2ac6fb8, 32'h428d49f9, 32'hc23b03d1, 32'hc234a245, 32'hc281d4f1, 32'h428696c5, 32'hc20a16eb, 32'h41d91728};
test_bias[4200:4200] = '{32'h42316b3f};
test_output[4200:4200] = '{32'hc2d01451};
test_input[33608:33615] = '{32'hc1241144, 32'h4211b933, 32'hc2ab3520, 32'hc0ef47da, 32'h423e915d, 32'hc126dc0d, 32'hc195097a, 32'hc15f446f};
test_weights[33608:33615] = '{32'hc22cb3bf, 32'h4173f4ff, 32'hc203289c, 32'h42b23760, 32'hc27aefe2, 32'h42075582, 32'hc2358b68, 32'hc289d705};
test_bias[4201:4201] = '{32'hc1a9d810};
test_output[4201:4201] = '{32'h44c5e6bc};
test_input[33616:33623] = '{32'hc1fbf3be, 32'hc2c2a964, 32'h41c0f606, 32'h41ede2b8, 32'hc23573ba, 32'hc2059f47, 32'h42c6d41e, 32'h429fb2a6};
test_weights[33616:33623] = '{32'hc16c6833, 32'hc28fd56e, 32'h4214dacc, 32'hc2acdfc2, 32'h423aed83, 32'hc2bd077a, 32'h426e54d6, 32'h401ba0ac};
test_bias[4202:4202] = '{32'h425d6a8f};
test_output[4202:4202] = '{32'h464b2add};
test_input[33624:33631] = '{32'h42502fd5, 32'hc28abf69, 32'h428c22b3, 32'h40b97859, 32'h4222589c, 32'h429e14a2, 32'h414bf23f, 32'h4269edb5};
test_weights[33624:33631] = '{32'hc1c44961, 32'h411bd3c8, 32'h413756dc, 32'h424a35de, 32'hc198e7ce, 32'h428e562c, 32'hc2096e07, 32'h4298827e};
test_bias[4203:4203] = '{32'h427c5288};
test_output[4203:4203] = '{32'h45fc6abd};
test_input[33632:33639] = '{32'hc2a77663, 32'hc29d32d6, 32'hc2820d44, 32'hc25c91ed, 32'h41d0242b, 32'h4283bea8, 32'hc2974f23, 32'h4236ba48};
test_weights[33632:33639] = '{32'h426b6da3, 32'h42a53c8b, 32'hc2194ab7, 32'h42a5021a, 32'hc1207b9e, 32'hc2bd3c93, 32'hc2a339e4, 32'hc2b4bf2e};
test_bias[4204:4204] = '{32'hc1adbd2b};
test_output[4204:4204] = '{32'hc68c39b2};
test_input[33640:33647] = '{32'hc2600d45, 32'h42a20d27, 32'hc22715b5, 32'hc14f9158, 32'h41fd9159, 32'h427d325f, 32'h415940cf, 32'hc1fb4a76};
test_weights[33640:33647] = '{32'hc05800a1, 32'hc257a61f, 32'hc2c2ffc6, 32'hc276ce99, 32'hc199bb1d, 32'h40b97cc9, 32'hc2b45c11, 32'hc0cad3cc};
test_bias[4205:4205] = '{32'h401341d1};
test_output[4205:4205] = '{32'hc40ed730};
test_input[33648:33655] = '{32'hc12756fb, 32'hc22c1fd3, 32'hc1a04b64, 32'hc270c511, 32'hc0357657, 32'hc1e67ba4, 32'h42a796fe, 32'hc2989b34};
test_weights[33648:33655] = '{32'h4259298f, 32'h41bab8e8, 32'h42619351, 32'h4280f8ee, 32'h42bfe006, 32'h429f9ac6, 32'hbca03777, 32'hc23138f4};
test_bias[4206:4206] = '{32'hc21b0561};
test_output[4206:4206] = '{32'hc5b5b4b9};
test_input[33656:33663] = '{32'h42a9a089, 32'h42b759d4, 32'h40d7c26e, 32'h4243ee74, 32'hc2aa7bab, 32'h4255ec1e, 32'h42aff76e, 32'h42c3ca93};
test_weights[33656:33663] = '{32'h42919950, 32'hc1a5ef99, 32'h42a9343c, 32'h424fa05f, 32'hc28c38eb, 32'h3f86eee6, 32'hc001d4fd, 32'h424b967d};
test_bias[4207:4207] = '{32'h42976baa};
test_output[4207:4207] = '{32'h468ef4c6};
test_input[33664:33671] = '{32'hc1b87303, 32'hc06a1acb, 32'hc2699ffd, 32'h41ba5bc2, 32'hc192f7c7, 32'hc285ab1e, 32'hc16cea84, 32'hc29927f9};
test_weights[33664:33671] = '{32'hc2be6d69, 32'h42841e33, 32'h420aeb94, 32'hc2491b6d, 32'h40e7b7ab, 32'h4138d165, 32'hc2945f9a, 32'h424fb6a0};
test_bias[4208:4208] = '{32'hc26ea6b4};
test_output[4208:4208] = '{32'hc59f0648};
test_input[33672:33679] = '{32'h428cf7c8, 32'h42c664af, 32'h42717262, 32'hc1ff4977, 32'h4177c863, 32'hc0fc4768, 32'h42515a67, 32'h40dc9e1f};
test_weights[33672:33679] = '{32'h4113f8d4, 32'hc1e2e38d, 32'h4223552b, 32'h41ec5b00, 32'h402835fd, 32'h42150bb3, 32'h420d81a6, 32'h40c13cdb};
test_bias[4209:4209] = '{32'h420be597};
test_output[4209:4209] = '{32'h4481732d};
test_input[33680:33687] = '{32'h42b1bbff, 32'hc2a7f7ec, 32'hc2b0f5e4, 32'hc265840d, 32'h41fcbd9d, 32'hc2366481, 32'h421fb5e0, 32'hc2001a9a};
test_weights[33680:33687] = '{32'h42842f1b, 32'h421bdda3, 32'h42513efb, 32'hc2ac5933, 32'hc232d0c2, 32'hc211c90b, 32'hc11a3699, 32'h417fd74b};
test_bias[4210:4210] = '{32'h41693052};
test_output[4210:4210] = '{32'h450ec1c4};
test_input[33688:33695] = '{32'hc29acf36, 32'h42037469, 32'h41c1cb70, 32'h420a8e49, 32'hc2943078, 32'hc2081cc2, 32'hc2a676ee, 32'h42846698};
test_weights[33688:33695] = '{32'hc2c24751, 32'hc1177d9f, 32'h4218ee99, 32'h41b25fb3, 32'h428c45e0, 32'h41cda378, 32'hc1c5b430, 32'hc2311209};
test_bias[4211:4211] = '{32'hc20a583a};
test_output[4211:4211] = '{32'h44f0d849};
test_input[33696:33703] = '{32'h42afd243, 32'h41a3e988, 32'hc29d7424, 32'hc28c1438, 32'h428bc8eb, 32'h428b0914, 32'h42c790a0, 32'hc18bc3db};
test_weights[33696:33703] = '{32'h4226f30c, 32'hc1cea86c, 32'hc2c3b5ab, 32'h4232ba49, 32'h42be2a42, 32'h42831069, 32'hc08b8b75, 32'h429cb84f};
test_bias[4212:4212] = '{32'h4281bfe2};
test_output[4212:4212] = '{32'h4686303c};
test_input[33704:33711] = '{32'h42119727, 32'h41c59c87, 32'h422ffdd6, 32'h4289516f, 32'h41bb2ef6, 32'h41bffee3, 32'hc29443c5, 32'h406fb469};
test_weights[33704:33711] = '{32'h42abe16c, 32'hc2a4934d, 32'h424de79e, 32'hc1b6e726, 32'hc28a8aaa, 32'h42870fc6, 32'hc2b5f2ad, 32'hc2484092};
test_bias[4213:4213] = '{32'h4125fcde};
test_output[4213:4213] = '{32'h46029591};
test_input[33712:33719] = '{32'h412b3792, 32'h422a964a, 32'h42b5bba5, 32'h4298519c, 32'hc2bb7f2f, 32'hc1479021, 32'hc163ed22, 32'h42663951};
test_weights[33712:33719] = '{32'h3fc9b720, 32'h4121aabb, 32'hc1ffd15e, 32'h42a0f5da, 32'h41dea00a, 32'h427ce671, 32'h42246e56, 32'hc24cd35a};
test_bias[4214:4214] = '{32'h429b9902};
test_output[4214:4214] = '{32'hc546d064};
test_input[33720:33727] = '{32'h418c7b54, 32'h4286e1a2, 32'h4253f7ca, 32'h42b355f1, 32'hc20b47b1, 32'hc187b6fe, 32'hc271f1ac, 32'hc227066a};
test_weights[33720:33727] = '{32'h423d69fd, 32'hc254b096, 32'hc23d19fb, 32'hc2b1fbdc, 32'h4210f793, 32'h42512387, 32'hc25a640f, 32'h41459e03};
test_bias[4215:4215] = '{32'h4214ed57};
test_output[4215:4215] = '{32'hc6445197};
test_input[33728:33735] = '{32'hc2935ef3, 32'hc241a51a, 32'h40b695fe, 32'hc1f4c100, 32'h4292e037, 32'hc03c2e70, 32'h42810ba1, 32'h42531e1c};
test_weights[33728:33735] = '{32'hc19f0a8c, 32'h426d45bf, 32'h4218f128, 32'h4129fb2e, 32'hc222a1b0, 32'hc1a17e9f, 32'hc1e54af7, 32'hc2254a32};
test_bias[4216:4216] = '{32'hc22446d5};
test_output[4216:4216] = '{32'hc604fdf8};
test_input[33736:33743] = '{32'h4241ed45, 32'hc2940638, 32'h4283495c, 32'hc1148d69, 32'h41108f2e, 32'h42a34bf6, 32'hc2b88c63, 32'h42245e47};
test_weights[33736:33743] = '{32'hc1a5e55f, 32'h42881d89, 32'h4235a970, 32'hc2c6f4ac, 32'h426e92df, 32'h42acd0b9, 32'h40cfc9da, 32'hc2bc3d33};
test_bias[4217:4217] = '{32'h42a8fcb3};
test_output[4217:4217] = '{32'h44864143};
test_input[33744:33751] = '{32'hc282c3d7, 32'hc1f00a51, 32'h426cd13c, 32'h4281d077, 32'h40a389df, 32'hc28418f2, 32'hc292344c, 32'hc26e7c3f};
test_weights[33744:33751] = '{32'h42c191e2, 32'hc287eb6e, 32'h42844feb, 32'hc2b48b4c, 32'hc0f543bf, 32'h42869ecb, 32'h4259ad56, 32'hc00ec584};
test_bias[4218:4218] = '{32'hc0aea06e};
test_output[4218:4218] = '{32'hc6639c11};
test_input[33752:33759] = '{32'hc2a0dd4b, 32'h42888119, 32'hc1348361, 32'h42640271, 32'h42603f06, 32'h42557e3d, 32'h40acee89, 32'hc1953594};
test_weights[33752:33759] = '{32'hc1d7b156, 32'h429f7863, 32'hc2479a57, 32'hc1db35ed, 32'hc2073db9, 32'h4056d7eb, 32'hc21ca062, 32'h4295da57};
test_bias[4219:4219] = '{32'hc161df44};
test_output[4219:4219] = '{32'h454c83db};
test_input[33760:33767] = '{32'hc277af39, 32'h428ea519, 32'hc1f43664, 32'h42515e44, 32'hc23963c6, 32'h41ee5125, 32'hc2b1bb1b, 32'h42626c89};
test_weights[33760:33767] = '{32'hc266a988, 32'hc110c987, 32'hc1f88325, 32'hc2a5b15d, 32'hc2bfe797, 32'hc293a323, 32'hc265d3d7, 32'hc2c3f630};
test_bias[4220:4220] = '{32'h42ad097c};
test_output[4220:4220] = '{32'h44b2efc3};
test_input[33768:33775] = '{32'h41be0b05, 32'hbf514932, 32'hc241dcb7, 32'hc24da361, 32'h4210dc70, 32'hc23a3442, 32'h41f74093, 32'h4180a03a};
test_weights[33768:33775] = '{32'hc2a6cd41, 32'hc2a0b61d, 32'hc0d46632, 32'h42bfdb35, 32'hc2b4278c, 32'h42b364b4, 32'h4231ef5a, 32'h4176bea6};
test_bias[4221:4221] = '{32'hc1a253b9};
test_output[4221:4221] = '{32'hc641226e};
test_input[33776:33783] = '{32'h42af29ab, 32'h421528b9, 32'h427f7b04, 32'hc235ed18, 32'h42af140f, 32'h425ce525, 32'hc26b8951, 32'hc24bd05a};
test_weights[33776:33783] = '{32'hc240993e, 32'h421f092d, 32'h41ef9d8b, 32'hc1a09e85, 32'hc2253882, 32'hc2a36a64, 32'h42abbea6, 32'hc1a942d2};
test_bias[4222:4222] = '{32'hc1532a74};
test_output[4222:4222] = '{32'hc63befaf};
test_input[33784:33791] = '{32'h429aa50d, 32'h42c45c62, 32'hc2075bd7, 32'hc21a65e1, 32'hc294e5a2, 32'h41fa9dce, 32'h422bebe7, 32'hc276ebe1};
test_weights[33784:33791] = '{32'h426e59d6, 32'h419fe765, 32'h426e4038, 32'h42a3d01b, 32'h42c0bccd, 32'hc1bf1f75, 32'h4170db55, 32'hc2a6faff};
test_bias[4223:4223] = '{32'h42a0a336};
test_output[4223:4223] = '{32'hc4223d1c};
test_input[33792:33799] = '{32'h4286b59d, 32'hc235f406, 32'h4231ec7b, 32'h424c7bd0, 32'h426f7ad7, 32'h41da1dd8, 32'h4292b067, 32'hc29b5e18};
test_weights[33792:33799] = '{32'h429330c3, 32'hc2747b92, 32'hc2c7c419, 32'h401ef690, 32'hc2c64ab6, 32'h42a1307c, 32'hc2a000b2, 32'hc1ea11df};
test_bias[4224:4224] = '{32'h42b3e391};
test_output[4224:4224] = '{32'hc56eded1};
test_input[33800:33807] = '{32'hc1eef505, 32'hc1669f36, 32'hc1cd86a1, 32'h41df8759, 32'hc136adbc, 32'h42ac5604, 32'hc1becd87, 32'h424216f4};
test_weights[33800:33807] = '{32'h413185a6, 32'hc13b0f87, 32'h41aa453c, 32'h3d7d1c50, 32'h4215b339, 32'h41d8ec22, 32'h42b62e20, 32'h42bb3aa2};
test_bias[4225:4225] = '{32'h423075fb};
test_output[4225:4225] = '{32'h4561f333};
test_input[33808:33815] = '{32'h42190d8b, 32'hc0e706c9, 32'hc2b0cc35, 32'hc277bb1d, 32'h426dd690, 32'hc1daab20, 32'h41c78055, 32'hc2c760c4};
test_weights[33808:33815] = '{32'h418c1b6b, 32'hbfb679b9, 32'h4297cbab, 32'h41ca72c7, 32'hc1da40fd, 32'h425a3f9e, 32'h3e6b98ec, 32'h420c6058};
test_bias[4226:4226] = '{32'hc2823886};
test_output[4226:4226] = '{32'hc65eee2a};
test_input[33816:33823] = '{32'hc29edff6, 32'h41874e95, 32'h42c77575, 32'hc2591fef, 32'h404ca571, 32'h429cc050, 32'hc29e8a42, 32'hc2178d1f};
test_weights[33816:33823] = '{32'h41c93afb, 32'h4103f2f0, 32'h41957aee, 32'hc285e79d, 32'h42b09d14, 32'hc2b85213, 32'hc2afd08d, 32'h421c5e93};
test_bias[4227:4227] = '{32'h428c2a88};
test_output[4227:4227] = '{32'h450cfa78};
test_input[33824:33831] = '{32'hc23c836a, 32'hc22f412b, 32'h423f0511, 32'hc1c8823d, 32'h42bf6ea7, 32'hc1c0fadd, 32'hc135806b, 32'h42546feb};
test_weights[33824:33831] = '{32'h42952535, 32'hc1407c5a, 32'h41cc44db, 32'h4241b0bc, 32'hc10344e0, 32'h42c4d24f, 32'h42c68f08, 32'hc2ae5cbb};
test_bias[4228:4228] = '{32'hc1aa7249};
test_output[4228:4228] = '{32'hc63a3a16};
test_input[33832:33839] = '{32'h4278370e, 32'h41a5a25f, 32'hc135acc4, 32'hc25b3fee, 32'h4262c3ee, 32'hc193be1d, 32'hc24212cb, 32'hc1d8bdad};
test_weights[33832:33839] = '{32'hc1df3193, 32'h428ed1a7, 32'h414b670f, 32'h4255c22f, 32'hc1b23357, 32'h42ba112d, 32'hc266af26, 32'hc172ca12};
test_bias[4229:4229] = '{32'hc1f15987};
test_output[4229:4229] = '{32'hc5438280};
test_input[33840:33847] = '{32'hc15b0823, 32'hc0d3c32b, 32'hc2ab4459, 32'hc21a22fe, 32'h41db7b27, 32'hc291855e, 32'h425f9c9b, 32'h4234b2fd};
test_weights[33840:33847] = '{32'h41d466c7, 32'h42256742, 32'h4245444a, 32'h42aba34a, 32'h41dd947f, 32'hc2b64a71, 32'h42759d27, 32'h42941472};
test_bias[4230:4230] = '{32'hc28ef66f};
test_output[4230:4230] = '{32'h45b952b2};
test_input[33848:33855] = '{32'h41b7fdc5, 32'h41cf5b31, 32'hc1818def, 32'hc181e90f, 32'hbf90e7f5, 32'hc2c79176, 32'h41f2417c, 32'hc0c5cbcf};
test_weights[33848:33855] = '{32'h4272d9f5, 32'h41f06557, 32'hc1855dae, 32'hc29a0170, 32'hc21e72c4, 32'hc0d739a7, 32'hc28ec9a8, 32'h42502c4e};
test_bias[4231:4231] = '{32'h4127d41b};
test_output[4231:4231] = '{32'h44f24db7};
test_input[33856:33863] = '{32'hc29f0090, 32'h42bb0cfa, 32'h42ad50e6, 32'h425628bb, 32'h41cd6a35, 32'h412a5bd4, 32'hc26838cf, 32'hc176fc6b};
test_weights[33856:33863] = '{32'hc297dbf7, 32'h42a47771, 32'h41308452, 32'hc225717b, 32'hc20ed797, 32'h42be680f, 32'hc0e2b97d, 32'hc2c2869e};
test_bias[4232:4232] = '{32'h3fdaf716};
test_output[4232:4232] = '{32'h466240a5};
test_input[33864:33871] = '{32'h42c28b5d, 32'hc27a751c, 32'h40b121fe, 32'h4256129b, 32'hc2c18595, 32'hc2b350ad, 32'h42af6d25, 32'hc232f58f};
test_weights[33864:33871] = '{32'h42924b3f, 32'h42b571b2, 32'h427284c4, 32'h414b0c4a, 32'hc2553168, 32'h4275dfdd, 32'hc2892d16, 32'hc2356264};
test_bias[4233:4233] = '{32'hc1b91a84};
test_output[4233:4233] = '{32'hc4ef5dfb};
test_input[33872:33879] = '{32'hc18f319f, 32'h42c15598, 32'hc1a56a5b, 32'hc2937404, 32'hc2814c17, 32'hc2b512b6, 32'h42b4126d, 32'hc1d34e60};
test_weights[33872:33879] = '{32'hc1fba7c6, 32'h419e0f87, 32'hc29b3e13, 32'hc25923d1, 32'hc22d5c68, 32'hc26614ea, 32'h429a83e1, 32'h4229c9dc};
test_bias[4234:4234] = '{32'hc2bc73e6};
test_output[4234:4234] = '{32'h46aa8cac};
test_input[33880:33887] = '{32'h42c23e60, 32'hc2918a3c, 32'hc2404584, 32'hc2a8bf41, 32'h42c375e0, 32'hc2b1ce94, 32'h42911abc, 32'hc0239a09};
test_weights[33880:33887] = '{32'h411226d9, 32'hc2a442c8, 32'hc26a9517, 32'hc234fea5, 32'hc2c3118c, 32'h427b4069, 32'h41cbc20a, 32'h4292856e};
test_bias[4235:4235] = '{32'hc1fb999e};
test_output[4235:4235] = '{32'h4156165d};
test_input[33888:33895] = '{32'h42943c6b, 32'h41b0428b, 32'hc22151f9, 32'hc2b2ae86, 32'h41a6e7c8, 32'hc24230c3, 32'hc1fc9ca8, 32'h42ae91a5};
test_weights[33888:33895] = '{32'h42706937, 32'hc293c4ee, 32'hc2019796, 32'hc2c5c884, 32'h41a67ed2, 32'h420e6839, 32'h4255637c, 32'hc28b551e};
test_bias[4236:4236] = '{32'h4194ad45};
test_output[4236:4236] = '{32'h457579ee};
test_input[33896:33903] = '{32'h42bcbb68, 32'h42a972d3, 32'h428eae84, 32'h42260820, 32'hc180610d, 32'h40a95da9, 32'h41c3c5cb, 32'h41dc9a23};
test_weights[33896:33903] = '{32'hc1e7d8f7, 32'hc2b3a02c, 32'h411d6b7f, 32'hc1f08810, 32'h427336f0, 32'hc1eb6fb9, 32'hc2a217dc, 32'h429ff49d};
test_bias[4237:4237] = '{32'h41a297fc};
test_output[4237:4237] = '{32'hc6380d5d};
test_input[33904:33911] = '{32'h42c58e8f, 32'hc09fa37d, 32'hbc7eaa3e, 32'h42b0f5bb, 32'h41feba97, 32'hc224aa55, 32'hc27c1eca, 32'h421605a2};
test_weights[33904:33911] = '{32'h425a1ee8, 32'hc0bdb043, 32'h42049d85, 32'hc020206a, 32'hc29e919b, 32'hc2472297, 32'h42bfd242, 32'hc2825561};
test_bias[4238:4238] = '{32'hc182a85d};
test_output[4238:4238] = '{32'hc56cab2c};
test_input[33912:33919] = '{32'h429eff16, 32'hc1298b66, 32'hc216edfa, 32'h429cbb48, 32'h42a123aa, 32'hc2867698, 32'hc205e88d, 32'h40a6732e};
test_weights[33912:33919] = '{32'h429a1ebe, 32'hc2aed98c, 32'hc1530b10, 32'h42c4275b, 32'h429e69d1, 32'h42595088, 32'h426ac341, 32'h4273fb47};
test_bias[4239:4239] = '{32'h42238767};
test_output[4239:4239] = '{32'h467f9a11};
test_input[33920:33927] = '{32'hc1f888d9, 32'hc21f1a29, 32'hc29d08bf, 32'hc2451a78, 32'h413d7488, 32'h42b39eda, 32'h41ddd464, 32'h42b77dcd};
test_weights[33920:33927] = '{32'hc26d48f1, 32'hc1956c19, 32'hc248b4c6, 32'h428f107d, 32'h423fe37e, 32'h41b0f61f, 32'h41da44bf, 32'hc2b8a08a};
test_bias[4240:4240] = '{32'hc16c3791};
test_output[4240:4240] = '{32'hc507c325};
test_input[33928:33935] = '{32'h421a3bd4, 32'hc2744022, 32'h420a4b43, 32'h41c987ca, 32'hc2249f49, 32'hc2c22782, 32'hc21b0ae7, 32'hc283ba4c};
test_weights[33928:33935] = '{32'hc29577d1, 32'hc1a500e5, 32'hc2b5aa9b, 32'h41fc1ef7, 32'h4282afd3, 32'h42b5fdea, 32'h42448e7e, 32'hc2c501a4};
test_bias[4241:4241] = '{32'hc2bb34d3};
test_output[4241:4241] = '{32'hc62be823};
test_input[33936:33943] = '{32'hc2a7246b, 32'hc2c6ea22, 32'hc103970a, 32'h427a3bab, 32'hc2c725ab, 32'hc1ccb010, 32'hc27c657a, 32'hc21569d6};
test_weights[33936:33943] = '{32'hc05988f2, 32'hc05ef0f6, 32'hc2a12ed4, 32'h41b3f269, 32'h42b6e090, 32'hc2b43444, 32'hc29d4260, 32'hc20cf94f};
test_bias[4242:4242] = '{32'hc04f7782};
test_output[4242:4242] = '{32'h4507fa20};
test_input[33944:33951] = '{32'hc2117bab, 32'hc257771c, 32'h4166ffe4, 32'h4270395b, 32'hc24a089e, 32'hc19e0d4c, 32'hc2908837, 32'hc256b12d};
test_weights[33944:33951] = '{32'hc2068eed, 32'h42a8737d, 32'h42030af7, 32'h4287cfad, 32'hc246888f, 32'hc2c1de6c, 32'h42800394, 32'h42077d85};
test_bias[4243:4243] = '{32'h422137aa};
test_output[4243:4243] = '{32'hc439e581};
test_input[33952:33959] = '{32'hc284353a, 32'hc2a9b719, 32'hc22ba43d, 32'hc13eabf4, 32'h42c7c934, 32'h42be8709, 32'h408f6c93, 32'h42b3294f};
test_weights[33952:33959] = '{32'h41e9ee3e, 32'hc252fb1b, 32'h41f57a5d, 32'hc2c64491, 32'hc2bfd645, 32'hc2ba833c, 32'hc19f59ad, 32'h4272181f};
test_bias[4244:4244] = '{32'h42b198fc};
test_output[4244:4244] = '{32'hc62632de};
test_input[33960:33967] = '{32'h42b8961a, 32'hc2bb3ebe, 32'hc25c0b2e, 32'hc1b95a6f, 32'h4266bea1, 32'h42831287, 32'h41062e56, 32'hc27b270a};
test_weights[33960:33967] = '{32'hc1f5add8, 32'h412e95e2, 32'h423e399b, 32'h414959bd, 32'hc1e8f226, 32'hc2c3385d, 32'h412ac78c, 32'h4298b062};
test_bias[4245:4245] = '{32'hc2813d01};
test_output[4245:4245] = '{32'hc69931d4};
test_input[33968:33975] = '{32'h42bddd8f, 32'h42a97afc, 32'hc2c473b3, 32'hc22035a8, 32'h41d05800, 32'hc2abd8a9, 32'h42a740a4, 32'h4195f404};
test_weights[33968:33975] = '{32'hc1bfed54, 32'hc2696be7, 32'h42003b5c, 32'h429024e6, 32'h41d61d26, 32'hc19e0996, 32'h402b339e, 32'hc2a8b209};
test_bias[4246:4246] = '{32'hc296d9c8};
test_output[4246:4246] = '{32'hc64021fc};
test_input[33976:33983] = '{32'h423a24f2, 32'h42bdbc8c, 32'h4213b7bb, 32'hc0d531dd, 32'h40eb6291, 32'h4198313e, 32'hc1b3ac65, 32'h424526fb};
test_weights[33976:33983] = '{32'hc103be71, 32'h422b873a, 32'h421f906b, 32'h41f01223, 32'hc282bede, 32'hc1061ad4, 32'h3f6af9f6, 32'h42013bc4};
test_bias[4247:4247] = '{32'hc2a4ab7e};
test_output[4247:4247] = '{32'h45b57ab9};
test_input[33984:33991] = '{32'hc1d5356d, 32'hc26a08e1, 32'h40d59aa9, 32'h42b0adcb, 32'hc284e324, 32'hc210eaaa, 32'h42ad925d, 32'hc2999572};
test_weights[33984:33991] = '{32'h42bda327, 32'h42307963, 32'hc207d8c7, 32'h41979d1a, 32'h424ba379, 32'h4270f652, 32'hc265600e, 32'h40287568};
test_bias[4248:4248] = '{32'h42a30d0a};
test_output[4248:4248] = '{32'hc65fccb3};
test_input[33992:33999] = '{32'hc276d50e, 32'hc240a22d, 32'h41fd4a89, 32'h42483677, 32'h424aa227, 32'h4227b355, 32'hc20acf37, 32'h42a1f4c7};
test_weights[33992:33999] = '{32'h417ddcb6, 32'hc2ab7a85, 32'h42c1f0a6, 32'h42a25819, 32'h42991b24, 32'h4207ad0c, 32'hc21857ab, 32'h42c6bbe1};
test_bias[4249:4249] = '{32'hc23a8dc9};
test_output[4249:4249] = '{32'h46c29191};
test_input[34000:34007] = '{32'hc0a8250c, 32'h42748bc0, 32'h415ee116, 32'h41aac99e, 32'h42317cd2, 32'hc27065bf, 32'h4049c78c, 32'hc24eb786};
test_weights[34000:34007] = '{32'h42a8dcf3, 32'hc1c066c8, 32'hc19251b1, 32'h41ec2ff5, 32'hc2a11916, 32'h41c12f39, 32'hc210c080, 32'h40a4f689};
test_bias[4250:4250] = '{32'h42848e62};
test_output[4250:4250] = '{32'hc5d6f0e3};
test_input[34008:34015] = '{32'hc2abad93, 32'hc2b9be72, 32'h41284526, 32'hc2921b79, 32'hc244ffa8, 32'h42aefccc, 32'h4238c1ce, 32'hc2a4d373};
test_weights[34008:34015] = '{32'h42a5865c, 32'hc1a4578d, 32'hc2a6c2ed, 32'hbd756261, 32'h42b6b452, 32'hc27cc7b8, 32'hc1a67888, 32'h4212e6f6};
test_bias[4251:4251] = '{32'hc1a31825};
test_output[4251:4251] = '{32'hc69d12b7};
test_input[34016:34023] = '{32'h4292c868, 32'h4290cb71, 32'hc2c619c4, 32'hc298fbd3, 32'hc2b67a5f, 32'hc25b8eea, 32'h42177715, 32'hc0122247};
test_weights[34016:34023] = '{32'h42aa5cb9, 32'h420c1630, 32'hc2304173, 32'hc200e9db, 32'h424aedad, 32'hc248791e, 32'hc2b7ae2b, 32'hc2081c84};
test_bias[4252:4252] = '{32'h42965f58};
test_output[4252:4252] = '{32'h4622b901};
test_input[34024:34031] = '{32'hc1ce048e, 32'hc19573a7, 32'hc1cebbad, 32'h4285fec7, 32'hc19efbec, 32'h428a5fe9, 32'hc25b3c09, 32'hc2b8ad4c};
test_weights[34024:34031] = '{32'hc2b5a641, 32'hc22230fc, 32'hc25d1081, 32'h424b3bb8, 32'hc25f8462, 32'hc2bc6a69, 32'h4190a00a, 32'hc2166607};
test_bias[4253:4253] = '{32'hc10c08b0};
test_output[4253:4253] = '{32'h459c0b83};
test_input[34032:34039] = '{32'h4191da0e, 32'hc1cd0b08, 32'h425fb922, 32'h41e146f1, 32'hc2bb89ae, 32'h42a49aa5, 32'h419bc726, 32'h40931ec2};
test_weights[34032:34039] = '{32'h41f4735f, 32'hc23abfee, 32'h42c32dee, 32'hc28a45e6, 32'h42823bba, 32'hc2bd31b3, 32'hc29d95a4, 32'h42ac1e79};
test_bias[4254:4254] = '{32'hc249e2c4};
test_output[4254:4254] = '{32'hc6195da3};
test_input[34040:34047] = '{32'hc2763fd3, 32'h42609be2, 32'h42be05d6, 32'hc1236193, 32'hc08702ae, 32'h42c7bd3b, 32'hc25b5e0e, 32'hc2a794a7};
test_weights[34040:34047] = '{32'h425bce42, 32'hbf63c263, 32'hc0411076, 32'hc2c18167, 32'hc2b00c3b, 32'h42b16ddc, 32'hc2b82617, 32'hc29cc8fe};
test_bias[4255:4255] = '{32'hc1f7f756};
test_output[4255:4255] = '{32'h468d4d9c};
test_input[34048:34055] = '{32'hc286bb1c, 32'h41c516d2, 32'h429b3466, 32'h40d92fa2, 32'h420dbf75, 32'hc25d460f, 32'hc28a2188, 32'h426886ef};
test_weights[34048:34055] = '{32'h41945940, 32'hc2872ae3, 32'h42a1d823, 32'h4128bbaf, 32'h418719f4, 32'h40396842, 32'h42091dbe, 32'h424c9909};
test_bias[4256:4256] = '{32'hc1d7d0d7};
test_output[4256:4256] = '{32'h458b31f9};
test_input[34056:34063] = '{32'h41d665eb, 32'h42953bc3, 32'hc284f1ea, 32'hc28c460e, 32'h42032939, 32'h41d76337, 32'hc1a20d7a, 32'h424164fd};
test_weights[34056:34063] = '{32'h3fac8f3b, 32'h42975641, 32'h40eacef1, 32'h41940361, 32'h42006a9c, 32'hc274e272, 32'hc2af8cbe, 32'h427826af};
test_bias[4257:4257] = '{32'h42857aba};
test_output[4257:4257] = '{32'h45fe8bca};
test_input[34064:34071] = '{32'h4289af86, 32'h42a9f100, 32'hbf130727, 32'h4254f995, 32'h42a18155, 32'hc1d03d32, 32'hc29bdd72, 32'h41cc1eff};
test_weights[34064:34071] = '{32'h42beb87d, 32'hc2842d9b, 32'hc20fec94, 32'hc269bfef, 32'hc2aee63e, 32'h42a0eca0, 32'h42b7acfc, 32'h408511ea};
test_bias[4258:4258] = '{32'hc265e92b};
test_output[4258:4258] = '{32'hc68fcc87};
test_input[34072:34079] = '{32'hc2b7d6f6, 32'hc2ac862f, 32'hc2764be6, 32'hc1a86a52, 32'h42a2d49b, 32'hc26c2271, 32'h41d2a404, 32'h42af6bec};
test_weights[34072:34079] = '{32'hc29a4183, 32'hc1adb099, 32'hc2b2ec18, 32'h42a8fb5c, 32'hc0b01599, 32'h41752512, 32'h4280fedc, 32'h42b5f360};
test_bias[4259:4259] = '{32'hc25314c9};
test_output[4259:4259] = '{32'h46a3c977};
test_input[34080:34087] = '{32'h411a1274, 32'h425337ec, 32'hc1294e07, 32'hc1e6d846, 32'hc26e866b, 32'h4217176f, 32'h42060daa, 32'hc0e3cf4b};
test_weights[34080:34087] = '{32'h41855a96, 32'hc1164690, 32'hc15e74b7, 32'h427c1fa7, 32'h426f6e57, 32'h41184631, 32'hc2c5db5d, 32'hc0614dda};
test_bias[4260:4260] = '{32'hc21b08ec};
test_output[4260:4260] = '{32'hc605888a};
test_input[34088:34095] = '{32'h410102de, 32'hc03579e8, 32'h42b1035d, 32'h42c7b094, 32'h428e5b7a, 32'h40faf28e, 32'h42490ba8, 32'hc1ddf913};
test_weights[34088:34095] = '{32'h429d905c, 32'hc2b1847b, 32'hc2c61ae8, 32'hc188d963, 32'hc22bb946, 32'hc18d6fe6, 32'hc13ee56f, 32'hc2424b92};
test_bias[4261:4261] = '{32'h4209f8d0};
test_output[4261:4261] = '{32'hc63b7eb5};
test_input[34096:34103] = '{32'h427d454a, 32'h427dd06a, 32'hc2b32f67, 32'h41567e53, 32'hc25f4d34, 32'hc22d9ee1, 32'h42c6dd54, 32'hc11544d6};
test_weights[34096:34103] = '{32'hc2b2c051, 32'hc2603db2, 32'hc13b5533, 32'h4298a5ca, 32'hc2892e87, 32'h41d0ceab, 32'hc241e6c3, 32'h428861a4};
test_bias[4262:4262] = '{32'h414e5e11};
test_output[4262:4262] = '{32'hc61a8cd2};
test_input[34104:34111] = '{32'h4253db39, 32'h4202a651, 32'hc2c6a634, 32'hc2aeeefb, 32'h4098c30f, 32'hc28722e8, 32'h4032a0e1, 32'hc26ff823};
test_weights[34104:34111] = '{32'hc1f2eef1, 32'h42a0b46b, 32'hc23c1a57, 32'h42c1cb8d, 32'hc1e6a0af, 32'h42c6dc74, 32'h4294a4e5, 32'h42c0d855};
test_bias[4263:4263] = '{32'hc23304d7};
test_output[4263:4263] = '{32'hc66e88f1};
test_input[34112:34119] = '{32'hc23702d0, 32'h42176d6d, 32'h42b2bc5b, 32'hc0bf1f0d, 32'h4292b859, 32'hc06de858, 32'hc252ebc6, 32'h41d6df22};
test_weights[34112:34119] = '{32'hc0acbccd, 32'hc29d4568, 32'hc0d838bb, 32'h3f8d41be, 32'hc246cac8, 32'h42be4830, 32'h42ae1c0a, 32'h423e9fbd};
test_bias[4264:4264] = '{32'h4282db62};
test_output[4264:4264] = '{32'hc6256387};
test_input[34120:34127] = '{32'h4277e457, 32'h42ae34c6, 32'h427666af, 32'hc1cf19bf, 32'hc2a2aaad, 32'hc15a633b, 32'hc1886748, 32'hc1a794c9};
test_weights[34120:34127] = '{32'hc0ff2b90, 32'hc2b0381d, 32'hc2bbb391, 32'hc2c3d40f, 32'h4245c44d, 32'hc2b5f003, 32'hc1da3f81, 32'h423bcf1f};
test_bias[4265:4265] = '{32'h4289569e};
test_output[4265:4265] = '{32'hc664d259};
test_input[34128:34135] = '{32'hc0f1e47b, 32'hc29caa31, 32'hc2853a1e, 32'h4171359b, 32'h422f03ed, 32'h41efac76, 32'h418b1e1b, 32'hc2a550d7};
test_weights[34128:34135] = '{32'h4188c85a, 32'h4148c9ba, 32'h413a5c10, 32'hc2bdf256, 32'hbe4068a5, 32'h423c5fba, 32'hc1a7a7d1, 32'h41d763c0};
test_bias[4266:4266] = '{32'hc05d87f8};
test_output[4266:4266] = '{32'hc58cf4da};
test_input[34136:34143] = '{32'h4289a267, 32'hc19d4aea, 32'h41246391, 32'hbf0d2fea, 32'h4238cd0d, 32'hc1939633, 32'h425b8c5d, 32'hc1c99223};
test_weights[34136:34143] = '{32'hc14e24b5, 32'hc214bc96, 32'hc2c24f9c, 32'h42a7611e, 32'hbdeee7a8, 32'h42b14fe7, 32'h427e5fc3, 32'h4221e646};
test_bias[4267:4267] = '{32'hc1e8cb78};
test_output[4267:4267] = '{32'hc3c7a6d1};
test_input[34144:34151] = '{32'h42c0a03b, 32'h42aefa26, 32'hc2c0df74, 32'h41ae2dbf, 32'h42c5f358, 32'hc1b3daa4, 32'h414a5b50, 32'h4207cb12};
test_weights[34144:34151] = '{32'h413f198b, 32'hc2b5462f, 32'h42216d03, 32'h42966e99, 32'h41f3e18e, 32'h42069418, 32'hc196375a, 32'hc282a332};
test_bias[4268:4268] = '{32'hc2b1d5ed};
test_output[4268:4268] = '{32'hc6119233};
test_input[34152:34159] = '{32'h416a0461, 32'h42a44726, 32'h4267fe7a, 32'hbf6c3fa0, 32'h42191a29, 32'hc1df7d20, 32'hc20b3a79, 32'h424a092e};
test_weights[34152:34159] = '{32'hc2071b53, 32'h42980f85, 32'hc25f72aa, 32'h42a7782e, 32'hc1e139fc, 32'hc2731016, 32'hc2330d65, 32'h4274154c};
test_bias[4269:4269] = '{32'h421492ad};
test_output[4269:4269] = '{32'h45f1990e};
test_input[34160:34167] = '{32'hc22dc483, 32'hc2ad181c, 32'hc23e63a4, 32'h4264534a, 32'h42b5c06a, 32'hc2c1513b, 32'hc141fd05, 32'h4214febe};
test_weights[34160:34167] = '{32'h42913ecb, 32'hc235a828, 32'hc211b853, 32'hc2a4f98f, 32'hc1aea5bd, 32'hc2c1be8f, 32'hc2ba39e7, 32'h428b0c70};
test_bias[4270:4270] = '{32'h422a3efb};
test_output[4270:4270] = '{32'h460bb796};
test_input[34168:34175] = '{32'h4224ccbe, 32'hc18397ad, 32'h420906d9, 32'h40545d9b, 32'hc28e3b6f, 32'hc21b48c5, 32'h414cd714, 32'h4123bc0e};
test_weights[34168:34175] = '{32'hc22e0249, 32'hc2b1b40e, 32'h41e4a8e7, 32'hc258123b, 32'h42a1d63e, 32'hc28a975c, 32'h412f53ba, 32'h4286c8bd};
test_bias[4271:4271] = '{32'hc268ea28};
test_output[4271:4271] = '{32'hc4e3f407};
test_input[34176:34183] = '{32'h4285c412, 32'h42765466, 32'hc2c71b3e, 32'h40ff3876, 32'h42b3eccf, 32'hc149cda6, 32'h412b75a3, 32'hc2c137eb};
test_weights[34176:34183] = '{32'hc2b0ef8d, 32'hc26582e4, 32'hc190c92a, 32'h42914337, 32'h427fd638, 32'hc2a6f934, 32'hc0ada0eb, 32'h407d70b8};
test_bias[4272:4272] = '{32'h41cbf3ce};
test_output[4272:4272] = '{32'hc4296f53};
test_input[34184:34191] = '{32'hc27624f7, 32'hc2ade10e, 32'h4228bd01, 32'h411cd19f, 32'h429fac1f, 32'hc1b5e613, 32'hc2a6ee19, 32'hc0255d94};
test_weights[34184:34191] = '{32'hc24dd8b8, 32'h41dabd82, 32'h428d983b, 32'hc1c3f141, 32'hc2ad9b3c, 32'hc1634b6b, 32'hc2b1cc65, 32'h427c128b};
test_bias[4273:4273] = '{32'hc28357ba};
test_output[4273:4273] = '{32'h4580c457};
test_input[34192:34199] = '{32'h42bc42b0, 32'h4291897d, 32'hc2b8de2c, 32'h42bc90d1, 32'hc201a1a7, 32'h42b0e100, 32'hc214ab57, 32'h42998722};
test_weights[34192:34199] = '{32'h429f96e7, 32'h4199cedc, 32'h4089daba, 32'hc286935d, 32'hc2bf907a, 32'hc22656ae, 32'hc11f40c4, 32'h4206f871};
test_bias[4274:4274] = '{32'hc0e4aecd};
test_output[4274:4274] = '{32'h458e19ea};
test_input[34200:34207] = '{32'hc2380f8c, 32'h42c73282, 32'hc1e2f2a3, 32'h41e9f20a, 32'h42ba6434, 32'hc12052f2, 32'h42672f39, 32'h429dbc9b};
test_weights[34200:34207] = '{32'h42a3e239, 32'hc25ea6b8, 32'hc2924898, 32'hc2053a0b, 32'hc2b2927e, 32'hc2b553ec, 32'h42502d82, 32'hc27a9634};
test_bias[4275:4275] = '{32'h42845a6b};
test_output[4275:4275] = '{32'hc688a9c7};
test_input[34208:34215] = '{32'h4210a15c, 32'h41c72be5, 32'hc2245e0f, 32'h42aed51d, 32'hc237b8e1, 32'h4294e3c3, 32'h4281011e, 32'hc27aa36f};
test_weights[34208:34215] = '{32'hc29b37aa, 32'hc2a6c08a, 32'hc1759f34, 32'hc28b8bc4, 32'hc16a3526, 32'h41a9b53b, 32'h42b787af, 32'hc284e913};
test_bias[4276:4276] = '{32'hc2935833};
test_output[4276:4276] = '{32'h44eed37f};
test_input[34216:34223] = '{32'h420a1790, 32'h4277b551, 32'hc1449c0c, 32'hc2a4024d, 32'h423d5a23, 32'h40ba28d4, 32'hc25f5c6b, 32'hbf7795da};
test_weights[34216:34223] = '{32'hc2a4aad2, 32'hc2b22c1c, 32'hc2138519, 32'h423c574e, 32'h4290b115, 32'hc2c048cf, 32'hc2c6b5c1, 32'h41586557};
test_bias[4277:4277] = '{32'h41c6b411};
test_output[4277:4277] = '{32'hc550e190};
test_input[34224:34231] = '{32'h4233f780, 32'hc22c3c9d, 32'hc29ed0cb, 32'h4289df72, 32'hc261ff94, 32'hc08de394, 32'hc229b22e, 32'h42bf9df9};
test_weights[34224:34231] = '{32'h40ba9519, 32'hc19d7f82, 32'h41c40273, 32'h4106ea62, 32'h4217018b, 32'hc2b49efb, 32'h42a19762, 32'hc0d12bbd};
test_bias[4278:4278] = '{32'hc1885ca1};
test_output[4278:4278] = '{32'hc5bd4de3};
test_input[34232:34239] = '{32'h429fb2b4, 32'hc23e5381, 32'h41a7eb56, 32'hc222d493, 32'hc2a8535a, 32'hc2b4abe2, 32'h428162b2, 32'hc2a439be};
test_weights[34232:34239] = '{32'hc1e8e9c8, 32'h427542ad, 32'hc101776b, 32'hc2b0b7f9, 32'hc179579b, 32'hc2066f42, 32'hc2c284f5, 32'hc0162568};
test_bias[4279:4279] = '{32'hc288fb8d};
test_output[4279:4279] = '{32'hc56335b7};
test_input[34240:34247] = '{32'h42b0ba7a, 32'hc1444a8e, 32'hc26c7273, 32'h41b71c08, 32'h3fb1312b, 32'h4186a135, 32'hc011e7f2, 32'h4254bade};
test_weights[34240:34247] = '{32'hc298b845, 32'h42aee996, 32'hc213192b, 32'hbe15eac9, 32'hc21b40b5, 32'hc18f1184, 32'hc112d3ef, 32'h4094e438};
test_bias[4280:4280] = '{32'hc2957e85};
test_output[4280:4280] = '{32'hc5b59821};
test_input[34248:34255] = '{32'hc25a6afc, 32'hc2b2a805, 32'hc27d9a6b, 32'h424e309a, 32'hc219c57d, 32'h413b8204, 32'h42b566cd, 32'h409a9a88};
test_weights[34248:34255] = '{32'hc1a8d18b, 32'hc275b38a, 32'h42810a24, 32'hc2a5072c, 32'h42585e70, 32'hc14fc534, 32'hc24acfdf, 32'hc2005b9e};
test_bias[4281:4281] = '{32'hc1a874ad};
test_output[4281:4281] = '{32'hc6081cf4};
test_input[34256:34263] = '{32'h41316222, 32'hc283f4ba, 32'h42493e55, 32'hc2a2f64a, 32'hc20888ce, 32'h4151560d, 32'h424cf505, 32'hc2c67609};
test_weights[34256:34263] = '{32'h41ee89e8, 32'h41ffb833, 32'hc256e0e7, 32'h4224570e, 32'hc23affd1, 32'h429049f4, 32'h423a35b2, 32'hc1a87afc};
test_bias[4282:4282] = '{32'hc20c31c6};
test_output[4282:4282] = '{32'hc454426c};
test_input[34264:34271] = '{32'h41919359, 32'h42738eec, 32'h41be9563, 32'h4245f469, 32'h4077e0cb, 32'hc09174b7, 32'h420a1920, 32'h42c36a52};
test_weights[34264:34271] = '{32'hc19f763a, 32'h4152f7b0, 32'h42a279e8, 32'hc27f638a, 32'hc299edd0, 32'h41df9cc0, 32'h42196f13, 32'hc28305d4};
test_bias[4283:4283] = '{32'h40eedeee};
test_output[4283:4283] = '{32'hc5c4349a};
test_input[34272:34279] = '{32'h4198a654, 32'h42a9c4e3, 32'h42a553d1, 32'hc127bb9a, 32'hc2608dc6, 32'hc2582680, 32'h4248f637, 32'h4127f426};
test_weights[34272:34279] = '{32'hc139a678, 32'h42af44a1, 32'hc12f1ffc, 32'hc2226cca, 32'h42ab4cd7, 32'h4076b413, 32'hc28fd00c, 32'hc2930f07};
test_bias[4284:4284] = '{32'hc2b6ba7c};
test_output[4284:4284] = '{32'hc52c2194};
test_input[34280:34287] = '{32'h414a921f, 32'hc227d47b, 32'h428c4437, 32'hc27465e8, 32'hc1de07c7, 32'h42a8ff5f, 32'hc28d9eae, 32'hc2ad91d5};
test_weights[34280:34287] = '{32'h41b9ceaa, 32'h402f6723, 32'hc230562e, 32'hc28dcc10, 32'hc201259f, 32'hc2adc487, 32'h42c77fdc, 32'h42c59aa4};
test_bias[4285:4285] = '{32'hc200952b};
test_output[4285:4285] = '{32'hc6a1b087};
test_input[34288:34295] = '{32'h40e638e9, 32'h42abada3, 32'h41ccf2ae, 32'hc270beb7, 32'hc0e045f9, 32'hc008caf3, 32'h42939df9, 32'h424ae609};
test_weights[34288:34295] = '{32'h42349b3b, 32'h42c01a47, 32'h42c171f4, 32'h4291c167, 32'hc29a8aef, 32'hc1a0cfcc, 32'hc2ad76fc, 32'hbecb1f4e};
test_bias[4286:4286] = '{32'h420dd215};
test_output[4286:4286] = '{32'h4456ede6};
test_input[34296:34303] = '{32'h4184ee51, 32'h4220be0c, 32'h425c885e, 32'hc15d46a7, 32'h424e863d, 32'hc18dd995, 32'hc2646318, 32'h420dd1ec};
test_weights[34296:34303] = '{32'hc1e62c09, 32'hc0918ab0, 32'hc2854512, 32'hc081e35d, 32'h4207116e, 32'h42457c85, 32'h42a901be, 32'h42167df7};
test_bias[4287:4287] = '{32'h425b5add};
test_output[4287:4287] = '{32'hc5d5f4dc};
test_input[34304:34311] = '{32'hc0de5fe9, 32'hc1fc1e60, 32'hc2248ac4, 32'h411dede6, 32'hc2152a9a, 32'h429460c0, 32'h42bdd248, 32'h41fc73c7};
test_weights[34304:34311] = '{32'h42b56667, 32'h42aaf1a0, 32'hc2ba413d, 32'h42b9920a, 32'hc28c6dd4, 32'h418710f5, 32'h4259ec15, 32'h4252bf65};
test_bias[4288:4288] = '{32'hc29d6405};
test_output[4288:4288] = '{32'h463c41bd};
test_input[34312:34319] = '{32'hc2bfe9ad, 32'h42c54f8e, 32'hc171c87f, 32'h418a5fa9, 32'hc19ac1c7, 32'h4228941d, 32'hc2c4b1be, 32'hc22b5a69};
test_weights[34312:34319] = '{32'h40a10fe2, 32'hc29346a2, 32'hc15684e7, 32'h422974ee, 32'hc28c2f92, 32'h41b6e025, 32'hc1c21d6e, 32'hc288ae21};
test_bias[4289:4289] = '{32'h408d4b50};
test_output[4289:4289] = '{32'h444e50d6};
test_input[34320:34327] = '{32'h42bd3e4f, 32'hc246f948, 32'h42c10d24, 32'h41a82420, 32'hc2b4c118, 32'h426d9213, 32'hc2b5304f, 32'hc2124126};
test_weights[34320:34327] = '{32'hc213f2f6, 32'h4243496a, 32'h428d1391, 32'hc1bafef8, 32'hc29314b4, 32'hc2233105, 32'hc1189d35, 32'h424b9627};
test_bias[4290:4290] = '{32'hbfaafa20};
test_output[4290:4290] = '{32'h4561e37a};
test_input[34328:34335] = '{32'hc1861873, 32'hc20a2d2d, 32'h420eea05, 32'h4006f4b2, 32'h40add016, 32'hc1ed0a0e, 32'hc2c4053b, 32'hc1a67a40};
test_weights[34328:34335] = '{32'hc293f87d, 32'h41ae5537, 32'h42bee823, 32'h422bbed3, 32'hc1e07746, 32'h42b28fcb, 32'h41a61388, 32'hc19c40c7};
test_bias[4291:4291] = '{32'h413c2c86};
test_output[4291:4291] = '{32'hc3d4f46e};
test_input[34336:34343] = '{32'hc1dc8bfd, 32'h42832716, 32'h42356790, 32'hc28ab15d, 32'h429385b8, 32'hc2a20d12, 32'hc232b06e, 32'hc2838a8f};
test_weights[34336:34343] = '{32'hc1463da3, 32'h423e6c04, 32'h4220ac70, 32'h42c1d2d4, 32'h4227a02f, 32'hc1ba5014, 32'hc2c43c97, 32'h41b17c37};
test_bias[4292:4292] = '{32'h42743f37};
test_output[4292:4292] = '{32'h45cbfdb3};
test_input[34344:34351] = '{32'hc19d8902, 32'h42a5a244, 32'hc2469864, 32'h4192be5b, 32'hc24f49be, 32'h428fdb5d, 32'h41827686, 32'h4250c7ae};
test_weights[34344:34351] = '{32'hc20ed905, 32'h405316b6, 32'hc216e06e, 32'h4232f930, 32'h423c7a0f, 32'h423f9edf, 32'hc2697893, 32'h4150fccf};
test_bias[4293:4293] = '{32'hbfabe121};
test_output[4293:4293] = '{32'h45899287};
test_input[34352:34359] = '{32'hc1801daa, 32'h41da8dcd, 32'h42604080, 32'h41e628f7, 32'h42aff2c7, 32'h4213c68b, 32'hc230b782, 32'h42c312ce};
test_weights[34352:34359] = '{32'hc2bef298, 32'h427b6592, 32'h41c87abf, 32'h4244a137, 32'h42a9a10a, 32'h4245066c, 32'h4284b8db, 32'hc27b244c};
test_bias[4294:4294] = '{32'h40e117aa};
test_output[4294:4294] = '{32'h45c4cdcf};
test_input[34360:34367] = '{32'hc22107fb, 32'hc297707c, 32'h42b130bc, 32'h417827e9, 32'hc2aae0e7, 32'hc282faaa, 32'h42b76ad1, 32'hc20e1d4b};
test_weights[34360:34367] = '{32'hc07feb91, 32'h42ad87d9, 32'h4180b306, 32'hc1c78d03, 32'hc224ca5c, 32'hc28cefc3, 32'hc210b518, 32'hc2bb00c8};
test_bias[4295:4295] = '{32'h42347c5b};
test_output[4295:4295] = '{32'h452fdbc2};
test_input[34368:34375] = '{32'hc28bd5ab, 32'h420f13eb, 32'hc2420480, 32'hc24919d7, 32'h422ea853, 32'h4211d290, 32'hc0e81e5f, 32'hc2754e48};
test_weights[34368:34375] = '{32'h4281c3bc, 32'hc25a4888, 32'hc23ed679, 32'h42221326, 32'h429e3667, 32'hc1b33908, 32'h409ab435, 32'h41934a7a};
test_bias[4296:4296] = '{32'hc2b5ee3a};
test_output[4296:4296] = '{32'hc596e871};
test_input[34376:34383] = '{32'h414810cf, 32'h42c15d60, 32'hc01f0793, 32'h42b45c5a, 32'hc2a30b80, 32'hc28f9d2e, 32'hc0e4e1f9, 32'hc28dd7be};
test_weights[34376:34383] = '{32'hc2c26519, 32'h4297f49d, 32'hc2bb7f51, 32'hc245ed0f, 32'h42811657, 32'h41f187d0, 32'hc0d5e6c4, 32'hc11f40e7};
test_bias[4297:4297] = '{32'h42a32255};
test_output[4297:4297] = '{32'hc592ab1a};
test_input[34384:34391] = '{32'hc25d7666, 32'hc1bee44d, 32'h3f85eafc, 32'h406aff9a, 32'hc239130c, 32'hc29b2ad4, 32'h42916235, 32'h425cd052};
test_weights[34384:34391] = '{32'h42039d0d, 32'h41a96c57, 32'h41e02ad8, 32'h3f76762f, 32'hc26aef6d, 32'hc28b5fa2, 32'h401cf48c, 32'hc2855086};
test_bias[4298:4298] = '{32'hc26f8c3e};
test_output[4298:4298] = '{32'h450dc8f8};
test_input[34392:34399] = '{32'h422bf11e, 32'hc25abe9f, 32'h417900b8, 32'hc19901d8, 32'h42252a87, 32'hc2413910, 32'h419436fc, 32'h42a2f3fb};
test_weights[34392:34399] = '{32'hc2b8c86a, 32'h42ac78f6, 32'h42395eec, 32'h41fb9113, 32'h42c48594, 32'hc2766906, 32'h42951ce8, 32'hc29585c9};
test_bias[4299:4299] = '{32'h4089cb1b};
test_output[4299:4299] = '{32'hc5c301c4};
test_input[34400:34407] = '{32'h421bbee6, 32'hc1ca1efc, 32'hc1e5113a, 32'hc1ee77a7, 32'h420388ea, 32'h4290745a, 32'hc21450f1, 32'hc215e58f};
test_weights[34400:34407] = '{32'hc2a213c1, 32'h4211e8a4, 32'hc24f6840, 32'h424b073e, 32'h42bb8649, 32'h41c6db95, 32'h415f974c, 32'h42981321};
test_bias[4300:4300] = '{32'h426113df};
test_output[4300:4300] = '{32'hc51e9f48};
test_input[34408:34415] = '{32'h42aeb9c8, 32'h419c8d4b, 32'h42a8a465, 32'h42baa1ac, 32'hc149512d, 32'h4235bd7a, 32'hc109ff78, 32'h42b250a7};
test_weights[34408:34415] = '{32'hc2a934ce, 32'hc1839ce4, 32'h42bc6578, 32'h42a7838a, 32'hc2a640c6, 32'hc1ec5e35, 32'hc2a69e16, 32'hc2a274b8};
test_bias[4301:4301] = '{32'hbfe72225};
test_output[4301:4301] = '{32'h4498f846};
test_input[34416:34423] = '{32'h427eabf1, 32'h42323d46, 32'hc200ba2e, 32'h411b6dfb, 32'h42498f7c, 32'h42978df0, 32'h42bfcdd5, 32'h41ed34f6};
test_weights[34416:34423] = '{32'hc165761a, 32'h42b8e674, 32'hc19704b5, 32'h41013f5e, 32'h4186564c, 32'h4295bc22, 32'hc27a9dc6, 32'hc1c022f0};
test_bias[4302:4302] = '{32'hc292b914};
test_output[4302:4302] = '{32'h45621b8a};
test_input[34424:34431] = '{32'hc2388d0a, 32'h4268578a, 32'h425c2a6d, 32'hc163a7fd, 32'h42774a5f, 32'h42bcd205, 32'hc2962c81, 32'h42358063};
test_weights[34424:34431] = '{32'h42c46bcf, 32'h415ad663, 32'hc2861873, 32'hc1e03376, 32'h423ee153, 32'h41f0586a, 32'hc29fb318, 32'h429c345e};
test_bias[4303:4303] = '{32'hc2a941dc};
test_output[4303:4303] = '{32'h4600547c};
test_input[34432:34439] = '{32'h420d0767, 32'h42553bba, 32'h42b204e0, 32'hc2a84feb, 32'hc1379c50, 32'h42ab36bc, 32'h41edb633, 32'h41feb81a};
test_weights[34432:34439] = '{32'h4257b6b5, 32'hc19cb917, 32'h42819c72, 32'h42b04fb0, 32'h42195f3e, 32'hc2bb405a, 32'h412ce3d0, 32'h425229f6};
test_bias[4304:4304] = '{32'hc1b77067};
test_output[4304:4304] = '{32'hc5e36ba4};
test_input[34440:34447] = '{32'hc22dc65e, 32'hc2c41f11, 32'hc1ad2acf, 32'h42bc9545, 32'hc292c920, 32'hc131d9e7, 32'h4282710c, 32'h428e4f8a};
test_weights[34440:34447] = '{32'hc273ba65, 32'hc28fe763, 32'hbebe5452, 32'hc2751b0c, 32'h42aa1052, 32'h429d7cd4, 32'h42c1fa02, 32'h421e9bf6};
test_bias[4305:4305] = '{32'h409aab56};
test_output[4305:4305] = '{32'h45ba873f};
test_input[34448:34455] = '{32'h4047d256, 32'h4206f93c, 32'hc26fe18c, 32'h42a515e7, 32'hc1e122fb, 32'h425f288c, 32'h42c53037, 32'hc1c66b49};
test_weights[34448:34455] = '{32'hc26fee8d, 32'h42a17435, 32'h4265e6e2, 32'h3e4b0bdb, 32'hc1293756, 32'h4214bd70, 32'hc20c7df6, 32'hc2aad04b};
test_bias[4306:4306] = '{32'h4234b4e4};
test_output[4306:4306] = '{32'h4332fbc0};
test_input[34456:34463] = '{32'h42b200cc, 32'h418d49de, 32'h42986b70, 32'hc2273321, 32'h428b832f, 32'h428fd3bf, 32'h416e0c45, 32'hc1dd82e7};
test_weights[34456:34463] = '{32'h42b44eff, 32'h3fe780ba, 32'h42321ac9, 32'h42a08c75, 32'h4288f2a3, 32'h421ae7c5, 32'hc27adbb7, 32'hc205896f};
test_bias[4307:4307] = '{32'hc227eb2f};
test_output[4307:4307] = '{32'h4673d1c2};
test_input[34464:34471] = '{32'hc2817a13, 32'h42acc5c0, 32'hc2350107, 32'hc26022e2, 32'hc20fb3ff, 32'hc18041c2, 32'hc2aa5bad, 32'h3e95b396};
test_weights[34464:34471] = '{32'h411b9307, 32'h42484884, 32'hc29ef498, 32'hc2c4f1f5, 32'hc1b296c3, 32'hc12fceb9, 32'hc1a14517, 32'hc1dca703};
test_bias[4308:4308] = '{32'h3fd4b7b8};
test_output[4308:4308] = '{32'h46722c48};
test_input[34472:34479] = '{32'hc2c263ac, 32'hc116418f, 32'h428c9d27, 32'h4243f022, 32'hc2839630, 32'hc256d203, 32'hc2933d8d, 32'hc2945489};
test_weights[34472:34479] = '{32'h414705c6, 32'h420a133a, 32'hc23ebd39, 32'h42aebd86, 32'h4079b9aa, 32'hc2b532ad, 32'h41cd015f, 32'h42ac06e3};
test_bias[4309:4309] = '{32'hc2b2d0e7};
test_output[4309:4309] = '{32'hc58801be};
test_input[34480:34487] = '{32'h428ecc0e, 32'h429188c8, 32'hc230df7f, 32'h4210e60b, 32'h4268fc85, 32'hc2b43b19, 32'hc201fff6, 32'hc20faac1};
test_weights[34480:34487] = '{32'h420bd51c, 32'h42400cbb, 32'hc2b910c8, 32'h40a64b92, 32'hc26c73d2, 32'hc2b8f291, 32'hc0126461, 32'hc2a0f774};
test_bias[4310:4310] = '{32'hc274738f};
test_output[4310:4310] = '{32'h468d1f59};
test_input[34488:34495] = '{32'hc142a7a7, 32'hc1a5980f, 32'h42897c9d, 32'h428784ef, 32'h42ab9739, 32'hc2b15be2, 32'h4248c566, 32'h3fa21cb4};
test_weights[34488:34495] = '{32'h42494243, 32'h421b979f, 32'h41d4e5a8, 32'hc2543e31, 32'h42b1f5ce, 32'h42812ad2, 32'h42c7dffc, 32'h42c57a05};
test_bias[4311:4311] = '{32'h427d2fce};
test_output[4311:4311] = '{32'h45758122};
test_input[34496:34503] = '{32'hc22a46bd, 32'h41931073, 32'hc214d5c7, 32'h428f6c99, 32'h42b8ce08, 32'hc261e450, 32'h41c9a825, 32'h421c15f9};
test_weights[34496:34503] = '{32'hc280ce7e, 32'hc2a2c16c, 32'hc23c76f9, 32'h42a47549, 32'hc2b40711, 32'hc26821b2, 32'h4286af96, 32'hc2c67956};
test_bias[4312:4312] = '{32'hc299edf2};
test_output[4312:4312] = '{32'h44c871ca};
test_input[34504:34511] = '{32'hc16886da, 32'h3ea7bfe2, 32'h424ad007, 32'h4237b23a, 32'hc282cbf6, 32'h4262b7be, 32'h42a6c109, 32'hc25f5ba6};
test_weights[34504:34511] = '{32'hc08506c2, 32'hc13f2635, 32'h41b30a8c, 32'hc2bcbca2, 32'h42970fa1, 32'h41d6a15e, 32'h417c5c40, 32'hc25c271d};
test_bias[4313:4313] = '{32'h428149c2};
test_output[4313:4313] = '{32'hc503c73b};
test_input[34512:34519] = '{32'hc298f44d, 32'h42a2fd21, 32'hc2365680, 32'h425e71fb, 32'hc2bb90be, 32'hc2ba6763, 32'hc271477c, 32'hc23ec8d9};
test_weights[34512:34519] = '{32'h42bb1182, 32'hc28075fd, 32'h42971634, 32'hc1b92727, 32'hc182581c, 32'hc2acbda7, 32'hbebde943, 32'h429d97e8};
test_bias[4314:4314] = '{32'hc20b32b4};
test_output[4314:4314] = '{32'hc630bca4};
test_input[34520:34527] = '{32'h40c9b213, 32'hc200d97b, 32'h427c47b8, 32'h4225b4fe, 32'h42abbc64, 32'h427d4852, 32'hc2b031c9, 32'h40eeed8a};
test_weights[34520:34527] = '{32'h423a6f7e, 32'hc2a2ddbc, 32'hc20973ec, 32'hc18d6d20, 32'h42023d52, 32'h42265fa8, 32'h4021cbc1, 32'hc282a8b0};
test_bias[4315:4315] = '{32'h42aa34c8};
test_output[4315:4315] = '{32'h4596abb4};
test_input[34528:34535] = '{32'hc2c6c52a, 32'h428b1629, 32'h42a0cd32, 32'h429dfcf2, 32'hc29d86c1, 32'hc2724919, 32'hc2899e55, 32'hc278b495};
test_weights[34528:34535] = '{32'hc29c38f9, 32'h4299c5f9, 32'h422b812b, 32'h42a8fac0, 32'hc262e17c, 32'h4267a51a, 32'hc2a19013, 32'hc17bfc9c};
test_bias[4316:4316] = '{32'h41b6df6e};
test_output[4316:4316] = '{32'h46f03f99};
test_input[34536:34543] = '{32'hc2c5c600, 32'hc279d2e1, 32'h4293f136, 32'hc271a5df, 32'hc1ff9b76, 32'hc29fe808, 32'hbec516bb, 32'h424c144d};
test_weights[34536:34543] = '{32'hc26a85ca, 32'h42a74a66, 32'h422f768d, 32'h420be2bd, 32'hc21b37fc, 32'hc2aa9b35, 32'hc1b35dd8, 32'hc235df7f};
test_bias[4317:4317] = '{32'hc2a055a1};
test_output[4317:4317] = '{32'h45e6744c};
test_input[34544:34551] = '{32'hc28cfc1a, 32'h42724646, 32'h42a21e11, 32'h4279b44c, 32'hc2202d8b, 32'h428eb286, 32'h42b24db4, 32'hc2614de5};
test_weights[34544:34551] = '{32'hc1d15a87, 32'h41b36724, 32'h423b3de3, 32'h3f7f2bd9, 32'h423d59c5, 32'hc10dccb4, 32'h4287fad3, 32'hc2175de6};
test_bias[4318:4318] = '{32'h4220d1ad};
test_output[4318:4318] = '{32'h46477320};
test_input[34552:34559] = '{32'hc2a9f832, 32'hc1d349f4, 32'h42a113e5, 32'hc175aea6, 32'h428f72be, 32'hc227f58c, 32'hc10a325f, 32'h423c7a19};
test_weights[34552:34559] = '{32'h424588db, 32'hc2614d6e, 32'h3f4a2c7a, 32'h4278be73, 32'hc1eb5793, 32'hc24a0991, 32'h428834fb, 32'hc2c77686};
test_bias[4319:4319] = '{32'h4278ff84};
test_output[4319:4319] = '{32'hc609bb5f};
test_input[34560:34567] = '{32'hc2403871, 32'hc26d1a31, 32'hbfe75dd6, 32'hc2778017, 32'h420348d8, 32'h42aabe98, 32'hc29bbba6, 32'hc1d96c89};
test_weights[34560:34567] = '{32'h42021bb6, 32'hc28fa4ca, 32'h41212d47, 32'hc2c3e600, 32'hc18a2a8d, 32'h425f2cd4, 32'h4264aabd, 32'h420b02e7};
test_bias[4320:4320] = '{32'h40d22bbb};
test_output[4320:4320] = '{32'h45ebbd64};
test_input[34568:34575] = '{32'hc2a2d3de, 32'hc1fea93e, 32'h4048789f, 32'hc1d0ff10, 32'hc2959e89, 32'hc111bf3c, 32'h40f5b6fc, 32'hc0ce1705};
test_weights[34568:34575] = '{32'h42916a1d, 32'hc223b7e4, 32'hc2bbdd85, 32'hbfcd1506, 32'hc2a04785, 32'hc2a69c24, 32'h40652a4e, 32'hc1570506};
test_bias[4321:4321] = '{32'h420c98f4};
test_output[4321:4321] = '{32'h44fe4ce7};
test_input[34576:34583] = '{32'hc1533cce, 32'h42affaf3, 32'h42a56288, 32'hc236972a, 32'h4049f5f0, 32'h42a6ddf3, 32'h42558389, 32'h414f1282};
test_weights[34576:34583] = '{32'h42c2077d, 32'h41a0519c, 32'h42ae442f, 32'h401bd311, 32'hc24c2b09, 32'h42af65fd, 32'hc264be5f, 32'h4254a0e7};
test_bias[4322:4322] = '{32'h423c9047};
test_output[4322:4322] = '{32'h4641fcc2};
test_input[34584:34591] = '{32'hc2b6df02, 32'h415c14a4, 32'hc29fcc1e, 32'hc29221f6, 32'h4123344a, 32'hc227df2d, 32'h4289771d, 32'h42458e66};
test_weights[34584:34591] = '{32'hc1143820, 32'h422f8f21, 32'h422ea80a, 32'hc2912b45, 32'hc06b1bce, 32'h413b497f, 32'h42854f0b, 32'hc1cdc888};
test_bias[4323:4323] = '{32'h427036a4};
test_output[4323:4323] = '{32'h45beddfa};
test_input[34592:34599] = '{32'h428c43cb, 32'h428c3764, 32'hc210b8c6, 32'h4212403d, 32'hc19977f9, 32'hc2b14990, 32'hc218971c, 32'h41903f61};
test_weights[34592:34599] = '{32'hc117273b, 32'hc13cb50b, 32'hc21ea40e, 32'hc25b73dc, 32'h429fb62d, 32'h42827466, 32'h42bd98ce, 32'h418516ea};
test_bias[4324:4324] = '{32'h41d7456f};
test_output[4324:4324] = '{32'hc645df38};
test_input[34600:34607] = '{32'hc25d69bd, 32'h4206ed18, 32'h42813b70, 32'h426d59db, 32'h42c2266b, 32'h42894024, 32'hc1b856e1, 32'hc2765e87};
test_weights[34600:34607] = '{32'hc24c2c26, 32'h42b27b14, 32'hc1918c7c, 32'h42a1e2c5, 32'h3f0c4ba3, 32'hc2b89f76, 32'hc26cf846, 32'hc2b9983d};
test_bias[4325:4325] = '{32'hc2529a79};
test_output[4325:4325] = '{32'h461f8554};
test_input[34608:34615] = '{32'h42355760, 32'hc2aacb2b, 32'hc1e0b976, 32'hc2aaa23e, 32'h421ac846, 32'hc0b77cc0, 32'hc281b971, 32'h4243362f};
test_weights[34608:34615] = '{32'hc2736915, 32'h42920a3d, 32'hc22fe140, 32'hc110be55, 32'hc272926b, 32'h427210d4, 32'hc0ae6f7a, 32'h41cfccb3};
test_bias[4326:4326] = '{32'hc1f83920};
test_output[4326:4326] = '{32'hc5fcd748};
test_input[34616:34623] = '{32'hc2c29d57, 32'h4286fa9b, 32'hc20a154f, 32'hc024c5a5, 32'hc1ed6c4f, 32'h405d2223, 32'h424dbf37, 32'hc25e5647};
test_weights[34616:34623] = '{32'hc2977a2a, 32'h42a9d898, 32'h4282c01e, 32'hc1b092a3, 32'hc0911cce, 32'hc262c76d, 32'hc2099c15, 32'h41f211f1};
test_bias[4327:4327] = '{32'hc232f1d1};
test_output[4327:4327] = '{32'h45e57ebf};
test_input[34624:34631] = '{32'hc27d2e3e, 32'h412eebde, 32'hc2a0fafb, 32'hc2265ccc, 32'hc246ae96, 32'h42319f43, 32'hc2321e5b, 32'h423350a4};
test_weights[34624:34631] = '{32'h42bb038f, 32'hc1cd5472, 32'hc2a991e7, 32'hc2b355a1, 32'h42af7a1d, 32'h42b998b6, 32'hc2051950, 32'hc2946da3};
test_bias[4328:4328] = '{32'h42247821};
test_output[4328:4328] = '{32'h451092eb};
test_input[34632:34639] = '{32'hc2153235, 32'hc154a77f, 32'hc042b32b, 32'h40ac4876, 32'hc2077a00, 32'h4262e650, 32'h40461712, 32'hc281f343};
test_weights[34632:34639] = '{32'h3ea16f95, 32'hc07da46d, 32'hc23312f1, 32'h427013ad, 32'h4257f59d, 32'hc1cc00ac, 32'h40b83355, 32'hc185619d};
test_bias[4329:4329] = '{32'hc2aacdd3};
test_output[4329:4329] = '{32'hc4dbe426};
test_input[34640:34647] = '{32'h42b56625, 32'hc21cd592, 32'hc191c170, 32'h42c1588f, 32'hc2970266, 32'hc1464db2, 32'hc2c42920, 32'h42c7ae35};
test_weights[34640:34647] = '{32'hc2c4c848, 32'h426f6146, 32'hc028da8c, 32'h42a250ed, 32'hc18d9ee6, 32'h40487699, 32'hc24ac0cb, 32'h4292ee51};
test_bias[4330:4330] = '{32'hc21d186f};
test_output[4330:4330] = '{32'h461f3109};
test_input[34648:34655] = '{32'hc288d410, 32'hc298eb2a, 32'h423bbfca, 32'hc2902153, 32'hc2926222, 32'hc2096e15, 32'h41b257c9, 32'hc2bd0ba6};
test_weights[34648:34655] = '{32'hc28b61bf, 32'h3fe205e9, 32'h42bfb464, 32'hc2adfb37, 32'hc1eb961b, 32'hc235c1be, 32'h42141667, 32'hc2b67a93};
test_bias[4331:4331] = '{32'h42538548};
test_output[4331:4331] = '{32'h46df97a5};
test_input[34656:34663] = '{32'hc2234529, 32'h42b25db7, 32'h427e354e, 32'h425b61ab, 32'h423e7948, 32'h4139c7fd, 32'hc290cd2b, 32'hc2b8e21a};
test_weights[34656:34663] = '{32'hc2a34a71, 32'hc26aafc5, 32'h4244552e, 32'h426985ec, 32'hc20a1851, 32'hc224dc22, 32'h4210510b, 32'hc2a4231a};
test_bias[4332:4332] = '{32'hc2b07f79};
test_output[4332:4332] = '{32'h45e08758};
test_input[34664:34671] = '{32'hc2a63d79, 32'hc24bb6c0, 32'hc2aec4d1, 32'hc1b34bc7, 32'hc22a2fd2, 32'hc2a250b7, 32'hc152fa65, 32'hc1afea2e};
test_weights[34664:34671] = '{32'hc0eb3048, 32'hc2691580, 32'hc24d6f86, 32'h42735dc7, 32'hc2b9a7af, 32'hc15d824f, 32'h418cf8c1, 32'h42bd7450};
test_bias[4333:4333] = '{32'hc2961312};
test_output[4333:4333] = '{32'h4612a688};
test_input[34672:34679] = '{32'h42976db3, 32'hc20b5d5b, 32'hc207d1b3, 32'h428c6b29, 32'h42106063, 32'h4285b37a, 32'hc21f8d69, 32'h4293adab};
test_weights[34672:34679] = '{32'h429d54aa, 32'h4205df91, 32'h4181c3e6, 32'h428d9747, 32'h42bfdfb2, 32'h42a523fb, 32'h410c164f, 32'h414eb998};
test_bias[4334:4334] = '{32'hc1eaa380};
test_output[4334:4334] = '{32'h46929fa9};
test_input[34680:34687] = '{32'h42c7fa5a, 32'h429bff07, 32'hc0c9bfc3, 32'h41100d80, 32'hc2ae35f0, 32'h42bc6b05, 32'hc28e142d, 32'hc2b1e268};
test_weights[34680:34687] = '{32'h42add2f0, 32'h42045824, 32'h427e9cd8, 32'h428e2380, 32'h42151515, 32'hc1279666, 32'h420d6284, 32'hc18c2dad};
test_bias[4335:4335] = '{32'hc1893c05};
test_output[4335:4335] = '{32'h45c51463};
test_input[34688:34695] = '{32'h42b21805, 32'h42613d73, 32'hc264da34, 32'hc255f8b7, 32'hc27247e9, 32'hc1ca3a3b, 32'hc2b66705, 32'hc2afcfee};
test_weights[34688:34695] = '{32'h41de185c, 32'hc2c089ec, 32'hc09dd5e4, 32'h40e389c2, 32'hc23de484, 32'h41c17efa, 32'hc28b0342, 32'hc1613989};
test_bias[4336:4336] = '{32'hc270e2a1};
test_output[4336:4336] = '{32'h45d26a91};
test_input[34696:34703] = '{32'hc2b3490a, 32'h4210ec1a, 32'hc2af6c2b, 32'h4235857d, 32'h41e2707d, 32'hc25a1e9e, 32'hc1aee813, 32'h42ad2902};
test_weights[34696:34703] = '{32'hc293e7dd, 32'h427849c0, 32'hc18af298, 32'h4157cf07, 32'h4212e576, 32'hc2b45ae9, 32'hc21d64c6, 32'h41987a17};
test_bias[4337:4337] = '{32'hc292e720};
test_output[4337:4337] = '{32'h46979f34};
test_input[34704:34711] = '{32'hc2aee9f6, 32'hbf6caf7f, 32'h41adadbd, 32'h42489f8e, 32'h420dfc38, 32'hc29f2f92, 32'h4217c774, 32'hc200350a};
test_weights[34704:34711] = '{32'h41e346a3, 32'hc26479fc, 32'hc245e46a, 32'hc2b445ae, 32'h42817a25, 32'h422e678b, 32'h41732a8b, 32'h42c52431};
test_bias[4338:4338] = '{32'hc0aebb87};
test_output[4338:4338] = '{32'hc6382cd4};
test_input[34712:34719] = '{32'h42a43abb, 32'hc12cbd81, 32'hc235cba4, 32'h42029777, 32'h42ac4ab0, 32'h429112bb, 32'h41a5f244, 32'h40dbb7da};
test_weights[34712:34719] = '{32'hc18e52e3, 32'hc2a92fef, 32'hc2845786, 32'h4171bd04, 32'h4238b6e8, 32'h42192a54, 32'hc0e640ab, 32'hc285a1bf};
test_bias[4339:4339] = '{32'hc102d6dd};
test_output[4339:4339] = '{32'h460e120c};
test_input[34720:34727] = '{32'hc1f2476d, 32'h4187aed7, 32'hc20360c2, 32'h41df5408, 32'hc2becb17, 32'h42b985ee, 32'h424808e5, 32'h41d20981};
test_weights[34720:34727] = '{32'h429151e6, 32'hc0b1f476, 32'hc27ddab0, 32'hc2a9fca4, 32'hc2547d09, 32'h42a66fa1, 32'hc1d924d3, 32'h42865370};
test_bias[4340:4340] = '{32'h42329a0d};
test_output[4340:4340] = '{32'h46267a94};
test_input[34728:34735] = '{32'hc1f33a12, 32'hc222e099, 32'hc2a2dfa0, 32'hc1c15f90, 32'h41cf85cf, 32'h429a5cf8, 32'h42a2f9a8, 32'h4289dde3};
test_weights[34728:34735] = '{32'hc280baf0, 32'hc2c1d587, 32'h42341833, 32'h42affe4f, 32'h428d8660, 32'hc230e4e0, 32'hc1d7a9ca, 32'h42707414};
test_bias[4341:4341] = '{32'hc24de6eb};
test_output[4341:4341] = '{32'h43d5d653};
test_input[34736:34743] = '{32'hc29ab58b, 32'hc130547a, 32'h426f911f, 32'hc2bb6ede, 32'h42a95fb6, 32'hc19e0abf, 32'h422a3163, 32'h41ed6152};
test_weights[34736:34743] = '{32'hc2190c78, 32'h41215bd5, 32'hc29f614b, 32'h4296fc7a, 32'hc2a2fe70, 32'hc24c2d3e, 32'h41dda5af, 32'h421c33e4};
test_bias[4342:4342] = '{32'h421bcf67};
test_output[4342:4342] = '{32'hc6438fb7};
test_input[34744:34751] = '{32'h4287161b, 32'hc283adc7, 32'h42c57e5e, 32'hc1145554, 32'hc24e10d9, 32'hc0f97a8d, 32'hc22222d3, 32'h4244e537};
test_weights[34744:34751] = '{32'hc2aa2db1, 32'h42870984, 32'hc2854d9b, 32'h42ab1d2a, 32'hc27f5a27, 32'h4282175d, 32'h4295231c, 32'hc296d918};
test_bias[4343:4343] = '{32'h428bf5a6};
test_output[4343:4343] = '{32'hc6a79614};
test_input[34752:34759] = '{32'h42bdff20, 32'h41e2a0ec, 32'hc21aafec, 32'hc139e026, 32'h41b85af5, 32'h425dd2ff, 32'hc274a3ba, 32'h424195e4};
test_weights[34752:34759] = '{32'hc095647e, 32'hc2b0cc70, 32'h421dc761, 32'h41f5210d, 32'hc189858b, 32'h42c0be1f, 32'h416535ef, 32'h424c5081};
test_bias[4344:4344] = '{32'hc0c15693};
test_output[4344:4344] = '{32'h44d59ef8};
test_input[34760:34767] = '{32'hc25de142, 32'hc2a6ffe7, 32'hc2aa8270, 32'hc2a0128e, 32'h4175eb27, 32'hc274e570, 32'h423774a0, 32'h4194d680};
test_weights[34760:34767] = '{32'h4297c962, 32'hc2aa52a8, 32'h42bb30f8, 32'hc27347c9, 32'hc272763b, 32'h42a64175, 32'h421f024f, 32'hc1275d61};
test_bias[4345:4345] = '{32'h422e2c46};
test_output[4345:4345] = '{32'hc58e7b9e};
test_input[34768:34775] = '{32'h41650f8f, 32'hc2080901, 32'h42ab4590, 32'hc1f4cfca, 32'h42a0e898, 32'hc271c4c8, 32'hc209af89, 32'hc2750ce3};
test_weights[34768:34775] = '{32'h411e21ec, 32'hc2452518, 32'h424c3194, 32'h3ecbb1c8, 32'hc28fe91f, 32'hc27c93a9, 32'hc2af6790, 32'hc28068ed};
test_bias[4346:4346] = '{32'hc20debfa};
test_output[4346:4346] = '{32'h462dc4ef};
test_input[34776:34783] = '{32'hc1577550, 32'hc286bcae, 32'hc2a374f9, 32'h424b754e, 32'hbf6f4211, 32'h41319a70, 32'hc2a9c7a2, 32'hc170b722};
test_weights[34776:34783] = '{32'hc2687b1b, 32'hc22adfb3, 32'hc228ab90, 32'hc0a3d7d4, 32'hc248ad75, 32'hc2b55d57, 32'hc0785c4a, 32'h4247525d};
test_bias[4347:4347] = '{32'h4201e7c5};
test_output[4347:4347] = '{32'h45abd73f};
test_input[34784:34791] = '{32'hc2bf5adc, 32'hc2782b59, 32'h42a308a2, 32'hc2968137, 32'hc27e2d5b, 32'hc2abf015, 32'h42c4b025, 32'hc1dcb8ee};
test_weights[34784:34791] = '{32'h427fd854, 32'hc227c26b, 32'h42204a4b, 32'h41d7296c, 32'hc2994718, 32'h412f79f8, 32'h40ec0c37, 32'h429e1e04};
test_bias[4348:4348] = '{32'hc1411d4d};
test_output[4348:4348] = '{32'h433848e0};
test_input[34792:34799] = '{32'hc1997f86, 32'h42547b2d, 32'h42600068, 32'hc23b1bfc, 32'hc106230f, 32'hc287384d, 32'hc2073f39, 32'hc2a13dc8};
test_weights[34792:34799] = '{32'hc19d8119, 32'h42bae9b0, 32'hc16b8e00, 32'hc162915b, 32'h429c2bc2, 32'hc2af0cae, 32'h42a5df65, 32'h426d4bca};
test_bias[4349:4349] = '{32'hc195d1b6};
test_output[4349:4349] = '{32'h453155b1};
test_input[34800:34807] = '{32'h42b472ba, 32'h409d052e, 32'h42bd556d, 32'hc2be1f26, 32'h426ea591, 32'hc231bb78, 32'hc247e2ce, 32'h42c62c25};
test_weights[34800:34807] = '{32'h421d1470, 32'h429fc139, 32'h42220d7f, 32'hc11424ba, 32'hc1b3bbf6, 32'hc2580650, 32'h42b7e675, 32'h423ab4e8};
test_bias[4350:4350] = '{32'hc2694d68};
test_output[4350:4350] = '{32'h46174618};
test_input[34808:34815] = '{32'h42171273, 32'hc241d18d, 32'hc224c8ee, 32'h4285ced8, 32'h4293087c, 32'hc222a5ac, 32'hc19f6ac8, 32'hc23db7a4};
test_weights[34808:34815] = '{32'hc2487a9a, 32'hc28b392d, 32'h42521943, 32'h428960dc, 32'h40e17743, 32'h41eac73f, 32'hc144641a, 32'h42c64771};
test_bias[4351:4351] = '{32'hc1fb7b33};
test_output[4351:4351] = '{32'hc49c8e3a};
test_input[34816:34823] = '{32'hc2047978, 32'hc295aad3, 32'h42041df5, 32'hc2bf046f, 32'h423824fc, 32'hc2ba26bf, 32'h425658a8, 32'hc2813597};
test_weights[34816:34823] = '{32'h4245d690, 32'h42bca46d, 32'h42c6d11b, 32'h40ca8a46, 32'hc122cbc8, 32'hc26b7238, 32'h418d65f0, 32'h40539f8d};
test_bias[4352:4352] = '{32'hc2a61eb5};
test_output[4352:4352] = '{32'hc3b27736};
test_input[34824:34831] = '{32'h417de4cb, 32'h423166dc, 32'h42a40cee, 32'h4234f45d, 32'h429a7bb5, 32'h416b5885, 32'hc1af2642, 32'hc2693d9d};
test_weights[34824:34831] = '{32'h42c4e282, 32'h42645a2d, 32'h40837982, 32'h41adbc5b, 32'h42b24935, 32'h42915bfe, 32'h41d4b656, 32'hc1879d80};
test_bias[4353:4353] = '{32'hc21fa82d};
test_output[4353:4353] = '{32'h465699e9};
test_input[34832:34839] = '{32'hc1b2c8df, 32'hc180d89e, 32'h428b709d, 32'hc1ffed93, 32'h422d23d4, 32'hc03d7519, 32'hc2337ed4, 32'h411e51ab};
test_weights[34832:34839] = '{32'hc2c60f0e, 32'hc18b44c2, 32'hc298754e, 32'hc1be26ac, 32'hc2b4f765, 32'h42814ad7, 32'hc273f786, 32'h42a4be68};
test_bias[4354:4354] = '{32'hc0d8bee9};
test_output[4354:4354] = '{32'hc523f834};
test_input[34840:34847] = '{32'hc1dc2054, 32'hc24daaa2, 32'h428704a0, 32'hc296a1c9, 32'h429c2792, 32'hc146323d, 32'hc2b0bf95, 32'h424431dc};
test_weights[34840:34847] = '{32'hc06d3379, 32'hc1863c15, 32'h42bf218e, 32'hc13ab3ed, 32'hc2b2d305, 32'h4299236a, 32'h422029f2, 32'hbf9da629};
test_bias[4355:4355] = '{32'h41776b18};
test_output[4355:4355] = '{32'hc5491f67};
test_input[34848:34855] = '{32'h428563e0, 32'hc298dca3, 32'h423137ca, 32'hc2c31034, 32'hc23a00be, 32'h4200eea5, 32'hc20048d4, 32'h4253eb94};
test_weights[34848:34855] = '{32'hc284f477, 32'h410da4fc, 32'hc28be308, 32'hc1c25776, 32'h42937733, 32'hc209bdd8, 32'hc2c2a201, 32'hc24a3bfe};
test_bias[4356:4356] = '{32'hc165e93a};
test_output[4356:4356] = '{32'hc61b7969};
test_input[34856:34863] = '{32'hc2422878, 32'h429a7043, 32'hc268270b, 32'hc298bbf9, 32'hc0f95fbe, 32'h42237012, 32'h42a73da8, 32'h42357b7f};
test_weights[34856:34863] = '{32'hc259c9df, 32'h425afe15, 32'h411c3e8d, 32'h41941c03, 32'hc25bd106, 32'hc2679de5, 32'h425d04e9, 32'h42811274};
test_bias[4357:4357] = '{32'h41699177};
test_output[4357:4357] = '{32'h46244cf6};
test_input[34864:34871] = '{32'hc169a9b7, 32'h4292817f, 32'h4217b98c, 32'hc1b6eed4, 32'h41ef4b1d, 32'hc26e3122, 32'h3fe4e987, 32'h4278ed2a};
test_weights[34864:34871] = '{32'h4078feae, 32'hc23a47d4, 32'h42066c84, 32'h4224c4aa, 32'hc22aadfd, 32'hc2b79828, 32'h41666a9c, 32'hc1e4c201};
test_bias[4358:4358] = '{32'h42aed554};
test_output[4358:4358] = '{32'hc418ef76};
test_input[34872:34879] = '{32'hc2babe6e, 32'h4255b7d0, 32'h428adb3f, 32'hc11264f4, 32'h4225d093, 32'hc20226fb, 32'h422b80d7, 32'hc2844952};
test_weights[34872:34879] = '{32'h408e97e3, 32'hc25df61b, 32'h41e2c5e3, 32'h418049a8, 32'hbe336a22, 32'hc22762c1, 32'hc190076d, 32'h42bb531a};
test_bias[4359:4359] = '{32'h42394d44};
test_output[4359:4359] = '{32'hc5deaf84};
test_input[34880:34887] = '{32'hc28377f2, 32'h415563a1, 32'h41a171f6, 32'h42470137, 32'h415ee19b, 32'h42c6c3c2, 32'h414a0d38, 32'h424507cd};
test_weights[34880:34887] = '{32'hc15c6306, 32'h41b31f50, 32'h412c834b, 32'hc28c68e3, 32'hc1e4aaf7, 32'hc26cf872, 32'h42b0a57c, 32'hc2c7d7c7};
test_bias[4360:4360] = '{32'hc2c491b8};
test_output[4360:4360] = '{32'hc63f9726};
test_input[34888:34895] = '{32'hbccc680d, 32'h41855691, 32'hc2c7ec35, 32'hc2a9736f, 32'hc2560bca, 32'hc19c5af8, 32'h42b85be3, 32'hc2b8248a};
test_weights[34888:34895] = '{32'h4274ffd7, 32'h42801adf, 32'hc138129a, 32'h421f05de, 32'hc1e47988, 32'h4229820c, 32'hc158b1ee, 32'h4245b468};
test_bias[4361:4361] = '{32'h42aec17c};
test_output[4361:4361] = '{32'hc5c0a036};
test_input[34896:34903] = '{32'h423557c6, 32'h4276bc5d, 32'h419c273e, 32'hc29689bd, 32'h4076883a, 32'h425a3885, 32'h428e002a, 32'h429d2a3f};
test_weights[34896:34903] = '{32'hc202997f, 32'hc27bfaf0, 32'hc28b4f67, 32'h40c6ec06, 32'h42b94859, 32'hc2af1d0a, 32'hc1e0394d, 32'hc2bf6515};
test_bias[4362:4362] = '{32'h4265f2e8};
test_output[4362:4362] = '{32'hc6a493ec};
test_input[34904:34911] = '{32'h42b53d95, 32'h41e1029b, 32'h404781f1, 32'hc20a5342, 32'h421b02a4, 32'h42203609, 32'hc126bf26, 32'hc18369a4};
test_weights[34904:34911] = '{32'hc275ea36, 32'hc1be8635, 32'h42568f96, 32'hc0ad0d7b, 32'h427cdff1, 32'hc211fb5e, 32'hc1fbad3e, 32'h4219cd5e};
test_bias[4363:4363] = '{32'hc2a9014d};
test_output[4363:4363] = '{32'hc5a53790};
test_input[34912:34919] = '{32'h42818652, 32'hc1e9a284, 32'hc08a54f1, 32'h42846e7a, 32'hc17bb04c, 32'hc2c2b63c, 32'hc24d4599, 32'h41208a2a};
test_weights[34912:34919] = '{32'hc29ad38b, 32'h3e36e8d1, 32'hc22c4cee, 32'h42717ac4, 32'h42a31e8f, 32'h42346bae, 32'h42b1f6bc, 32'h429ac1dc};
test_bias[4364:4364] = '{32'hc2495a96};
test_output[4364:4364] = '{32'hc621b64a};
test_input[34920:34927] = '{32'hc2a09107, 32'hc2a6938a, 32'hc205ec7c, 32'h4216e6f5, 32'h421ae8c0, 32'hc26f05ea, 32'hc215e418, 32'h42c4058f};
test_weights[34920:34927] = '{32'hc2a5741e, 32'h42024761, 32'h42827c72, 32'h40ca0048, 32'hc29fd334, 32'hc1788ed1, 32'hc046201c, 32'h4291a338};
test_bias[4365:4365] = '{32'h40afb625};
test_output[4365:4365] = '{32'h45dd1572};
test_input[34928:34935] = '{32'h41788c22, 32'hc25cccd3, 32'hc1bf557f, 32'h41c805d5, 32'h4236861b, 32'hc236c46c, 32'hc2344f53, 32'h4265e0c4};
test_weights[34928:34935] = '{32'h41649aae, 32'hc20bc9e7, 32'h422bdf8b, 32'hc1d0b220, 32'h413a9654, 32'hc2019c19, 32'h427ed186, 32'h421ba9b4};
test_bias[4366:4366] = '{32'hc28cd317};
test_output[4366:4366] = '{32'h44de464b};
test_input[34936:34943] = '{32'h42aeda7c, 32'h41fc0fa8, 32'h42246669, 32'h42273a04, 32'hc0f951f4, 32'h40af9f8b, 32'hc291b42d, 32'h415a55d1};
test_weights[34936:34943] = '{32'h428fc33d, 32'h42aacf5e, 32'h427458fa, 32'h40952d64, 32'h3f33cb06, 32'h4272cfbf, 32'h42822174, 32'h418a2c22};
test_bias[4367:4367] = '{32'h418f9d2b};
test_output[4367:4367] = '{32'h45eb1014};
test_input[34944:34951] = '{32'h428d451f, 32'hc2764143, 32'h40ff68f0, 32'hc1e44668, 32'h423aea99, 32'h4292b467, 32'hc26b9ee9, 32'hc27e9496};
test_weights[34944:34951] = '{32'h42893574, 32'hc1eff50a, 32'h427b1ddf, 32'h420914e7, 32'h42678c6c, 32'hc25d5c5e, 32'h41dc038a, 32'h42c6f70c};
test_bias[4368:4368] = '{32'h4292d9e2};
test_output[4368:4368] = '{32'hc53c8d1c};
test_input[34952:34959] = '{32'hc2c175e7, 32'hc2acdc49, 32'hc22496e7, 32'hc0337696, 32'hc1e92a41, 32'hc2ad911b, 32'h420933e0, 32'hc299ad6c};
test_weights[34952:34959] = '{32'hc12a8191, 32'hc29b2219, 32'hc2617c27, 32'hc2b9d93b, 32'h429ee213, 32'hc2941d72, 32'h424a752e, 32'h42822c7e};
test_bias[4369:4369] = '{32'hc2a549bd};
test_output[4369:4369] = '{32'h462d1b83};
test_input[34960:34967] = '{32'h42788ccb, 32'hc28a6c43, 32'hc296532b, 32'h420429ed, 32'hc1dc54aa, 32'h40da1585, 32'hc1db6a07, 32'hc1e91f5f};
test_weights[34960:34967] = '{32'hc1937872, 32'hc251703a, 32'hc246be9a, 32'hc27e4086, 32'h42af918c, 32'hc28e8d4e, 32'hc2ba44bc, 32'hc248f1be};
test_bias[4370:4370] = '{32'hc2af6f69};
test_output[4370:4370] = '{32'h45a09f33};
test_input[34968:34975] = '{32'h42154277, 32'hc1a2c0e7, 32'hc1f91f8a, 32'hc28bfb9b, 32'h42845aaa, 32'h41ce5f31, 32'h419c3a1c, 32'h41209159};
test_weights[34968:34975] = '{32'h420a3a5b, 32'hc2994e7d, 32'hc260be31, 32'hc2a89e3d, 32'hc2934e90, 32'hbf318fe1, 32'h42b5f49b, 32'h4270f55a};
test_bias[4371:4371] = '{32'h42487b75};
test_output[4371:4371] = '{32'h45fb35e3};
test_input[34976:34983] = '{32'hc2970279, 32'hc2bce403, 32'hc2a79549, 32'h41b32363, 32'hc22f0503, 32'hc29a357a, 32'hc28edc23, 32'hc294df88};
test_weights[34976:34983] = '{32'hc18ee96e, 32'hc17c671c, 32'hc2ba7f9f, 32'hc2c608bf, 32'h426d17e1, 32'hc2c1d0d6, 32'h42084115, 32'h41d5ec3d};
test_bias[4372:4372] = '{32'h429c49b2};
test_output[4372:4372] = '{32'h460c2032};
test_input[34984:34991] = '{32'h427f3c9c, 32'h42814054, 32'h41e5dbbc, 32'hc1483e5f, 32'h42af57bf, 32'h420df34c, 32'hc2b89a0b, 32'h4270b6f3};
test_weights[34984:34991] = '{32'h423d1e2b, 32'h422c07d6, 32'h41c02e69, 32'hc2407087, 32'h4180d2cf, 32'hc2578337, 32'h42c1d01c, 32'hc28a451c};
test_bias[4373:4373] = '{32'h42add199};
test_output[4373:4373] = '{32'hc5c8ede5};
test_input[34992:34999] = '{32'hc290936e, 32'hc21e61ad, 32'h408bdffb, 32'h42487d48, 32'h42b45260, 32'h420fdb91, 32'h40f1ae61, 32'hbfc23775};
test_weights[34992:34999] = '{32'hc2acf6fb, 32'hc25cc7bb, 32'h4293331d, 32'h4278d7ea, 32'h42c0e498, 32'hc2beb89f, 32'hc1088649, 32'h42c3d7c3};
test_bias[4374:4374] = '{32'hc2b8dbc6};
test_output[4374:4374] = '{32'h46838b42};
test_input[35000:35007] = '{32'hc2add74b, 32'h42031954, 32'hc1fac53b, 32'hc1d93278, 32'hc25e42d3, 32'hc22d7a23, 32'hc22b119b, 32'h421307ec};
test_weights[35000:35007] = '{32'h42accfa4, 32'h42a8dd76, 32'hc2c5180c, 32'h421b797d, 32'hc12252d8, 32'hc1c8a390, 32'h425de6cd, 32'hc2925ca9};
test_bias[4375:4375] = '{32'h4095b35a};
test_output[4375:4375] = '{32'hc5bf1df3};
test_input[35008:35015] = '{32'hc2c0d0cd, 32'hc2a0ad65, 32'h42479a7b, 32'h4223afc2, 32'h425e1f20, 32'h42280c52, 32'hc22a1806, 32'h4212a7b6};
test_weights[35008:35015] = '{32'h42bb599c, 32'hc2c02430, 32'hc25ad80f, 32'hc22f99a8, 32'hc213a043, 32'hc1ae2f21, 32'h420b2ce1, 32'hc11a1486};
test_bias[4376:4376] = '{32'hc28a5b90};
test_output[4376:4376] = '{32'hc627457a};
test_input[35016:35023] = '{32'h42837ce7, 32'h425e330b, 32'hc29ceb24, 32'h42315534, 32'h41a6e128, 32'h420e4d10, 32'hc2aee477, 32'h42763aab};
test_weights[35016:35023] = '{32'hc1f6e70a, 32'h42425c36, 32'hc28d0caf, 32'h4283760a, 32'h414cc6c8, 32'hc2ae0002, 32'hc1ea96b0, 32'h42421867};
test_bias[4377:4377] = '{32'h41009b76};
test_output[4377:4377] = '{32'h463922c5};
test_input[35024:35031] = '{32'h4148a733, 32'h41f9f1b6, 32'hc2a543c5, 32'hc2646118, 32'h424429b4, 32'hbe2cbe76, 32'hc2c431bb, 32'hc2114650};
test_weights[35024:35031] = '{32'h42b5baaa, 32'h42c09025, 32'h429cda58, 32'hc1da1f65, 32'h413bed29, 32'hc2a3a22a, 32'hc2858ec1, 32'h3f0ee9e5};
test_bias[4378:4378] = '{32'h422b06ab};
test_output[4378:4378] = '{32'h45c79714};
test_input[35032:35039] = '{32'hc2a9ca5f, 32'h414b0a06, 32'hc2c7fb9b, 32'hc23d1e42, 32'hc05c3ab0, 32'h423c6876, 32'h4258d5bf, 32'h4127b7bd};
test_weights[35032:35039] = '{32'hc0fa099b, 32'h4288e917, 32'hc2c6cc8e, 32'h40fc23c0, 32'hc1a8f6f4, 32'hc18836a3, 32'hc092aa22, 32'h4124378b};
test_bias[4379:4379] = '{32'hc296ab20};
test_output[4379:4379] = '{32'h461ea45c};
test_input[35040:35047] = '{32'hc1dfb209, 32'h41deb89d, 32'hc242c3b5, 32'h42494be8, 32'hc07985f0, 32'hc1b67a09, 32'h42b6a1eb, 32'h427ed0ab};
test_weights[35040:35047] = '{32'h42265274, 32'h419b46ec, 32'h42934009, 32'hc284bc08, 32'h420aa578, 32'h4290242c, 32'hc193d291, 32'hc1d255eb};
test_bias[4380:4380] = '{32'h41aae320};
test_output[4380:4380] = '{32'hc645ebde};
test_input[35048:35055] = '{32'h4209b899, 32'h426b2847, 32'h4249079d, 32'hc11eb464, 32'h41cbebc6, 32'hc2aab1f6, 32'hc2627227, 32'hc2813171};
test_weights[35048:35055] = '{32'h42a375ea, 32'h42228aa3, 32'h4207590d, 32'h42b100c9, 32'hc12da178, 32'h4266254e, 32'h42a4bb58, 32'h42798b85};
test_bias[4381:4381] = '{32'h4279213b};
test_output[4381:4381] = '{32'hc5f380b7};
test_input[35056:35063] = '{32'hc2263c59, 32'hc21fca2a, 32'hc245fd35, 32'h41e27aa1, 32'hc29477cd, 32'hc29164e6, 32'h41897965, 32'h41c7ac9a};
test_weights[35056:35063] = '{32'hc1bc7f9e, 32'h41921ec6, 32'hc2387408, 32'h422d3dfa, 32'hc20c5851, 32'hc27ec3ea, 32'h41e54e11, 32'hc1314faa};
test_bias[4382:4382] = '{32'hc1916eef};
test_output[4382:4382] = '{32'h462edae7};
test_input[35064:35071] = '{32'hc2331651, 32'h42bd248d, 32'hc1554ec7, 32'h4256e83d, 32'h3fa50fa8, 32'hc273228c, 32'hc2b19319, 32'hc22e23f9};
test_weights[35064:35071] = '{32'hc2075014, 32'h42a331d8, 32'h4130175f, 32'hc11b2c51, 32'hc09f6f3c, 32'hc29647c7, 32'h3ee97821, 32'hc2a5b522};
test_bias[4383:4383] = '{32'h42a75680};
test_output[4383:4383] = '{32'h46830d4c};
test_input[35072:35079] = '{32'hc2463428, 32'hc11c2279, 32'h421a8e39, 32'hc27ef962, 32'hc285a979, 32'h421540d3, 32'h428f4db0, 32'hc254bda7};
test_weights[35072:35079] = '{32'h4199e074, 32'h42a866f3, 32'hc1308446, 32'h4200e02b, 32'hc1fb2b53, 32'hc25a3239, 32'hc26f6bea, 32'h41489bed};
test_bias[4384:4384] = '{32'h41ca826a};
test_output[4384:4384] = '{32'hc60e88e2};
test_input[35080:35087] = '{32'h42c179a6, 32'hc2718c38, 32'hc215ef7e, 32'hc2993991, 32'hc28ce2c2, 32'h426016c5, 32'hc1049b72, 32'hc21bb6f9};
test_weights[35080:35087] = '{32'h42801edf, 32'hc25dab75, 32'h4185e181, 32'hc18fdd44, 32'hc113a18d, 32'hc23550cf, 32'hc0ba07d3, 32'hc24ad5da};
test_bias[4385:4385] = '{32'h420bb52c};
test_output[4385:4385] = '{32'h4623768d};
test_input[35088:35095] = '{32'h42460049, 32'hc2b5e768, 32'hc2b965a4, 32'hc24c1a05, 32'hc1613cfa, 32'hc1bfcabd, 32'h409b4be7, 32'hc25b7445};
test_weights[35088:35095] = '{32'hc2788a97, 32'h429a2dd5, 32'h42afa46a, 32'hc2c765e9, 32'hc09cca84, 32'h428df9bc, 32'h424ca5f0, 32'h428a9fa7};
test_bias[4386:4386] = '{32'h415e56b4};
test_output[4386:4386] = '{32'hc68f1482};
test_input[35096:35103] = '{32'hc22796e2, 32'hc280036f, 32'hc279188e, 32'h421b18e7, 32'hc2c7d5ad, 32'h41eb9840, 32'hc1156b67, 32'h42a14164};
test_weights[35096:35103] = '{32'hc1ec2856, 32'h419d1fab, 32'h40aef5d0, 32'h415f9a3e, 32'hc0a83f57, 32'hc206d6e3, 32'h417f4fbe, 32'h42b89b39};
test_bias[4387:4387] = '{32'h422e425f};
test_output[4387:4387] = '{32'h45dc5355};
test_input[35104:35111] = '{32'h42c53740, 32'h428bfd85, 32'h3ffd783b, 32'h4107889c, 32'hc2add199, 32'hc2bf2f36, 32'hc2baa45f, 32'h40bd5481};
test_weights[35104:35111] = '{32'h42bddee6, 32'h4275b6f8, 32'h428106a7, 32'h42c415b5, 32'h429b5be6, 32'h426dc9a0, 32'hc2203b7c, 32'h427893ff};
test_bias[4388:4388] = '{32'h423a76d9};
test_output[4388:4388] = '{32'h45c61150};
test_input[35112:35119] = '{32'h4037876c, 32'hc0b1adbe, 32'hc2114df7, 32'h429a1714, 32'h42c08371, 32'hc2824584, 32'hc1b4dfb0, 32'hc2a97036};
test_weights[35112:35119] = '{32'hc269f189, 32'hbd29e08f, 32'h421d9e28, 32'h41f70b7a, 32'hc1acef86, 32'hc1e933ad, 32'h42883dda, 32'hc2369636};
test_bias[4389:4389] = '{32'hc28a6708};
test_output[4389:4389] = '{32'h45328093};
test_input[35120:35127] = '{32'h4284c3a0, 32'h429f4c6c, 32'h40ba31de, 32'h4183c672, 32'h42503911, 32'h41c752af, 32'h422ce414, 32'h4250e044};
test_weights[35120:35127] = '{32'h41fa576f, 32'hc2ab5cec, 32'hbf5207d3, 32'hc2126d05, 32'hc2af0232, 32'h41e97998, 32'h4216ee29, 32'hc27c2d29};
test_bias[4390:4390] = '{32'hc2325b51};
test_output[4390:4390] = '{32'hc62a22c2};
test_input[35128:35135] = '{32'hc2346066, 32'h4228025f, 32'h42b6b2ec, 32'h422c7612, 32'hc21c69c7, 32'h41ed95bf, 32'hc2c5068a, 32'h42776c94};
test_weights[35128:35135] = '{32'h42c5fc49, 32'h424fce48, 32'h3f9704d6, 32'hc24101f9, 32'h429dee3c, 32'h421f1274, 32'hc21eaae8, 32'hc28dde1e};
test_bias[4391:4391] = '{32'hc28d3d49};
test_output[4391:4391] = '{32'hc5d1bf43};
test_input[35136:35143] = '{32'hc2043f65, 32'h4295bab0, 32'hc2c7b12e, 32'h426eec03, 32'hc22ca907, 32'h3fe22bdb, 32'hc2b8b0b1, 32'h4105a0bf};
test_weights[35136:35143] = '{32'h42a50dae, 32'hc1d6eb2c, 32'h41b03924, 32'hc2532ac6, 32'h427dff91, 32'hc2b1caba, 32'hc1bf85f9, 32'hc22d023b};
test_bias[4392:4392] = '{32'h42545eed};
test_output[4392:4392] = '{32'hc62d3f2a};
test_input[35144:35151] = '{32'hc23ef48c, 32'h42409d48, 32'hc1dce0ba, 32'h42a14bb8, 32'h41d7d2b1, 32'h42231bfa, 32'h42b7a464, 32'h41aedecb};
test_weights[35144:35151] = '{32'h41049b91, 32'hc203b928, 32'h42960094, 32'h4238436c, 32'hc2835f5f, 32'hc2a2f2b1, 32'h425e8919, 32'hc2b50b3a};
test_bias[4393:4393] = '{32'hc0d2249e};
test_output[4393:4393] = '{32'hc510450b};
test_input[35152:35159] = '{32'h419e8a61, 32'h427e8d4d, 32'hc274c628, 32'hc27e56ec, 32'h42b22ed5, 32'h4252975a, 32'h3d9ecb1a, 32'h428f598f};
test_weights[35152:35159] = '{32'h4284313e, 32'h41665366, 32'hc233fe81, 32'hc183ce48, 32'h42b55013, 32'hc08f68cc, 32'h42437f6e, 32'hc25e80d5};
test_bias[4394:4394] = '{32'hbfda058f};
test_output[4394:4394] = '{32'h461a6c3f};
test_input[35160:35167] = '{32'h42665556, 32'hc24fb798, 32'hc2c6134f, 32'hc2c0a98b, 32'hc1db74bd, 32'h42a639fb, 32'hc1ca2580, 32'h427e5bf6};
test_weights[35160:35167] = '{32'hc2a3a164, 32'hc20033d1, 32'h42bcd4cc, 32'hc24ce8ef, 32'hc217f03a, 32'hc29c8706, 32'h422224b6, 32'h427bc760};
test_bias[4395:4395] = '{32'hc1ba5102};
test_output[4395:4395] = '{32'hc61bc9a6};
test_input[35168:35175] = '{32'hc180a35b, 32'h424e6fa8, 32'h42260c2e, 32'hc223b065, 32'h408a1b82, 32'hc2995284, 32'hc164648a, 32'h424b82a7};
test_weights[35168:35175] = '{32'hc05ad5cd, 32'hc1f22c6b, 32'h40d4b006, 32'h420db7c0, 32'hc13158f9, 32'hc2afbc27, 32'h4261fbc8, 32'hc259517b};
test_bias[4396:4396] = '{32'hc2b858e6};
test_output[4396:4396] = '{32'h43ac12a2};
test_input[35176:35183] = '{32'h42871211, 32'hc2c1a680, 32'hc281a4fe, 32'h4204f659, 32'h42c0c74b, 32'h423d139f, 32'h42c6ec36, 32'h3fec38f0};
test_weights[35176:35183] = '{32'h42939ece, 32'h424e76bf, 32'hc0ffe837, 32'h427b2edc, 32'hc20ed263, 32'hc23ec4df, 32'h41431b69, 32'hc217422a};
test_bias[4397:4397] = '{32'h42a5a676};
test_output[4397:4397] = '{32'hc4eaa910};
test_input[35184:35191] = '{32'hc25b6a29, 32'h423c064c, 32'hc0cb9a73, 32'h4283ea65, 32'hc2a613eb, 32'hc2a0bc36, 32'hc263a995, 32'hc2487c5e};
test_weights[35184:35191] = '{32'h41e8c141, 32'hc26ef558, 32'h423d51d3, 32'hc1cd7f26, 32'hc28c2679, 32'h4217c8a9, 32'h41db7661, 32'hc28b2cbb};
test_bias[4398:4398] = '{32'h425c0c8d};
test_output[4398:4398] = '{32'hc4ce14d8};
test_input[35192:35199] = '{32'hc27c843d, 32'h426fbf33, 32'hc2a73e03, 32'h42a4d3df, 32'h41571d54, 32'hc1cff388, 32'h429d8bea, 32'hc193ee23};
test_weights[35192:35199] = '{32'h4268c395, 32'h41885558, 32'hc292cf1f, 32'h42a59d5d, 32'hc2b97271, 32'hc2c2f864, 32'hc02c1226, 32'h42c64943};
test_bias[4399:4399] = '{32'h41c049da};
test_output[4399:4399] = '{32'h4615a370};
test_input[35200:35207] = '{32'h42abe75d, 32'hc2111c94, 32'hc0889c0d, 32'hc2019967, 32'hc24b9c07, 32'h4104da5d, 32'hc262c9e2, 32'h4226f6c1};
test_weights[35200:35207] = '{32'h4267f997, 32'h41e313cc, 32'h429b9e7c, 32'h427f57b2, 32'h42223077, 32'h42859a70, 32'h4283e05c, 32'hc28a61e1};
test_bias[4400:4400] = '{32'h42b62642};
test_output[4400:4400] = '{32'hc5cad292};
test_input[35208:35215] = '{32'hc24c41ad, 32'hc2c67959, 32'h4229e127, 32'hc25823f9, 32'h424ccd6b, 32'hc171018e, 32'h40e464cd, 32'hc26125d5};
test_weights[35208:35215] = '{32'hc2600e17, 32'h42be4981, 32'h419446a9, 32'hc28389f1, 32'h4232ea2f, 32'hc2394160, 32'h415cc1d3, 32'h41f951f7};
test_bias[4401:4401] = '{32'h4299c1c1};
test_output[4401:4401] = '{32'hc44fe19d};
test_input[35216:35223] = '{32'hc2959043, 32'h40fe848b, 32'hc10618e2, 32'h42a276eb, 32'hc2b47285, 32'h41ba5066, 32'hc2929612, 32'hc28899f4};
test_weights[35216:35223] = '{32'hc04bd872, 32'hc218f26a, 32'h428036ff, 32'h40ab15ce, 32'hc2323206, 32'hc186e0eb, 32'hc0607812, 32'h4015ecd1};
test_bias[4402:4402] = '{32'hc1c46468};
test_output[4402:4402] = '{32'h455ca4c5};
test_input[35224:35231] = '{32'hc2523429, 32'hc28e0d06, 32'hc185205a, 32'hc29d07d3, 32'hc265e267, 32'h420195e9, 32'h42a48487, 32'h42c20a7d};
test_weights[35224:35231] = '{32'hc209ab36, 32'h421eb275, 32'h42afb159, 32'hc126764a, 32'h41aca5ba, 32'h4267ecf2, 32'h424ac823, 32'h42406db6};
test_bias[4403:4403] = '{32'h4249394a};
test_output[4403:4403] = '{32'h45f5fdf5};
test_input[35232:35239] = '{32'hc2a1761b, 32'h42c56ab1, 32'h4215c2cc, 32'hc23cc22a, 32'h413a0876, 32'h42b8f812, 32'hc1fda617, 32'h40836ced};
test_weights[35232:35239] = '{32'h41562d0d, 32'hc2055701, 32'hc2c1443d, 32'h42a8b061, 32'hc1de8d7d, 32'hc2951708, 32'hc1188e8d, 32'h421e3ba2};
test_bias[4404:4404] = '{32'h422a569d};
test_output[4404:4404] = '{32'hc691ef35};
test_input[35240:35247] = '{32'h4206425e, 32'h41564076, 32'h41ef29e0, 32'h42821ab4, 32'h4125deff, 32'h42c5c2af, 32'h418e4558, 32'hc1d1e466};
test_weights[35240:35247] = '{32'h42bad08e, 32'hc1e6fc0d, 32'h42aa8081, 32'hc18d7440, 32'h415f5b11, 32'h400fe5d6, 32'h42812e54, 32'h427a060f};
test_bias[4405:4405] = '{32'hc2b487f0};
test_output[4405:4405] = '{32'h4575c745};
test_input[35248:35255] = '{32'hc139e908, 32'hc2a657ad, 32'h429b6ca3, 32'h4208109a, 32'h42708c0d, 32'hc1996387, 32'h4237b472, 32'hc0500243};
test_weights[35248:35255] = '{32'h4152a9e9, 32'hc20737bf, 32'hc2260fc0, 32'h423419ef, 32'hc2155f35, 32'hc14ee361, 32'h428f3731, 32'h42623006};
test_bias[4406:4406] = '{32'h42228fba};
test_output[4406:4406] = '{32'h4503fae1};
test_input[35256:35263] = '{32'hc2a473e6, 32'h4206790a, 32'hc22e67e1, 32'h40511cec, 32'h4267d2fa, 32'h41e47eb6, 32'h42270dc5, 32'h428fb75d};
test_weights[35256:35263] = '{32'h41fa6d81, 32'hc1c2d04a, 32'h425ea927, 32'hc25d4de5, 32'hc2c5f7b5, 32'h404ace2f, 32'h4236c765, 32'hc282c28a};
test_bias[4407:4407] = '{32'h42925d85};
test_output[4407:4407] = '{32'hc6606cdd};
test_input[35264:35271] = '{32'hc29e59a2, 32'hc29f024d, 32'hc2b3e2a8, 32'hc236955a, 32'hc25c0d5c, 32'hc2bbcb64, 32'h41147b8c, 32'hc2b4be64};
test_weights[35264:35271] = '{32'h40904581, 32'h429cce43, 32'hc29d98ef, 32'hc2644528, 32'hc0d1efbf, 32'h42c2e5d8, 32'h42c7537c, 32'hc204e7ad};
test_bias[4408:4408] = '{32'hc24f6f2b};
test_output[4408:4408] = '{32'hc4e27328};
test_input[35272:35279] = '{32'hc18419b1, 32'h429d7c5c, 32'h40eed76d, 32'h3f55d278, 32'h421dbbaa, 32'hc1c5aec2, 32'h3f27b988, 32'hc16e20a6};
test_weights[35272:35279] = '{32'h421b7561, 32'hc19ac07e, 32'h406552c2, 32'hc2587dcb, 32'hc14bd01f, 32'h428cb94a, 32'hc21a8114, 32'h42a23171};
test_bias[4409:4409] = '{32'hc2426b70};
test_output[4409:4409] = '{32'hc5b24a20};
test_input[35280:35287] = '{32'hc2460024, 32'h427b4a91, 32'h42321463, 32'hc0b45c51, 32'h420379e9, 32'h42c38ec2, 32'hc2328f33, 32'h429b2aa7};
test_weights[35280:35287] = '{32'h422a5de0, 32'h402b8f4e, 32'h41c61d53, 32'hc2c7674d, 32'hc2a3c307, 32'hc2c41d5e, 32'h423893bf, 32'h4258d0aa};
test_bias[4410:4410] = '{32'hc2b278cb};
test_output[4410:4410] = '{32'hc6240a16};
test_input[35288:35295] = '{32'h42548659, 32'hc24dd45e, 32'h42a736ae, 32'hc25eed86, 32'hc1924758, 32'hc252c27e, 32'hc19c1779, 32'h42810796};
test_weights[35288:35295] = '{32'hc190c8be, 32'hc14f5c54, 32'hc2330a74, 32'h4298dd1a, 32'hc2a6d2f4, 32'h4293641a, 32'hc2c288c9, 32'h4242fb56};
test_bias[4411:4411] = '{32'hc18c2f41};
test_output[4411:4411] = '{32'hc5afeaea};
test_input[35296:35303] = '{32'hc19ffa8e, 32'hc1e1af3b, 32'h4220a013, 32'h42aefe3d, 32'hc2bb25f9, 32'hc26b3c0b, 32'h423b8266, 32'hc2131cd4};
test_weights[35296:35303] = '{32'hc22e7ba5, 32'h41340781, 32'hc293b581, 32'hc28a7864, 32'hc296501e, 32'h40ea8082, 32'hc2525edb, 32'hc22709b4};
test_bias[4412:4412] = '{32'h42369a6f};
test_output[4412:4412] = '{32'hc52bedaf};
test_input[35304:35311] = '{32'h4298c808, 32'h429e5ad7, 32'h429de369, 32'hc2449e3d, 32'hc0a064b9, 32'hc1e6dfd7, 32'h41e98af6, 32'h42b361f5};
test_weights[35304:35311] = '{32'h40dd7962, 32'h422e27ee, 32'h42ba13df, 32'hc28d1c99, 32'hc1abcb88, 32'hc0da6687, 32'h4297b6f1, 32'h4274a373};
test_bias[4413:4413] = '{32'hc28fa877};
test_output[4413:4413] = '{32'h46b1838b};
test_input[35312:35319] = '{32'hc1a74c58, 32'hc230645f, 32'h42beeb34, 32'hc2335ba5, 32'hc00db39d, 32'h4299e5a6, 32'h4279cd82, 32'h429c27d3};
test_weights[35312:35319] = '{32'h40a529fa, 32'hc2839e86, 32'hc1280eb0, 32'hc281619f, 32'h408111af, 32'h429b91d2, 32'h42a4f3dd, 32'h41b67730};
test_bias[4414:4414] = '{32'h42281857};
test_output[4414:4414] = '{32'h4689d468};
test_input[35320:35327] = '{32'hc1e5d376, 32'hc2c5af3a, 32'h429a80fb, 32'h42b17a46, 32'h414c087f, 32'hc270fd69, 32'hc2204ce5, 32'hc208d2c1};
test_weights[35320:35327] = '{32'hc25d571b, 32'hc1f05b84, 32'hc21012aa, 32'hc11e0eed, 32'h40a6ab87, 32'h424d8ccf, 32'h41579597, 32'h42c1113e};
test_bias[4415:4415] = '{32'hc20fe45e};
test_output[4415:4415] = '{32'hc5bbb9ec};
test_input[35328:35335] = '{32'hc21047e4, 32'hc223dea3, 32'h4226770f, 32'hc2b8b1cc, 32'h4228fcd9, 32'h410877b4, 32'hc2422971, 32'hc190a9c3};
test_weights[35328:35335] = '{32'h4294e740, 32'h42276e48, 32'hc287320b, 32'h41f7f76f, 32'h424817e2, 32'hc25a984b, 32'h42b2ab7e, 32'h42878746};
test_bias[4416:4416] = '{32'h419ccaa8};
test_output[4416:4416] = '{32'hc65a4afd};
test_input[35336:35343] = '{32'hc20c00a7, 32'h406ef5f9, 32'h41f39e2b, 32'hc1ec3776, 32'h42793027, 32'hc2afb1b8, 32'h4194b5cd, 32'hc270d6d0};
test_weights[35336:35343] = '{32'h424cc73b, 32'hc00760bd, 32'hc23550c0, 32'h429fba3e, 32'hc2a3fea1, 32'hc285ab25, 32'h42865561, 32'h415cc472};
test_bias[4417:4417] = '{32'hc156689d};
test_output[4417:4417] = '{32'hc58896ec};
test_input[35344:35351] = '{32'hc2769898, 32'h42ba8981, 32'h428fb572, 32'hc2566e20, 32'hc26df7eb, 32'hc20688de, 32'hc28497cd, 32'hc08a81da};
test_weights[35344:35351] = '{32'hc26255a1, 32'hc27e5534, 32'h42028a5d, 32'h4287c80f, 32'h42c5c851, 32'hc286e3bc, 32'hc140ae7b, 32'h42b0cb53};
test_bias[4418:4418] = '{32'hc252e0d4};
test_output[4418:4418] = '{32'hc5da6206};
test_input[35352:35359] = '{32'hc0a35655, 32'h42c58dad, 32'hc1eee2f5, 32'hc0dce62e, 32'h42292997, 32'hc2455628, 32'h425947b8, 32'h414089eb};
test_weights[35352:35359] = '{32'h424280a7, 32'hc11140c9, 32'hc0f0c60d, 32'h41a68f9a, 32'hc11094ed, 32'hc2686db0, 32'h4271cd64, 32'hc1374ef6};
test_bias[4419:4419] = '{32'h42565d66};
test_output[4419:4419] = '{32'h45905f8a};
test_input[35360:35367] = '{32'h40a8ac61, 32'hc2bd5036, 32'h42249a73, 32'hc2961350, 32'h42a293f4, 32'h42a66c13, 32'h428cb832, 32'hc2add681};
test_weights[35360:35367] = '{32'hc23130f5, 32'hc26665ba, 32'h40d93b40, 32'h41b14e46, 32'h425cb993, 32'hc1309e9c, 32'h429c36f2, 32'h4280ba80};
test_bias[4420:4420] = '{32'h417cf346};
test_output[4420:4420] = '{32'h45e4b7be};
test_input[35368:35375] = '{32'h42290037, 32'h41da9b35, 32'h42b9c61b, 32'hc2b37175, 32'h41b8b7ab, 32'h41078aff, 32'h420661c7, 32'h423eab0c};
test_weights[35368:35375] = '{32'h42ad7090, 32'h421a8e35, 32'h41b279b2, 32'hc2a66b78, 32'hc26d69d3, 32'h41f703f3, 32'hc17db483, 32'h420578f0};
test_bias[4421:4421] = '{32'h42bcad96};
test_output[4421:4421] = '{32'h465f743c};
test_input[35376:35383] = '{32'h41186d67, 32'hc2bc8458, 32'h429bbf94, 32'hbfed48b1, 32'h410b4df1, 32'hc272533a, 32'hc213b223, 32'hc2a23391};
test_weights[35376:35383] = '{32'hc0316eb0, 32'h41a8b410, 32'h42a0f141, 32'h42301678, 32'hc22c970a, 32'hc2bc653a, 32'h419ce769, 32'h41b2d02b};
test_bias[4422:4422] = '{32'h411549a7};
test_output[4422:4422] = '{32'h45d9f206};
test_input[35384:35391] = '{32'hc1e425c2, 32'hc2a1affc, 32'h41a4309a, 32'h414e6286, 32'hc2a16dbb, 32'hc2a22c5a, 32'hc274a0cf, 32'h424c7c90};
test_weights[35384:35391] = '{32'hc226e1c1, 32'hc224b30d, 32'h4233f118, 32'h4148e643, 32'hc21f803b, 32'h42c6ea14, 32'hc1f1f9d5, 32'h41ea851b};
test_bias[4423:4423] = '{32'hc0a87982};
test_output[4423:4423] = '{32'h45802666};
test_input[35392:35399] = '{32'hc2218fe7, 32'h41e50051, 32'hc2163c37, 32'hc2325da8, 32'hc2248252, 32'h42c0cc62, 32'hc25cab7b, 32'h4013ee6a};
test_weights[35392:35399] = '{32'hc1c12b50, 32'hc25127dc, 32'hc29a0eba, 32'hc242c078, 32'h42aa1d40, 32'h402d26bd, 32'h429c54e8, 32'h42461fb5};
test_bias[4424:4424] = '{32'h423be98b};
test_output[4424:4424] = '{32'hc531d6ec};
test_input[35400:35407] = '{32'hc1adac15, 32'h429853da, 32'hc27fc4ae, 32'h428b1a84, 32'h428bb98a, 32'hc289802f, 32'hc1b48f32, 32'hc29de9af};
test_weights[35400:35407] = '{32'hc0fbc222, 32'hc2882c88, 32'hc221f184, 32'h4263831a, 32'hc26613a5, 32'h420327c8, 32'h429798f0, 32'h416e1a06};
test_bias[4425:4425] = '{32'h40500b01};
test_output[4425:4425] = '{32'hc5ee4b59};
test_input[35408:35415] = '{32'h42c68176, 32'h42c55a02, 32'hbf6a076c, 32'hc202c1cb, 32'h4261460b, 32'hc03ba37f, 32'h41748bfc, 32'h42a1d687};
test_weights[35408:35415] = '{32'h423be0fb, 32'h42a442b7, 32'h4292935b, 32'hc1cbe0dd, 32'hc296a7e2, 32'hc17ee7e0, 32'h42402219, 32'h428a2efc};
test_bias[4426:4426] = '{32'hc24166ac};
test_output[4426:4426] = '{32'h4673f4eb};
test_input[35416:35423] = '{32'hc2071ce5, 32'hc2c40002, 32'h41b54ebb, 32'h42af4fd7, 32'h4260b178, 32'h421742b1, 32'hc2309ac4, 32'h42a010a9};
test_weights[35416:35423] = '{32'h41c36e9b, 32'hc2a259ee, 32'hc2c10fd5, 32'hc2911e88, 32'h420af008, 32'hc2835805, 32'h42b4e4a0, 32'hc1facd3d};
test_bias[4427:4427] = '{32'hc214261f};
test_output[4427:4427] = '{32'hc604a663};
test_input[35424:35431] = '{32'h40e608af, 32'hc295c9b9, 32'h423719dd, 32'hc268429a, 32'h424399dd, 32'h427c63a3, 32'hc0c930de, 32'h41c4de26};
test_weights[35424:35431] = '{32'hc29af20e, 32'hc2825644, 32'h428debaf, 32'h429503fc, 32'hc2af457a, 32'h422c8ced, 32'h427257ca, 32'hc277abde};
test_bias[4428:4428] = '{32'h42bcd0d5};
test_output[4428:4428] = '{32'hc3000305};
test_input[35432:35439] = '{32'hc28435bd, 32'h4294f369, 32'h424dd24a, 32'hc291614e, 32'hc2841386, 32'h42816295, 32'h42ad131b, 32'hc2b2df8b};
test_weights[35432:35439] = '{32'hc23d9b13, 32'hc2245904, 32'hc227720b, 32'hc1bc9118, 32'hc24400f2, 32'h418a75d8, 32'h41dadd92, 32'hc1e7476e};
test_bias[4429:4429] = '{32'hc296f754};
test_output[4429:4429] = '{32'h460a8865};
test_input[35440:35447] = '{32'h420ebe73, 32'h42a187f6, 32'h42b4cc38, 32'hc1e714c9, 32'h410173cc, 32'h428ff264, 32'hc2998cd7, 32'h421b292a};
test_weights[35440:35447] = '{32'h42bad5dc, 32'h4291071f, 32'hc104e580, 32'h40c8cfd2, 32'hc2733d20, 32'h426a8030, 32'hbf11c246, 32'h426f49bf};
test_bias[4430:4430] = '{32'hc1af4d77};
test_output[4430:4430] = '{32'h465fdfe5};
test_input[35448:35455] = '{32'h3f6fb36a, 32'hc25acd1b, 32'h427e70fb, 32'hc2169cdd, 32'hc26f6054, 32'h41e416eb, 32'hc29cd704, 32'hc2461d14};
test_weights[35448:35455] = '{32'h41aaa083, 32'h4205723b, 32'h423347c4, 32'h405a3fc8, 32'hc1e15d72, 32'h42bd7018, 32'hc21a8f73, 32'h41a0adab};
test_bias[4431:4431] = '{32'h425e6119};
test_output[4431:4431] = '{32'h45e7189d};
test_input[35456:35463] = '{32'h42c11398, 32'hc2a3cfe7, 32'hc2abb1c0, 32'h3eb0010d, 32'hc26f177e, 32'h4203fd40, 32'hc172c6f7, 32'h42c23b7f};
test_weights[35456:35463] = '{32'h41932f2a, 32'hc297fb53, 32'h4195f0b0, 32'h42b93350, 32'h42a0c9d8, 32'h425d39c4, 32'hc2339261, 32'hc2046447};
test_bias[4432:4432] = '{32'hc1942fec};
test_output[4432:4432] = '{32'h445ebca6};
test_input[35464:35471] = '{32'hc21dd47a, 32'h41094fa5, 32'hc2378840, 32'h42b02b49, 32'h42686dad, 32'h427c764a, 32'hc20bc0e6, 32'h40f4c379};
test_weights[35464:35471] = '{32'hc1d3b94d, 32'hc233d9b9, 32'h42bd4a22, 32'h41df458f, 32'hc21e1b9f, 32'hc2c6959c, 32'h41a9a991, 32'h41edf8c5};
test_bias[4433:4433] = '{32'hc146d8e8};
test_output[4433:4433] = '{32'hc6212d93};
test_input[35472:35479] = '{32'h428e13c0, 32'h41f59ada, 32'hc1164714, 32'h429380b4, 32'hc1e19487, 32'hbfe98a55, 32'hc2b8e8cd, 32'h421233ae};
test_weights[35472:35479] = '{32'h429ab33a, 32'hbf9e529b, 32'h42536ad9, 32'hbe1ca169, 32'h3fe468b0, 32'h425ecf38, 32'hc26ffd05, 32'h42905f73};
test_bias[4434:4434] = '{32'hc275102e};
test_output[4434:4434] = '{32'h4649e59d};
test_input[35480:35487] = '{32'h4029a418, 32'hc1bf850d, 32'h4228bfa9, 32'h4287a82e, 32'hc2898b5d, 32'hc2b0af39, 32'hc280db93, 32'hc244546c};
test_weights[35480:35487] = '{32'hc0544206, 32'h412251bc, 32'hc2336bd2, 32'h418853a0, 32'h4057d988, 32'hc2c52e29, 32'h41d75adf, 32'h4283582b};
test_bias[4435:4435] = '{32'h420315d3};
test_output[4435:4435] = '{32'h45204a3c};
test_input[35488:35495] = '{32'h4253b6a0, 32'h42bdc5f7, 32'h423963fa, 32'h41b41a42, 32'h425c31e1, 32'hc22a2291, 32'hc28c6751, 32'hc2b083ec};
test_weights[35488:35495] = '{32'h408e2471, 32'h424a4ef5, 32'h4165355a, 32'hc208d697, 32'hc266a528, 32'h424ee8de, 32'hc1dacc46, 32'hc2359417};
test_bias[4436:4436] = '{32'h42739318};
test_output[4436:4436] = '{32'h45ad27cc};
test_input[35496:35503] = '{32'h420b53ea, 32'hc2a3b038, 32'hc1a34fa0, 32'hc27f8417, 32'h40863576, 32'hc22c1302, 32'hc281bd72, 32'hc21b8b0d};
test_weights[35496:35503] = '{32'h42845c42, 32'h425d78df, 32'hc26ec9be, 32'h42c08991, 32'hc250d44d, 32'h41982215, 32'hc246ad34, 32'h42568b00};
test_bias[4437:4437] = '{32'h42952ff7};
test_output[4437:4437] = '{32'hc5da3aa3};
test_input[35504:35511] = '{32'h42c72089, 32'h4293aafc, 32'hc21acab5, 32'hc22b0341, 32'hc240aeb0, 32'h4193b2a2, 32'h3f9b8c4e, 32'hc0d92d6d};
test_weights[35504:35511] = '{32'hc267c453, 32'hc189873d, 32'h41251c76, 32'h42998ed0, 32'h4232a3b7, 32'hc1073e5f, 32'h42ae72c0, 32'h4240f5ca};
test_bias[4438:4438] = '{32'h42acab54};
test_output[4438:4438] = '{32'hc64da9db};
test_input[35512:35519] = '{32'h42c0bec6, 32'hc24fb8ff, 32'h423b4348, 32'hc08e06a8, 32'h41b2b5f8, 32'hc2b13052, 32'h42a0e0b1, 32'hc29b5735};
test_weights[35512:35519] = '{32'h4218405f, 32'hc22a109a, 32'h4281caba, 32'h42a9fb17, 32'h42bacaee, 32'h422438b1, 32'h42aeedcb, 32'hc10f349e};
test_bias[4439:4439] = '{32'h428de5fa};
test_output[4439:4439] = '{32'h46670f39};
test_input[35520:35527] = '{32'hc0a037bf, 32'hc29e5a71, 32'h42b29116, 32'hc27e3026, 32'h4083de26, 32'hc19c2f40, 32'h4218cbca, 32'hc2523b86};
test_weights[35520:35527] = '{32'hc2c51ed4, 32'hc24f377a, 32'h420251e2, 32'h42be2af0, 32'hc1890228, 32'h416e299c, 32'h4249078f, 32'h3fd69271};
test_bias[4440:4440] = '{32'hc2353e01};
test_output[4440:4440] = '{32'h45346e4a};
test_input[35528:35535] = '{32'hc143d5a7, 32'h4247d985, 32'hc1d632a8, 32'h42a405c8, 32'h42c67278, 32'h4219ed96, 32'hc295c2b8, 32'h42c38715};
test_weights[35528:35535] = '{32'hc269bb88, 32'hc225e073, 32'h428b4d27, 32'h42903989, 32'h40477bf4, 32'h42584585, 32'h4221cd6b, 32'hc27285f0};
test_bias[4441:4441] = '{32'h4271147a};
test_output[4441:4441] = '{32'hc56e5d10};
test_input[35536:35543] = '{32'hbf8e71b0, 32'hc2161135, 32'hc2c5c973, 32'hc18a2130, 32'h42b89633, 32'h42015033, 32'hc1d45f71, 32'hc26065d4};
test_weights[35536:35543] = '{32'hbf2c3b4b, 32'h42418863, 32'hc2acccc9, 32'h42668ad9, 32'h427755fd, 32'h40048e89, 32'hc19cdb0f, 32'hc2bfccb4};
test_bias[4442:4442] = '{32'hc1e14623};
test_output[4442:4442] = '{32'h4687c9cc};
test_input[35544:35551] = '{32'hbe9c9b0f, 32'hc2801a72, 32'hc1e1098f, 32'hc297055c, 32'h426c3898, 32'h42afa2e1, 32'h42c79e1d, 32'h42997e83};
test_weights[35544:35551] = '{32'h41911c50, 32'h42183451, 32'h428078f0, 32'hc2b58dc1, 32'h42265916, 32'hc1678abb, 32'hc1aa9dc4, 32'h419732aa};
test_bias[4443:4443] = '{32'hc28217d7};
test_output[4443:4443] = '{32'h453e6c97};
test_input[35552:35559] = '{32'h4240624c, 32'h428bc0c1, 32'h429fa067, 32'h421f7f88, 32'hc287d185, 32'hc21ba254, 32'hc2b315f8, 32'h42325f08};
test_weights[35552:35559] = '{32'h4220cec0, 32'hc2ad8d40, 32'hc299bdb5, 32'hc285820f, 32'h406df4b9, 32'hc1f5da10, 32'hc1139bf6, 32'hc25dde42};
test_bias[4444:4444] = '{32'hc2056ec2};
test_output[4444:4444] = '{32'hc6558261};
test_input[35560:35567] = '{32'hc2545b4d, 32'hc2c2a9c1, 32'h428cfb6a, 32'hc120a652, 32'h4287bfc8, 32'h41658b63, 32'hc21fac6e, 32'hc247b8cf};
test_weights[35560:35567] = '{32'h424ffbd2, 32'hc2bd5a76, 32'hc2ad6fcb, 32'hc2890dfe, 32'h422840c8, 32'h42a3bf22, 32'hc11573e8, 32'hc21d4003};
test_bias[4445:4445] = '{32'h4068113b};
test_output[4445:4445] = '{32'h45e7367a};
test_input[35568:35575] = '{32'hc2333107, 32'hc15f47a8, 32'h42a350c6, 32'h42aabd62, 32'h3fa3208c, 32'hc275874c, 32'h4260e29f, 32'hc289ce08};
test_weights[35568:35575] = '{32'h4099493a, 32'hc209d419, 32'hc2bf699a, 32'hc21392ee, 32'hc1ab8c94, 32'hc27b4d3d, 32'hc2ba0eab, 32'h42ba04a8};
test_bias[4446:4446] = '{32'h42bb6483};
test_output[4446:4446] = '{32'hc68fdd04};
test_input[35576:35583] = '{32'h42508108, 32'hc29cb975, 32'hc2016304, 32'h416b8d2b, 32'hc2a26d2e, 32'hc171b6bf, 32'hc2093572, 32'h42a035d8};
test_weights[35576:35583] = '{32'hc12672cf, 32'hc0db271f, 32'hc26c5502, 32'hc24483e1, 32'h42ae9649, 32'h4241987b, 32'hc1ab30f6, 32'h423aa300};
test_bias[4447:4447] = '{32'h401a183c};
test_output[4447:4447] = '{32'hc5074370};
test_input[35584:35591] = '{32'h41e52ef3, 32'h4230cc04, 32'hc1ff133f, 32'h42133ed3, 32'h4215a3a8, 32'h42b67520, 32'hc2ab635d, 32'hc2c5799e};
test_weights[35584:35591] = '{32'h4241077e, 32'h41b4eb13, 32'h428571ce, 32'h421df57e, 32'h420a5856, 32'h422dd290, 32'h427e07a8, 32'hc024ee2b};
test_bias[4448:4448] = '{32'hbfcd61b5};
test_output[4448:4448] = '{32'h44de2663};
test_input[35592:35599] = '{32'hbf3c2721, 32'hc1fa07eb, 32'h42943276, 32'h422848eb, 32'hc0fa3df5, 32'hc12ad198, 32'h422a3b7e, 32'h42c697be};
test_weights[35592:35599] = '{32'h41808805, 32'hc2992009, 32'hbfa7a2bf, 32'h4200d258, 32'h41ae750b, 32'h428eef6a, 32'hc2bd32e1, 32'hc0b6a856};
test_bias[4449:4449] = '{32'hc2c58cf0};
test_output[4449:4449] = '{32'hc4f843e5};
test_input[35600:35607] = '{32'hc15d07db, 32'h4299323f, 32'hc0927a78, 32'h4238f0ca, 32'hc0ba3d7b, 32'hc28dad59, 32'hc2284619, 32'hc2747269};
test_weights[35600:35607] = '{32'h40da0137, 32'hc2679846, 32'h429f9871, 32'h42a8e71d, 32'h41bd7689, 32'hc1f37876, 32'hc1a9bbcf, 32'hbf16b1c4};
test_bias[4450:4450] = '{32'hbf32608e};
test_output[4450:4450] = '{32'h44f4861a};
test_input[35608:35615] = '{32'hc2c1bd31, 32'h41726dc5, 32'hc23db1e6, 32'hc28d0df9, 32'hc27d5393, 32'hbf72aa3b, 32'hc2011d4b, 32'hc0dd37b2};
test_weights[35608:35615] = '{32'hc1ad0bca, 32'h4190832a, 32'h42222b1c, 32'h420bc73b, 32'h40f96804, 32'h42aefcfb, 32'h42a3d924, 32'hc0b03fef};
test_bias[4451:4451] = '{32'hc287b0f7};
test_output[4451:4451] = '{32'hc5a4a6c3};
test_input[35616:35623] = '{32'h4131ce7f, 32'h41be22c6, 32'h4278a1bd, 32'hc2b94c91, 32'hc1e8ef2b, 32'h4113e0d8, 32'h427149f2, 32'h40f1c80c};
test_weights[35616:35623] = '{32'hc27cf6f5, 32'hc02cf52b, 32'hc2bf4fc0, 32'h42701716, 32'hc294119d, 32'hbe857420, 32'h4236d25f, 32'hc2abb6ec};
test_bias[4452:4452] = '{32'h425988b0};
test_output[4452:4452] = '{32'hc5f8af1b};
test_input[35624:35631] = '{32'hc19798b1, 32'hc20b93c6, 32'h427791af, 32'hc26871e6, 32'h418affec, 32'hc1193e4b, 32'h427d881d, 32'hc2396c63};
test_weights[35624:35631] = '{32'hc27195c4, 32'h41327624, 32'hc2076928, 32'h42a82994, 32'h42173884, 32'h42bd8487, 32'hc29ad2e3, 32'h42167783};
test_bias[4453:4453] = '{32'hc232c286};
test_output[4453:4453] = '{32'hc64dcf00};
test_input[35632:35639] = '{32'hc263f9f9, 32'h4268ea09, 32'hc22f5acb, 32'hc27d4c71, 32'h4106303e, 32'hc092df80, 32'hc2baa521, 32'hc11f7ff5};
test_weights[35632:35639] = '{32'hc29368be, 32'hc284dadd, 32'hc23cf836, 32'hc22b6832, 32'hc1290311, 32'hc2ae0e62, 32'h42389ee9, 32'hc243201b};
test_bias[4454:4454] = '{32'hc22b671c};
test_output[4454:4454] = '{32'h44c38abb};
test_input[35640:35647] = '{32'hc2a9ae7d, 32'hc2a32fb8, 32'hc2b13815, 32'hc2b37533, 32'h41120f32, 32'h4243e53f, 32'h42735f5e, 32'hc2b2d004};
test_weights[35640:35647] = '{32'h429a4ae5, 32'h422f3cab, 32'h4294136f, 32'h412e4e81, 32'hc2c4788f, 32'hc1b4747a, 32'h4286332b, 32'hc0a2dde2};
test_bias[4455:4455] = '{32'hc22ac3a4};
test_output[4455:4455] = '{32'hc66cf0e0};
test_input[35648:35655] = '{32'h42bc2a48, 32'h41e289f1, 32'h423175eb, 32'h41d45146, 32'h4269040a, 32'hc2c089bf, 32'hc294569c, 32'h42413279};
test_weights[35648:35655] = '{32'h421b79c4, 32'hc28e6fa3, 32'h41fdbd04, 32'h4185b57d, 32'h4203d0f0, 32'hc266b33f, 32'hc1c4e97d, 32'hc0fbe55c};
test_bias[4456:4456] = '{32'hc2320fe3};
test_output[4456:4456] = '{32'h46412f3a};
test_input[35656:35663] = '{32'hc26c6606, 32'hbef5fd92, 32'h42c7c22a, 32'hc25aed75, 32'hc2be2d43, 32'hc2b3f18c, 32'h42c43aa6, 32'h42418871};
test_weights[35656:35663] = '{32'hc26e0de6, 32'h423dd3fe, 32'hc29e14b4, 32'h42a993a9, 32'hc05b232c, 32'hc2c2c65c, 32'h42b8ba3f, 32'hc29617c1};
test_bias[4457:4457] = '{32'hc2b286e3};
test_output[4457:4457] = '{32'h45a867dd};
test_input[35664:35671] = '{32'hc1d00bdc, 32'h428e7373, 32'h42555869, 32'hc14d27cf, 32'h4291599e, 32'h4276686c, 32'h42b41e54, 32'h42a28f88};
test_weights[35664:35671] = '{32'h428e94cd, 32'hc2a51188, 32'hc208123d, 32'h4271de85, 32'hc188891a, 32'hc0e6e97f, 32'h42231b78, 32'hc1035d29};
test_bias[4458:4458] = '{32'h4213bcbd};
test_output[4458:4458] = '{32'hc60c1499};
test_input[35672:35679] = '{32'h41ef98b9, 32'hc2b3cc19, 32'hc24a60a5, 32'hc2678e49, 32'h426289f2, 32'hc29c682a, 32'hc25250b5, 32'h419bb406};
test_weights[35672:35679] = '{32'h418c5de5, 32'hc2675537, 32'hc1948803, 32'hc093c62b, 32'h424a5502, 32'hc22819ff, 32'h4193abb9, 32'h42173977};
test_bias[4459:4459] = '{32'h429ba3b1};
test_output[4459:4459] = '{32'h4649f6b6};
test_input[35680:35687] = '{32'h42ba502e, 32'h418f1030, 32'h41eb70f6, 32'hc28a889c, 32'h42643c2f, 32'hc280310f, 32'hc16cf11e, 32'hc1aa90e7};
test_weights[35680:35687] = '{32'hc2842a33, 32'hc262e5a6, 32'hc1b9e6a1, 32'h41a35ecb, 32'hc2222c8a, 32'hc2863683, 32'h42001dd9, 32'hc2693665};
test_bias[4460:4460] = '{32'h41ff1db2};
test_output[4460:4460] = '{32'hc5ca8251};
test_input[35688:35695] = '{32'hc2afcc44, 32'h42a7ad72, 32'h4265b913, 32'h42bd2d4c, 32'h4283e73d, 32'h42801ee1, 32'h40f22118, 32'h40a0a5c8};
test_weights[35688:35695] = '{32'h42ad8fde, 32'hc204210a, 32'hbf3805b3, 32'h4227180b, 32'hc2957672, 32'hc12e5512, 32'h42b8bd8b, 32'hc1ef11b4};
test_bias[4461:4461] = '{32'hc28525df};
test_output[4461:4461] = '{32'hc635be9b};
test_input[35696:35703] = '{32'hc1ef92cb, 32'hc2682056, 32'hc1e76ea4, 32'hc1936316, 32'h42793032, 32'h414658ae, 32'hc21b17f8, 32'hc22f4019};
test_weights[35696:35703] = '{32'h412c3f9e, 32'hc19d5579, 32'h41e177cc, 32'h41f33425, 32'h418e556f, 32'h42b4fabd, 32'hc12c4024, 32'hc2a7815e};
test_bias[4462:4462] = '{32'hc2b49200};
test_output[4462:4462] = '{32'h45b13197};
test_input[35704:35711] = '{32'h422303a2, 32'h42bb55a5, 32'h42a7d546, 32'h426e4b4b, 32'hc23a945e, 32'hc24fb623, 32'h427a272c, 32'hc106637b};
test_weights[35704:35711] = '{32'h42051fe3, 32'hc1c05517, 32'hc2790104, 32'h427c297c, 32'h41ca335a, 32'h4194c37f, 32'h42c198a5, 32'hc0442770};
test_bias[4463:4463] = '{32'h41409da3};
test_output[4463:4463] = '{32'h44c5dbc8};
test_input[35712:35719] = '{32'hc293d609, 32'h42b5f2cc, 32'h41f47b74, 32'hc2a0211e, 32'hc24c77f5, 32'hc29cfd58, 32'h420356e6, 32'hc191d234};
test_weights[35712:35719] = '{32'hc1893adc, 32'h4299daeb, 32'h42a1daa9, 32'hc2a61bcd, 32'h425f5b98, 32'hc235cd18, 32'h4226fcf2, 32'hc2b7384f};
test_bias[4464:4464] = '{32'h3efcac3b};
test_output[4464:4464] = '{32'h46a52f38};
test_input[35720:35727] = '{32'hc1f6a194, 32'hc2a58d06, 32'h4204ae31, 32'h41c9648b, 32'h4188feaa, 32'h41e40913, 32'hc18d74c7, 32'h42a94068};
test_weights[35720:35727] = '{32'h42b69d69, 32'h40d98a6a, 32'h4291f8f0, 32'h4290fa66, 32'h429da179, 32'h4257237c, 32'h427787c5, 32'h42be3229};
test_bias[4465:4465] = '{32'hc2604867};
test_output[4465:4465] = '{32'h4626619d};
test_input[35728:35735] = '{32'h425b164c, 32'h42b36d00, 32'h42c0d189, 32'hc268daab, 32'hc2bb46fb, 32'hc0b8a2c8, 32'h40c874db, 32'h4192ade1};
test_weights[35728:35735] = '{32'hc20501be, 32'h429b4035, 32'hc2ab8b58, 32'hc29f9204, 32'hc29ee643, 32'h42b433d2, 32'h423ec44d, 32'h42c6abf9};
test_bias[4466:4466] = '{32'h40e2d100};
test_output[4466:4466] = '{32'h462513c4};
test_input[35736:35743] = '{32'h4117672b, 32'h41c47202, 32'h421860a5, 32'h426ce4b7, 32'hc28616e1, 32'hc1e15037, 32'h421f4cfe, 32'h42c26a81};
test_weights[35736:35743] = '{32'h42b2140c, 32'h420f5670, 32'h4237b5f0, 32'h42509537, 32'h42a567f0, 32'hc2bbbb4d, 32'h423973aa, 32'hc2c5232f};
test_bias[4467:4467] = '{32'hc2c3f1d0};
test_output[4467:4467] = '{32'hc582706e};
test_input[35744:35751] = '{32'hc2580235, 32'hc27a3e73, 32'hc1e5997d, 32'hc2399bb9, 32'h408f4f90, 32'hc2169795, 32'h41e82b2b, 32'h42c16e67};
test_weights[35744:35751] = '{32'h4213e391, 32'h41291866, 32'hc243dd97, 32'hc28a4131, 32'h411dd155, 32'h422727c4, 32'h42278b15, 32'hc1d6b013};
test_bias[4468:4468] = '{32'hc1c33527};
test_output[4468:4468] = '{32'hc474899a};
test_input[35752:35759] = '{32'hc1cbc23a, 32'hc289f307, 32'h41ff15e0, 32'h425ff43d, 32'hc1f896ab, 32'hc1a354b4, 32'h42bbad6d, 32'h42bf0948};
test_weights[35752:35759] = '{32'hc22dbf06, 32'h40aadbf5, 32'hc2b65854, 32'h418ca889, 32'hc0e7a69b, 32'h427f3c6f, 32'hc2444769, 32'hc201ce92};
test_bias[4469:4469] = '{32'h3fbe8337};
test_output[4469:4469] = '{32'hc61bb556};
test_input[35760:35767] = '{32'h42b9a473, 32'hc1994cff, 32'hc1df76a4, 32'hc2a8c621, 32'hc27754fd, 32'hc201c9d3, 32'h41ab6719, 32'hc18d4111};
test_weights[35760:35767] = '{32'h429c12e3, 32'h41ba5134, 32'h413d78d2, 32'h42914f62, 32'hc264ea5a, 32'h42a31513, 32'h41da7b5e, 32'hc1caa2d7};
test_bias[4470:4470] = '{32'hc2bb6fe4};
test_output[4470:4470] = '{32'h45076c61};
test_input[35768:35775] = '{32'h42a47567, 32'h41a053d6, 32'hc2c500b4, 32'h42140b09, 32'h42b651ae, 32'hc2855d5b, 32'h4278a36b, 32'h419e06bf};
test_weights[35768:35775] = '{32'h421fa5b3, 32'h42975ed3, 32'h4291e587, 32'hc25c62cc, 32'hc1c157aa, 32'hc29c4af0, 32'hc2c25994, 32'hc190bc5b};
test_bias[4471:4471] = '{32'hc20f18b6};
test_output[4471:4471] = '{32'hc5f55cc5};
test_input[35776:35783] = '{32'hc2b92e5f, 32'h415f4299, 32'h428260f7, 32'hc1e0f67b, 32'hc2afb18b, 32'h4237424e, 32'hc2afe863, 32'hc21dc85d};
test_weights[35776:35783] = '{32'hc1acfc54, 32'h412ba2a7, 32'h41cbb785, 32'hc2b7227a, 32'hc2bcb25f, 32'h41cfde48, 32'h42c4e2b9, 32'h411610c3};
test_bias[4472:4472] = '{32'hc022abf4};
test_output[4472:4472] = '{32'h45d5934f};
test_input[35784:35791] = '{32'h4240b4c7, 32'h428cdaf2, 32'h42301e03, 32'hc29e7e5e, 32'hc229509a, 32'h41ce02a3, 32'hc29be411, 32'h42102291};
test_weights[35784:35791] = '{32'hc116e340, 32'hc27fb68b, 32'hc2104970, 32'h42c78060, 32'h4239fbdd, 32'hc2977328, 32'hc283a959, 32'h420f5961};
test_bias[4473:4473] = '{32'h4246b60b};
test_output[4473:4473] = '{32'hc639deb4};
test_input[35792:35799] = '{32'h4209bbd6, 32'hc1c7dcff, 32'h42943705, 32'hc20a8a16, 32'h428db9ae, 32'hc1b27194, 32'h42971ff2, 32'h4281513d};
test_weights[35792:35799] = '{32'hc28587d7, 32'hc21e9b44, 32'hc1b07684, 32'h42089ae8, 32'h42104982, 32'hc2923e4e, 32'h42a72b1c, 32'h40652ca7};
test_bias[4474:4474] = '{32'h4280c76b};
test_output[4474:4474] = '{32'h45d0889d};
test_input[35800:35807] = '{32'hc2bcbf47, 32'h42b69ea8, 32'h42bfffdc, 32'h42b234a4, 32'h420f5a92, 32'h42a4f617, 32'hc16d922f, 32'h42977452};
test_weights[35800:35807] = '{32'hc2b49e57, 32'h421d92c0, 32'hc2a41fa5, 32'h42b5c06f, 32'hc1769b60, 32'h42adb183, 32'hc267ef4d, 32'hc1aa9cb5};
test_bias[4475:4475] = '{32'hc2c2ee36};
test_output[4475:4475] = '{32'h468d64f4};
test_input[35808:35815] = '{32'h42915220, 32'hc2af3f0d, 32'hc28248fc, 32'h414f4bdd, 32'h41b051eb, 32'h427e6a7f, 32'hc0c1bc2a, 32'hc2680c95};
test_weights[35808:35815] = '{32'hc1cce3f2, 32'hc28fef61, 32'h42b8f902, 32'hc2bd8e6b, 32'h42886a55, 32'hc22d156f, 32'hc21c9d8d, 32'h41941974};
test_bias[4476:4476] = '{32'h42364f68};
test_output[4476:4476] = '{32'hc5977f0c};
test_input[35816:35823] = '{32'h42076ac1, 32'h4227ff2f, 32'hbf50643c, 32'h42195064, 32'hc2bee0c3, 32'hc224ede4, 32'hc24ea26e, 32'hc2a8093a};
test_weights[35816:35823] = '{32'hc2a5b431, 32'h40daee75, 32'h421c4b5d, 32'hc1c47f1e, 32'h4224dd1b, 32'h4228bcf1, 32'h416c2097, 32'hc29015fd};
test_bias[4477:4477] = '{32'h3fe56a63};
test_output[4477:4477] = '{32'hc571f6e6};
test_input[35824:35831] = '{32'hc13c69e1, 32'hc1ff27c9, 32'hc08a8918, 32'h4262e667, 32'h42ab3511, 32'h423a3453, 32'hc22d67ab, 32'h42a65515};
test_weights[35824:35831] = '{32'h4278891b, 32'hc22f3b49, 32'hc211f430, 32'hc2672033, 32'hc2c3e5a7, 32'h418f0ac1, 32'hc1414ab9, 32'hc25fc69b};
test_bias[4478:4478] = '{32'hc24460f0};
test_output[4478:4478] = '{32'hc65da246};
test_input[35832:35839] = '{32'h4211df62, 32'h41893c76, 32'hc2c43f27, 32'hc18df265, 32'h428b02f3, 32'hc2692fcc, 32'h422e7717, 32'hc21ed5ae};
test_weights[35832:35839] = '{32'h41583e1f, 32'hbef000e8, 32'h422016aa, 32'hc2462533, 32'hc2b4b712, 32'hc2817a78, 32'h428af319, 32'hc2c1cb14};
test_bias[4479:4479] = '{32'hc199b1a9};
test_output[4479:4479] = '{32'h44dfa11f};
test_input[35840:35847] = '{32'hc294e621, 32'hc2baffe3, 32'hc2092526, 32'hc0906279, 32'hc28742fb, 32'hc2ad6a4e, 32'hc20d95dc, 32'h4299fe1c};
test_weights[35840:35847] = '{32'h42b49dc0, 32'h423de0cd, 32'h405be11c, 32'h42b9e90c, 32'h41ac0b62, 32'h4297a5a6, 32'h41d00b75, 32'h4282d88a};
test_bias[4480:4480] = '{32'h429ef9bf};
test_output[4480:4480] = '{32'hc672ae66};
test_input[35848:35855] = '{32'hc1e252c4, 32'hc2506a11, 32'hc2b42640, 32'hc28cf6a3, 32'hc24fcbfc, 32'h41f8b0a4, 32'h422523b6, 32'h426ba163};
test_weights[35848:35855] = '{32'h40e67a30, 32'h411a8d9a, 32'hc2571775, 32'hc2a9d53b, 32'h4291d7c7, 32'h4230b7b5, 32'h42bd55d5, 32'hc1d6c922};
test_bias[4481:4481] = '{32'h41b15a47};
test_output[4481:4481] = '{32'h461d1ec0};
test_input[35856:35863] = '{32'h4295f0e5, 32'hc2b58ccf, 32'h41bee096, 32'hc0e16dc9, 32'h42c5561a, 32'h423b44f0, 32'h428a1268, 32'h429534fc};
test_weights[35856:35863] = '{32'h414392f7, 32'h421f00b0, 32'hc16118b3, 32'h42ae74d4, 32'hc2468dc2, 32'h427f3e34, 32'h42372d57, 32'h42890d5c};
test_bias[4482:4482] = '{32'hc283461c};
test_output[4482:4482] = '{32'h4525fad6};
test_input[35864:35871] = '{32'h424598e2, 32'hc230d296, 32'hc23cdf9d, 32'h42706de0, 32'hc1d29865, 32'h42bbcb26, 32'hc196ddaa, 32'hc18a571f};
test_weights[35864:35871] = '{32'h42b2c5b4, 32'hc22d160d, 32'hc21fe2f1, 32'h418de2c3, 32'hc2237d95, 32'hc0bd4de0, 32'hc26155c9, 32'hc20539a8};
test_bias[4483:4483] = '{32'hc2786831};
test_output[4483:4483] = '{32'h4631ca55};
test_input[35872:35879] = '{32'hc11873ff, 32'h41127e5c, 32'h423a71a5, 32'h4275a040, 32'hc17221d1, 32'h42a3f050, 32'hbe73968c, 32'h42152fc2};
test_weights[35872:35879] = '{32'hc1a072a2, 32'hc28c5232, 32'h42929b00, 32'hc1b774ea, 32'h4281d2b2, 32'h42c610b1, 32'hc2bca584, 32'hc256bb64};
test_bias[4484:4484] = '{32'hc2b2a305};
test_output[4484:4484] = '{32'h45cefbf3};
test_input[35880:35887] = '{32'h422e3efa, 32'h42a38602, 32'h425bd1f8, 32'h3f3d82ba, 32'hc2111e00, 32'hc1d61fff, 32'h42bf7f83, 32'hc29a2141};
test_weights[35880:35887] = '{32'h429c99e0, 32'h423f3b01, 32'hc2b73f94, 32'h42a158b6, 32'hc26cdcc6, 32'hc2928f04, 32'hc1ad4c28, 32'h42a95a47};
test_bias[4485:4485] = '{32'hc2892a12};
test_output[4485:4485] = '{32'hc50a6647};
test_input[35888:35895] = '{32'hc157a9c9, 32'hc202632b, 32'h4247d1c8, 32'hc2600863, 32'h410acd5f, 32'h4203cd23, 32'hc1e4b2f7, 32'h42836c8c};
test_weights[35888:35895] = '{32'hc1300c6e, 32'hc22f0171, 32'hc1c3deb0, 32'h42c63154, 32'hc11ac3f3, 32'hc1bcab0d, 32'hc250d6ee, 32'h4250612e};
test_bias[4486:4486] = '{32'h411d5970};
test_output[4486:4486] = '{32'hc48dc5c5};
test_input[35896:35903] = '{32'h4256a607, 32'hc2a305d4, 32'h4203a138, 32'hc2aab544, 32'h41eec62b, 32'hc26edd2b, 32'hc236a0ee, 32'hc20bcbfe};
test_weights[35896:35903] = '{32'h41e61eeb, 32'hc168113a, 32'h42597890, 32'h4290be45, 32'hc2bf47ee, 32'h4201edbe, 32'hc279344e, 32'h428135d3};
test_bias[4487:4487] = '{32'h42566341};
test_output[4487:4487] = '{32'hc5b5c29d};
test_input[35904:35911] = '{32'hc24e5076, 32'hc26af78f, 32'h4288a1d4, 32'hc0d0a5d3, 32'h422691fc, 32'hc26aefef, 32'h411ae7c9, 32'h42b5f3a8};
test_weights[35904:35911] = '{32'h428349ec, 32'h42a733bb, 32'h428e3f63, 32'h40432b41, 32'hc299f6e5, 32'hc17ee9f9, 32'h42a0bde0, 32'h427cc544};
test_bias[4488:4488] = '{32'h42625dc6};
test_output[4488:4488] = '{32'h445602a3};
test_input[35912:35919] = '{32'hc2b3d4b3, 32'hc200a0a2, 32'h42bd0c4e, 32'h41db826a, 32'h42962d83, 32'h41c89293, 32'hc18da1f1, 32'h428f6537};
test_weights[35912:35919] = '{32'hc1053abf, 32'hc2958293, 32'hc2bfb30e, 32'h42b9ea66, 32'h42788759, 32'h42b0dcf7, 32'hc1da8b48, 32'h426f5b11};
test_bias[4489:4489] = '{32'h4197c288};
test_output[4489:4489] = '{32'h4601fa75};
test_input[35920:35927] = '{32'h42c5c3a4, 32'hc28fb133, 32'h420a6fe4, 32'h42840748, 32'hc299e3e8, 32'h3fd0f85b, 32'hc28dff37, 32'hc2b1edf0};
test_weights[35920:35927] = '{32'h4295280f, 32'h41e0a36f, 32'h42bee7ab, 32'hc2b1b752, 32'h42c6e50d, 32'hc18180ae, 32'hc09a93c5, 32'hc2aa9a58};
test_bias[4490:4490] = '{32'h428596d2};
test_output[4490:4490] = '{32'h4542ad55};
test_input[35928:35935] = '{32'h4264c652, 32'hc29ca3e5, 32'hc20b59aa, 32'hc203b59a, 32'hc2033d83, 32'hc14bd33e, 32'hc1aa91df, 32'hc240cf95};
test_weights[35928:35935] = '{32'hc1f47f51, 32'h419a7ed0, 32'h42c6bffc, 32'h428f7c7e, 32'h4113243a, 32'h4049b308, 32'hc272fe04, 32'hc1c0e35d};
test_bias[4491:4491] = '{32'hc23ec7b8};
test_output[4491:4491] = '{32'hc5db473a};
test_input[35936:35943] = '{32'hc275b341, 32'h41b9e6de, 32'hc034000a, 32'hc2c61e07, 32'hc1b3e9ef, 32'hc2759547, 32'hc12472ac, 32'hc2b13c4a};
test_weights[35936:35943] = '{32'h4277814a, 32'hc184f97a, 32'hc0435fc5, 32'hc1acae93, 32'hc223d79e, 32'h428b09f0, 32'hc2004afb, 32'h4224cc41};
test_bias[4492:4492] = '{32'hc209f7c9};
test_output[4492:4492] = '{32'hc6089c5c};
test_input[35944:35951] = '{32'h422ac4cb, 32'hc1a21bce, 32'h42594497, 32'h40318fa3, 32'h42194449, 32'h418cd657, 32'h411c27e5, 32'h4284fd60};
test_weights[35944:35951] = '{32'h4282abcf, 32'hc2bdbe3a, 32'hc2991a9a, 32'hc2961ef2, 32'h42bfc450, 32'h40df6d80, 32'h4230debf, 32'h429447f2};
test_bias[4493:4493] = '{32'hc28d8dac};
test_output[4493:4493] = '{32'h4613641d};
test_input[35952:35959] = '{32'hc29f6e9a, 32'hc2846e35, 32'h40deb25a, 32'hc28f0b1e, 32'h4235a68c, 32'hc28f20d1, 32'hbf7e1949, 32'hc191bdd3};
test_weights[35952:35959] = '{32'hc002f528, 32'h427dfde2, 32'h42264e23, 32'hc29e3402, 32'hc1e01398, 32'h41f1ce00, 32'hc0c1bb72, 32'hc11714bd};
test_bias[4494:4494] = '{32'hbf892a87};
test_output[4494:4494] = '{32'hc4a91619};
test_input[35960:35967] = '{32'hc29f4bb8, 32'h42a935b9, 32'h414d9480, 32'h42042ef7, 32'hc25141cd, 32'h42644dd9, 32'hc26ccf35, 32'hc2057bb9};
test_weights[35960:35967] = '{32'hc2805a2c, 32'h422d366c, 32'h41efde05, 32'hc205883c, 32'h424474ae, 32'h42827614, 32'h40f0592c, 32'h422ec674};
test_bias[4495:4495] = '{32'hc22fa332};
test_output[4495:4495] = '{32'h45e30271};
test_input[35968:35975] = '{32'hc29934e5, 32'hc2305603, 32'hc25d96df, 32'hbfdd9802, 32'h421199ef, 32'hc2467c9c, 32'h42b1c091, 32'h42b67c1f};
test_weights[35968:35975] = '{32'hc281f87f, 32'hc06f8855, 32'h41e3b49f, 32'h412ca4be, 32'h425ab9de, 32'hc140c70d, 32'hc2264e9e, 32'hc1949677};
test_bias[4496:4496] = '{32'h42473f9d};
test_output[4496:4496] = '{32'h4446f6f3};
test_input[35976:35983] = '{32'hc241411a, 32'h42bc957d, 32'hc248c95d, 32'hc1aff148, 32'hc2a5ce49, 32'hc2b29a78, 32'h42b22330, 32'hc2861aa7};
test_weights[35976:35983] = '{32'hc282e28e, 32'h41cd3d80, 32'hc28c6d16, 32'h426ade70, 32'hc2a4431e, 32'hc2889c89, 32'hc2adfec4, 32'h4291ea94};
test_bias[4497:4497] = '{32'hc2a97b89};
test_output[4497:4497] = '{32'h45f9e934};
test_input[35984:35991] = '{32'h4073ee1d, 32'hc1b6686b, 32'h41742505, 32'hc22cd074, 32'hc1d63795, 32'hc13cc5a1, 32'h428e99bd, 32'h41a4b778};
test_weights[35984:35991] = '{32'hc2082621, 32'hc17cfd01, 32'hbfa05dbd, 32'h42a595e5, 32'hc2a5bbed, 32'h42afd295, 32'h42c5000f, 32'hc25f8360};
test_bias[4498:4498] = '{32'hc1880eef};
test_output[4498:4498] = '{32'h456580b3};
test_input[35992:35999] = '{32'hc1d2f95a, 32'hc288132e, 32'h4253a3b3, 32'h42bc50ea, 32'h4298933e, 32'h420d2318, 32'hc284d879, 32'hc2723cf3};
test_weights[35992:35999] = '{32'h42bbcae0, 32'hc12168a0, 32'hc28570ee, 32'hc2319302, 32'h42818ea7, 32'h42a49d62, 32'hc19cca8d, 32'hc02bf46e};
test_bias[4499:4499] = '{32'h42519d0d};
test_output[4499:4499] = '{32'hc309240e};
test_input[36000:36007] = '{32'hc2114490, 32'h41e904f1, 32'hc2c5cb7d, 32'hc2a813b8, 32'hc208b9ca, 32'hc2b9f005, 32'hc2786ab9, 32'h42b44ffe};
test_weights[36000:36007] = '{32'h41439147, 32'hbfe31dee, 32'h4152be01, 32'hc2581537, 32'h404ba94d, 32'hc13f4640, 32'hc13a5d1c, 32'h42a45f73};
test_bias[4500:4500] = '{32'h4280d8e3};
test_output[4500:4500] = '{32'h463a96b2};
test_input[36008:36015] = '{32'hc2924012, 32'h4232bfe2, 32'h428c5322, 32'hc28818da, 32'hc0ea2f10, 32'hc29348e1, 32'h41ca6398, 32'h42ad638a};
test_weights[36008:36015] = '{32'h427845a9, 32'h4265f667, 32'h42b4dcec, 32'hc2a732a3, 32'hc25a5b29, 32'h4292d99e, 32'hc2c1c323, 32'h4290953d};
test_bias[4501:4501] = '{32'hc251f53b};
test_output[4501:4501] = '{32'h4609d0aa};
test_input[36016:36023] = '{32'hc20808f6, 32'h40ae91ed, 32'hc24fc311, 32'h41ec612b, 32'hc200d4de, 32'h42987e96, 32'hc22c4df0, 32'h4268e5d2};
test_weights[36016:36023] = '{32'hc233fc1a, 32'hc09a2004, 32'hc1f193c6, 32'h42147c88, 32'h42282e1f, 32'hc23f4725, 32'h420181bd, 32'hc29a4818};
test_bias[4502:4502] = '{32'hc266e243};
test_output[4502:4502] = '{32'hc5d3b6d6};
test_input[36024:36031] = '{32'hc2a2f683, 32'hc1b277d6, 32'h417c6842, 32'hc12b2c2e, 32'hc260616a, 32'hc1eb198d, 32'hc2604b1a, 32'hc2245ca9};
test_weights[36024:36031] = '{32'h42c59c3f, 32'h415e8bf0, 32'h41422219, 32'h4091ae27, 32'hc28d4563, 32'hc206aa7d, 32'h42b25efc, 32'h42a847ba};
test_bias[4503:4503] = '{32'hc1c4fe71};
test_output[4503:4503] = '{32'hc637966e};
test_input[36032:36039] = '{32'hc2a2ff4e, 32'hc280c8a7, 32'h4218d57b, 32'hc0c74d6d, 32'h419e55bd, 32'h4007eee5, 32'hc2a4a775, 32'hc2a1b77e};
test_weights[36032:36039] = '{32'hc20cba0f, 32'hc2afe979, 32'h41664565, 32'h42205c1e, 32'hc2a62f5d, 32'h41bd9dfb, 32'h41eb1e1d, 32'hc0a3e47e};
test_bias[4504:4504] = '{32'h40f2bdf1};
test_output[4504:4504] = '{32'h45a3b86c};
test_input[36040:36047] = '{32'h42a28880, 32'h41c80d24, 32'h41bbd72b, 32'hc14df390, 32'hc28bcd90, 32'h40e08ca4, 32'h428bcde2, 32'hc1e55f5a};
test_weights[36040:36047] = '{32'h4205db54, 32'hc29184ea, 32'hc28df2cc, 32'h423072c3, 32'hc22492e9, 32'h41fd72f8, 32'hc2c6fccd, 32'h427462dc};
test_bias[4505:4505] = '{32'hc234f0cc};
test_output[4505:4505] = '{32'hc5da5db8};
test_input[36048:36055] = '{32'hc13b6513, 32'h428e995a, 32'hc2a3dd2c, 32'hc18492a8, 32'h421e04a4, 32'hbff6209a, 32'h4248327c, 32'hc2b9e465};
test_weights[36048:36055] = '{32'h40afec87, 32'h40b868df, 32'hc23e77f3, 32'hc2073d5e, 32'hc0b81a12, 32'hc08c3acf, 32'hc29b17ba, 32'h3ed387e1};
test_bias[4506:4506] = '{32'hc2669ad5};
test_output[4506:4506] = '{32'h441906b4};
test_input[36056:36063] = '{32'h4269c461, 32'hc1e71f52, 32'hc2202895, 32'hc21f6042, 32'hc2a4ed94, 32'hc256e60d, 32'h42add98d, 32'h41264ef6};
test_weights[36056:36063] = '{32'h41e3a931, 32'h42109ffb, 32'h42a3e779, 32'h4295064f, 32'hc2192ebe, 32'h418ebcad, 32'h428c968b, 32'h427bc3a7};
test_bias[4507:4507] = '{32'hc2832523};
test_output[4507:4507] = '{32'h454c2c19};
test_input[36064:36071] = '{32'hc0ad0c8a, 32'h42bc4c01, 32'hc02b4a59, 32'h42a09678, 32'h421409dc, 32'h4267da25, 32'h42b8951d, 32'h42adb17a};
test_weights[36064:36071] = '{32'hc1a06dc4, 32'hc26cebe4, 32'hc2706c2d, 32'h4108232b, 32'hc2af4b61, 32'h42c2ebe2, 32'hc2be690c, 32'h42c157da};
test_bias[4508:4508] = '{32'h41f35c55};
test_output[4508:4508] = '{32'hc5213334};
test_input[36072:36079] = '{32'hc23380c2, 32'hc1301c3a, 32'hc28a621f, 32'h4217b53b, 32'hc271754c, 32'h429340d7, 32'h4207143a, 32'hc107c328};
test_weights[36072:36079] = '{32'hc2219236, 32'h42c516b7, 32'h42bf1bad, 32'hc237d844, 32'hc25254b3, 32'hc244482e, 32'hc296ccae, 32'h4253198a};
test_bias[4509:4509] = '{32'hc2bede36};
test_output[4509:4509] = '{32'hc62e4bd2};
test_input[36080:36087] = '{32'h419116cc, 32'h40cab3ba, 32'hc275ff8e, 32'hb9b2d7fb, 32'h42707e05, 32'h42a362c2, 32'hc232f7d6, 32'hc29a2380};
test_weights[36080:36087] = '{32'h42c169b8, 32'hc12e74e5, 32'h426679a0, 32'hc270c38e, 32'hc25cf4ab, 32'hc1b56887, 32'hc188d12b, 32'hc119e05e};
test_bias[4510:4510] = '{32'hc24289b3};
test_output[4510:4510] = '{32'hc5ae346e};
test_input[36088:36095] = '{32'hc2045b69, 32'hc12acc80, 32'hc2b01c48, 32'h429e1521, 32'hc2b2619e, 32'h41e8c2d8, 32'h41e5af3b, 32'hc2a8ee0a};
test_weights[36088:36095] = '{32'h4040529c, 32'hc256f0d9, 32'hc21276c0, 32'h4188153d, 32'h427394c7, 32'h42a08202, 32'hc29ae074, 32'hc2033dcf};
test_bias[4511:4511] = '{32'h4283aa63};
test_output[4511:4511] = '{32'h452007fe};
test_input[36096:36103] = '{32'h42a64ae7, 32'h3eb8ee1f, 32'hc2c31379, 32'h423b3621, 32'hc1967094, 32'hc255e4d6, 32'h42a92969, 32'hc27d302d};
test_weights[36096:36103] = '{32'h429a8d8d, 32'h42020b79, 32'h42c5f7c1, 32'h411957b0, 32'hc23fc2fa, 32'h413c5a23, 32'hc20cc55d, 32'h42896eaa};
test_bias[4512:4512] = '{32'h41d94482};
test_output[4512:4512] = '{32'hc619107c};
test_input[36104:36111] = '{32'hc2367b68, 32'h42c00a3d, 32'hc1125719, 32'h428070e9, 32'h41711a7f, 32'hc2723e5b, 32'hc2c4d07b, 32'h428db4af};
test_weights[36104:36111] = '{32'hc1bcc439, 32'hc21f1bbb, 32'h4285d6c3, 32'h42c10621, 32'hc25b0bee, 32'h42ad2233, 32'h423dad9d, 32'hc1cb2234};
test_bias[4513:4513] = '{32'hc0fe6b1c};
test_output[4513:4513] = '{32'hc61788ae};
test_input[36112:36119] = '{32'hc296af5f, 32'h416b50fc, 32'h42a0e4c7, 32'hc02c524e, 32'h413f25e9, 32'hc2ae2081, 32'h42a31be3, 32'h42aea60a};
test_weights[36112:36119] = '{32'h4289467c, 32'h424e4cb9, 32'h422616dc, 32'hc25952b6, 32'h429362d6, 32'h42bde052, 32'hc29b473c, 32'h42a51a63};
test_bias[4514:4514] = '{32'h42336a3d};
test_output[4514:4514] = '{32'hc5e6ed25};
test_input[36120:36127] = '{32'h410d0441, 32'hc261bbab, 32'hc21b32f0, 32'h42bc23c7, 32'h4234ef2a, 32'h41b7982a, 32'h41e659f3, 32'h40ba1c8b};
test_weights[36120:36127] = '{32'h420b51ab, 32'hc21fc402, 32'h41c620e9, 32'h427a2cd5, 32'hc243b156, 32'hc213475b, 32'h42198311, 32'h41dc88f3};
test_bias[4515:4515] = '{32'hc280785a};
test_output[4515:4515] = '{32'h45afd60f};
test_input[36128:36135] = '{32'h429f0a30, 32'hc2c2cd43, 32'h42390a67, 32'h41ea54e1, 32'hc2a09b37, 32'h42915611, 32'hc1902a22, 32'h4225a81a};
test_weights[36128:36135] = '{32'hc1f6894e, 32'hc0af09f4, 32'h403a4455, 32'h42988faa, 32'h428bf6d9, 32'hc12e352a, 32'h41c77d7b, 32'hc2b8bfa9};
test_bias[4516:4516] = '{32'hc211e5c2};
test_output[4516:4516] = '{32'hc6207ce5};
test_input[36136:36143] = '{32'h4294424c, 32'h4202c803, 32'hc1c983ec, 32'hc0c85d48, 32'h40a03841, 32'h42900baa, 32'hc2aa7802, 32'hc0c95f02};
test_weights[36136:36143] = '{32'h42b5d3af, 32'h42800d3d, 32'h41e0a584, 32'hc2a83bac, 32'h41b83ccb, 32'h429d54ec, 32'hc2b35ea2, 32'hc22c461e};
test_bias[4517:4517] = '{32'h4289c3df};
test_output[4517:4517] = '{32'h46af227a};
test_input[36144:36151] = '{32'hc283b148, 32'hc27c7192, 32'h41e6dbd2, 32'hc192de47, 32'h4287abda, 32'h42919eb3, 32'hc2183d0a, 32'hc2a1e992};
test_weights[36144:36151] = '{32'h4068e0d3, 32'h41ff9eb3, 32'h418fccbe, 32'hc20e7af6, 32'hc226dd08, 32'h4244a808, 32'h4002a85c, 32'hc1cbe8ec};
test_bias[4518:4518] = '{32'h41d808d5};
test_output[4518:4518] = '{32'h44d1e2b4};
test_input[36152:36159] = '{32'hc28cc73f, 32'h42012100, 32'hc1797369, 32'hc21d6704, 32'h428ca454, 32'hc2bf6673, 32'hc13c4ee2, 32'hc293c0bd};
test_weights[36152:36159] = '{32'hc2c0cd20, 32'h425132cc, 32'h428e558c, 32'hc2134205, 32'hc2c5b5d3, 32'hc24e93a9, 32'h42b80522, 32'hc247f15d};
test_bias[4519:4519] = '{32'h41d06a67};
test_output[4519:4519] = '{32'h46137eee};
test_input[36160:36167] = '{32'h42b9d5ac, 32'hc1c9d524, 32'hc274eb29, 32'hc2967173, 32'h41949053, 32'hc20d2cc0, 32'hc2999dd6, 32'h429a947f};
test_weights[36160:36167] = '{32'h427fb521, 32'h4219acd3, 32'hc1185f0c, 32'h42699dad, 32'hc28877a8, 32'hbf7bea27, 32'h42a4c687, 32'hc2112688};
test_bias[4520:4520] = '{32'hc16c2e74};
test_output[4520:4520] = '{32'hc6100d8c};
test_input[36168:36175] = '{32'h42979944, 32'h41e0040a, 32'h4221056e, 32'h41d804b9, 32'h41467616, 32'hc0cc191b, 32'h42b6adc3, 32'hc10ad212};
test_weights[36168:36175] = '{32'hc29647a9, 32'h40fa8257, 32'h40ca2dd9, 32'hc1a8ccd7, 32'h423f8124, 32'hc21f322c, 32'hc25ab7cb, 32'h42a1b85e};
test_bias[4521:4521] = '{32'h4180e132};
test_output[4521:4521] = '{32'hc625ffad};
test_input[36176:36183] = '{32'hc265af4e, 32'hc2a24c66, 32'h421eddc6, 32'h42625d25, 32'h42929559, 32'h42b6d283, 32'h42c77b17, 32'h4140dfe5};
test_weights[36176:36183] = '{32'hc26245c9, 32'hc214862d, 32'hc1d7a131, 32'h42813f68, 32'hc2a53b55, 32'hc1bec810, 32'h429207d8, 32'h42a38089};
test_bias[4522:4522] = '{32'h428d5e0f};
test_output[4522:4522] = '{32'h460bdee3};
test_input[36184:36191] = '{32'hc288c7a9, 32'h42517ee1, 32'hc2bdcd85, 32'h42575470, 32'hc29f501c, 32'h427d486b, 32'h41a3132a, 32'hc2994d2c};
test_weights[36184:36191] = '{32'hc2b94446, 32'hc2bd9d82, 32'h4235a1b0, 32'hc23b77fc, 32'h42a54c0f, 32'hc254697d, 32'hc2290eec, 32'h429fe232};
test_bias[4523:4523] = '{32'hc1e12f34};
test_output[4523:4523] = '{32'hc6af3398};
test_input[36192:36199] = '{32'h428d096c, 32'hc2c51e99, 32'hc257582e, 32'hc0a53df7, 32'hc2393460, 32'hc286eef4, 32'h41d98954, 32'h42c0c5b5};
test_weights[36192:36199] = '{32'h40c34341, 32'hc0d428ae, 32'hc276c89c, 32'h42b41927, 32'hc2a75659, 32'h42b203ff, 32'hc2888d58, 32'hc1d103b2};
test_bias[4524:4524] = '{32'h4101e823};
test_output[4524:4524] = '{32'hc51fd997};
test_input[36200:36207] = '{32'h42a6e604, 32'h4221b3b0, 32'h41abe98c, 32'h3e9efe2b, 32'h42677b06, 32'h41b99491, 32'hc22598ce, 32'h40e5fc00};
test_weights[36200:36207] = '{32'h42ae3a53, 32'h4103f6ee, 32'hbfccdcb7, 32'h42a8d737, 32'h426b2c14, 32'hc2a4b24b, 32'hc278320c, 32'h42990898};
test_bias[4525:4525] = '{32'h42868d17};
test_output[4525:4525] = '{32'h463fc396};
test_input[36208:36215] = '{32'hbe651f9f, 32'h411e9e15, 32'h4155dd79, 32'hc17a1f38, 32'hc0fb2c42, 32'h427cf868, 32'h42803c1f, 32'hc29f68b0};
test_weights[36208:36215] = '{32'h42a13412, 32'h416a3828, 32'hc297ff66, 32'h41c7f4e7, 32'h4272f9d0, 32'hc1c5c9a5, 32'h41ad2a35, 32'hc21eb44e};
test_bias[4526:4526] = '{32'h41d7c7b0};
test_output[4526:4526] = '{32'h449d2af7};
test_input[36216:36223] = '{32'h421b7f39, 32'h41b28135, 32'hc2591320, 32'h417e2f00, 32'h428d6c9d, 32'hc1e7f715, 32'h4240689b, 32'hc2301dd9};
test_weights[36216:36223] = '{32'hc2a36364, 32'h42a8f26b, 32'hc2a3600a, 32'h4189a800, 32'hc28c1f9d, 32'h42a60d3b, 32'h42a82b25, 32'h40c5a62d};
test_bias[4527:4527] = '{32'h4295e22b};
test_output[4527:4527] = '{32'hc2c4f178};
test_input[36224:36231] = '{32'hc00d5271, 32'hc2261ddf, 32'h42b759e7, 32'h40ac9209, 32'hc1746105, 32'hc2404cf5, 32'h4201dfad, 32'hc28bff64};
test_weights[36224:36231] = '{32'hc0a7d7d8, 32'hc27c8343, 32'h42c7a2a1, 32'h418cb835, 32'hc121affe, 32'h41a9788c, 32'h4291dbfa, 32'hc28adfdc};
test_bias[4528:4528] = '{32'hc1f61607};
test_output[4528:4528] = '{32'h468e4918};
test_input[36232:36239] = '{32'hc12f2bd0, 32'h408d55ef, 32'hc244f8b4, 32'hc24a16fe, 32'hc2aceef9, 32'h42b31cb2, 32'hc2516c84, 32'hc2b7b194};
test_weights[36232:36239] = '{32'hc289d1a9, 32'hc1286b36, 32'hc2c78818, 32'hc23b4e76, 32'h4215cf4a, 32'hc2a130b8, 32'hc221229f, 32'hc2447ff6};
test_bias[4529:4529] = '{32'hc250f85a};
test_output[4529:4529] = '{32'h45801931};
test_input[36240:36247] = '{32'hc2a22938, 32'h42357346, 32'hc28fa63b, 32'hc2068d7c, 32'hc280aff6, 32'hc2155bce, 32'hc28ef67c, 32'hc1de17a7};
test_weights[36240:36247] = '{32'h427f9ea6, 32'hc2ae6fd0, 32'h42564bb5, 32'h418fedf2, 32'h42a10fde, 32'h428625ef, 32'hc11bd7b5, 32'hc278639c};
test_bias[4530:4530] = '{32'hc284ad30};
test_output[4530:4530] = '{32'hc693d6c2};
test_input[36248:36255] = '{32'hc0ac9eea, 32'h413db8f9, 32'hc2a3cd2a, 32'hc2bd349c, 32'hc281080f, 32'hc1f3b237, 32'hc20e1647, 32'h42af8b6a};
test_weights[36248:36255] = '{32'h42564717, 32'h4214a553, 32'hc1b5d660, 32'h421cc08f, 32'hc2bd319d, 32'hc2a60571, 32'hc2883ee9, 32'h41a95045};
test_bias[4531:4531] = '{32'h42a56670};
test_output[4531:4531] = '{32'h46308726};
test_input[36256:36263] = '{32'h4274b273, 32'h41805180, 32'h40a71b06, 32'hc257b922, 32'hc298253c, 32'hc1fcacfd, 32'hc1b4925e, 32'h42c18450};
test_weights[36256:36263] = '{32'h415ec432, 32'h422057bc, 32'h413298ac, 32'h42b583e0, 32'h42bf9276, 32'hc28cf477, 32'hc28a69ee, 32'h3f062657};
test_bias[4532:4532] = '{32'hc29cb721};
test_output[4532:4532] = '{32'hc5d69f50};
test_input[36264:36271] = '{32'h4239f6f7, 32'h4248795c, 32'h422badd3, 32'h42a2c179, 32'h4289ea93, 32'hc2116d4b, 32'hc188d9c9, 32'h41ec7a8b};
test_weights[36264:36271] = '{32'h425ae90a, 32'hc18b9af6, 32'h428ddbd8, 32'h4275c822, 32'h4274dd24, 32'h40cbc4c9, 32'h4274651a, 32'hc27f9f21};
test_bias[4533:4533] = '{32'hc211353f};
test_output[4533:4533] = '{32'h4627b68b};
test_input[36272:36279] = '{32'hc1c636e1, 32'hc2a65424, 32'hc220ccdc, 32'h4286b7e2, 32'hc28818cb, 32'hc181de72, 32'h410ab53b, 32'hc2a4c159};
test_weights[36272:36279] = '{32'hc2b19fb0, 32'hc260f0de, 32'hc2343dab, 32'hc2ada84d, 32'hc0219e57, 32'hc1c227c6, 32'hc1c61f3d, 32'hc2be50bf};
test_bias[4534:4534] = '{32'hc2b277cb};
test_output[4534:4534] = '{32'h462af2db};
test_input[36280:36287] = '{32'h429b08f5, 32'h42743842, 32'hc2b27f2c, 32'hc20c1182, 32'hc2631eeb, 32'h4286c8b1, 32'hc2b99830, 32'hc011127c};
test_weights[36280:36287] = '{32'hc2b718fd, 32'hc27721de, 32'h425215ec, 32'hc2bcc99d, 32'h42bb233e, 32'h41e41f90, 32'hc2ab97f6, 32'hc1fb732e};
test_bias[4535:4535] = '{32'h4291665c};
test_output[4535:4535] = '{32'hc5eb82c0};
test_input[36288:36295] = '{32'h4292d5dc, 32'hc24fbab4, 32'hc2956001, 32'h42a427a2, 32'h42c6f533, 32'hc0d66cb2, 32'h42bdcb68, 32'hc19443f3};
test_weights[36288:36295] = '{32'hc257f67a, 32'hc1bc4c1f, 32'h42553754, 32'h427146c9, 32'hc2922e57, 32'h42bb3871, 32'hc2c268ec, 32'hc184dd24};
test_bias[4536:4536] = '{32'hbf0816c8};
test_output[4536:4536] = '{32'hc6913690};
test_input[36296:36303] = '{32'hc2baa3cd, 32'h42956632, 32'h41c770e4, 32'h420067dc, 32'hc2a0469e, 32'hc28cd524, 32'h411030d9, 32'hc2038a2e};
test_weights[36296:36303] = '{32'hc2a5e4e6, 32'hc23afe38, 32'h40fe70e2, 32'hc16c87a7, 32'h4220e234, 32'hc29c4ed3, 32'hc20b29f7, 32'hc0b0d3a4};
test_bias[4537:4537] = '{32'hc0f7490f};
test_output[4537:4537] = '{32'h45bf0605};
test_input[36304:36311] = '{32'h42264706, 32'hc24c8059, 32'hc229a2d7, 32'hc28960f1, 32'h4266032b, 32'h429aa9b9, 32'hc1c6a64f, 32'h429dffeb};
test_weights[36304:36311] = '{32'h4034fd8e, 32'hc04e4234, 32'hc1c69505, 32'hc25038b7, 32'h42a7d310, 32'h4246f516, 32'hc28a6fb6, 32'h42a5d964};
test_bias[4538:4538] = '{32'h41a036bd};
test_output[4538:4538] = '{32'h46aae048};
test_input[36312:36319] = '{32'h4202233c, 32'h405feaed, 32'hc2c6dc06, 32'h42c0ad67, 32'h41af391c, 32'hc29a300d, 32'hc21c9781, 32'h41fc2ae5};
test_weights[36312:36319] = '{32'hc285a40a, 32'hc2c72beb, 32'h42be28bd, 32'h420486e0, 32'hc2bc43b5, 32'h41b0393f, 32'hc2bb7325, 32'hc29dab44};
test_bias[4539:4539] = '{32'hc2b0a1b5};
test_output[4539:4539] = '{32'hc632e16e};
test_input[36320:36327] = '{32'h40e4be18, 32'h429f5977, 32'h421c09ba, 32'hc23e98a3, 32'h42c1e246, 32'h401d5293, 32'hc2aa5b01, 32'h41d38652};
test_weights[36320:36327] = '{32'h42434e71, 32'h42b60921, 32'h419d7cfb, 32'h42ad85af, 32'hc1febb48, 32'hc2a217eb, 32'hc1ce1951, 32'h42916582};
test_bias[4540:4540] = '{32'hc29a3cda};
test_output[4540:4540] = '{32'h459be131};
test_input[36328:36335] = '{32'hc0f9c051, 32'h428f3baa, 32'hc2b31234, 32'hc2675f82, 32'h4283bb76, 32'hc2ad9037, 32'h40d260ae, 32'hc2a4a0d1};
test_weights[36328:36335] = '{32'h42740e34, 32'hc24daff3, 32'hc02918f5, 32'h4111315a, 32'h42bef8d0, 32'hc22100b7, 32'h429792ef, 32'h42c19a75};
test_bias[4541:4541] = '{32'h42a767c3};
test_output[4541:4541] = '{32'hc5003105};
test_input[36336:36343] = '{32'h42821ee5, 32'h4298d7f3, 32'hc28fd2be, 32'hc1eefbfb, 32'h41e03c0b, 32'h41c490d3, 32'hc292593f, 32'h41c78e97};
test_weights[36336:36343] = '{32'hc103e92c, 32'h42bc9ac8, 32'h4244ffc1, 32'hc246d62b, 32'h4000084b, 32'hc2c4ecbf, 32'h426bb871, 32'h421486d0};
test_bias[4542:4542] = '{32'hc191464b};
test_output[4542:4542] = '{32'hc49033b1};
test_input[36344:36351] = '{32'h42b54511, 32'h41b83a7f, 32'hc2937000, 32'hc1343e5a, 32'h42c1fc02, 32'h420d05da, 32'hc2909f2d, 32'hc238d74c};
test_weights[36344:36351] = '{32'h42354855, 32'h427f02d9, 32'hc1b8e8a8, 32'h4267b9a4, 32'h42a332a5, 32'h425bfadd, 32'hc27723ac, 32'h42adec1c};
test_bias[4543:4543] = '{32'hc2332eee};
test_output[4543:4543] = '{32'h4683e9aa};
test_input[36352:36359] = '{32'h41d6c36f, 32'h42a0e647, 32'h40f9c62a, 32'h42305ccb, 32'hc27e23b7, 32'h4272e151, 32'hc26737f0, 32'hc1f38f82};
test_weights[36352:36359] = '{32'h425037ee, 32'h41ac9f2b, 32'hbed30bf5, 32'hc267eaeb, 32'h421724c3, 32'h42c46a95, 32'hc2a68e55, 32'h42367bd9};
test_bias[4544:4544] = '{32'h42929e6f};
test_output[4544:4544] = '{32'h45ee93f6};
test_input[36360:36367] = '{32'h41da9976, 32'h42c0fc80, 32'hc27ada1d, 32'h42c662c3, 32'h4284f1f0, 32'hc28bd203, 32'hc1c221eb, 32'h428238e3};
test_weights[36360:36367] = '{32'hc2bdf5ee, 32'hc1907bf5, 32'hc20bd697, 32'hc2b6c2db, 32'hc20a8305, 32'h4251fdec, 32'h41e2bcb8, 32'hc29b659f};
test_bias[4545:4545] = '{32'h422b092e};
test_output[4545:4545] = '{32'hc6b2cbd9};
test_input[36368:36375] = '{32'hbe1d5ac8, 32'hc1f3aa6b, 32'hc273514b, 32'h42a3ef81, 32'hc1407af4, 32'h427735b0, 32'h42bc034f, 32'hc2892ad3};
test_weights[36368:36375] = '{32'h40e3c044, 32'h426c21b0, 32'hc23057bf, 32'h420a0175, 32'h4102e9d9, 32'h419fc448, 32'h41adc17d, 32'hc1823153};
test_bias[4546:4546] = '{32'h41fd8b49};
test_output[4546:4546] = '{32'h45fb1ff8};
test_input[36376:36383] = '{32'h421d3d7e, 32'hc2b8f60b, 32'h42af1129, 32'hc164ee61, 32'h3f7ca8c3, 32'hc158dbb6, 32'hc21a8311, 32'hc1560bc4};
test_weights[36376:36383] = '{32'hc253d414, 32'hc29cd8c3, 32'hc230f59a, 32'hc0fec79c, 32'h42b82d11, 32'h41331778, 32'hc28de281, 32'h42c7d171};
test_bias[4547:4547] = '{32'h42917cc5};
test_output[4547:4547] = '{32'h4530c0d8};
test_input[36384:36391] = '{32'hc2759473, 32'hc2a6153b, 32'hc2025f85, 32'h4242ac1d, 32'hc246dc77, 32'h42c19bce, 32'hc284930e, 32'hc29d1c0e};
test_weights[36384:36391] = '{32'h42a7cb32, 32'hc29673d1, 32'h428f6f6b, 32'hc05ec3b9, 32'hc2afa679, 32'h40ef9d7f, 32'h429b3887, 32'h41374f8c};
test_bias[4548:4548] = '{32'hc0c62d55};
test_output[4548:4548] = '{32'hc514281f};
test_input[36392:36399] = '{32'h3f2559eb, 32'h41a1229c, 32'h41ad1c53, 32'hc1ae8f49, 32'h40e812fc, 32'hc0b46b92, 32'hc27bb152, 32'hc2858eef};
test_weights[36392:36399] = '{32'h422ccb84, 32'h4287175d, 32'hc28d7b7c, 32'h41b12bb5, 32'hc117c64b, 32'h42973714, 32'h41f4840a, 32'h425071f2};
test_bias[4549:4549] = '{32'hc2096311};
test_output[4549:4549] = '{32'hc5ccf16a};
test_input[36400:36407] = '{32'hc139e297, 32'h42aa2c7c, 32'hc26b0497, 32'h42965ec2, 32'hc2194290, 32'h413923c6, 32'hc18e56ba, 32'hc275084a};
test_weights[36400:36407] = '{32'hc216659b, 32'hc293c628, 32'hc26a479e, 32'hc2a82bd4, 32'hc2a4d8e3, 32'hc283fd9d, 32'h421f8643, 32'hc09f9297};
test_bias[4550:4550] = '{32'h41d99858};
test_output[4550:4550] = '{32'hc5d1c9cd};
test_input[36408:36415] = '{32'hc26b3032, 32'hc2384d8e, 32'h42c63740, 32'hc27cb228, 32'h418fd887, 32'h42a12c99, 32'hc260859d, 32'hc08d4fa5};
test_weights[36408:36415] = '{32'h4142c19a, 32'h42865d08, 32'hc2687067, 32'h410bcd6f, 32'h41def4e2, 32'hc29b00b7, 32'h41049615, 32'h4286859d};
test_bias[4551:4551] = '{32'h42218b5f};
test_output[4551:4551] = '{32'hc6819913};
test_input[36416:36423] = '{32'hc21a8239, 32'hc2821192, 32'h425c5827, 32'hc1cc143f, 32'h42b1490e, 32'h405980b1, 32'h4243d1b4, 32'hc2a5e873};
test_weights[36416:36423] = '{32'hc22ffef5, 32'h4235c083, 32'h4049cc6d, 32'hc2225177, 32'hc0088e71, 32'hc22aa348, 32'hc180a13f, 32'hc23d5112};
test_bias[4552:4552] = '{32'hc2808ad1};
test_output[4552:4552] = '{32'h45286070};
test_input[36424:36431] = '{32'h41e20739, 32'hc2ba7ff3, 32'hc0964480, 32'h41f4c4ec, 32'hc2ba26b3, 32'h4271da97, 32'h42bd8583, 32'hc2a331c1};
test_weights[36424:36431] = '{32'hc1530f19, 32'h41a3310d, 32'h42c17680, 32'h408fee51, 32'hc1c823be, 32'hc2b0261f, 32'hc20ca716, 32'h42acc30f};
test_bias[4553:4553] = '{32'hc26b64b5};
test_output[4553:4553] = '{32'hc67a6eb0};
test_input[36432:36439] = '{32'hc27d7103, 32'hc2bffd0c, 32'h421887ed, 32'h4296951f, 32'h42140bc4, 32'h41c14ddf, 32'hc261ffee, 32'h42892460};
test_weights[36432:36439] = '{32'h422a95df, 32'h42a6fe2a, 32'hc1a2421c, 32'h410558c0, 32'h41f953d9, 32'hc2068b0a, 32'hc201015d, 32'hc2a965f2};
test_bias[4554:4554] = '{32'h3ea61032};
test_output[4554:4554] = '{32'hc662af47};
test_input[36440:36447] = '{32'h415003ed, 32'h42be69e2, 32'hc2a2b017, 32'h428b4a6e, 32'hc242f527, 32'h42a7cceb, 32'h42600333, 32'hc2c24649};
test_weights[36440:36447] = '{32'hc27d1c2a, 32'h42a55037, 32'hc2a26b6c, 32'h42ba0ae6, 32'h428eb117, 32'hc235984b, 32'hc2aafb67, 32'h42bef276};
test_bias[4555:4555] = '{32'hc2b2a2f9};
test_output[4555:4555] = '{32'hc4a346aa};
test_input[36448:36455] = '{32'hc2261b1a, 32'h417e212f, 32'h42b13fbe, 32'h4207a0a7, 32'hc1b87c7b, 32'hc2b01ba5, 32'h42b5883b, 32'h4116b3d2};
test_weights[36448:36455] = '{32'hc1c0805b, 32'hc2c4c518, 32'h4207764d, 32'h42a7eace, 32'h4278e1d1, 32'h4274d203, 32'hc2449ff0, 32'h42ba76f4};
test_bias[4556:4556] = '{32'hc0e01d43};
test_output[4556:4556] = '{32'hc5a050de};
test_input[36456:36463] = '{32'h4290c3b5, 32'h3fd05572, 32'h42c6c959, 32'h41d91ba4, 32'hc2426170, 32'hc252b71f, 32'h40162c43, 32'h4182a67c};
test_weights[36456:36463] = '{32'hc2a07c15, 32'h42b4d4b5, 32'h4154ed74, 32'h425727ca, 32'hc237bcfb, 32'h40756cc7, 32'h42004f0b, 32'hc27c7222};
test_bias[4557:4557] = '{32'hc2a6e390};
test_output[4557:4557] = '{32'hc4ebe57c};
test_input[36464:36471] = '{32'h40f21578, 32'h4214b023, 32'h42555cac, 32'hc0dd838c, 32'h424c2232, 32'hc296f86f, 32'h42a30d24, 32'hc2a8d224};
test_weights[36464:36471] = '{32'h429a4429, 32'h4226bf06, 32'h42abb8a8, 32'hc2b05b96, 32'hc28bb14c, 32'h42b64b54, 32'hc0f9205a, 32'h40a273bd};
test_bias[4558:4558] = '{32'hc22ee472};
test_output[4558:4558] = '{32'hc58422c2};
test_input[36472:36479] = '{32'hc18cabe7, 32'hbfa4a065, 32'h420065fe, 32'hc29f0c15, 32'hc212ac74, 32'hc20b86ad, 32'h4261927c, 32'hc21ea3b4};
test_weights[36472:36479] = '{32'h424e0490, 32'hc279d0e7, 32'h42c4f6c5, 32'h42317b86, 32'h42c590dc, 32'h3ea953fc, 32'hc1deda9d, 32'h417ad306};
test_bias[4559:4559] = '{32'h4195dc21};
test_output[4559:4559] = '{32'hc5dac23a};
test_input[36480:36487] = '{32'h41fb956e, 32'h41250104, 32'h42561aca, 32'hc25bde15, 32'hc2a1329b, 32'h4104cd85, 32'hc2982665, 32'hc21ed5fe};
test_weights[36480:36487] = '{32'h42995f03, 32'hc0f08df4, 32'h42b389a7, 32'h428c0af2, 32'h41d21947, 32'h42b02c27, 32'h41ba0039, 32'hc1644f13};
test_bias[4560:4560] = '{32'h40cd9be0};
test_output[4560:4560] = '{32'h44313aa3};
test_input[36488:36495] = '{32'hc28f0ddf, 32'h40c1c779, 32'hc1ac6539, 32'h422810af, 32'h420f5974, 32'h42c334e8, 32'hc185bd52, 32'hc279e8a4};
test_weights[36488:36495] = '{32'h41dab904, 32'h4234a60a, 32'h42475bdb, 32'hc1b67351, 32'hc24dead8, 32'hc1a872bc, 32'h3ff49c0a, 32'h41b6a5a5};
test_bias[4561:4561] = '{32'h40e8124d};
test_output[4561:4561] = '{32'hc60da5e2};
test_input[36496:36503] = '{32'h422519c8, 32'hc275aeda, 32'hc11fff1b, 32'h42214ed8, 32'hc2b2ce9f, 32'h42bad598, 32'hc20c406a, 32'h4220e381};
test_weights[36496:36503] = '{32'h429424e1, 32'h412097c6, 32'hc299d1c7, 32'h41f3cc20, 32'hc1f48abb, 32'hc202826c, 32'hc29159bc, 32'hc294ff2f};
test_bias[4562:4562] = '{32'h428520cf};
test_output[4562:4562] = '{32'h4569e136};
test_input[36504:36511] = '{32'hc23411c9, 32'hc2a0493d, 32'hc29a032f, 32'hc27fc14b, 32'hc1ed42fa, 32'h42432c8e, 32'h416b1055, 32'h4222332a};
test_weights[36504:36511] = '{32'hc2658447, 32'hc0799dd8, 32'h41d5b465, 32'h41d62c05, 32'h41af9cd4, 32'hc04a1d07, 32'hc1e13312, 32'hc29fcc0e};
test_bias[4563:4563] = '{32'h42b0d4c2};
test_output[4563:4563] = '{32'hc5a3daa0};
test_input[36512:36519] = '{32'hc1fea03d, 32'hc2b11f38, 32'hc245cda1, 32'h42b8198e, 32'h4283ec9d, 32'h429e2d31, 32'h428afa4f, 32'h426d4217};
test_weights[36512:36519] = '{32'hc216ffb4, 32'h4189410d, 32'hc25cbe4e, 32'h4264237e, 32'h423999f4, 32'h4237ad1b, 32'hc24bb22d, 32'hc185f903};
test_bias[4564:4564] = '{32'hc21a8454};
test_output[4564:4564] = '{32'h4618db56};
test_input[36520:36527] = '{32'hc264e65f, 32'hc1354c29, 32'h4239257a, 32'hc198aff8, 32'h427e78c1, 32'h41c977a2, 32'h42b6af08, 32'h3fba5984};
test_weights[36520:36527] = '{32'hc1f9906b, 32'hc261209f, 32'h41bf035e, 32'h417c2711, 32'h4274a60f, 32'h41d2c1c6, 32'hbf9437d7, 32'hc2bd5074};
test_bias[4565:4565] = '{32'h428ed624};
test_output[4565:4565] = '{32'h45edcca3};
test_input[36528:36535] = '{32'h42a8ad16, 32'hc0d234a3, 32'h42a10075, 32'h41c32772, 32'h410dc1da, 32'hc01d27fe, 32'hc27944a9, 32'hc1c8920f};
test_weights[36528:36535] = '{32'h42b97250, 32'hc2844775, 32'hc2c04456, 32'hc2278708, 32'hc25e5f10, 32'h427d0eee, 32'h42818562, 32'hc29c2f2b};
test_bias[4566:4566] = '{32'hc17569ea};
test_output[4566:4566] = '{32'hc54aefc3};
test_input[36536:36543] = '{32'hc2afc527, 32'h42b4dfe0, 32'hc253ff0e, 32'h41cddf7d, 32'hc288f9c4, 32'h420846b6, 32'hc24ac5e9, 32'h42a72927};
test_weights[36536:36543] = '{32'h418d3507, 32'hc2a093ed, 32'h424d04e2, 32'hc2b903e1, 32'h42a7892d, 32'hc26e2c8c, 32'h42532bcf, 32'hc2bf818d};
test_bias[4567:4567] = '{32'h42bb9dbd};
test_output[4567:4567] = '{32'hc6fc0931};
test_input[36544:36551] = '{32'h42867f30, 32'hc18bada9, 32'h41f81c78, 32'h42ab3700, 32'h425035f2, 32'h41b6f621, 32'hc0047351, 32'hc1e038a9};
test_weights[36544:36551] = '{32'hc2a6cf23, 32'hc1ad7ded, 32'hc2a97c89, 32'hc1a2c343, 32'hc23e1593, 32'hc2c05d2a, 32'hc22b1c96, 32'hbfc2e6d4};
test_bias[4568:4568] = '{32'h42246ac1};
test_output[4568:4568] = '{32'hc65c5466};
test_input[36552:36559] = '{32'h422bfcf5, 32'h42a5d82d, 32'hc2075c79, 32'h42383e5e, 32'hc2b9360a, 32'h42a3cdc8, 32'hc2411ca9, 32'hc2a84478};
test_weights[36552:36559] = '{32'h41f722e1, 32'h42ae10d6, 32'h40fafd5b, 32'hc21001f2, 32'h42803228, 32'h4282ef46, 32'h41b39647, 32'h42b81da3};
test_bias[4569:4569] = '{32'h41c3cffb};
test_output[4569:4569] = '{32'hc52c4dd4};
test_input[36560:36567] = '{32'hc2b014dc, 32'h42bef1f4, 32'h408d7f32, 32'h42c757cb, 32'hc274b7e7, 32'h41db93cb, 32'h42851ce7, 32'hc2954fba};
test_weights[36560:36567] = '{32'h42b224c4, 32'hc29ed33b, 32'h42babac9, 32'h415d734d, 32'hc2a7f3da, 32'h417a2ac6, 32'h422ed23e, 32'hc28a69e5};
test_bias[4570:4570] = '{32'hc1fe25c2};
test_output[4570:4570] = '{32'hc1a5f1be};
test_input[36568:36575] = '{32'hc122b3fc, 32'hc1b8a1fc, 32'h4253e3f4, 32'h4211ffb3, 32'hc2856ed5, 32'h42c48e51, 32'hc24a5f6b, 32'hc22e1f38};
test_weights[36568:36575] = '{32'hc1ebb5b6, 32'h42b77190, 32'h4243dc80, 32'hc20838fd, 32'hc2b26671, 32'h420c632d, 32'h41d9dc1d, 32'h427f8730};
test_bias[4571:4571] = '{32'h42b33c12};
test_output[4571:4571] = '{32'h4598078f};
test_input[36576:36583] = '{32'hc29b3579, 32'hc2319337, 32'h41d7e98d, 32'h4263c789, 32'hc281a8b6, 32'h42adae73, 32'h41ecb0c1, 32'h42a1b6f4};
test_weights[36576:36583] = '{32'hc2bafd7a, 32'hc280f406, 32'hc1b8a821, 32'h42aabd72, 32'h424b3b0c, 32'hc2b65f4e, 32'h41c509b2, 32'hc06434bf};
test_bias[4572:4572] = '{32'hc2c12058};
test_output[4572:4572] = '{32'h4559fbac};
test_input[36584:36591] = '{32'hc2c446be, 32'hc2b44009, 32'h40a1102b, 32'h4217d4c8, 32'h4253302f, 32'hc294dc01, 32'hc2a858cf, 32'h4222c2ca};
test_weights[36584:36591] = '{32'h4282e5e4, 32'h4187871f, 32'hc1c6990b, 32'hc27ffa57, 32'hc286caf2, 32'h4184c43e, 32'hc18a364f, 32'h42955af2};
test_bias[4573:4573] = '{32'hc2865a3b};
test_output[4573:4573] = '{32'hc629defa};
test_input[36592:36599] = '{32'hc261e900, 32'hc173af18, 32'hc26fc05d, 32'hc1069b23, 32'h3f96a05f, 32'h4277c67f, 32'hc1db1cda, 32'hc2b3b8f9};
test_weights[36592:36599] = '{32'hc130477e, 32'h42607981, 32'hc245c5ec, 32'hc213e5b1, 32'hc2ae3bd2, 32'hc1c5877e, 32'hc2b8ffea, 32'h41caca98};
test_bias[4574:4574] = '{32'h41f58b6d};
test_output[4574:4574] = '{32'h44d40ddb};
test_input[36600:36607] = '{32'hc2c589c1, 32'h4278e4f0, 32'h4280f244, 32'hc2828556, 32'hc254c62e, 32'hc239ef20, 32'hc210867f, 32'h42a04206};
test_weights[36600:36607] = '{32'h427ac9a5, 32'h41bb7937, 32'hc2a22520, 32'hc1dad4d8, 32'h429a44cc, 32'h418df410, 32'h41c4b064, 32'h42af0931};
test_bias[4575:4575] = '{32'h42c1cf31};
test_output[4575:4575] = '{32'hc5d7165b};
test_input[36608:36615] = '{32'hc188f0b9, 32'h41beb7c4, 32'hc0b0455b, 32'hc1a83ec6, 32'hc25be2ac, 32'hc28837f6, 32'hc28385e9, 32'hc28dff37};
test_weights[36608:36615] = '{32'hc257e2cf, 32'hc1d2222f, 32'h41b0c70e, 32'hc15e1d84, 32'h4297b8ff, 32'h4186f33d, 32'h42599987, 32'hc2a97280};
test_bias[4576:4576] = '{32'hc0d60aa3};
test_output[4576:4576] = '{32'hc517415e};
test_input[36616:36623] = '{32'hc21256de, 32'hc1ec6ecb, 32'hc129142b, 32'hc0bb1e31, 32'hc20911f8, 32'hc2ad2349, 32'hbfb2cafc, 32'h41f67de2};
test_weights[36616:36623] = '{32'h4033809e, 32'hc24d0005, 32'hc1f17e91, 32'h427ed4ea, 32'h42a4f1ca, 32'hc2928915, 32'hc19566c6, 32'h3fa0504a};
test_bias[4577:4577] = '{32'h42914f52};
test_output[4577:4577] = '{32'h459ca365};
test_input[36624:36631] = '{32'h41db4400, 32'hc1f106c9, 32'h4270c0e2, 32'h42c7b439, 32'h429519f5, 32'h423ff5d0, 32'h425e2e6d, 32'h41a809eb};
test_weights[36624:36631] = '{32'hc2b987b4, 32'hc2aa487e, 32'hc26f90cc, 32'h418e99bc, 32'h41853747, 32'hc10ddba6, 32'h42088ccc, 32'hc19d96e9};
test_bias[4578:4578] = '{32'hc1b88654};
test_output[4578:4578] = '{32'h43ec83b7};
test_input[36632:36639] = '{32'hc243de88, 32'h41515f73, 32'h42aacd2e, 32'hc2181f42, 32'h41c0a021, 32'h4259d149, 32'h42b80a1a, 32'h4258c42d};
test_weights[36632:36639] = '{32'h40b37ab0, 32'h427bdb1c, 32'hc0718df7, 32'h41329010, 32'hc294d887, 32'hc1e05d79, 32'h42954bd8, 32'h413a2918};
test_bias[4579:4579] = '{32'h40c9ffda};
test_output[4579:4579] = '{32'h457954b0};
test_input[36640:36647] = '{32'h417f2b0e, 32'h428b70fd, 32'hc2112bfc, 32'hc11bbdd0, 32'hc1c022ef, 32'h42ad2817, 32'hc281b562, 32'hc257beb1};
test_weights[36640:36647] = '{32'hc2b4b39b, 32'hc0d33c9b, 32'hc23aac94, 32'hc21ee427, 32'h42c39612, 32'h3f8f3a31, 32'h427c0395, 32'h4204374c};
test_bias[4580:4580] = '{32'hc19b0ae6};
test_output[4580:4580] = '{32'hc5f8c688};
test_input[36648:36655] = '{32'h41ae4019, 32'h42a36d55, 32'hc0a371f3, 32'h42b08919, 32'h419bbdb6, 32'h4292b77a, 32'hc264188b, 32'h42980794};
test_weights[36648:36655] = '{32'h42bcba70, 32'h428fc7fb, 32'h41ba6288, 32'h4292d60e, 32'h4271fc9b, 32'hc04637bf, 32'hc27e4f03, 32'hc2611d10};
test_bias[4581:4581] = '{32'h422a3fd0};
test_output[4581:4581] = '{32'h46649f1d};
test_input[36656:36663] = '{32'h422d9d59, 32'hc284ab56, 32'h3f4c8a05, 32'h42b04a8c, 32'h42611fe8, 32'h41d9f217, 32'h42754a16, 32'hc27b8130};
test_weights[36656:36663] = '{32'hc2bbc277, 32'hc253848d, 32'hc27232d7, 32'h42987e22, 32'h426dae94, 32'h41a67db7, 32'hc2375fa3, 32'hc170d11a};
test_bias[4582:4582] = '{32'h42c10726};
test_output[4582:4582] = '{32'h4600e11e};
test_input[36664:36671] = '{32'hc197a995, 32'h429358f0, 32'h4219f161, 32'h4210e116, 32'hc279b7a4, 32'hc21ecdda, 32'h42297c28, 32'hc262d6fc};
test_weights[36664:36671] = '{32'hc2a75698, 32'h429f264d, 32'h416fcc97, 32'h42b5394c, 32'h42418283, 32'hc2ad6015, 32'h4231d23b, 32'h419a70fa};
test_bias[4583:4583] = '{32'hc18017c5};
test_output[4583:4583] = '{32'h464356f6};
test_input[36672:36679] = '{32'h41b662bc, 32'h3fe7c471, 32'h42257641, 32'hc1c3887b, 32'hc123d9df, 32'hc0ac4743, 32'h414ffea5, 32'h429b0da0};
test_weights[36672:36679] = '{32'h40829739, 32'hc2819abe, 32'h41fe8610, 32'h4216db4f, 32'h41dec706, 32'hc242fde6, 32'hc13c9d6c, 32'hc2327dad};
test_bias[4584:4584] = '{32'hc1aafc9d};
test_output[4584:4584] = '{32'hc54d6d49};
test_input[36680:36687] = '{32'h425e237c, 32'h42a45de3, 32'hc1a16f4e, 32'hc298738e, 32'h4290b5e4, 32'hc21a7269, 32'h424d66cf, 32'hc283526c};
test_weights[36680:36687] = '{32'hc1408dce, 32'h42418307, 32'hc18e457e, 32'hc257898f, 32'h42a4e61a, 32'h42322b9f, 32'h4181522e, 32'hc2402bc2};
test_bias[4585:4585] = '{32'h4182b23d};
test_output[4585:4585] = '{32'h467a5202};
test_input[36688:36695] = '{32'h429b5a6b, 32'h4238190a, 32'hc2a16576, 32'h41979f47, 32'hc1cc464f, 32'h4214a8fb, 32'hc260fb85, 32'h41e6bf80};
test_weights[36688:36695] = '{32'h418f11c7, 32'h423b8e9e, 32'h41de9244, 32'h421690e9, 32'hc2a89222, 32'hc0b31d0c, 32'hc220e0f8, 32'hc2a16176};
test_bias[4586:4586] = '{32'h41a1d82f};
test_output[4586:4586] = '{32'h4574aa36};
test_input[36696:36703] = '{32'h3eef767e, 32'hc216516d, 32'h4294194d, 32'hc2889499, 32'h4204dc38, 32'hc298d7f0, 32'h42887883, 32'h42b41f74};
test_weights[36696:36703] = '{32'hc29576d8, 32'hc2acd99f, 32'h4266966a, 32'h42aad2ec, 32'h425ebe66, 32'h41d0746c, 32'hc253a9a1, 32'hc2c35ef4};
test_bias[4587:4587] = '{32'hc215fa42};
test_output[4587:4587] = '{32'hc62aeb51};
test_input[36704:36711] = '{32'hc1acfd78, 32'hc0e29f42, 32'hc2bf95ec, 32'h42a19d2c, 32'h42a6c48d, 32'h427ed130, 32'hc28f4bed, 32'hc1f918b0};
test_weights[36704:36711] = '{32'h42ab75e4, 32'hc19f476e, 32'hc1a3e140, 32'hc2b7ab52, 32'hc09b3667, 32'h418a3a34, 32'hc2315653, 32'h4235b2a0};
test_bias[4588:4588] = '{32'h428c019f};
test_output[4588:4588] = '{32'hc5911816};
test_input[36712:36719] = '{32'hc259d97c, 32'h4091d448, 32'h418ab038, 32'hc28d792c, 32'h42af095f, 32'h4218a285, 32'h4279c5d3, 32'h403a3f94};
test_weights[36712:36719] = '{32'hc299a282, 32'hc1d373fb, 32'hc1154c6f, 32'hc28071a7, 32'h42260f23, 32'hc2bac5ae, 32'h410c2d19, 32'hc287df0a};
test_bias[4589:4589] = '{32'hc0c96fa7};
test_output[4589:4589] = '{32'h460a64ac};
test_input[36720:36727] = '{32'h42a8c7b6, 32'h42c6b06e, 32'h42850a2c, 32'hc27d8424, 32'h4261f4ba, 32'h421a36b6, 32'hc1e9eaf9, 32'h42637614};
test_weights[36720:36727] = '{32'h41824e5a, 32'hc1e22147, 32'hc28d4edc, 32'h42adc4bd, 32'hc1d164b7, 32'h420e1969, 32'h42a33823, 32'h4256f559};
test_bias[4590:4590] = '{32'h3fbe3aae};
test_output[4590:4590] = '{32'hc62d176e};
test_input[36728:36735] = '{32'hc26b42d0, 32'h428fbe96, 32'h429020a2, 32'h42035eea, 32'h41ccc162, 32'h42557211, 32'hc25e0063, 32'h428ac3b3};
test_weights[36728:36735] = '{32'hc23be657, 32'h41914cd3, 32'hc2aed5d9, 32'h40a7b27c, 32'h42667527, 32'h40d51c63, 32'hc2b080e5, 32'h42765d4d};
test_bias[4591:4591] = '{32'hc19b43bd};
test_output[4591:4591] = '{32'h460b6a64};
test_input[36736:36743] = '{32'h4103bce6, 32'hc24c34a5, 32'hc22fca5e, 32'hc1bd5b82, 32'h425bee82, 32'h4128b55d, 32'h41ebdfd3, 32'h42adb78f};
test_weights[36736:36743] = '{32'h423cf35a, 32'hc2a13ff2, 32'h41d19e0c, 32'h422bcc57, 32'h413e5434, 32'h4289a878, 32'hc1e9610e, 32'hc2bb5db8};
test_bias[4592:4592] = '{32'h41eeba21};
test_output[4592:4592] = '{32'hc5a4169a};
test_input[36744:36751] = '{32'hc2c2b402, 32'h42490adc, 32'h41887dde, 32'h42a0b5c9, 32'hc1dc9ee7, 32'h424a93c3, 32'h4220b8e9, 32'h4231ac27};
test_weights[36744:36751] = '{32'hc189bdad, 32'hc13d71ea, 32'hc23badf6, 32'h40a0778f, 32'hc24789b0, 32'hc176ab78, 32'hc2a73594, 32'h413694bc};
test_bias[4593:4593] = '{32'hc10b9038};
test_output[4593:4593] = '{32'hc4c5d771};
test_input[36752:36759] = '{32'h42996f93, 32'h414dba65, 32'hc27bc108, 32'h424f6563, 32'hc2c2ed3f, 32'hc2656572, 32'hc2a6d49e, 32'h4293c8e1};
test_weights[36752:36759] = '{32'h4206e6f4, 32'hc0514531, 32'hc27bc939, 32'hc238189f, 32'h42c328e2, 32'h40f58100, 32'hc2389899, 32'hc2b5d01a};
test_bias[4594:4594] = '{32'hc1dd32c4};
test_output[4594:4594] = '{32'hc6085454};
test_input[36760:36767] = '{32'hc16d72d2, 32'hc289c0e5, 32'hc0ed6532, 32'h42c6abd8, 32'hc2adf533, 32'hc092de97, 32'hc2bae544, 32'h41cb9a52};
test_weights[36760:36767] = '{32'h4223fb99, 32'hc26d9a6a, 32'h41bf703e, 32'hc2012b76, 32'hc271e369, 32'hc295f6cc, 32'hc2b3df90, 32'h40bbb232};
test_bias[4595:4595] = '{32'h428d7a31};
test_output[4595:4595] = '{32'h465fd7d3};
test_input[36768:36775] = '{32'h429c67f6, 32'h42bc5ea4, 32'h4207a623, 32'hc11ea6e7, 32'hc29f5c40, 32'hc1049d3e, 32'h4251d2da, 32'hc242344c};
test_weights[36768:36775] = '{32'hc1cb80ad, 32'h4214d2e7, 32'hc238ca62, 32'hc083a4da, 32'hc24301d2, 32'h42930e73, 32'h42b6bf72, 32'h421e767f};
test_bias[4596:4596] = '{32'h4218d8a6};
test_output[4596:4596] = '{32'h45c0e0c4};
test_input[36776:36783] = '{32'hc2971f8b, 32'h4299a296, 32'hc292e6d4, 32'h418dc244, 32'hc1f60695, 32'hc283fe62, 32'h42a1fbc8, 32'hc262620d};
test_weights[36776:36783] = '{32'h4208d464, 32'hc1d27210, 32'hc29a227b, 32'h428c18ac, 32'hc2904a20, 32'hc1dc7404, 32'h41536dd2, 32'h42a0fa8b};
test_bias[4597:4597] = '{32'h42bddca0};
test_output[4597:4597] = '{32'h4537f8f8};
test_input[36784:36791] = '{32'hc1a5b8df, 32'h3e3c238f, 32'h411d50d9, 32'h42a1e72e, 32'hc29c3030, 32'hc2898438, 32'h415cabc7, 32'hc21da0b5};
test_weights[36784:36791] = '{32'hc21b8a50, 32'hbfb72a2f, 32'hc1f25a55, 32'hc0545af0, 32'hc2bb339a, 32'h42bee45f, 32'h411a7b4e, 32'h3e303c44};
test_bias[4598:4598] = '{32'h420729d6};
test_output[4598:4598] = '{32'h448f3dd0};
test_input[36792:36799] = '{32'h4188616a, 32'hc0b29d2b, 32'hc2463319, 32'hc0a14285, 32'hc2019f82, 32'h429a4284, 32'hc28dfa5a, 32'h428f04bf};
test_weights[36792:36799] = '{32'hc24038cd, 32'hc22b82e5, 32'h427d4234, 32'h42a65c71, 32'h42bde00d, 32'hc267f1a4, 32'hc16ce289, 32'h4269fd21};
test_bias[4599:4599] = '{32'hc2accdb4};
test_output[4599:4599] = '{32'hc5cc4cb0};
test_input[36800:36807] = '{32'h415b3d2a, 32'h42afcfaf, 32'h4210ff3a, 32'hc28c9e1b, 32'h424ed6ed, 32'hc288ff4f, 32'h42a99049, 32'h428fac15};
test_weights[36800:36807] = '{32'h427dd9ef, 32'h42b96616, 32'h4234ae75, 32'hc0c9869b, 32'hc2852360, 32'h42b5e4bd, 32'hc299898f, 32'h4280c358};
test_bias[4600:4600] = '{32'hc29de8b2};
test_output[4600:4600] = '{32'hc406042a};
test_input[36808:36815] = '{32'h41ed914a, 32'hbfc10ce6, 32'h418dd906, 32'hc1ab1d39, 32'h426bd6bc, 32'hc243441b, 32'h41d0a0ad, 32'h422e140d};
test_weights[36808:36815] = '{32'h428bb833, 32'hc2bdee5f, 32'h42a0f270, 32'h41b0e293, 32'hbfb85612, 32'hc229b547, 32'h40a189fa, 32'h4259fe5d};
test_bias[4601:4601] = '{32'h41fae945};
test_output[4601:4601] = '{32'h45f065ae};
test_input[36816:36823] = '{32'h42b218f8, 32'h41babd7c, 32'h418c3efa, 32'hc2954120, 32'hc2c19c8b, 32'h426c45e9, 32'h4280b4dd, 32'h41b1fbd9};
test_weights[36816:36823] = '{32'h412d4e51, 32'h4272c0e6, 32'hc218db1d, 32'hbfbc2b9e, 32'h415c625a, 32'hc2891c9c, 32'hc2a2694b, 32'h429f1a43};
test_bias[4602:4602] = '{32'h41e5792d};
test_output[4602:4602] = '{32'hc5da69e9};
test_input[36824:36831] = '{32'hc2488156, 32'hc2908647, 32'h41a205e3, 32'hc1878c66, 32'h415a5a43, 32'h3f111866, 32'h4157a1ce, 32'h41ba07f3};
test_weights[36824:36831] = '{32'hc29c200f, 32'h4284a08d, 32'h418a7666, 32'h40222c72, 32'hc1b7a839, 32'h4292d3b5, 32'h3f3b7286, 32'hc28b8c7f};
test_bias[4603:4603] = '{32'hc284b31c};
test_output[4603:4603] = '{32'hc51da131};
test_input[36832:36839] = '{32'hc28494c8, 32'h42c1c6f5, 32'h421fc863, 32'hc200b67b, 32'h41c40b12, 32'hc183603f, 32'h420d4aa8, 32'hc241cbac};
test_weights[36832:36839] = '{32'hc1b84a70, 32'h41a2d9b7, 32'hbfdcbcf1, 32'hc2c4cbcd, 32'h42be709a, 32'h423f4aaa, 32'hc28e5e96, 32'h423556bf};
test_bias[4604:4604] = '{32'h42b9a7d4};
test_output[4604:4604] = '{32'h455c6c94};
test_input[36840:36847] = '{32'hbf018a99, 32'hc2236b97, 32'h416d1eec, 32'hc2babc84, 32'h42bb2fda, 32'h4241893c, 32'hc2b72f95, 32'h422aa8aa};
test_weights[36840:36847] = '{32'hbfcfe80a, 32'hc286d47c, 32'h40dc00cb, 32'h4014e917, 32'h42907bf5, 32'hc2336c25, 32'hc18c64a6, 32'h42ba3eb7};
test_bias[4605:4605] = '{32'h427dbb7a};
test_output[4605:4605] = '{32'h46492aa7};
test_input[36848:36855] = '{32'hc2c07503, 32'hc0bce161, 32'hc2bc842f, 32'h4217a324, 32'hc0bc3218, 32'hc00fba17, 32'h41b36a42, 32'h40832bae};
test_weights[36848:36855] = '{32'hc1c749d2, 32'h4263ef1b, 32'h42825ec3, 32'hc272ae57, 32'hc2a9ef25, 32'hc267d7e6, 32'h41911025, 32'hc232685f};
test_bias[4606:4606] = '{32'hc1ded8d1};
test_output[4606:4606] = '{32'hc5adac52};
test_input[36856:36863] = '{32'hc2754377, 32'h4220e3c1, 32'hc27ded87, 32'h41912c3b, 32'hc2af50d0, 32'h42932281, 32'hc2a7107a, 32'h4259d74e};
test_weights[36856:36863] = '{32'h42a5af86, 32'h4286d449, 32'h429d304a, 32'hc260abc8, 32'h4244d605, 32'h4173ef6e, 32'hc1abd654, 32'h4260300a};
test_bias[4607:4607] = '{32'h423a28b0};
test_output[4607:4607] = '{32'hc5d09b50};
test_input[36864:36871] = '{32'h428d003d, 32'hc2b3db04, 32'h4230d717, 32'hc201d9b7, 32'h4258eeac, 32'hc2a432f7, 32'h41a90b25, 32'h40494e5d};
test_weights[36864:36871] = '{32'hbe404cdc, 32'h409af9c1, 32'h3e3262dd, 32'hc262c171, 32'h42842668, 32'hc22e4e86, 32'h425b038b, 32'hc1dee9a8};
test_bias[4608:4608] = '{32'hc299efa5};
test_output[4608:4608] = '{32'h46154292};
test_input[36872:36879] = '{32'hc214e298, 32'h42c2a655, 32'h41632790, 32'hc1b4ff8a, 32'h4235a663, 32'hc22cd2b0, 32'hbfd04547, 32'h41b3f45a};
test_weights[36872:36879] = '{32'hc18f93e9, 32'h41c98e7d, 32'hc2bce70f, 32'h4192fb7e, 32'hc24ad4f1, 32'hc1de61af, 32'hc2826c80, 32'hc2b64a87};
test_bias[4609:4609] = '{32'h4148c78c};
test_output[4609:4609] = '{32'hc4d0bcba};
test_input[36880:36887] = '{32'hc205f776, 32'h413dff78, 32'h424baf97, 32'hc20557d2, 32'hc1e359ce, 32'h42ab879a, 32'hc1948d68, 32'h42b81501};
test_weights[36880:36887] = '{32'h41a61525, 32'h42a5672c, 32'hc28e4b10, 32'hc1a97f28, 32'h425b0162, 32'hc0faa687, 32'h4170adcf, 32'hc2bab912};
test_bias[4610:4610] = '{32'h4275fa5c};
test_output[4610:4610] = '{32'hc65591fc};
test_input[36888:36895] = '{32'h426e6f97, 32'hc2a47205, 32'h41ceb64b, 32'h40e63e7e, 32'h42a436a3, 32'h425472a3, 32'h41d1fc57, 32'h421f125b};
test_weights[36888:36895] = '{32'hc15b6abc, 32'hc1a0e37e, 32'hc213dad2, 32'h428ce11c, 32'hc1fb8d64, 32'h42201e8a, 32'hc27432f6, 32'h419a556a};
test_bias[4611:4611] = '{32'hc20592be};
test_output[4611:4611] = '{32'hc46a200d};
test_input[36896:36903] = '{32'hc1b3e9fc, 32'h411fa74d, 32'hc2c5b85f, 32'h426d7012, 32'h41826fad, 32'hc2c35372, 32'hc283eaac, 32'hbfc9c496};
test_weights[36896:36903] = '{32'h422907f7, 32'h422cade7, 32'hc1ed30a3, 32'hc214a569, 32'hc1828e7f, 32'hc2a6f18f, 32'h420065ef, 32'h424162a3};
test_bias[4612:4612] = '{32'h413ee558};
test_output[4612:4612] = '{32'h45b8b0f3};
test_input[36904:36911] = '{32'hc2156272, 32'hc0cb1ee4, 32'h42b30eec, 32'h429ef7d1, 32'hc211df74, 32'hc2acb1f9, 32'hc29a9afb, 32'hc218c4b5};
test_weights[36904:36911] = '{32'hc098d199, 32'h42a5c570, 32'hc2c1295a, 32'h42acd620, 32'h4278ee5a, 32'h4294db72, 32'hc21cafe9, 32'h426d5e0d};
test_bias[4613:4613] = '{32'h42805a21};
test_output[4613:4613] = '{32'hc61c304a};
test_input[36912:36919] = '{32'hc16464e0, 32'hc1e2d3b8, 32'h42480890, 32'h4130aa1a, 32'hc2ba39e5, 32'h419192c9, 32'hc20691ac, 32'h41cd672d};
test_weights[36912:36919] = '{32'hc1a3beb6, 32'hc23e01b0, 32'hc286084a, 32'h41523a69, 32'hc17479e7, 32'hc28c52d4, 32'h42b996f3, 32'h421027c9};
test_bias[4614:4614] = '{32'hc1bec715};
test_output[4614:4614] = '{32'hc56399d3};
test_input[36920:36927] = '{32'h42374d91, 32'h4256af7c, 32'hc188e2c8, 32'hc240b382, 32'h42848eb0, 32'hc2badee1, 32'hc094ced4, 32'h428229f4};
test_weights[36920:36927] = '{32'h42a77cf1, 32'hc29ab0dd, 32'h4218867d, 32'h4280ffaf, 32'hc1df617d, 32'hc294db4f, 32'hc2aa4e94, 32'hc205643e};
test_bias[4615:4615] = '{32'h42b4dccb};
test_output[4615:4615] = '{32'hc4236d0a};
test_input[36928:36935] = '{32'h4274b13b, 32'hc213e310, 32'h4238f7c9, 32'h412c688d, 32'h4217b819, 32'hc2023453, 32'hc065aee7, 32'h42b8ced0};
test_weights[36928:36935] = '{32'h42519c34, 32'hc2ab6151, 32'hc1e3c444, 32'h41fd23ac, 32'h42bb0165, 32'hc2a45260, 32'h423114e1, 32'h4109dc52};
test_bias[4616:4616] = '{32'hc1a67332};
test_output[4616:4616] = '{32'h463f2e73};
test_input[36936:36943] = '{32'hc1fcd459, 32'hc2a122f3, 32'hc1828326, 32'h4251339f, 32'h41b6ef5e, 32'h4235a25a, 32'h42174dfd, 32'hc27caee0};
test_weights[36936:36943] = '{32'h42a5ecb7, 32'hc205358b, 32'h42196a31, 32'hc294039f, 32'h4277d614, 32'h42ac0b4c, 32'hc29aa4a3, 32'hc18273af};
test_bias[4617:4617] = '{32'h42b7f7c9};
test_output[4617:4617] = '{32'hc464b763};
test_input[36944:36951] = '{32'hc28f60d5, 32'h41cb5d5e, 32'hc234e049, 32'h424d7fec, 32'hc233c564, 32'hc21e0cb9, 32'hc23fa7be, 32'h428dabcb};
test_weights[36944:36951] = '{32'h41d97c1d, 32'hc1b573e4, 32'h42bf72ba, 32'h41eb87e2, 32'h3fe6a67e, 32'hc20f69b6, 32'h403c9491, 32'h41d7c141};
test_bias[4618:4618] = '{32'hc107a58d};
test_output[4618:4618] = '{32'hc50c519d};
test_input[36952:36959] = '{32'h41263e93, 32'hc1a5c3d5, 32'h42a3e37e, 32'h422742eb, 32'h4123a436, 32'hc23f4f46, 32'h42852a63, 32'hc266b99a};
test_weights[36952:36959] = '{32'h429981b7, 32'h42a4b4f6, 32'hc2648d2e, 32'h42955b9a, 32'h429e981c, 32'h429696a0, 32'h422e9faf, 32'hc29f5a2a};
test_bias[4619:4619] = '{32'h4264c4ab};
test_output[4619:4619] = '{32'h450fd4f6};
test_input[36960:36967] = '{32'h3fcc2c7e, 32'hc2481f48, 32'hc2b7a052, 32'hc29ecc68, 32'h42685799, 32'h429afe5e, 32'hc2c6b06b, 32'h41389c47};
test_weights[36960:36967] = '{32'h42abb729, 32'hc28113a8, 32'h42bc9d08, 32'h42bb8eba, 32'hc2c331fd, 32'hc2ab6421, 32'hc2c41127, 32'h411fb632};
test_bias[4620:4620] = '{32'h429306a3};
test_output[4620:4620] = '{32'hc66c444c};
test_input[36968:36975] = '{32'hc194731a, 32'hc1cf8633, 32'h428c010d, 32'hc0201d0b, 32'h4236ad86, 32'hc2c293a4, 32'h4195f15f, 32'hc192b5f8};
test_weights[36968:36975] = '{32'hc2af243a, 32'h42a0210b, 32'hc2965f76, 32'h4287669c, 32'hc29078a8, 32'h422bd885, 32'h425c9f3d, 32'h42c54af7};
test_bias[4621:4621] = '{32'hc299a121};
test_output[4621:4621] = '{32'hc65e1cea};
test_input[36976:36983] = '{32'h420e5649, 32'h427e1792, 32'h42b0b306, 32'h414a4077, 32'hc0dec441, 32'hc1c68c11, 32'h4254ec70, 32'h40b7d111};
test_weights[36976:36983] = '{32'hc26d04e6, 32'hc1284e15, 32'hc29bc7bb, 32'hc1a5c502, 32'hc285089b, 32'h40de6a1c, 32'h41cf9df5, 32'h41ad9709};
test_bias[4622:4622] = '{32'h41c92797};
test_output[4622:4622] = '{32'hc5fd1380};
test_input[36984:36991] = '{32'hc13f03b7, 32'h4202ef25, 32'h41caf0a0, 32'hc0ecb40c, 32'hc215adbe, 32'h41fe1959, 32'hc27ccb38, 32'h4202dc23};
test_weights[36984:36991] = '{32'h41254cd9, 32'h4129740f, 32'hc1e92f76, 32'hc1b9711a, 32'hc270e9bc, 32'h40b3c7c1, 32'hc195d98d, 32'h423a16a4};
test_bias[4623:4623] = '{32'h42554812};
test_output[4623:4623] = '{32'h45977502};
test_input[36992:36999] = '{32'h41c7a13b, 32'h42c7eec7, 32'hc0ccbcdc, 32'hc1a19dee, 32'h42053135, 32'h428ea051, 32'h4236e977, 32'hc22ff475};
test_weights[36992:36999] = '{32'hc22d3cbc, 32'h428c0602, 32'hc2960d13, 32'hc2ad5887, 32'hc238429e, 32'h42c0f16d, 32'hc2aa5b78, 32'hc1fe0523};
test_bias[4624:4624] = '{32'h4121f625};
test_output[4624:4624] = '{32'h462bfae0};
test_input[37000:37007] = '{32'hc2567c46, 32'h4286a1c7, 32'hc289de73, 32'h42a8b48a, 32'h4245d0b3, 32'h4126a558, 32'h42203bf0, 32'hc224b34e};
test_weights[37000:37007] = '{32'hc2368227, 32'h428e67f4, 32'hc1438bc9, 32'h42c1bbcf, 32'hc21ec091, 32'hc2457dcd, 32'hc243a32f, 32'hc27c952d};
test_bias[4625:4625] = '{32'hc10adc96};
test_output[4625:4625] = '{32'h46612135};
test_input[37008:37015] = '{32'hc233f451, 32'h421a1114, 32'hc2a6c048, 32'hc2b22929, 32'h426ef803, 32'h42c21d58, 32'h42c20d9e, 32'h42ab40f5};
test_weights[37008:37015] = '{32'hc23443ab, 32'hc16e1834, 32'hc29cb975, 32'hc282de0d, 32'h429fd422, 32'hc0b26ccd, 32'h4247322a, 32'hc2b74184};
test_bias[4626:4626] = '{32'hc1bf7f86};
test_output[4626:4626] = '{32'h466a8f3c};
test_input[37016:37023] = '{32'hc2bd2d9d, 32'hc283c23a, 32'h42092be3, 32'h41fe7a26, 32'hc18fb92e, 32'hc2a668a3, 32'hc2385307, 32'hc15722bd};
test_weights[37016:37023] = '{32'h42b2b5a3, 32'hc2023741, 32'hc28951ca, 32'hc2950f37, 32'h4252d835, 32'hc27e4251, 32'h41164e82, 32'hc25c07cb};
test_bias[4627:4627] = '{32'hc25165d8};
test_output[4627:4627] = '{32'hc5c92303};
test_input[37024:37031] = '{32'hc299c8d4, 32'hc2a5fca2, 32'h428d3ec7, 32'hc1891115, 32'h428a5fe8, 32'h4217e0c8, 32'h4270c6eb, 32'h4251a28a};
test_weights[37024:37031] = '{32'hc0ce307c, 32'h429b2df7, 32'hc28c06d1, 32'h428cd781, 32'hc2a40efa, 32'h421e4233, 32'hc2c1918f, 32'h42698ffb};
test_bias[4628:4628] = '{32'h40f2f0da};
test_output[4628:4628] = '{32'hc694a491};
test_input[37032:37039] = '{32'hc20b16c8, 32'hc203dde4, 32'h427c705d, 32'h404f022e, 32'h42b44d71, 32'h427a3bf3, 32'hc29358d1, 32'hc0a6bbe5};
test_weights[37032:37039] = '{32'hc2007810, 32'h428649c5, 32'h42a5e165, 32'hc1a786bd, 32'h410ff393, 32'h423b7b87, 32'hc15cfba1, 32'h4097f281};
test_bias[4629:4629] = '{32'hc26fddbd};
test_output[4629:4629] = '{32'h4608a7cb};
test_input[37040:37047] = '{32'h42a8124d, 32'h42767c0e, 32'h415c5e48, 32'h42b38e09, 32'h3e9527c1, 32'hc2a1d3d2, 32'h42a8f1ab, 32'h4252c442};
test_weights[37040:37047] = '{32'h403e7f91, 32'hc27b17ca, 32'hc1e51848, 32'hc24b79ee, 32'hc232bd6d, 32'hc2530926, 32'hc286a684, 32'h4260fb1e};
test_bias[4630:4630] = '{32'h429cbca9};
test_output[4630:4630] = '{32'hc5d9c407};
test_input[37048:37055] = '{32'hc2b47e11, 32'h429881bc, 32'hc1de7dcb, 32'h42100516, 32'hc1ad0d70, 32'hc21cff0c, 32'hc2a5c963, 32'hc2157631};
test_weights[37048:37055] = '{32'h42297b72, 32'hc2543402, 32'hc28e14e2, 32'h4055ceca, 32'h4290362b, 32'h415b38a9, 32'h42655e81, 32'h4277c3e1};
test_bias[4631:4631] = '{32'hc2202904};
test_output[4631:4631] = '{32'hc66a0983};
test_input[37056:37063] = '{32'h42b8ceb2, 32'hc18e1c6f, 32'hc2a2d63e, 32'hc282369d, 32'h40ff0ebd, 32'hc180f62d, 32'hc2af780a, 32'hc2588296};
test_weights[37056:37063] = '{32'hc143d5f6, 32'h408d8e88, 32'hc118d53b, 32'h422dbd2f, 32'h417a8136, 32'h42718232, 32'h41dc6f0c, 32'h42b56fad};
test_bias[4632:4632] = '{32'hc2b67a0b};
test_output[4632:4632] = '{32'hc6341d30};
test_input[37064:37071] = '{32'h42969e87, 32'hc2a7e017, 32'hc216ee94, 32'hc2a1e18c, 32'h41c1ffac, 32'h42b30312, 32'h4297a30c, 32'h428b6d46};
test_weights[37064:37071] = '{32'h428e9726, 32'hc1861ff7, 32'h42baaa37, 32'h42623026, 32'h4238c1b4, 32'hc1b2c9d3, 32'h42197ee2, 32'h4225ef24};
test_bias[4633:4633] = '{32'hc22d024f};
test_output[4633:4633] = '{32'h455e3bb7};
test_input[37072:37079] = '{32'h42c37e74, 32'h422e05c3, 32'hc217e37c, 32'h41b4de4f, 32'hc288b044, 32'h41ce6822, 32'h4275c2da, 32'h4253a6c0};
test_weights[37072:37079] = '{32'hc2a343c3, 32'hc24e447b, 32'h41bed432, 32'hc27bb3a9, 32'h42afc14e, 32'h3f15b852, 32'hc1e9c1bd, 32'hc19ebd91};
test_bias[4634:4634] = '{32'hc1b4fa50};
test_output[4634:4634] = '{32'hc6a743ac};
test_input[37080:37087] = '{32'h424d1d6e, 32'h417d98df, 32'h42409c9a, 32'h42797147, 32'h427b1dd8, 32'hc28cfcaa, 32'hc2b5c24a, 32'hc158a726};
test_weights[37080:37087] = '{32'h42b125b9, 32'hc2bbd483, 32'hc28dbe1c, 32'hc1be04bd, 32'h413f2722, 32'h42072dbc, 32'hc1e0b9a9, 32'h429d1159};
test_bias[4635:4635] = '{32'h42a3cba0};
test_output[4635:4635] = '{32'hc4edac6f};
test_input[37088:37095] = '{32'h421c52b2, 32'hc1ce8de1, 32'h42845d3a, 32'hc182e8b7, 32'h4251ae24, 32'h422e3709, 32'hc2a3cbe1, 32'hc2b5e13e};
test_weights[37088:37095] = '{32'h42a2fea9, 32'hc21b2f89, 32'hc1d1e38c, 32'h428208e6, 32'hc23f0ba8, 32'hc2956256, 32'h42415dde, 32'h42acf016};
test_bias[4636:4636] = '{32'h42630e21};
test_output[4636:4636] = '{32'hc67c20c1};
test_input[37096:37103] = '{32'h418db3de, 32'hc296c9a4, 32'hc2ab5e3f, 32'hc2870395, 32'h42594322, 32'h4298e31c, 32'h42705718, 32'h4281a807};
test_weights[37096:37103] = '{32'h429f96b7, 32'h42a13881, 32'hc2bdfa8b, 32'h4246a896, 32'hc299cc5d, 32'hc0a83c00, 32'hc289433b, 32'hc28c0120};
test_bias[4637:4637] = '{32'hc2b54946};
test_output[4637:4637] = '{32'hc64e63d6};
test_input[37104:37111] = '{32'hc1e31175, 32'hc2a28926, 32'hc172bbc8, 32'hc01569cd, 32'hc26faf76, 32'hc2b930ee, 32'hc1ff906b, 32'hc18b6086};
test_weights[37104:37111] = '{32'hc289b1da, 32'hc1d66c08, 32'hc2a1c561, 32'h42a570ab, 32'hc28fa9cd, 32'hc29d606a, 32'h417a0fbc, 32'h42200a1e};
test_bias[4638:4638] = '{32'h408ecee3};
test_output[4638:4638] = '{32'h4673338e};
test_input[37112:37119] = '{32'hc20ff3df, 32'hbf964197, 32'hc17739b9, 32'hc2ba8b3f, 32'h416e754b, 32'hc2903002, 32'hc275f802, 32'hc0d569dd};
test_weights[37112:37119] = '{32'h4292cb82, 32'hc1ab2016, 32'h423ecf3e, 32'hc2b3ddda, 32'h40cf513a, 32'h41fdd84a, 32'h42b1fa70, 32'hc12bc4ee};
test_bias[4639:4639] = '{32'h42056bc5};
test_output[4639:4639] = '{32'hc51db5bf};
test_input[37120:37127] = '{32'hc1288f04, 32'hc10da618, 32'hc2992fb8, 32'h41126686, 32'hc2b298e7, 32'hc101cce8, 32'h42bc5f53, 32'h40edf73d};
test_weights[37120:37127] = '{32'hc219d212, 32'hc1b227a9, 32'hc2287a50, 32'hc12fcb78, 32'h40defa3c, 32'h424b3efb, 32'h429658e5, 32'hc270cae1};
test_bias[4640:4640] = '{32'hc1d478c2};
test_output[4640:4640] = '{32'h46114dd2};
test_input[37128:37135] = '{32'hc2b8f68f, 32'hc205482f, 32'h424a81f5, 32'h42ad3ef0, 32'h422328f4, 32'hc2b64b92, 32'hc2852500, 32'hc1497c4e};
test_weights[37128:37135] = '{32'h426978e1, 32'h4141d022, 32'hc2413337, 32'hc1aa3303, 32'h428be87a, 32'h42a906e0, 32'h4239c977, 32'hc23db498};
test_bias[4641:4641] = '{32'hc25d4c4f};
test_output[4641:4641] = '{32'hc688a362};
test_input[37136:37143] = '{32'hc236e8be, 32'hc294ac41, 32'h427b024d, 32'h42aa1baf, 32'h421c6509, 32'hc28c0026, 32'hc2b79603, 32'h4282f3b3};
test_weights[37136:37143] = '{32'h4225350b, 32'h42b78d4b, 32'h425baf85, 32'h42609767, 32'h4227af42, 32'hc23b538c, 32'h421dbcec, 32'h4186932e};
test_bias[4642:4642] = '{32'hc23aaba8};
test_output[4642:4642] = '{32'h44e8eba4};
test_input[37144:37151] = '{32'h42bfd89b, 32'h41ce2992, 32'h41bdeb61, 32'hc180307f, 32'h4125ec7c, 32'h42aa12a5, 32'h419dc664, 32'h426b8b97};
test_weights[37144:37151] = '{32'hc24a84a5, 32'h429fa2ad, 32'hc2b377f3, 32'h416cace1, 32'h4211b815, 32'h428930c6, 32'h420406d1, 32'h428361be};
test_bias[4643:4643] = '{32'h423e2657};
test_output[4643:4643] = '{32'h45af55ef};
test_input[37152:37159] = '{32'h41bbc387, 32'h419b335c, 32'h42081f92, 32'h4272cda7, 32'hc29393bd, 32'hc200a617, 32'hc09b5583, 32'hc1988604};
test_weights[37152:37159] = '{32'hc2af6d63, 32'h40d63bcf, 32'h42297f63, 32'h400f07f6, 32'hbf531c7f, 32'h41d1ddad, 32'h42a4528e, 32'h42118987};
test_bias[4644:4644] = '{32'h405e9e06};
test_output[4644:4644] = '{32'hc50af019};
test_input[37160:37167] = '{32'h421d289d, 32'hc28f6394, 32'h429030db, 32'h41fa0fea, 32'hc1f7a2b6, 32'h4224c0bb, 32'h4199a3a8, 32'hc28cb6df};
test_weights[37160:37167] = '{32'hc01dd550, 32'hc27297c8, 32'h427e0770, 32'hc25e0333, 32'h4284f06e, 32'hc0d694f8, 32'hc259388b, 32'h42b5d0e5};
test_bias[4645:4645] = '{32'hc2bbe152};
test_output[4645:4645] = '{32'hc52d3b15};
test_input[37168:37175] = '{32'hc20e0b6b, 32'h422a04ca, 32'h410455ae, 32'h3fd2773b, 32'hc2b9b184, 32'hc253548e, 32'h429aa11d, 32'hc2bef903};
test_weights[37168:37175] = '{32'hc06d209a, 32'h41d675c7, 32'h41b1ab41, 32'h4278df02, 32'h4196683a, 32'h4145e9b4, 32'hbfecf9c2, 32'h4280ae89};
test_bias[4646:4646] = '{32'h40ca941e};
test_output[4646:4646] = '{32'hc5de94c3};
test_input[37176:37183] = '{32'hc2ba5f63, 32'h40518ac5, 32'hc2b10801, 32'hc2b7da3d, 32'h41b776b1, 32'hc25f344c, 32'hc09922d1, 32'h42a284ef};
test_weights[37176:37183] = '{32'hc1f1615f, 32'h4291ab69, 32'hc2908efb, 32'h42a72008, 32'hc2a6db5c, 32'h412e5435, 32'h42b4156f, 32'hc217dbde};
test_bias[4647:4647] = '{32'hc23ba399};
test_output[4647:4647] = '{32'hc586ed4a};
test_input[37184:37191] = '{32'h420a722c, 32'h42307f95, 32'hc291116d, 32'h42abbc56, 32'hc295dd81, 32'hc204c8d1, 32'hc042bd90, 32'h42a2f671};
test_weights[37184:37191] = '{32'hc2152485, 32'h42a53016, 32'hc2c76f45, 32'hc21170b3, 32'hc2a80da2, 32'h4202fa15, 32'hc21e13da, 32'h41874a1d};
test_bias[4648:4648] = '{32'hc189ca92};
test_output[4648:4648] = '{32'h464d8bea};
test_input[37192:37199] = '{32'h42808f60, 32'hc2b5791b, 32'hc2867008, 32'h41e2a34c, 32'h42415534, 32'hc221d127, 32'h42141485, 32'hc29f08aa};
test_weights[37192:37199] = '{32'h42a2dc47, 32'hc113ae68, 32'h4243bed9, 32'hc22ee167, 32'h424d6a68, 32'hc2257f84, 32'h42551b92, 32'h4224a322};
test_bias[4649:4649] = '{32'hc088851a};
test_output[4649:4649] = '{32'h45895709};
test_input[37200:37207] = '{32'hc1a51495, 32'h42a151fb, 32'h415b8ba2, 32'hc2c125a9, 32'h41fbd197, 32'h41b84b10, 32'hc24b887d, 32'h42adf147};
test_weights[37200:37207] = '{32'hc284ef80, 32'hc2c7861b, 32'hc2583557, 32'h42873d48, 32'hc28f0a90, 32'hc21c3892, 32'hc15c7be9, 32'hc016e6b4};
test_bias[4650:4650] = '{32'hc2b320fa};
test_output[4650:4650] = '{32'hc682673e};
test_input[37208:37215] = '{32'h42a4a09f, 32'h41b47d51, 32'hc26b5f59, 32'h4283923a, 32'hc2be4fa5, 32'h42432709, 32'h42a9aeea, 32'hc2412bdd};
test_weights[37208:37215] = '{32'hc1721d08, 32'hc274c3d4, 32'h424a4a9c, 32'hc241ef5f, 32'hc0fa245d, 32'hc28cb067, 32'hc21dd503, 32'h4283af31};
test_bias[4651:4651] = '{32'h4286cf5b};
test_output[4651:4651] = '{32'hc68c2751};
test_input[37216:37223] = '{32'hc2aa47a5, 32'hc240d9a1, 32'h420c271a, 32'hc215ff58, 32'h420191d2, 32'hc1e18026, 32'hc2966464, 32'hc2a579f5};
test_weights[37216:37223] = '{32'h428b646b, 32'h42ae65ad, 32'h4271b145, 32'hc1f7517b, 32'h42aaa536, 32'hc28b3360, 32'hc2b73a6b, 32'h429665e0};
test_bias[4652:4652] = '{32'h427dd1cb};
test_output[4652:4652] = '{32'hc4afa88f};
test_input[37224:37231] = '{32'h42b64702, 32'hc2b8dad7, 32'hc2af3b50, 32'hc285074c, 32'hc290d484, 32'h41d3acda, 32'hc28e160d, 32'h42691ef7};
test_weights[37224:37231] = '{32'hc1025812, 32'hc2876760, 32'hc2a5787c, 32'hc1a47155, 32'hc20f7a57, 32'hc2ba8a5d, 32'hc2c32cdb, 32'hc2b62ddf};
test_bias[4653:4653] = '{32'hc1b93117};
test_output[4653:4653] = '{32'h4677d776};
test_input[37232:37239] = '{32'h41d07cd4, 32'h4276b617, 32'h42a1e2d0, 32'hc2a14740, 32'h410d9a31, 32'hc2a9a696, 32'hc11b8db6, 32'hc2529d73};
test_weights[37232:37239] = '{32'h4276127c, 32'h42395f33, 32'h42c54044, 32'hc24d60a6, 32'h41c0d617, 32'h425cf141, 32'hc1b4efd0, 32'h42a605ae};
test_bias[4654:4654] = '{32'hc1e1ee1b};
test_output[4654:4654] = '{32'h45f7edb3};
test_input[37240:37247] = '{32'h41f19223, 32'hc29acfb0, 32'hc2203f91, 32'hc2b9e908, 32'hc0e79f70, 32'h3d2ad7b2, 32'hc225807b, 32'h42924c2f};
test_weights[37240:37247] = '{32'hc2189ea5, 32'h425e91bb, 32'hc001dc26, 32'h42b0d54e, 32'hc20f4c22, 32'hc25415c7, 32'h41ab0a2a, 32'hc24d067a};
test_bias[4655:4655] = '{32'hc29bae7c};
test_output[4655:4655] = '{32'hc68d06b4};
test_input[37248:37255] = '{32'hc297b294, 32'h429fb306, 32'h41a761e4, 32'h4048f2c7, 32'hc1c5f2ce, 32'h4244cc70, 32'hc2480682, 32'h4284ac48};
test_weights[37248:37255] = '{32'h42abff71, 32'hc1599227, 32'h427dc6ea, 32'hc244cfe0, 32'h42780da9, 32'h422bf029, 32'hc25aef30, 32'h4086dac0};
test_bias[4656:4656] = '{32'hc2a187e1};
test_output[4656:4656] = '{32'hc536791f};
test_input[37256:37263] = '{32'h408ce2b1, 32'hc01405c8, 32'h4289bda0, 32'hc0d89663, 32'hc1a722a3, 32'hc285b70c, 32'hc1b3fb90, 32'hc21006a3};
test_weights[37256:37263] = '{32'h41946c71, 32'hc24eb897, 32'hc15b3f30, 32'hc286922f, 32'h427373fd, 32'hc2448363, 32'hc1b7a3a7, 32'hc0f1d803};
test_bias[4657:4657] = '{32'h426707c2};
test_output[4657:4657] = '{32'h4520c42d};
test_input[37264:37271] = '{32'h4098ce65, 32'hc29025ab, 32'h42aafd5d, 32'h42b29573, 32'h42983285, 32'hc1dff6c3, 32'h42a8d094, 32'hc2a62835};
test_weights[37264:37271] = '{32'hc28039ad, 32'h42b48f24, 32'h42bc2cf6, 32'h41bcb301, 32'hc2186979, 32'hc24997a2, 32'hc1d7b47d, 32'hc194a8aa};
test_bias[4658:4658] = '{32'hc28f4018};
test_output[4658:4658] = '{32'h44829c27};
test_input[37272:37279] = '{32'hc2c37835, 32'h4000ba8e, 32'h42748a63, 32'h42b58ee0, 32'h418d3df8, 32'h42c70c0a, 32'h42bd16da, 32'h42bc7884};
test_weights[37272:37279] = '{32'hc2a70c12, 32'hc2500fac, 32'h418462b0, 32'hc206ec4a, 32'hc28355d6, 32'hc18ab9b7, 32'hc18059e9, 32'hc2c4c022};
test_bias[4659:4659] = '{32'h409fb75e};
test_output[4659:4659] = '{32'hc5ef5a96};
test_input[37280:37287] = '{32'h40fb92fa, 32'h42932506, 32'h4185eb2c, 32'h423f2197, 32'h42ab537e, 32'hc277c8b5, 32'hc22261dd, 32'hbf83e7ab};
test_weights[37280:37287] = '{32'h41d90773, 32'h41c87c84, 32'h420a2320, 32'hc2216f70, 32'h42b1e360, 32'hc2ad6425, 32'hc29ecd53, 32'h423b8e5a};
test_bias[4660:4660] = '{32'h41aa9807};
test_output[4660:4660] = '{32'h4683f968};
test_input[37288:37295] = '{32'h3ff4a838, 32'h429eed0c, 32'hc28001f4, 32'hc21a175f, 32'hc239b0a1, 32'hc2c653d4, 32'hc1f8266c, 32'hc25387ee};
test_weights[37288:37295] = '{32'hc0e0ea10, 32'h40b3d2dc, 32'hc277aa65, 32'hc1b88703, 32'hc1a17695, 32'h4262e731, 32'hc26556cb, 32'hc20fdfe9};
test_bias[4661:4661] = '{32'hc2705a3c};
test_output[4661:4661] = '{32'h4583c6c4};
test_input[37296:37303] = '{32'hc12a165e, 32'h4220040e, 32'hc1c94f1d, 32'hc2c65275, 32'hc29e26ac, 32'hc269b669, 32'h42438252, 32'h42993244};
test_weights[37296:37303] = '{32'h420b6325, 32'hc0debd86, 32'hc1cbdf49, 32'hc27cd3b1, 32'hc29e7335, 32'h4089f15b, 32'hc26be791, 32'hc2b79c5e};
test_bias[4662:4662] = '{32'h42bf2abd};
test_output[4662:4662] = '{32'h45195c85};
test_input[37304:37311] = '{32'hc1b38ae3, 32'h42748198, 32'hc2674d0c, 32'hc2a43648, 32'hc23a9b2c, 32'hc20328af, 32'h4240e5f1, 32'hc27d320f};
test_weights[37304:37311] = '{32'hc2af41aa, 32'hc29eff5a, 32'h408a26c2, 32'hc19be9c0, 32'hc287b33a, 32'hc29d345d, 32'hc282597a, 32'h4283a3f5};
test_bias[4663:4663] = '{32'h3f1a9d0e};
test_output[4663:4663] = '{32'hc5424708};
test_input[37312:37319] = '{32'h4239187f, 32'h41850779, 32'hc1e77c8c, 32'h4296cb10, 32'hc273e85b, 32'h42a324ab, 32'hc17472a2, 32'hc27530d0};
test_weights[37312:37319] = '{32'h42c0f001, 32'h41f64512, 32'hc0d936c4, 32'hc1ac4a66, 32'h41aee263, 32'h41b9e030, 32'hc1f03774, 32'hc1e1ed53};
test_bias[4664:4664] = '{32'h3f1a88fc};
test_output[4664:4664] = '{32'h45c4ea29};
test_input[37320:37327] = '{32'h423b8794, 32'h42c3f408, 32'h42359548, 32'h41d03ca6, 32'hc1db4f58, 32'hc235e572, 32'h42a5f54c, 32'hc19053d4};
test_weights[37320:37327] = '{32'h41dca8fb, 32'h42647aff, 32'hbf1b0513, 32'h41f07d95, 32'hc2c091c1, 32'hc2833efd, 32'h425c0c79, 32'h42b4d68c};
test_bias[4665:4665] = '{32'h42083482};
test_output[4665:4665] = '{32'h467daf9d};
test_input[37328:37335] = '{32'hc19c2786, 32'h425a9a45, 32'hc245f1c8, 32'hc1ecbf26, 32'h42a762d9, 32'h42af7757, 32'hc15493a2, 32'h41da85e2};
test_weights[37328:37335] = '{32'h42bb1a01, 32'hc200672c, 32'h424fbb52, 32'h41f4aafd, 32'h420d8d27, 32'h424cb353, 32'h42872bcb, 32'hc28d65bb};
test_bias[4666:4666] = '{32'h41c2be63};
test_output[4666:4666] = '{32'hc5168b19};
test_input[37336:37343] = '{32'h41aee322, 32'hc0d89ddf, 32'h429e147b, 32'hc029cb4f, 32'hc1ccadc7, 32'h42948eb3, 32'hc1d92b7f, 32'hc2bb0a54};
test_weights[37336:37343] = '{32'hc2a6f765, 32'hc2b0b416, 32'h428d1254, 32'h4165fb8b, 32'h42034643, 32'hc2764e92, 32'h428b1314, 32'h41a41b4f};
test_bias[4667:4667] = '{32'h41d3dcbc};
test_output[4667:4667] = '{32'hc598983a};
test_input[37344:37351] = '{32'h41fae6ed, 32'hc259b39f, 32'hc2c3b2c4, 32'hc2b6cd7d, 32'hc25c704a, 32'h412eb695, 32'h419fe078, 32'hc0eb0696};
test_weights[37344:37351] = '{32'hc29d096e, 32'h42a18080, 32'h4064a581, 32'hc1dab528, 32'hc12cb347, 32'h415714e4, 32'h429e0dac, 32'hc2953d5b};
test_bias[4668:4668] = '{32'hc24c17d0};
test_output[4668:4668] = '{32'hc4ec4958};
test_input[37352:37359] = '{32'hc104cac6, 32'hc1d8dd1f, 32'h42b1015d, 32'h41f7c099, 32'hc2628b94, 32'h405a9700, 32'h42835d89, 32'hc18589e1};
test_weights[37352:37359] = '{32'h41e5ce10, 32'hc12101ed, 32'hc2c45990, 32'hc2902510, 32'hc1a0df0c, 32'h41a8a741, 32'h42a8ef73, 32'h414a17d3};
test_bias[4669:4669] = '{32'hc23e38b4};
test_output[4669:4669] = '{32'hc5890e76};
test_input[37360:37367] = '{32'h42b1d82c, 32'hc2b8b827, 32'hc23f5c08, 32'h40e49831, 32'hc128ee65, 32'h42985f01, 32'hc0473410, 32'hc2281f43};
test_weights[37360:37367] = '{32'h42949ffd, 32'hc2306e7b, 32'hc24a58e3, 32'h42472cba, 32'hc0f2656d, 32'h42bd3b10, 32'hc2868e6d, 32'h429cd457};
test_bias[4670:4670] = '{32'hc05258ea};
test_output[4670:4670] = '{32'h4689f067};
test_input[37368:37375] = '{32'hc2799962, 32'hc2061a4d, 32'hc1023654, 32'hc1f9940e, 32'hbeebdcd5, 32'h42205454, 32'h4203f973, 32'h42c77216};
test_weights[37368:37375] = '{32'hbe857bd4, 32'h4296527f, 32'hc205b04d, 32'h414a5ef1, 32'h42a82aaa, 32'hc1b93cc5, 32'hc2be108c, 32'hc20e71f9};
test_bias[4671:4671] = '{32'hc2ad3c76};
test_output[4671:4671] = '{32'hc621f942};
test_input[37376:37383] = '{32'hc271a8c4, 32'hc247ba59, 32'h415a07fb, 32'h426aa60b, 32'h4281d245, 32'hc2b13310, 32'hc0c55104, 32'hc24520d6};
test_weights[37376:37383] = '{32'h425cf73b, 32'hc2b9c26a, 32'hc2c43ded, 32'h405c248b, 32'hc098c4b0, 32'h41d70387, 32'hc23e95a1, 32'h40e16b9a};
test_bias[4672:4672] = '{32'h4268e427};
test_output[4672:4672] = '{32'hc51d9575};
test_input[37384:37391] = '{32'h40cf1619, 32'hc24b93e4, 32'hc2c6ce5e, 32'hc226cdec, 32'hc22959ba, 32'h429b1aac, 32'hc2043ffd, 32'h418cd9f5};
test_weights[37384:37391] = '{32'hc27cb26f, 32'hc0c63124, 32'h42bc4da4, 32'hc29eee32, 32'h42c26202, 32'hc2833480, 32'h421b7f0c, 32'hc258c322};
test_bias[4673:4673] = '{32'h421d4a5a};
test_output[4673:4673] = '{32'hc6890a9e};
test_input[37392:37399] = '{32'h42bef2ba, 32'hc28dd68d, 32'h42404b29, 32'hc21a27fd, 32'h425b73ad, 32'h42bd9756, 32'hc27d55b5, 32'h42140a44};
test_weights[37392:37399] = '{32'hc135459b, 32'h42bc4892, 32'h4251be4f, 32'h41c6c261, 32'h42ade719, 32'h42c53325, 32'h422b4a57, 32'h42b45abd};
test_bias[4674:4674] = '{32'hc2835a9a};
test_output[4674:4674] = '{32'h46048847};
test_input[37400:37407] = '{32'h41863756, 32'hc0c93ad5, 32'hc22e3285, 32'h42305b68, 32'hbff783cd, 32'h42720de8, 32'h428e4677, 32'hc2b7e9da};
test_weights[37400:37407] = '{32'hc2a61686, 32'hc08a9598, 32'hc2003718, 32'h428431c4, 32'hc1796e3c, 32'hc2448803, 32'h42a59864, 32'h41427408};
test_bias[4675:4675] = '{32'hc2ba6981};
test_output[4675:4675] = '{32'h45924248};
test_input[37408:37415] = '{32'hc0c07da6, 32'hc206e049, 32'h42c1159e, 32'hc2719865, 32'hc141ffd9, 32'h42691460, 32'hbf8cce17, 32'hc2b9dcb6};
test_weights[37408:37415] = '{32'hc1d95182, 32'hc2276fbd, 32'hc2bb43c1, 32'h4281acbf, 32'h428fa168, 32'h41c31448, 32'hc2b3bb01, 32'h424a18ca};
test_bias[4676:4676] = '{32'h413a447c};
test_output[4676:4676] = '{32'hc670dd61};
test_input[37416:37423] = '{32'hc1927c2c, 32'hc298846a, 32'hc2ab1913, 32'h423c5896, 32'hc2c58ca5, 32'hc1b8a031, 32'hc24bf4d1, 32'h42046477};
test_weights[37416:37423] = '{32'hc2348972, 32'hc2a6aea1, 32'hc0c8ae2a, 32'h4266833c, 32'hc282eb1d, 32'hc1fccd57, 32'hc2b37908, 32'h42195775};
test_bias[4677:4677] = '{32'hc24cb90b};
test_output[4677:4677] = '{32'h46b6f845};
test_input[37424:37431] = '{32'h41730d95, 32'h41cecc5f, 32'hc1e05727, 32'hc20074bb, 32'hc280625b, 32'h42acb78e, 32'h4242f67b, 32'hc2806434};
test_weights[37424:37431] = '{32'hc2663edb, 32'hc2a01d09, 32'h42440355, 32'hc1bf59bd, 32'h429c5cfd, 32'h42366f57, 32'hc0b0ca7b, 32'h428d6b09};
test_bias[4678:4678] = '{32'h42990b9d};
test_output[4678:4678] = '{32'hc6124743};
test_input[37432:37439] = '{32'hc29cc969, 32'hc2690891, 32'hc2580d5f, 32'hc23e42bf, 32'h40dad800, 32'h41ded8f1, 32'h426678a0, 32'h42541961};
test_weights[37432:37439] = '{32'h41857b5e, 32'hc29556c4, 32'h419a1625, 32'h41a04a58, 32'hc2a2ee38, 32'h42804251, 32'h420784f7, 32'h41727b8d};
test_bias[4679:4679] = '{32'h4254a36d};
test_output[4679:4679] = '{32'h459ef6bb};
test_input[37440:37447] = '{32'h409984b7, 32'hc18de239, 32'h422e94d4, 32'h424fb349, 32'h40f303e7, 32'h41818d11, 32'hc2ae0aea, 32'hc29cef34};
test_weights[37440:37447] = '{32'h428e4514, 32'hc26b12ce, 32'hc28a119a, 32'hc2b3f738, 32'h428e3bc1, 32'hc2014b26, 32'h421df8d0, 32'h4293f40d};
test_bias[4680:4680] = '{32'hc1b17094};
test_output[4680:4680] = '{32'hc672f373};
test_input[37448:37455] = '{32'hc2951b86, 32'hc1b5d8d6, 32'h42b63f20, 32'h42ae7d27, 32'hc271aaa0, 32'hc2279853, 32'hc268a453, 32'h42c328f7};
test_weights[37448:37455] = '{32'h41782f2f, 32'hc1d72778, 32'hc2471278, 32'hc2600bdc, 32'h41f166b0, 32'h42539adb, 32'hc25f6786, 32'hc237fc64};
test_bias[4681:4681] = '{32'hc1dee69e};
test_output[4681:4681] = '{32'hc66ea925};
test_input[37456:37463] = '{32'h42bfd190, 32'h429098a2, 32'h41dbbad9, 32'hc256c590, 32'hc29dce05, 32'hc194dec6, 32'hc2739702, 32'h4294a00c};
test_weights[37456:37463] = '{32'h423d8175, 32'hc18a3862, 32'h420a2c6b, 32'h4228b79f, 32'hc2b54c9c, 32'h424247b0, 32'h42ab9eac, 32'hc2c1d6a8};
test_bias[4682:4682] = '{32'h414e9839};
test_output[4682:4682] = '{32'hc582dcf6};
test_input[37464:37471] = '{32'hc28c3548, 32'h413494b8, 32'hc2b5d37b, 32'hc27b18ad, 32'hc2b5ea52, 32'hc283407d, 32'hc14031a2, 32'hc10b957f};
test_weights[37464:37471] = '{32'h429ef421, 32'hc280d364, 32'hc2af5c28, 32'hc28059d6, 32'h42a96ada, 32'hc22438af, 32'h41a30801, 32'hc21effb9};
test_bias[4683:4683] = '{32'hc2704975};
test_output[4683:4683] = '{32'h44371ef5};
test_input[37472:37479] = '{32'h4298255f, 32'h41fc880b, 32'h42471669, 32'h4285e301, 32'hc2c56f8d, 32'hc1c19308, 32'h41ccb92b, 32'hc1cadaa1};
test_weights[37472:37479] = '{32'hc277fd2c, 32'hc28c5a35, 32'hc1151c56, 32'hc119cec2, 32'h42849b35, 32'h40972435, 32'hc07630b4, 32'hc2869219};
test_bias[4684:4684] = '{32'h4280a921};
test_output[4684:4684] = '{32'hc64b89d5};
test_input[37480:37487] = '{32'h427fecd8, 32'h420696da, 32'h41d52f60, 32'h428573a5, 32'h425892d7, 32'hc2aebd84, 32'hc2301478, 32'hc2a0081a};
test_weights[37480:37487] = '{32'h428ab0c8, 32'h423af0ad, 32'hc207cedd, 32'h41dd4bf4, 32'h42665124, 32'hc2334ffe, 32'hc1695128, 32'hc2a48058};
test_bias[4685:4685] = '{32'h42b54109};
test_output[4685:4685] = '{32'h46a664cc};
test_input[37488:37495] = '{32'hc20224a8, 32'hc2b4d172, 32'h42b94f5b, 32'h41d78cac, 32'hc2a884c2, 32'hc26d88d4, 32'hc270086d, 32'hc279d222};
test_weights[37488:37495] = '{32'hc2ab0e68, 32'h42b23fa7, 32'h41aeb2d5, 32'h4283cc05, 32'hc0e26a88, 32'h41ec494a, 32'h422c9ef1, 32'hc20f7890};
test_bias[4686:4686] = '{32'h415a0c5b};
test_output[4686:4686] = '{32'hc5399b70};
test_input[37496:37503] = '{32'hc2bd314f, 32'hc193044b, 32'hc288eb54, 32'h42aba968, 32'h409d8a67, 32'hc1a2bee4, 32'h4293531c, 32'h423228d4};
test_weights[37496:37503] = '{32'h42bc11e9, 32'hc209cae7, 32'hc2a048d1, 32'hc2781d2b, 32'h42a487b9, 32'h41f53d19, 32'hc1d50ea2, 32'h42a8f79a};
test_bias[4687:4687] = '{32'h421ab4d6};
test_output[4687:4687] = '{32'hc5ca74be};
test_input[37504:37511] = '{32'hc2097b9e, 32'hc19ad009, 32'hc29a062c, 32'h42a9b08f, 32'h427ad1f2, 32'h428fa4da, 32'hc283b807, 32'hc2019dc2};
test_weights[37504:37511] = '{32'hc277d500, 32'h42947805, 32'h42b72009, 32'h421bf3d0, 32'hc2315a75, 32'h41109762, 32'h422ff948, 32'h40aee9ea};
test_bias[4688:4688] = '{32'h429b64d8};
test_output[4688:4688] = '{32'hc5ff93e5};
test_input[37512:37519] = '{32'h421aac57, 32'hc19d5c68, 32'h4298de8b, 32'h42736778, 32'h41bae9ea, 32'h408a450c, 32'h421e410f, 32'h41e097b0};
test_weights[37512:37519] = '{32'h42377e4f, 32'h418b4330, 32'h41cba5cf, 32'hc2bceac9, 32'h42a9eb6d, 32'hc1624d32, 32'h4206f135, 32'hc249462d};
test_bias[4689:4689] = '{32'hc278a73c};
test_output[4689:4689] = '{32'hc412bd77};
test_input[37520:37527] = '{32'hc2958f41, 32'hc296b892, 32'hc1fb1fe0, 32'h4245d8a8, 32'h423893c7, 32'hc29428a3, 32'hc2b911ed, 32'hc299b07a};
test_weights[37520:37527] = '{32'hc29fb7c0, 32'h40142e9f, 32'h418f4ae6, 32'h4294f142, 32'h428251ab, 32'h42770369, 32'hc225d6e6, 32'h42b4700c};
test_bias[4690:4690] = '{32'hbfc77e9b};
test_output[4690:4690] = '{32'h4584e5ec};
test_input[37528:37535] = '{32'hc23f593a, 32'hc247a14e, 32'h42281143, 32'h412592ab, 32'hc24a07e3, 32'hc21bd261, 32'hc18eb56b, 32'h41ffbd26};
test_weights[37528:37535] = '{32'hc038b7d8, 32'hc0b17a28, 32'hc2b42b70, 32'hc2a0d08b, 32'h429d6231, 32'h42aad577, 32'h42b3a6ed, 32'h41f87a46};
test_bias[4691:4691] = '{32'hc0ac01b6};
test_output[4691:4691] = '{32'hc63d5c90};
test_input[37536:37543] = '{32'hc293c8bd, 32'hc101e642, 32'h429a195a, 32'h3f597c1d, 32'h3f8c7d2b, 32'h42870d4d, 32'hc1a5cba0, 32'h422f18c6};
test_weights[37536:37543] = '{32'h429eaf36, 32'hc2c7e8d9, 32'h42435573, 32'hc217b922, 32'hc19b5bbd, 32'hc29a6b63, 32'hc1cc71dd, 32'hc2835a12};
test_bias[4692:4692] = '{32'hc0b95670};
test_output[4692:4692] = '{32'hc60b2bc3};
test_input[37544:37551] = '{32'h426663cc, 32'hc0de710a, 32'hc0b36ae8, 32'h41d8d9bb, 32'hc1bb3ba6, 32'hc25d8f93, 32'hc14762a0, 32'hc28cb994};
test_weights[37544:37551] = '{32'hc26fbb33, 32'h42be15b8, 32'hc2a87fa7, 32'hc1183f04, 32'h424f19bb, 32'h428e3501, 32'h42a071b0, 32'h425543b4};
test_bias[4693:4693] = '{32'h410fea6e};
test_output[4693:4693] = '{32'hc6577a2f};
test_input[37552:37559] = '{32'h42c2c93a, 32'hc2149e53, 32'h429c13cd, 32'h42347d79, 32'hc2a4e3c5, 32'hc245eb52, 32'h41cd311e, 32'h4227f81c};
test_weights[37552:37559] = '{32'hc28edad9, 32'hc1dee79b, 32'h417d26c0, 32'h424c7cc0, 32'h41aa6d58, 32'hc2632990, 32'h4074bfe8, 32'hc23f2183};
test_bias[4694:4694] = '{32'hc2c28589};
test_output[4694:4694] = '{32'hc5503de2};
test_input[37560:37567] = '{32'h3e038625, 32'h4205b0b3, 32'h42959a37, 32'h4279ceb5, 32'h3f3913a2, 32'h418cbc8f, 32'h4247bf2d, 32'h4241b51d};
test_weights[37560:37567] = '{32'h42222beb, 32'h4036b4b3, 32'h41a3f3fa, 32'h42b7645d, 32'h3fe68c0d, 32'hc182d59a, 32'h42c219fe, 32'h419a2d54};
test_bias[4695:4695] = '{32'hc23d9825};
test_output[4695:4695] = '{32'h4648184e};
test_input[37568:37575] = '{32'h42ad890e, 32'h42b17ec9, 32'h42329c62, 32'hc2a6ac0d, 32'h42bbe974, 32'hc12cb231, 32'h4257718f, 32'h4292835e};
test_weights[37568:37575] = '{32'h41ecc044, 32'h42a86bbf, 32'h426ddb8f, 32'hc03d5411, 32'hc2091e41, 32'hc29f4951, 32'hc29ce850, 32'hc250c275};
test_bias[4696:4696] = '{32'h4220918c};
test_output[4696:4696] = '{32'h4520d353};
test_input[37576:37583] = '{32'hc2a90cc8, 32'hc16ad9ed, 32'hc1e61bcc, 32'h3f9e148f, 32'h41c89beb, 32'h425a32ce, 32'h42a31430, 32'hc1897ed6};
test_weights[37576:37583] = '{32'h4297392e, 32'hc2308f01, 32'hc19486ba, 32'h425e70e0, 32'h428b7c80, 32'h41dfb432, 32'h421ca467, 32'hc29675fc};
test_bias[4697:4697] = '{32'h4268f3f1};
test_output[4697:4697] = '{32'h452761ea};
test_input[37584:37591] = '{32'hc28ce016, 32'hc25ad0db, 32'hc2c5491c, 32'hc1fc0320, 32'h42ad4b64, 32'h4253bfcb, 32'h42436673, 32'hc2a4324b};
test_weights[37584:37591] = '{32'h42aa4f9b, 32'h4286081d, 32'h4286e6be, 32'h42bc925c, 32'hc2b0dc6e, 32'h420baa1a, 32'h42163da6, 32'hc25a8d5b};
test_bias[4698:4698] = '{32'hc29a1537};
test_output[4698:4698] = '{32'hc6935494};
test_input[37592:37599] = '{32'h423350ed, 32'hc2374c01, 32'hc203e6d3, 32'hc12a6305, 32'h41e6fe12, 32'hc27633d4, 32'hc24cfc6b, 32'h42ac1292};
test_weights[37592:37599] = '{32'hc0a32421, 32'h4269ca00, 32'h4223259a, 32'h429d6fd6, 32'hbf475065, 32'hc2718037, 32'h4299eedd, 32'h428fd851};
test_bias[4699:4699] = '{32'h420b4db4};
test_output[4699:4699] = '{32'h445c8405};
test_input[37600:37607] = '{32'h4183a11b, 32'h42ab6fe5, 32'h421f74c1, 32'hc0c05ace, 32'hc297db72, 32'h42a9ae66, 32'hc0eb50e0, 32'h42b0fe26};
test_weights[37600:37607] = '{32'h4294e323, 32'hc2708acc, 32'hc2646118, 32'h422f37bb, 32'h420b2919, 32'hc293bf13, 32'hc299785f, 32'h41df168d};
test_bias[4700:4700] = '{32'h42bec401};
test_output[4700:4700] = '{32'hc63f6af7};
test_input[37608:37615] = '{32'hc2c43f8b, 32'hc11be486, 32'h4264dd5e, 32'h42930e88, 32'h4299ec33, 32'h4260d007, 32'h41ffef5b, 32'h42329f26};
test_weights[37608:37615] = '{32'hc2b29ee9, 32'h42c3a639, 32'hc1f62afc, 32'hc20f36ea, 32'hc2b1bace, 32'hc20e45b3, 32'hc16f8977, 32'hc2868424};
test_bias[4701:4701] = '{32'h429d8a71};
test_output[4701:4701] = '{32'hc609e284};
test_input[37616:37623] = '{32'hc06af23f, 32'hc218cf06, 32'hc13a36dc, 32'hc2023359, 32'h41ef52ea, 32'h4231429d, 32'h42c73c05, 32'hc2a74a10};
test_weights[37616:37623] = '{32'hc294111a, 32'hc2b99634, 32'h3fe2c432, 32'hc2c41c63, 32'h419019d3, 32'hbfb4e564, 32'hc1ddee0f, 32'hc1eef135};
test_bias[4702:4702] = '{32'h42c23e0a};
test_output[4702:4702] = '{32'h45e3ff48};
test_input[37624:37631] = '{32'h401e30aa, 32'h429d33d0, 32'hc2983a16, 32'h401f6a64, 32'hc27f9357, 32'hc1cc5749, 32'h426e0fa5, 32'hbdbc85ec};
test_weights[37624:37631] = '{32'hc22219cd, 32'hc2063309, 32'hc16a842c, 32'hc2aa4e9b, 32'h42b34fcd, 32'h42c277b6, 32'hc086dec9, 32'hc2b04f6b};
test_bias[4703:4703] = '{32'hc0ea5930};
test_output[4703:4703] = '{32'hc620df52};
test_input[37632:37639] = '{32'hc2aa18fa, 32'h42a9b9e9, 32'hc29debd6, 32'h428e36e2, 32'hc1b3c51f, 32'h4278f7ba, 32'hc2800728, 32'hc248cdce};
test_weights[37632:37639] = '{32'h426e382b, 32'h42b83088, 32'h40db08e2, 32'h41b13c3f, 32'hc17476e1, 32'hc16a1103, 32'hbf272e34, 32'hc29c567c};
test_bias[4704:4704] = '{32'h429de803};
test_output[4704:4704] = '{32'h45e2f7a3};
test_input[37640:37647] = '{32'hc2c2ac2d, 32'hc2ba357c, 32'hc2851af1, 32'h42b99f0b, 32'hc2892333, 32'h42acf34d, 32'hc2beb8fa, 32'hc1fa3f50};
test_weights[37640:37647] = '{32'h42328283, 32'hc06144a0, 32'h41c5f7bb, 32'hc29acccd, 32'h4289b94c, 32'hc0871577, 32'h4264a3f7, 32'hc29e339a};
test_bias[4705:4705] = '{32'h425905c2};
test_output[4705:4705] = '{32'hc6a2ef62};
test_input[37648:37655] = '{32'hc2aa3c1d, 32'h41cec28c, 32'hc2c27fcb, 32'h415e5545, 32'hc2ab2858, 32'hc1542c26, 32'hc274b475, 32'hc0b4d081};
test_weights[37648:37655] = '{32'hc2a47af2, 32'hc10cd296, 32'h42959438, 32'h423bad61, 32'hc2ab9c1b, 32'hc27a82e2, 32'hc2aa818b, 32'hc1e52352};
test_bias[4706:4706] = '{32'h424b04c7};
test_output[4706:4706] = '{32'h4656e3d3};
test_input[37656:37663] = '{32'h41a191a0, 32'h425f2af6, 32'h42245b13, 32'h42a91799, 32'hc2b55594, 32'hc2c3122f, 32'h42ab0551, 32'hc162baba};
test_weights[37656:37663] = '{32'hc21d04a1, 32'h418aa843, 32'h4293d6a1, 32'hc205c3ae, 32'h42c10c2b, 32'h422f1eaf, 32'hc1e7b72e, 32'h42bb3d2f};
test_bias[4707:4707] = '{32'h42a4afe7};
test_output[4707:4707] = '{32'hc67f9a2b};
test_input[37664:37671] = '{32'h41c53616, 32'hc2567dea, 32'hc114b278, 32'h4100c860, 32'hc2b664f4, 32'h4187fd34, 32'h415457e1, 32'h42b7d200};
test_weights[37664:37671] = '{32'h42973601, 32'hc20c26f8, 32'hc27db08f, 32'hc29a07bf, 32'h427e8549, 32'hc230efa9, 32'h416f3974, 32'hc1c9b41b};
test_bias[4708:4708] = '{32'h41d3ee75};
test_output[4708:4708] = '{32'hc59a3874};
test_input[37672:37679] = '{32'hc2357f2f, 32'h40c02970, 32'hc2b805c7, 32'h4162a426, 32'hc11ff885, 32'hc21729dd, 32'h42b27967, 32'h4237f55d};
test_weights[37672:37679] = '{32'h42502617, 32'hc15871f3, 32'hc1d03bb4, 32'h422eaffe, 32'h42bba853, 32'h41a817cc, 32'hc2c79881, 32'h409c377e};
test_bias[4709:4709] = '{32'h423f6f30};
test_output[4709:4709] = '{32'hc6190908};
test_input[37680:37687] = '{32'h429a8194, 32'h429c68eb, 32'hc268aa38, 32'h42b794f7, 32'hc293bab0, 32'h41dba71b, 32'h42b21960, 32'hc21f3abc};
test_weights[37680:37687] = '{32'h428f8c43, 32'h40bfaf35, 32'hc1d16a87, 32'h42a07298, 32'hc2862015, 32'h42c3cf3b, 32'h42ad99e5, 32'h41a345b1};
test_bias[4710:4710] = '{32'hc1dab532};
test_output[4710:4710] = '{32'h46e5ee42};
test_input[37688:37695] = '{32'h42bcc36b, 32'hc1d870aa, 32'h42276794, 32'hc2c13221, 32'hc291498c, 32'hc2a8f783, 32'hc1b501b9, 32'h42525b46};
test_weights[37688:37695] = '{32'h42b965d5, 32'hc20dddc1, 32'h42609e27, 32'h425e5992, 32'h409127cc, 32'hc222e737, 32'h4238c868, 32'h42928692};
test_bias[4711:4711] = '{32'hc21e74c0};
test_output[4711:4711] = '{32'h46446103};
test_input[37696:37703] = '{32'h4277c9d8, 32'hc117de6d, 32'hc29ce496, 32'hc118bf54, 32'h4231f97e, 32'hc26f9e3c, 32'hc2733f09, 32'h427c2f29};
test_weights[37696:37703] = '{32'hc16d7917, 32'hc261ce77, 32'hc1a69fb1, 32'h429ea2bd, 32'h425144fa, 32'h42594109, 32'hc00153a4, 32'hc0ea17ce};
test_bias[4712:4712] = '{32'hbfdfbd1d};
test_output[4712:4712] = '{32'hc441361d};
test_input[37704:37711] = '{32'h42c6aa3a, 32'hc2ad764e, 32'h42945400, 32'hc2866201, 32'hc2350229, 32'h4126dfe1, 32'h427f38c0, 32'h4272ed6f};
test_weights[37704:37711] = '{32'h41f7fc87, 32'hc22527e7, 32'hc1681a43, 32'h41bf9805, 32'hc2bf49f2, 32'h4281b4a9, 32'h42960698, 32'h427028a3};
test_bias[4713:4713] = '{32'h42134b8e};
test_output[4713:4713] = '{32'h46885208};
test_input[37712:37719] = '{32'h410fc5d4, 32'h423e1cb3, 32'h42bd8663, 32'hc2810eea, 32'hc1835727, 32'hc1ad6e3e, 32'h42592a14, 32'h418b491c};
test_weights[37712:37719] = '{32'hc06d999c, 32'hc2a4448e, 32'h4226abbe, 32'hc21ae23e, 32'hc29875b8, 32'h42607ba7, 32'hc246220e, 32'h42bf6cda};
test_bias[4714:4714] = '{32'h42a2b3f4};
test_output[4714:4714] = '{32'h44c87287};
test_input[37720:37727] = '{32'hc1a3719e, 32'h42031659, 32'h42be2bec, 32'h4118ac32, 32'h42bf5a42, 32'hc2b80792, 32'h4157faf4, 32'h429bfc93};
test_weights[37720:37727] = '{32'h420142a8, 32'h420552e4, 32'hc2bb0d45, 32'h411c335a, 32'hc1e394dc, 32'hc28811cb, 32'h41ab5a77, 32'h42372f41};
test_bias[4715:4715] = '{32'h4135f810};
test_output[4715:4715] = '{32'hc46f3fac};
test_input[37728:37735] = '{32'h425b0fdc, 32'h41c3d885, 32'h42acc4f3, 32'h4271707e, 32'h42232a6e, 32'h41afb043, 32'h413620cf, 32'h418405e1};
test_weights[37728:37735] = '{32'h41a5dc32, 32'h4179ebd6, 32'h4226dc27, 32'h418bcd55, 32'h41de3a5e, 32'hc1926b17, 32'h4288a0e7, 32'h42a0d4cc};
test_bias[4716:4716] = '{32'h42453f4b};
test_output[4716:4716] = '{32'h460d9577};
test_input[37736:37743] = '{32'h3eac25f0, 32'hc142c7fb, 32'h41a7a6ca, 32'h4216c227, 32'h4257c389, 32'h3fe2e83f, 32'h41a7f184, 32'h42a2a51b};
test_weights[37736:37743] = '{32'h41c9b4a7, 32'hc16bcf11, 32'hc15e30d5, 32'h3e75d91e, 32'hc2a71ecc, 32'h4189fd35, 32'hc2bd4a96, 32'hc2acb4c1};
test_bias[4717:4717] = '{32'hc27b195c};
test_output[4717:4717] = '{32'hc6552bae};
test_input[37744:37751] = '{32'hc2c15e35, 32'hc29ca0cc, 32'hc25067b5, 32'h41992f75, 32'h429ab575, 32'h424b5a2b, 32'h42b21006, 32'hc2811dac};
test_weights[37744:37751] = '{32'h42579e00, 32'h429f0520, 32'h42933a1f, 32'h423862b7, 32'hc206e73e, 32'h4257ad26, 32'h40b0cc7b, 32'h40b5cc16};
test_bias[4718:4718] = '{32'hc22ea253};
test_output[4718:4718] = '{32'hc65d8570};
test_input[37752:37759] = '{32'hc2c1ea03, 32'h41c684c8, 32'h421a1b0e, 32'h420a3692, 32'hc2199fd6, 32'h429c79c4, 32'hc2ae3401, 32'h42260785};
test_weights[37752:37759] = '{32'hc2c6a2a4, 32'h41e530c3, 32'hc182710c, 32'hc239d372, 32'hc236e7e3, 32'hc2c42214, 32'h42a09168, 32'hc212e6b4};
test_bias[4719:4719] = '{32'hc2a7468e};
test_output[4719:4719] = '{32'hc5c85137};
test_input[37760:37767] = '{32'h415b0d0c, 32'hc29c93a6, 32'hc2bf0b0d, 32'hc2836894, 32'h4219f4ef, 32'h42b20375, 32'hc2298147, 32'hc26fc708};
test_weights[37760:37767] = '{32'hc29c8df8, 32'h42a2d586, 32'h42b2dd66, 32'hc27c2bd9, 32'h3ff5c799, 32'hc288a59a, 32'h40d60fa6, 32'hc2acf530};
test_bias[4720:4720] = '{32'hc29f1769};
test_output[4720:4720] = '{32'hc64ba2a4};
test_input[37768:37775] = '{32'hc1f18225, 32'hc2a641fe, 32'h41a0bc34, 32'hc2831813, 32'h4216e5ae, 32'h428fe07d, 32'h42816f8f, 32'h4281f6d8};
test_weights[37768:37775] = '{32'hc28289ec, 32'h4272119d, 32'hc1dbf913, 32'hc255d8bc, 32'hc2c1dc6b, 32'hc2900551, 32'hbf1d4806, 32'hc271cae2};
test_bias[4721:4721] = '{32'h41362665};
test_output[4721:4721] = '{32'hc64997b0};
test_input[37776:37783] = '{32'h42a9295e, 32'hc2c6b52f, 32'hc24f2dc1, 32'h42be4399, 32'hc1919c7a, 32'hc2839dfd, 32'h423ef3b6, 32'hc2471a54};
test_weights[37776:37783] = '{32'hc286e6ab, 32'hc0cdfc29, 32'hc22c0289, 32'hc1a46428, 32'h42190bd9, 32'h42683772, 32'h4291dd5e, 32'hc26ad291};
test_bias[4722:4722] = '{32'h421d0bd8};
test_output[4722:4722] = '{32'hc5332e38};
test_input[37784:37791] = '{32'h428849e9, 32'h42996bb6, 32'hbf0dce56, 32'h4112e46c, 32'hc12c8cc8, 32'hc2ad19a9, 32'h41abff42, 32'hc26ab656};
test_weights[37784:37791] = '{32'h42c45d60, 32'hc28e63e8, 32'h421d483b, 32'hc245dc60, 32'h4136c078, 32'hc29c5797, 32'h3da52ca6, 32'h429ae488};
test_bias[4723:4723] = '{32'h40b13996};
test_output[4723:4723] = '{32'h4532aaae};
test_input[37792:37799] = '{32'hc1e9f4e9, 32'h42950532, 32'h4216a897, 32'hc26f0ec8, 32'hc28c697b, 32'h423bc56f, 32'hc2aee985, 32'h41d53f35};
test_weights[37792:37799] = '{32'h4263712a, 32'h42c4010a, 32'hc17fe0f3, 32'hc28ff7ef, 32'h42877ef6, 32'h407dc59d, 32'h415ba39f, 32'hc2508ab1};
test_bias[4724:4724] = '{32'h42a782ee};
test_output[4724:4724] = '{32'h450d658a};
test_input[37800:37807] = '{32'h41e994bb, 32'hc2818aaa, 32'h403f0ab5, 32'h422b7806, 32'h41d97ca4, 32'hc1bf1876, 32'hc286b86f, 32'h424cf90b};
test_weights[37800:37807] = '{32'hc2609747, 32'h4172d2ac, 32'h40c38487, 32'h41a6ef52, 32'h4297ac6d, 32'hc1f8c260, 32'hc2931dd1, 32'h4265c0dc};
test_bias[4725:4725] = '{32'hc265c771};
test_output[4725:4725] = '{32'h460b9e67};
test_input[37808:37815] = '{32'h422c4143, 32'hc26c4616, 32'h42182d52, 32'h428d0a74, 32'hc04d2583, 32'hc28b5267, 32'h422b45fb, 32'h429170d2};
test_weights[37808:37815] = '{32'hc28032ea, 32'hc24dcb91, 32'hc2822064, 32'h420d13cf, 32'hc16185be, 32'h42a0d36b, 32'h4276e5ee, 32'h42140674};
test_bias[4726:4726] = '{32'hc27cd7a4};
test_output[4726:4726] = '{32'h409e5674};
test_input[37816:37823] = '{32'h426e7912, 32'hc1dbf4a5, 32'hc26d7c3c, 32'hc22d32a5, 32'hc2b0f7a6, 32'h425f647b, 32'hc1b005ce, 32'hc28dc66f};
test_weights[37816:37823] = '{32'hc1fd7fa9, 32'h415b21a5, 32'h429fde71, 32'hc186601b, 32'h42861dc5, 32'h417ae8ec, 32'hc0e00ad5, 32'hc2659641};
test_bias[4727:4727] = '{32'hc1e5aad3};
test_output[4727:4727] = '{32'hc5df5f47};
test_input[37824:37831] = '{32'hc20374bf, 32'h418ff110, 32'hc29eac38, 32'hc18b1ae3, 32'h42ab4e9e, 32'h42775757, 32'h4296328e, 32'hc1c5fd6c};
test_weights[37824:37831] = '{32'hc246d7ba, 32'hc1b25bf4, 32'h408b55e9, 32'h42244d5e, 32'hc22c888b, 32'h42014802, 32'hc1bc3ee1, 32'h428e66b9};
test_bias[4728:4728] = '{32'h41765c11};
test_output[4728:4728] = '{32'hc59d67c6};
test_input[37832:37839] = '{32'h404cf7ce, 32'hc1f10c4d, 32'hc134e2f6, 32'h428113cc, 32'h4286e3b6, 32'hc295aa21, 32'h413e2494, 32'hbcd42ed1};
test_weights[37832:37839] = '{32'hc1694341, 32'h41d19fa2, 32'h429ae22e, 32'hc25cd502, 32'h42386ebc, 32'h3fd568e6, 32'h41761114, 32'h4184ec66};
test_bias[4729:4729] = '{32'hc28ea923};
test_output[4729:4729] = '{32'hc5082c88};
test_input[37840:37847] = '{32'hc206f74c, 32'hc291218a, 32'h42b7327b, 32'hc2c029a2, 32'h42938fe2, 32'hc28a8ffe, 32'hc0d642b9, 32'hc1254f10};
test_weights[37840:37847] = '{32'hc1d5d33e, 32'hc23030c8, 32'h417738d4, 32'hc08bcda7, 32'hc1351754, 32'h41b09af6, 32'h42a11a1f, 32'hc1e017c7};
test_bias[4730:4730] = '{32'h41ea7bae};
test_output[4730:4730] = '{32'h4551428a};
test_input[37848:37855] = '{32'h427bd115, 32'hc2c13469, 32'h4235f80b, 32'hc1fe4668, 32'h4240c307, 32'hc2816d26, 32'hc26cc24e, 32'h41774d63};
test_weights[37848:37855] = '{32'h417b4249, 32'hc130b36f, 32'h4288d0b2, 32'h40790b4d, 32'hc1875b26, 32'hc2be8cb1, 32'hc2bb7335, 32'hc14ef7fb};
test_bias[4731:4731] = '{32'hc28cca43};
test_output[4731:4731] = '{32'h4674dcd3};
test_input[37856:37863] = '{32'h416aa2fd, 32'h42c027bf, 32'hc1c12ce0, 32'h409536c7, 32'hc2c129f7, 32'hc2328e06, 32'hc2715e57, 32'hc2684cff};
test_weights[37856:37863] = '{32'hc28d2d04, 32'hc1dbb1f7, 32'hc206fa7f, 32'hc28076ae, 32'hc132523b, 32'h429eb5b0, 32'hc06ae6f3, 32'hc160df3e};
test_bias[4732:4732] = '{32'hc2168d65};
test_output[4732:4732] = '{32'hc590811d};
test_input[37864:37871] = '{32'hc2b0d7ee, 32'h429dcd12, 32'hc29bdef7, 32'h42a6ac43, 32'hc2a11c03, 32'hc2a00cd1, 32'h4292df2c, 32'h42947244};
test_weights[37864:37871] = '{32'hc2c0aa5e, 32'hc213944e, 32'h42816d4a, 32'h427721e6, 32'hc2b47d15, 32'h42b0c701, 32'hc258c8e8, 32'h426639b9};
test_bias[4733:4733] = '{32'h42002a79};
test_output[4733:4733] = '{32'h45c2c4d9};
test_input[37872:37879] = '{32'hc244d999, 32'h42a9a3f6, 32'h42be988f, 32'hc2a3b592, 32'hc2918aeb, 32'hc2894bc5, 32'h429c0fd9, 32'hc22c65b3};
test_weights[37872:37879] = '{32'hc204dba4, 32'h41b75116, 32'h422553d2, 32'h414ad3fd, 32'hc2bd60c1, 32'h4299ee76, 32'hc2988b96, 32'hc2c0fa3a};
test_bias[4734:4734] = '{32'hc260f138};
test_output[4734:4734] = '{32'h45c2e9b7};
test_input[37880:37887] = '{32'hc195c96b, 32'h42ab499a, 32'h40dfa5b3, 32'hc1bdb9ab, 32'h42b5d718, 32'hc2c52976, 32'hc2b11bbe, 32'h42b1f37f};
test_weights[37880:37887] = '{32'hc0982a77, 32'hc204461a, 32'h42b0da7c, 32'hc172effc, 32'h4224e7cd, 32'h41395245, 32'h42a4912c, 32'h4200f970};
test_bias[4735:4735] = '{32'hc2bc4a5a};
test_output[4735:4735] = '{32'hc56564b6};
test_input[37888:37895] = '{32'hc16dbfb7, 32'h427595c0, 32'hc2b6e48b, 32'hc16e265e, 32'h429ce21e, 32'hc299e5e8, 32'hc18f3c20, 32'hc21752bd};
test_weights[37888:37895] = '{32'hc2958954, 32'hc28e9627, 32'h41b28fd6, 32'hc24e2eed, 32'h4105ba89, 32'h41ed7294, 32'h42a4f9cf, 32'h425e9f89};
test_bias[4736:4736] = '{32'hc285fd26};
test_output[4736:4736] = '{32'hc61966d2};
test_input[37896:37903] = '{32'h428c825c, 32'h42ab8a42, 32'hc104c371, 32'hc25ba84f, 32'h4264841f, 32'hc14013a0, 32'hc21a26e3, 32'hc29d5a4a};
test_weights[37896:37903] = '{32'h4114cf56, 32'hc22589ef, 32'hc1d218c6, 32'hc2a25a3e, 32'hc23b1c08, 32'h42ba1315, 32'hbf3dca8a, 32'hc265521d};
test_bias[4737:4737] = '{32'hc11e8932};
test_output[4737:4737] = '{32'h451d774a};
test_input[37904:37911] = '{32'h42550cba, 32'h416779a5, 32'hc251be76, 32'hc2b8343c, 32'h4263715d, 32'hc19b261c, 32'h3f755aa9, 32'h424a59d8};
test_weights[37904:37911] = '{32'hc2869574, 32'hc28afe95, 32'h4177b1f1, 32'h426a0279, 32'h41ff06be, 32'h42aae5bb, 32'hc2a77208, 32'h40e7cec4};
test_bias[4738:4738] = '{32'h41f4a494};
test_output[4738:4738] = '{32'hc62134ff};
test_input[37912:37919] = '{32'h42676116, 32'hc2206bcb, 32'hc2328841, 32'hc2826ccf, 32'hc2467426, 32'hc293ef36, 32'hc2c57a54, 32'h4002b350};
test_weights[37912:37919] = '{32'hc22a404e, 32'hc2ae81f1, 32'hc20c101e, 32'hc2668ec4, 32'hc26dfff0, 32'hc0960922, 32'h42b47c70, 32'h421751f1};
test_bias[4739:4739] = '{32'h42880257};
test_output[4739:4739] = '{32'h445f21f7};
test_input[37920:37927] = '{32'hc216a402, 32'hc2a05637, 32'hc2afe05a, 32'hc2219ed8, 32'h4173a351, 32'h428163a6, 32'hc2b8f77a, 32'hc1dbe7c6};
test_weights[37920:37927] = '{32'hc2a144bf, 32'hc29295e2, 32'h42a14f1d, 32'h41ea4dac, 32'h42ba0525, 32'hc1f3d0ed, 32'h421707a9, 32'hc2c5f26d};
test_bias[4740:4740] = '{32'h42284dc3};
test_output[4740:4740] = '{32'hc4220c98};
test_input[37928:37935] = '{32'h42b8e0c5, 32'h42b64ad7, 32'hc2ace7be, 32'h42c64254, 32'hc29be4f5, 32'h41d82baa, 32'h41b56b21, 32'h41fd6b25};
test_weights[37928:37935] = '{32'hc290be2d, 32'h42aa376f, 32'hc1e05d7f, 32'hc2ae71f7, 32'hc2859e38, 32'hc2453ceb, 32'h408df10b, 32'h42bd6cbb};
test_bias[4741:4741] = '{32'hc2c6cd74};
test_output[4741:4741] = '{32'h44d7471c};
test_input[37936:37943] = '{32'hbfb603fa, 32'h429c3fa9, 32'h4140e5fa, 32'hc2953bdb, 32'h4250cc20, 32'hc290c49a, 32'hc0e7ca89, 32'h426844a9};
test_weights[37936:37943] = '{32'h429f691e, 32'hc21a3309, 32'h42473f4d, 32'hc2be529e, 32'h428e9e47, 32'h4205332d, 32'h418fcd6d, 32'hc21ca5a1};
test_bias[4742:4742] = '{32'hc29c6744};
test_output[4742:4742] = '{32'h4554da7d};
test_input[37944:37951] = '{32'hc1fa00d3, 32'hc2574e70, 32'h42993126, 32'hc25c4ed1, 32'hc2a06af2, 32'h425a7cce, 32'h4248818e, 32'hc2acce50};
test_weights[37944:37951] = '{32'h428143ea, 32'h425707b6, 32'hc2090ef4, 32'h421a8cc7, 32'h3fdaa1bc, 32'hc2c0633c, 32'h416e0419, 32'hc2aa325c};
test_bias[4743:4743] = '{32'h42715b25};
test_output[4743:4743] = '{32'hc5d793b9};
test_input[37952:37959] = '{32'h4287fb6b, 32'hc29a35c4, 32'h4292c512, 32'h419449c5, 32'h429d59f5, 32'h4257004e, 32'h42bba230, 32'hc231fe77};
test_weights[37952:37959] = '{32'h42729029, 32'h429632d7, 32'h425c05e8, 32'hc19114e0, 32'hc0fd0bc8, 32'h4296f786, 32'h42888365, 32'hc2602513};
test_bias[4744:4744] = '{32'h40e0d090};
test_output[4744:4744] = '{32'h466090e2};
test_input[37960:37967] = '{32'h426ba582, 32'h42559551, 32'hc26d4b7d, 32'hc11ac85e, 32'hc2b1af46, 32'hc1062799, 32'h42c699e5, 32'h421ac0f5};
test_weights[37960:37967] = '{32'h42981e17, 32'hc2b4fd93, 32'hc265173b, 32'hc2897dbb, 32'h40b8f29c, 32'hc220a000, 32'hc2acd365, 32'hc2585eab};
test_bias[4745:4745] = '{32'hc2872e56};
test_output[4745:4745] = '{32'hc5e134fc};
test_input[37968:37975] = '{32'hc241b57d, 32'h42bc0581, 32'hc0863ef8, 32'h42889a48, 32'h4294e166, 32'h425798a5, 32'hc21c39b4, 32'hc20a5871};
test_weights[37968:37975] = '{32'hc23ef02e, 32'h4282d313, 32'hc1a22fe4, 32'hc2a708b8, 32'hc2b37c0b, 32'hc260a498, 32'h42bcdb54, 32'h42648604};
test_bias[4746:4746] = '{32'h428bf406};
test_output[4746:4746] = '{32'hc642ae74};
test_input[37976:37983] = '{32'hc2165837, 32'hc1771dcf, 32'hc2790896, 32'h4280a915, 32'hc2c13698, 32'hc289d708, 32'hc21f4824, 32'h421b5c5a};
test_weights[37976:37983] = '{32'hc1feea8a, 32'h429d6644, 32'hc2502b6c, 32'hc18f4bb6, 32'hc1868c2b, 32'h4258ff77, 32'hc1bd261b, 32'hc28e38fa};
test_bias[4747:4747] = '{32'h4186b9d4};
test_output[4747:4747] = '{32'hc4e6f8d9};
test_input[37984:37991] = '{32'hc2bd73cc, 32'hc2b57add, 32'hc26024a9, 32'hc2210fa1, 32'hc1bd24ce, 32'h4214f2f2, 32'h4071f535, 32'h42a8a77e};
test_weights[37984:37991] = '{32'hc03b1655, 32'hc18761e6, 32'hc1da0257, 32'hc296bc21, 32'h412e7cef, 32'h4231ef44, 32'h41b37088, 32'h422a8a60};
test_bias[4748:4748] = '{32'hc1aa5df3};
test_output[4748:4748] = '{32'h46329e7e};
test_input[37992:37999] = '{32'h4243e00b, 32'hc02f0661, 32'h422e2a09, 32'hc239fa62, 32'h401789b4, 32'h42493619, 32'h427aede2, 32'h4198c155};
test_weights[37992:37999] = '{32'hc2054265, 32'h425ede84, 32'h428d47c0, 32'h41b4eeaf, 32'hc2b44de5, 32'hc1af8a80, 32'hc1df681c, 32'hc2c011a6};
test_bias[4749:4749] = '{32'hc293092c};
test_output[4749:4749] = '{32'hc593ff1a};
test_input[38000:38007] = '{32'h41f0839b, 32'h428444ce, 32'hc2767720, 32'h421f10ec, 32'h4278028f, 32'h428c05e2, 32'h41be136b, 32'h4251ff3a};
test_weights[38000:38007] = '{32'h42b92343, 32'h40dd7f71, 32'h4161a96a, 32'hc297c692, 32'h42408e31, 32'h429b4922, 32'hc230696a, 32'hc2bfef21};
test_bias[4750:4750] = '{32'h425ebec0};
test_output[4750:4750] = '{32'h44da069b};
test_input[38008:38015] = '{32'hc2971244, 32'h42437351, 32'hc206ab84, 32'h422aa129, 32'h42c59f7e, 32'hc1a9b1ac, 32'h42b03415, 32'h42894e9d};
test_weights[38008:38015] = '{32'hc29ef192, 32'h41c98035, 32'h42070857, 32'hc293ba97, 32'hc2bcd416, 32'hc2360c69, 32'h412a2f27, 32'hc2a2b534};
test_bias[4751:4751] = '{32'h423b9e48};
test_output[4751:4751] = '{32'hc61c8b21};
test_input[38016:38023] = '{32'h42b68a2f, 32'h428b3efd, 32'h41d45c5a, 32'hc1c9ba04, 32'h42990f28, 32'h429b80ee, 32'h420cb543, 32'h41ef2748};
test_weights[38016:38023] = '{32'hc2770180, 32'hc202d2d3, 32'h4290c7e1, 32'h419d226e, 32'hc25fad9d, 32'hc2ab7751, 32'h42acbd2d, 32'h4290872d};
test_bias[4752:4752] = '{32'hc1ea933b};
test_output[4752:4752] = '{32'hc63f9c24};
test_input[38024:38031] = '{32'hc2a8a66b, 32'h4293574f, 32'h422489db, 32'h421bf080, 32'hc27e87e6, 32'h42a7f328, 32'hc20917c6, 32'hc220b5f8};
test_weights[38024:38031] = '{32'hc12fee57, 32'hc2b67078, 32'h426974a4, 32'h42b4e159, 32'h4208817d, 32'h410f435d, 32'h42c5fb03, 32'hc289540e};
test_bias[4753:4753] = '{32'hc22792d9};
test_output[4753:4753] = '{32'hc4f53d04};
test_input[38032:38039] = '{32'h4294ec81, 32'h426b9307, 32'h425f564f, 32'hc13abda4, 32'hc1f94683, 32'hc2172764, 32'hc2abe0fd, 32'h4212d12e};
test_weights[38032:38039] = '{32'h4282941e, 32'h41fbd0f8, 32'h42450414, 32'h42832947, 32'hc23c76a3, 32'hc293d3d0, 32'hc2577fb2, 32'hc28b4344};
test_bias[4754:4754] = '{32'h42b02d40};
test_output[4754:4754] = '{32'h466c4dec};
test_input[38040:38047] = '{32'hc2249f98, 32'hc2ac1668, 32'h4296438a, 32'h4283c674, 32'h42a10241, 32'hc2b27f29, 32'h42c0d619, 32'h426edd82};
test_weights[38040:38047] = '{32'hc1be2f98, 32'hc2c6b5fd, 32'h428d7822, 32'h42982043, 32'h3f2803c7, 32'hc21cdcc6, 32'hc1a472c9, 32'hc2912636};
test_bias[4755:4755] = '{32'h42acd9e0};
test_output[4755:4755] = '{32'h4686315f};
test_input[38048:38055] = '{32'h427cba7d, 32'h41b10bf3, 32'h412e86aa, 32'hc21102bc, 32'h420f828f, 32'h42c77080, 32'h40d59023, 32'hc2c6fd77};
test_weights[38048:38055] = '{32'h4253a469, 32'hc2b7330a, 32'h42509ecd, 32'hc2882d8c, 32'h428fe61b, 32'h429f35f5, 32'hc2100bef, 32'h4197ead4};
test_bias[4756:4756] = '{32'hc240b3ae};
test_output[4756:4756] = '{32'h46465b57};
test_input[38056:38063] = '{32'h418d2972, 32'h4214e777, 32'hc2b0e926, 32'hc2bc4970, 32'hc2c2a949, 32'h3fdf86f2, 32'h410ac2c1, 32'hc29f3df1};
test_weights[38056:38063] = '{32'hc2460f93, 32'hc293f23c, 32'h41b7c646, 32'h4292009e, 32'hc27f934e, 32'hc01167ec, 32'h42b6f823, 32'hc15f06cc};
test_bias[4757:4757] = '{32'hc248cecb};
test_output[4757:4757] = '{32'hc58b80ac};
test_input[38064:38071] = '{32'h41bb1a54, 32'h41ef1a77, 32'hc1ba6daa, 32'hc28846c0, 32'hc20c5912, 32'hc1b8b75f, 32'hc10562f0, 32'h4189a94b};
test_weights[38064:38071] = '{32'h424a6a0e, 32'h4200670b, 32'hc2c2fd4c, 32'h428b17bb, 32'hc1a099a0, 32'hc25c9a73, 32'h423bcf2d, 32'hc1c8f58b};
test_bias[4758:4758] = '{32'h4148b0db};
test_output[4758:4758] = '{32'h4452b219};
test_input[38072:38079] = '{32'h423dce80, 32'h4282af25, 32'h4296e36f, 32'h422599ab, 32'hc2762830, 32'h415d816c, 32'hc2b59d1b, 32'hc1e08283};
test_weights[38072:38079] = '{32'h42278e88, 32'hc231c372, 32'h41c79f4a, 32'hc0cf10a8, 32'h41de1e73, 32'hc27353ae, 32'h41b43e2c, 32'hc0fb9762};
test_bias[4759:4759] = '{32'h4297fa38};
test_output[4759:4759] = '{32'hc5611903};
test_input[38080:38087] = '{32'h421b6636, 32'h425c81da, 32'hc198ac5d, 32'h4191bbae, 32'hc2af9989, 32'h4192430b, 32'hc100a03a, 32'h42910d3a};
test_weights[38080:38087] = '{32'h413e2a29, 32'hc271c6cc, 32'h42a1204f, 32'hc2131354, 32'h4264ea91, 32'h42be09c0, 32'h4248148a, 32'hc1be931f};
test_bias[4760:4760] = '{32'hc25113c9};
test_output[4760:4760] = '{32'hc624ccdf};
test_input[38088:38095] = '{32'hc1b10aec, 32'hc1a29542, 32'h41d2bf74, 32'hc2bd4072, 32'h41e1d1e4, 32'h4179c50e, 32'h421748c2, 32'hc29498ff};
test_weights[38088:38095] = '{32'hc2a3298d, 32'hc1eca10d, 32'h428e4cec, 32'h423e893b, 32'h41f6482b, 32'hc28b08a2, 32'h4004bc95, 32'hc1dc0ff2};
test_bias[4761:4761] = '{32'h424c238e};
test_output[4761:4761] = '{32'h44d85134};
test_input[38096:38103] = '{32'h40510869, 32'h40ca595f, 32'hc2762fbb, 32'hc20ecae2, 32'h421d63fa, 32'hc1e3e6d4, 32'h420851bd, 32'h429edd40};
test_weights[38096:38103] = '{32'h41dd3dda, 32'h42656ab8, 32'h4058d939, 32'h4225ea37, 32'hc1d6809f, 32'h42572429, 32'h42623e2d, 32'h41f62657};
test_bias[4762:4762] = '{32'hc0d308df};
test_output[4762:4762] = '{32'h4407614a};
test_input[38104:38111] = '{32'h426e62cf, 32'hc27ed519, 32'hc28991f9, 32'hc15ea174, 32'h41899cc6, 32'hc2667841, 32'hc06f0cf3, 32'hc2225dbc};
test_weights[38104:38111] = '{32'h42a93d8b, 32'h42656a77, 32'h423479ff, 32'h4249fc64, 32'h420b74a6, 32'h41e503c3, 32'h42c20921, 32'h422674e4};
test_bias[4763:4763] = '{32'hc26b252c};
test_output[4763:4763] = '{32'hc5ae484c};
test_input[38112:38119] = '{32'hc28ac108, 32'hc2bc9176, 32'hc2a55564, 32'h41a47c32, 32'hc1ef920e, 32'h4261dff7, 32'h419b5073, 32'hc2a0dd11};
test_weights[38112:38119] = '{32'h42a2bb0f, 32'h41f408e3, 32'hc1d7fd3a, 32'h40ce8968, 32'h428d918c, 32'h413aefa3, 32'hc116ebc2, 32'hc0ffab45};
test_bias[4764:4764] = '{32'h41a47a6d};
test_output[4764:4764] = '{32'hc5df0247};
test_input[38120:38127] = '{32'h42b069a8, 32'h41a756f4, 32'hc19acb22, 32'h427176ee, 32'h42416f27, 32'hc2b22397, 32'hc2acb638, 32'hc253b3d7};
test_weights[38120:38127] = '{32'h4099f6d7, 32'h41b2ad73, 32'hc289b8da, 32'hc26544e5, 32'h4298233e, 32'h425a4c3c, 32'hc2035ff8, 32'h42867160};
test_bias[4765:4765] = '{32'hc2ab7061};
test_output[4765:4765] = '{32'hc5499964};
test_input[38128:38135] = '{32'h429d86ca, 32'hc1d22cde, 32'h40889be5, 32'hc2a30100, 32'hc2a08b32, 32'h40c1b6c6, 32'hc2866225, 32'h40eeac7e};
test_weights[38128:38135] = '{32'h422223c8, 32'h42299ff2, 32'h420713a8, 32'hc2948bec, 32'hc25c2389, 32'h4106848f, 32'h410d72aa, 32'hc2292630};
test_bias[4766:4766] = '{32'h40ebd16c};
test_output[4766:4766] = '{32'h46390afa};
test_input[38136:38143] = '{32'h429ba252, 32'hc2459982, 32'hc2700b67, 32'hc1c27934, 32'h4164368a, 32'hc20323a9, 32'h42bfc59e, 32'h42a8ffc5};
test_weights[38136:38143] = '{32'hc1c6379f, 32'hc22687d8, 32'h42670680, 32'h42ab4a40, 32'h427aaa15, 32'h4122cd8c, 32'hc12fbf56, 32'hc1844fb0};
test_bias[4767:4767] = '{32'hc240f4c2};
test_output[4767:4767] = '{32'hc5e5f17d};
test_input[38144:38151] = '{32'h42495821, 32'hc23b9ddb, 32'h4260c093, 32'h41f0d4a3, 32'hc2b07ea1, 32'h42a5ee4f, 32'hc129476b, 32'h42c22f54};
test_weights[38144:38151] = '{32'h42465954, 32'hc1a1ad32, 32'h4217e2ed, 32'h41c0663b, 32'h425a879b, 32'hc292dc0b, 32'hc2276274, 32'hc16ee4cd};
test_bias[4768:4768] = '{32'hc2068074};
test_output[4768:4768] = '{32'hc5b0a312};
test_input[38152:38159] = '{32'h42a39f39, 32'h4086a31c, 32'h4181dbf8, 32'hc20c52fb, 32'h40f80334, 32'h42910316, 32'h428db93f, 32'hc2c30055};
test_weights[38152:38159] = '{32'h42c292a1, 32'h42aeef22, 32'h428ce5cd, 32'h41ada106, 32'hc28a0d03, 32'hc14ed0ff, 32'h42173257, 32'h42adab07};
test_bias[4769:4769] = '{32'h41028fc9};
test_output[4769:4769] = '{32'h44b62c58};
test_input[38160:38167] = '{32'h4284a48f, 32'h429d17e2, 32'h42b05f73, 32'h421f0583, 32'hc1e6f8c9, 32'hc27a63b8, 32'h41a05605, 32'hc0feb604};
test_weights[38160:38167] = '{32'hc2b6a02f, 32'hc24bde90, 32'hc1102198, 32'h426301ff, 32'hc2aff098, 32'hc2a44449, 32'hc2b8bd0c, 32'h416446d4};
test_bias[4770:4770] = '{32'hc219b5cc};
test_output[4770:4770] = '{32'hc53679e0};
test_input[38168:38175] = '{32'h3f0f2b5c, 32'hc0f9353f, 32'h41924336, 32'hc2a41797, 32'h42acc4e3, 32'hc2be03ca, 32'hbfb8d2bf, 32'hc1374908};
test_weights[38168:38175] = '{32'hc0b618e1, 32'hc225970a, 32'hc2a07150, 32'h42799b6e, 32'hc27f22ca, 32'hc200c450, 32'h41a20570, 32'h42bb3973};
test_bias[4771:4771] = '{32'hc20eb62c};
test_output[4771:4771] = '{32'hc61a003e};
test_input[38176:38183] = '{32'hc2776358, 32'hc2a4561a, 32'h42797992, 32'hc286cd87, 32'hc1120de7, 32'h41ddc0f6, 32'hc2af8da0, 32'hc217fb55};
test_weights[38176:38183] = '{32'hc234d320, 32'hc2ad33ef, 32'h41865c55, 32'h42c7feda, 32'hc26bfd8b, 32'hc2a09e05, 32'hc1d952a0, 32'h423f4cc4};
test_bias[4772:4772] = '{32'h428823b5};
test_output[4772:4772] = '{32'h4545f204};
test_input[38184:38191] = '{32'h416acd9f, 32'h42a828f9, 32'h412482c9, 32'hc2811964, 32'hc2ba58ad, 32'h42c77869, 32'hc2b3af9c, 32'hc11335e7};
test_weights[38184:38191] = '{32'hc2aa7166, 32'h42b55c80, 32'h421dcd31, 32'h41d09fb0, 32'hc2c6627a, 32'h41fbd7f5, 32'hc2811201, 32'h42569458};
test_bias[4773:4773] = '{32'hbf4b1fac};
test_output[4773:4773] = '{32'h46b1fb14};
test_input[38192:38199] = '{32'hc29dd53a, 32'hc21f3c39, 32'h4270da63, 32'h41b1c29a, 32'h429ceab0, 32'h40251a55, 32'hc18cf7bd, 32'hc1d28b46};
test_weights[38192:38199] = '{32'h411bcc51, 32'hc14fa56b, 32'h414f6a1e, 32'hc20ca8b5, 32'hc2b0fb08, 32'h40fa8341, 32'hc298e465, 32'hc20d2a8f};
test_bias[4774:4774] = '{32'h4298e07e};
test_output[4774:4774] = '{32'hc596b74a};
test_input[38200:38207] = '{32'h428c6acb, 32'h4208eba6, 32'h403a6b28, 32'h42036ceb, 32'h4252d6e8, 32'h42bd5872, 32'hc2a7d94d, 32'hc255e018};
test_weights[38200:38207] = '{32'h428d4d6b, 32'h42b76f54, 32'h41d31d8a, 32'h42b04f62, 32'h426d0363, 32'h41c25226, 32'hc268f770, 32'h4234e3a5};
test_bias[4775:4775] = '{32'h4139a31b};
test_output[4775:4775] = '{32'h46944300};
test_input[38208:38215] = '{32'hc2a6dbe4, 32'h4298e2b0, 32'hc2c07612, 32'hc2a16dc2, 32'h4200bb02, 32'hc082b719, 32'hbfca5eb1, 32'h429e53f3};
test_weights[38208:38215] = '{32'h424259d1, 32'hc2acbd03, 32'hc2917c0e, 32'h413257d8, 32'h4285d80f, 32'hc28c1f22, 32'h4214a3d9, 32'h417081d0};
test_bias[4776:4776] = '{32'h42a891e5};
test_output[4776:4776] = '{32'hc4610ae3};
test_input[38216:38223] = '{32'h4263fcbd, 32'hc1107bed, 32'hc2a36173, 32'hc2b41489, 32'h429683e0, 32'h4127f2aa, 32'hc26151a0, 32'h42c3c40e};
test_weights[38216:38223] = '{32'h41bc6240, 32'hc2b76623, 32'hc29f971e, 32'hc22ba544, 32'hc2be814d, 32'hc266a43d, 32'h4264c0d1, 32'h429d4102};
test_bias[4777:4777] = '{32'h41970e16};
test_output[4777:4777] = '{32'h4610e1dd};
test_input[38224:38231] = '{32'hc1971e04, 32'h42c42f30, 32'hc1bb0a59, 32'hc223838f, 32'h420717dd, 32'hc2b2be0d, 32'hc114d989, 32'h42b343ba};
test_weights[38224:38231] = '{32'h40ce8bd2, 32'hc251d2f1, 32'h40ce4362, 32'hc2acb3bb, 32'hc223cc8d, 32'hc1667c60, 32'hc21aeff6, 32'h41838699};
test_bias[4778:4778] = '{32'h41bdc4f0};
test_output[4778:4778] = '{32'hc2fc494e};
test_input[38232:38239] = '{32'h42b69c51, 32'hc23ae759, 32'hc0e020e5, 32'h413eb6d7, 32'hc289fcb3, 32'hc1d58a75, 32'h42968341, 32'h40debe5e};
test_weights[38232:38239] = '{32'hc1ad9801, 32'h42b6ad6e, 32'h42810b55, 32'hc1cbdf23, 32'hc2b0578c, 32'h426cfa21, 32'hbf93bf84, 32'h4289cedb};
test_bias[4779:4779] = '{32'h4208f4b7};
test_output[4779:4779] = '{32'hc501bf94};
test_input[38240:38247] = '{32'hc1b1c59a, 32'hc1be379d, 32'hc257ff70, 32'hc272159d, 32'hc1e815c6, 32'hc2376cab, 32'h422dc51e, 32'h4201910d};
test_weights[38240:38247] = '{32'h429f3fba, 32'hc25833dc, 32'hc27db5bb, 32'h42879aba, 32'hc279da56, 32'h41f42d30, 32'h41aa2ac7, 32'h422c95d0};
test_bias[4780:4780] = '{32'h41df2b1a};
test_output[4780:4780] = '{32'h44c7ec85};
test_input[38248:38255] = '{32'h41877f88, 32'h42be1f2e, 32'h42be0e71, 32'hc2c0e7f8, 32'hc15b0cd7, 32'hc034722f, 32'hc26c8430, 32'hc153813c};
test_weights[38248:38255] = '{32'h41fd9046, 32'h428e9438, 32'h428264b2, 32'h41c7355d, 32'hc2ad2099, 32'h427ae63d, 32'h4155b7b9, 32'hc2594607};
test_bias[4781:4781] = '{32'h42b557cf};
test_output[4781:4781] = '{32'h463d9a50};
test_input[38256:38263] = '{32'h4281e614, 32'hc2b567d2, 32'h42a018ea, 32'h41dc27e1, 32'h42aba0ef, 32'hc2bbcd45, 32'hc1a0e797, 32'h429fa3fa};
test_weights[38256:38263] = '{32'h42ad5bd0, 32'hc0a8cab5, 32'hc232c02d, 32'h4211bbe1, 32'hc29d86c2, 32'h42588755, 32'hc29cfef2, 32'h4266cafc};
test_bias[4782:4782] = '{32'h4244ea79};
test_output[4782:4782] = '{32'hc501ae03};
test_input[38264:38271] = '{32'h42b9d707, 32'h4266bc17, 32'hc26dccf2, 32'h427cc028, 32'hc17a246a, 32'h429665e4, 32'h4275a90d, 32'h416cd35c};
test_weights[38264:38271] = '{32'h4206dfd6, 32'h41c8349e, 32'h42bea41b, 32'h41b8b1c2, 32'hc27eb511, 32'h421a90af, 32'hc187f388, 32'hc19a1a24};
test_bias[4783:4783] = '{32'hc2b4aa04};
test_output[4783:4783] = '{32'h45322dae};
test_input[38272:38279] = '{32'h426e69e8, 32'h429dd3e4, 32'h41ffc4c4, 32'hc24d15e5, 32'hc23ec479, 32'h420f88e7, 32'hc1a606ee, 32'h42bc6e9e};
test_weights[38272:38279] = '{32'hc2862ac3, 32'hc2985808, 32'hc2949aec, 32'hc1922495, 32'h418d051d, 32'hc2018591, 32'hc26c2250, 32'h4189af5c};
test_bias[4784:4784] = '{32'h4196d1d6};
test_output[4784:4784] = '{32'hc62565c9};
test_input[38280:38287] = '{32'hc1b08f99, 32'hc26c0bf4, 32'h424b16e3, 32'hc292cb6d, 32'hc21e8008, 32'hc28f4188, 32'h4211baf1, 32'h41ea923f};
test_weights[38280:38287] = '{32'h42459ef7, 32'hc1e65376, 32'hc2652e94, 32'hc1f6583f, 32'hc115874c, 32'h424981d3, 32'h420d3862, 32'hc216ce17};
test_bias[4785:4785] = '{32'h428b8a79};
test_output[4785:4785] = '{32'hc53d3c93};
test_input[38288:38295] = '{32'hc22d0e79, 32'hc280462d, 32'h42bf8d2f, 32'hc2be5583, 32'h4208ff62, 32'h41e84adb, 32'h42b6127d, 32'h428a26c9};
test_weights[38288:38295] = '{32'hc2b9b4e2, 32'hc2c7a5ea, 32'h3fa2544f, 32'h412835c6, 32'h427765d0, 32'hc0b05dc5, 32'hc23bebb1, 32'h42aabc4f};
test_bias[4786:4786] = '{32'hc24ee1dd};
test_output[4786:4786] = '{32'h464c2c69};
test_input[38296:38303] = '{32'hc0904380, 32'hc21ccfa4, 32'h4285a798, 32'h42c5f1d0, 32'hc24b3bd4, 32'h422379e8, 32'hc262357a, 32'h41ac842d};
test_weights[38296:38303] = '{32'h4233a36f, 32'hc2ac3954, 32'h42321022, 32'h3ec8c9ca, 32'hc1adc2fd, 32'hc1158d18, 32'hc22bbab3, 32'hc194a037};
test_bias[4787:4787] = '{32'h40e3ddb9};
test_output[4787:4787] = '{32'h460bbc19};
test_input[38304:38311] = '{32'h42666c4f, 32'hc23a4ebc, 32'h4278e05c, 32'h4239e154, 32'h418290a0, 32'hc1db938b, 32'h41bf1e68, 32'hc25563f8};
test_weights[38304:38311] = '{32'hc2aac57e, 32'hc1833f40, 32'h429f04ac, 32'h428d90c3, 32'h421e110f, 32'h414a0057, 32'hc20ea36e, 32'hc082c2e7};
test_bias[4788:4788] = '{32'h4254e15e};
test_output[4788:4788] = '{32'h456d76a3};
test_input[38312:38319] = '{32'h428bc9b5, 32'hc29cc6b0, 32'hc2ac7c2e, 32'h42081c6f, 32'h424495dc, 32'hc1c0160d, 32'h4245e72a, 32'h42969576};
test_weights[38312:38319] = '{32'hc22e49b2, 32'hc2c2ceef, 32'h42b19038, 32'h42c48257, 32'hc2a1bf77, 32'hc2609cf6, 32'h4269a8ab, 32'h412b5128};
test_bias[4789:4789] = '{32'hc24038f8};
test_output[4789:4789] = '{32'h44a24c61};
test_input[38320:38327] = '{32'hc21b6112, 32'hc280f22f, 32'h424a1618, 32'hc242e9f3, 32'h41c79888, 32'hc2c66bac, 32'h42b11f66, 32'hbd7a9f54};
test_weights[38320:38327] = '{32'hc26ce0c0, 32'hc2c07272, 32'h41fac912, 32'hc2b8edc6, 32'h42c4a390, 32'hc2bfda57, 32'hbf00c4ca, 32'h4192277b};
test_bias[4790:4790] = '{32'hc07431c3};
test_output[4790:4790] = '{32'h46cf240e};
test_input[38328:38335] = '{32'hc10c75f9, 32'h4287f2cc, 32'h429ba1db, 32'h3fb9b291, 32'h41c299a1, 32'hc20927b6, 32'h41897e7a, 32'hc283dc95};
test_weights[38328:38335] = '{32'hbeffbaf1, 32'h426f60d7, 32'hc1290782, 32'hc208fedc, 32'h42610528, 32'h42b4b15d, 32'hc0a1b2a4, 32'hc24c36aa};
test_bias[4791:4791] = '{32'h41458260};
test_output[4791:4791] = '{32'h4594d44a};
test_input[38336:38343] = '{32'hc261a068, 32'hc21d6f3f, 32'hc2802a87, 32'h41a66e2b, 32'hc2b892d4, 32'hc18d0e97, 32'hc08bb1fe, 32'hc236dee3};
test_weights[38336:38343] = '{32'hc2b181ea, 32'h42844c48, 32'h42c0895b, 32'hc2a0349f, 32'h42a10f8b, 32'hc2240ee2, 32'h42af2d16, 32'h406a9422};
test_bias[4792:4792] = '{32'h4216d981};
test_output[4792:4792] = '{32'hc645b719};
test_input[38344:38351] = '{32'hc14057bf, 32'h3ee50348, 32'hc298f64b, 32'hc2c60dc2, 32'hc2a7e9ea, 32'h42a803bb, 32'hc21ebdd0, 32'hc220f040};
test_weights[38344:38351] = '{32'h428edb7a, 32'hc172a935, 32'hc2078a81, 32'hc2a25fb6, 32'h4291a2c7, 32'hc2a19a24, 32'hc26611ed, 32'h414319fa};
test_bias[4793:4793] = '{32'h426394b1};
test_output[4793:4793] = '{32'hc4a0d7ec};
test_input[38352:38359] = '{32'hc22e574d, 32'h417a8db6, 32'h424a455e, 32'h42c5dbf7, 32'hc1963b42, 32'h425bc8be, 32'h417b13f3, 32'h425f200d};
test_weights[38352:38359] = '{32'h423c3129, 32'h42142d75, 32'hc29b3d8e, 32'h418df7d6, 32'h42168115, 32'h41f43e47, 32'hc12767f8, 32'hc1b6de90};
test_bias[4794:4794] = '{32'hc25bf832};
test_output[4794:4794] = '{32'hc5821a54};
test_input[38360:38367] = '{32'h42add667, 32'h411ff925, 32'hc2412e4a, 32'hc15492e6, 32'hc1a08d50, 32'hc1a49d3b, 32'hc2890cc0, 32'hc231f0f6};
test_weights[38360:38367] = '{32'hc1ac5d60, 32'h41436242, 32'hc0f64f22, 32'h42c4b45d, 32'h41a62be1, 32'hc2418487, 32'hc2bb6a81, 32'hc1c456ca};
test_bias[4795:4795] = '{32'hc083b240};
test_output[4795:4795] = '{32'h45a8d057};
test_input[38368:38375] = '{32'h41ae95e3, 32'hc2a13d3b, 32'h42b91b33, 32'h41c4e56c, 32'h42b160dc, 32'hc18db2f2, 32'hc27db13c, 32'hc2934ff1};
test_weights[38368:38375] = '{32'hc28ceb43, 32'hc22399c5, 32'h42c3c426, 32'hc2a9c419, 32'h4298faf2, 32'hc1b99155, 32'hc2795726, 32'h42ad8abb};
test_bias[4796:4796] = '{32'h418b0548};
test_output[4796:4796] = '{32'h46530132};
test_input[38376:38383] = '{32'h4285a53c, 32'h427422d4, 32'h4187cf4e, 32'hc1858384, 32'h42c4678e, 32'h4294f69e, 32'hc02093a8, 32'hc2b7f195};
test_weights[38376:38383] = '{32'hbf94ca5f, 32'h415f5b94, 32'h42b83369, 32'h41b353de, 32'hc0eb632a, 32'h42981e67, 32'hc292e0ce, 32'hc2a14267};
test_bias[4797:4797] = '{32'h42c78d67};
test_output[4797:4797] = '{32'h46643883};
test_input[38384:38391] = '{32'h427d0e30, 32'hc28ebb77, 32'h42ae2910, 32'h4259b011, 32'h42b4eb77, 32'hc2933f4d, 32'hc2922356, 32'hc1e442d8};
test_weights[38384:38391] = '{32'h4295e22f, 32'h42599e79, 32'h42c0697b, 32'hc2b4931c, 32'h410b2bcb, 32'h427e1fce, 32'hc2b92da3, 32'hc28a619d};
test_bias[4798:4798] = '{32'hc248810e};
test_output[4798:4798] = '{32'h460e858d};
test_input[38392:38399] = '{32'hc24746e2, 32'hc2b8f220, 32'h412065fe, 32'hc29b4981, 32'h4287cf6e, 32'hc2a81edb, 32'h42466a47, 32'h428a87a5};
test_weights[38392:38399] = '{32'hc28e4b8e, 32'h421bc65c, 32'h4143ade7, 32'h4242ba5c, 32'h4295e6d4, 32'hc138233c, 32'h42c1e532, 32'h42c5f22c};
test_bias[4799:4799] = '{32'h42210838};
test_output[4799:4799] = '{32'h465b7e5b};
test_input[38400:38407] = '{32'h41c79419, 32'hc1279ff6, 32'hc226bf30, 32'h42865d68, 32'hc22ea087, 32'hc24f04a3, 32'h4295a057, 32'hc17f8ca5};
test_weights[38400:38407] = '{32'hc1e192ec, 32'hc20f5701, 32'h421d078d, 32'h40d208d8, 32'h42611d93, 32'h42b2381f, 32'hc1c80a9f, 32'h42bc031d};
test_bias[4800:4800] = '{32'h423dc7f9};
test_output[4800:4800] = '{32'hc63a343e};
test_input[38408:38415] = '{32'hc206ba57, 32'h4259d77e, 32'hc2c73e37, 32'h4250ffd3, 32'h42696ff5, 32'h42b1c48d, 32'h40620d71, 32'hc2acd3ce};
test_weights[38408:38415] = '{32'h423b6313, 32'h42843202, 32'hc1cfe51e, 32'hbe8f7b69, 32'hc29ab05a, 32'hc2beddc8, 32'h42a218a4, 32'hc1e8e077};
test_bias[4801:4801] = '{32'h4248888a};
test_output[4801:4801] = '{32'hc5ad62c2};
test_input[38416:38423] = '{32'h41a72c93, 32'h42b9a49d, 32'hc1a71bf7, 32'hc257eda1, 32'h42090f90, 32'h3fe55a94, 32'h41373aea, 32'hc29c3986};
test_weights[38416:38423] = '{32'hc2a768c5, 32'h42ae7096, 32'hc2929377, 32'hc1b896dc, 32'hc1ff5fd9, 32'hc13a34d3, 32'h416de5fc, 32'hc293e31e};
test_bias[4802:4802] = '{32'h41fb4a4c};
test_output[4802:4802] = '{32'h465a8872};
test_input[38424:38431] = '{32'hc29bf33f, 32'hc2432ac5, 32'hc2695cf4, 32'h42457813, 32'h42418010, 32'hc2c2a4f3, 32'h42a62408, 32'h428a44d9};
test_weights[38424:38431] = '{32'hc2af7223, 32'hc1e130e5, 32'h420099ee, 32'h4293125b, 32'hc2be7cd6, 32'h41a53cfd, 32'h427d3579, 32'h42ab4faf};
test_bias[4803:4803] = '{32'h42533081};
test_output[4803:4803] = '{32'h4663dee6};
test_input[38432:38439] = '{32'h41f70a9e, 32'hc1bf70ac, 32'h4061f6b4, 32'h421d3462, 32'hc115c8d2, 32'h42a2e6e4, 32'hc19408d9, 32'hc2c0c415};
test_weights[38432:38439] = '{32'hc1d3444a, 32'h3f8e9efb, 32'hc2868601, 32'hc2999e03, 32'hc2b24c37, 32'h426788c5, 32'hc28fd8e6, 32'hc211246c};
test_bias[4804:4804] = '{32'hc28a4738};
test_output[4804:4804] = '{32'h45c2100c};
test_input[38440:38447] = '{32'h42909ee8, 32'hc2089fac, 32'hc2890bb0, 32'hc2becc5c, 32'hc25949fe, 32'h42829876, 32'hc28de810, 32'hc27de300};
test_weights[38440:38447] = '{32'h42c3ac3f, 32'h41aaf6db, 32'hc286d17e, 32'hc2bcf9eb, 32'hc28ab44a, 32'hc28f945a, 32'hc138c095, 32'hc19dc38c};
test_bias[4805:4805] = '{32'h42b1662f};
test_output[4805:4805] = '{32'h46a5c24e};
test_input[38448:38455] = '{32'hc2af1879, 32'h4145a1d1, 32'h421be106, 32'h4288f494, 32'h421fbb0c, 32'hc284addb, 32'hc2ab054f, 32'hc286d172};
test_weights[38448:38455] = '{32'hc2a64229, 32'hc1b99b76, 32'h426c887d, 32'h429752d0, 32'h42b6f1bd, 32'hc1fbeef7, 32'hc189a9a4, 32'h428bfc34};
test_bias[4806:4806] = '{32'hc21aeafc};
test_output[4806:4806] = '{32'h46844a6a};
test_input[38456:38463] = '{32'hc23e1502, 32'hc29afe85, 32'h41e8454b, 32'h42099a10, 32'hc23e6a0f, 32'h42772145, 32'hc2ac6b1c, 32'h426dcd1f};
test_weights[38456:38463] = '{32'hc13a1c2f, 32'hc2040e67, 32'hc1e93a01, 32'hc0f42e33, 32'h427716cd, 32'hc2934352, 32'hc1ac458f, 32'h42ab6400};
test_bias[4807:4807] = '{32'hc2a96971};
test_output[4807:4807] = '{32'h44ac5ddc};
test_input[38464:38471] = '{32'h4256271e, 32'hc1940c05, 32'h42c5fe3f, 32'hc253aef3, 32'h42be22a6, 32'hc20d4060, 32'h41d0b8ff, 32'hc1d08903};
test_weights[38464:38471] = '{32'h429ce1de, 32'h4192962a, 32'hc04445db, 32'hc2a0ab8a, 32'hc252cb44, 32'hc16dfe79, 32'hc1cfb854, 32'hc2aef662};
test_bias[4808:4808] = '{32'h42b7251e};
test_output[4808:4808] = '{32'h459cd135};
test_input[38472:38479] = '{32'hc2b9d8ab, 32'hc295cc1e, 32'hc20a5d1f, 32'h4234edc6, 32'h3ff66e3b, 32'hc23ba440, 32'h4211fd4f, 32'h428fa677};
test_weights[38472:38479] = '{32'hc21a29af, 32'h417eb079, 32'h425681dd, 32'hc0238bc9, 32'hc1a53bf8, 32'hc2bf1204, 32'h42777503, 32'h429cd5e7};
test_bias[4809:4809] = '{32'hc1db215d};
test_output[4809:4809] = '{32'h4646ccba};
test_input[38480:38487] = '{32'h4298506e, 32'h423e4e06, 32'h42be6ab7, 32'hc0039f86, 32'hc24be771, 32'hc2c63782, 32'h413b583e, 32'hc201c00a};
test_weights[38480:38487] = '{32'hc299f0a9, 32'hc29bd0ed, 32'hc1bd1f62, 32'hc2a0f6ba, 32'h42a4dcfd, 32'hc2768b57, 32'h429fbc78, 32'h425a84c5};
test_bias[4810:4810] = '{32'h42b9c9b5};
test_output[4810:4810] = '{32'hc623ebee};
test_input[38488:38495] = '{32'h429124f0, 32'hc2a8a398, 32'h41a6a868, 32'h414463c3, 32'hc0fd5448, 32'hc1029f53, 32'h41e54f75, 32'h426bc134};
test_weights[38488:38495] = '{32'hc238ff3b, 32'hc28a6819, 32'hc2a244d6, 32'h42af499e, 32'h4291d469, 32'hc2a403e5, 32'hc29862e3, 32'hc1bb5da0};
test_bias[4811:4811] = '{32'h42346019};
test_output[4811:4811] = '{32'hc4c3554c};
test_input[38496:38503] = '{32'h429fbe79, 32'hc29967c1, 32'hc29ec935, 32'h41f843b6, 32'h41b70684, 32'hc0066bb0, 32'h424e9bbf, 32'hc222d566};
test_weights[38496:38503] = '{32'hc2acb327, 32'hc227232c, 32'h42b92a6a, 32'h41c0a010, 32'h42583f9a, 32'h42c41efa, 32'h42482cbb, 32'hc2a9e8b6};
test_bias[4812:4812] = '{32'h42be0942};
test_output[4812:4812] = '{32'hc54360e3};
test_input[38504:38511] = '{32'hc20a6302, 32'hc2100e03, 32'hc2b2a8ee, 32'h41ce527a, 32'hc2b2f2b9, 32'hbfe1df9f, 32'h428c8333, 32'hc28bfbdb};
test_weights[38504:38511] = '{32'hc2235ee0, 32'h4229d224, 32'hc22fe0a3, 32'hc2b6b84e, 32'h423f5c42, 32'hc214da74, 32'hc232b5c3, 32'h42560727};
test_bias[4813:4813] = '{32'h421b62cb};
test_output[4813:4813] = '{32'hc61610ea};
test_input[38512:38519] = '{32'hc296cbd6, 32'hc207c054, 32'h429b1971, 32'hc0976588, 32'h42a97d3a, 32'h40ef96f9, 32'h4230e7b9, 32'h42c284d3};
test_weights[38512:38519] = '{32'hc2a66a48, 32'hc1e89be9, 32'hc1e1112d, 32'h4196257f, 32'hbf444a53, 32'h41b61271, 32'hc2a34487, 32'h4259505c};
test_bias[4814:4814] = '{32'h41ca9719};
test_output[4814:4814] = '{32'h45d45246};
test_input[38520:38527] = '{32'hc2ba004a, 32'h4208bcd1, 32'h42849700, 32'h42a132e3, 32'hc29b2af9, 32'h413b34df, 32'h420319ea, 32'hc290d215};
test_weights[38520:38527] = '{32'hc1fdafa6, 32'h42bb12c8, 32'hc2438380, 32'h42c1a6a2, 32'h4287b797, 32'h42976ddb, 32'hc2aff216, 32'hc29a2e46};
test_bias[4815:4815] = '{32'h42c42a15};
test_output[4815:4815] = '{32'h460ea158};
test_input[38528:38535] = '{32'h40b33587, 32'h4167bdf2, 32'hc294c582, 32'h42adb544, 32'h42226e7b, 32'hbfd65b41, 32'h42936210, 32'h41569ad4};
test_weights[38528:38535] = '{32'hc2745b67, 32'hc20ed27e, 32'h42351b50, 32'hc213b493, 32'h41701cfd, 32'hc2455cb7, 32'hc0c744a3, 32'h42208cb5};
test_bias[4816:4816] = '{32'hc12daa4e};
test_output[4816:4816] = '{32'hc5d08e1e};
test_input[38536:38543] = '{32'h41891261, 32'h42b6827d, 32'h4214f15e, 32'h42732457, 32'h419dae77, 32'hc1b62cd7, 32'h4293ba18, 32'hc21c4aca};
test_weights[38536:38543] = '{32'h4290b0e3, 32'hc08618f8, 32'h426a6eae, 32'h41b890f4, 32'hc2adb651, 32'hc29ba14a, 32'hbf220623, 32'hc25137d8};
test_bias[4817:4817] = '{32'h427141c2};
test_output[4817:4817] = '{32'h45ccf92f};
test_input[38544:38551] = '{32'hc0ed11f9, 32'h42a72aee, 32'hc205594e, 32'h40f4b9d8, 32'h4298627e, 32'hc2b6a533, 32'hc2573865, 32'h42b39262};
test_weights[38544:38551] = '{32'hc2c1a60e, 32'hc0d29412, 32'hc2c03a37, 32'h40aa5fd4, 32'hc25a0262, 32'hc2476ff4, 32'hc1f4514c, 32'hc24ee38b};
test_bias[4818:4818] = '{32'hc0ad45b2};
test_output[4818:4818] = '{32'h4449a939};
test_input[38552:38559] = '{32'hc2688f71, 32'h4199beb4, 32'hc19c3862, 32'h42a0a458, 32'hc29af750, 32'h4263c5d2, 32'h416da34f, 32'hc17cad3c};
test_weights[38552:38559] = '{32'h428bf45e, 32'hc13005b8, 32'h4243ab1d, 32'hc2048f0a, 32'hc2ba8d02, 32'h42c25802, 32'hc232385c, 32'h42861e5d};
test_bias[4819:4819] = '{32'h4249eafa};
test_output[4819:4819] = '{32'h454794bf};
test_input[38560:38567] = '{32'h41fd5a22, 32'h428a4a17, 32'h3f34e255, 32'hc158bbf0, 32'h42867915, 32'h40605216, 32'h42a87007, 32'hc2275139};
test_weights[38560:38567] = '{32'h3d73c3dd, 32'hc2ab661b, 32'hc28cd47a, 32'h4281c13e, 32'h4286e80f, 32'hc24c827a, 32'h429cad0b, 32'h42aa6607};
test_bias[4820:4820] = '{32'h42a1638e};
test_output[4820:4820] = '{32'h441a8a59};
test_input[38568:38575] = '{32'hc248ec00, 32'hc291643f, 32'h412f15e8, 32'hc20db356, 32'hc2ac87bb, 32'h42bd347c, 32'hc2832298, 32'hc28e028f};
test_weights[38568:38575] = '{32'hc1a85675, 32'hc16bb96e, 32'h41da6330, 32'h42649b01, 32'hc22780cf, 32'h41e16478, 32'hc27c5456, 32'hc2bb9089};
test_bias[4821:4821] = '{32'h404ba244};
test_output[4821:4821] = '{32'h46888c69};
test_input[38576:38583] = '{32'h429c7bc2, 32'hc15c9762, 32'h41c36c3c, 32'hc29b6d89, 32'h422896e1, 32'hc2382746, 32'hc28925b7, 32'h4280c85c};
test_weights[38576:38583] = '{32'hc156bb0b, 32'hc27ee8a5, 32'h429cf102, 32'hc1767020, 32'h42774b1f, 32'hc22c651f, 32'hc2c19d1b, 32'hc28ca232};
test_bias[4822:4822] = '{32'hc22a4acd};
test_output[4822:4822] = '{32'h46160147};
test_input[38584:38591] = '{32'hc29a7b77, 32'hc26b9368, 32'h42bceef7, 32'hc24e3c3a, 32'h4231c0c8, 32'hc2487f39, 32'hc1f480d6, 32'h428c076b};
test_weights[38584:38591] = '{32'h4265e849, 32'h42b0b03b, 32'h4291382d, 32'h42681826, 32'hc1ef1389, 32'hc1c06594, 32'h42810388, 32'hc26d10bc};
test_bias[4823:4823] = '{32'hc237d125};
test_output[4823:4823] = '{32'hc63c81dd};
test_input[38592:38599] = '{32'h41fdf72f, 32'hc1d744ac, 32'hc286c8da, 32'hc2a0ba9e, 32'hc294e440, 32'h4253bb2a, 32'h428513b7, 32'h421efd1e};
test_weights[38592:38599] = '{32'hc28f3357, 32'hc29196ca, 32'hc078cda0, 32'hc21331dd, 32'h4280a448, 32'hc2493ff8, 32'hc2b9a68c, 32'h42aa0926};
test_bias[4824:4824] = '{32'hc279b962};
test_output[4824:4824] = '{32'hc5e7715d};
test_input[38600:38607] = '{32'hc1ccf4d0, 32'hc1c352e3, 32'hc243f7a7, 32'hc1c6adea, 32'hc2283c4b, 32'hc23390d5, 32'hc15e9231, 32'hc298fa31};
test_weights[38600:38607] = '{32'h42a9c399, 32'h42413a22, 32'h41acaf21, 32'h414f8b9b, 32'hc2496377, 32'hc1beb1dd, 32'hc1eb2dc4, 32'hc2809659};
test_bias[4825:4825] = '{32'hc2b602f6};
test_output[4825:4825] = '{32'h456698c3};
test_input[38608:38615] = '{32'hc28c145e, 32'hc1aeb61c, 32'h412e0de9, 32'hc28706a2, 32'hc1ef8d47, 32'h41a039e9, 32'h4273243b, 32'h41f5c5c3};
test_weights[38608:38615] = '{32'h41753bd3, 32'hc2bbe0a4, 32'hc2144392, 32'hc063b89c, 32'h4184dd35, 32'hc198fadc, 32'h424b99a8, 32'hc1fec094};
test_bias[4826:4826] = '{32'hc28c77d1};
test_output[4826:4826] = '{32'h44f78531};
test_input[38616:38623] = '{32'hc2639586, 32'h428a1a5a, 32'h4232d811, 32'h41467bd5, 32'h42a4f476, 32'h4295e419, 32'hc26f40e7, 32'h429893d8};
test_weights[38616:38623] = '{32'h41d13bb1, 32'h42211fab, 32'h4183204b, 32'h4214f872, 32'hc24d808c, 32'h4209a5bd, 32'h40b4f4d4, 32'hc2839214};
test_bias[4827:4827] = '{32'h4278443b};
test_output[4827:4827] = '{32'hc58b875c};
test_input[38624:38631] = '{32'h42559f98, 32'hc28a415b, 32'hc2c5cf46, 32'h40ce1f54, 32'h428b5109, 32'h41828091, 32'h42b5a74e, 32'h41c9f1cb};
test_weights[38624:38631] = '{32'h4120646a, 32'hc2625062, 32'h41c6d4a5, 32'hc1f9be97, 32'h42001b09, 32'h42ae5210, 32'h42b71780, 32'hc18790d1};
test_bias[4828:4828] = '{32'hc2215198};
test_output[4828:4828] = '{32'h464f9ada};
test_input[38632:38639] = '{32'hc1ac96ca, 32'hc2b7ecaf, 32'h41c56762, 32'h4294158e, 32'h4161f5bd, 32'hc237640f, 32'h42c00ce7, 32'hc2c75b2e};
test_weights[38632:38639] = '{32'h40b3d6b1, 32'h41c4fca6, 32'h41f7b376, 32'h429aa5b4, 32'hc22d9e51, 32'hc2a29a8e, 32'h40a2fed0, 32'h4222f1f5};
test_bias[4829:4829] = '{32'h42a96c99};
test_output[4829:4829] = '{32'h4569364d};
test_input[38640:38647] = '{32'h422919b1, 32'h41731f1f, 32'hc2858999, 32'hc2bda370, 32'hc2314e91, 32'h41c4eed6, 32'h41efeb88, 32'hc2c1526e};
test_weights[38640:38647] = '{32'h425a114d, 32'h428171e6, 32'h42aa74f8, 32'hbda0fd48, 32'h42801903, 32'hc20e9193, 32'h420c5c84, 32'hc2c3e34e};
test_bias[4830:4830] = '{32'hc29d57c8};
test_output[4830:4830] = '{32'h45874ce3};
test_input[38648:38655] = '{32'h41a76f1f, 32'h41115dc7, 32'h423bb8a1, 32'h429bd89c, 32'h424efb34, 32'hc18ca1d7, 32'hc1cac756, 32'h428c2256};
test_weights[38648:38655] = '{32'h42c1b1f3, 32'hc2516f21, 32'hc18f8d9a, 32'hc2b33f61, 32'hc2a7a159, 32'h3f8c1ba1, 32'h4212d32f, 32'h42b1fa0d};
test_bias[4831:4831] = '{32'hc22df9e3};
test_output[4831:4831] = '{32'hc5a7cd4b};
test_input[38656:38663] = '{32'h428006a8, 32'h42531cc7, 32'hc2a1792a, 32'hc2ace5a7, 32'hc2bcda0c, 32'hc15f2fa0, 32'hc291c032, 32'h41a0a32d};
test_weights[38656:38663] = '{32'h421144d2, 32'hc2608237, 32'h419603ef, 32'hc23cbaad, 32'h4224764e, 32'h41ef1470, 32'h40ace27b, 32'h429009ff};
test_bias[4832:4832] = '{32'hc21a84d0};
test_output[4832:4832] = '{32'hc4a9c325};
test_input[38664:38671] = '{32'h428089e6, 32'h42a5dc1a, 32'h41b81f50, 32'h428691ef, 32'h42baeb11, 32'hc217ce68, 32'h429d1127, 32'h423e7d26};
test_weights[38664:38671] = '{32'h4218544e, 32'hc18a9a50, 32'hc25bd89d, 32'h40c776d4, 32'h410cf415, 32'h42b5dbee, 32'h42778e97, 32'hc2c160b6};
test_bias[4833:4833] = '{32'h428ff403};
test_output[4833:4833] = '{32'hc5056946};
test_input[38672:38679] = '{32'hc2c4b1e6, 32'h4163efbc, 32'hc294f6a4, 32'hc2308db4, 32'hc27a8685, 32'hc2523f43, 32'hc23298b9, 32'h4233f608};
test_weights[38672:38679] = '{32'hc2c5fafb, 32'h42c36a59, 32'hc21749a4, 32'h4255cb9f, 32'hc2781bad, 32'h418e8556, 32'h4143a443, 32'hc2a2ac2f};
test_bias[4834:4834] = '{32'h41282360};
test_output[4834:4834] = '{32'h46218bbe};
test_input[38680:38687] = '{32'hc229327f, 32'h418a0b94, 32'h4284014e, 32'h429b6f98, 32'h42230472, 32'h42800b9d, 32'h3fc01043, 32'hc2af18c3};
test_weights[38680:38687] = '{32'hc1fef04e, 32'h42a33b5d, 32'h414ba287, 32'h429d9b55, 32'h4287f0a9, 32'hc288995c, 32'h425ff2b4, 32'h424048d5};
test_bias[4835:4835] = '{32'h42bc50c5};
test_output[4835:4835] = '{32'h457f7bd9};
test_input[38688:38695] = '{32'hc29e99c0, 32'hc1c12334, 32'h425fc8a5, 32'h429279a1, 32'hc187c2d2, 32'h42480587, 32'hc29c3088, 32'hc1f948e9};
test_weights[38688:38695] = '{32'hc2589482, 32'h42b875a2, 32'h404ec779, 32'hc2b3fa04, 32'hc26bcc45, 32'h42b670ba, 32'h429c8230, 32'hc28d3c61};
test_bias[4836:4836] = '{32'hc290cfad};
test_output[4836:4836] = '{32'hc52cbf4f};
test_input[38696:38703] = '{32'hc1acd55b, 32'h41106cd5, 32'hc1dffe6d, 32'h421b04fe, 32'hc272bb15, 32'hc2a9b011, 32'hc1249c1e, 32'h427bb216};
test_weights[38696:38703] = '{32'hc2ba8d74, 32'h41ea8cbd, 32'hc2b30047, 32'h4222ea7b, 32'hc1d2ff72, 32'h3fbf096e, 32'hc12f2170, 32'hc280a243};
test_bias[4837:4837] = '{32'hc2a4a489};
test_output[4837:4837] = '{32'h456ed46e};
test_input[38704:38711] = '{32'hc18db5d5, 32'hc006a19c, 32'hc2b9470b, 32'hc0093a1f, 32'hc2077b18, 32'hc293d034, 32'h421beabf, 32'hc21e2744};
test_weights[38704:38711] = '{32'h42931bf4, 32'h4228b598, 32'h429351a3, 32'h409a6181, 32'h42abea5f, 32'hc12bfc6c, 32'h42c76410, 32'hc2b75532};
test_bias[4838:4838] = '{32'h4212a45f};
test_output[4838:4838] = '{32'hc52eba49};
test_input[38712:38719] = '{32'hc22d0bd5, 32'h428f0739, 32'h428309e6, 32'h3f3e6c49, 32'h42284c8c, 32'hc2315062, 32'hc227df37, 32'h42c654fa};
test_weights[38712:38719] = '{32'hc2642aa3, 32'h42abe41b, 32'h4288f748, 32'h428b4347, 32'h42c6e42c, 32'h4276d692, 32'hc2847123, 32'h42093bdd};
test_bias[4839:4839] = '{32'hc29d1f81};
test_output[4839:4839] = '{32'h46a1c08b};
test_input[38720:38727] = '{32'hc1a7922a, 32'hc2582494, 32'hc234cea8, 32'h410a9f72, 32'hc1e05e96, 32'h4293a808, 32'hc20269ff, 32'h4291fcb6};
test_weights[38720:38727] = '{32'hc167e65f, 32'h4211861f, 32'hc2665a55, 32'h422bed51, 32'h429a940c, 32'hc090606f, 32'hc208f7dc, 32'hc24be5f4};
test_bias[4840:4840] = '{32'hc27f936b};
test_output[4840:4840] = '{32'hc570fdbe};
test_input[38728:38735] = '{32'hc1e2efcf, 32'hbf89bf35, 32'h40894b5d, 32'h410820db, 32'h4267e8bd, 32'h41fc466d, 32'hc23ffac4, 32'h415b3bc2};
test_weights[38728:38735] = '{32'h426e0482, 32'hc23e93a0, 32'h428805c8, 32'h42c7fbec, 32'h4245dce2, 32'hc2a74747, 32'h42802d34, 32'hc19d8b52};
test_bias[4841:4841] = '{32'h4297a7a3};
test_output[4841:4841] = '{32'hc55cdb43};
test_input[38736:38743] = '{32'h429be9c0, 32'hc18234e0, 32'hc0e150a7, 32'h428eb374, 32'hc2072455, 32'hc27905c8, 32'hc087f14d, 32'hc00a656a};
test_weights[38736:38743] = '{32'h4289c0bb, 32'hc2b3bff8, 32'hbfa54b04, 32'hc1d15dd2, 32'h424f54f5, 32'h419f6f5a, 32'hc1dd12da, 32'h428c2b3e};
test_bias[4842:4842] = '{32'h42a57952};
test_output[4842:4842] = '{32'h44fdd388};
test_input[38744:38751] = '{32'hc2b78421, 32'hc1aa6814, 32'h42664989, 32'h4234dc8e, 32'h42ae0427, 32'hc189ba8b, 32'h421451ab, 32'hc24f5175};
test_weights[38744:38751] = '{32'hc2a8b76a, 32'h4201a9c6, 32'h4235daa3, 32'h41dcff40, 32'hc2665935, 32'hc24680a3, 32'h4148e15e, 32'h42c712f2};
test_bias[4843:4843] = '{32'hc2bdc0b2};
test_output[4843:4843] = '{32'h44f681cc};
test_input[38752:38759] = '{32'hc241c63d, 32'hc29ba0e6, 32'hc1f9d6a0, 32'h418d2388, 32'hc2672f9c, 32'h42ac06e3, 32'h412a8d4b, 32'h427e5a10};
test_weights[38752:38759] = '{32'h40f45359, 32'hc22ab6f0, 32'h422fd984, 32'h41c84b3f, 32'hc263f7d8, 32'h4282e30f, 32'hc18a2e44, 32'h428a8359};
test_bias[4844:4844] = '{32'h42532ae9};
test_output[4844:4844] = '{32'h466dbdab};
test_input[38760:38767] = '{32'hc2be0674, 32'hc272558d, 32'h425af7c6, 32'h42c7547e, 32'h4177dcdf, 32'hc29e776c, 32'h408b2756, 32'hc29f4e3d};
test_weights[38760:38767] = '{32'h42bc8ab3, 32'h41945b77, 32'h41f21cc2, 32'hc27a559d, 32'hc2a12f6e, 32'h426c4b25, 32'h42817c96, 32'hc25d06fc};
test_bias[4845:4845] = '{32'h3da6f1cf};
test_output[4845:4845] = '{32'hc6788cc9};
test_input[38768:38775] = '{32'hc20c9c88, 32'hc2c2db51, 32'h40bff9ad, 32'hc2bca586, 32'h421563d1, 32'hc2248923, 32'hc25fd351, 32'hc10872d6};
test_weights[38768:38775] = '{32'h42223215, 32'h41ac8288, 32'h42a9d4ec, 32'h42c761ff, 32'hc2964c23, 32'h41831d93, 32'hc28bfeb8, 32'hc06cf5c7};
test_bias[4846:4846] = '{32'h40891cfb};
test_output[4846:4846] = '{32'hc63ab0ed};
test_input[38776:38783] = '{32'hc285f2e4, 32'hc2bd5935, 32'h4237217d, 32'h422305a7, 32'hc1d6ed42, 32'h426f2fa8, 32'hc1413300, 32'hc1932f02};
test_weights[38776:38783] = '{32'h41f6cffc, 32'hc28b72f5, 32'hc2a862ca, 32'h42b60d49, 32'h4187daeb, 32'hc2903fff, 32'h4151c4ed, 32'h4287119b};
test_bias[4847:4847] = '{32'h4206c4ff};
test_output[4847:4847] = '{32'hc4da42d6};
test_input[38784:38791] = '{32'hc2c26c38, 32'h42a8c026, 32'h426e1f4d, 32'hc0a98ca0, 32'hc2acc341, 32'h4127cb79, 32'h41947707, 32'h41324a8d};
test_weights[38784:38791] = '{32'hc29e8726, 32'h42a05dba, 32'hc2761b86, 32'h3ecdac07, 32'h41445b8f, 32'hc1c4a3e4, 32'h42bd6196, 32'h41954cb8};
test_bias[4848:4848] = '{32'hc1ba4523};
test_output[4848:4848] = '{32'h4632982f};
test_input[38792:38799] = '{32'h423e6719, 32'h41c0d640, 32'h42c76773, 32'hc29466c5, 32'h4297a8ad, 32'hc2a2b5c2, 32'hc28381c4, 32'hc2a4c70d};
test_weights[38792:38799] = '{32'h426ed266, 32'h42b4e01e, 32'h42738f6a, 32'hc245db22, 32'h4053eb89, 32'h42bdd63f, 32'h42ad54ae, 32'hc1c9997f};
test_bias[4849:4849] = '{32'h4269460c};
test_output[4849:4849] = '{32'h4569013d};
test_input[38800:38807] = '{32'h42587cde, 32'hc2b7c1db, 32'h42b2edb0, 32'hc1fb2218, 32'h41f8ea5a, 32'hc2874763, 32'hc1f9836b, 32'h4269a43f};
test_weights[38800:38807] = '{32'h4270a1a9, 32'hc2af5208, 32'h42c560b6, 32'h42c40a69, 32'h4288a651, 32'h42b7ee34, 32'hc26b3851, 32'hc28048dc};
test_bias[4850:4850] = '{32'hc25cb4ee};
test_output[4850:4850] = '{32'h462bdf38};
test_input[38808:38815] = '{32'hc2a57920, 32'hc12dd42e, 32'h420775d4, 32'h4277cbd0, 32'h428871bc, 32'h41f88e9b, 32'hc1b0ede2, 32'hc1b4c5c0};
test_weights[38808:38815] = '{32'hc2ba7423, 32'hc29d5570, 32'h40b16780, 32'hc29d1486, 32'hc2c0986e, 32'h417b7870, 32'h429b5782, 32'h413d4e2e};
test_bias[4851:4851] = '{32'h4297b349};
test_output[4851:4851] = '{32'hc580234c};
test_input[38816:38823] = '{32'h42506da6, 32'h42ad6582, 32'h42871051, 32'hc1825d35, 32'hc1faca21, 32'hc11a8525, 32'hc2864ca4, 32'hc1ef26f0};
test_weights[38816:38823] = '{32'h42c6d4be, 32'h419e285b, 32'h42295353, 32'hc299b92b, 32'h425caaa2, 32'hc23e9347, 32'h41efe8a0, 32'h42c20b56};
test_bias[4852:4852] = '{32'hc282424e};
test_output[4852:4852] = '{32'h4594a79b};
test_input[38824:38831] = '{32'h42c5ee75, 32'h41467726, 32'h4102266a, 32'h42b9d5df, 32'h41c84aed, 32'h4159f454, 32'hc2622c1b, 32'h408def0f};
test_weights[38824:38831] = '{32'h42270a6e, 32'hc065bb30, 32'h42887822, 32'hc2244d11, 32'hc2bc7fe7, 32'h42a1ef9d, 32'hc22d9042, 32'h42c088ab};
test_bias[4853:4853] = '{32'hc26e50c9};
test_output[4853:4853] = '{32'h45156daa};
test_input[38832:38839] = '{32'h428b3ad8, 32'hc212c130, 32'hc1b3a19a, 32'h411c5d5c, 32'hc25b67e7, 32'h418c0ea9, 32'hc24da2a3, 32'h41c61dc0};
test_weights[38832:38839] = '{32'h41744d66, 32'hc2524512, 32'h42b0a5a2, 32'hc203bf21, 32'h429a5658, 32'hc00c7642, 32'h409bd615, 32'h420a5293};
test_bias[4854:4854] = '{32'h41ed181e};
test_output[4854:4854] = '{32'hc5385199};
test_input[38840:38847] = '{32'h42200baa, 32'hc113536c, 32'hc2c6e34a, 32'h41c3b17d, 32'hc2aa3a9b, 32'h42b4899f, 32'h429b64b1, 32'h41d47f0a};
test_weights[38840:38847] = '{32'h41ec8942, 32'hc24dd2f6, 32'hc2abc43f, 32'h425b4dc8, 32'hc2094702, 32'hc2c4c00d, 32'h42b711c1, 32'hc299047d};
test_bias[4855:4855] = '{32'h4240793e};
test_output[4855:4855] = '{32'h46274ce5};
test_input[38848:38855] = '{32'hc2878a7f, 32'hc0f94ef3, 32'h4238766e, 32'hc28e5a78, 32'hc2bbbc4e, 32'h42726180, 32'h4272c120, 32'hc20a25c0};
test_weights[38848:38855] = '{32'hc2aa12e4, 32'hc2819a3d, 32'hc294f480, 32'hc2c2c3f5, 32'hc18d96fd, 32'hc283c8af, 32'hc285f752, 32'h4164a163};
test_bias[4856:4856] = '{32'h42a4fc20};
test_output[4856:4856] = '{32'h4538d213};
test_input[38856:38863] = '{32'hc26fbb13, 32'hc2504070, 32'h4289440d, 32'h41a4d86e, 32'h428b3a34, 32'hc15e197c, 32'hc0462f7b, 32'h429cdcab};
test_weights[38856:38863] = '{32'h42af75b2, 32'h410fa4bb, 32'hc0b49cad, 32'h425f465c, 32'hc2c6be74, 32'h42886054, 32'h4240a491, 32'hc1f59cd5};
test_bias[4857:4857] = '{32'hc2101fa8};
test_output[4857:4857] = '{32'hc670ef29};
test_input[38864:38871] = '{32'hc2706206, 32'h42c0d5d6, 32'hc0542eeb, 32'h42c058ee, 32'hc09db649, 32'h42c239a1, 32'h41010c4c, 32'hc2a157ed};
test_weights[38864:38871] = '{32'hc25ba8ed, 32'h4266d95e, 32'hc09abd88, 32'h4299104b, 32'h4262e111, 32'hc1b4adb7, 32'hc285e896, 32'h421619ca};
test_bias[4858:4858] = '{32'hc283a06f};
test_output[4858:4858] = '{32'h461e5c97};
test_input[38872:38879] = '{32'hc2aa4472, 32'hc25435a8, 32'hc291829e, 32'hc2453377, 32'hc26cb2e2, 32'h42bca90d, 32'hc266d57f, 32'h4199babb};
test_weights[38872:38879] = '{32'h424713a9, 32'hc29fbcef, 32'h41d8e467, 32'h42900bc7, 32'hc201f3d6, 32'hc22de708, 32'hc2a60482, 32'h425984d4};
test_bias[4859:4859] = '{32'h4256d0e9};
test_output[4859:4859] = '{32'hc4e294be};
test_input[38880:38887] = '{32'h41c92bd4, 32'h4282ce9d, 32'h424e29d1, 32'hc1c1f96e, 32'h42713271, 32'h42932a9c, 32'h4293b272, 32'h42c54028};
test_weights[38880:38887] = '{32'hc2c6f5e4, 32'h41863092, 32'hc2936abe, 32'hc2b80344, 32'hc1a3ec59, 32'h42800b61, 32'h41bfb245, 32'hc2a69c32};
test_bias[4860:4860] = '{32'hc1c6a0de};
test_output[4860:4860] = '{32'hc5ba83f9};
test_input[38888:38895] = '{32'h421383ae, 32'h42aca33f, 32'hc14d9328, 32'h42c6bad7, 32'hc20cf8dd, 32'h4224b7c3, 32'hc26da9cc, 32'hc289e012};
test_weights[38888:38895] = '{32'hc1d5abbd, 32'hc254b246, 32'hc1bf8661, 32'h424b7b73, 32'h4278e135, 32'hc2b14c96, 32'hc289b0b5, 32'h42739a7f};
test_bias[4861:4861] = '{32'h416ba1e3};
test_output[4861:4861] = '{32'hc5c0288e};
test_input[38896:38903] = '{32'hc1dbf709, 32'hc21fdc08, 32'hc12e3045, 32'hc2c67631, 32'h421e35bc, 32'hc26cbd1b, 32'h4093bafc, 32'h41fd3c32};
test_weights[38896:38903] = '{32'hc2a3159e, 32'h4284b7d2, 32'hc2af9c04, 32'h41395f14, 32'hc2355f0f, 32'h4286773e, 32'h41ba9617, 32'h40d40c32};
test_bias[4862:4862] = '{32'h40e36c61};
test_output[4862:4862] = '{32'hc5bd1e1e};
test_input[38904:38911] = '{32'h40fc7353, 32'h41ff3e1d, 32'hc222ffc3, 32'h426c218e, 32'h41d7bfd2, 32'hc22f3f54, 32'hc21197d1, 32'hc2c17d71};
test_weights[38904:38911] = '{32'h4288eeb2, 32'h42aedb84, 32'h40a31550, 32'h41d0084a, 32'h42a157be, 32'h4235833e, 32'hc1e97e9e, 32'hc12ecf98};
test_bias[4863:4863] = '{32'h42420ce8};
test_output[4863:4863] = '{32'h45db22df};
test_input[38912:38919] = '{32'hc285ee70, 32'hc2809019, 32'hc090c526, 32'h42729259, 32'h428bd8c9, 32'hc2a28127, 32'h41ce9e3a, 32'h41f66023};
test_weights[38912:38919] = '{32'h4245e60f, 32'hc26a597a, 32'h417fb87a, 32'hc110e26d, 32'hc2151776, 32'h427e1e37, 32'h42aa6820, 32'hc2292228};
test_bias[4864:4864] = '{32'h41b584fb};
test_output[4864:4864] = '{32'hc5db3c94};
test_input[38920:38927] = '{32'h3fe8bbd2, 32'h42a52e3b, 32'h425ea095, 32'h42c45d20, 32'hc276a5e8, 32'hc1961e2d, 32'h423d674f, 32'h4195eb32};
test_weights[38920:38927] = '{32'hc2a1589c, 32'h40ad2a3d, 32'h428b2641, 32'hc215bbf4, 32'h41fa34c6, 32'hc2ac098f, 32'h41f469d0, 32'hc13d5e9f};
test_bias[4865:4865] = '{32'hc28e5077};
test_output[4865:4865] = '{32'h44a7115d};
test_input[38928:38935] = '{32'hc1953103, 32'hc27c8bdf, 32'h42b23324, 32'hc22178bf, 32'hc2ae0624, 32'hc2b35ac1, 32'hc2c16893, 32'h423884ca};
test_weights[38928:38935] = '{32'hc2246404, 32'hc239acf8, 32'hc197989c, 32'hc1139b86, 32'h42368939, 32'h41b7d8e6, 32'hc109e56d, 32'h426e503c};
test_bias[4866:4866] = '{32'h41c6bbdf};
test_output[4866:4866] = '{32'hc22f1de8};
test_input[38936:38943] = '{32'hc2126aff, 32'h40ab981c, 32'hc261ac0b, 32'hc24206a7, 32'h42b502d6, 32'hc2082d06, 32'h42b7a188, 32'hc2899f4b};
test_weights[38936:38943] = '{32'hc1f1d067, 32'h4134223f, 32'hc21c3625, 32'h411136b5, 32'h424d3937, 32'hc2197095, 32'hc2a37d82, 32'hc2834e0e};
test_bias[4867:4867] = '{32'h41989471};
test_output[4867:4867] = '{32'h45b8b3ba};
test_input[38944:38951] = '{32'h42667fb1, 32'h4299f38b, 32'hc2a7a07c, 32'h42af33b6, 32'h427091cc, 32'h41b69619, 32'hc1bb98de, 32'hc230c18f};
test_weights[38944:38951] = '{32'h425af1a3, 32'h42509895, 32'hc259bb80, 32'h42672fff, 32'hc1311bf6, 32'h428c1fac, 32'hc203051a, 32'h42ac29be};
test_bias[4868:4868] = '{32'h42173f83};
test_output[4868:4868] = '{32'h466623f7};
test_input[38952:38959] = '{32'hc284ee9f, 32'h429788e5, 32'h429762c5, 32'hc2c51e2a, 32'h425dea33, 32'h4185e712, 32'h41d7f6da, 32'hc2c32588};
test_weights[38952:38959] = '{32'hc22e7b2d, 32'hc1eb6784, 32'hc2b335a6, 32'h41ea437f, 32'h427cd32c, 32'hc08093a2, 32'hc2525235, 32'hbcdf28ee};
test_bias[4869:4869] = '{32'hc2379604};
test_output[4869:4869] = '{32'hc5db70c2};
test_input[38960:38967] = '{32'h42ba2ee1, 32'hc284c1f0, 32'h42851463, 32'hc1bf055d, 32'h42008b5f, 32'h4214c9cf, 32'h429238d8, 32'h42053801};
test_weights[38960:38967] = '{32'h4205ab9e, 32'h42c2978e, 32'hc1b77786, 32'h41c17623, 32'hc1801de9, 32'h42aacc16, 32'h40b5c804, 32'hc220224f};
test_bias[4870:4870] = '{32'h429e42ee};
test_output[4870:4870] = '{32'hc562bd28};
test_input[38968:38975] = '{32'hc17fe221, 32'h4218eeae, 32'h42780a01, 32'hc17a7f0a, 32'hc22c5d7d, 32'hc29c17cd, 32'h41c817c9, 32'hc2c16e81};
test_weights[38968:38975] = '{32'h4252002b, 32'hc1b2c10c, 32'hc1c2475b, 32'hc2a1830a, 32'h404a0c36, 32'h4214a666, 32'h41d21cd1, 32'hc2b8b70d};
test_bias[4871:4871] = '{32'hc1e247d5};
test_output[4871:4871] = '{32'h458f68fc};
test_input[38976:38983] = '{32'h4294e998, 32'h41f19ffb, 32'hc291cce2, 32'hc22b7ed9, 32'hc2a40bc7, 32'hc157f713, 32'hc26058f2, 32'hc215383a};
test_weights[38976:38983] = '{32'h424bb969, 32'h42981085, 32'h429d36cc, 32'hc09d94a6, 32'h42881daa, 32'hc1e83bf0, 32'hc1958824, 32'h42ae8d11};
test_bias[4872:4872] = '{32'h42af4e24};
test_output[4872:4872] = '{32'hc5d2a8a7};
test_input[38984:38991] = '{32'h416fc006, 32'hc26ef1f1, 32'h4112fde7, 32'h4241f9a7, 32'h41b48353, 32'h4177bec7, 32'h42583bde, 32'h42c30ec4};
test_weights[38984:38991] = '{32'hc2b38eb3, 32'hc281b4cf, 32'h429b27f4, 32'hc26e4018, 32'hc21da2ea, 32'h429f71a7, 32'hc21eef58, 32'h4254968c};
test_bias[4873:4873] = '{32'h42a02e48};
test_output[4873:4873] = '{32'h456e5ccf};
test_input[38992:38999] = '{32'h421a893b, 32'h4285e02a, 32'hc2b53913, 32'hc21eb87e, 32'h411b63df, 32'hc27e17b3, 32'h4253e994, 32'h4218d7cd};
test_weights[38992:38999] = '{32'h428a3075, 32'h4233f5e4, 32'h42acf686, 32'hc2b9c6fd, 32'hc246d0ae, 32'hc214babc, 32'hc2331066, 32'hc1b40614};
test_bias[4874:4874] = '{32'h4101a3c6};
test_output[4874:4874] = '{32'h433a6b3d};
test_input[39000:39007] = '{32'hc29c505f, 32'h42b85ec4, 32'h41671c65, 32'hc262f848, 32'hc25378f1, 32'h4079a4e4, 32'h42535fae, 32'h4271932a};
test_weights[39000:39007] = '{32'hc288086e, 32'h42962c38, 32'h419a1fd1, 32'hc0fd7d44, 32'hc1ea89a9, 32'h4185791c, 32'hc2358610, 32'h42baee19};
test_bias[4875:4875] = '{32'hc2b28985};
test_output[4875:4875] = '{32'h468a93e4};
test_input[39008:39015] = '{32'h422c4b0a, 32'h42166a4d, 32'hc24b133c, 32'h4019be1f, 32'h40dd5e2f, 32'h424d3240, 32'h420793f2, 32'hc233f9ca};
test_weights[39008:39015] = '{32'h4169e79d, 32'h42b7a621, 32'hc238a207, 32'h428ac3f7, 32'h4273787c, 32'hc01f2c68, 32'hc196acc7, 32'h424188ae};
test_bias[4876:4876] = '{32'hc20c9679};
test_output[4876:4876] = '{32'h457c3b3a};
test_input[39016:39023] = '{32'hc2778415, 32'h42b126dd, 32'h401a5724, 32'h41f24d6a, 32'h4222b275, 32'hc046e1b0, 32'h41be4da7, 32'h4008d72b};
test_weights[39016:39023] = '{32'hc25379aa, 32'hc27ee62c, 32'h412d4270, 32'hc282623f, 32'hc27e9b22, 32'hbde40ad9, 32'hc27da863, 32'hc0fefceb};
test_bias[4877:4877] = '{32'h4156894f};
test_output[4877:4877] = '{32'hc60398b3};
test_input[39024:39031] = '{32'h414bd461, 32'h41def27f, 32'hc2450268, 32'hc1f441b2, 32'hc2277b28, 32'hc23277d4, 32'hc2850cdb, 32'hc219f9e0};
test_weights[39024:39031] = '{32'hc2184b46, 32'h42396d93, 32'h42556405, 32'h41667477, 32'hc27b123d, 32'hc1bb49c1, 32'h429829d7, 32'hc1d0a0fc};
test_bias[4878:4878] = '{32'h41dec1e8};
test_output[4878:4878] = '{32'hc5239656};
test_input[39032:39039] = '{32'h4274e617, 32'hc1567952, 32'h428eaeb9, 32'h427a33cc, 32'h4227c117, 32'h42ae2222, 32'hc2843253, 32'h4224b505};
test_weights[39032:39039] = '{32'h425235c9, 32'hc28123cb, 32'hc2464166, 32'h4272657f, 32'hc0bcb433, 32'hc022035f, 32'hc0804ef0, 32'hc2bb28e2};
test_bias[4879:4879] = '{32'hc2abd7e6};
test_output[4879:4879] = '{32'h4343af12};
test_input[39040:39047] = '{32'hc0bc37a9, 32'hc279f5db, 32'hc1ae64a6, 32'hc2831c11, 32'h42a717b5, 32'h41462af9, 32'hc290312f, 32'hc296be3b};
test_weights[39040:39047] = '{32'h41fa7880, 32'h42996d02, 32'h42694b53, 32'h4266bce9, 32'h428540c2, 32'h42666990, 32'hc1f47cba, 32'hc20d5aac};
test_bias[4880:4880] = '{32'hc15ff83a};
test_output[4880:4880] = '{32'h4489baaf};
test_input[39048:39055] = '{32'h42012b83, 32'hc220408d, 32'h42b465a3, 32'hc1bde427, 32'h427aa1d3, 32'hc14b86a8, 32'h42b03f9b, 32'hc280f696};
test_weights[39048:39055] = '{32'hc2a37014, 32'hc1bc0979, 32'h42af00dc, 32'hc232e62b, 32'hc24fecf5, 32'hc26ff0d5, 32'hc11df7e7, 32'hc260a851};
test_bias[4881:4881] = '{32'hc27bc094};
test_output[4881:4881] = '{32'h45e8db92};
test_input[39056:39063] = '{32'h4118f242, 32'hc0badc16, 32'hbfc0a926, 32'h424767e6, 32'hc1bf1d29, 32'h40fb65a6, 32'h41541a53, 32'hc2565de6};
test_weights[39056:39063] = '{32'hc23ef6ea, 32'h429589ae, 32'h42b6d557, 32'h421c46f7, 32'hc2c4a401, 32'h40220ad6, 32'hc18fbf61, 32'hc2ba7392};
test_bias[4882:4882] = '{32'h42a70676};
test_output[4882:4882] = '{32'h45fdf9cf};
test_input[39064:39071] = '{32'hc2be36d5, 32'hc2a01d8c, 32'h42a295d6, 32'h427c8720, 32'h42277952, 32'h422db32f, 32'hc2b843d9, 32'h419b1348};
test_weights[39064:39071] = '{32'hc288e4fb, 32'hc22c1531, 32'hc287e343, 32'hc2bc2d2b, 32'hc2a0fc32, 32'h41ba6869, 32'hc285d2f0, 32'hc265bb1b};
test_bias[4883:4883] = '{32'h424b979c};
test_output[4883:4883] = '{32'h449a5834};
test_input[39072:39079] = '{32'h41130bb5, 32'h40bbbe61, 32'h42baec29, 32'h41731484, 32'hc1e674eb, 32'h425fc013, 32'hc290928d, 32'hc26aac5b};
test_weights[39072:39079] = '{32'hc1ce57ac, 32'hc2069842, 32'h420d77a0, 32'h421ad54b, 32'hc26d2b15, 32'h42a4dbde, 32'h425da2c8, 32'hc261a3cf};
test_bias[4884:4884] = '{32'hc2550a03};
test_output[4884:4884] = '{32'h460d138e};
test_input[39080:39087] = '{32'hc29822e4, 32'hc25fe9bd, 32'hc2754b59, 32'h413f7792, 32'h41b5db2e, 32'h42b7f517, 32'h41340844, 32'h4295ac1f};
test_weights[39080:39087] = '{32'h42255101, 32'hc2587795, 32'h4192b127, 32'h42838fb9, 32'h410af278, 32'hc0999d0c, 32'hc21ac69e, 32'hc1c9b0a6};
test_bias[4885:4885] = '{32'h40edf721};
test_output[4885:4885] = '{32'hc53c2899};
test_input[39088:39095] = '{32'h40820def, 32'h429130c2, 32'h4193be4a, 32'h42bd5183, 32'hc2160c45, 32'h42a64dab, 32'hc1bb4e42, 32'h4292e07f};
test_weights[39088:39095] = '{32'hc2a00616, 32'h420208b1, 32'hc1b49cf1, 32'hc2a4430c, 32'hc2c38acd, 32'hc287268a, 32'hc126d037, 32'hc2b78711};
test_bias[4886:4886] = '{32'h42a54df5};
test_output[4886:4886] = '{32'hc662e112};
test_input[39096:39103] = '{32'h41c012b8, 32'hc2b82bfe, 32'h420c6e91, 32'hc256a7ba, 32'h42ae82dd, 32'h428e3aa2, 32'h42079ff4, 32'hc1bba831};
test_weights[39096:39103] = '{32'h41a0a936, 32'hc1f9a2e0, 32'h42c08e94, 32'hc15c9058, 32'hbfb5b1c6, 32'h42b05aeb, 32'h425babe3, 32'h42b83a3e};
test_bias[4887:4887] = '{32'hc104e2b8};
test_output[4887:4887] = '{32'h46500dcc};
test_input[39104:39111] = '{32'hc193856a, 32'h42643b6e, 32'h413c5c71, 32'h418d4bac, 32'h42399b66, 32'hbff0b23a, 32'h41f63225, 32'hc26e0c6b};
test_weights[39104:39111] = '{32'hc2a21cb6, 32'hc28811ed, 32'h42991ed3, 32'h42c29985, 32'h41fa6075, 32'hc1d50fac, 32'h427b104e, 32'hc2041365};
test_bias[4888:4888] = '{32'hc28fb032};
test_output[4888:4888] = '{32'h45adbd33};
test_input[39112:39119] = '{32'hc226137c, 32'hc23b0140, 32'hc291ce4c, 32'h4241f7f8, 32'h420498a9, 32'hc184113c, 32'hc2bf8c5c, 32'h418a4a28};
test_weights[39112:39119] = '{32'h429e38c6, 32'h4298a298, 32'h426eb5bb, 32'hc10a2440, 32'h42bc8156, 32'h410f311e, 32'h42c3aeac, 32'h424960f3};
test_bias[4889:4889] = '{32'hc147daf2};
test_output[4889:4889] = '{32'hc6860c39};
test_input[39120:39127] = '{32'hc2814ca1, 32'h428d37fd, 32'h42987ccf, 32'h42366c45, 32'hc24861ea, 32'h42854255, 32'hc0ca3fa5, 32'h42a9d2d0};
test_weights[39120:39127] = '{32'hc242890a, 32'hc20e34f6, 32'hc2c2840f, 32'h423103b7, 32'h4298fbf8, 32'h425318f0, 32'h4102b38e, 32'h42b87775};
test_bias[4890:4890] = '{32'h425a18ad};
test_output[4890:4890] = '{32'h452c3c88};
test_input[39128:39135] = '{32'hc2aa0f94, 32'hc232fdc6, 32'hc2c63163, 32'h4257dbb6, 32'h42540f5e, 32'hc2292d02, 32'hc2c7adc2, 32'hc0134a13};
test_weights[39128:39135] = '{32'hc24c1d1e, 32'h42a729c5, 32'h3fb0ce47, 32'hc299b344, 32'hc17b2f2a, 32'h4274ce4d, 32'hc1e0224d, 32'h4288cca4};
test_bias[4891:4891] = '{32'h42867ffd};
test_output[4891:4891] = '{32'hc5897752};
test_input[39136:39143] = '{32'hc2928065, 32'h408d97bc, 32'hc1ec5660, 32'hc28585a8, 32'h41073c3d, 32'hc0c536f3, 32'hc24796ba, 32'hc2c6fa98};
test_weights[39136:39143] = '{32'hc29b68d5, 32'hc2bf77a0, 32'h41bbd8f5, 32'hc2ae771e, 32'hc1aad511, 32'hc28feab9, 32'hc2aeadf8, 32'h4257c038};
test_bias[4892:4892] = '{32'hc285aca5};
test_output[4892:4892] = '{32'h4615c94f};
test_input[39144:39151] = '{32'h42a97168, 32'h42b0910e, 32'h42ad4fa3, 32'hc1bbcbc8, 32'hc24754db, 32'hc04ad2ce, 32'hc0c1b395, 32'h4180c4e2};
test_weights[39144:39151] = '{32'h42aeb531, 32'hc2a7ba00, 32'hc2136c4f, 32'hc297f2be, 32'hc19e8490, 32'h423d91d9, 32'hc280eac2, 32'hc1ff8696};
test_bias[4893:4893] = '{32'hc1b6b7f1};
test_output[4893:4893] = '{32'hc434b518};
test_input[39152:39159] = '{32'h425eeab6, 32'hc2a7661d, 32'hc20c046b, 32'h426ba763, 32'hc1cf9211, 32'hc2add3a7, 32'h42963a04, 32'hc0629925};
test_weights[39152:39159] = '{32'hc2831b9d, 32'h4232f327, 32'hc1d435b7, 32'hc2aa2971, 32'h410bd275, 32'h42918a90, 32'hc246df6b, 32'h419d4752};
test_bias[4894:4894] = '{32'hc1622ee6};
test_output[4894:4894] = '{32'hc6aab6bf};
test_input[39160:39167] = '{32'h42306aa7, 32'hc29616b3, 32'hc1efde1d, 32'h4246e028, 32'h4208d4a9, 32'hc10383f3, 32'h4209d8de, 32'h4287c08e};
test_weights[39160:39167] = '{32'h42c3ca95, 32'hc243ed65, 32'hc2669539, 32'h42176c3b, 32'h425e6943, 32'hc0aca82a, 32'h41bb534c, 32'hc27ab054};
test_bias[4895:4895] = '{32'hc10e6d4c};
test_output[4895:4895] = '{32'h461db9e0};
test_input[39168:39175] = '{32'hc2a645de, 32'h42c01d10, 32'h42ac6fb3, 32'h42937ac8, 32'hc24d2552, 32'h41d38ba4, 32'h42af3a85, 32'hc2bcb4cf};
test_weights[39168:39175] = '{32'hc2a4e17b, 32'h42a52ed5, 32'hc2c2995c, 32'h42c4c779, 32'h41fa87d3, 32'hc277b656, 32'h403e8495, 32'h3fab4971};
test_bias[4896:4896] = '{32'hc171ced4};
test_output[4896:4896] = '{32'h4624851a};
test_input[39176:39183] = '{32'hc23d7d20, 32'h4271efab, 32'h42bc0229, 32'hbec97ca8, 32'h42b57c50, 32'h42785d55, 32'h428578e0, 32'hc20cd91a};
test_weights[39176:39183] = '{32'h4193ded9, 32'h42ade3e2, 32'h41cc1419, 32'hc29ed0d0, 32'h42aca285, 32'h42115e70, 32'h42b85ccc, 32'hc2473348};
test_bias[4897:4897] = '{32'hc2580e86};
test_output[4897:4897] = '{32'h46c1620e};
test_input[39184:39191] = '{32'hc2375f1c, 32'hc218dd3e, 32'h423b94d4, 32'h42b6f102, 32'hc2bc4ede, 32'hc28a31f7, 32'hc2c25b30, 32'hc20570a8};
test_weights[39184:39191] = '{32'h4135b5a0, 32'h4296e0a1, 32'h428e5518, 32'h41886bcc, 32'h422f651b, 32'hc1b5f1b2, 32'h41918df0, 32'hc29f22b5};
test_bias[4898:4898] = '{32'hc278c78a};
test_output[4898:4898] = '{32'hc36f5ea2};
test_input[39192:39199] = '{32'hc2649a84, 32'h42a2890c, 32'h420904ca, 32'hc2932e3e, 32'h420db7a6, 32'hc2263a1e, 32'h42c1faba, 32'hc1a062b9};
test_weights[39192:39199] = '{32'h42378ffc, 32'hc214882e, 32'hc20c7d05, 32'hc079d621, 32'h427f6f28, 32'hc2343b4d, 32'h41c4868c, 32'hc2bb1145};
test_bias[4899:4899] = '{32'h41f74df2};
test_output[4899:4899] = '{32'h44e96d75};
test_input[39200:39207] = '{32'h419c8320, 32'h421bc7ff, 32'h429d8af6, 32'h41d5d5b6, 32'hc2bed21b, 32'hc21a1837, 32'hc251bdd8, 32'hc1c62ed3};
test_weights[39200:39207] = '{32'h41ab0218, 32'h42b5435d, 32'h4276145d, 32'hc2c7ea66, 32'h41c83162, 32'h42c33fb3, 32'hc2990114, 32'h425415a7};
test_bias[4900:4900] = '{32'h418db212};
test_output[4900:4900] = '{32'h452814ff};
test_input[39208:39215] = '{32'hc282f811, 32'h424465bb, 32'h4257421b, 32'hc0c904e7, 32'h4226811b, 32'h429de45e, 32'hc2b30976, 32'hc290f36e};
test_weights[39208:39215] = '{32'hc08c80b0, 32'h42373807, 32'hc1a14090, 32'hc2180532, 32'hc0fb6f69, 32'h4201d99d, 32'hc2aa2751, 32'h42a006d3};
test_bias[4901:4901] = '{32'h424c5d10};
test_output[4901:4901] = '{32'h45b51243};
test_input[39216:39223] = '{32'h429e71c3, 32'hc2c4b958, 32'hc1d47e0d, 32'hc22af4d4, 32'hbf87a14e, 32'hc19b4acd, 32'h42a08979, 32'h42a68278};
test_weights[39216:39223] = '{32'h4128c64e, 32'hc2b72ded, 32'h4293038c, 32'h4138b07c, 32'h41acc439, 32'hc2be7bb3, 32'hc26c8dfb, 32'h414ccfe9};
test_bias[4902:4902] = '{32'h41bd3ecd};
test_output[4902:4902] = '{32'h45adf903};
test_input[39224:39231] = '{32'h4203bd2b, 32'hc2b8fb1d, 32'h41919a10, 32'hc23a292c, 32'hc2a569b5, 32'hc1ccae4d, 32'hc2525c2c, 32'hc243dfea};
test_weights[39224:39231] = '{32'hc181c3e8, 32'h42617383, 32'h4294ad1c, 32'h42aa9ee1, 32'h42aa6976, 32'h4225b938, 32'h418d3fb4, 32'hc2955b08};
test_bias[4903:4903] = '{32'h425acc65};
test_output[4903:4903] = '{32'hc655e2c8};
test_input[39232:39239] = '{32'h429fc98f, 32'hc13d4c7b, 32'hc1cf4680, 32'h424cd03f, 32'h420a1657, 32'h415012a0, 32'h427a20a6, 32'hc252d3cf};
test_weights[39232:39239] = '{32'h41c1a178, 32'h4295ec8a, 32'hc2953b32, 32'h42505df2, 32'hc28c2fa4, 32'hc0cb4891, 32'h42100614, 32'hc1909cfd};
test_bias[4904:4904] = '{32'hc29838a1};
test_output[4904:4904] = '{32'h45c4097b};
test_input[39240:39247] = '{32'h4147b39d, 32'h416ed5e8, 32'h42bb20b9, 32'hc24554c6, 32'hc2bfcfe5, 32'hc2bc162d, 32'h40e337b7, 32'hc0620a56};
test_weights[39240:39247] = '{32'hc2b17d99, 32'h411c3426, 32'h42ad8195, 32'hc160b7ef, 32'h409839da, 32'h4284c683, 32'h40f73332, 32'h42ada4fc};
test_bias[4905:4905] = '{32'hc1e65499};
test_output[4905:4905] = '{32'h4458f0e9};
test_input[39248:39255] = '{32'hc29305a6, 32'h40fffe03, 32'h42b22310, 32'hc2b14258, 32'h4249b360, 32'h42be4f74, 32'hc2438ea3, 32'hc1bba356};
test_weights[39248:39255] = '{32'hc23e1fe0, 32'hc21074b5, 32'hc2b5a1c2, 32'hbe7e7d83, 32'hc259b040, 32'hc24d59eb, 32'h40faa036, 32'h423ece47};
test_bias[4906:4906] = '{32'hc2140112};
test_output[4906:4906] = '{32'hc65b36be};
test_input[39256:39263] = '{32'hbf7794a7, 32'h4284c1cc, 32'h422e4bb9, 32'hc240ffa8, 32'h422d9a7b, 32'h42a7512a, 32'h4250985d, 32'h429cac6b};
test_weights[39256:39263] = '{32'h42a6d6ce, 32'h42991fd4, 32'hc21ace21, 32'h42bcf2f5, 32'hc1136eac, 32'h42a589b0, 32'hc2171b09, 32'h42c4c044};
test_bias[4907:4907] = '{32'hbe7a6c18};
test_output[4907:4907] = '{32'h462c250b};
test_input[39264:39271] = '{32'hc2160f97, 32'h425dcfef, 32'hc22767ef, 32'h42bff040, 32'h3dcf922a, 32'h40647ab5, 32'hc1338b9c, 32'hc29eb758};
test_weights[39264:39271] = '{32'h4247a5cc, 32'h41574e8b, 32'hc2602968, 32'hc2c3f301, 32'h426ad943, 32'hc0f22da6, 32'hc29f4d9c, 32'h415995a2};
test_bias[4908:4908] = '{32'hc2287c0b};
test_output[4908:4908] = '{32'hc603bfed};
test_input[39272:39279] = '{32'h418dc941, 32'h421630af, 32'hc0757741, 32'hc291ef74, 32'h42859d42, 32'hc237cd89, 32'hc17e7a7e, 32'hc29a2f7d};
test_weights[39272:39279] = '{32'hc2520de1, 32'hc2c05994, 32'hc297aa93, 32'hc29e87df, 32'h42aeab6d, 32'hc2b5c33a, 32'h427a7c4b, 32'h428482ea};
test_bias[4909:4909] = '{32'h3fab7b72};
test_output[4909:4909] = '{32'h45aa07e3};
test_input[39280:39287] = '{32'hc25b9e49, 32'h42590ae4, 32'hc29aae88, 32'hc27ac106, 32'hc25d1b3f, 32'h425b396a, 32'hc241e30d, 32'h42843c9b};
test_weights[39280:39287] = '{32'h420d549c, 32'hc280cd4b, 32'hc2801a96, 32'h41d80fe8, 32'hc14883ee, 32'hc20c784d, 32'hc1d6df33, 32'h4122947a};
test_bias[4910:4910] = '{32'h40a4bc5d};
test_output[4910:4910] = '{32'hc4b253ef};
test_input[39288:39295] = '{32'hc18f1d3c, 32'hc2c044e0, 32'h42b07d2b, 32'h4268bd23, 32'hc1cef999, 32'hc2b61a8b, 32'h4295a36d, 32'hc187f41d};
test_weights[39288:39295] = '{32'h4106b11a, 32'h42c37580, 32'hc29ee6d1, 32'h4236ae04, 32'h42c0172c, 32'hc2c5926d, 32'hc222e76b, 32'h4282c311};
test_bias[4911:4911] = '{32'h42b253c3};
test_output[4911:4911] = '{32'hc6330b4a};
test_input[39296:39303] = '{32'h41bba6e6, 32'h41b73361, 32'hc2858654, 32'hc257ed26, 32'h428be02d, 32'h415279d6, 32'h4295b4d2, 32'h42462dc0};
test_weights[39296:39303] = '{32'h41b4e1b8, 32'hc19e0e7b, 32'hc131be88, 32'hc2809ca6, 32'hc2b8082b, 32'h42645e63, 32'hc2b29782, 32'hc2b56166};
test_bias[4912:4912] = '{32'h42400635};
test_output[4912:4912] = '{32'hc643aaf5};
test_input[39304:39311] = '{32'hc173da7e, 32'hc28da6c9, 32'h42303970, 32'h426ae305, 32'h42a4eae5, 32'h41bbd35b, 32'hc2baadcc, 32'hc1a7aa66};
test_weights[39304:39311] = '{32'hc2a36f98, 32'hc2c188ba, 32'hc2175fac, 32'hc296607a, 32'h412a04ba, 32'h425577d5, 32'hc15dce87, 32'hc085c0dd};
test_bias[4913:4913] = '{32'hc2aaea82};
test_output[4913:4913] = '{32'h45aa0f3f};
test_input[39312:39319] = '{32'h41852958, 32'hc2ab7b62, 32'h42a7f968, 32'hc15a4090, 32'h4252bf68, 32'hc2b40a99, 32'h418201d7, 32'h41de9539};
test_weights[39312:39319] = '{32'hc2c1d3be, 32'hc20ec860, 32'h42973533, 32'h4202c576, 32'hc230c2d5, 32'h416b2d0b, 32'hc2a931e1, 32'h411e789d};
test_bias[4914:4914] = '{32'h416d3359};
test_output[4914:4914] = '{32'h452376e1};
test_input[39320:39327] = '{32'hc1db774a, 32'hc1892e7b, 32'h41af57e6, 32'hc25ffa01, 32'hbfcb689b, 32'hc2a49f71, 32'h42906362, 32'h428db724};
test_weights[39320:39327] = '{32'h41c59ff2, 32'hc23fe09b, 32'h42936aa6, 32'h3f8f1d66, 32'hc2bf8ff6, 32'hc236c0c7, 32'h42395869, 32'hc244b092};
test_bias[4915:4915] = '{32'hc11309a9};
test_output[4915:4915] = '{32'h45aab3a0};
test_input[39328:39335] = '{32'hc281304b, 32'h4295916d, 32'hc1e004e0, 32'h422ef408, 32'h428c6435, 32'hc214d954, 32'h4139b9c5, 32'h42553344};
test_weights[39328:39335] = '{32'hc2b11f87, 32'hc1cc0b99, 32'h4278482a, 32'h4227431d, 32'h3f3081bf, 32'h42ae8fd1, 32'h42ab50cf, 32'h428a7672};
test_bias[4916:4916] = '{32'hc094a270};
test_output[4916:4916] = '{32'h45a8413b};
test_input[39336:39343] = '{32'hc2aa9933, 32'h42140066, 32'hc1bea231, 32'h4266b7a1, 32'hc25e5051, 32'hbfe6f472, 32'h413844ad, 32'hc28ecd83};
test_weights[39336:39343] = '{32'h41d5794d, 32'h41f645b8, 32'hc194ddec, 32'h42ab1966, 32'h42b51691, 32'hc22cb6ad, 32'h4212ebc4, 32'hc185ad7f};
test_bias[4917:4917] = '{32'h428bc158};
test_output[4917:4917] = '{32'h447315e1};
test_input[39344:39351] = '{32'hc2816511, 32'h40aa6de7, 32'hc29e30fc, 32'hc28db014, 32'hc22daefb, 32'hc28e1c39, 32'h416d519c, 32'hc118bccb};
test_weights[39344:39351] = '{32'h42a6acb5, 32'h42351f8e, 32'hc19aa952, 32'h428ac338, 32'h420a0ccd, 32'h4288b786, 32'hc2bc32e9, 32'h427c8c48};
test_bias[4918:4918] = '{32'hc247ae20};
test_output[4918:4918] = '{32'hc6845995};
test_input[39352:39359] = '{32'h41f8fca8, 32'h407a42de, 32'hc20d104f, 32'h42915642, 32'h42a7b63a, 32'h42969d2b, 32'h4191524c, 32'h42b192f5};
test_weights[39352:39359] = '{32'h425cf4a2, 32'h429afc94, 32'h42b77f6f, 32'hc1a8446b, 32'hc2772c6c, 32'h42b9f78d, 32'hc147d4cd, 32'hc1bc851b};
test_bias[4919:4919] = '{32'h42ac6a08};
test_output[4919:4919] = '{32'hc5452328};
test_input[39360:39367] = '{32'h41fe4890, 32'h4147a109, 32'hc29f702d, 32'hc1dbfa10, 32'h41b6c287, 32'h42471778, 32'h42398cc4, 32'h4253feb5};
test_weights[39360:39367] = '{32'hc25f0541, 32'hc25ff951, 32'hc2ae5899, 32'hc2b8d250, 32'h425d9d08, 32'h42ab86e3, 32'hc2b7c585, 32'hc29e0069};
test_bias[4920:4920] = '{32'h429a00bd};
test_output[4920:4920] = '{32'h4582ad46};
test_input[39368:39375] = '{32'hc20444a4, 32'h42bb3440, 32'hc25eb088, 32'hc2207485, 32'h42be6c1e, 32'hc2406539, 32'hc285b60a, 32'h41b53439};
test_weights[39368:39375] = '{32'hc2807ccd, 32'h42b0507b, 32'hc26aee69, 32'hc146a1b9, 32'hbf3c297b, 32'h420b0f5f, 32'hc2c41a48, 32'hc204f749};
test_bias[4921:4921] = '{32'h413f76bc};
test_output[4921:4921] = '{32'h468e5000};
test_input[39376:39383] = '{32'h421d5889, 32'h42121f0a, 32'h426a4d5b, 32'hc1c7d229, 32'hc25c02e0, 32'hc1851853, 32'hc29f0b8c, 32'hc25b092f};
test_weights[39376:39383] = '{32'hc1e690cd, 32'h428fcf22, 32'hc13c8972, 32'hbf7a701f, 32'h424d7021, 32'hc11ba372, 32'hc2a8282f, 32'hc25e6fed};
test_bias[4922:4922] = '{32'h429f9f67};
test_output[4922:4922] = '{32'h45f9395c};
test_input[39384:39391] = '{32'h428635f0, 32'hc2342ea7, 32'h415a02c5, 32'hc2848baa, 32'hc20fc3d5, 32'hc1d5b38d, 32'hc2119c31, 32'hc2a592c7};
test_weights[39384:39391] = '{32'h413dda2a, 32'hc23ae829, 32'h429f29e1, 32'hc02b632e, 32'h41b19f2a, 32'h4290cf5c, 32'hc2adddd6, 32'h42729763};
test_bias[4923:4923] = '{32'h424cab05};
test_output[4923:4923] = '{32'hc3bb241b};
test_input[39392:39399] = '{32'hbf965e23, 32'hc2bf6eec, 32'hc1629852, 32'hc29f0d4c, 32'hc2c30a1a, 32'hbed6f8ff, 32'hc0cfb0c8, 32'h42b29349};
test_weights[39392:39399] = '{32'h428243a3, 32'h41d0958e, 32'h41e78546, 32'h42450fa8, 32'h42233470, 32'h42b031a8, 32'hc040dc40, 32'hc2807e15};
test_bias[4924:4924] = '{32'h41991d52};
test_output[4924:4924] = '{32'hc681caf2};
test_input[39400:39407] = '{32'h417ea6c4, 32'hc207b0e4, 32'hc20db4ad, 32'h4256c637, 32'hc239d805, 32'h4281992d, 32'h41df9814, 32'h4120fb7d};
test_weights[39400:39407] = '{32'h41adc8ae, 32'h4241c85a, 32'hc181d01b, 32'h42a34e54, 32'h42c7a640, 32'h42c052e3, 32'hc109cc70, 32'h42586e01};
test_bias[4925:4925] = '{32'h42a70aea};
test_output[4925:4925] = '{32'h45b04f15};
test_input[39408:39415] = '{32'h42701afe, 32'hc2735437, 32'hc22727e5, 32'hc2662e9f, 32'h42a860b9, 32'h42435a42, 32'hc2a93330, 32'hc0eac037};
test_weights[39408:39415] = '{32'h4272cfcf, 32'hc1f9daa3, 32'h4271af8f, 32'hc28ceb56, 32'h423c693b, 32'h42a4b267, 32'h41e343ee, 32'h421ff7e2};
test_bias[4926:4926] = '{32'h429003bb};
test_output[4926:4926] = '{32'h46424fbc};
test_input[39416:39423] = '{32'hc2c2b5b8, 32'hc2c51eee, 32'h4295fae7, 32'hc294b5a0, 32'hc269514a, 32'hc240cc0e, 32'h41bbcaba, 32'hc29b18ba};
test_weights[39416:39423] = '{32'hc197af57, 32'hc29603b1, 32'hc221b0d1, 32'h4143a310, 32'h427add1b, 32'hc232365a, 32'h41f7882e, 32'hc185d940};
test_bias[4927:4927] = '{32'hc2b20677};
test_output[4927:4927] = '{32'h45b2d1b5};
test_input[39424:39431] = '{32'hc2b8d0dd, 32'hc27ab8f3, 32'h42a0fa16, 32'h427a8964, 32'h4143d9b7, 32'hc2bfe0fb, 32'h40e98f3c, 32'hc2c77f5a};
test_weights[39424:39431] = '{32'hc20f00f0, 32'h40431c06, 32'hc1c997a3, 32'h420661a2, 32'h3fadb3b6, 32'hc0a3a698, 32'hc287a9bf, 32'hc29fdd97};
test_bias[4928:4928] = '{32'h41857412};
test_output[4928:4928] = '{32'h462eda72};
test_input[39432:39439] = '{32'h3f509185, 32'h428c5ce9, 32'hc1c34b88, 32'hc2398e04, 32'hc2331c83, 32'hc1d8ec64, 32'h42bbc4fb, 32'h42832901};
test_weights[39432:39439] = '{32'hc2a1799d, 32'h424fb9d6, 32'h42b1479b, 32'hc29ee19d, 32'hc26c6ac5, 32'h42c26f26, 32'h42a19a43, 32'hc19985ae};
test_bias[4929:4929] = '{32'h4233602d};
test_output[4929:4929] = '{32'h46336bd8};
test_input[39440:39447] = '{32'hc2b8c03f, 32'hc2961640, 32'h41d54136, 32'hc25f69b1, 32'hc107e015, 32'hc2a95c34, 32'hc196c695, 32'h428ff649};
test_weights[39440:39447] = '{32'hc18121d4, 32'hc29e189e, 32'h42b84bc7, 32'hc2864685, 32'h4290d893, 32'hc245aae3, 32'hc25049ed, 32'h4272cf28};
test_bias[4930:4930] = '{32'h42485ae2};
test_output[4930:4930] = '{32'h46b08fb5};
test_input[39448:39455] = '{32'h41fda14d, 32'h42270dcc, 32'hc127a35b, 32'hc29f0d7d, 32'hc2a05c74, 32'h4189d2f1, 32'h420e35fb, 32'hc124aee3};
test_weights[39448:39455] = '{32'h420b38d9, 32'h42c51b40, 32'hc19caefc, 32'h428040e2, 32'h41be154d, 32'hc131c9c4, 32'hc1ed0b64, 32'hc1ca0864};
test_bias[4931:4931] = '{32'hc10a328f};
test_output[4931:4931] = '{32'hc520de08};
test_input[39456:39463] = '{32'h429a8968, 32'hc2361cfe, 32'h42870bd2, 32'hc268aa46, 32'h426393ad, 32'hc0fcede6, 32'hc29d322c, 32'h42832cc1};
test_weights[39456:39463] = '{32'h42a27644, 32'hc21de425, 32'h42bd250e, 32'hc2827a29, 32'hc2324185, 32'h420422b2, 32'hbfe7b41e, 32'h417bbfe0};
test_bias[4932:4932] = '{32'hc2bbdcde};
test_output[4932:4932] = '{32'h46813404};
test_input[39464:39471] = '{32'h42c08392, 32'h3ffeab0b, 32'hc267e544, 32'h4239bda8, 32'h4213cd41, 32'hc27d7dd4, 32'h4257b0af, 32'h4288e162};
test_weights[39464:39471] = '{32'hc1076a38, 32'h429a797f, 32'hc2a8c299, 32'h42548022, 32'hc2737632, 32'hc2a78d8f, 32'hc2af402c, 32'h419b0960};
test_bias[4933:4933] = '{32'h4233411f};
test_output[4933:4933] = '{32'h45c8206a};
test_input[39472:39479] = '{32'h42895cb1, 32'hc2bad06e, 32'hc20fdb69, 32'hc289d9ac, 32'hc292aba4, 32'h426c50be, 32'h42bc278d, 32'h40d56caa};
test_weights[39472:39479] = '{32'h40d5367c, 32'h42badfa5, 32'hc284cf11, 32'h41e2c3d4, 32'hc2ad4ea8, 32'hc174c8ed, 32'h429f0ea5, 32'h41d424c5};
test_bias[4934:4934] = '{32'h426c301c};
test_output[4934:4934] = '{32'h45a6a88f};
test_input[39480:39487] = '{32'h42bbc074, 32'hc1130e05, 32'hc2765768, 32'hc21b82f4, 32'h41e89f3a, 32'hc25b2aa3, 32'hc2140a86, 32'h417ec582};
test_weights[39480:39487] = '{32'hc24ffdde, 32'h4207ebd8, 32'hc1d095b2, 32'hc2bf76a9, 32'h42276953, 32'h40a606b4, 32'hc264eb50, 32'hc2c01b38};
test_bias[4935:4935] = '{32'h42248c6e};
test_output[4935:4935] = '{32'h44d40bda};
test_input[39488:39495] = '{32'h424f4174, 32'hc2b8a26a, 32'h4191d627, 32'hc28d517f, 32'hc291d28c, 32'h42957932, 32'h42899a38, 32'h42880e38};
test_weights[39488:39495] = '{32'hc2ab2337, 32'h426f7d17, 32'hc20d605d, 32'hc1a6893b, 32'hc22f7c52, 32'h42310e3b, 32'hc155fea5, 32'hc1070309};
test_bias[4936:4936] = '{32'hc2867f1f};
test_output[4936:4936] = '{32'hc582e734};
test_input[39496:39503] = '{32'h42a6107c, 32'h420772a9, 32'h42b05934, 32'hc219ad8e, 32'hc2be7943, 32'h42a120d6, 32'h426c048b, 32'h4105d0fd};
test_weights[39496:39503] = '{32'hc2c7b9db, 32'h42ac95ec, 32'hc2a224d8, 32'h423c0203, 32'h42825845, 32'h41a6dad8, 32'hc2a191c9, 32'hc099afea};
test_bias[4937:4937] = '{32'hc23cd40f};
test_output[4937:4937] = '{32'hc6b93129};
test_input[39504:39511] = '{32'hc1e1aac1, 32'h42c70121, 32'h4289bf6c, 32'hc2aa14e0, 32'h420573e2, 32'hc2b41f0b, 32'hc1bccff7, 32'h42c3a026};
test_weights[39504:39511] = '{32'hc1c82740, 32'h402afb1f, 32'h423b6e33, 32'h42b1073d, 32'hc22a57db, 32'hc2c16bf6, 32'h4269ac01, 32'h42808b1b};
test_bias[4938:4938] = '{32'h3fb7631b};
test_output[4938:4938] = '{32'h460a9765};
test_input[39512:39519] = '{32'hc25493a6, 32'h423efc97, 32'hc1b83224, 32'hc29941e6, 32'h41ee9e9c, 32'hc2648d96, 32'h42327313, 32'h4284a203};
test_weights[39512:39519] = '{32'h428cf452, 32'h419527b1, 32'hc276e580, 32'h42bfe8b0, 32'hc2290e4b, 32'hc1405dc5, 32'hc206b565, 32'hc1c738ee};
test_bias[4939:4939] = '{32'h42648222};
test_output[4939:4939] = '{32'hc642a571};
test_input[39520:39527] = '{32'h421a4a47, 32'hc20b150a, 32'hc29c81b3, 32'h42080ff0, 32'h400ddbdf, 32'h4295053f, 32'hc2a9c2fe, 32'h41a976ff};
test_weights[39520:39527] = '{32'h423d5c0f, 32'hc134d48e, 32'hc2be1471, 32'h4209f3e8, 32'hc191a2b0, 32'h41ea9e40, 32'hc20292d0, 32'hc28f70c6};
test_bias[4940:4940] = '{32'hc28c49a0};
test_output[4940:4940] = '{32'h465d2e2e};
test_input[39528:39535] = '{32'h423a057d, 32'h42b5cb3d, 32'hc280d0f4, 32'hc081fc61, 32'hc1af19ad, 32'h42a19b4b, 32'h40eb5d05, 32'h41b5c0ee};
test_weights[39528:39535] = '{32'hbe8aa948, 32'hc2559273, 32'hc2589bb3, 32'h40f0a05f, 32'h41b1179a, 32'hc2970c4e, 32'hc2b84d85, 32'h41de0d99};
test_bias[4941:4941] = '{32'hc21d26d7};
test_output[4941:4941] = '{32'hc5fc911c};
test_input[39536:39543] = '{32'hc2843168, 32'h4228c263, 32'hc29f6b8c, 32'hbf6f441d, 32'hc2b4bf6e, 32'h41c0ee2c, 32'hc1c7adf8, 32'hc232c1b3};
test_weights[39536:39543] = '{32'hc2a22017, 32'hc29e995a, 32'hc2652655, 32'hc1e5d264, 32'hc222d669, 32'h42292d48, 32'hc29a42ec, 32'hc1ed59f6};
test_bias[4942:4942] = '{32'h41d4d6aa};
test_output[4942:4942] = '{32'h4663d912};
test_input[39544:39551] = '{32'hc28d314c, 32'h3e49a31d, 32'h42802768, 32'h42a6f0ad, 32'h42946a8b, 32'h42964a58, 32'hc22e558c, 32'h42238862};
test_weights[39544:39551] = '{32'hc29e6575, 32'hc2402aeb, 32'h41ec2df5, 32'h429d7e93, 32'h40a997ba, 32'hc2bac343, 32'h42a4d4d6, 32'hc2af2086};
test_bias[4943:4943] = '{32'h413b41df};
test_output[4943:4943] = '{32'h43832e83};
test_input[39552:39559] = '{32'hc2bad0fd, 32'h42b62a21, 32'hc2821739, 32'h42731739, 32'h42b0fa80, 32'hc29e66e3, 32'hc2a53c03, 32'hc24adcc9};
test_weights[39552:39559] = '{32'h42b0e1db, 32'h417eaa5d, 32'h42762a7f, 32'h42a7bfca, 32'hc288b5ac, 32'hc290396a, 32'hc2185e41, 32'h4236d95c};
test_bias[4944:4944] = '{32'hc26806f2};
test_output[4944:4944] = '{32'hc5a51d9f};
test_input[39560:39567] = '{32'h42c4fbb9, 32'h41cbd84c, 32'hc2b8dfdb, 32'hc1cb570c, 32'h42192863, 32'hc183ea3c, 32'hc2b0a5da, 32'hc27af3a4};
test_weights[39560:39567] = '{32'h41c726df, 32'hc18b6f31, 32'hc2b425f2, 32'hc28006b4, 32'hc241ad57, 32'hc175b6e5, 32'h420d9c2a, 32'hc2b8d77f};
test_bias[4945:4945] = '{32'hc221f795};
test_output[4945:4945] = '{32'h464afcc5};
test_input[39568:39575] = '{32'h4287dad5, 32'hc27631c6, 32'hc27ee0b9, 32'hc15d8d44, 32'hc22f9f4a, 32'hc211393d, 32'hc1ed649c, 32'hc2c69956};
test_weights[39568:39575] = '{32'h42683fac, 32'h416fe516, 32'hc1d1dd3e, 32'hc029b756, 32'hc27c626c, 32'hc0c77186, 32'h4156eb29, 32'h4249baef};
test_bias[4946:4946] = '{32'h42b727aa};
test_output[4946:4946] = '{32'h4516b11b};
test_input[39576:39583] = '{32'h42bb5f80, 32'hc2598c43, 32'h4201d5b7, 32'h428f3942, 32'h42c60697, 32'hc29c00aa, 32'hc1468c11, 32'hbe61cdc9};
test_weights[39576:39583] = '{32'h41a8eb49, 32'hc2a6faf3, 32'h4219963e, 32'h428e0bf6, 32'hc2c00898, 32'hc2a404de, 32'hc1bf8370, 32'hc1f2d024};
test_bias[4947:4947] = '{32'h421b12df};
test_output[4947:4947] = '{32'h461d8f6b};
test_input[39584:39591] = '{32'hc2af9da1, 32'h42c39e5e, 32'hc2aa938a, 32'h40f0e3fe, 32'h42c77118, 32'h40667a38, 32'hc110b140, 32'hc23436b8};
test_weights[39584:39591] = '{32'h423e2528, 32'hc28733ce, 32'h4253e85a, 32'hc0d34e99, 32'h4193d846, 32'hc28f2ca2, 32'h41e00f44, 32'hc2b57242};
test_bias[4948:4948] = '{32'hc21a242f};
test_output[4948:4948] = '{32'hc61bd5ad};
test_input[39592:39599] = '{32'hc276939e, 32'h418b5c37, 32'h41cb5005, 32'hc2728bc7, 32'hc2b6323e, 32'hc21e246f, 32'hc276f008, 32'hc243abd6};
test_weights[39592:39599] = '{32'h3fc4eba8, 32'hc0c1ea4e, 32'hc28b275d, 32'h4248268b, 32'hc21772f2, 32'hc29923b0, 32'h4275c4cb, 32'h42a9a524};
test_bias[4949:4949] = '{32'hc1788a8c};
test_output[4949:4949] = '{32'hc5caa25a};
test_input[39600:39607] = '{32'hc28ddf6c, 32'hc2c21df0, 32'h427a9dfc, 32'h423499db, 32'hc1a774c4, 32'h4248b771, 32'h41e17d96, 32'h42bccf1f};
test_weights[39600:39607] = '{32'hc25e55ce, 32'hc28494b0, 32'hc12ae7b2, 32'h400cad08, 32'h40986730, 32'h42bc4bbf, 32'h422636f7, 32'hc2aa3a61};
test_bias[4950:4950] = '{32'h429761e8};
test_output[4950:4950] = '{32'h45eeda84};
test_input[39608:39615] = '{32'h4283d486, 32'h425c4ea0, 32'h425ba653, 32'h42083980, 32'hc29b106c, 32'h4297021e, 32'hc2a51021, 32'h3fd793d8};
test_weights[39608:39615] = '{32'h42bbbe30, 32'h42593860, 32'h42a30c47, 32'h419f01e0, 32'h3fd3862a, 32'hc2a5f229, 32'hc2538852, 32'h42aa2de6};
test_bias[4951:4951] = '{32'hc257cb58};
test_output[4951:4951] = '{32'h4641a41b};
test_input[39616:39623] = '{32'hc29fcbbe, 32'h410f4b08, 32'h42348d6f, 32'hc24a9278, 32'h424b8d12, 32'h42246b3c, 32'hc2772c25, 32'hc27d4a3e};
test_weights[39616:39623] = '{32'h42149919, 32'h422f2f7f, 32'hc206ebb9, 32'h42b5518f, 32'hc23c315d, 32'h41fcfadd, 32'hc26708fb, 32'hc1bef044};
test_bias[4952:4952] = '{32'hc287a5f6};
test_output[4952:4952] = '{32'hc5951b9f};
test_input[39624:39631] = '{32'h42c5cf0b, 32'hc2880a31, 32'hc2484f70, 32'h40ec1097, 32'h418a334b, 32'h41b6d27d, 32'h425aaa7d, 32'hc247d858};
test_weights[39624:39631] = '{32'hc2842758, 32'h4268e3d4, 32'hc29fa7ca, 32'hc1f59e89, 32'hc288ec5c, 32'hc1f1dd25, 32'hc25cbbec, 32'hc0e81936};
test_bias[4953:4953] = '{32'hc298631e};
test_output[4953:4953] = '{32'hc6310259};
test_input[39632:39639] = '{32'hc27bd0c0, 32'hc0dba5e6, 32'h3f468036, 32'h424f2122, 32'h41b45617, 32'hc0afa2ba, 32'h4148ab54, 32'hc2022a12};
test_weights[39632:39639] = '{32'h42aae4dd, 32'h42217b04, 32'h42909ae3, 32'h41b5a285, 32'hc146de1b, 32'hc19cff3b, 32'h41f72516, 32'h41f03d54};
test_bias[4954:4954] = '{32'h41ece387};
test_output[4954:4954] = '{32'hc5a1296e};
test_input[39640:39647] = '{32'hc25c4aa1, 32'hc09e4e00, 32'hc1bfb84a, 32'h4270143a, 32'h412410fe, 32'h418bef39, 32'h41891b5b, 32'hc29021fc};
test_weights[39640:39647] = '{32'h406921a8, 32'hc2a34971, 32'hc2af9639, 32'hc153fa15, 32'hc2a6e56e, 32'hc09937e0, 32'hc134fb84, 32'h427b00c7};
test_bias[4955:4955] = '{32'hc281e14a};
test_output[4955:4955] = '{32'hc583831b};
test_input[39648:39655] = '{32'hc27bb440, 32'h41dbae23, 32'h41845cec, 32'h42ac377e, 32'hc2ba9187, 32'hc1c93c93, 32'h41b9fff3, 32'hc1a75656};
test_weights[39648:39655] = '{32'hc250e536, 32'hc1f44646, 32'h42441fd5, 32'h41814c7a, 32'h42bd04f3, 32'h4258b6c7, 32'hc202911d, 32'hc2a16a3a};
test_bias[4956:4956] = '{32'hc2c67c2b};
test_output[4956:4956] = '{32'hc592d2fc};
test_input[39656:39663] = '{32'h41b24696, 32'hc279337e, 32'h422e3651, 32'h41e8c48c, 32'hc21a9e2c, 32'h40a2eefe, 32'hc2b5aa07, 32'h4284b310};
test_weights[39656:39663] = '{32'h4258f9d7, 32'hc23631f2, 32'hc2a4b221, 32'h423797fa, 32'h421f66f0, 32'hc18d5e33, 32'h42061d05, 32'hc1880757};
test_bias[4957:4957] = '{32'hc13139d6};
test_output[4957:4957] = '{32'hc57b3a0c};
test_input[39664:39671] = '{32'h42be45ad, 32'hc23ec0d3, 32'h40d06ca5, 32'h423c678b, 32'h41a3298a, 32'h422063e2, 32'hc194de6b, 32'h42a9461d};
test_weights[39664:39671] = '{32'hc2a37f5e, 32'hc2733a7c, 32'hc29f76a1, 32'h4280987a, 32'h4265b23e, 32'h3fd8fa8f, 32'hc1aa93f6, 32'h41b4ad9a};
test_bias[4958:4958] = '{32'h42b12530};
test_output[4958:4958] = '{32'h449e7721};
test_input[39672:39679] = '{32'hc10f1e40, 32'h42a38288, 32'hc2834996, 32'h4284a14c, 32'hc2386b4a, 32'hc2bc9498, 32'h424afd8f, 32'h429338ca};
test_weights[39672:39679] = '{32'hc2af3e3d, 32'hc2ba0535, 32'hc274f41d, 32'h429dd8ee, 32'h42680c04, 32'hc287d202, 32'h419d0c2b, 32'hc2b8f07d};
test_bias[4959:4959] = '{32'h40a83366};
test_output[4959:4959] = '{32'h43b26842};
test_input[39680:39687] = '{32'hc28474b5, 32'h42222327, 32'hc2c1049e, 32'hc2aedbe2, 32'h41c2e702, 32'h42c3a7aa, 32'hbf3b425d, 32'hc1c210f9};
test_weights[39680:39687] = '{32'h429158ec, 32'hc2843063, 32'hc1ce64a4, 32'h3f4885cc, 32'hc1ae6bcb, 32'hc2a2fb1c, 32'h41b4adbb, 32'hc2a62b08};
test_bias[4960:4960] = '{32'hc269c007};
test_output[4960:4960] = '{32'hc635c5ab};
test_input[39688:39695] = '{32'h42afcdcf, 32'h42b3f8f0, 32'hc20da2d4, 32'hc2106906, 32'hc2ae8d2b, 32'h428e19b6, 32'hc2c325e2, 32'h4294af67};
test_weights[39688:39695] = '{32'hc2896647, 32'h42139ea7, 32'h422f26b2, 32'h42baafef, 32'h4067672b, 32'hc0ba2b50, 32'hbeca28e3, 32'hc1cdd9e2};
test_bias[4961:4961] = '{32'h42c146cc};
test_output[4961:4961] = '{32'hc61e8419};
test_input[39696:39703] = '{32'hc2b43f69, 32'hc1a00f1b, 32'hc0df6d4a, 32'h423a3b3e, 32'hc1e00929, 32'h40e05999, 32'h4205ed93, 32'h42c22f29};
test_weights[39696:39703] = '{32'hc15f429c, 32'h41758d4e, 32'hc2bd6b93, 32'hc119b9aa, 32'hc2a8dda9, 32'hc251ee6b, 32'h42a81e70, 32'hc219b8f8};
test_bias[4962:4962] = '{32'h41e384c2};
test_output[4962:4962] = '{32'h450e09f2};
test_input[39704:39711] = '{32'h426b17f4, 32'h421ac382, 32'hc1d4c1f7, 32'h422a4b32, 32'h41931bfe, 32'h421d665b, 32'hc2a250de, 32'hc28d7d51};
test_weights[39704:39711] = '{32'h42156a99, 32'h427fa91e, 32'h4221887c, 32'h41bfa386, 32'h422984d7, 32'hc2b16a19, 32'h40ab3d30, 32'h3ea263a7};
test_bias[4963:4963] = '{32'h42552b83};
test_output[4963:4963] = '{32'h44bb6ed7};
test_input[39712:39719] = '{32'h4244a6df, 32'h42c2fe49, 32'hc2c18a37, 32'h41832e62, 32'hc23bd201, 32'h42b6aaa2, 32'h41358420, 32'hc2a3b2dc};
test_weights[39712:39719] = '{32'h42600a06, 32'hc27eee76, 32'hc2bddcf1, 32'hc22929a4, 32'hc1c717d5, 32'hc034137f, 32'hc2ac87f0, 32'hc2a5f55e};
test_bias[4964:4964] = '{32'hc1db1237};
test_output[4964:4964] = '{32'h463748f3};
test_input[39720:39727] = '{32'hc2953675, 32'hc135955c, 32'h4201ec81, 32'hc2388350, 32'hc2acea2c, 32'hc2ae7107, 32'h42b01177, 32'h42ae7667};
test_weights[39720:39727] = '{32'hc29a8be9, 32'h42a9f90f, 32'hc050ad23, 32'hc2c3be90, 32'hbfef7f3a, 32'hc1fa29aa, 32'hc2271186, 32'h41e190ba};
test_bias[4965:4965] = '{32'h42c06852};
test_output[4965:4965] = '{32'h462b855d};
test_input[39728:39735] = '{32'h4122ca05, 32'h41d0ceb1, 32'hc1c3b9fe, 32'h4207460b, 32'hc2593dd2, 32'hc2b49f67, 32'h4275be42, 32'h418a4880};
test_weights[39728:39735] = '{32'h428280a2, 32'hc28d0ffa, 32'h41e071af, 32'hc2617740, 32'hc28bbe36, 32'h410e9666, 32'h4005837c, 32'hc2bcd01a};
test_bias[4966:4966] = '{32'h425755a5};
test_output[4966:4966] = '{32'hc50b59aa};
test_input[39736:39743] = '{32'h41d35598, 32'hc29aea90, 32'h4293310b, 32'h40fcc06c, 32'h42632b5d, 32'hc2aac674, 32'h41dc27ed, 32'h4280e7e1};
test_weights[39736:39743] = '{32'hc25060f2, 32'hc29c1e3c, 32'h429cb6db, 32'hc283d0eb, 32'h428efd6a, 32'h40aa29e8, 32'h40b8da06, 32'h41c99a75};
test_bias[4967:4967] = '{32'h42252586};
test_output[4967:4967] = '{32'h466fcc79};
test_input[39744:39751] = '{32'hc1d67060, 32'hc0808cc8, 32'h428745ce, 32'hc24859ba, 32'hc2c607ee, 32'hc1f7371b, 32'h420f8073, 32'hc221d93e};
test_weights[39744:39751] = '{32'h42b87e0b, 32'h42b7049e, 32'hc23590ea, 32'h429d94fc, 32'hc2bdcdb4, 32'h41bdb498, 32'h4245078b, 32'h4282a9e8};
test_bias[4968:4968] = '{32'h4112eb40};
test_output[4968:4968] = '{32'hc500c049};
test_input[39752:39759] = '{32'hc29f1cd4, 32'hc1502001, 32'h41cf9522, 32'h42280b6e, 32'hc28862cb, 32'h417dd0d9, 32'h429b27ad, 32'hc18969c3};
test_weights[39752:39759] = '{32'hc26fa10a, 32'h41828977, 32'hc15ae348, 32'hc18205d3, 32'hc296e40b, 32'h41850065, 32'h4293668b, 32'h42751e21};
test_bias[4969:4969] = '{32'h421a7452};
test_output[4969:4969] = '{32'h4654f049};
test_input[39760:39767] = '{32'h4240b278, 32'hc2a0934e, 32'hc2c6edd5, 32'h40a60711, 32'hc2847e54, 32'hc2b9222c, 32'hc1839f98, 32'hc2b8f824};
test_weights[39760:39767] = '{32'h3f27a481, 32'hc2ab61a2, 32'h42a45f42, 32'hc257a87e, 32'h42c180d0, 32'hc189dd8d, 32'hc2c4b9cc, 32'h42c2b4b4};
test_bias[4970:4970] = '{32'hc0bd480e};
test_output[4970:4970] = '{32'hc656d158};
test_input[39768:39775] = '{32'hc204f569, 32'h417d9075, 32'hc271089a, 32'h41c7d7c7, 32'hc11e667b, 32'hc2b39455, 32'hc28589d2, 32'h42760362};
test_weights[39768:39775] = '{32'h41e33670, 32'h4294ef66, 32'h3fa5bb26, 32'hc0cd515f, 32'hc2a3a7b3, 32'h420225c9, 32'hc286b12e, 32'hc2a9bb59};
test_bias[4971:4971] = '{32'hc25c43b5};
test_output[4971:4971] = '{32'hc534b8eb};
test_input[39776:39783] = '{32'hc2c08e2f, 32'h429315ad, 32'h42a999e7, 32'h4172d1d5, 32'h4197ee22, 32'h41e4954e, 32'h41a80985, 32'h425c8b15};
test_weights[39776:39783] = '{32'hc2b7b80b, 32'h420272ba, 32'h411ea06b, 32'hc2a1660b, 32'hc2a74242, 32'hc24cbc00, 32'h421cff01, 32'h4283a1d5};
test_bias[4972:4972] = '{32'h425407a1};
test_output[4972:4972] = '{32'h464067cc};
test_input[39784:39791] = '{32'hc21009bd, 32'hc280a741, 32'hc21cd1fa, 32'h42ab2498, 32'h421546c8, 32'h40bffe01, 32'hc1c02871, 32'h41ea48b5};
test_weights[39784:39791] = '{32'hc226798b, 32'h41abd433, 32'h429235ab, 32'h4203abc4, 32'h423f2ced, 32'h422057c2, 32'h42c54e50, 32'hc22197d0};
test_bias[4973:4973] = '{32'h420b1328};
test_output[4973:4973] = '{32'hc4b24151};
test_input[39792:39799] = '{32'h41760be4, 32'h42c25c77, 32'hc25f0332, 32'h42057b46, 32'hc28cfe5b, 32'h42b2ee92, 32'hc293107c, 32'h4284e1c7};
test_weights[39792:39799] = '{32'hc2234a91, 32'h42855366, 32'h41aae4eb, 32'hc149a057, 32'h42a13042, 32'h420f0f1f, 32'h4232c485, 32'h4136e120};
test_bias[4974:4974] = '{32'hc200322b};
test_output[4974:4974] = '{32'hc4487150};
test_input[39800:39807] = '{32'hc2c69603, 32'h42b1160c, 32'hc04021e1, 32'h4238c00f, 32'hc297455a, 32'h416ff99c, 32'hc2800e83, 32'hc18286e1};
test_weights[39800:39807] = '{32'h41b3c89b, 32'hc2c72bdd, 32'hc2a799f5, 32'hc1a42ee7, 32'hc2a89c7f, 32'h4290789e, 32'hc1eb0e02, 32'h413dd224};
test_bias[4975:4975] = '{32'h4285e5a4};
test_output[4975:4975] = '{32'hc51e2c92};
test_input[39808:39815] = '{32'h422a1793, 32'hc17dd026, 32'h42bbdda1, 32'h42ad5d49, 32'h418aa72d, 32'hc2b4a677, 32'hc2685f79, 32'hc20f5ef2};
test_weights[39808:39815] = '{32'hc2afa725, 32'h41c178bf, 32'hc1fc2513, 32'h40a2af9c, 32'h41aac265, 32'hc29c397c, 32'h425bd42d, 32'h4221d0d6};
test_bias[4976:4976] = '{32'hc19d1c0b};
test_output[4976:4976] = '{32'hc5722ffe};
test_input[39816:39823] = '{32'hc279628a, 32'h4213c40d, 32'h42b630a8, 32'hc24597f6, 32'h423dac2b, 32'h42affbd9, 32'h42815ff0, 32'hc1b28624};
test_weights[39816:39823] = '{32'hc255002c, 32'h4209b634, 32'h424c9cfe, 32'hc18c8804, 32'hc1de3f01, 32'hc2ab06fd, 32'hc1c9a449, 32'h42287ac6};
test_bias[4977:4977] = '{32'hc06d8ff9};
test_output[4977:4977] = '{32'hc4a212c7};
test_input[39824:39831] = '{32'h422564cc, 32'h4218dfc8, 32'hc272c66f, 32'hc2b96fae, 32'h420371c8, 32'hc2b3887b, 32'hc2b38cb9, 32'hc277d59a};
test_weights[39824:39831] = '{32'h40cddb22, 32'h42a460a3, 32'hc2c2c51f, 32'h4278cd26, 32'hc22e81fa, 32'h4293a895, 32'hc0a2350d, 32'h4258c04f};
test_bias[4978:4978] = '{32'hc13b5085};
test_output[4978:4978] = '{32'hc5e80303};
test_input[39832:39839] = '{32'hc28e2ef1, 32'hc2b76ec0, 32'h415265dc, 32'h427f758f, 32'h41f8a49a, 32'h4270b9e7, 32'hc29cd468, 32'hc294da2c};
test_weights[39832:39839] = '{32'hc161af7a, 32'hc2105339, 32'hc2b4a1db, 32'h42a97d51, 32'h418e121b, 32'h42a7e4c9, 32'hc2836d0f, 32'hc1f2b035};
test_bias[4979:4979] = '{32'h42b20fa5};
test_output[4979:4979] = '{32'h46a9108e};
test_input[39840:39847] = '{32'h4284fcf4, 32'h429370b4, 32'h41b3de20, 32'h424d3a40, 32'h42110756, 32'hc2282ecd, 32'hc23a607b, 32'hc0cfd2ed};
test_weights[39840:39847] = '{32'h42bd4ff9, 32'hc2698525, 32'h41478c1f, 32'hc025d712, 32'hc13e09ff, 32'hc13534a6, 32'h4210002e, 32'hc238d823};
test_bias[4980:4980] = '{32'hc215e74e};
test_output[4980:4980] = '{32'h44402204};
test_input[39848:39855] = '{32'h41c964f1, 32'hc2967bd6, 32'hc2810158, 32'h42959bad, 32'hc0d9e0b3, 32'hbf8a9d04, 32'hc2a47c33, 32'h420490e8};
test_weights[39848:39855] = '{32'hc2b244a6, 32'h4227c168, 32'h418a1dc1, 32'h41848f0a, 32'hc2985e86, 32'hc29cd855, 32'h419bd424, 32'h4299b1e5};
test_bias[4981:4981] = '{32'hc205513e};
test_output[4981:4981] = '{32'hc56ae60d};
test_input[39856:39863] = '{32'hc254cc8b, 32'h428758c9, 32'hc2bf624a, 32'hc1866d19, 32'hc2387c81, 32'hc1235996, 32'h428e35cb, 32'h421ed924};
test_weights[39856:39863] = '{32'hc212dbd3, 32'h426f0214, 32'hc214492b, 32'h42406990, 32'h41860b76, 32'hc2c7b7f5, 32'h42aba273, 32'h42798b11};
test_bias[4982:4982] = '{32'h40258c3d};
test_output[4982:4982] = '{32'h46893995};
test_input[39864:39871] = '{32'h411746be, 32'h41de99fa, 32'h428c2836, 32'h42acc3d5, 32'hc23152f6, 32'hc2b84f33, 32'hc29b1825, 32'hc243dbe9};
test_weights[39864:39871] = '{32'h42a5040c, 32'h408daaae, 32'hc2022a8f, 32'h41c189b4, 32'h41d8fd00, 32'h42251d06, 32'hc255e5c2, 32'hc1f5904a};
test_bias[4983:4983] = '{32'h41ac47d2};
test_output[4983:4983] = '{32'h44ac3042};
test_input[39872:39879] = '{32'h41a900b2, 32'h4241d5ad, 32'hc237d091, 32'h4248bcc6, 32'hc1e70f6d, 32'h407fc416, 32'hc1f5d599, 32'hc272793a};
test_weights[39872:39879] = '{32'hc2adf54e, 32'hbf4a9fe8, 32'h425485e8, 32'hc2914cf9, 32'hbf8f8d2b, 32'h411edb18, 32'h42c4c193, 32'hbff6a80c};
test_bias[4984:4984] = '{32'hc20f57a8};
test_output[4984:4984] = '{32'hc629454e};
test_input[39880:39887] = '{32'h4281def0, 32'hc253c3ee, 32'hc23d0ecd, 32'h40ed2c26, 32'h3e17e50c, 32'hc0acee58, 32'h42818286, 32'h419597bc};
test_weights[39880:39887] = '{32'hc21ab87c, 32'h425b2cb2, 32'hc2b1b595, 32'hc1a4998e, 32'h42a4a790, 32'hc19f2ffe, 32'h42b164e1, 32'h420b08e5};
test_bias[4985:4985] = '{32'h4011d1ac};
test_output[4985:4985] = '{32'h45a0f147};
test_input[39888:39895] = '{32'hc12174de, 32'h4214ec5b, 32'h40b91219, 32'h428bf3ed, 32'h3fcbd66a, 32'hc215ab85, 32'h4269856e, 32'h426b39d9};
test_weights[39888:39895] = '{32'hc2856e23, 32'hc29437be, 32'hc272e665, 32'hc2b3d6a5, 32'hc1d96e68, 32'hc29a3cb6, 32'hc015744d, 32'hc21104d6};
test_bias[4986:4986] = '{32'hc2275e28};
test_output[4986:4986] = '{32'hc60014e0};
test_input[39896:39903] = '{32'h42013b55, 32'h423c8835, 32'hc2b27cc3, 32'h42b6a4a0, 32'hc2ab0754, 32'h411ad8ef, 32'h4063303a, 32'hc21b84f9};
test_weights[39896:39903] = '{32'h4228d679, 32'h42c5011a, 32'h4199fc2a, 32'hc294a0c1, 32'hbfe43364, 32'hc29caaa7, 32'hc2430400, 32'hc24b6440};
test_bias[4987:4987] = '{32'h42ad138f};
test_output[4987:4987] = '{32'hc497a1cc};
test_input[39904:39911] = '{32'h4230e18c, 32'h42872830, 32'hc2a75d7e, 32'hc2bcdb4b, 32'hc28bfb0a, 32'hc2c459df, 32'h41aa39f7, 32'hc169ab2a};
test_weights[39904:39911] = '{32'hc2713ce4, 32'hc2902e7d, 32'h42012bba, 32'hc1249f59, 32'hc23939e0, 32'h42b7ee81, 32'hc206332b, 32'hc2b1c3f6};
test_bias[4988:4988] = '{32'hc1f1c467};
test_output[4988:4988] = '{32'hc6629d23};
test_input[39912:39919] = '{32'hc23b72d3, 32'h42a34697, 32'hc2ab86da, 32'h4252f9bf, 32'h41fa36b6, 32'hc2b64224, 32'h420c3591, 32'h41f9e2c2};
test_weights[39912:39919] = '{32'hc20fc73f, 32'h42a023bf, 32'hc19fba31, 32'hc1a9f5b7, 32'h4284620d, 32'h42b99b60, 32'h423b165b, 32'hc2b513d5};
test_bias[4989:4989] = '{32'h42acd703};
test_output[4989:4989] = '{32'h44a57e9f};
test_input[39920:39927] = '{32'hc2477fc7, 32'h42aaac84, 32'hc26d66c3, 32'hc2b4d736, 32'h420a401d, 32'hc2656d49, 32'hc21fedc9, 32'hc2617a46};
test_weights[39920:39927] = '{32'h425d2d6f, 32'hc1054495, 32'hc213fd86, 32'h42aa8f3a, 32'hc2a23e92, 32'h410d688b, 32'hc2c40158, 32'hc29de5c7};
test_bias[4990:4990] = '{32'hc0424fda};
test_output[4990:4990] = '{32'hc5758e23};
test_input[39928:39935] = '{32'h415102f1, 32'h4190af1c, 32'h4275d427, 32'h42a63bb0, 32'h42bcdb5b, 32'h42b28df8, 32'hbeb5c2b0, 32'h4291831f};
test_weights[39928:39935] = '{32'hc2b1da77, 32'hc266a1e9, 32'hc22b7c21, 32'h41996d16, 32'h42b1e1e9, 32'hc21e9a8b, 32'hc0da91d4, 32'hc238bc5f};
test_bias[4991:4991] = '{32'hc12a9e0a};
test_output[4991:4991] = '{32'hc4db5d02};
test_input[39936:39943] = '{32'h415515e9, 32'hc13629ad, 32'h40fd7559, 32'h426ec2b4, 32'hc1bf9c64, 32'h4108a684, 32'hc205db9f, 32'h42ba51d9};
test_weights[39936:39943] = '{32'h42a6fab1, 32'h41ea2a73, 32'h428874cd, 32'h42791356, 32'hbfb03db8, 32'hc1e945c1, 32'h42a77318, 32'h4238e56f};
test_bias[4992:4992] = '{32'h42adaeac};
test_output[4992:4992] = '{32'h45c858c5};
test_input[39944:39951] = '{32'h41f02661, 32'h4156c9ec, 32'h41d92c3d, 32'h42b56d46, 32'hc2c60089, 32'h4213bd4f, 32'h42b6b287, 32'h42359eac};
test_weights[39944:39951] = '{32'hc2695cec, 32'hc288923a, 32'hc1854fc0, 32'h420f8018, 32'h41837c5e, 32'hc207340d, 32'h42a6264f, 32'h41e44d86};
test_bias[4993:4993] = '{32'hc26783af};
test_output[4993:4993] = '{32'h45be2870};
test_input[39952:39959] = '{32'h426551c7, 32'h428f4987, 32'h41969d8e, 32'h426d199c, 32'hc273c2e8, 32'hc21a9d3d, 32'h423a3e53, 32'h40d49c62};
test_weights[39952:39959] = '{32'hc2af6664, 32'h428273be, 32'h41217aaa, 32'hc220e3c8, 32'h41ed636c, 32'h40c7cac0, 32'h428dec59, 32'hc03e19a2};
test_bias[4994:4994] = '{32'h423b5fdf};
test_output[4994:4994] = '{32'hc49e6f60};
test_input[39960:39967] = '{32'h41c26c20, 32'h41d41dd9, 32'hc28567bc, 32'hc26b6872, 32'h419c4abc, 32'hc2a47937, 32'h4138a7fa, 32'hc2b68cd0};
test_weights[39960:39967] = '{32'h41a9d801, 32'h428ef0d8, 32'hc24a6184, 32'h42aa6588, 32'h42b25a90, 32'hc14b85e0, 32'hc26e44ad, 32'h42a0395f};
test_bias[4995:4995] = '{32'hc2940543};
test_output[4995:4995] = '{32'hc58d0dcb};
test_input[39968:39975] = '{32'h421a052f, 32'h419a0434, 32'h4200607e, 32'hc2c59c4f, 32'h41c1146d, 32'hc14ca9af, 32'h421c66cd, 32'hc2bb5199};
test_weights[39968:39975] = '{32'h41a2525d, 32'h41c2fc80, 32'h4286caa0, 32'h422b26a5, 32'h42969535, 32'hc2c16d29, 32'hc20183e9, 32'hc215dbe1};
test_bias[4996:4996] = '{32'h42acfbf3};
test_output[4996:4996] = '{32'h458ecc25};
test_input[39976:39983] = '{32'h426691d7, 32'h42168c09, 32'hc29f2dd0, 32'hc24ed376, 32'h425c09ee, 32'h428f44d9, 32'h42a97fbd, 32'hc27049cc};
test_weights[39976:39983] = '{32'h42b423fe, 32'h41fbd77d, 32'h416f31f6, 32'h4083b060, 32'h41ea85b1, 32'hc12ebd3a, 32'h4207d21f, 32'h42a5b965};
test_bias[4997:4997] = '{32'h4159d659};
test_output[4997:4997] = '{32'h45685f39};
test_input[39984:39991] = '{32'hc1b6c7b0, 32'h42a157ab, 32'h42c6a789, 32'h42803655, 32'h42a6919e, 32'hc29e5c99, 32'hc17ada86, 32'hc2b59825};
test_weights[39984:39991] = '{32'h42c65105, 32'hc26fa768, 32'hc246c253, 32'h42161aec, 32'h41913783, 32'hc282d64a, 32'h42417014, 32'hc2a947a1};
test_bias[4998:4998] = '{32'h42a281cf};
test_output[4998:4998] = '{32'h457e71ba};
test_input[39992:39999] = '{32'hc25ef94d, 32'hc19db57d, 32'hc26f2ce2, 32'hc056d127, 32'h4178bfbd, 32'h42bd7c29, 32'h4279519c, 32'h424d1800};
test_weights[39992:39999] = '{32'h4226a0ed, 32'h4289b091, 32'hc198665f, 32'hc2a3e206, 32'h42705384, 32'h42738dec, 32'h421bda13, 32'hc2a3430b};
test_bias[4999:4999] = '{32'hc1d1235c};
test_output[4999:4999] = '{32'h4525e899};
end
`endif
