`ifndef RELU_BACKWARD_TEST_H
`define RELU_BACKWARD_TEST_H
reg [31:0] test_input [40000];
reg [31:0] test_output [40000];
initial begin
test_input[0:7] = '{32'hc2aa9e3b, 32'hc29ecd98, 32'h413c290a, 32'hc26338d9, 32'h4262616e, 32'h415184cf, 32'h4259a8b7, 32'h425d6264};
test_output[0:7] = '{32'h0, 32'h0, 32'h413c290a, 32'h0, 32'h4262616e, 32'h415184cf, 32'h4259a8b7, 32'h425d6264};
test_input[8:15] = '{32'hc1cff7a3, 32'h40a3448f, 32'hc218eb3b, 32'hc2a6dbdd, 32'hc18ef5ea, 32'hc1865a77, 32'h41907e01, 32'hc23b80fe};
test_output[8:15] = '{32'h0, 32'h40a3448f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41907e01, 32'h0};
test_input[16:23] = '{32'h4254a8d8, 32'h42c0c677, 32'h42a58d77, 32'h429a65a1, 32'h4110fdac, 32'hc1f10f9a, 32'hc277a7c0, 32'h4239e583};
test_output[16:23] = '{32'h4254a8d8, 32'h42c0c677, 32'h42a58d77, 32'h429a65a1, 32'h4110fdac, 32'h0, 32'h0, 32'h4239e583};
test_input[24:31] = '{32'hc1cbf83f, 32'hc26e8608, 32'hc2a0cc73, 32'hc20d7cb4, 32'h42a5a983, 32'h414df76a, 32'hc2b8584b, 32'hc2802167};
test_output[24:31] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a5a983, 32'h414df76a, 32'h0, 32'h0};
test_input[32:39] = '{32'h4292f4c9, 32'h41ec38ca, 32'h41319bd1, 32'h42793455, 32'h41b1dc0c, 32'h4285afc3, 32'hbfe28fac, 32'h4064cf6c};
test_output[32:39] = '{32'h4292f4c9, 32'h41ec38ca, 32'h41319bd1, 32'h42793455, 32'h41b1dc0c, 32'h4285afc3, 32'h0, 32'h4064cf6c};
test_input[40:47] = '{32'hc1be1d79, 32'hc1620cdc, 32'h4297ee44, 32'h42ab9ea5, 32'hc1ac1f82, 32'hc24fb63f, 32'h4270b571, 32'hc26aa4ab};
test_output[40:47] = '{32'h0, 32'h0, 32'h4297ee44, 32'h42ab9ea5, 32'h0, 32'h0, 32'h4270b571, 32'h0};
test_input[48:55] = '{32'h4057b918, 32'hc282802d, 32'hc1bac092, 32'h42b2b885, 32'hc20c0260, 32'hc26436f7, 32'hc211c5c5, 32'hc28b82d4};
test_output[48:55] = '{32'h4057b918, 32'h0, 32'h0, 32'h42b2b885, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[56:63] = '{32'hc22b111b, 32'hc17b86d2, 32'h414b8cbe, 32'h42878f82, 32'hc2043d41, 32'h41e2a73e, 32'h42a762f3, 32'hc2bbef36};
test_output[56:63] = '{32'h0, 32'h0, 32'h414b8cbe, 32'h42878f82, 32'h0, 32'h41e2a73e, 32'h42a762f3, 32'h0};
test_input[64:71] = '{32'hc2908579, 32'hc28e4536, 32'hc1c7e7a2, 32'h42a3f09f, 32'hc1d07a07, 32'hc29c70a1, 32'hc146a510, 32'h428e0417};
test_output[64:71] = '{32'h0, 32'h0, 32'h0, 32'h42a3f09f, 32'h0, 32'h0, 32'h0, 32'h428e0417};
test_input[72:79] = '{32'h42b44818, 32'hc2a56070, 32'h42abdbe7, 32'hc1f37f3a, 32'h4202f012, 32'h42a40359, 32'h42560d32, 32'h4131a01c};
test_output[72:79] = '{32'h42b44818, 32'h0, 32'h42abdbe7, 32'h0, 32'h4202f012, 32'h42a40359, 32'h42560d32, 32'h4131a01c};
test_input[80:87] = '{32'h42626601, 32'hc2b36543, 32'h41e670e1, 32'h42af3f72, 32'hc246ed80, 32'hc1530158, 32'h42ba7175, 32'hc1edee39};
test_output[80:87] = '{32'h42626601, 32'h0, 32'h41e670e1, 32'h42af3f72, 32'h0, 32'h0, 32'h42ba7175, 32'h0};
test_input[88:95] = '{32'hc2b662aa, 32'hc182312d, 32'hc1bfc27f, 32'h428f7b92, 32'hc252900f, 32'h42bce958, 32'hbeb930a4, 32'h42908127};
test_output[88:95] = '{32'h0, 32'h0, 32'h0, 32'h428f7b92, 32'h0, 32'h42bce958, 32'h0, 32'h42908127};
test_input[96:103] = '{32'h41ece1f9, 32'h3f0f0fe7, 32'hc297f6ba, 32'hc2c6785e, 32'hc2aa2a45, 32'h42a4efbb, 32'h42a97dc7, 32'h4224dbd5};
test_output[96:103] = '{32'h41ece1f9, 32'h3f0f0fe7, 32'h0, 32'h0, 32'h0, 32'h42a4efbb, 32'h42a97dc7, 32'h4224dbd5};
test_input[104:111] = '{32'h4284156d, 32'h41d1249b, 32'h4265240a, 32'h41b70b53, 32'h42171f35, 32'h4146f466, 32'h42a35443, 32'h420c930c};
test_output[104:111] = '{32'h4284156d, 32'h41d1249b, 32'h4265240a, 32'h41b70b53, 32'h42171f35, 32'h4146f466, 32'h42a35443, 32'h420c930c};
test_input[112:119] = '{32'h427b18a3, 32'h4026b437, 32'hc28d6844, 32'hc250cb25, 32'h414f5512, 32'h41e8e082, 32'hc191f30a, 32'h428a0ae0};
test_output[112:119] = '{32'h427b18a3, 32'h4026b437, 32'h0, 32'h0, 32'h414f5512, 32'h41e8e082, 32'h0, 32'h428a0ae0};
test_input[120:127] = '{32'h424e43ea, 32'hc2745f05, 32'hc1c936b3, 32'h42830cfb, 32'hc2bf7e5d, 32'hc1bd1e5a, 32'h410e77bc, 32'h4258c85b};
test_output[120:127] = '{32'h424e43ea, 32'h0, 32'h0, 32'h42830cfb, 32'h0, 32'h0, 32'h410e77bc, 32'h4258c85b};
test_input[128:135] = '{32'hc2b33754, 32'h42295c10, 32'h40ebe94d, 32'h41330ce9, 32'h428bcaa3, 32'hc0420868, 32'h40e46688, 32'hc28f0594};
test_output[128:135] = '{32'h0, 32'h42295c10, 32'h40ebe94d, 32'h41330ce9, 32'h428bcaa3, 32'h0, 32'h40e46688, 32'h0};
test_input[136:143] = '{32'hc27ec275, 32'hc29bc867, 32'h4259d663, 32'h42bc1b0a, 32'hc2c16279, 32'hc1f9fda7, 32'hc1aa0f22, 32'h41dd4b37};
test_output[136:143] = '{32'h0, 32'h0, 32'h4259d663, 32'h42bc1b0a, 32'h0, 32'h0, 32'h0, 32'h41dd4b37};
test_input[144:151] = '{32'hc218a030, 32'h4186bc8d, 32'h421f3d36, 32'h424e4c30, 32'hc2c14d86, 32'h42aa6b0c, 32'hc1f9f8a1, 32'hc22abd9b};
test_output[144:151] = '{32'h0, 32'h4186bc8d, 32'h421f3d36, 32'h424e4c30, 32'h0, 32'h42aa6b0c, 32'h0, 32'h0};
test_input[152:159] = '{32'h41f527a9, 32'hc1b0ae32, 32'h4085c07e, 32'hc1a46b8d, 32'hc25ef2a6, 32'h42b1e8e6, 32'hc1f7eb81, 32'h4288a705};
test_output[152:159] = '{32'h41f527a9, 32'h0, 32'h4085c07e, 32'h0, 32'h0, 32'h42b1e8e6, 32'h0, 32'h4288a705};
test_input[160:167] = '{32'hc2b5e281, 32'h41267fb6, 32'h42bc2e61, 32'hc2a924ef, 32'hc239d352, 32'hc10b5f39, 32'h425683a4, 32'h4261f227};
test_output[160:167] = '{32'h0, 32'h41267fb6, 32'h42bc2e61, 32'h0, 32'h0, 32'h0, 32'h425683a4, 32'h4261f227};
test_input[168:175] = '{32'h42902f40, 32'h40784bd0, 32'h4165ab51, 32'h4230666b, 32'hc2bc90f5, 32'h427fa24b, 32'hc2c48a0c, 32'hc2a87a56};
test_output[168:175] = '{32'h42902f40, 32'h40784bd0, 32'h4165ab51, 32'h4230666b, 32'h0, 32'h427fa24b, 32'h0, 32'h0};
test_input[176:183] = '{32'h41a113be, 32'h4291730b, 32'h42b113b6, 32'hc0d17a49, 32'hc23a8cb0, 32'hc172ddce, 32'h422f62c6, 32'hc1fc94a4};
test_output[176:183] = '{32'h41a113be, 32'h4291730b, 32'h42b113b6, 32'h0, 32'h0, 32'h0, 32'h422f62c6, 32'h0};
test_input[184:191] = '{32'hc1d97f87, 32'h42477287, 32'h41d48d0b, 32'h420d9f40, 32'h42935ce4, 32'h41702a83, 32'h424cda1e, 32'h40a4fe41};
test_output[184:191] = '{32'h0, 32'h42477287, 32'h41d48d0b, 32'h420d9f40, 32'h42935ce4, 32'h41702a83, 32'h424cda1e, 32'h40a4fe41};
test_input[192:199] = '{32'h421b8fa9, 32'h42b79626, 32'h42743b01, 32'hc2100ee2, 32'hc1823cb1, 32'h417222f0, 32'h42b99e92, 32'h423cb971};
test_output[192:199] = '{32'h421b8fa9, 32'h42b79626, 32'h42743b01, 32'h0, 32'h0, 32'h417222f0, 32'h42b99e92, 32'h423cb971};
test_input[200:207] = '{32'hc1f7beb1, 32'hc2894246, 32'hc28955a0, 32'h42c618f9, 32'h428f60a0, 32'h428a9143, 32'h42beaf86, 32'h41e6f67d};
test_output[200:207] = '{32'h0, 32'h0, 32'h0, 32'h42c618f9, 32'h428f60a0, 32'h428a9143, 32'h42beaf86, 32'h41e6f67d};
test_input[208:215] = '{32'hc1bba88e, 32'hc2b11498, 32'hc2b95cb4, 32'hc24232c2, 32'hc23a8eaa, 32'hc1541205, 32'h42910e13, 32'h425b77c4};
test_output[208:215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42910e13, 32'h425b77c4};
test_input[216:223] = '{32'h40ae4984, 32'hc23920f0, 32'h42a50820, 32'hc278ab86, 32'hc17cdf30, 32'h429e0cd1, 32'h421920ea, 32'h429e25a4};
test_output[216:223] = '{32'h40ae4984, 32'h0, 32'h42a50820, 32'h0, 32'h0, 32'h429e0cd1, 32'h421920ea, 32'h429e25a4};
test_input[224:231] = '{32'h42a21fac, 32'hc1f90d44, 32'hc15ae6e2, 32'hc2a8481d, 32'h42129c25, 32'hc206b595, 32'hc2a2c9e4, 32'h41d2b35d};
test_output[224:231] = '{32'h42a21fac, 32'h0, 32'h0, 32'h0, 32'h42129c25, 32'h0, 32'h0, 32'h41d2b35d};
test_input[232:239] = '{32'hc19aa1e1, 32'hc21dfc1b, 32'hc2aa9149, 32'h41b0551f, 32'h427a004d, 32'hc2970c02, 32'h40fe2bc6, 32'h4213baae};
test_output[232:239] = '{32'h0, 32'h0, 32'h0, 32'h41b0551f, 32'h427a004d, 32'h0, 32'h40fe2bc6, 32'h4213baae};
test_input[240:247] = '{32'h41a4c2be, 32'hc28ceb5f, 32'hc27aa785, 32'hc285193b, 32'h41b3e653, 32'hc006630c, 32'hc2150cbc, 32'hc280b507};
test_output[240:247] = '{32'h41a4c2be, 32'h0, 32'h0, 32'h0, 32'h41b3e653, 32'h0, 32'h0, 32'h0};
test_input[248:255] = '{32'h42c7ab35, 32'h41ed1875, 32'hc289de73, 32'h42c59e12, 32'hc195b70a, 32'h41fa8562, 32'h428c568b, 32'hc2ad779c};
test_output[248:255] = '{32'h42c7ab35, 32'h41ed1875, 32'h0, 32'h42c59e12, 32'h0, 32'h41fa8562, 32'h428c568b, 32'h0};
test_input[256:263] = '{32'hc2b26376, 32'h42821947, 32'h3c29f453, 32'hbf686431, 32'h42ab2af2, 32'hc21a8dcf, 32'hc0c30c1a, 32'hc2b88dce};
test_output[256:263] = '{32'h0, 32'h42821947, 32'h3c29f453, 32'h0, 32'h42ab2af2, 32'h0, 32'h0, 32'h0};
test_input[264:271] = '{32'h4270165a, 32'hc230e01e, 32'hc1df0ed6, 32'h429e18b7, 32'h40c04b59, 32'h42801c00, 32'h42a60af8, 32'hc2bbfac1};
test_output[264:271] = '{32'h4270165a, 32'h0, 32'h0, 32'h429e18b7, 32'h40c04b59, 32'h42801c00, 32'h42a60af8, 32'h0};
test_input[272:279] = '{32'hc2bf4db5, 32'hc20ce4e1, 32'hc184ce3a, 32'hc2759e97, 32'hc24ebf28, 32'hc2058e58, 32'h428dc2d1, 32'hc296df91};
test_output[272:279] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428dc2d1, 32'h0};
test_input[280:287] = '{32'h42ba37e8, 32'hc0969884, 32'hc285f573, 32'hc29bd632, 32'h40852593, 32'h429fd762, 32'hc1ce807d, 32'h425f4522};
test_output[280:287] = '{32'h42ba37e8, 32'h0, 32'h0, 32'h0, 32'h40852593, 32'h429fd762, 32'h0, 32'h425f4522};
test_input[288:295] = '{32'h4281b5a4, 32'h42b10b99, 32'h422a35c4, 32'h42975492, 32'h41f5d5c9, 32'hc1864295, 32'hc23c30e7, 32'hc2a0c9d7};
test_output[288:295] = '{32'h4281b5a4, 32'h42b10b99, 32'h422a35c4, 32'h42975492, 32'h41f5d5c9, 32'h0, 32'h0, 32'h0};
test_input[296:303] = '{32'h42a78afd, 32'h420532ea, 32'hc29a8621, 32'hc2aeacf3, 32'hc23e54a0, 32'hbf689c13, 32'hc2b9f3f6, 32'hc25d6334};
test_output[296:303] = '{32'h42a78afd, 32'h420532ea, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[304:311] = '{32'hc1f75f6e, 32'h425967d0, 32'hc2b3b182, 32'hc1898241, 32'h424a6476, 32'h401580db, 32'h42b3bdae, 32'h4266dd7c};
test_output[304:311] = '{32'h0, 32'h425967d0, 32'h0, 32'h0, 32'h424a6476, 32'h401580db, 32'h42b3bdae, 32'h4266dd7c};
test_input[312:319] = '{32'hc2ac3190, 32'h42a701fb, 32'h42003b1f, 32'h42c767df, 32'hc29ac175, 32'h41df788f, 32'hc262e90c, 32'h42439788};
test_output[312:319] = '{32'h0, 32'h42a701fb, 32'h42003b1f, 32'h42c767df, 32'h0, 32'h41df788f, 32'h0, 32'h42439788};
test_input[320:327] = '{32'h413fb449, 32'hbfdc93ef, 32'hc28754ac, 32'hc25db43d, 32'h413b64fb, 32'hc17d0be9, 32'h4260d166, 32'h420c87f0};
test_output[320:327] = '{32'h413fb449, 32'h0, 32'h0, 32'h0, 32'h413b64fb, 32'h0, 32'h4260d166, 32'h420c87f0};
test_input[328:335] = '{32'h4001b997, 32'h427cbf1a, 32'hc217efbc, 32'h417e5c9e, 32'hc24278d8, 32'hc1db22a6, 32'h4008855b, 32'h42bfcb0d};
test_output[328:335] = '{32'h4001b997, 32'h427cbf1a, 32'h0, 32'h417e5c9e, 32'h0, 32'h0, 32'h4008855b, 32'h42bfcb0d};
test_input[336:343] = '{32'h42a3b123, 32'hc2c0b28b, 32'hc283a924, 32'hc2acffae, 32'hc265c545, 32'hc2939f2f, 32'h42ab88a3, 32'h42713fed};
test_output[336:343] = '{32'h42a3b123, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ab88a3, 32'h42713fed};
test_input[344:351] = '{32'h42a86802, 32'h426f5d07, 32'h426d1ceb, 32'h42bb731a, 32'hc2ac2252, 32'h41749afd, 32'h427a44f6, 32'h42a0e842};
test_output[344:351] = '{32'h42a86802, 32'h426f5d07, 32'h426d1ceb, 32'h42bb731a, 32'h0, 32'h41749afd, 32'h427a44f6, 32'h42a0e842};
test_input[352:359] = '{32'hc185d0e4, 32'hc25dd38d, 32'hc2003745, 32'h426695f8, 32'hc2adfcae, 32'hc2b42c25, 32'h429cf484, 32'hc2023887};
test_output[352:359] = '{32'h0, 32'h0, 32'h0, 32'h426695f8, 32'h0, 32'h0, 32'h429cf484, 32'h0};
test_input[360:367] = '{32'hc2b85163, 32'hc14198c1, 32'h427991ae, 32'h41a8dbb7, 32'hc29ea65b, 32'hc19fa0f4, 32'h41c35b9c, 32'hc288e3b1};
test_output[360:367] = '{32'h0, 32'h0, 32'h427991ae, 32'h41a8dbb7, 32'h0, 32'h0, 32'h41c35b9c, 32'h0};
test_input[368:375] = '{32'h41a59d0e, 32'hc2801ef7, 32'h4291950e, 32'hbf3591a5, 32'h42b605f7, 32'h42a3f23f, 32'h4281b63d, 32'h41e5ea37};
test_output[368:375] = '{32'h41a59d0e, 32'h0, 32'h4291950e, 32'h0, 32'h42b605f7, 32'h42a3f23f, 32'h4281b63d, 32'h41e5ea37};
test_input[376:383] = '{32'hc25a977c, 32'h42c113f3, 32'hc2ace622, 32'h4244c43a, 32'h414eefe2, 32'h423b0224, 32'hc285b74b, 32'hc1af5388};
test_output[376:383] = '{32'h0, 32'h42c113f3, 32'h0, 32'h4244c43a, 32'h414eefe2, 32'h423b0224, 32'h0, 32'h0};
test_input[384:391] = '{32'h423edbcd, 32'hc257bf6b, 32'hc234c1db, 32'h42a1806e, 32'h4207deb0, 32'h4229bfaa, 32'hc2ac778c, 32'hc1d9eebc};
test_output[384:391] = '{32'h423edbcd, 32'h0, 32'h0, 32'h42a1806e, 32'h4207deb0, 32'h4229bfaa, 32'h0, 32'h0};
test_input[392:399] = '{32'h424901ed, 32'h418fd37b, 32'hc09d799b, 32'h429693fd, 32'hc220c4ec, 32'h4243d11f, 32'hc22ee56d, 32'hc272a99b};
test_output[392:399] = '{32'h424901ed, 32'h418fd37b, 32'h0, 32'h429693fd, 32'h0, 32'h4243d11f, 32'h0, 32'h0};
test_input[400:407] = '{32'h41237ffb, 32'h4249489d, 32'hc21ff29c, 32'h42be218f, 32'hc28c3e1b, 32'h42bdbe13, 32'hc28768a5, 32'hc1db990e};
test_output[400:407] = '{32'h41237ffb, 32'h4249489d, 32'h0, 32'h42be218f, 32'h0, 32'h42bdbe13, 32'h0, 32'h0};
test_input[408:415] = '{32'h4298cd08, 32'h426751ed, 32'h41971b12, 32'h422c6333, 32'h4217f0bc, 32'h4251c54c, 32'h4161627a, 32'hc2c54b3f};
test_output[408:415] = '{32'h4298cd08, 32'h426751ed, 32'h41971b12, 32'h422c6333, 32'h4217f0bc, 32'h4251c54c, 32'h4161627a, 32'h0};
test_input[416:423] = '{32'hc25862c2, 32'hc18c78fb, 32'hc2837d59, 32'h418d4b6e, 32'h4196f8bf, 32'h42b3b42c, 32'hc2bd3d33, 32'hc2650635};
test_output[416:423] = '{32'h0, 32'h0, 32'h0, 32'h418d4b6e, 32'h4196f8bf, 32'h42b3b42c, 32'h0, 32'h0};
test_input[424:431] = '{32'hc25c6a9b, 32'h42b00cc9, 32'h411854f3, 32'h420f0ac9, 32'hc21cd78e, 32'hc2bc17d6, 32'h428126c1, 32'hc2aa025b};
test_output[424:431] = '{32'h0, 32'h42b00cc9, 32'h411854f3, 32'h420f0ac9, 32'h0, 32'h0, 32'h428126c1, 32'h0};
test_input[432:439] = '{32'hc23ea219, 32'hc2ab2975, 32'h41a98a82, 32'h423c9953, 32'h42699572, 32'h41a863f8, 32'h426d9990, 32'hc1ebee53};
test_output[432:439] = '{32'h0, 32'h0, 32'h41a98a82, 32'h423c9953, 32'h42699572, 32'h41a863f8, 32'h426d9990, 32'h0};
test_input[440:447] = '{32'hc281b9f8, 32'h429c2015, 32'h4118f676, 32'hc195770a, 32'hc1cd081c, 32'h426c49a0, 32'h42bebbd2, 32'hc1c695d0};
test_output[440:447] = '{32'h0, 32'h429c2015, 32'h4118f676, 32'h0, 32'h0, 32'h426c49a0, 32'h42bebbd2, 32'h0};
test_input[448:455] = '{32'h4295b8cc, 32'h42bd772e, 32'h3fee3d48, 32'h4292ff52, 32'h423f2275, 32'hc1ece1bc, 32'hc28737f0, 32'h42aa1426};
test_output[448:455] = '{32'h4295b8cc, 32'h42bd772e, 32'h3fee3d48, 32'h4292ff52, 32'h423f2275, 32'h0, 32'h0, 32'h42aa1426};
test_input[456:463] = '{32'hc1cb0eb0, 32'h4232104b, 32'h426219cc, 32'h411ce222, 32'h4252753c, 32'h428628ea, 32'h423ae094, 32'h42a0f74f};
test_output[456:463] = '{32'h0, 32'h4232104b, 32'h426219cc, 32'h411ce222, 32'h4252753c, 32'h428628ea, 32'h423ae094, 32'h42a0f74f};
test_input[464:471] = '{32'hc22c4ab0, 32'h42b5e77f, 32'h410b24fa, 32'h4287dc70, 32'hc25264c7, 32'hc232f6a6, 32'hc19e0f13, 32'hc2c358ee};
test_output[464:471] = '{32'h0, 32'h42b5e77f, 32'h410b24fa, 32'h4287dc70, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[472:479] = '{32'h41d5ac62, 32'hc2241377, 32'hc21f4acb, 32'hc2b45799, 32'hc2968d86, 32'h425ff225, 32'h42c22911, 32'h42141c4b};
test_output[472:479] = '{32'h41d5ac62, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425ff225, 32'h42c22911, 32'h42141c4b};
test_input[480:487] = '{32'hc29e496d, 32'h428a32dc, 32'h421a5870, 32'hc223019d, 32'hc28d5736, 32'h4215f996, 32'hc2c1cd85, 32'hc23990f0};
test_output[480:487] = '{32'h0, 32'h428a32dc, 32'h421a5870, 32'h0, 32'h0, 32'h4215f996, 32'h0, 32'h0};
test_input[488:495] = '{32'hc2169d14, 32'h41a94804, 32'hc265b235, 32'hc25664c7, 32'hc11ba843, 32'hc2898756, 32'h42ad1f5b, 32'hc1d76e83};
test_output[488:495] = '{32'h0, 32'h41a94804, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ad1f5b, 32'h0};
test_input[496:503] = '{32'h420076ef, 32'hc2654539, 32'hc286e008, 32'h4227582e, 32'h41bcdea7, 32'hc2872960, 32'h42c1d2fe, 32'h4261f6ec};
test_output[496:503] = '{32'h420076ef, 32'h0, 32'h0, 32'h4227582e, 32'h41bcdea7, 32'h0, 32'h42c1d2fe, 32'h4261f6ec};
test_input[504:511] = '{32'hc2562bf7, 32'hc281fc0d, 32'hc1a30dc6, 32'h404b8f5b, 32'hc2ac8dd6, 32'hc2b178ca, 32'h4261f2cb, 32'hc1b0730d};
test_output[504:511] = '{32'h0, 32'h0, 32'h0, 32'h404b8f5b, 32'h0, 32'h0, 32'h4261f2cb, 32'h0};
test_input[512:519] = '{32'h42371237, 32'h42a140a6, 32'h42349225, 32'hc25b463f, 32'h40439ca8, 32'h42abfcb2, 32'hc230d2cd, 32'hc2c603fb};
test_output[512:519] = '{32'h42371237, 32'h42a140a6, 32'h42349225, 32'h0, 32'h40439ca8, 32'h42abfcb2, 32'h0, 32'h0};
test_input[520:527] = '{32'h42c105b7, 32'h42c571ab, 32'hc297979e, 32'h41c626d1, 32'h41d88d5d, 32'h41a28e04, 32'hc049f74d, 32'h4266ae86};
test_output[520:527] = '{32'h42c105b7, 32'h42c571ab, 32'h0, 32'h41c626d1, 32'h41d88d5d, 32'h41a28e04, 32'h0, 32'h4266ae86};
test_input[528:535] = '{32'h41c65b2f, 32'h42229802, 32'h410c2ec3, 32'hc2c6cc7b, 32'hc29d2d79, 32'h3e913020, 32'h42aaaf84, 32'h42a61dcc};
test_output[528:535] = '{32'h41c65b2f, 32'h42229802, 32'h410c2ec3, 32'h0, 32'h0, 32'h3e913020, 32'h42aaaf84, 32'h42a61dcc};
test_input[536:543] = '{32'hc01f9712, 32'h4253de9b, 32'hbfce53dc, 32'h4078a3ee, 32'h4239a613, 32'h41265326, 32'hc060ff1e, 32'hc2bad15f};
test_output[536:543] = '{32'h0, 32'h4253de9b, 32'h0, 32'h4078a3ee, 32'h4239a613, 32'h41265326, 32'h0, 32'h0};
test_input[544:551] = '{32'h4220deba, 32'hc02f6e9c, 32'hc2a95457, 32'hc299f8cd, 32'hc1b1cad4, 32'h42654450, 32'hc27b578b, 32'h42785b98};
test_output[544:551] = '{32'h4220deba, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42654450, 32'h0, 32'h42785b98};
test_input[552:559] = '{32'hc2ba181c, 32'hc2a8270f, 32'hc1b26e00, 32'h4160011d, 32'hc2bca110, 32'hc2025f4d, 32'hc255a627, 32'h41de8cb8};
test_output[552:559] = '{32'h0, 32'h0, 32'h0, 32'h4160011d, 32'h0, 32'h0, 32'h0, 32'h41de8cb8};
test_input[560:567] = '{32'h41be4357, 32'h415cf364, 32'h426e1451, 32'hc23409de, 32'h4215b4a5, 32'hc227ab11, 32'h428500ff, 32'h428e4ea9};
test_output[560:567] = '{32'h41be4357, 32'h415cf364, 32'h426e1451, 32'h0, 32'h4215b4a5, 32'h0, 32'h428500ff, 32'h428e4ea9};
test_input[568:575] = '{32'h42667b54, 32'hc292e975, 32'hc26cb216, 32'hc224b5d5, 32'h418d5cab, 32'hc2c70be5, 32'hc2a52bf2, 32'h42a11f15};
test_output[568:575] = '{32'h42667b54, 32'h0, 32'h0, 32'h0, 32'h418d5cab, 32'h0, 32'h0, 32'h42a11f15};
test_input[576:583] = '{32'hc2a81502, 32'hc293bbf1, 32'hc0cb6264, 32'h411220b4, 32'hc28c8534, 32'hc22ed2d2, 32'h42559117, 32'h41d4803c};
test_output[576:583] = '{32'h0, 32'h0, 32'h0, 32'h411220b4, 32'h0, 32'h0, 32'h42559117, 32'h41d4803c};
test_input[584:591] = '{32'h42b8071c, 32'h42c42afa, 32'h428ba01a, 32'hc2115d51, 32'hc281fafb, 32'h3ea2931a, 32'hc2a998ba, 32'h429d8fcf};
test_output[584:591] = '{32'h42b8071c, 32'h42c42afa, 32'h428ba01a, 32'h0, 32'h0, 32'h3ea2931a, 32'h0, 32'h429d8fcf};
test_input[592:599] = '{32'h40f9a081, 32'hc1ffb83f, 32'hc2be7292, 32'h416d88a5, 32'h40c0dcd2, 32'h4286f97a, 32'h4275d120, 32'h41f36cfe};
test_output[592:599] = '{32'h40f9a081, 32'h0, 32'h0, 32'h416d88a5, 32'h40c0dcd2, 32'h4286f97a, 32'h4275d120, 32'h41f36cfe};
test_input[600:607] = '{32'h41949a79, 32'h428a4bdf, 32'h42b85170, 32'h42c19bd7, 32'hc24c6228, 32'h42b3a32e, 32'hc29f1650, 32'hc20d50f8};
test_output[600:607] = '{32'h41949a79, 32'h428a4bdf, 32'h42b85170, 32'h42c19bd7, 32'h0, 32'h42b3a32e, 32'h0, 32'h0};
test_input[608:615] = '{32'hc273726e, 32'hc2c0b6c0, 32'h429bcdee, 32'hc194d549, 32'h422b50bb, 32'h42a9b175, 32'hc27942f0, 32'hc1423f57};
test_output[608:615] = '{32'h0, 32'h0, 32'h429bcdee, 32'h0, 32'h422b50bb, 32'h42a9b175, 32'h0, 32'h0};
test_input[616:623] = '{32'hc203164c, 32'hc2a95033, 32'h40f2a7c3, 32'hc1b179ff, 32'h4287826b, 32'h41028ef0, 32'hc20a80d1, 32'hc28cdb1d};
test_output[616:623] = '{32'h0, 32'h0, 32'h40f2a7c3, 32'h0, 32'h4287826b, 32'h41028ef0, 32'h0, 32'h0};
test_input[624:631] = '{32'hc1c126c3, 32'hc24901f3, 32'hc1f4169c, 32'h425b4254, 32'h42b777c3, 32'hc28db9c5, 32'h40775069, 32'h426952fb};
test_output[624:631] = '{32'h0, 32'h0, 32'h0, 32'h425b4254, 32'h42b777c3, 32'h0, 32'h40775069, 32'h426952fb};
test_input[632:639] = '{32'hc2651020, 32'h41ee8f57, 32'h428861c8, 32'hc1d92ac4, 32'hc2adf545, 32'hc27aa74a, 32'h42b3c0db, 32'hc2bae340};
test_output[632:639] = '{32'h0, 32'h41ee8f57, 32'h428861c8, 32'h0, 32'h0, 32'h0, 32'h42b3c0db, 32'h0};
test_input[640:647] = '{32'h4247660c, 32'h423bb1eb, 32'hc1e1f07f, 32'h41be189e, 32'h429d323c, 32'h42a8c775, 32'hc29bf2d9, 32'hc27ead09};
test_output[640:647] = '{32'h4247660c, 32'h423bb1eb, 32'h0, 32'h41be189e, 32'h429d323c, 32'h42a8c775, 32'h0, 32'h0};
test_input[648:655] = '{32'hc23d16e1, 32'h41611119, 32'h4238654e, 32'hc2928705, 32'hc2175cab, 32'hc241e5e5, 32'hc12e92d2, 32'h42897ae6};
test_output[648:655] = '{32'h0, 32'h41611119, 32'h4238654e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42897ae6};
test_input[656:663] = '{32'hc2a82304, 32'h423020dd, 32'h419d4448, 32'hc282685d, 32'hc18fab82, 32'hc2b67d89, 32'h42151176, 32'hc151257f};
test_output[656:663] = '{32'h0, 32'h423020dd, 32'h419d4448, 32'h0, 32'h0, 32'h0, 32'h42151176, 32'h0};
test_input[664:671] = '{32'hc1860a51, 32'h41e8fb95, 32'h4225b1c3, 32'hc287bcde, 32'h4275135e, 32'hc2c506b6, 32'h4235ca7b, 32'h41360a43};
test_output[664:671] = '{32'h0, 32'h41e8fb95, 32'h4225b1c3, 32'h0, 32'h4275135e, 32'h0, 32'h4235ca7b, 32'h41360a43};
test_input[672:679] = '{32'h42a02249, 32'h4191ec05, 32'h41bfd341, 32'hc0d3ef1c, 32'hc21874a8, 32'hc2bd95f9, 32'hc2424d3a, 32'h4218f574};
test_output[672:679] = '{32'h42a02249, 32'h4191ec05, 32'h41bfd341, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4218f574};
test_input[680:687] = '{32'hc23a7207, 32'hc1ae246e, 32'hc2ae2974, 32'hc217c5fa, 32'hc23df11e, 32'h42bf1932, 32'h42a144e8, 32'hc29be6ac};
test_output[680:687] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bf1932, 32'h42a144e8, 32'h0};
test_input[688:695] = '{32'hbe4d30d3, 32'hc2ba5aaf, 32'h42957238, 32'hbd23ac14, 32'h42563a6d, 32'hc15629ed, 32'h409f2928, 32'h41125277};
test_output[688:695] = '{32'h0, 32'h0, 32'h42957238, 32'h0, 32'h42563a6d, 32'h0, 32'h409f2928, 32'h41125277};
test_input[696:703] = '{32'h40cb619a, 32'hc28d61c9, 32'h42c64930, 32'h41153f8c, 32'h4216b73b, 32'h4028724a, 32'hc22de293, 32'h420874b3};
test_output[696:703] = '{32'h40cb619a, 32'h0, 32'h42c64930, 32'h41153f8c, 32'h4216b73b, 32'h4028724a, 32'h0, 32'h420874b3};
test_input[704:711] = '{32'hc26a498b, 32'hc181307e, 32'hc27eb7d8, 32'h42463e14, 32'hbf78e833, 32'h41860bbd, 32'hc284a223, 32'h42a692e0};
test_output[704:711] = '{32'h0, 32'h0, 32'h0, 32'h42463e14, 32'h0, 32'h41860bbd, 32'h0, 32'h42a692e0};
test_input[712:719] = '{32'hc2667d42, 32'h421133e8, 32'h429ee74c, 32'h423c2bcf, 32'h426a0a25, 32'h41cfef06, 32'h40a764a8, 32'hc2a93885};
test_output[712:719] = '{32'h0, 32'h421133e8, 32'h429ee74c, 32'h423c2bcf, 32'h426a0a25, 32'h41cfef06, 32'h40a764a8, 32'h0};
test_input[720:727] = '{32'h429bd78d, 32'hc2807f9d, 32'h422fd05a, 32'hc295669a, 32'hc2468170, 32'h422f3f33, 32'h42198282, 32'h41f41a87};
test_output[720:727] = '{32'h429bd78d, 32'h0, 32'h422fd05a, 32'h0, 32'h0, 32'h422f3f33, 32'h42198282, 32'h41f41a87};
test_input[728:735] = '{32'hc2934e20, 32'hc1c15838, 32'hc14d989d, 32'hc2896a28, 32'h41b3cb40, 32'hc1ffd129, 32'h429267cb, 32'h428b8b4a};
test_output[728:735] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41b3cb40, 32'h0, 32'h429267cb, 32'h428b8b4a};
test_input[736:743] = '{32'hc09b2e01, 32'h42bdfe16, 32'h4261832a, 32'hc2a48d50, 32'hc2c39e7a, 32'h3f9671aa, 32'hc1c2279e, 32'hc2204b6f};
test_output[736:743] = '{32'h0, 32'h42bdfe16, 32'h4261832a, 32'h0, 32'h0, 32'h3f9671aa, 32'h0, 32'h0};
test_input[744:751] = '{32'hc21a2390, 32'h42bb2997, 32'h40f3bb3d, 32'h42078fb7, 32'hc1a9a90e, 32'hc0374bb6, 32'h42aeb78b, 32'h4210d9f4};
test_output[744:751] = '{32'h0, 32'h42bb2997, 32'h40f3bb3d, 32'h42078fb7, 32'h0, 32'h0, 32'h42aeb78b, 32'h4210d9f4};
test_input[752:759] = '{32'hc18802d9, 32'hc2269064, 32'h426a4ef2, 32'hc2084dad, 32'h42bd7dec, 32'hc23026cb, 32'h429a15b0, 32'h4234d29b};
test_output[752:759] = '{32'h0, 32'h0, 32'h426a4ef2, 32'h0, 32'h42bd7dec, 32'h0, 32'h429a15b0, 32'h4234d29b};
test_input[760:767] = '{32'hc198682a, 32'h429db1cd, 32'hc169bf04, 32'h41dab148, 32'hc21859da, 32'h429b162c, 32'h42b5dd18, 32'h4295ac46};
test_output[760:767] = '{32'h0, 32'h429db1cd, 32'h0, 32'h41dab148, 32'h0, 32'h429b162c, 32'h42b5dd18, 32'h4295ac46};
test_input[768:775] = '{32'h426965d9, 32'hc27cc2a2, 32'hc1c76751, 32'h42b5cdba, 32'hc2877429, 32'hc23bc460, 32'hc28f4d14, 32'h425f6815};
test_output[768:775] = '{32'h426965d9, 32'h0, 32'h0, 32'h42b5cdba, 32'h0, 32'h0, 32'h0, 32'h425f6815};
test_input[776:783] = '{32'hc08ebafa, 32'hc26e1c77, 32'h427fcb5b, 32'h429dd50e, 32'hc29414d5, 32'hc2ac79bc, 32'h42783f03, 32'hc0dc7ea5};
test_output[776:783] = '{32'h0, 32'h0, 32'h427fcb5b, 32'h429dd50e, 32'h0, 32'h0, 32'h42783f03, 32'h0};
test_input[784:791] = '{32'hc289a88e, 32'h42bcd4a8, 32'hc1892313, 32'h41a7c120, 32'h4189634c, 32'h41296818, 32'hc21fee4a, 32'hc212aa7e};
test_output[784:791] = '{32'h0, 32'h42bcd4a8, 32'h0, 32'h41a7c120, 32'h4189634c, 32'h41296818, 32'h0, 32'h0};
test_input[792:799] = '{32'hc18e4260, 32'hc19f9499, 32'hc1e8c9b3, 32'hc2a901ae, 32'h42197400, 32'hc22dd673, 32'hc28424cf, 32'h41e48fb1};
test_output[792:799] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42197400, 32'h0, 32'h0, 32'h41e48fb1};
test_input[800:807] = '{32'hc2b68916, 32'h414c477f, 32'hc26f4fa5, 32'hc193de14, 32'hc2859821, 32'hbf66e474, 32'hc211f0d3, 32'h4211c232};
test_output[800:807] = '{32'h0, 32'h414c477f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4211c232};
test_input[808:815] = '{32'hc0036c83, 32'h41ce7034, 32'hc29c3f81, 32'hc1d972ce, 32'h42961c25, 32'h40100884, 32'h42b91ca8, 32'h418d462b};
test_output[808:815] = '{32'h0, 32'h41ce7034, 32'h0, 32'h0, 32'h42961c25, 32'h40100884, 32'h42b91ca8, 32'h418d462b};
test_input[816:823] = '{32'hc1e7efe7, 32'hc2a66e24, 32'h423becb6, 32'hc2b08624, 32'hc248bb77, 32'h41d4d1d2, 32'hc2278296, 32'hc2a4dfa3};
test_output[816:823] = '{32'h0, 32'h0, 32'h423becb6, 32'h0, 32'h0, 32'h41d4d1d2, 32'h0, 32'h0};
test_input[824:831] = '{32'h42bbb923, 32'h420692f6, 32'hc20ee53f, 32'h41d16c15, 32'h41e959b2, 32'h428a1374, 32'hc2780213, 32'hc297aa19};
test_output[824:831] = '{32'h42bbb923, 32'h420692f6, 32'h0, 32'h41d16c15, 32'h41e959b2, 32'h428a1374, 32'h0, 32'h0};
test_input[832:839] = '{32'hc298248a, 32'hc22f20f4, 32'hc229b6ae, 32'hc24b0451, 32'h42b36c17, 32'hc1b7f811, 32'hc21f4361, 32'h427e1a0c};
test_output[832:839] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42b36c17, 32'h0, 32'h0, 32'h427e1a0c};
test_input[840:847] = '{32'hc292caf4, 32'h424ac2b8, 32'h429fa468, 32'hc2aa34fb, 32'h41657dbd, 32'h42821031, 32'h41171684, 32'h419473b1};
test_output[840:847] = '{32'h0, 32'h424ac2b8, 32'h429fa468, 32'h0, 32'h41657dbd, 32'h42821031, 32'h41171684, 32'h419473b1};
test_input[848:855] = '{32'hc2647335, 32'hc281cdda, 32'hc2b24508, 32'h3dd10245, 32'h428eca2e, 32'hc21dee76, 32'hc29ff40c, 32'h409def7f};
test_output[848:855] = '{32'h0, 32'h0, 32'h0, 32'h3dd10245, 32'h428eca2e, 32'h0, 32'h0, 32'h409def7f};
test_input[856:863] = '{32'hc2260ddc, 32'hc19e2f0c, 32'hc2182eeb, 32'h4207aa8c, 32'hc2699613, 32'hc226e956, 32'hc2bb6667, 32'h42ac05cd};
test_output[856:863] = '{32'h0, 32'h0, 32'h0, 32'h4207aa8c, 32'h0, 32'h0, 32'h0, 32'h42ac05cd};
test_input[864:871] = '{32'h42b5de97, 32'h42b1ae63, 32'h4283475a, 32'hc21b5457, 32'hc157cfce, 32'hc266bc30, 32'h419e835b, 32'hc1ff6013};
test_output[864:871] = '{32'h42b5de97, 32'h42b1ae63, 32'h4283475a, 32'h0, 32'h0, 32'h0, 32'h419e835b, 32'h0};
test_input[872:879] = '{32'hc29d3e77, 32'hc240c35c, 32'h41aa412c, 32'h421d37cd, 32'hc2165564, 32'h4215434d, 32'hc1716be4, 32'hc1e5dd27};
test_output[872:879] = '{32'h0, 32'h0, 32'h41aa412c, 32'h421d37cd, 32'h0, 32'h4215434d, 32'h0, 32'h0};
test_input[880:887] = '{32'hc13547d8, 32'hc2a34560, 32'hc23dad1d, 32'hc2b4104a, 32'h429988db, 32'hc29531ef, 32'h422c3940, 32'h428b121c};
test_output[880:887] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429988db, 32'h0, 32'h422c3940, 32'h428b121c};
test_input[888:895] = '{32'hc23c7fe4, 32'h42716445, 32'hc2859c3b, 32'h41e238c0, 32'hc1dd2f69, 32'hc261f42c, 32'hc2c3c928, 32'h4249070a};
test_output[888:895] = '{32'h0, 32'h42716445, 32'h0, 32'h41e238c0, 32'h0, 32'h0, 32'h0, 32'h4249070a};
test_input[896:903] = '{32'h4239d6a3, 32'hc292a840, 32'hc25c9f47, 32'h42b99393, 32'h42b43a2b, 32'hc09ce125, 32'hc2313be5, 32'h42c06446};
test_output[896:903] = '{32'h4239d6a3, 32'h0, 32'h0, 32'h42b99393, 32'h42b43a2b, 32'h0, 32'h0, 32'h42c06446};
test_input[904:911] = '{32'hc2b8eace, 32'h41e790f9, 32'h4268e489, 32'h41c37eec, 32'h41d80f23, 32'hc25047af, 32'h4117fada, 32'h427ca390};
test_output[904:911] = '{32'h0, 32'h41e790f9, 32'h4268e489, 32'h41c37eec, 32'h41d80f23, 32'h0, 32'h4117fada, 32'h427ca390};
test_input[912:919] = '{32'hc212d1fc, 32'h425823d8, 32'hc28c7a04, 32'hc1f3a383, 32'h420ca9ee, 32'h428f63da, 32'h4238b3d9, 32'hc26f37ef};
test_output[912:919] = '{32'h0, 32'h425823d8, 32'h0, 32'h0, 32'h420ca9ee, 32'h428f63da, 32'h4238b3d9, 32'h0};
test_input[920:927] = '{32'h4249e992, 32'h428b7505, 32'h3fd63bff, 32'h3f2ce973, 32'hc24ee77a, 32'hc2a9ec44, 32'hc2c7d92a, 32'h4297e03f};
test_output[920:927] = '{32'h4249e992, 32'h428b7505, 32'h3fd63bff, 32'h3f2ce973, 32'h0, 32'h0, 32'h0, 32'h4297e03f};
test_input[928:935] = '{32'h4239b4d5, 32'h421792da, 32'h425ad132, 32'h41ea8d28, 32'h4229a8ef, 32'hc256c6c3, 32'h429364d5, 32'h42b9e817};
test_output[928:935] = '{32'h4239b4d5, 32'h421792da, 32'h425ad132, 32'h41ea8d28, 32'h4229a8ef, 32'h0, 32'h429364d5, 32'h42b9e817};
test_input[936:943] = '{32'hc0fc2332, 32'h42bb4568, 32'h3ff5d5f8, 32'hc2bb3b6b, 32'hc1eb15f0, 32'hc24e5d7f, 32'hc26c0545, 32'h425664b8};
test_output[936:943] = '{32'h0, 32'h42bb4568, 32'h3ff5d5f8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425664b8};
test_input[944:951] = '{32'h4282da67, 32'hc2626904, 32'hc1146324, 32'hc295df96, 32'h41a15f4f, 32'hc2b143f5, 32'hc289752e, 32'h42a86bcf};
test_output[944:951] = '{32'h4282da67, 32'h0, 32'h0, 32'h0, 32'h41a15f4f, 32'h0, 32'h0, 32'h42a86bcf};
test_input[952:959] = '{32'h41bf090d, 32'h42c4b4c2, 32'h400c15ca, 32'hc26f927a, 32'hc201c74c, 32'h420efd6a, 32'hc20e2b9f, 32'h41f7eb7b};
test_output[952:959] = '{32'h41bf090d, 32'h42c4b4c2, 32'h400c15ca, 32'h0, 32'h0, 32'h420efd6a, 32'h0, 32'h41f7eb7b};
test_input[960:967] = '{32'hc1888025, 32'hc24cefdd, 32'hc23a1d5f, 32'hc1ae081c, 32'h41e0eb4c, 32'h428e530d, 32'h4252b771, 32'h426d8e2d};
test_output[960:967] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41e0eb4c, 32'h428e530d, 32'h4252b771, 32'h426d8e2d};
test_input[968:975] = '{32'h42c53549, 32'h421e63a8, 32'h42756344, 32'h429c6486, 32'h421b2bab, 32'h42b58355, 32'hc24baa08, 32'h422a0598};
test_output[968:975] = '{32'h42c53549, 32'h421e63a8, 32'h42756344, 32'h429c6486, 32'h421b2bab, 32'h42b58355, 32'h0, 32'h422a0598};
test_input[976:983] = '{32'hc052d856, 32'hc2b775b4, 32'hc2c5937b, 32'hc1e2e3f2, 32'hc06e616b, 32'h41a73735, 32'hc186aeff, 32'h426695de};
test_output[976:983] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41a73735, 32'h0, 32'h426695de};
test_input[984:991] = '{32'hc287b57d, 32'h4203d191, 32'hc2bc2f9d, 32'h42810342, 32'hc22518dc, 32'h42c199ac, 32'h418775d4, 32'h41484aae};
test_output[984:991] = '{32'h0, 32'h4203d191, 32'h0, 32'h42810342, 32'h0, 32'h42c199ac, 32'h418775d4, 32'h41484aae};
test_input[992:999] = '{32'h428bed88, 32'h42885c3a, 32'h41bf0a45, 32'hc21b7cb3, 32'h42ac8b6b, 32'hc20bde31, 32'h42a71a7b, 32'h4211eb09};
test_output[992:999] = '{32'h428bed88, 32'h42885c3a, 32'h41bf0a45, 32'h0, 32'h42ac8b6b, 32'h0, 32'h42a71a7b, 32'h4211eb09};
test_input[1000:1007] = '{32'hc1c2b8d4, 32'h41073999, 32'hc28c9700, 32'h4215a32b, 32'hc1992a31, 32'hc05ae673, 32'hc0f4bb07, 32'h42acfd24};
test_output[1000:1007] = '{32'h0, 32'h41073999, 32'h0, 32'h4215a32b, 32'h0, 32'h0, 32'h0, 32'h42acfd24};
test_input[1008:1015] = '{32'h42bdc735, 32'hc1aa379d, 32'h423949b9, 32'h40cf884e, 32'h4286b120, 32'h427f5948, 32'h3f53e7e5, 32'h4187d8d8};
test_output[1008:1015] = '{32'h42bdc735, 32'h0, 32'h423949b9, 32'h40cf884e, 32'h4286b120, 32'h427f5948, 32'h3f53e7e5, 32'h4187d8d8};
test_input[1016:1023] = '{32'hc20b2714, 32'hc2b3cfcf, 32'h4281e3fd, 32'h42530f72, 32'hc2bd0d14, 32'hc2041484, 32'hc2c34bbd, 32'h41a42bbe};
test_output[1016:1023] = '{32'h0, 32'h0, 32'h4281e3fd, 32'h42530f72, 32'h0, 32'h0, 32'h0, 32'h41a42bbe};
test_input[1024:1031] = '{32'hc2886be9, 32'h4158a8df, 32'h4280b73a, 32'hc298f991, 32'hc28afc77, 32'hc13ee71e, 32'h429d9fe4, 32'h4293b450};
test_output[1024:1031] = '{32'h0, 32'h4158a8df, 32'h4280b73a, 32'h0, 32'h0, 32'h0, 32'h429d9fe4, 32'h4293b450};
test_input[1032:1039] = '{32'hc17ed412, 32'h424da220, 32'h4221e2e2, 32'hc237a641, 32'hc25e47d9, 32'h42a9cee0, 32'h409743ff, 32'hc298c3af};
test_output[1032:1039] = '{32'h0, 32'h424da220, 32'h4221e2e2, 32'h0, 32'h0, 32'h42a9cee0, 32'h409743ff, 32'h0};
test_input[1040:1047] = '{32'h42b33a4c, 32'hc2873827, 32'h41d21ed6, 32'h4293bd39, 32'h42b387c7, 32'hc252d4dc, 32'hc29a273c, 32'hc221795a};
test_output[1040:1047] = '{32'h42b33a4c, 32'h0, 32'h41d21ed6, 32'h4293bd39, 32'h42b387c7, 32'h0, 32'h0, 32'h0};
test_input[1048:1055] = '{32'h4195ddfc, 32'hc26809c9, 32'hc1e78ab9, 32'h42597168, 32'h41a4c520, 32'h4216f05d, 32'hc2837d86, 32'hc25c336a};
test_output[1048:1055] = '{32'h4195ddfc, 32'h0, 32'h0, 32'h42597168, 32'h41a4c520, 32'h4216f05d, 32'h0, 32'h0};
test_input[1056:1063] = '{32'h42091a4c, 32'hc2b2f4a9, 32'h426d5595, 32'hc28d4ccc, 32'h41ffc7b1, 32'h41867eb6, 32'hc2987155, 32'h41047122};
test_output[1056:1063] = '{32'h42091a4c, 32'h0, 32'h426d5595, 32'h0, 32'h41ffc7b1, 32'h41867eb6, 32'h0, 32'h41047122};
test_input[1064:1071] = '{32'hc29301da, 32'hc291c568, 32'hc29ea864, 32'h42af1065, 32'hc2a1f81d, 32'h42491b92, 32'h412a2ebc, 32'h3fb96890};
test_output[1064:1071] = '{32'h0, 32'h0, 32'h0, 32'h42af1065, 32'h0, 32'h42491b92, 32'h412a2ebc, 32'h3fb96890};
test_input[1072:1079] = '{32'h42b06bc5, 32'h415de815, 32'hc2321228, 32'h419518f1, 32'hc1baf21d, 32'hc214461b, 32'h41dc3a7e, 32'hc23b488c};
test_output[1072:1079] = '{32'h42b06bc5, 32'h415de815, 32'h0, 32'h419518f1, 32'h0, 32'h0, 32'h41dc3a7e, 32'h0};
test_input[1080:1087] = '{32'h409f0f8b, 32'h422bc23e, 32'hc23486b3, 32'hc2402c34, 32'h42c5e44e, 32'hc24d8bfc, 32'hc23081e4, 32'hc20d5731};
test_output[1080:1087] = '{32'h409f0f8b, 32'h422bc23e, 32'h0, 32'h0, 32'h42c5e44e, 32'h0, 32'h0, 32'h0};
test_input[1088:1095] = '{32'h42416dc4, 32'hc2b70c8a, 32'h42b0c8df, 32'h42bf4610, 32'hc1893822, 32'h42aaf3ca, 32'h4283c85c, 32'h42afe2fa};
test_output[1088:1095] = '{32'h42416dc4, 32'h0, 32'h42b0c8df, 32'h42bf4610, 32'h0, 32'h42aaf3ca, 32'h4283c85c, 32'h42afe2fa};
test_input[1096:1103] = '{32'hc2aa8046, 32'hbf80f233, 32'hc206bbae, 32'h4256975d, 32'hc125f88a, 32'h42c4be5f, 32'hc2c12ede, 32'hc101d5a5};
test_output[1096:1103] = '{32'h0, 32'h0, 32'h0, 32'h4256975d, 32'h0, 32'h42c4be5f, 32'h0, 32'h0};
test_input[1104:1111] = '{32'hc2b9582c, 32'hc224802b, 32'hc2b2247a, 32'hc209b6ea, 32'h42c1fb52, 32'hbf073716, 32'hc1b1a953, 32'hc25a7996};
test_output[1104:1111] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42c1fb52, 32'h0, 32'h0, 32'h0};
test_input[1112:1119] = '{32'h42b3c0c2, 32'hc233ab85, 32'hc288beff, 32'hc29f4f02, 32'h41a82ef2, 32'h4294eafa, 32'h422d44db, 32'hc1a1e91e};
test_output[1112:1119] = '{32'h42b3c0c2, 32'h0, 32'h0, 32'h0, 32'h41a82ef2, 32'h4294eafa, 32'h422d44db, 32'h0};
test_input[1120:1127] = '{32'h428aa01b, 32'h424ba5a7, 32'h42486e65, 32'hc2837d42, 32'h423d98b8, 32'hc1dc6b10, 32'hc2a68c62, 32'h42745dba};
test_output[1120:1127] = '{32'h428aa01b, 32'h424ba5a7, 32'h42486e65, 32'h0, 32'h423d98b8, 32'h0, 32'h0, 32'h42745dba};
test_input[1128:1135] = '{32'hc0aecbe9, 32'hc1e55d93, 32'h42028366, 32'h42336ae9, 32'hc1337cd5, 32'hc2323fb0, 32'h4259aa85, 32'h42b263fc};
test_output[1128:1135] = '{32'h0, 32'h0, 32'h42028366, 32'h42336ae9, 32'h0, 32'h0, 32'h4259aa85, 32'h42b263fc};
test_input[1136:1143] = '{32'hc1d0fce3, 32'hc02b2ac0, 32'h429c851c, 32'hc27ffae0, 32'h423bfa8a, 32'h426d384c, 32'h42ac5248, 32'hc1787728};
test_output[1136:1143] = '{32'h0, 32'h0, 32'h429c851c, 32'h0, 32'h423bfa8a, 32'h426d384c, 32'h42ac5248, 32'h0};
test_input[1144:1151] = '{32'hc2959af1, 32'hc25a7b92, 32'h42448dfa, 32'hc29e9827, 32'h4189e52d, 32'h42074751, 32'hc28ce805, 32'hc27dd216};
test_output[1144:1151] = '{32'h0, 32'h0, 32'h42448dfa, 32'h0, 32'h4189e52d, 32'h42074751, 32'h0, 32'h0};
test_input[1152:1159] = '{32'h42000bdf, 32'h427bd1f2, 32'h427945dd, 32'h42a5a45e, 32'h422155e0, 32'hc28e13f4, 32'hc1e55706, 32'hc2848728};
test_output[1152:1159] = '{32'h42000bdf, 32'h427bd1f2, 32'h427945dd, 32'h42a5a45e, 32'h422155e0, 32'h0, 32'h0, 32'h0};
test_input[1160:1167] = '{32'hc24cab42, 32'h422c3385, 32'h428f9ff0, 32'hc1c21bb9, 32'h4255defb, 32'h4202cbe5, 32'h42bd8ae6, 32'hbea4fb17};
test_output[1160:1167] = '{32'h0, 32'h422c3385, 32'h428f9ff0, 32'h0, 32'h4255defb, 32'h4202cbe5, 32'h42bd8ae6, 32'h0};
test_input[1168:1175] = '{32'hc2b7f846, 32'h40d7f3ec, 32'hc26e09dc, 32'h413e3f47, 32'h4236bacf, 32'hc1b400d5, 32'hc0958b06, 32'hc2b10980};
test_output[1168:1175] = '{32'h0, 32'h40d7f3ec, 32'h0, 32'h413e3f47, 32'h4236bacf, 32'h0, 32'h0, 32'h0};
test_input[1176:1183] = '{32'h42a23b5a, 32'hc1fdbf05, 32'h429421b9, 32'h4275f349, 32'h4197e295, 32'h42b0ecb8, 32'hc29fd1f9, 32'h415da9e7};
test_output[1176:1183] = '{32'h42a23b5a, 32'h0, 32'h429421b9, 32'h4275f349, 32'h4197e295, 32'h42b0ecb8, 32'h0, 32'h415da9e7};
test_input[1184:1191] = '{32'h425bbf69, 32'h42ac9d33, 32'hc2350e50, 32'h42312767, 32'hc1cdfa08, 32'h41959f70, 32'h429207e1, 32'hc2355198};
test_output[1184:1191] = '{32'h425bbf69, 32'h42ac9d33, 32'h0, 32'h42312767, 32'h0, 32'h41959f70, 32'h429207e1, 32'h0};
test_input[1192:1199] = '{32'h42862841, 32'hc1dcc27e, 32'hc2bbb57a, 32'h42a94eb0, 32'hc1d19b8b, 32'hc247a06a, 32'hc19cf394, 32'hc1a2326f};
test_output[1192:1199] = '{32'h42862841, 32'h0, 32'h0, 32'h42a94eb0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1200:1207] = '{32'hc1c4fae6, 32'h4242ee31, 32'h407c4e7c, 32'h42b48e50, 32'h422a7ca2, 32'hc0f626ad, 32'hc2bdf0de, 32'hc2848ff9};
test_output[1200:1207] = '{32'h0, 32'h4242ee31, 32'h407c4e7c, 32'h42b48e50, 32'h422a7ca2, 32'h0, 32'h0, 32'h0};
test_input[1208:1215] = '{32'hc2217de7, 32'hc2b8065d, 32'h4154560c, 32'h41d8bead, 32'hc1efafa9, 32'h42aebf01, 32'hc29ea254, 32'h42ab1b22};
test_output[1208:1215] = '{32'h0, 32'h0, 32'h4154560c, 32'h41d8bead, 32'h0, 32'h42aebf01, 32'h0, 32'h42ab1b22};
test_input[1216:1223] = '{32'h420cbd44, 32'hbfa43caa, 32'hc2a1552f, 32'hc1e2656f, 32'h42144835, 32'hc28b2b63, 32'hc26e61a7, 32'hc232ee42};
test_output[1216:1223] = '{32'h420cbd44, 32'h0, 32'h0, 32'h0, 32'h42144835, 32'h0, 32'h0, 32'h0};
test_input[1224:1231] = '{32'hc29b038d, 32'hc19452ff, 32'hc1a4336e, 32'hc253852e, 32'h427371f7, 32'hc2434a65, 32'hc1d51662, 32'h4187f81d};
test_output[1224:1231] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h427371f7, 32'h0, 32'h0, 32'h4187f81d};
test_input[1232:1239] = '{32'h41f71ac5, 32'hc2adc9d0, 32'hc2693773, 32'hc24f5243, 32'hc22b02e7, 32'hc0e3b0d1, 32'h426a47d3, 32'h42c71975};
test_output[1232:1239] = '{32'h41f71ac5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426a47d3, 32'h42c71975};
test_input[1240:1247] = '{32'h42110cfe, 32'h424c6869, 32'hc118e0c4, 32'hc1b93168, 32'h42c10f4e, 32'h42aa0993, 32'hc14f8652, 32'h41c89671};
test_output[1240:1247] = '{32'h42110cfe, 32'h424c6869, 32'h0, 32'h0, 32'h42c10f4e, 32'h42aa0993, 32'h0, 32'h41c89671};
test_input[1248:1255] = '{32'h3f160043, 32'h41852ce7, 32'h425ee9b7, 32'h421a3e19, 32'hc29f6b21, 32'h41cc4148, 32'hc0372ab7, 32'hc223a563};
test_output[1248:1255] = '{32'h3f160043, 32'h41852ce7, 32'h425ee9b7, 32'h421a3e19, 32'h0, 32'h41cc4148, 32'h0, 32'h0};
test_input[1256:1263] = '{32'h423b0d92, 32'hc12a4067, 32'hc1d39960, 32'h42c4c8f5, 32'h421e7651, 32'h421101e4, 32'h40e4930a, 32'h428b53b6};
test_output[1256:1263] = '{32'h423b0d92, 32'h0, 32'h0, 32'h42c4c8f5, 32'h421e7651, 32'h421101e4, 32'h40e4930a, 32'h428b53b6};
test_input[1264:1271] = '{32'hc2641001, 32'h4291dea2, 32'hbdcc8e87, 32'hc219fd85, 32'hc131092d, 32'hc2a69ac9, 32'hc29edbe2, 32'hc2b70fe1};
test_output[1264:1271] = '{32'h0, 32'h4291dea2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1272:1279] = '{32'h42865712, 32'h41b6d9ad, 32'h3f70ac13, 32'hc243d9a9, 32'h4281a762, 32'hc1e8ba3b, 32'h4259ea44, 32'h424e5406};
test_output[1272:1279] = '{32'h42865712, 32'h41b6d9ad, 32'h3f70ac13, 32'h0, 32'h4281a762, 32'h0, 32'h4259ea44, 32'h424e5406};
test_input[1280:1287] = '{32'h42b37541, 32'h42b3ed4b, 32'hc2a5f3c4, 32'h41bd4b35, 32'h42936012, 32'hc1496256, 32'h4295c665, 32'hc2530e6d};
test_output[1280:1287] = '{32'h42b37541, 32'h42b3ed4b, 32'h0, 32'h41bd4b35, 32'h42936012, 32'h0, 32'h4295c665, 32'h0};
test_input[1288:1295] = '{32'h423a59c9, 32'h424bf00c, 32'hc29dc783, 32'h4252b7d2, 32'hc28625be, 32'h42bb96a4, 32'hc230d468, 32'h4285b4fa};
test_output[1288:1295] = '{32'h423a59c9, 32'h424bf00c, 32'h0, 32'h4252b7d2, 32'h0, 32'h42bb96a4, 32'h0, 32'h4285b4fa};
test_input[1296:1303] = '{32'h4233dcd6, 32'hc1434419, 32'h425379ae, 32'h41e796fe, 32'hc06fad86, 32'h4218dc83, 32'h422058a8, 32'h42a8f7f4};
test_output[1296:1303] = '{32'h4233dcd6, 32'h0, 32'h425379ae, 32'h41e796fe, 32'h0, 32'h4218dc83, 32'h422058a8, 32'h42a8f7f4};
test_input[1304:1311] = '{32'h41a376f8, 32'h419af1bb, 32'hc282cbfc, 32'h41a90c60, 32'hc15e41ee, 32'hc11d16c2, 32'h42b5bba1, 32'h41ef2c52};
test_output[1304:1311] = '{32'h41a376f8, 32'h419af1bb, 32'h0, 32'h41a90c60, 32'h0, 32'h0, 32'h42b5bba1, 32'h41ef2c52};
test_input[1312:1319] = '{32'hc2173280, 32'h42090450, 32'hc19fbee0, 32'h428871cf, 32'h422d5d60, 32'h42b92e49, 32'h42349281, 32'h424ca049};
test_output[1312:1319] = '{32'h0, 32'h42090450, 32'h0, 32'h428871cf, 32'h422d5d60, 32'h42b92e49, 32'h42349281, 32'h424ca049};
test_input[1320:1327] = '{32'hc2834cca, 32'h401ef372, 32'hc25e9849, 32'h420a7195, 32'h4010bf4c, 32'h42a50766, 32'hc2c77e7e, 32'hc0e0c466};
test_output[1320:1327] = '{32'h0, 32'h401ef372, 32'h0, 32'h420a7195, 32'h4010bf4c, 32'h42a50766, 32'h0, 32'h0};
test_input[1328:1335] = '{32'h42b4aca9, 32'h42bb55f4, 32'hc28661bd, 32'hc21f82a5, 32'hc26f533e, 32'h42ba70b0, 32'h42a8d4e5, 32'hc23a3923};
test_output[1328:1335] = '{32'h42b4aca9, 32'h42bb55f4, 32'h0, 32'h0, 32'h0, 32'h42ba70b0, 32'h42a8d4e5, 32'h0};
test_input[1336:1343] = '{32'hc0a518a9, 32'h421f18d9, 32'hc1c38086, 32'h42215e5c, 32'hc245d5d8, 32'hc2720fd2, 32'hc2a742e1, 32'h411a6570};
test_output[1336:1343] = '{32'h0, 32'h421f18d9, 32'h0, 32'h42215e5c, 32'h0, 32'h0, 32'h0, 32'h411a6570};
test_input[1344:1351] = '{32'hc1c66279, 32'hc2933ea7, 32'hc1481981, 32'hc2294ba7, 32'h428ba7c0, 32'h40c74274, 32'hc1eaee21, 32'hc25f35eb};
test_output[1344:1351] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h428ba7c0, 32'h40c74274, 32'h0, 32'h0};
test_input[1352:1359] = '{32'h407da726, 32'hc1a204d4, 32'hc25e9878, 32'h40e87592, 32'hc1cbaf37, 32'hc2648aa4, 32'h42b5f360, 32'h424aba9f};
test_output[1352:1359] = '{32'h407da726, 32'h0, 32'h0, 32'h40e87592, 32'h0, 32'h0, 32'h42b5f360, 32'h424aba9f};
test_input[1360:1367] = '{32'h40cce56b, 32'hc2797767, 32'hc1da0f15, 32'hc2483a19, 32'hc248d481, 32'h4291c95a, 32'hc248837c, 32'h425663fa};
test_output[1360:1367] = '{32'h40cce56b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4291c95a, 32'h0, 32'h425663fa};
test_input[1368:1375] = '{32'h4290ad55, 32'hc2585312, 32'hc2c384df, 32'hc2c3e8a6, 32'h4251c331, 32'h429ce6cb, 32'hc1c4715f, 32'hc17a3289};
test_output[1368:1375] = '{32'h4290ad55, 32'h0, 32'h0, 32'h0, 32'h4251c331, 32'h429ce6cb, 32'h0, 32'h0};
test_input[1376:1383] = '{32'h420cb6c3, 32'h42bc5973, 32'h41f127e5, 32'h418588bd, 32'hc2080276, 32'hc1f256c8, 32'h3ff2ed8e, 32'h419c86d2};
test_output[1376:1383] = '{32'h420cb6c3, 32'h42bc5973, 32'h41f127e5, 32'h418588bd, 32'h0, 32'h0, 32'h3ff2ed8e, 32'h419c86d2};
test_input[1384:1391] = '{32'hc29ea078, 32'hc29cae1f, 32'hc27a1d16, 32'hc12c1a7a, 32'hc2011cf9, 32'hc26b1237, 32'hc2b9e8d9, 32'h4268db60};
test_output[1384:1391] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4268db60};
test_input[1392:1399] = '{32'h41d3809d, 32'hc293fc5e, 32'hc2a3c0aa, 32'hc27a8c0f, 32'hc2c6715b, 32'h42c56a95, 32'hc23dd5c5, 32'h420e44ed};
test_output[1392:1399] = '{32'h41d3809d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c56a95, 32'h0, 32'h420e44ed};
test_input[1400:1407] = '{32'h42057529, 32'hc24c3077, 32'hc24e7575, 32'h42c53730, 32'hc224ea05, 32'hc2009c1f, 32'hc2852858, 32'h426fd227};
test_output[1400:1407] = '{32'h42057529, 32'h0, 32'h0, 32'h42c53730, 32'h0, 32'h0, 32'h0, 32'h426fd227};
test_input[1408:1415] = '{32'hc29b569a, 32'h42552ab0, 32'hc2596280, 32'h416cfed2, 32'h42c5ff29, 32'hc23cedee, 32'hc296d712, 32'hc2a9d89e};
test_output[1408:1415] = '{32'h0, 32'h42552ab0, 32'h0, 32'h416cfed2, 32'h42c5ff29, 32'h0, 32'h0, 32'h0};
test_input[1416:1423] = '{32'hc2b5dff7, 32'h42c5063e, 32'hc2855f00, 32'hc24ae0ad, 32'hc2153f5c, 32'hc2c2e322, 32'h42447d82, 32'hc1efdd65};
test_output[1416:1423] = '{32'h0, 32'h42c5063e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42447d82, 32'h0};
test_input[1424:1431] = '{32'hc29fe5b2, 32'h41c393ab, 32'h41ec6242, 32'hc1348d44, 32'h4194a14e, 32'hc25e4853, 32'hc262a5a9, 32'h426ed35d};
test_output[1424:1431] = '{32'h0, 32'h41c393ab, 32'h41ec6242, 32'h0, 32'h4194a14e, 32'h0, 32'h0, 32'h426ed35d};
test_input[1432:1439] = '{32'hc2ad880e, 32'hc2c52308, 32'hc124455c, 32'hc29bd430, 32'hc222a643, 32'h422b939d, 32'h425b53a0, 32'h3f60b924};
test_output[1432:1439] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422b939d, 32'h425b53a0, 32'h3f60b924};
test_input[1440:1447] = '{32'hc182b30c, 32'h40cef2a0, 32'hc2adb210, 32'h420ffa33, 32'hc14c5709, 32'h406e2b2f, 32'hc242ac74, 32'hc26eb16b};
test_output[1440:1447] = '{32'h0, 32'h40cef2a0, 32'h0, 32'h420ffa33, 32'h0, 32'h406e2b2f, 32'h0, 32'h0};
test_input[1448:1455] = '{32'hc2aff8f7, 32'h423c1140, 32'hc2c1e5b6, 32'hc22230e6, 32'hc28b23b8, 32'h42b7076e, 32'h423d6f00, 32'h42231d99};
test_output[1448:1455] = '{32'h0, 32'h423c1140, 32'h0, 32'h0, 32'h0, 32'h42b7076e, 32'h423d6f00, 32'h42231d99};
test_input[1456:1463] = '{32'h429caa96, 32'h428fa536, 32'hc2855c8a, 32'h429dc95d, 32'h42817593, 32'hc1a419bd, 32'hc04d6cd5, 32'h42a2a8e9};
test_output[1456:1463] = '{32'h429caa96, 32'h428fa536, 32'h0, 32'h429dc95d, 32'h42817593, 32'h0, 32'h0, 32'h42a2a8e9};
test_input[1464:1471] = '{32'hc26ddcff, 32'h428a4e89, 32'hc28a2025, 32'hc203bdb6, 32'h41837064, 32'h42c3e0e1, 32'h3fed610d, 32'hc2a74e69};
test_output[1464:1471] = '{32'h0, 32'h428a4e89, 32'h0, 32'h0, 32'h41837064, 32'h42c3e0e1, 32'h3fed610d, 32'h0};
test_input[1472:1479] = '{32'h42110381, 32'hc16b8321, 32'h42285430, 32'hc2b062a5, 32'h42b5a921, 32'hc1056647, 32'hc2ae0fe7, 32'h420ce00e};
test_output[1472:1479] = '{32'h42110381, 32'h0, 32'h42285430, 32'h0, 32'h42b5a921, 32'h0, 32'h0, 32'h420ce00e};
test_input[1480:1487] = '{32'h4268818a, 32'hc27c7051, 32'hc226d71c, 32'h4290f121, 32'h429f7765, 32'hc2c73994, 32'h42b02840, 32'h425361d6};
test_output[1480:1487] = '{32'h4268818a, 32'h0, 32'h0, 32'h4290f121, 32'h429f7765, 32'h0, 32'h42b02840, 32'h425361d6};
test_input[1488:1495] = '{32'h42784b6c, 32'h423d7d2e, 32'hc223451a, 32'hc12f9556, 32'h40cf9f33, 32'h42921037, 32'h41880c7f, 32'h42b79776};
test_output[1488:1495] = '{32'h42784b6c, 32'h423d7d2e, 32'h0, 32'h0, 32'h40cf9f33, 32'h42921037, 32'h41880c7f, 32'h42b79776};
test_input[1496:1503] = '{32'h420d79d9, 32'h4218e02a, 32'h41c20efd, 32'hc28f6a5c, 32'h4248f688, 32'hc2b58581, 32'hbf9337c0, 32'h41829d70};
test_output[1496:1503] = '{32'h420d79d9, 32'h4218e02a, 32'h41c20efd, 32'h0, 32'h4248f688, 32'h0, 32'h0, 32'h41829d70};
test_input[1504:1511] = '{32'h4289c2a6, 32'hc2a674dd, 32'hc26ef840, 32'hc1ac983a, 32'hc23998d9, 32'h42519c1e, 32'h428c0bd2, 32'h4203d8f3};
test_output[1504:1511] = '{32'h4289c2a6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42519c1e, 32'h428c0bd2, 32'h4203d8f3};
test_input[1512:1519] = '{32'hc247bb2a, 32'hc2c77ea5, 32'hc25e2bbb, 32'hc236e2c8, 32'h42836126, 32'hc1cee5e0, 32'hc19811b9, 32'h420c219c};
test_output[1512:1519] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42836126, 32'h0, 32'h0, 32'h420c219c};
test_input[1520:1527] = '{32'h420f9ce3, 32'h42a8c031, 32'h4266d655, 32'h41e36851, 32'hc2105288, 32'hc0848ae6, 32'h42c03569, 32'hc12e4942};
test_output[1520:1527] = '{32'h420f9ce3, 32'h42a8c031, 32'h4266d655, 32'h41e36851, 32'h0, 32'h0, 32'h42c03569, 32'h0};
test_input[1528:1535] = '{32'h427e37cd, 32'hc21d7115, 32'h4287ac4a, 32'hc25cbf99, 32'hc24b2d08, 32'h422442d1, 32'h42147f9e, 32'hc29e1278};
test_output[1528:1535] = '{32'h427e37cd, 32'h0, 32'h4287ac4a, 32'h0, 32'h0, 32'h422442d1, 32'h42147f9e, 32'h0};
test_input[1536:1543] = '{32'h42bf83a8, 32'hc2636e2f, 32'h42217d24, 32'hc21e75d0, 32'h416f248d, 32'hc249c14a, 32'h42145103, 32'hc2796776};
test_output[1536:1543] = '{32'h42bf83a8, 32'h0, 32'h42217d24, 32'h0, 32'h416f248d, 32'h0, 32'h42145103, 32'h0};
test_input[1544:1551] = '{32'hc204b48c, 32'hc2416480, 32'h402601ac, 32'h42a4a97c, 32'hc1b9dce1, 32'hc29c0c1e, 32'hc1f0bccc, 32'hc2be1114};
test_output[1544:1551] = '{32'h0, 32'h0, 32'h402601ac, 32'h42a4a97c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1552:1559] = '{32'h41f8d66d, 32'h4206c6d7, 32'hc2c4195a, 32'hc28ed800, 32'hc21e6cb3, 32'h423edc45, 32'h42bf1b5b, 32'h42147a3e};
test_output[1552:1559] = '{32'h41f8d66d, 32'h4206c6d7, 32'h0, 32'h0, 32'h0, 32'h423edc45, 32'h42bf1b5b, 32'h42147a3e};
test_input[1560:1567] = '{32'h42c1e2ad, 32'hc23f98b6, 32'h420f2d46, 32'hc1e0c13e, 32'h4244ea76, 32'h423bc68e, 32'hc24de981, 32'hc1e66ba5};
test_output[1560:1567] = '{32'h42c1e2ad, 32'h0, 32'h420f2d46, 32'h0, 32'h4244ea76, 32'h423bc68e, 32'h0, 32'h0};
test_input[1568:1575] = '{32'h414c0086, 32'hc22cb992, 32'h42beb571, 32'hc197763d, 32'hc232cb91, 32'hc2c2ff20, 32'h4254180e, 32'h42a4aaf4};
test_output[1568:1575] = '{32'h414c0086, 32'h0, 32'h42beb571, 32'h0, 32'h0, 32'h0, 32'h4254180e, 32'h42a4aaf4};
test_input[1576:1583] = '{32'hc2c69127, 32'hc2a5a6a3, 32'hc2515a49, 32'h41f37cf1, 32'h3fb40b5e, 32'h4230342b, 32'h42bbdfe0, 32'hc293735f};
test_output[1576:1583] = '{32'h0, 32'h0, 32'h0, 32'h41f37cf1, 32'h3fb40b5e, 32'h4230342b, 32'h42bbdfe0, 32'h0};
test_input[1584:1591] = '{32'hc00382a1, 32'h41056a0f, 32'hc1cf20bc, 32'h42c7d341, 32'hc2c118e9, 32'hc2281c36, 32'h42a0ecb5, 32'hc28ac29a};
test_output[1584:1591] = '{32'h0, 32'h41056a0f, 32'h0, 32'h42c7d341, 32'h0, 32'h0, 32'h42a0ecb5, 32'h0};
test_input[1592:1599] = '{32'hc26591f3, 32'hc1c63321, 32'hc284aa93, 32'h42c70fe5, 32'h414b567f, 32'hc24cbe9e, 32'h42b8cd42, 32'h41b1e5a1};
test_output[1592:1599] = '{32'h0, 32'h0, 32'h0, 32'h42c70fe5, 32'h414b567f, 32'h0, 32'h42b8cd42, 32'h41b1e5a1};
test_input[1600:1607] = '{32'hc2604fac, 32'h42aae8e7, 32'h427723a1, 32'hc2487d61, 32'hc1c2a0f4, 32'h423b4e89, 32'hc0460950, 32'h425745c8};
test_output[1600:1607] = '{32'h0, 32'h42aae8e7, 32'h427723a1, 32'h0, 32'h0, 32'h423b4e89, 32'h0, 32'h425745c8};
test_input[1608:1615] = '{32'h41b4ce09, 32'h41b530d1, 32'h4209e66c, 32'hc2b29a42, 32'h42b08cc3, 32'hc21ea319, 32'hc20d2108, 32'h4043db75};
test_output[1608:1615] = '{32'h41b4ce09, 32'h41b530d1, 32'h4209e66c, 32'h0, 32'h42b08cc3, 32'h0, 32'h0, 32'h4043db75};
test_input[1616:1623] = '{32'h42ba661e, 32'hc21ed7f6, 32'h4272434b, 32'h4276bad1, 32'h411f2c87, 32'h40f65bb8, 32'hc1acaa6c, 32'hc293641e};
test_output[1616:1623] = '{32'h42ba661e, 32'h0, 32'h4272434b, 32'h4276bad1, 32'h411f2c87, 32'h40f65bb8, 32'h0, 32'h0};
test_input[1624:1631] = '{32'h42b67167, 32'h42851e06, 32'hc2b4143f, 32'h42631a68, 32'h426d5c79, 32'hc28cf574, 32'h4091c912, 32'hc2808105};
test_output[1624:1631] = '{32'h42b67167, 32'h42851e06, 32'h0, 32'h42631a68, 32'h426d5c79, 32'h0, 32'h4091c912, 32'h0};
test_input[1632:1639] = '{32'hc2459c73, 32'hc2151f8f, 32'hc29429fe, 32'h42c02cc3, 32'h41a6aeb4, 32'hc101f73a, 32'h42ab2144, 32'h417565d6};
test_output[1632:1639] = '{32'h0, 32'h0, 32'h0, 32'h42c02cc3, 32'h41a6aeb4, 32'h0, 32'h42ab2144, 32'h417565d6};
test_input[1640:1647] = '{32'h4182a07f, 32'h3fb3126a, 32'hc1cbea3c, 32'h42b74726, 32'h42132f3b, 32'hc21496f7, 32'hc1dd2a70, 32'h423f9b65};
test_output[1640:1647] = '{32'h4182a07f, 32'h3fb3126a, 32'h0, 32'h42b74726, 32'h42132f3b, 32'h0, 32'h0, 32'h423f9b65};
test_input[1648:1655] = '{32'hc2594c4d, 32'h4278fbdf, 32'h41cb293b, 32'h42a0d3de, 32'h4297cbc6, 32'h42869284, 32'hc283b2e8, 32'hc28aecb3};
test_output[1648:1655] = '{32'h0, 32'h4278fbdf, 32'h41cb293b, 32'h42a0d3de, 32'h4297cbc6, 32'h42869284, 32'h0, 32'h0};
test_input[1656:1663] = '{32'h42bc1215, 32'hc2a75210, 32'h41808ad8, 32'hc29fd035, 32'hbf7c7121, 32'h41b1a46b, 32'hc2ae6cf2, 32'h4239a5f0};
test_output[1656:1663] = '{32'h42bc1215, 32'h0, 32'h41808ad8, 32'h0, 32'h0, 32'h41b1a46b, 32'h0, 32'h4239a5f0};
test_input[1664:1671] = '{32'h421fb137, 32'hc1a44298, 32'h41b1b9a5, 32'h4258cbc4, 32'h403cbd06, 32'h41ce10e4, 32'h429a32a9, 32'h414201b4};
test_output[1664:1671] = '{32'h421fb137, 32'h0, 32'h41b1b9a5, 32'h4258cbc4, 32'h403cbd06, 32'h41ce10e4, 32'h429a32a9, 32'h414201b4};
test_input[1672:1679] = '{32'h42829af9, 32'h41056273, 32'hc188a2b0, 32'h4272feb0, 32'hc236bbe2, 32'h42b0b2f6, 32'hc2109696, 32'h41a4d4e2};
test_output[1672:1679] = '{32'h42829af9, 32'h41056273, 32'h0, 32'h4272feb0, 32'h0, 32'h42b0b2f6, 32'h0, 32'h41a4d4e2};
test_input[1680:1687] = '{32'h4254953e, 32'hc265e269, 32'hc19543ed, 32'hc25c3978, 32'h422d0977, 32'hc10b463b, 32'h420b90ed, 32'h40492e76};
test_output[1680:1687] = '{32'h4254953e, 32'h0, 32'h0, 32'h0, 32'h422d0977, 32'h0, 32'h420b90ed, 32'h40492e76};
test_input[1688:1695] = '{32'h41ef33b8, 32'hc2b1de94, 32'h427b6652, 32'h4228edc0, 32'hc2ba45aa, 32'hc15605fc, 32'hc2af2d0b, 32'hc1efae5f};
test_output[1688:1695] = '{32'h41ef33b8, 32'h0, 32'h427b6652, 32'h4228edc0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[1696:1703] = '{32'hc0d9e6f6, 32'h427698e2, 32'h417a3766, 32'hc10a7d16, 32'hc265d8e4, 32'h418c0adb, 32'hc20454f2, 32'hc2ab120b};
test_output[1696:1703] = '{32'h0, 32'h427698e2, 32'h417a3766, 32'h0, 32'h0, 32'h418c0adb, 32'h0, 32'h0};
test_input[1704:1711] = '{32'h428ef448, 32'h42c28d25, 32'h426a54fb, 32'hc11f288e, 32'h42c292d0, 32'h42c0f6c9, 32'hc10bc873, 32'h4298d5ee};
test_output[1704:1711] = '{32'h428ef448, 32'h42c28d25, 32'h426a54fb, 32'h0, 32'h42c292d0, 32'h42c0f6c9, 32'h0, 32'h4298d5ee};
test_input[1712:1719] = '{32'h407e1cf0, 32'h41842dcc, 32'h41c2d0e4, 32'h41ea428b, 32'h42557499, 32'hc27956af, 32'hc19b3602, 32'hc100b9ef};
test_output[1712:1719] = '{32'h407e1cf0, 32'h41842dcc, 32'h41c2d0e4, 32'h41ea428b, 32'h42557499, 32'h0, 32'h0, 32'h0};
test_input[1720:1727] = '{32'hc1ea4b23, 32'hc29f3360, 32'hc2b26d54, 32'hc27348ac, 32'h40a4699f, 32'h4284ee95, 32'hc244142a, 32'hc23b5c7d};
test_output[1720:1727] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40a4699f, 32'h4284ee95, 32'h0, 32'h0};
test_input[1728:1735] = '{32'hc1869601, 32'hc24b76a8, 32'h4295b68f, 32'h415642f7, 32'h429f03da, 32'hc22a8e86, 32'hc26a672e, 32'hc2bd2bb1};
test_output[1728:1735] = '{32'h0, 32'h0, 32'h4295b68f, 32'h415642f7, 32'h429f03da, 32'h0, 32'h0, 32'h0};
test_input[1736:1743] = '{32'hc2ae1dce, 32'hc18b1965, 32'h40f9850d, 32'hc2ae4741, 32'hc245d00d, 32'hc1a9720b, 32'hc24eb60a, 32'h42577694};
test_output[1736:1743] = '{32'h0, 32'h0, 32'h40f9850d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42577694};
test_input[1744:1751] = '{32'h4262fa2b, 32'h426a9884, 32'hc155a282, 32'hc26ec6fd, 32'h42689c51, 32'h414b7eba, 32'h41c701cd, 32'h42c754ca};
test_output[1744:1751] = '{32'h4262fa2b, 32'h426a9884, 32'h0, 32'h0, 32'h42689c51, 32'h414b7eba, 32'h41c701cd, 32'h42c754ca};
test_input[1752:1759] = '{32'h41225690, 32'h4257c0da, 32'hc2968886, 32'h3edf38f0, 32'h4185e34f, 32'hc28496d7, 32'hc006ae31, 32'h40d4168a};
test_output[1752:1759] = '{32'h41225690, 32'h4257c0da, 32'h0, 32'h3edf38f0, 32'h4185e34f, 32'h0, 32'h0, 32'h40d4168a};
test_input[1760:1767] = '{32'hc0185ed7, 32'h422280a8, 32'h423bea6f, 32'h42bf4727, 32'h42a5b406, 32'hc00f5678, 32'hc14cd685, 32'hc29576f2};
test_output[1760:1767] = '{32'h0, 32'h422280a8, 32'h423bea6f, 32'h42bf4727, 32'h42a5b406, 32'h0, 32'h0, 32'h0};
test_input[1768:1775] = '{32'h42a3df63, 32'hc1b62895, 32'h42a4b94f, 32'hc219a55a, 32'hc27fa611, 32'h4299eb46, 32'h42b28630, 32'h42a9ed3b};
test_output[1768:1775] = '{32'h42a3df63, 32'h0, 32'h42a4b94f, 32'h0, 32'h0, 32'h4299eb46, 32'h42b28630, 32'h42a9ed3b};
test_input[1776:1783] = '{32'hc1e63ead, 32'h42b8c810, 32'h413cca20, 32'h425745ac, 32'hc216d8c7, 32'h4207fb1b, 32'hc28e8964, 32'hc1c59446};
test_output[1776:1783] = '{32'h0, 32'h42b8c810, 32'h413cca20, 32'h425745ac, 32'h0, 32'h4207fb1b, 32'h0, 32'h0};
test_input[1784:1791] = '{32'hc2925caf, 32'h41496a39, 32'hc1b1dbc5, 32'h41729fe1, 32'h410e2868, 32'hc2baa8b0, 32'hc26bd208, 32'hc2ad4d5c};
test_output[1784:1791] = '{32'h0, 32'h41496a39, 32'h0, 32'h41729fe1, 32'h410e2868, 32'h0, 32'h0, 32'h0};
test_input[1792:1799] = '{32'hc29ce0f2, 32'h427b12c4, 32'hc272c40a, 32'hc1aad8ff, 32'hc267c688, 32'hc2c783dd, 32'h423a3d50, 32'hc2bcb2f1};
test_output[1792:1799] = '{32'h0, 32'h427b12c4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423a3d50, 32'h0};
test_input[1800:1807] = '{32'hc29f2d41, 32'h411376a9, 32'h4208da15, 32'h41f278cb, 32'h3ff11298, 32'hc28ddfdd, 32'h41a5cb1d, 32'hc23e0c6b};
test_output[1800:1807] = '{32'h0, 32'h411376a9, 32'h4208da15, 32'h41f278cb, 32'h3ff11298, 32'h0, 32'h41a5cb1d, 32'h0};
test_input[1808:1815] = '{32'h42a72b70, 32'hc255c317, 32'h42b691fb, 32'h42b60eb8, 32'hc273de32, 32'h421a0b2e, 32'hc2b9217f, 32'hc18f22f2};
test_output[1808:1815] = '{32'h42a72b70, 32'h0, 32'h42b691fb, 32'h42b60eb8, 32'h0, 32'h421a0b2e, 32'h0, 32'h0};
test_input[1816:1823] = '{32'h42892d84, 32'hc234a25a, 32'hc2c05c65, 32'h425d1fbb, 32'hc218e076, 32'hc2baae08, 32'h421405d3, 32'hc2b8e334};
test_output[1816:1823] = '{32'h42892d84, 32'h0, 32'h0, 32'h425d1fbb, 32'h0, 32'h0, 32'h421405d3, 32'h0};
test_input[1824:1831] = '{32'hc236d1d3, 32'hc22fa531, 32'hc1cbac3a, 32'h428aed54, 32'h42a82507, 32'hc2ba63f6, 32'h42ba1a8b, 32'h4170174e};
test_output[1824:1831] = '{32'h0, 32'h0, 32'h0, 32'h428aed54, 32'h42a82507, 32'h0, 32'h42ba1a8b, 32'h4170174e};
test_input[1832:1839] = '{32'h42633952, 32'h41d15a11, 32'h41a5a7ff, 32'hc1be21c5, 32'hc2a6cc66, 32'hc226a51b, 32'hc19f8849, 32'h4296a3a4};
test_output[1832:1839] = '{32'h42633952, 32'h41d15a11, 32'h41a5a7ff, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4296a3a4};
test_input[1840:1847] = '{32'h422c43ff, 32'h42c1d200, 32'h421f206b, 32'hc2068ff6, 32'hc22cd125, 32'h41392bd1, 32'hc22497c6, 32'h41db1ae6};
test_output[1840:1847] = '{32'h422c43ff, 32'h42c1d200, 32'h421f206b, 32'h0, 32'h0, 32'h41392bd1, 32'h0, 32'h41db1ae6};
test_input[1848:1855] = '{32'h42acb7a2, 32'h42882644, 32'hc2475f1e, 32'h41d3d1ce, 32'hc2836669, 32'h42be8a4f, 32'hc1e4ca7f, 32'h428cac66};
test_output[1848:1855] = '{32'h42acb7a2, 32'h42882644, 32'h0, 32'h41d3d1ce, 32'h0, 32'h42be8a4f, 32'h0, 32'h428cac66};
test_input[1856:1863] = '{32'hc29669ec, 32'hc2a340e6, 32'hc2ac31a9, 32'h414bb1b3, 32'h41c7971b, 32'hc213ddb6, 32'h417031d9, 32'hc25c5146};
test_output[1856:1863] = '{32'h0, 32'h0, 32'h0, 32'h414bb1b3, 32'h41c7971b, 32'h0, 32'h417031d9, 32'h0};
test_input[1864:1871] = '{32'hc2c3b6fd, 32'hc13693f3, 32'h3f44640b, 32'hc292bbda, 32'h42b181fc, 32'hc2656d55, 32'hc07e34ef, 32'h42a9b820};
test_output[1864:1871] = '{32'h0, 32'h0, 32'h3f44640b, 32'h0, 32'h42b181fc, 32'h0, 32'h0, 32'h42a9b820};
test_input[1872:1879] = '{32'h42737ba3, 32'h4185e8a6, 32'hc29c5c40, 32'h409409cb, 32'hc1e6cada, 32'h409e1efc, 32'hc115e0bd, 32'h4081be5b};
test_output[1872:1879] = '{32'h42737ba3, 32'h4185e8a6, 32'h0, 32'h409409cb, 32'h0, 32'h409e1efc, 32'h0, 32'h4081be5b};
test_input[1880:1887] = '{32'h41c453b2, 32'hc15161fd, 32'h41c904e3, 32'hc20803f7, 32'hc2c518c7, 32'h429101c7, 32'h41660b12, 32'h4150a419};
test_output[1880:1887] = '{32'h41c453b2, 32'h0, 32'h41c904e3, 32'h0, 32'h0, 32'h429101c7, 32'h41660b12, 32'h4150a419};
test_input[1888:1895] = '{32'hc298eb34, 32'h42c4a294, 32'hc18e9dd9, 32'h42a886e4, 32'h42b601dc, 32'h42862163, 32'hc2638227, 32'hc2078166};
test_output[1888:1895] = '{32'h0, 32'h42c4a294, 32'h0, 32'h42a886e4, 32'h42b601dc, 32'h42862163, 32'h0, 32'h0};
test_input[1896:1903] = '{32'h426829f3, 32'hc1890b17, 32'h4171d4b9, 32'h42689b4f, 32'h41853696, 32'h42c61549, 32'h421aa420, 32'hc2328779};
test_output[1896:1903] = '{32'h426829f3, 32'h0, 32'h4171d4b9, 32'h42689b4f, 32'h41853696, 32'h42c61549, 32'h421aa420, 32'h0};
test_input[1904:1911] = '{32'hc1e8d565, 32'h4293b6d0, 32'hc2be018e, 32'hc1a953e6, 32'h418b96f0, 32'hc1ce85ec, 32'hc2bcd656, 32'hc2a2fd17};
test_output[1904:1911] = '{32'h0, 32'h4293b6d0, 32'h0, 32'h0, 32'h418b96f0, 32'h0, 32'h0, 32'h0};
test_input[1912:1919] = '{32'hc26da6fd, 32'h42723d71, 32'h420bb755, 32'hc2b9b5b5, 32'h418e6e6e, 32'hc21af964, 32'hc2beefbc, 32'hc251dc82};
test_output[1912:1919] = '{32'h0, 32'h42723d71, 32'h420bb755, 32'h0, 32'h418e6e6e, 32'h0, 32'h0, 32'h0};
test_input[1920:1927] = '{32'h4287a45f, 32'hc2149e24, 32'h42563a2d, 32'hc0b6e803, 32'h42a6e5c2, 32'h42a898a8, 32'hc1adc305, 32'hc143c642};
test_output[1920:1927] = '{32'h4287a45f, 32'h0, 32'h42563a2d, 32'h0, 32'h42a6e5c2, 32'h42a898a8, 32'h0, 32'h0};
test_input[1928:1935] = '{32'h3fcbf284, 32'h429b4565, 32'h41f02a98, 32'h41ebee80, 32'hc2a2d063, 32'hc298800d, 32'h42534a5c, 32'h424a9541};
test_output[1928:1935] = '{32'h3fcbf284, 32'h429b4565, 32'h41f02a98, 32'h41ebee80, 32'h0, 32'h0, 32'h42534a5c, 32'h424a9541};
test_input[1936:1943] = '{32'h426ed222, 32'hc16e0302, 32'h42455f65, 32'hc25a7914, 32'h42c13440, 32'hc2c2e0ed, 32'hc284ec59, 32'h429c904b};
test_output[1936:1943] = '{32'h426ed222, 32'h0, 32'h42455f65, 32'h0, 32'h42c13440, 32'h0, 32'h0, 32'h429c904b};
test_input[1944:1951] = '{32'h4261c953, 32'hc2bf42c3, 32'h41b032de, 32'h42981e89, 32'h42b6ea21, 32'hc247578b, 32'h420109a2, 32'h421a6018};
test_output[1944:1951] = '{32'h4261c953, 32'h0, 32'h41b032de, 32'h42981e89, 32'h42b6ea21, 32'h0, 32'h420109a2, 32'h421a6018};
test_input[1952:1959] = '{32'h40bc3e1c, 32'h42068482, 32'hc15ced72, 32'hc2891235, 32'h4151dc81, 32'h42b94711, 32'hc1bfcd2f, 32'h427e48ec};
test_output[1952:1959] = '{32'h40bc3e1c, 32'h42068482, 32'h0, 32'h0, 32'h4151dc81, 32'h42b94711, 32'h0, 32'h427e48ec};
test_input[1960:1967] = '{32'hc23a4bc5, 32'hc16fac98, 32'h41bf779b, 32'h41a5e2cd, 32'hc2c4b5fc, 32'h423afdf1, 32'hc1c29ffe, 32'hc27975bc};
test_output[1960:1967] = '{32'h0, 32'h0, 32'h41bf779b, 32'h41a5e2cd, 32'h0, 32'h423afdf1, 32'h0, 32'h0};
test_input[1968:1975] = '{32'hc17f836a, 32'hc2b8f0c9, 32'h4215cdf6, 32'hc1a4e106, 32'hc2332e82, 32'h42918eb3, 32'hc29d1179, 32'h42a672ab};
test_output[1968:1975] = '{32'h0, 32'h0, 32'h4215cdf6, 32'h0, 32'h0, 32'h42918eb3, 32'h0, 32'h42a672ab};
test_input[1976:1983] = '{32'hc0df540c, 32'h428b8c07, 32'hc28223f3, 32'hc265f46c, 32'h400fa202, 32'h4256e505, 32'hc1289ffa, 32'hc25d8ba5};
test_output[1976:1983] = '{32'h0, 32'h428b8c07, 32'h0, 32'h0, 32'h400fa202, 32'h4256e505, 32'h0, 32'h0};
test_input[1984:1991] = '{32'hc2aca166, 32'h4218bb72, 32'hc218ee60, 32'hc15f2f0e, 32'hc218056d, 32'h416f6081, 32'h420150d7, 32'h419978d5};
test_output[1984:1991] = '{32'h0, 32'h4218bb72, 32'h0, 32'h0, 32'h0, 32'h416f6081, 32'h420150d7, 32'h419978d5};
test_input[1992:1999] = '{32'hc28db701, 32'h429616a9, 32'hc233b43c, 32'h429e836d, 32'hc25055db, 32'hc253e07c, 32'hc253ed82, 32'hc2c2bc2c};
test_output[1992:1999] = '{32'h0, 32'h429616a9, 32'h0, 32'h429e836d, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2000:2007] = '{32'h429a970f, 32'hc1d06f6b, 32'hc2858a3b, 32'h42b4fed1, 32'hc2314e9e, 32'h4205eef3, 32'h42b61d45, 32'hc0879070};
test_output[2000:2007] = '{32'h429a970f, 32'h0, 32'h0, 32'h42b4fed1, 32'h0, 32'h4205eef3, 32'h42b61d45, 32'h0};
test_input[2008:2015] = '{32'h40583e08, 32'hc21d65c2, 32'h422ca14d, 32'h422b70e4, 32'h419261b7, 32'h422b3bcb, 32'h4144ceb4, 32'hc201630e};
test_output[2008:2015] = '{32'h40583e08, 32'h0, 32'h422ca14d, 32'h422b70e4, 32'h419261b7, 32'h422b3bcb, 32'h4144ceb4, 32'h0};
test_input[2016:2023] = '{32'hc23e30ec, 32'h42701d07, 32'hc2a21c30, 32'h424d32c7, 32'hc28bc11f, 32'hc249874e, 32'h428ca908, 32'h42b4790b};
test_output[2016:2023] = '{32'h0, 32'h42701d07, 32'h0, 32'h424d32c7, 32'h0, 32'h0, 32'h428ca908, 32'h42b4790b};
test_input[2024:2031] = '{32'hc183c108, 32'hc2c529f5, 32'hc0931944, 32'hc23942d4, 32'h42474a4b, 32'h42b290c8, 32'hc2a0046f, 32'hc2346b4f};
test_output[2024:2031] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42474a4b, 32'h42b290c8, 32'h0, 32'h0};
test_input[2032:2039] = '{32'hc23937bd, 32'h42af013a, 32'hc28dc7ee, 32'h419a2e33, 32'h42181e70, 32'h40d20939, 32'hc2a9b0a6, 32'hc2965a56};
test_output[2032:2039] = '{32'h0, 32'h42af013a, 32'h0, 32'h419a2e33, 32'h42181e70, 32'h40d20939, 32'h0, 32'h0};
test_input[2040:2047] = '{32'h42bb0509, 32'h42abcd67, 32'hc2498c4a, 32'hc247ceca, 32'h42978ae8, 32'hc2a48cd2, 32'h410ab0e2, 32'h429f08ba};
test_output[2040:2047] = '{32'h42bb0509, 32'h42abcd67, 32'h0, 32'h0, 32'h42978ae8, 32'h0, 32'h410ab0e2, 32'h429f08ba};
test_input[2048:2055] = '{32'h42a44f24, 32'h4217e210, 32'h41ec2b33, 32'hc288dac2, 32'hc24696f4, 32'h42b0c493, 32'h4108b6ef, 32'hc20ff51d};
test_output[2048:2055] = '{32'h42a44f24, 32'h4217e210, 32'h41ec2b33, 32'h0, 32'h0, 32'h42b0c493, 32'h4108b6ef, 32'h0};
test_input[2056:2063] = '{32'hc15ae7f0, 32'h42a0fab8, 32'hc2881262, 32'hc0f57c7e, 32'h41b91322, 32'hc27f656b, 32'h41efbfd4, 32'hc2c7c628};
test_output[2056:2063] = '{32'h0, 32'h42a0fab8, 32'h0, 32'h0, 32'h41b91322, 32'h0, 32'h41efbfd4, 32'h0};
test_input[2064:2071] = '{32'hc21543dd, 32'h42aa2ece, 32'hc28ac1f4, 32'h41bb21d8, 32'hc2b6bd04, 32'h42a3fdd7, 32'h4291ffef, 32'hc21f8a76};
test_output[2064:2071] = '{32'h0, 32'h42aa2ece, 32'h0, 32'h41bb21d8, 32'h0, 32'h42a3fdd7, 32'h4291ffef, 32'h0};
test_input[2072:2079] = '{32'hc2bd7546, 32'hc18c3a75, 32'hc28cf028, 32'h42a69821, 32'hc1ee4197, 32'hc271c93e, 32'hc20a0312, 32'hc1968d5c};
test_output[2072:2079] = '{32'h0, 32'h0, 32'h0, 32'h42a69821, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2080:2087] = '{32'h3e9cea82, 32'h42714995, 32'h425de75f, 32'h41ed976c, 32'hc29fb389, 32'h4210adce, 32'h42c55257, 32'hc29561c8};
test_output[2080:2087] = '{32'h3e9cea82, 32'h42714995, 32'h425de75f, 32'h41ed976c, 32'h0, 32'h4210adce, 32'h42c55257, 32'h0};
test_input[2088:2095] = '{32'h42bd0503, 32'h408e0bba, 32'hc147670f, 32'h4197275a, 32'hc0ced294, 32'h41a78f62, 32'h429b94c5, 32'hc204ad65};
test_output[2088:2095] = '{32'h42bd0503, 32'h408e0bba, 32'h0, 32'h4197275a, 32'h0, 32'h41a78f62, 32'h429b94c5, 32'h0};
test_input[2096:2103] = '{32'h4214c166, 32'hc1745c24, 32'h41abceeb, 32'h422c5a03, 32'h419bd915, 32'hc28fa4f8, 32'h412ac054, 32'h42a784a4};
test_output[2096:2103] = '{32'h4214c166, 32'h0, 32'h41abceeb, 32'h422c5a03, 32'h419bd915, 32'h0, 32'h412ac054, 32'h42a784a4};
test_input[2104:2111] = '{32'h41474131, 32'hc29d4214, 32'h3f3d74ea, 32'hc2bd630a, 32'hc2bacc0e, 32'hc24eef56, 32'h427248e2, 32'h4046368f};
test_output[2104:2111] = '{32'h41474131, 32'h0, 32'h3f3d74ea, 32'h0, 32'h0, 32'h0, 32'h427248e2, 32'h4046368f};
test_input[2112:2119] = '{32'h428eb493, 32'hc290e08d, 32'h4268ad49, 32'hc276a91b, 32'hc283b652, 32'h41ac0cdf, 32'h4299165d, 32'h40f3236e};
test_output[2112:2119] = '{32'h428eb493, 32'h0, 32'h4268ad49, 32'h0, 32'h0, 32'h41ac0cdf, 32'h4299165d, 32'h40f3236e};
test_input[2120:2127] = '{32'hc19d072c, 32'hc2884783, 32'h4206767f, 32'hc294e8a8, 32'hc27d2452, 32'hc283a446, 32'hc23e4ef8, 32'h41152c0a};
test_output[2120:2127] = '{32'h0, 32'h0, 32'h4206767f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41152c0a};
test_input[2128:2135] = '{32'hc0c6d6cd, 32'h42b25f55, 32'hc270d271, 32'h424bf73d, 32'h4282a8c4, 32'hc099bc96, 32'hc1687294, 32'h42bb1883};
test_output[2128:2135] = '{32'h0, 32'h42b25f55, 32'h0, 32'h424bf73d, 32'h4282a8c4, 32'h0, 32'h0, 32'h42bb1883};
test_input[2136:2143] = '{32'hc2bc0027, 32'hc295a788, 32'h42921193, 32'h41e30ab7, 32'h42a15277, 32'h4107f35f, 32'hc1d4d815, 32'hc273790b};
test_output[2136:2143] = '{32'h0, 32'h0, 32'h42921193, 32'h41e30ab7, 32'h42a15277, 32'h4107f35f, 32'h0, 32'h0};
test_input[2144:2151] = '{32'h4219460c, 32'hc27736fd, 32'hc2a12186, 32'hc2c3af57, 32'h41981412, 32'hc25a9e47, 32'hc26c9d0b, 32'hc2285f58};
test_output[2144:2151] = '{32'h4219460c, 32'h0, 32'h0, 32'h0, 32'h41981412, 32'h0, 32'h0, 32'h0};
test_input[2152:2159] = '{32'h42a0bb47, 32'h42a0b549, 32'h42a9a840, 32'h4273277d, 32'h422fbbb7, 32'hc238d9f7, 32'h420cc830, 32'hc2b0557f};
test_output[2152:2159] = '{32'h42a0bb47, 32'h42a0b549, 32'h42a9a840, 32'h4273277d, 32'h422fbbb7, 32'h0, 32'h420cc830, 32'h0};
test_input[2160:2167] = '{32'h41097753, 32'hc2a30c32, 32'hc16508e8, 32'h4232f95a, 32'h414061da, 32'h42c5a7c6, 32'h40274f71, 32'h42a930cd};
test_output[2160:2167] = '{32'h41097753, 32'h0, 32'h0, 32'h4232f95a, 32'h414061da, 32'h42c5a7c6, 32'h40274f71, 32'h42a930cd};
test_input[2168:2175] = '{32'hc294d0d1, 32'h42c1c5a2, 32'hc24c5086, 32'h3fa38686, 32'hc1754907, 32'h42444bdc, 32'h420e306a, 32'hc188db6f};
test_output[2168:2175] = '{32'h0, 32'h42c1c5a2, 32'h0, 32'h3fa38686, 32'h0, 32'h42444bdc, 32'h420e306a, 32'h0};
test_input[2176:2183] = '{32'h41cc0bd1, 32'hc01314b7, 32'hc2290e9c, 32'h42aaa4ad, 32'h42c3186c, 32'h40cb95b2, 32'h4292a35a, 32'hc21370f2};
test_output[2176:2183] = '{32'h41cc0bd1, 32'h0, 32'h0, 32'h42aaa4ad, 32'h42c3186c, 32'h40cb95b2, 32'h4292a35a, 32'h0};
test_input[2184:2191] = '{32'h423b211b, 32'h4293e3bf, 32'h3f2a341d, 32'hc28991fa, 32'hc2329125, 32'hc2c36986, 32'hc22389eb, 32'hc1ba2154};
test_output[2184:2191] = '{32'h423b211b, 32'h4293e3bf, 32'h3f2a341d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2192:2199] = '{32'h428900e4, 32'h42af49c9, 32'hc2c1ff0a, 32'h42a8102a, 32'h420eadd2, 32'h42b7936a, 32'h4109726e, 32'hc2677d82};
test_output[2192:2199] = '{32'h428900e4, 32'h42af49c9, 32'h0, 32'h42a8102a, 32'h420eadd2, 32'h42b7936a, 32'h4109726e, 32'h0};
test_input[2200:2207] = '{32'hc136f675, 32'hc2b6ef7f, 32'h427fdf6e, 32'h42bc4b47, 32'h428d574b, 32'h4106e8b6, 32'h42b2a434, 32'hc29f0068};
test_output[2200:2207] = '{32'h0, 32'h0, 32'h427fdf6e, 32'h42bc4b47, 32'h428d574b, 32'h4106e8b6, 32'h42b2a434, 32'h0};
test_input[2208:2215] = '{32'hc27d3e38, 32'hc2ad6f95, 32'hc2ae6e7d, 32'hc0555c5b, 32'h42b656b1, 32'h4248f44e, 32'hc1a61b02, 32'h41bafae1};
test_output[2208:2215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42b656b1, 32'h4248f44e, 32'h0, 32'h41bafae1};
test_input[2216:2223] = '{32'hc1b3c814, 32'hc1a95a9a, 32'hc23a517f, 32'h42b3952d, 32'h41ba1106, 32'hc1c9c7af, 32'hc28be144, 32'h42a1d49f};
test_output[2216:2223] = '{32'h0, 32'h0, 32'h0, 32'h42b3952d, 32'h41ba1106, 32'h0, 32'h0, 32'h42a1d49f};
test_input[2224:2231] = '{32'h41a84f82, 32'hc1aa6253, 32'h4192374c, 32'hc240686a, 32'h42464518, 32'hbffb0908, 32'hc2c5533d, 32'h429360fa};
test_output[2224:2231] = '{32'h41a84f82, 32'h0, 32'h4192374c, 32'h0, 32'h42464518, 32'h0, 32'h0, 32'h429360fa};
test_input[2232:2239] = '{32'h42209162, 32'h40cf390d, 32'h41c7caf0, 32'hc110b127, 32'hc28f3cc6, 32'h4289bdfd, 32'hc20a0061, 32'h4227d65e};
test_output[2232:2239] = '{32'h42209162, 32'h40cf390d, 32'h41c7caf0, 32'h0, 32'h0, 32'h4289bdfd, 32'h0, 32'h4227d65e};
test_input[2240:2247] = '{32'hc28f8266, 32'hc23bc973, 32'h428b1d1a, 32'hc2a6e958, 32'hc2185935, 32'hc0b1f2ba, 32'hc1cc50ef, 32'h42c36025};
test_output[2240:2247] = '{32'h0, 32'h0, 32'h428b1d1a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c36025};
test_input[2248:2255] = '{32'h423495bf, 32'hc29c5d23, 32'hc21b9faf, 32'hc2b7c898, 32'h4230d052, 32'hc2a10625, 32'h41be7c08, 32'hc0c6c57b};
test_output[2248:2255] = '{32'h423495bf, 32'h0, 32'h0, 32'h0, 32'h4230d052, 32'h0, 32'h41be7c08, 32'h0};
test_input[2256:2263] = '{32'hc0848b95, 32'h424e73b0, 32'hc113294e, 32'hc0b4f5e4, 32'h428f3898, 32'h426955d9, 32'h428dd202, 32'h42241c08};
test_output[2256:2263] = '{32'h0, 32'h424e73b0, 32'h0, 32'h0, 32'h428f3898, 32'h426955d9, 32'h428dd202, 32'h42241c08};
test_input[2264:2271] = '{32'h409e5983, 32'hc28bf201, 32'h41dd6c84, 32'h40fbe9c6, 32'h3ece8016, 32'h4253fb68, 32'hc26d21ae, 32'h428fb514};
test_output[2264:2271] = '{32'h409e5983, 32'h0, 32'h41dd6c84, 32'h40fbe9c6, 32'h3ece8016, 32'h4253fb68, 32'h0, 32'h428fb514};
test_input[2272:2279] = '{32'h429ff555, 32'h42712623, 32'h42c7b2d6, 32'h3f8289a5, 32'h426ce0bb, 32'hc2b8ec80, 32'h42b863fa, 32'h42a6bf1a};
test_output[2272:2279] = '{32'h429ff555, 32'h42712623, 32'h42c7b2d6, 32'h3f8289a5, 32'h426ce0bb, 32'h0, 32'h42b863fa, 32'h42a6bf1a};
test_input[2280:2287] = '{32'h42bb29a8, 32'h42718017, 32'hc29e095f, 32'hc2610735, 32'hc28bc959, 32'h4283334b, 32'h42795fdc, 32'h4296e6fd};
test_output[2280:2287] = '{32'h42bb29a8, 32'h42718017, 32'h0, 32'h0, 32'h0, 32'h4283334b, 32'h42795fdc, 32'h4296e6fd};
test_input[2288:2295] = '{32'h419db6da, 32'h4273e69a, 32'h42ab0829, 32'hc273ee3e, 32'h42960a29, 32'hc20ed4bd, 32'h421623c2, 32'hc19ee62b};
test_output[2288:2295] = '{32'h419db6da, 32'h4273e69a, 32'h42ab0829, 32'h0, 32'h42960a29, 32'h0, 32'h421623c2, 32'h0};
test_input[2296:2303] = '{32'hc20e67a2, 32'hbebde9e5, 32'hc267e844, 32'hc21b7157, 32'h421247d4, 32'h420f2c80, 32'hc28d22dc, 32'h42abafa8};
test_output[2296:2303] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h421247d4, 32'h420f2c80, 32'h0, 32'h42abafa8};
test_input[2304:2311] = '{32'hc272aff7, 32'hc1191ea1, 32'hc2589ae2, 32'h41aa9ab7, 32'hc25913ba, 32'h4183b8e5, 32'hc28cca92, 32'hc19fdb84};
test_output[2304:2311] = '{32'h0, 32'h0, 32'h0, 32'h41aa9ab7, 32'h0, 32'h4183b8e5, 32'h0, 32'h0};
test_input[2312:2319] = '{32'hc27323a7, 32'h40edad0c, 32'h423cb31a, 32'h4286048d, 32'h4236865b, 32'h427b9fba, 32'hbe1c1658, 32'hc21ac8b4};
test_output[2312:2319] = '{32'h0, 32'h40edad0c, 32'h423cb31a, 32'h4286048d, 32'h4236865b, 32'h427b9fba, 32'h0, 32'h0};
test_input[2320:2327] = '{32'hc2a3f012, 32'h424a8b8b, 32'hc29b6ad4, 32'h429dc358, 32'h4286a007, 32'hc1b2c8d4, 32'h4294014c, 32'hc2795259};
test_output[2320:2327] = '{32'h0, 32'h424a8b8b, 32'h0, 32'h429dc358, 32'h4286a007, 32'h0, 32'h4294014c, 32'h0};
test_input[2328:2335] = '{32'h42ab10eb, 32'h4253387b, 32'h42a8648b, 32'h42a26921, 32'h4282a976, 32'hc22a02db, 32'hc1540a6f, 32'h418063a0};
test_output[2328:2335] = '{32'h42ab10eb, 32'h4253387b, 32'h42a8648b, 32'h42a26921, 32'h4282a976, 32'h0, 32'h0, 32'h418063a0};
test_input[2336:2343] = '{32'h4179e1b0, 32'hc237ff38, 32'h424259ef, 32'h41b6a994, 32'h42a95652, 32'hc2b14d94, 32'h427f2873, 32'hc2a338a2};
test_output[2336:2343] = '{32'h4179e1b0, 32'h0, 32'h424259ef, 32'h41b6a994, 32'h42a95652, 32'h0, 32'h427f2873, 32'h0};
test_input[2344:2351] = '{32'hc20048a0, 32'hc20d6c60, 32'h425facc6, 32'hc1bf5b2e, 32'h42b36727, 32'h422d5186, 32'hc1799450, 32'hc209fa76};
test_output[2344:2351] = '{32'h0, 32'h0, 32'h425facc6, 32'h0, 32'h42b36727, 32'h422d5186, 32'h0, 32'h0};
test_input[2352:2359] = '{32'hc2081888, 32'hc2817b2a, 32'h42ab54a9, 32'h42223523, 32'h41edc91b, 32'h4289b215, 32'hc2a68f68, 32'hc2b33b49};
test_output[2352:2359] = '{32'h0, 32'h0, 32'h42ab54a9, 32'h42223523, 32'h41edc91b, 32'h4289b215, 32'h0, 32'h0};
test_input[2360:2367] = '{32'h41c8a158, 32'hc1f35fe7, 32'hc2b0e467, 32'hc2b5a6c4, 32'hc10f3a08, 32'h401bb4dc, 32'hc0a46e36, 32'h42584a03};
test_output[2360:2367] = '{32'h41c8a158, 32'h0, 32'h0, 32'h0, 32'h0, 32'h401bb4dc, 32'h0, 32'h42584a03};
test_input[2368:2375] = '{32'hc2252285, 32'h42b27194, 32'hc1141f86, 32'h41b75c7d, 32'hc1fb5f50, 32'h42bce873, 32'h42987bf5, 32'hc27fea72};
test_output[2368:2375] = '{32'h0, 32'h42b27194, 32'h0, 32'h41b75c7d, 32'h0, 32'h42bce873, 32'h42987bf5, 32'h0};
test_input[2376:2383] = '{32'hbf254987, 32'h417abe2f, 32'h42c2d856, 32'hc0debb9d, 32'h41e2ac41, 32'h41181586, 32'hc277d189, 32'h42693a19};
test_output[2376:2383] = '{32'h0, 32'h417abe2f, 32'h42c2d856, 32'h0, 32'h41e2ac41, 32'h41181586, 32'h0, 32'h42693a19};
test_input[2384:2391] = '{32'h41be953a, 32'h41f6f669, 32'hc293619e, 32'h42b378c4, 32'hc230f57e, 32'h42c215bd, 32'hc29e6c31, 32'hc1ff4cd0};
test_output[2384:2391] = '{32'h41be953a, 32'h41f6f669, 32'h0, 32'h42b378c4, 32'h0, 32'h42c215bd, 32'h0, 32'h0};
test_input[2392:2399] = '{32'h42278b1c, 32'hbf4c3ef2, 32'h4249cd6e, 32'hc26cde35, 32'h421a524a, 32'hc2ae1573, 32'h41feda41, 32'hc2b8e18d};
test_output[2392:2399] = '{32'h42278b1c, 32'h0, 32'h4249cd6e, 32'h0, 32'h421a524a, 32'h0, 32'h41feda41, 32'h0};
test_input[2400:2407] = '{32'h4294ac10, 32'hc1b892fe, 32'hc2a52fbb, 32'h4182bb32, 32'h428b8ef1, 32'hc27c2471, 32'hc249110f, 32'h4243cf09};
test_output[2400:2407] = '{32'h4294ac10, 32'h0, 32'h0, 32'h4182bb32, 32'h428b8ef1, 32'h0, 32'h0, 32'h4243cf09};
test_input[2408:2415] = '{32'h424354fb, 32'h4248c526, 32'h42055fcc, 32'hc1e4e5fe, 32'hc2147fd9, 32'hc101199c, 32'hc25b01e1, 32'h41f90e64};
test_output[2408:2415] = '{32'h424354fb, 32'h4248c526, 32'h42055fcc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f90e64};
test_input[2416:2423] = '{32'h425823ed, 32'hc0c51c86, 32'hc20b0358, 32'h42b1711c, 32'hc2bd36ef, 32'hc0ce3cf2, 32'h4270ce7a, 32'hc2417124};
test_output[2416:2423] = '{32'h425823ed, 32'h0, 32'h0, 32'h42b1711c, 32'h0, 32'h0, 32'h4270ce7a, 32'h0};
test_input[2424:2431] = '{32'hc2bf0ab8, 32'h41c14058, 32'h415b9173, 32'hc2379a6e, 32'h420fb1d7, 32'h425d22d3, 32'h425f3fcb, 32'h42366d21};
test_output[2424:2431] = '{32'h0, 32'h41c14058, 32'h415b9173, 32'h0, 32'h420fb1d7, 32'h425d22d3, 32'h425f3fcb, 32'h42366d21};
test_input[2432:2439] = '{32'hc2be8bc6, 32'h428192b7, 32'h42afb250, 32'h42b08e51, 32'hc26b31e4, 32'hc12665e9, 32'h42ad1cc9, 32'h423cd8af};
test_output[2432:2439] = '{32'h0, 32'h428192b7, 32'h42afb250, 32'h42b08e51, 32'h0, 32'h0, 32'h42ad1cc9, 32'h423cd8af};
test_input[2440:2447] = '{32'hc215ef37, 32'hc1de1c10, 32'hc0450d1a, 32'h3e1d58b8, 32'h427e13a9, 32'h41d6c95e, 32'h41a181d4, 32'hc1bc7eb6};
test_output[2440:2447] = '{32'h0, 32'h0, 32'h0, 32'h3e1d58b8, 32'h427e13a9, 32'h41d6c95e, 32'h41a181d4, 32'h0};
test_input[2448:2455] = '{32'hc255cedc, 32'hc1311ca1, 32'hc239378e, 32'hc12d21d4, 32'hc2189473, 32'hc1a2161e, 32'h4255daf6, 32'h4280874b};
test_output[2448:2455] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4255daf6, 32'h4280874b};
test_input[2456:2463] = '{32'h42887aa3, 32'h429fc0e8, 32'hc2b085e0, 32'h41d7bb51, 32'hc25f5b7e, 32'h42c3618f, 32'hbfe064d4, 32'h42447668};
test_output[2456:2463] = '{32'h42887aa3, 32'h429fc0e8, 32'h0, 32'h41d7bb51, 32'h0, 32'h42c3618f, 32'h0, 32'h42447668};
test_input[2464:2471] = '{32'hc2b86068, 32'hc27f8057, 32'hc221527f, 32'hc24ad589, 32'h424e5255, 32'h42a3f0d1, 32'hc1387e69, 32'h40f7ada7};
test_output[2464:2471] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h424e5255, 32'h42a3f0d1, 32'h0, 32'h40f7ada7};
test_input[2472:2479] = '{32'hc2b9b397, 32'hc211de6c, 32'hc1d22ea2, 32'hc2b7a11c, 32'hc1e45ab8, 32'hc2b86dbd, 32'hc2093d37, 32'hc1ce57aa};
test_output[2472:2479] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2480:2487] = '{32'hc139739c, 32'h429a20c9, 32'h428c4721, 32'hc2bf22a0, 32'h42b6f301, 32'hc083237b, 32'hc2ac6bbd, 32'h42a963b4};
test_output[2480:2487] = '{32'h0, 32'h429a20c9, 32'h428c4721, 32'h0, 32'h42b6f301, 32'h0, 32'h0, 32'h42a963b4};
test_input[2488:2495] = '{32'h4221dd75, 32'hc153c89b, 32'hc1673ddb, 32'hc208ae5c, 32'hc28fcfde, 32'h42731fe6, 32'hc27b7887, 32'hc1afa689};
test_output[2488:2495] = '{32'h4221dd75, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42731fe6, 32'h0, 32'h0};
test_input[2496:2503] = '{32'hc28cb4f8, 32'h41993a40, 32'h412b6ede, 32'hc13bc3ef, 32'h42826582, 32'hc25c0682, 32'hc16f490e, 32'h428be3b2};
test_output[2496:2503] = '{32'h0, 32'h41993a40, 32'h412b6ede, 32'h0, 32'h42826582, 32'h0, 32'h0, 32'h428be3b2};
test_input[2504:2511] = '{32'h41fc3f63, 32'h42819f97, 32'h429a5963, 32'h4293a5b8, 32'h42a05573, 32'hc2144978, 32'hc200423c, 32'hc1c27188};
test_output[2504:2511] = '{32'h41fc3f63, 32'h42819f97, 32'h429a5963, 32'h4293a5b8, 32'h42a05573, 32'h0, 32'h0, 32'h0};
test_input[2512:2519] = '{32'hc1add886, 32'hc2be640a, 32'h42c2af9b, 32'hc1f80ec1, 32'hc2b8562b, 32'h42c331dd, 32'h41a42e15, 32'hc26c909a};
test_output[2512:2519] = '{32'h0, 32'h0, 32'h42c2af9b, 32'h0, 32'h0, 32'h42c331dd, 32'h41a42e15, 32'h0};
test_input[2520:2527] = '{32'h424d5f1a, 32'hc13c7e3d, 32'h416efe15, 32'h42ae54ec, 32'hc2627ec9, 32'hc2a17218, 32'hc28b557a, 32'h420872ce};
test_output[2520:2527] = '{32'h424d5f1a, 32'h0, 32'h416efe15, 32'h42ae54ec, 32'h0, 32'h0, 32'h0, 32'h420872ce};
test_input[2528:2535] = '{32'h428a77cd, 32'h42210b17, 32'h4024696a, 32'hc1d202f1, 32'h420cdc4e, 32'hc21bdbca, 32'h41e3eb1f, 32'h427c752a};
test_output[2528:2535] = '{32'h428a77cd, 32'h42210b17, 32'h4024696a, 32'h0, 32'h420cdc4e, 32'h0, 32'h41e3eb1f, 32'h427c752a};
test_input[2536:2543] = '{32'h41179dcb, 32'hc1e72d6e, 32'hc2abdefc, 32'hc261f580, 32'hc2bdeeee, 32'hc29e7f37, 32'hc26885a5, 32'h4220ed40};
test_output[2536:2543] = '{32'h41179dcb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4220ed40};
test_input[2544:2551] = '{32'hc27e6ace, 32'h41b87b95, 32'h429ef73e, 32'hc2973fef, 32'h42340c5b, 32'hc2a29f74, 32'hc2536ea6, 32'hc12669ab};
test_output[2544:2551] = '{32'h0, 32'h41b87b95, 32'h429ef73e, 32'h0, 32'h42340c5b, 32'h0, 32'h0, 32'h0};
test_input[2552:2559] = '{32'hc236227e, 32'hc20d07e2, 32'hc25d8248, 32'h41ccf80b, 32'h4217cef0, 32'h4284ce22, 32'hc1d39834, 32'h41e1b9d4};
test_output[2552:2559] = '{32'h0, 32'h0, 32'h0, 32'h41ccf80b, 32'h4217cef0, 32'h4284ce22, 32'h0, 32'h41e1b9d4};
test_input[2560:2567] = '{32'hc071899a, 32'h420ce3dd, 32'hc1bacf18, 32'h41852a04, 32'hc1a8dac5, 32'h42b346c8, 32'hc1d4e456, 32'h422a97a6};
test_output[2560:2567] = '{32'h0, 32'h420ce3dd, 32'h0, 32'h41852a04, 32'h0, 32'h42b346c8, 32'h0, 32'h422a97a6};
test_input[2568:2575] = '{32'hc27c2bec, 32'h4267e2af, 32'h42ada625, 32'hc25b485d, 32'h41951e16, 32'hc29f2edf, 32'hc00dfd46, 32'hc2a0b4d1};
test_output[2568:2575] = '{32'h0, 32'h4267e2af, 32'h42ada625, 32'h0, 32'h41951e16, 32'h0, 32'h0, 32'h0};
test_input[2576:2583] = '{32'h4170f79a, 32'hc1065e96, 32'hc20464a1, 32'hc1cb1d80, 32'hc1909c6f, 32'h42ae0003, 32'h426bc533, 32'h4293433c};
test_output[2576:2583] = '{32'h4170f79a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ae0003, 32'h426bc533, 32'h4293433c};
test_input[2584:2591] = '{32'hc29f3fa7, 32'h426b227d, 32'hc28fc22b, 32'h425f579f, 32'hc290de60, 32'hc2c21a6a, 32'h4275d0f8, 32'hc176c1fa};
test_output[2584:2591] = '{32'h0, 32'h426b227d, 32'h0, 32'h425f579f, 32'h0, 32'h0, 32'h4275d0f8, 32'h0};
test_input[2592:2599] = '{32'hc210b841, 32'h410f4e5f, 32'h42af3a5f, 32'h42724aac, 32'h42b0df8d, 32'h42c08c63, 32'hc27fb780, 32'hc188587b};
test_output[2592:2599] = '{32'h0, 32'h410f4e5f, 32'h42af3a5f, 32'h42724aac, 32'h42b0df8d, 32'h42c08c63, 32'h0, 32'h0};
test_input[2600:2607] = '{32'h410a2238, 32'hc27dec6e, 32'hc2934ab9, 32'h40e4b65a, 32'h42c0583b, 32'h4100c3eb, 32'hc26b72bd, 32'h4295fca5};
test_output[2600:2607] = '{32'h410a2238, 32'h0, 32'h0, 32'h40e4b65a, 32'h42c0583b, 32'h4100c3eb, 32'h0, 32'h4295fca5};
test_input[2608:2615] = '{32'h4218826a, 32'h41be0847, 32'hc2ab053e, 32'h41ce4338, 32'hc23e0f14, 32'hc1cafa8f, 32'hc2bb11d2, 32'hc22e5954};
test_output[2608:2615] = '{32'h4218826a, 32'h41be0847, 32'h0, 32'h41ce4338, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2616:2623] = '{32'h425bc336, 32'h419e94fc, 32'hc224c80a, 32'h3f4945aa, 32'h42005109, 32'h41d667ee, 32'h40b77aca, 32'hc29b9d94};
test_output[2616:2623] = '{32'h425bc336, 32'h419e94fc, 32'h0, 32'h3f4945aa, 32'h42005109, 32'h41d667ee, 32'h40b77aca, 32'h0};
test_input[2624:2631] = '{32'hc2ad1d82, 32'h413cba5e, 32'h41d717ee, 32'h422e0e5c, 32'hc24f0b68, 32'hc0dbafa1, 32'hc1fd3237, 32'h40d790d6};
test_output[2624:2631] = '{32'h0, 32'h413cba5e, 32'h41d717ee, 32'h422e0e5c, 32'h0, 32'h0, 32'h0, 32'h40d790d6};
test_input[2632:2639] = '{32'h429c181d, 32'hc289268e, 32'h41109a02, 32'h410fd275, 32'h41fb33d5, 32'hc222b430, 32'h423aca58, 32'h426115c1};
test_output[2632:2639] = '{32'h429c181d, 32'h0, 32'h41109a02, 32'h410fd275, 32'h41fb33d5, 32'h0, 32'h423aca58, 32'h426115c1};
test_input[2640:2647] = '{32'hc2982c7c, 32'hc155cd8b, 32'h429a6925, 32'h423b8ff3, 32'h426a73a1, 32'h429d7977, 32'h414d2f8d, 32'h42441a0c};
test_output[2640:2647] = '{32'h0, 32'h0, 32'h429a6925, 32'h423b8ff3, 32'h426a73a1, 32'h429d7977, 32'h414d2f8d, 32'h42441a0c};
test_input[2648:2655] = '{32'h422d74e8, 32'h414e95fc, 32'h415d8040, 32'h42628b21, 32'h402b7332, 32'hc258c644, 32'h42c2961e, 32'hbfccd0ac};
test_output[2648:2655] = '{32'h422d74e8, 32'h414e95fc, 32'h415d8040, 32'h42628b21, 32'h402b7332, 32'h0, 32'h42c2961e, 32'h0};
test_input[2656:2663] = '{32'hc2947d0c, 32'h42a8ec0d, 32'h42c45e05, 32'h4240601f, 32'h429e3f3a, 32'h42bbc9a6, 32'h3ff87cf8, 32'hc28db940};
test_output[2656:2663] = '{32'h0, 32'h42a8ec0d, 32'h42c45e05, 32'h4240601f, 32'h429e3f3a, 32'h42bbc9a6, 32'h3ff87cf8, 32'h0};
test_input[2664:2671] = '{32'h42ab035a, 32'hc228e46a, 32'h40cf134d, 32'hc265099b, 32'hc260c670, 32'h41151ec1, 32'hc29012d8, 32'hc2c0a646};
test_output[2664:2671] = '{32'h42ab035a, 32'h0, 32'h40cf134d, 32'h0, 32'h0, 32'h41151ec1, 32'h0, 32'h0};
test_input[2672:2679] = '{32'hc20715c2, 32'h413eeea3, 32'h423133eb, 32'h429f6cf0, 32'hc25d98aa, 32'h41ef8a70, 32'hc2287cac, 32'hc1644472};
test_output[2672:2679] = '{32'h0, 32'h413eeea3, 32'h423133eb, 32'h429f6cf0, 32'h0, 32'h41ef8a70, 32'h0, 32'h0};
test_input[2680:2687] = '{32'hc279d1c7, 32'hc27bd0ce, 32'hc287efcd, 32'hc2b52ca6, 32'hc2882a16, 32'h428960c2, 32'h42841d31, 32'h4268856f};
test_output[2680:2687] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428960c2, 32'h42841d31, 32'h4268856f};
test_input[2688:2695] = '{32'h41583a41, 32'h4279d240, 32'hc22deb93, 32'hc1d4d955, 32'hbfd13d83, 32'h4293e4c3, 32'h424d89ea, 32'hc29aba95};
test_output[2688:2695] = '{32'h41583a41, 32'h4279d240, 32'h0, 32'h0, 32'h0, 32'h4293e4c3, 32'h424d89ea, 32'h0};
test_input[2696:2703] = '{32'hc2799839, 32'hc224eb8c, 32'hc16a7924, 32'hc2b01504, 32'h426a33f4, 32'h427d4421, 32'h42794413, 32'h42312c3f};
test_output[2696:2703] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h426a33f4, 32'h427d4421, 32'h42794413, 32'h42312c3f};
test_input[2704:2711] = '{32'h42a94f76, 32'h42553532, 32'h4187ac5c, 32'hc208b6f1, 32'h412745e2, 32'hc016fec7, 32'h42571e65, 32'h41f80483};
test_output[2704:2711] = '{32'h42a94f76, 32'h42553532, 32'h4187ac5c, 32'h0, 32'h412745e2, 32'h0, 32'h42571e65, 32'h41f80483};
test_input[2712:2719] = '{32'h42a14e0c, 32'h4229c99b, 32'h4286e2ee, 32'hc274a194, 32'hc21a9f0c, 32'h412a158d, 32'h42224939, 32'hbffba290};
test_output[2712:2719] = '{32'h42a14e0c, 32'h4229c99b, 32'h4286e2ee, 32'h0, 32'h0, 32'h412a158d, 32'h42224939, 32'h0};
test_input[2720:2727] = '{32'h4230858c, 32'h42054b57, 32'hc250d4cc, 32'hc2c2f9b9, 32'h42b10c1b, 32'h42c69584, 32'h41096f27, 32'hc1dbf160};
test_output[2720:2727] = '{32'h4230858c, 32'h42054b57, 32'h0, 32'h0, 32'h42b10c1b, 32'h42c69584, 32'h41096f27, 32'h0};
test_input[2728:2735] = '{32'hc20194b3, 32'h4286a8f5, 32'hc1b0b761, 32'h41e8e507, 32'hc2880675, 32'hc2c6bfab, 32'hc298d035, 32'hc281a816};
test_output[2728:2735] = '{32'h0, 32'h4286a8f5, 32'h0, 32'h41e8e507, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2736:2743] = '{32'hc1a1e9e9, 32'h42b493d1, 32'hc28650d5, 32'hc27e8c9b, 32'h41e203d6, 32'h41ea1448, 32'h42094d8c, 32'hc2afa0c2};
test_output[2736:2743] = '{32'h0, 32'h42b493d1, 32'h0, 32'h0, 32'h41e203d6, 32'h41ea1448, 32'h42094d8c, 32'h0};
test_input[2744:2751] = '{32'hc2c3d106, 32'hc14482d3, 32'hc0bdebb7, 32'h41a583a5, 32'hc1acd18b, 32'h428aaefa, 32'h42b3897a, 32'hc18c50d5};
test_output[2744:2751] = '{32'h0, 32'h0, 32'h0, 32'h41a583a5, 32'h0, 32'h428aaefa, 32'h42b3897a, 32'h0};
test_input[2752:2759] = '{32'h424f872e, 32'hc2627f28, 32'hc2602dc8, 32'h42a7803c, 32'h4268fceb, 32'h426a6ca8, 32'hc2995647, 32'h4118630c};
test_output[2752:2759] = '{32'h424f872e, 32'h0, 32'h0, 32'h42a7803c, 32'h4268fceb, 32'h426a6ca8, 32'h0, 32'h4118630c};
test_input[2760:2767] = '{32'hc19b73e0, 32'hc26a8aac, 32'hc27178ef, 32'h41d97672, 32'hc231739a, 32'h41a7e483, 32'hc16fb7d7, 32'hc28c24f0};
test_output[2760:2767] = '{32'h0, 32'h0, 32'h0, 32'h41d97672, 32'h0, 32'h41a7e483, 32'h0, 32'h0};
test_input[2768:2775] = '{32'h42873909, 32'hc283bec4, 32'h4268129a, 32'hc29f1130, 32'hc1b6b7ac, 32'h428d5f95, 32'hc2888983, 32'h41bfc4db};
test_output[2768:2775] = '{32'h42873909, 32'h0, 32'h4268129a, 32'h0, 32'h0, 32'h428d5f95, 32'h0, 32'h41bfc4db};
test_input[2776:2783] = '{32'h426a1ca4, 32'hc27f5322, 32'h41918976, 32'hc27a26b4, 32'hc210a92b, 32'h42819ff5, 32'hc13b6543, 32'h42435c48};
test_output[2776:2783] = '{32'h426a1ca4, 32'h0, 32'h41918976, 32'h0, 32'h0, 32'h42819ff5, 32'h0, 32'h42435c48};
test_input[2784:2791] = '{32'hc2918a50, 32'h41e4694e, 32'hc13669fc, 32'hc2b81969, 32'hc2bd8cbf, 32'hc1dddc0e, 32'hc2c32e01, 32'hc1a9edff};
test_output[2784:2791] = '{32'h0, 32'h41e4694e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[2792:2799] = '{32'hc0a01810, 32'hc1b38a39, 32'hc189fa57, 32'h4208329a, 32'h42aa2823, 32'hc2948e53, 32'h42bf7524, 32'hc225b685};
test_output[2792:2799] = '{32'h0, 32'h0, 32'h0, 32'h4208329a, 32'h42aa2823, 32'h0, 32'h42bf7524, 32'h0};
test_input[2800:2807] = '{32'h429cfa47, 32'hc25d0564, 32'hc2c78687, 32'h4289eb86, 32'h40d128b9, 32'h415c9a29, 32'h3fec2121, 32'h419c6cf9};
test_output[2800:2807] = '{32'h429cfa47, 32'h0, 32'h0, 32'h4289eb86, 32'h40d128b9, 32'h415c9a29, 32'h3fec2121, 32'h419c6cf9};
test_input[2808:2815] = '{32'hc1edc8aa, 32'hc2c1ba5e, 32'hc23f1b8a, 32'hc288644b, 32'h415b1505, 32'h41b61370, 32'hc2c78a6b, 32'hc203855a};
test_output[2808:2815] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h415b1505, 32'h41b61370, 32'h0, 32'h0};
test_input[2816:2823] = '{32'h4272972d, 32'h41861764, 32'hc2bec4c2, 32'h42b16d5a, 32'hc2c10a5b, 32'hc273f389, 32'hc29ae9e5, 32'h4168d0b6};
test_output[2816:2823] = '{32'h4272972d, 32'h41861764, 32'h0, 32'h42b16d5a, 32'h0, 32'h0, 32'h0, 32'h4168d0b6};
test_input[2824:2831] = '{32'hc29e0653, 32'hc22c919e, 32'hc126db12, 32'h42823513, 32'h426c4ebf, 32'h42a55b3b, 32'hc28e413b, 32'hc2c77292};
test_output[2824:2831] = '{32'h0, 32'h0, 32'h0, 32'h42823513, 32'h426c4ebf, 32'h42a55b3b, 32'h0, 32'h0};
test_input[2832:2839] = '{32'h4106b4f8, 32'h428e81a0, 32'hc2827651, 32'h42be18f9, 32'hc0eb8b81, 32'hc27cee6b, 32'hc107b45b, 32'h419377e8};
test_output[2832:2839] = '{32'h4106b4f8, 32'h428e81a0, 32'h0, 32'h42be18f9, 32'h0, 32'h0, 32'h0, 32'h419377e8};
test_input[2840:2847] = '{32'hc2012070, 32'hc24c822d, 32'hc254cdac, 32'hc065eaee, 32'h42aecbc0, 32'h40fece88, 32'hc2a0ea6b, 32'h41c088a3};
test_output[2840:2847] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42aecbc0, 32'h40fece88, 32'h0, 32'h41c088a3};
test_input[2848:2855] = '{32'hc2b369e0, 32'h413c38a0, 32'h4214f550, 32'hc28fed3f, 32'hc28742e7, 32'h4242780f, 32'hc23a0301, 32'hc263879f};
test_output[2848:2855] = '{32'h0, 32'h413c38a0, 32'h4214f550, 32'h0, 32'h0, 32'h4242780f, 32'h0, 32'h0};
test_input[2856:2863] = '{32'hc19372cd, 32'h413a422e, 32'h420bf5c2, 32'h4294e665, 32'hc2b8aa6b, 32'hc28187eb, 32'h42866870, 32'h425d5388};
test_output[2856:2863] = '{32'h0, 32'h413a422e, 32'h420bf5c2, 32'h4294e665, 32'h0, 32'h0, 32'h42866870, 32'h425d5388};
test_input[2864:2871] = '{32'hc1ce31a7, 32'h404c0ef7, 32'h42921a56, 32'h42b3918c, 32'hc2c08bcc, 32'hc2be84e4, 32'hc1af6789, 32'h41ed03d3};
test_output[2864:2871] = '{32'h0, 32'h404c0ef7, 32'h42921a56, 32'h42b3918c, 32'h0, 32'h0, 32'h0, 32'h41ed03d3};
test_input[2872:2879] = '{32'h42b9a064, 32'hc26f45d0, 32'hc20d8dc7, 32'h422af8b7, 32'h41c56a21, 32'hc16a2ef4, 32'h427bdf36, 32'h41bbcc84};
test_output[2872:2879] = '{32'h42b9a064, 32'h0, 32'h0, 32'h422af8b7, 32'h41c56a21, 32'h0, 32'h427bdf36, 32'h41bbcc84};
test_input[2880:2887] = '{32'hc26b41dc, 32'hc297070b, 32'h429979b8, 32'h42919675, 32'hc238b6d5, 32'hc158ac25, 32'h402ab915, 32'hc2505a99};
test_output[2880:2887] = '{32'h0, 32'h0, 32'h429979b8, 32'h42919675, 32'h0, 32'h0, 32'h402ab915, 32'h0};
test_input[2888:2895] = '{32'hc1508812, 32'h428c26f9, 32'h4176ea61, 32'hc2a4c28c, 32'hc29f064f, 32'h408ab123, 32'h41c46b76, 32'hc219e547};
test_output[2888:2895] = '{32'h0, 32'h428c26f9, 32'h4176ea61, 32'h0, 32'h0, 32'h408ab123, 32'h41c46b76, 32'h0};
test_input[2896:2903] = '{32'hc2ae1d90, 32'h42bdb76d, 32'hc1f108ab, 32'hc2c024e6, 32'h4284c471, 32'hc2a6a510, 32'hc2361b82, 32'hbf3ee124};
test_output[2896:2903] = '{32'h0, 32'h42bdb76d, 32'h0, 32'h0, 32'h4284c471, 32'h0, 32'h0, 32'h0};
test_input[2904:2911] = '{32'h4081faf6, 32'hc236b6d5, 32'hc2a6cffd, 32'hc1456f90, 32'h42c0340f, 32'hc2484d03, 32'h4031c25a, 32'h42c7ca23};
test_output[2904:2911] = '{32'h4081faf6, 32'h0, 32'h0, 32'h0, 32'h42c0340f, 32'h0, 32'h4031c25a, 32'h42c7ca23};
test_input[2912:2919] = '{32'hc0a33d81, 32'hc220d600, 32'hc2bf25f4, 32'h42b7f231, 32'hc2b22c8e, 32'hc2afbe01, 32'h42257b9f, 32'hc2931811};
test_output[2912:2919] = '{32'h0, 32'h0, 32'h0, 32'h42b7f231, 32'h0, 32'h0, 32'h42257b9f, 32'h0};
test_input[2920:2927] = '{32'hc28f8ad8, 32'h41eec1d1, 32'h41d65663, 32'hc26021bb, 32'hc2b473ef, 32'h4298b8f8, 32'hc2aa433f, 32'hc2a8a68d};
test_output[2920:2927] = '{32'h0, 32'h41eec1d1, 32'h41d65663, 32'h0, 32'h0, 32'h4298b8f8, 32'h0, 32'h0};
test_input[2928:2935] = '{32'hc28bb5a4, 32'hc141a38f, 32'hc284a845, 32'hc2c6e10b, 32'hc2b6fa7d, 32'h4018bea5, 32'h41341d4a, 32'hc20ae399};
test_output[2928:2935] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4018bea5, 32'h41341d4a, 32'h0};
test_input[2936:2943] = '{32'h4205e6a3, 32'hc2b1f075, 32'hc2b35249, 32'hc196c61f, 32'hc2a2963e, 32'hc1b1182d, 32'h41458ad6, 32'h4249e3df};
test_output[2936:2943] = '{32'h4205e6a3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41458ad6, 32'h4249e3df};
test_input[2944:2951] = '{32'hc2a1f12a, 32'hc2acc3ad, 32'h429dc395, 32'h424e0cae, 32'hc142b200, 32'h428ddd02, 32'h4189974b, 32'hc2ba511d};
test_output[2944:2951] = '{32'h0, 32'h0, 32'h429dc395, 32'h424e0cae, 32'h0, 32'h428ddd02, 32'h4189974b, 32'h0};
test_input[2952:2959] = '{32'h42292418, 32'h4299a7e9, 32'h421c08c8, 32'hc27a6f9d, 32'h42377fd7, 32'h42c24abe, 32'h421c4aa5, 32'hc1c27013};
test_output[2952:2959] = '{32'h42292418, 32'h4299a7e9, 32'h421c08c8, 32'h0, 32'h42377fd7, 32'h42c24abe, 32'h421c4aa5, 32'h0};
test_input[2960:2967] = '{32'h42001138, 32'h426749d5, 32'h422bb38b, 32'hc281f067, 32'h41efbefe, 32'hc21ae276, 32'hc285b80c, 32'hc28eb334};
test_output[2960:2967] = '{32'h42001138, 32'h426749d5, 32'h422bb38b, 32'h0, 32'h41efbefe, 32'h0, 32'h0, 32'h0};
test_input[2968:2975] = '{32'hc289f178, 32'hc2348d22, 32'h41105471, 32'h4237c7f5, 32'hc2c7d7cb, 32'h4229a4e7, 32'hc288cc63, 32'hc2b8e646};
test_output[2968:2975] = '{32'h0, 32'h0, 32'h41105471, 32'h4237c7f5, 32'h0, 32'h4229a4e7, 32'h0, 32'h0};
test_input[2976:2983] = '{32'h429dae84, 32'hc13143e9, 32'h429ddfa1, 32'h423e5ebd, 32'hc25ff42d, 32'hc22d01ff, 32'h42001b47, 32'h423fbb49};
test_output[2976:2983] = '{32'h429dae84, 32'h0, 32'h429ddfa1, 32'h423e5ebd, 32'h0, 32'h0, 32'h42001b47, 32'h423fbb49};
test_input[2984:2991] = '{32'hc2c22988, 32'hc21fd08b, 32'hc299cb6c, 32'h422ece8c, 32'h429950be, 32'h421a5515, 32'hc2846f23, 32'hc20b9cba};
test_output[2984:2991] = '{32'h0, 32'h0, 32'h0, 32'h422ece8c, 32'h429950be, 32'h421a5515, 32'h0, 32'h0};
test_input[2992:2999] = '{32'h418237c2, 32'hc076f8dc, 32'hc1c597ef, 32'h421c593e, 32'hc29f659d, 32'hc0e95891, 32'hc23fcddd, 32'hc2883be0};
test_output[2992:2999] = '{32'h418237c2, 32'h0, 32'h0, 32'h421c593e, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3000:3007] = '{32'h40a3e65d, 32'hc1709012, 32'hc1ff65af, 32'hc2562adc, 32'hc295d70a, 32'h428d3731, 32'h4244c1a1, 32'hc2a9a061};
test_output[3000:3007] = '{32'h40a3e65d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428d3731, 32'h4244c1a1, 32'h0};
test_input[3008:3015] = '{32'h3f6461c3, 32'hc10d5d01, 32'hc243a2f2, 32'h41fd70f0, 32'h429cfa61, 32'hc0fbb77f, 32'h429e8386, 32'hc1569cb5};
test_output[3008:3015] = '{32'h3f6461c3, 32'h0, 32'h0, 32'h41fd70f0, 32'h429cfa61, 32'h0, 32'h429e8386, 32'h0};
test_input[3016:3023] = '{32'hc29bf235, 32'hc1846c90, 32'h42a324b3, 32'h42aa8ef8, 32'hc24f9241, 32'hc1baa1c3, 32'hc27fdeb2, 32'h42aed5bf};
test_output[3016:3023] = '{32'h0, 32'h0, 32'h42a324b3, 32'h42aa8ef8, 32'h0, 32'h0, 32'h0, 32'h42aed5bf};
test_input[3024:3031] = '{32'h4248b7b1, 32'hc28e46d0, 32'hc2031d0b, 32'hc2a14835, 32'hc2401ff0, 32'h42a0b04d, 32'hc25b3340, 32'hc1996c72};
test_output[3024:3031] = '{32'h4248b7b1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a0b04d, 32'h0, 32'h0};
test_input[3032:3039] = '{32'h403cbf7e, 32'h42b87194, 32'h42699bc9, 32'h42b6e612, 32'h41ce1402, 32'hc223c255, 32'hc1d08337, 32'hc28df24f};
test_output[3032:3039] = '{32'h403cbf7e, 32'h42b87194, 32'h42699bc9, 32'h42b6e612, 32'h41ce1402, 32'h0, 32'h0, 32'h0};
test_input[3040:3047] = '{32'h4208b337, 32'hc242d517, 32'h4292f231, 32'hc260f883, 32'hc0a3ea72, 32'h42bc0261, 32'h42ad08b6, 32'h425b691f};
test_output[3040:3047] = '{32'h4208b337, 32'h0, 32'h4292f231, 32'h0, 32'h0, 32'h42bc0261, 32'h42ad08b6, 32'h425b691f};
test_input[3048:3055] = '{32'h42889b38, 32'h42a0cb29, 32'h4290b7bc, 32'hc22fd98d, 32'h42b7c505, 32'hc127fbab, 32'hc2319c5d, 32'hbf32b3fd};
test_output[3048:3055] = '{32'h42889b38, 32'h42a0cb29, 32'h4290b7bc, 32'h0, 32'h42b7c505, 32'h0, 32'h0, 32'h0};
test_input[3056:3063] = '{32'hc2afcdc8, 32'h3f9bb32b, 32'hc2b9a20c, 32'hc2a43bae, 32'h42a6a1bc, 32'h41b9dc21, 32'hc1f58106, 32'h4117d699};
test_output[3056:3063] = '{32'h0, 32'h3f9bb32b, 32'h0, 32'h0, 32'h42a6a1bc, 32'h41b9dc21, 32'h0, 32'h4117d699};
test_input[3064:3071] = '{32'hc1cbe7d4, 32'h421362f9, 32'h412623f0, 32'hc2aa3fe0, 32'h41191eb4, 32'hc1671e04, 32'h41759d34, 32'hc2256f6e};
test_output[3064:3071] = '{32'h0, 32'h421362f9, 32'h412623f0, 32'h0, 32'h41191eb4, 32'h0, 32'h41759d34, 32'h0};
test_input[3072:3079] = '{32'h424cfa84, 32'h42636cfa, 32'hc2c2e52f, 32'hc2122840, 32'h4215f95f, 32'hc2af1a79, 32'hc1998ebe, 32'hc2598093};
test_output[3072:3079] = '{32'h424cfa84, 32'h42636cfa, 32'h0, 32'h0, 32'h4215f95f, 32'h0, 32'h0, 32'h0};
test_input[3080:3087] = '{32'h412e23fa, 32'hc0ef0c92, 32'h4268ab38, 32'hc0846831, 32'h4106008b, 32'hc1aea6d4, 32'h4273f32c, 32'h40bee56f};
test_output[3080:3087] = '{32'h412e23fa, 32'h0, 32'h4268ab38, 32'h0, 32'h4106008b, 32'h0, 32'h4273f32c, 32'h40bee56f};
test_input[3088:3095] = '{32'h4208c305, 32'h420cd974, 32'hc1b13236, 32'hc17eab19, 32'hc20a2e3f, 32'h429b52f5, 32'h4144252c, 32'hc2242056};
test_output[3088:3095] = '{32'h4208c305, 32'h420cd974, 32'h0, 32'h0, 32'h0, 32'h429b52f5, 32'h4144252c, 32'h0};
test_input[3096:3103] = '{32'hc1152d44, 32'hc261bdd6, 32'hc1d4b1ad, 32'hc2465527, 32'hc092e9f5, 32'hc1c4e9d1, 32'h42060c3a, 32'hc2b78bdb};
test_output[3096:3103] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42060c3a, 32'h0};
test_input[3104:3111] = '{32'hc29a2895, 32'hc2ac8d29, 32'h425a3881, 32'h4225a264, 32'h427b88fa, 32'hc20a4ea0, 32'hc28fbb8a, 32'h429e5a95};
test_output[3104:3111] = '{32'h0, 32'h0, 32'h425a3881, 32'h4225a264, 32'h427b88fa, 32'h0, 32'h0, 32'h429e5a95};
test_input[3112:3119] = '{32'hc081a574, 32'hc28d3731, 32'hc21fd3fc, 32'h42448966, 32'hc2b93780, 32'hc2a4555d, 32'h42a54119, 32'hbfa1670a};
test_output[3112:3119] = '{32'h0, 32'h0, 32'h0, 32'h42448966, 32'h0, 32'h0, 32'h42a54119, 32'h0};
test_input[3120:3127] = '{32'hc2a0a40f, 32'h423693d5, 32'hc2a85763, 32'hc260801f, 32'hc210787d, 32'h42765fbe, 32'hc2312e4a, 32'hc2b32bbc};
test_output[3120:3127] = '{32'h0, 32'h423693d5, 32'h0, 32'h0, 32'h0, 32'h42765fbe, 32'h0, 32'h0};
test_input[3128:3135] = '{32'hc1b0e69d, 32'h4209c030, 32'hc2b02874, 32'hc193b56b, 32'hc22b87a4, 32'hc27315b8, 32'h4237d615, 32'hbf9c11bb};
test_output[3128:3135] = '{32'h0, 32'h4209c030, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4237d615, 32'h0};
test_input[3136:3143] = '{32'hc1a065fa, 32'hc21edd2b, 32'hc2c128cc, 32'h425c58d9, 32'h41b9a9ec, 32'h42a973d1, 32'h4297a51c, 32'hc227a317};
test_output[3136:3143] = '{32'h0, 32'h0, 32'h0, 32'h425c58d9, 32'h41b9a9ec, 32'h42a973d1, 32'h4297a51c, 32'h0};
test_input[3144:3151] = '{32'h421a6987, 32'hc1abfd52, 32'hc1c9290f, 32'h4224639a, 32'h4100dfb1, 32'h42ac86a5, 32'h426b03b8, 32'h4295b4b6};
test_output[3144:3151] = '{32'h421a6987, 32'h0, 32'h0, 32'h4224639a, 32'h4100dfb1, 32'h42ac86a5, 32'h426b03b8, 32'h4295b4b6};
test_input[3152:3159] = '{32'h41869dfe, 32'h4247f0c8, 32'hc24c1eb1, 32'h424a1f31, 32'hc27ffb04, 32'hc280ad9d, 32'h4199448a, 32'h42a1dd71};
test_output[3152:3159] = '{32'h41869dfe, 32'h4247f0c8, 32'h0, 32'h424a1f31, 32'h0, 32'h0, 32'h4199448a, 32'h42a1dd71};
test_input[3160:3167] = '{32'h41ca98f2, 32'h424497ab, 32'hc29acb63, 32'hc2b8a767, 32'h428678f4, 32'h41af4408, 32'h4085c954, 32'h426609aa};
test_output[3160:3167] = '{32'h41ca98f2, 32'h424497ab, 32'h0, 32'h0, 32'h428678f4, 32'h41af4408, 32'h4085c954, 32'h426609aa};
test_input[3168:3175] = '{32'h42bbd107, 32'hc16dedba, 32'h41d1d11c, 32'h422ef82d, 32'h4286d3ca, 32'hc29c498e, 32'h4177eb4d, 32'hc20528b9};
test_output[3168:3175] = '{32'h42bbd107, 32'h0, 32'h41d1d11c, 32'h422ef82d, 32'h4286d3ca, 32'h0, 32'h4177eb4d, 32'h0};
test_input[3176:3183] = '{32'h42aed780, 32'hc11e2abe, 32'hc1bff399, 32'h4111fa1e, 32'h4203b855, 32'hc2bf843a, 32'hc286534c, 32'h42b726c2};
test_output[3176:3183] = '{32'h42aed780, 32'h0, 32'h0, 32'h4111fa1e, 32'h4203b855, 32'h0, 32'h0, 32'h42b726c2};
test_input[3184:3191] = '{32'hc297b963, 32'hc1c2c196, 32'hc2abddf1, 32'h42002454, 32'h4154903d, 32'hc1b0a755, 32'h42aeace5, 32'hc28443a5};
test_output[3184:3191] = '{32'h0, 32'h0, 32'h0, 32'h42002454, 32'h4154903d, 32'h0, 32'h42aeace5, 32'h0};
test_input[3192:3199] = '{32'h42c5b9c7, 32'h42b42c07, 32'h409b7d65, 32'h4253f011, 32'hc2c79c8d, 32'h42c46d1d, 32'hc294e330, 32'hc095415e};
test_output[3192:3199] = '{32'h42c5b9c7, 32'h42b42c07, 32'h409b7d65, 32'h4253f011, 32'h0, 32'h42c46d1d, 32'h0, 32'h0};
test_input[3200:3207] = '{32'h428d4bb8, 32'h41ccd589, 32'hc28911c9, 32'hc07f377a, 32'hc2216c05, 32'h41fd8df0, 32'hc124ab92, 32'h42c312fa};
test_output[3200:3207] = '{32'h428d4bb8, 32'h41ccd589, 32'h0, 32'h0, 32'h0, 32'h41fd8df0, 32'h0, 32'h42c312fa};
test_input[3208:3215] = '{32'hc231d05a, 32'h41051e88, 32'hc20070e6, 32'h405b45e5, 32'hc269e669, 32'h42b427d0, 32'h4291dd46, 32'h429a3e57};
test_output[3208:3215] = '{32'h0, 32'h41051e88, 32'h0, 32'h405b45e5, 32'h0, 32'h42b427d0, 32'h4291dd46, 32'h429a3e57};
test_input[3216:3223] = '{32'hc287c1a4, 32'h42155b86, 32'h41f2efd2, 32'hc274e201, 32'hc1b10078, 32'hc24fc6ff, 32'h4073b742, 32'h422f97f4};
test_output[3216:3223] = '{32'h0, 32'h42155b86, 32'h41f2efd2, 32'h0, 32'h0, 32'h0, 32'h4073b742, 32'h422f97f4};
test_input[3224:3231] = '{32'hc282cb4f, 32'hc1c7aa0d, 32'h420b3751, 32'hc29c5d3f, 32'h428d0c6d, 32'h42277b19, 32'h4242c355, 32'hc20a31e4};
test_output[3224:3231] = '{32'h0, 32'h0, 32'h420b3751, 32'h0, 32'h428d0c6d, 32'h42277b19, 32'h4242c355, 32'h0};
test_input[3232:3239] = '{32'h421ee448, 32'hc1d16329, 32'hc26e19d5, 32'h42917654, 32'h42315c5f, 32'hc24b223f, 32'hc2450194, 32'h428ce634};
test_output[3232:3239] = '{32'h421ee448, 32'h0, 32'h0, 32'h42917654, 32'h42315c5f, 32'h0, 32'h0, 32'h428ce634};
test_input[3240:3247] = '{32'h422e481d, 32'h428c7886, 32'hc2a2e050, 32'h4229bfd0, 32'hc29d1b2f, 32'h41d8dac2, 32'h41fa302b, 32'h423b0ed6};
test_output[3240:3247] = '{32'h422e481d, 32'h428c7886, 32'h0, 32'h4229bfd0, 32'h0, 32'h41d8dac2, 32'h41fa302b, 32'h423b0ed6};
test_input[3248:3255] = '{32'hbfbe7fd7, 32'h4100a723, 32'h418677db, 32'h4285a529, 32'hc23e9ecd, 32'hc22228a6, 32'hc2969519, 32'h428de3f4};
test_output[3248:3255] = '{32'h0, 32'h4100a723, 32'h418677db, 32'h4285a529, 32'h0, 32'h0, 32'h0, 32'h428de3f4};
test_input[3256:3263] = '{32'h41de3768, 32'h422b9c83, 32'hc1c5c6d6, 32'h40391a38, 32'hc19ccb05, 32'hc2216af2, 32'h42b1378d, 32'hc29e5540};
test_output[3256:3263] = '{32'h41de3768, 32'h422b9c83, 32'h0, 32'h40391a38, 32'h0, 32'h0, 32'h42b1378d, 32'h0};
test_input[3264:3271] = '{32'hc1e3c195, 32'h4217bf2a, 32'hc201cc62, 32'hc2a816d5, 32'h4254bf57, 32'hc0c85c2e, 32'h42c08839, 32'hc27901a4};
test_output[3264:3271] = '{32'h0, 32'h4217bf2a, 32'h0, 32'h0, 32'h4254bf57, 32'h0, 32'h42c08839, 32'h0};
test_input[3272:3279] = '{32'h42767434, 32'h42a435b6, 32'hc2893e90, 32'h42b82f72, 32'h424fc316, 32'hc2094a51, 32'h40bf1422, 32'h41788ac2};
test_output[3272:3279] = '{32'h42767434, 32'h42a435b6, 32'h0, 32'h42b82f72, 32'h424fc316, 32'h0, 32'h40bf1422, 32'h41788ac2};
test_input[3280:3287] = '{32'hc226a161, 32'h42205c9f, 32'h4227150d, 32'h41c538a2, 32'hc24aaa0b, 32'h409132ca, 32'hc28a2ef8, 32'h4218db70};
test_output[3280:3287] = '{32'h0, 32'h42205c9f, 32'h4227150d, 32'h41c538a2, 32'h0, 32'h409132ca, 32'h0, 32'h4218db70};
test_input[3288:3295] = '{32'hc1bf0597, 32'hc2b611d9, 32'hc29c4f28, 32'h42a69343, 32'h41e938d0, 32'h41fe8289, 32'h421131ef, 32'h42c695ad};
test_output[3288:3295] = '{32'h0, 32'h0, 32'h0, 32'h42a69343, 32'h41e938d0, 32'h41fe8289, 32'h421131ef, 32'h42c695ad};
test_input[3296:3303] = '{32'hc1e8c546, 32'hc28399b6, 32'hc2ba8f44, 32'hc28ec3ec, 32'h42a826f9, 32'h422c117f, 32'hc1302eeb, 32'h4258bd3d};
test_output[3296:3303] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a826f9, 32'h422c117f, 32'h0, 32'h4258bd3d};
test_input[3304:3311] = '{32'hc2955ca0, 32'hc2bb0d24, 32'hc258cad0, 32'hc28c056c, 32'hc209ac8c, 32'hc0d38efe, 32'h427edf03, 32'hc20ade20};
test_output[3304:3311] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427edf03, 32'h0};
test_input[3312:3319] = '{32'h427adb3e, 32'h4245318b, 32'h423ce276, 32'h3ff268eb, 32'h42baf1d5, 32'h429f726e, 32'h425dbf80, 32'h4109867a};
test_output[3312:3319] = '{32'h427adb3e, 32'h4245318b, 32'h423ce276, 32'h3ff268eb, 32'h42baf1d5, 32'h429f726e, 32'h425dbf80, 32'h4109867a};
test_input[3320:3327] = '{32'hc19c3ff4, 32'h428b4d9d, 32'h427cbf4e, 32'h42a1d429, 32'hc2748745, 32'hc28411e7, 32'h42ac235f, 32'hc1dab201};
test_output[3320:3327] = '{32'h0, 32'h428b4d9d, 32'h427cbf4e, 32'h42a1d429, 32'h0, 32'h0, 32'h42ac235f, 32'h0};
test_input[3328:3335] = '{32'h41de6144, 32'h41a1dbee, 32'h415ef2f1, 32'h42b92a99, 32'h4265393f, 32'hc1dcf339, 32'hc26a1b3f, 32'hc248c92a};
test_output[3328:3335] = '{32'h41de6144, 32'h41a1dbee, 32'h415ef2f1, 32'h42b92a99, 32'h4265393f, 32'h0, 32'h0, 32'h0};
test_input[3336:3343] = '{32'h41dbc76e, 32'h42077363, 32'hc1b12606, 32'h41185ed2, 32'h41fef6f5, 32'h423ba4f1, 32'h42ac34a7, 32'hc1eb9f08};
test_output[3336:3343] = '{32'h41dbc76e, 32'h42077363, 32'h0, 32'h41185ed2, 32'h41fef6f5, 32'h423ba4f1, 32'h42ac34a7, 32'h0};
test_input[3344:3351] = '{32'hc236a714, 32'hc20ee065, 32'h41fbc32b, 32'hc28988db, 32'h421c6de8, 32'h424f3448, 32'h42953f14, 32'h419a5b63};
test_output[3344:3351] = '{32'h0, 32'h0, 32'h41fbc32b, 32'h0, 32'h421c6de8, 32'h424f3448, 32'h42953f14, 32'h419a5b63};
test_input[3352:3359] = '{32'hc209555c, 32'h4255ab51, 32'hc194620b, 32'hc211f7c9, 32'h42964a60, 32'hc29a981b, 32'hc29d2b64, 32'hc261f60a};
test_output[3352:3359] = '{32'h0, 32'h4255ab51, 32'h0, 32'h0, 32'h42964a60, 32'h0, 32'h0, 32'h0};
test_input[3360:3367] = '{32'h427a18e8, 32'h41f9d746, 32'h42a4eda8, 32'h40317e46, 32'hc299bf70, 32'h4250e71e, 32'hc26fa638, 32'h42056957};
test_output[3360:3367] = '{32'h427a18e8, 32'h41f9d746, 32'h42a4eda8, 32'h40317e46, 32'h0, 32'h4250e71e, 32'h0, 32'h42056957};
test_input[3368:3375] = '{32'hc29c0204, 32'hc1fe1244, 32'hc19cf3f6, 32'h42226e71, 32'h4260142d, 32'h4272f9c4, 32'h41b07cf3, 32'h42bc88ad};
test_output[3368:3375] = '{32'h0, 32'h0, 32'h0, 32'h42226e71, 32'h4260142d, 32'h4272f9c4, 32'h41b07cf3, 32'h42bc88ad};
test_input[3376:3383] = '{32'h422cd142, 32'hc23d9539, 32'h428d8b38, 32'h425f7206, 32'hc2a397a1, 32'hc2a1e889, 32'h42989609, 32'h42a50a2a};
test_output[3376:3383] = '{32'h422cd142, 32'h0, 32'h428d8b38, 32'h425f7206, 32'h0, 32'h0, 32'h42989609, 32'h42a50a2a};
test_input[3384:3391] = '{32'hc222f833, 32'hc200bf1b, 32'hc2acf52a, 32'h4096bae0, 32'h41f4f4f6, 32'h4278b2d8, 32'h42b248b4, 32'h42ba89b0};
test_output[3384:3391] = '{32'h0, 32'h0, 32'h0, 32'h4096bae0, 32'h41f4f4f6, 32'h4278b2d8, 32'h42b248b4, 32'h42ba89b0};
test_input[3392:3399] = '{32'hc2abccfb, 32'hc1e1b177, 32'hc257b327, 32'hc1ca0c55, 32'hc246063c, 32'h428fb75e, 32'hc2522796, 32'hc18bdee1};
test_output[3392:3399] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428fb75e, 32'h0, 32'h0};
test_input[3400:3407] = '{32'h42a5ac52, 32'h424677b3, 32'h423cc510, 32'hc298b4ff, 32'hc29aa802, 32'hc294a666, 32'h4240e851, 32'h429cd7c7};
test_output[3400:3407] = '{32'h42a5ac52, 32'h424677b3, 32'h423cc510, 32'h0, 32'h0, 32'h0, 32'h4240e851, 32'h429cd7c7};
test_input[3408:3415] = '{32'hc1528da4, 32'hc2281a84, 32'hc27e3a1d, 32'hc2bf46b5, 32'hc2c13e00, 32'h426327d9, 32'hc26e439c, 32'h425c2d8c};
test_output[3408:3415] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426327d9, 32'h0, 32'h425c2d8c};
test_input[3416:3423] = '{32'h42281f76, 32'h42c71ff5, 32'h3f43116a, 32'h4259444f, 32'h42770b13, 32'hc2619b2a, 32'hc290ee7e, 32'h41cf4e66};
test_output[3416:3423] = '{32'h42281f76, 32'h42c71ff5, 32'h3f43116a, 32'h4259444f, 32'h42770b13, 32'h0, 32'h0, 32'h41cf4e66};
test_input[3424:3431] = '{32'h4222d532, 32'hc2bf19a9, 32'hc00786d5, 32'hc28fa13f, 32'hc12078c7, 32'hc281a3c8, 32'h42a1e4e9, 32'hc03001e1};
test_output[3424:3431] = '{32'h4222d532, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a1e4e9, 32'h0};
test_input[3432:3439] = '{32'hc1c9cce5, 32'h42b308a0, 32'hc0fe6c0b, 32'hc0e4510d, 32'hc0c8b86a, 32'h40d37ef3, 32'hc2c6f501, 32'hc299bc4c};
test_output[3432:3439] = '{32'h0, 32'h42b308a0, 32'h0, 32'h0, 32'h0, 32'h40d37ef3, 32'h0, 32'h0};
test_input[3440:3447] = '{32'h426d5760, 32'hc0da0f4f, 32'hc2a59700, 32'h42621584, 32'h42b13960, 32'hc2971c8d, 32'hc2951fc9, 32'hc21b319a};
test_output[3440:3447] = '{32'h426d5760, 32'h0, 32'h0, 32'h42621584, 32'h42b13960, 32'h0, 32'h0, 32'h0};
test_input[3448:3455] = '{32'hc217044e, 32'h41ccc896, 32'hc29bb461, 32'h429b667e, 32'h413a6d57, 32'h42ae6070, 32'h40262276, 32'h429ff438};
test_output[3448:3455] = '{32'h0, 32'h41ccc896, 32'h0, 32'h429b667e, 32'h413a6d57, 32'h42ae6070, 32'h40262276, 32'h429ff438};
test_input[3456:3463] = '{32'h429bdadd, 32'h40cc9b63, 32'hc2c42f14, 32'hc2a77c62, 32'h423a8218, 32'h42abbb55, 32'h419017cf, 32'hc0aa6aa5};
test_output[3456:3463] = '{32'h429bdadd, 32'h40cc9b63, 32'h0, 32'h0, 32'h423a8218, 32'h42abbb55, 32'h419017cf, 32'h0};
test_input[3464:3471] = '{32'h42b14552, 32'hc1416ab4, 32'h4222837c, 32'hc253ab0a, 32'h41b1641d, 32'h429c8076, 32'h428c0bbc, 32'h428e5645};
test_output[3464:3471] = '{32'h42b14552, 32'h0, 32'h4222837c, 32'h0, 32'h41b1641d, 32'h429c8076, 32'h428c0bbc, 32'h428e5645};
test_input[3472:3479] = '{32'hc0a4b6e4, 32'h42a4f691, 32'h41277590, 32'h42029207, 32'hc21084cc, 32'h3dcfcd01, 32'hc2934d0c, 32'hc150a45b};
test_output[3472:3479] = '{32'h0, 32'h42a4f691, 32'h41277590, 32'h42029207, 32'h0, 32'h3dcfcd01, 32'h0, 32'h0};
test_input[3480:3487] = '{32'hc223d54f, 32'h42b588af, 32'hc285c54c, 32'h418070e1, 32'h4191dd53, 32'h42896b21, 32'h42c22ae5, 32'h42691881};
test_output[3480:3487] = '{32'h0, 32'h42b588af, 32'h0, 32'h418070e1, 32'h4191dd53, 32'h42896b21, 32'h42c22ae5, 32'h42691881};
test_input[3488:3495] = '{32'h4294c05a, 32'hc2b6b03a, 32'h42a135d8, 32'h421b0da8, 32'hc2c59bb0, 32'h4218ce02, 32'hc16a2689, 32'hc180762c};
test_output[3488:3495] = '{32'h4294c05a, 32'h0, 32'h42a135d8, 32'h421b0da8, 32'h0, 32'h4218ce02, 32'h0, 32'h0};
test_input[3496:3503] = '{32'h421d74b2, 32'hc27e0126, 32'h42a407a7, 32'hc242597f, 32'hc256d075, 32'hbff416d0, 32'h4110c93a, 32'h41cb3585};
test_output[3496:3503] = '{32'h421d74b2, 32'h0, 32'h42a407a7, 32'h0, 32'h0, 32'h0, 32'h4110c93a, 32'h41cb3585};
test_input[3504:3511] = '{32'hc24c8983, 32'h41e5a1cc, 32'hc1cd9a2b, 32'h42566e9c, 32'hc13490ea, 32'h42b08ae8, 32'h41ce7f34, 32'hc190d039};
test_output[3504:3511] = '{32'h0, 32'h41e5a1cc, 32'h0, 32'h42566e9c, 32'h0, 32'h42b08ae8, 32'h41ce7f34, 32'h0};
test_input[3512:3519] = '{32'hc2544b78, 32'h421aec5b, 32'h419c3ac6, 32'h40c21311, 32'h42c3ab31, 32'h4162e638, 32'h424d456e, 32'hc29dbe51};
test_output[3512:3519] = '{32'h0, 32'h421aec5b, 32'h419c3ac6, 32'h40c21311, 32'h42c3ab31, 32'h4162e638, 32'h424d456e, 32'h0};
test_input[3520:3527] = '{32'hc2016757, 32'h41d49845, 32'h41df7833, 32'h420805bc, 32'h413876cf, 32'hc21c5c35, 32'h429e00dd, 32'hc186691b};
test_output[3520:3527] = '{32'h0, 32'h41d49845, 32'h41df7833, 32'h420805bc, 32'h413876cf, 32'h0, 32'h429e00dd, 32'h0};
test_input[3528:3535] = '{32'hc29db028, 32'hc2113c1a, 32'h428837b7, 32'h42a31c02, 32'h4280386d, 32'h41591554, 32'h4243c8c1, 32'h418d732a};
test_output[3528:3535] = '{32'h0, 32'h0, 32'h428837b7, 32'h42a31c02, 32'h4280386d, 32'h41591554, 32'h4243c8c1, 32'h418d732a};
test_input[3536:3543] = '{32'hc2c14ed4, 32'hc1e434b6, 32'h4218af61, 32'hc1d6fc27, 32'h3fbf08bb, 32'hc25dba70, 32'h4182f6cb, 32'hc1c1e2ba};
test_output[3536:3543] = '{32'h0, 32'h0, 32'h4218af61, 32'h0, 32'h3fbf08bb, 32'h0, 32'h4182f6cb, 32'h0};
test_input[3544:3551] = '{32'hc22c7e08, 32'h422fb706, 32'hc2aa3fc3, 32'h4285ca1c, 32'hbfccd5ff, 32'h41bfd608, 32'hc18ee8c7, 32'h41e73957};
test_output[3544:3551] = '{32'h0, 32'h422fb706, 32'h0, 32'h4285ca1c, 32'h0, 32'h41bfd608, 32'h0, 32'h41e73957};
test_input[3552:3559] = '{32'hc2a17344, 32'h42651b9a, 32'hc2004300, 32'hc282d265, 32'h40cf89f3, 32'h4200ef53, 32'h413c4b03, 32'h40e51e87};
test_output[3552:3559] = '{32'h0, 32'h42651b9a, 32'h0, 32'h0, 32'h40cf89f3, 32'h4200ef53, 32'h413c4b03, 32'h40e51e87};
test_input[3560:3567] = '{32'hc29f8e9f, 32'hc27d034e, 32'hc2643c54, 32'h4173c41b, 32'hc15156bc, 32'h42402fd2, 32'h426e2955, 32'h421db5aa};
test_output[3560:3567] = '{32'h0, 32'h0, 32'h0, 32'h4173c41b, 32'h0, 32'h42402fd2, 32'h426e2955, 32'h421db5aa};
test_input[3568:3575] = '{32'h3fc1f73b, 32'hc2ba417a, 32'hc297c189, 32'h41f931d0, 32'hc1954e4c, 32'hc2c58c72, 32'hc2bf9ff2, 32'hc1aa86af};
test_output[3568:3575] = '{32'h3fc1f73b, 32'h0, 32'h0, 32'h41f931d0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3576:3583] = '{32'hc267c4d8, 32'h41f1b324, 32'h4187c397, 32'hc21d562d, 32'h42632754, 32'h422c0366, 32'h41df3e89, 32'hc1ab63ba};
test_output[3576:3583] = '{32'h0, 32'h41f1b324, 32'h4187c397, 32'h0, 32'h42632754, 32'h422c0366, 32'h41df3e89, 32'h0};
test_input[3584:3591] = '{32'h4297223c, 32'hc23e75df, 32'hc29a8458, 32'h42bbc85e, 32'hc27bc2cf, 32'h429e1988, 32'hc2a5148f, 32'hc206e900};
test_output[3584:3591] = '{32'h4297223c, 32'h0, 32'h0, 32'h42bbc85e, 32'h0, 32'h429e1988, 32'h0, 32'h0};
test_input[3592:3599] = '{32'h407dabc8, 32'h419db049, 32'h41b72053, 32'h41194489, 32'hc2707e76, 32'h413ee42a, 32'hc26feb6a, 32'hc2371306};
test_output[3592:3599] = '{32'h407dabc8, 32'h419db049, 32'h41b72053, 32'h41194489, 32'h0, 32'h413ee42a, 32'h0, 32'h0};
test_input[3600:3607] = '{32'hc2b61f0a, 32'h42a76b43, 32'hc2bc07cc, 32'h429fc08e, 32'h42794dcb, 32'hc28ec9fa, 32'h42054a3a, 32'h42ba24b2};
test_output[3600:3607] = '{32'h0, 32'h42a76b43, 32'h0, 32'h429fc08e, 32'h42794dcb, 32'h0, 32'h42054a3a, 32'h42ba24b2};
test_input[3608:3615] = '{32'h42842801, 32'hc0571357, 32'h42ad6b79, 32'h40718ca4, 32'hc293af89, 32'h41ce2d98, 32'h4290dedd, 32'h42742f53};
test_output[3608:3615] = '{32'h42842801, 32'h0, 32'h42ad6b79, 32'h40718ca4, 32'h0, 32'h41ce2d98, 32'h4290dedd, 32'h42742f53};
test_input[3616:3623] = '{32'hc2c58ace, 32'h42886376, 32'h4214df48, 32'h427daa7e, 32'hc2a1f174, 32'hc2482237, 32'hc22e9ecc, 32'hc2242cc8};
test_output[3616:3623] = '{32'h0, 32'h42886376, 32'h4214df48, 32'h427daa7e, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3624:3631] = '{32'h422ef8e7, 32'h424229fc, 32'h41f06310, 32'hc10f935d, 32'hc16ff248, 32'h4263b688, 32'hc077aa28, 32'hc2bbe51c};
test_output[3624:3631] = '{32'h422ef8e7, 32'h424229fc, 32'h41f06310, 32'h0, 32'h0, 32'h4263b688, 32'h0, 32'h0};
test_input[3632:3639] = '{32'h4297a4fa, 32'hc2a7b13c, 32'h42c707ac, 32'hc27291a5, 32'hc19e3111, 32'hc11885de, 32'hc165cf53, 32'hc230a05b};
test_output[3632:3639] = '{32'h4297a4fa, 32'h0, 32'h42c707ac, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3640:3647] = '{32'hc1b62d7f, 32'h41eadbd0, 32'hc24d843c, 32'hc16bb5e3, 32'hc2880bb7, 32'h423927b1, 32'h4248bbce, 32'hc2b956b0};
test_output[3640:3647] = '{32'h0, 32'h41eadbd0, 32'h0, 32'h0, 32'h0, 32'h423927b1, 32'h4248bbce, 32'h0};
test_input[3648:3655] = '{32'h42b78f50, 32'h42b94c1d, 32'hc2882dfa, 32'h41d21bed, 32'h424ec123, 32'hbf96a85b, 32'hc18fd8dd, 32'hc1c279a5};
test_output[3648:3655] = '{32'h42b78f50, 32'h42b94c1d, 32'h0, 32'h41d21bed, 32'h424ec123, 32'h0, 32'h0, 32'h0};
test_input[3656:3663] = '{32'h426d7f34, 32'h41b71c63, 32'h4195a1e0, 32'hc2c227a2, 32'hc2bdde5c, 32'hc237a1b3, 32'h42574cfe, 32'hc1aba620};
test_output[3656:3663] = '{32'h426d7f34, 32'h41b71c63, 32'h4195a1e0, 32'h0, 32'h0, 32'h0, 32'h42574cfe, 32'h0};
test_input[3664:3671] = '{32'h41cc247f, 32'h421d79ce, 32'h42232c43, 32'hc2bbbcac, 32'hc2b9165f, 32'h422fe374, 32'hc0a0dffa, 32'hc16f45e4};
test_output[3664:3671] = '{32'h41cc247f, 32'h421d79ce, 32'h42232c43, 32'h0, 32'h0, 32'h422fe374, 32'h0, 32'h0};
test_input[3672:3679] = '{32'h41f000a6, 32'hc220b9fd, 32'hc273fe23, 32'hc2c43d02, 32'hc2bdb41c, 32'h41ff56f9, 32'hc225a8b6, 32'h42014c36};
test_output[3672:3679] = '{32'h41f000a6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ff56f9, 32'h0, 32'h42014c36};
test_input[3680:3687] = '{32'hc2953693, 32'hc2140f20, 32'h417019cd, 32'hc1c72faa, 32'hc2a059ac, 32'hc1db30ee, 32'h421993a0, 32'hc288775d};
test_output[3680:3687] = '{32'h0, 32'h0, 32'h417019cd, 32'h0, 32'h0, 32'h0, 32'h421993a0, 32'h0};
test_input[3688:3695] = '{32'h428d3397, 32'hc2bc352b, 32'hc2b88d51, 32'hc244f8d2, 32'hc0585509, 32'hc29a5d4a, 32'h42c0705d, 32'h4285b7c8};
test_output[3688:3695] = '{32'h428d3397, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c0705d, 32'h4285b7c8};
test_input[3696:3703] = '{32'hc1ca8369, 32'hc27a6139, 32'hc223ca8d, 32'h42a78865, 32'hbf80d5ff, 32'hc2c600d6, 32'h42961010, 32'hc28b0df2};
test_output[3696:3703] = '{32'h0, 32'h0, 32'h0, 32'h42a78865, 32'h0, 32'h0, 32'h42961010, 32'h0};
test_input[3704:3711] = '{32'hc2962ad3, 32'hc2be224e, 32'h42c4166b, 32'h41f5a3ac, 32'hc2bc5ce2, 32'h41d1dfe2, 32'h424e610d, 32'hc211a0df};
test_output[3704:3711] = '{32'h0, 32'h0, 32'h42c4166b, 32'h41f5a3ac, 32'h0, 32'h41d1dfe2, 32'h424e610d, 32'h0};
test_input[3712:3719] = '{32'hc2a00a31, 32'hc24891f3, 32'hc2825f4f, 32'h42bbd38c, 32'hc24a358f, 32'h411b96d4, 32'hc2723266, 32'hc2a21b32};
test_output[3712:3719] = '{32'h0, 32'h0, 32'h0, 32'h42bbd38c, 32'h0, 32'h411b96d4, 32'h0, 32'h0};
test_input[3720:3727] = '{32'hc14aa3a4, 32'hc1c12076, 32'h42234aed, 32'h4195cc56, 32'h428ec8ea, 32'h41b3d1be, 32'h3f6254a7, 32'h41cc8a23};
test_output[3720:3727] = '{32'h0, 32'h0, 32'h42234aed, 32'h4195cc56, 32'h428ec8ea, 32'h41b3d1be, 32'h3f6254a7, 32'h41cc8a23};
test_input[3728:3735] = '{32'h4255f5aa, 32'hc24aea60, 32'hc2b217db, 32'h429a38f3, 32'hc2858055, 32'hc23f2b21, 32'hc1a0968e, 32'hc2429cff};
test_output[3728:3735] = '{32'h4255f5aa, 32'h0, 32'h0, 32'h429a38f3, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3736:3743] = '{32'hc28953c0, 32'h3e569009, 32'h41bdf7d4, 32'hc2ad3be3, 32'h426178c1, 32'h414e3969, 32'h418a4315, 32'h42a33793};
test_output[3736:3743] = '{32'h0, 32'h3e569009, 32'h41bdf7d4, 32'h0, 32'h426178c1, 32'h414e3969, 32'h418a4315, 32'h42a33793};
test_input[3744:3751] = '{32'hc1acd78b, 32'h42ad373a, 32'hc23d5694, 32'h4231bea0, 32'hc218c8c6, 32'h414a532a, 32'hc0464fdf, 32'hc2292674};
test_output[3744:3751] = '{32'h0, 32'h42ad373a, 32'h0, 32'h4231bea0, 32'h0, 32'h414a532a, 32'h0, 32'h0};
test_input[3752:3759] = '{32'h41a6c9e2, 32'h429ad02b, 32'hc22645cc, 32'h410daa6c, 32'h4224ce62, 32'h41f9edf4, 32'h429d1165, 32'h41228c1a};
test_output[3752:3759] = '{32'h41a6c9e2, 32'h429ad02b, 32'h0, 32'h410daa6c, 32'h4224ce62, 32'h41f9edf4, 32'h429d1165, 32'h41228c1a};
test_input[3760:3767] = '{32'hc28db224, 32'hc2922b9f, 32'h419585c4, 32'hc1fa7641, 32'h421ef765, 32'h4219f54e, 32'hc2057f0f, 32'hc2b2ac08};
test_output[3760:3767] = '{32'h0, 32'h0, 32'h419585c4, 32'h0, 32'h421ef765, 32'h4219f54e, 32'h0, 32'h0};
test_input[3768:3775] = '{32'h417d3ba7, 32'h42b3cb63, 32'h41954c19, 32'h42b2720f, 32'hc216fb57, 32'h42202801, 32'h41d31977, 32'hc2541c52};
test_output[3768:3775] = '{32'h417d3ba7, 32'h42b3cb63, 32'h41954c19, 32'h42b2720f, 32'h0, 32'h42202801, 32'h41d31977, 32'h0};
test_input[3776:3783] = '{32'h42c26c05, 32'h4281287b, 32'h427d5f7a, 32'hc23f01ba, 32'hc28ff467, 32'hc2411dda, 32'h4218bd42, 32'hc11a0ca1};
test_output[3776:3783] = '{32'h42c26c05, 32'h4281287b, 32'h427d5f7a, 32'h0, 32'h0, 32'h0, 32'h4218bd42, 32'h0};
test_input[3784:3791] = '{32'hc1cb7133, 32'hc272deb0, 32'hbf9d1851, 32'h428f67f2, 32'hc0ea7ebe, 32'hc28179a9, 32'h42a3728e, 32'hc256a439};
test_output[3784:3791] = '{32'h0, 32'h0, 32'h0, 32'h428f67f2, 32'h0, 32'h0, 32'h42a3728e, 32'h0};
test_input[3792:3799] = '{32'hc247699e, 32'h42954a31, 32'hc147ea9e, 32'hc285b1d4, 32'h42931d1c, 32'hc26fd98e, 32'h41b1613e, 32'hc22a4845};
test_output[3792:3799] = '{32'h0, 32'h42954a31, 32'h0, 32'h0, 32'h42931d1c, 32'h0, 32'h41b1613e, 32'h0};
test_input[3800:3807] = '{32'h4176ec09, 32'h42c795af, 32'hc2864a49, 32'h4236c1d2, 32'hc27289d2, 32'h4292760c, 32'hc26f5c72, 32'hc279db54};
test_output[3800:3807] = '{32'h4176ec09, 32'h42c795af, 32'h0, 32'h4236c1d2, 32'h0, 32'h4292760c, 32'h0, 32'h0};
test_input[3808:3815] = '{32'h426a8ea4, 32'h41c1f28c, 32'h42091863, 32'h42ab219a, 32'hc2450d86, 32'hc288e7fa, 32'hc255da13, 32'h4274e8f7};
test_output[3808:3815] = '{32'h426a8ea4, 32'h41c1f28c, 32'h42091863, 32'h42ab219a, 32'h0, 32'h0, 32'h0, 32'h4274e8f7};
test_input[3816:3823] = '{32'h42bcf5db, 32'h42343f18, 32'hc183be2f, 32'hc2b5f414, 32'h42b2d721, 32'h424be821, 32'h4145cb97, 32'h42c3ff5f};
test_output[3816:3823] = '{32'h42bcf5db, 32'h42343f18, 32'h0, 32'h0, 32'h42b2d721, 32'h424be821, 32'h4145cb97, 32'h42c3ff5f};
test_input[3824:3831] = '{32'hc275833a, 32'hc2ac66cf, 32'h4269a996, 32'hc25de479, 32'hc1fd1588, 32'hc28ce018, 32'h42556948, 32'hc2bb108d};
test_output[3824:3831] = '{32'h0, 32'h0, 32'h4269a996, 32'h0, 32'h0, 32'h0, 32'h42556948, 32'h0};
test_input[3832:3839] = '{32'h4070a207, 32'h421f42a7, 32'h41f26a5a, 32'hc2069af9, 32'hc26518c5, 32'h41af9f8a, 32'hc253bc9c, 32'h42425e73};
test_output[3832:3839] = '{32'h4070a207, 32'h421f42a7, 32'h41f26a5a, 32'h0, 32'h0, 32'h41af9f8a, 32'h0, 32'h42425e73};
test_input[3840:3847] = '{32'h415ff117, 32'hc20b7d27, 32'hc2966eb3, 32'h42b5ab8f, 32'hc2244b93, 32'h41e71b57, 32'h426dfa8e, 32'hc22e196e};
test_output[3840:3847] = '{32'h415ff117, 32'h0, 32'h0, 32'h42b5ab8f, 32'h0, 32'h41e71b57, 32'h426dfa8e, 32'h0};
test_input[3848:3855] = '{32'hc2888104, 32'h4293bb43, 32'hc251c915, 32'h42938c3d, 32'h426e22fd, 32'hc031c5f8, 32'h42c0eedc, 32'h4259bbf7};
test_output[3848:3855] = '{32'h0, 32'h4293bb43, 32'h0, 32'h42938c3d, 32'h426e22fd, 32'h0, 32'h42c0eedc, 32'h4259bbf7};
test_input[3856:3863] = '{32'h424a627d, 32'hc26dde48, 32'h42197790, 32'h412beee3, 32'h4250e6d2, 32'h4295a7df, 32'hc0618d8f, 32'hc2aa16ba};
test_output[3856:3863] = '{32'h424a627d, 32'h0, 32'h42197790, 32'h412beee3, 32'h4250e6d2, 32'h4295a7df, 32'h0, 32'h0};
test_input[3864:3871] = '{32'hc21f1df7, 32'h414194a3, 32'hc1faac69, 32'h423d1e39, 32'hc2b31a10, 32'hc265729c, 32'hc1b46e37, 32'h4195636f};
test_output[3864:3871] = '{32'h0, 32'h414194a3, 32'h0, 32'h423d1e39, 32'h0, 32'h0, 32'h0, 32'h4195636f};
test_input[3872:3879] = '{32'h42b77433, 32'hc1e26d46, 32'hc2309936, 32'hc11fdeeb, 32'hc254cb7d, 32'hc200cf39, 32'h42a8a512, 32'h429aa6eb};
test_output[3872:3879] = '{32'h42b77433, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a8a512, 32'h429aa6eb};
test_input[3880:3887] = '{32'hc251b1ae, 32'hc286f3e6, 32'h424817a8, 32'hc2591f0e, 32'h41c2055c, 32'hc0e06e88, 32'hc117aebf, 32'h429f8ee1};
test_output[3880:3887] = '{32'h0, 32'h0, 32'h424817a8, 32'h0, 32'h41c2055c, 32'h0, 32'h0, 32'h429f8ee1};
test_input[3888:3895] = '{32'h42563a4c, 32'hc1a642bf, 32'h427d239b, 32'hc2a88612, 32'hc0d5bbde, 32'hc0579820, 32'h4182c358, 32'h429063b9};
test_output[3888:3895] = '{32'h42563a4c, 32'h0, 32'h427d239b, 32'h0, 32'h0, 32'h0, 32'h4182c358, 32'h429063b9};
test_input[3896:3903] = '{32'hc172b9be, 32'h41951b3a, 32'h41f1fa1d, 32'h42396708, 32'h4271551a, 32'h425f729d, 32'h42abdd7d, 32'hc24cefe4};
test_output[3896:3903] = '{32'h0, 32'h41951b3a, 32'h41f1fa1d, 32'h42396708, 32'h4271551a, 32'h425f729d, 32'h42abdd7d, 32'h0};
test_input[3904:3911] = '{32'h4259eca0, 32'h42c2c1e1, 32'hc29b3876, 32'hc1455ea7, 32'hc1a5b1c1, 32'h4294585b, 32'h4295af1f, 32'hc277936e};
test_output[3904:3911] = '{32'h4259eca0, 32'h42c2c1e1, 32'h0, 32'h0, 32'h0, 32'h4294585b, 32'h4295af1f, 32'h0};
test_input[3912:3919] = '{32'hc18f90ce, 32'hc22945d4, 32'h424f6c39, 32'hc2b3336b, 32'h4287d836, 32'h424e48bd, 32'hc112a3cc, 32'hc09de112};
test_output[3912:3919] = '{32'h0, 32'h0, 32'h424f6c39, 32'h0, 32'h4287d836, 32'h424e48bd, 32'h0, 32'h0};
test_input[3920:3927] = '{32'hc12fc79e, 32'hc21cdb37, 32'h428fe60f, 32'hc1d14fa5, 32'h42a0000e, 32'h429418bf, 32'hc11a1a0e, 32'hc297dd33};
test_output[3920:3927] = '{32'h0, 32'h0, 32'h428fe60f, 32'h0, 32'h42a0000e, 32'h429418bf, 32'h0, 32'h0};
test_input[3928:3935] = '{32'h42b32164, 32'h41b877f6, 32'h4138a926, 32'hc1ed46e2, 32'hc247fe22, 32'h40e3052e, 32'h42bdfeae, 32'h42935796};
test_output[3928:3935] = '{32'h42b32164, 32'h41b877f6, 32'h4138a926, 32'h0, 32'h0, 32'h40e3052e, 32'h42bdfeae, 32'h42935796};
test_input[3936:3943] = '{32'h42af0ae1, 32'hc268da6c, 32'hc28fd990, 32'h425206dd, 32'hbf9e24a3, 32'hc2a28c33, 32'hc2b57c37, 32'hc23d0961};
test_output[3936:3943] = '{32'h42af0ae1, 32'h0, 32'h0, 32'h425206dd, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[3944:3951] = '{32'h41332621, 32'h42b27275, 32'hc2a9ad68, 32'hc29b862d, 32'hc2a2fd02, 32'h42767e48, 32'hc1ea5f9e, 32'hc2850d94};
test_output[3944:3951] = '{32'h41332621, 32'h42b27275, 32'h0, 32'h0, 32'h0, 32'h42767e48, 32'h0, 32'h0};
test_input[3952:3959] = '{32'h42b1da34, 32'hc2a26400, 32'h42531bc1, 32'h4204e754, 32'hc28bced3, 32'hc2a7b22c, 32'hc1caadab, 32'h4283e048};
test_output[3952:3959] = '{32'h42b1da34, 32'h0, 32'h42531bc1, 32'h4204e754, 32'h0, 32'h0, 32'h0, 32'h4283e048};
test_input[3960:3967] = '{32'h4200bb06, 32'hc2bc1d18, 32'h423f7a10, 32'h42988018, 32'h4279b7b2, 32'h42ae5e6d, 32'h42581600, 32'hc0a52d8e};
test_output[3960:3967] = '{32'h4200bb06, 32'h0, 32'h423f7a10, 32'h42988018, 32'h4279b7b2, 32'h42ae5e6d, 32'h42581600, 32'h0};
test_input[3968:3975] = '{32'h42a57959, 32'hc1756e70, 32'hc2afc14a, 32'hc00beaf0, 32'h42907466, 32'h42247aab, 32'h42bad1d2, 32'hc28610eb};
test_output[3968:3975] = '{32'h42a57959, 32'h0, 32'h0, 32'h0, 32'h42907466, 32'h42247aab, 32'h42bad1d2, 32'h0};
test_input[3976:3983] = '{32'hc26be9b0, 32'hc28249fa, 32'hc29b7ec0, 32'hc2acd756, 32'h4234a264, 32'hc2afe16b, 32'h423821d2, 32'h42198393};
test_output[3976:3983] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4234a264, 32'h0, 32'h423821d2, 32'h42198393};
test_input[3984:3991] = '{32'h42aec205, 32'h42c5b79a, 32'h41b2730b, 32'hc2a9c894, 32'hc2ad45f8, 32'hc278e936, 32'hc29e638a, 32'h42c0743b};
test_output[3984:3991] = '{32'h42aec205, 32'h42c5b79a, 32'h41b2730b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c0743b};
test_input[3992:3999] = '{32'h42370b7d, 32'h40852a81, 32'h42137bcb, 32'hc15e99a6, 32'h429b98cc, 32'hc2850dca, 32'h4241b451, 32'hc15835bd};
test_output[3992:3999] = '{32'h42370b7d, 32'h40852a81, 32'h42137bcb, 32'h0, 32'h429b98cc, 32'h0, 32'h4241b451, 32'h0};
test_input[4000:4007] = '{32'h40e313d4, 32'hc29b1b9c, 32'h42b29784, 32'h41b93504, 32'h41177cc9, 32'h410c0c5a, 32'hc07e1cc7, 32'h425fa8da};
test_output[4000:4007] = '{32'h40e313d4, 32'h0, 32'h42b29784, 32'h41b93504, 32'h41177cc9, 32'h410c0c5a, 32'h0, 32'h425fa8da};
test_input[4008:4015] = '{32'hc268d108, 32'hc29273e4, 32'hc200df37, 32'hc234ff26, 32'hc2b3b49b, 32'h429f3d3a, 32'hc1fabace, 32'hc293777b};
test_output[4008:4015] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429f3d3a, 32'h0, 32'h0};
test_input[4016:4023] = '{32'hc27cadfb, 32'hc2a28907, 32'h42b68238, 32'h42783bf6, 32'hc2af1939, 32'hc281af3c, 32'hc0ccff64, 32'h42afad0a};
test_output[4016:4023] = '{32'h0, 32'h0, 32'h42b68238, 32'h42783bf6, 32'h0, 32'h0, 32'h0, 32'h42afad0a};
test_input[4024:4031] = '{32'h41b21369, 32'h42370d5f, 32'hc226bb9d, 32'hc147566c, 32'h428b5440, 32'hc2913ebe, 32'h42244c99, 32'h41a5a535};
test_output[4024:4031] = '{32'h41b21369, 32'h42370d5f, 32'h0, 32'h0, 32'h428b5440, 32'h0, 32'h42244c99, 32'h41a5a535};
test_input[4032:4039] = '{32'hc2afad87, 32'h421422eb, 32'h424a085f, 32'hc2450e0d, 32'hc29f2d93, 32'hc100506f, 32'hc0476ee7, 32'h42ad0b83};
test_output[4032:4039] = '{32'h0, 32'h421422eb, 32'h424a085f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ad0b83};
test_input[4040:4047] = '{32'h425432e9, 32'h420c0cb1, 32'h3fd4e62a, 32'hc2b69c02, 32'hc23089f8, 32'hc1ee7953, 32'hc2989bcb, 32'h42a0f6fd};
test_output[4040:4047] = '{32'h425432e9, 32'h420c0cb1, 32'h3fd4e62a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a0f6fd};
test_input[4048:4055] = '{32'h41c835b5, 32'hc20d0db9, 32'hc26114a3, 32'h42b49c5a, 32'hc250ce90, 32'hc22d255d, 32'h427580a7, 32'hc0ea0a10};
test_output[4048:4055] = '{32'h41c835b5, 32'h0, 32'h0, 32'h42b49c5a, 32'h0, 32'h0, 32'h427580a7, 32'h0};
test_input[4056:4063] = '{32'h40b38a2f, 32'h42c0c7f9, 32'h4213e4a4, 32'hc2001367, 32'hc2b52f6a, 32'h426b0582, 32'hc2bef386, 32'h4242b833};
test_output[4056:4063] = '{32'h40b38a2f, 32'h42c0c7f9, 32'h4213e4a4, 32'h0, 32'h0, 32'h426b0582, 32'h0, 32'h4242b833};
test_input[4064:4071] = '{32'h41c5f04a, 32'h4215f209, 32'hc2012a98, 32'hc0c86001, 32'h424bdc6f, 32'hc2897736, 32'h4278579a, 32'h41b4a662};
test_output[4064:4071] = '{32'h41c5f04a, 32'h4215f209, 32'h0, 32'h0, 32'h424bdc6f, 32'h0, 32'h4278579a, 32'h41b4a662};
test_input[4072:4079] = '{32'hc2b99c0b, 32'hc174afb1, 32'h41fa8341, 32'hc2a04837, 32'hc01eddbf, 32'hc2b2ef28, 32'hc050a496, 32'h42874bed};
test_output[4072:4079] = '{32'h0, 32'h0, 32'h41fa8341, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42874bed};
test_input[4080:4087] = '{32'hc2aab316, 32'hc2b651d1, 32'h427baacd, 32'h4077ed3f, 32'hc2776c37, 32'hc23570a0, 32'h4270107d, 32'hc2822004};
test_output[4080:4087] = '{32'h0, 32'h0, 32'h427baacd, 32'h4077ed3f, 32'h0, 32'h0, 32'h4270107d, 32'h0};
test_input[4088:4095] = '{32'h4215890a, 32'hc23b305a, 32'h41d517de, 32'hc2523922, 32'hc286ade3, 32'h427457c7, 32'h41e27d46, 32'hc2b75fc4};
test_output[4088:4095] = '{32'h4215890a, 32'h0, 32'h41d517de, 32'h0, 32'h0, 32'h427457c7, 32'h41e27d46, 32'h0};
test_input[4096:4103] = '{32'hc2b7da01, 32'hbf0956d9, 32'hc1d13efa, 32'hc284e8b1, 32'h41f2b16a, 32'h41c575d2, 32'hc113f185, 32'h42354c06};
test_output[4096:4103] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41f2b16a, 32'h41c575d2, 32'h0, 32'h42354c06};
test_input[4104:4111] = '{32'hc285c5e6, 32'hc2c73168, 32'hc2980d26, 32'h42b9aec9, 32'h42271022, 32'hc28d9bb4, 32'h41efab24, 32'hc28d4b26};
test_output[4104:4111] = '{32'h0, 32'h0, 32'h0, 32'h42b9aec9, 32'h42271022, 32'h0, 32'h41efab24, 32'h0};
test_input[4112:4119] = '{32'h42bbd704, 32'hc2b4e951, 32'h416903cd, 32'h42114e6e, 32'hc1459792, 32'hc106d71a, 32'h420cac43, 32'hc1884202};
test_output[4112:4119] = '{32'h42bbd704, 32'h0, 32'h416903cd, 32'h42114e6e, 32'h0, 32'h0, 32'h420cac43, 32'h0};
test_input[4120:4127] = '{32'hc2a349dc, 32'hc2611105, 32'h40a57283, 32'hc2c6872a, 32'hc26b6241, 32'h401c0a9b, 32'hc21e9327, 32'h42898688};
test_output[4120:4127] = '{32'h0, 32'h0, 32'h40a57283, 32'h0, 32'h0, 32'h401c0a9b, 32'h0, 32'h42898688};
test_input[4128:4135] = '{32'hc2c32a07, 32'hc2199534, 32'h420b788c, 32'h426b71b0, 32'h420a3b40, 32'hc29999a6, 32'h41fe8ee4, 32'h428a11fc};
test_output[4128:4135] = '{32'h0, 32'h0, 32'h420b788c, 32'h426b71b0, 32'h420a3b40, 32'h0, 32'h41fe8ee4, 32'h428a11fc};
test_input[4136:4143] = '{32'h42981a04, 32'h424aac45, 32'hc29b5642, 32'h422b9cb5, 32'hc22d25b4, 32'hc1dcb0d9, 32'h42a99c51, 32'hc281d142};
test_output[4136:4143] = '{32'h42981a04, 32'h424aac45, 32'h0, 32'h422b9cb5, 32'h0, 32'h0, 32'h42a99c51, 32'h0};
test_input[4144:4151] = '{32'hc0d4db80, 32'h41085f14, 32'h418b1894, 32'hc22b6809, 32'h427dc687, 32'hc1a1fd1c, 32'hc2300fea, 32'h41e90fb5};
test_output[4144:4151] = '{32'h0, 32'h41085f14, 32'h418b1894, 32'h0, 32'h427dc687, 32'h0, 32'h0, 32'h41e90fb5};
test_input[4152:4159] = '{32'h424357c1, 32'h4193c841, 32'hc1d7a015, 32'h41ec4060, 32'h405fdaff, 32'h425c15dd, 32'h4190845c, 32'hc234acdf};
test_output[4152:4159] = '{32'h424357c1, 32'h4193c841, 32'h0, 32'h41ec4060, 32'h405fdaff, 32'h425c15dd, 32'h4190845c, 32'h0};
test_input[4160:4167] = '{32'h42241042, 32'hc25db353, 32'hc28e42e4, 32'hc1268fc8, 32'h42b71865, 32'hc1f64dbf, 32'hc2c402e5, 32'h42256eed};
test_output[4160:4167] = '{32'h42241042, 32'h0, 32'h0, 32'h0, 32'h42b71865, 32'h0, 32'h0, 32'h42256eed};
test_input[4168:4175] = '{32'h423a475f, 32'h42b61bf5, 32'h4285104b, 32'hc2a24dbb, 32'hbfdae69d, 32'hc2067fba, 32'h41cf076a, 32'h421d7833};
test_output[4168:4175] = '{32'h423a475f, 32'h42b61bf5, 32'h4285104b, 32'h0, 32'h0, 32'h0, 32'h41cf076a, 32'h421d7833};
test_input[4176:4183] = '{32'hc26da4e3, 32'hc2073032, 32'hc1bbdec4, 32'hc2893fa3, 32'h41ad0166, 32'hc1f19bc8, 32'h416b33b3, 32'h42477d32};
test_output[4176:4183] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41ad0166, 32'h0, 32'h416b33b3, 32'h42477d32};
test_input[4184:4191] = '{32'h4143a8fd, 32'hc268e3c9, 32'hc2892259, 32'hc2ae132d, 32'h422a6e5e, 32'h429e00f5, 32'hc21cc78a, 32'hc2b08c6a};
test_output[4184:4191] = '{32'h4143a8fd, 32'h0, 32'h0, 32'h0, 32'h422a6e5e, 32'h429e00f5, 32'h0, 32'h0};
test_input[4192:4199] = '{32'h4266ae66, 32'h42bc99b6, 32'hc06250d6, 32'hc253de92, 32'h42b5eb9b, 32'h42a74370, 32'h419a1b7b, 32'hc1817a2d};
test_output[4192:4199] = '{32'h4266ae66, 32'h42bc99b6, 32'h0, 32'h0, 32'h42b5eb9b, 32'h42a74370, 32'h419a1b7b, 32'h0};
test_input[4200:4207] = '{32'hc21f5338, 32'h4282f8c5, 32'h41331b3f, 32'hc0b93e9e, 32'h42c0106a, 32'h412da933, 32'h424aff07, 32'h429ce011};
test_output[4200:4207] = '{32'h0, 32'h4282f8c5, 32'h41331b3f, 32'h0, 32'h42c0106a, 32'h412da933, 32'h424aff07, 32'h429ce011};
test_input[4208:4215] = '{32'h41f04a46, 32'hc1bbbccf, 32'h425ff4dc, 32'h425bc4ec, 32'hc19f14b3, 32'hc2a8d2e9, 32'h428e4389, 32'hc21898a5};
test_output[4208:4215] = '{32'h41f04a46, 32'h0, 32'h425ff4dc, 32'h425bc4ec, 32'h0, 32'h0, 32'h428e4389, 32'h0};
test_input[4216:4223] = '{32'h42b9bca2, 32'hc2b7ba23, 32'h4106a58a, 32'hc1fd2585, 32'h42115821, 32'h42bea497, 32'hc290b020, 32'hc27374a9};
test_output[4216:4223] = '{32'h42b9bca2, 32'h0, 32'h4106a58a, 32'h0, 32'h42115821, 32'h42bea497, 32'h0, 32'h0};
test_input[4224:4231] = '{32'hc1816982, 32'hc28fbfa7, 32'hc280abee, 32'h41c58e70, 32'hc262bf1e, 32'hc26369c6, 32'h42856fc1, 32'h41dbc7a0};
test_output[4224:4231] = '{32'h0, 32'h0, 32'h0, 32'h41c58e70, 32'h0, 32'h0, 32'h42856fc1, 32'h41dbc7a0};
test_input[4232:4239] = '{32'h3f10c5b3, 32'h4292a82c, 32'h4256b9d0, 32'hc12fd8de, 32'h41556b8a, 32'h427ee171, 32'hc1cba36e, 32'hc258e399};
test_output[4232:4239] = '{32'h3f10c5b3, 32'h4292a82c, 32'h4256b9d0, 32'h0, 32'h41556b8a, 32'h427ee171, 32'h0, 32'h0};
test_input[4240:4247] = '{32'h41e7648b, 32'h4246ff0a, 32'hc1e63efd, 32'hc2835ab1, 32'h42a56afb, 32'hc2a40df8, 32'h4283a26f, 32'hc23334f3};
test_output[4240:4247] = '{32'h41e7648b, 32'h4246ff0a, 32'h0, 32'h0, 32'h42a56afb, 32'h0, 32'h4283a26f, 32'h0};
test_input[4248:4255] = '{32'hc208f7b2, 32'h4201c651, 32'h41b981d0, 32'hc2908e5f, 32'hc2ab6ddb, 32'hc24cd928, 32'h42930954, 32'h426f45e4};
test_output[4248:4255] = '{32'h0, 32'h4201c651, 32'h41b981d0, 32'h0, 32'h0, 32'h0, 32'h42930954, 32'h426f45e4};
test_input[4256:4263] = '{32'hc2a13112, 32'hc29a001c, 32'h4190d264, 32'hc291f3b9, 32'h42ad9f67, 32'h41816d49, 32'hc2b98a24, 32'h42ac03d1};
test_output[4256:4263] = '{32'h0, 32'h0, 32'h4190d264, 32'h0, 32'h42ad9f67, 32'h41816d49, 32'h0, 32'h42ac03d1};
test_input[4264:4271] = '{32'h4294bda3, 32'h42697287, 32'hc15477b2, 32'h41cbe503, 32'h420800d0, 32'h41e8428b, 32'h426e4950, 32'h42650685};
test_output[4264:4271] = '{32'h4294bda3, 32'h42697287, 32'h0, 32'h41cbe503, 32'h420800d0, 32'h41e8428b, 32'h426e4950, 32'h42650685};
test_input[4272:4279] = '{32'h428ab04b, 32'h422b593d, 32'hc21ed4e3, 32'h42043f7c, 32'hc277395e, 32'hc225a898, 32'h42a7878f, 32'hc29e64e2};
test_output[4272:4279] = '{32'h428ab04b, 32'h422b593d, 32'h0, 32'h42043f7c, 32'h0, 32'h0, 32'h42a7878f, 32'h0};
test_input[4280:4287] = '{32'h41abd704, 32'h427564f1, 32'h415b45fe, 32'hc246d0f9, 32'hc234fece, 32'h42ae67df, 32'hc1b636c3, 32'h41984091};
test_output[4280:4287] = '{32'h41abd704, 32'h427564f1, 32'h415b45fe, 32'h0, 32'h0, 32'h42ae67df, 32'h0, 32'h41984091};
test_input[4288:4295] = '{32'hc26a80a3, 32'h42bce936, 32'h42b2da4d, 32'h42823ec0, 32'hc22c8fb6, 32'h417c5ff5, 32'hc221cabf, 32'hc29cb2a6};
test_output[4288:4295] = '{32'h0, 32'h42bce936, 32'h42b2da4d, 32'h42823ec0, 32'h0, 32'h417c5ff5, 32'h0, 32'h0};
test_input[4296:4303] = '{32'h42a7ab1e, 32'h42409d56, 32'hc26757f1, 32'h4281c6e9, 32'h42338f39, 32'h4281f7a4, 32'h4225c1cb, 32'hc128fc46};
test_output[4296:4303] = '{32'h42a7ab1e, 32'h42409d56, 32'h0, 32'h4281c6e9, 32'h42338f39, 32'h4281f7a4, 32'h4225c1cb, 32'h0};
test_input[4304:4311] = '{32'h4214a7d6, 32'h42b3e20f, 32'hc1c63a58, 32'hc1bc094f, 32'h42946f06, 32'h42322a76, 32'hc23988a2, 32'h42af8d2a};
test_output[4304:4311] = '{32'h4214a7d6, 32'h42b3e20f, 32'h0, 32'h0, 32'h42946f06, 32'h42322a76, 32'h0, 32'h42af8d2a};
test_input[4312:4319] = '{32'h42bdb3b8, 32'h42439940, 32'hc110e7fb, 32'h423eb819, 32'hc2a618a4, 32'hc2397335, 32'hc1b5fcd7, 32'hc1192ff0};
test_output[4312:4319] = '{32'h42bdb3b8, 32'h42439940, 32'h0, 32'h423eb819, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4320:4327] = '{32'hc2a44c7a, 32'hc24f5337, 32'h414180f5, 32'hc242a4ae, 32'h41e76f09, 32'hc2444b78, 32'hc1d37cb9, 32'h42a9baca};
test_output[4320:4327] = '{32'h0, 32'h0, 32'h414180f5, 32'h0, 32'h41e76f09, 32'h0, 32'h0, 32'h42a9baca};
test_input[4328:4335] = '{32'hc216ec5a, 32'hc1592cec, 32'hc20fbeb1, 32'hc2723c81, 32'hc0793bf1, 32'hc28c1e4e, 32'hc2343444, 32'h42c2c749};
test_output[4328:4335] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c2c749};
test_input[4336:4343] = '{32'hc279ced4, 32'hc1a4a5ba, 32'h419cd66d, 32'hc1196769, 32'h42c62bd2, 32'hc20d293c, 32'hc18becc8, 32'h4202bf34};
test_output[4336:4343] = '{32'h0, 32'h0, 32'h419cd66d, 32'h0, 32'h42c62bd2, 32'h0, 32'h0, 32'h4202bf34};
test_input[4344:4351] = '{32'h42a46004, 32'hc2849ee7, 32'hc257a568, 32'h41ab1cc8, 32'h40a8b965, 32'h420ad031, 32'h42985bd7, 32'h4197694f};
test_output[4344:4351] = '{32'h42a46004, 32'h0, 32'h0, 32'h41ab1cc8, 32'h40a8b965, 32'h420ad031, 32'h42985bd7, 32'h4197694f};
test_input[4352:4359] = '{32'hc2940a4a, 32'hc1902ed3, 32'h40a0eccb, 32'hc0e6a1c5, 32'h4235880a, 32'h419e6bfe, 32'h4287ccea, 32'h41dcf060};
test_output[4352:4359] = '{32'h0, 32'h0, 32'h40a0eccb, 32'h0, 32'h4235880a, 32'h419e6bfe, 32'h4287ccea, 32'h41dcf060};
test_input[4360:4367] = '{32'h4261b8fa, 32'hc1b3a96f, 32'hc2bd5c8c, 32'hc1dcf21b, 32'hc1be2a14, 32'h42b7d596, 32'h4278e027, 32'hc29ad42b};
test_output[4360:4367] = '{32'h4261b8fa, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b7d596, 32'h4278e027, 32'h0};
test_input[4368:4375] = '{32'hc0c08938, 32'hc1a15304, 32'h41a656be, 32'hc1702c9d, 32'hc22b5771, 32'h4259d86a, 32'h417adc4d, 32'h426d341a};
test_output[4368:4375] = '{32'h0, 32'h0, 32'h41a656be, 32'h0, 32'h0, 32'h4259d86a, 32'h417adc4d, 32'h426d341a};
test_input[4376:4383] = '{32'hc2bfba06, 32'h426c3946, 32'hc29462fd, 32'h424a75f7, 32'hc144ef6a, 32'hc2afe1ec, 32'hc293c1be, 32'hc2038ca2};
test_output[4376:4383] = '{32'h0, 32'h426c3946, 32'h0, 32'h424a75f7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4384:4391] = '{32'hc292b5b9, 32'h425f61a8, 32'hc2b263dc, 32'hc2b52f6c, 32'hc2c78c57, 32'hc21cfdbc, 32'hc093c474, 32'hc0e2a2f9};
test_output[4384:4391] = '{32'h0, 32'h425f61a8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4392:4399] = '{32'h4261f681, 32'h42831eaa, 32'h424c6d63, 32'hc17d2077, 32'h40bd5564, 32'h42093d0f, 32'hc262e0f8, 32'h42899a6f};
test_output[4392:4399] = '{32'h4261f681, 32'h42831eaa, 32'h424c6d63, 32'h0, 32'h40bd5564, 32'h42093d0f, 32'h0, 32'h42899a6f};
test_input[4400:4407] = '{32'h42b013aa, 32'hc16836db, 32'h3fd67dd9, 32'hc2866397, 32'h4224af32, 32'h429d7b9d, 32'hc11463a2, 32'h428ea3a5};
test_output[4400:4407] = '{32'h42b013aa, 32'h0, 32'h3fd67dd9, 32'h0, 32'h4224af32, 32'h429d7b9d, 32'h0, 32'h428ea3a5};
test_input[4408:4415] = '{32'h42c7e5ec, 32'h42b42420, 32'h41c8db6f, 32'hc1b5d53b, 32'hc2ad95de, 32'hc2987491, 32'h420693da, 32'hc212bbc7};
test_output[4408:4415] = '{32'h42c7e5ec, 32'h42b42420, 32'h41c8db6f, 32'h0, 32'h0, 32'h0, 32'h420693da, 32'h0};
test_input[4416:4423] = '{32'hc2864c4e, 32'hc28ab78b, 32'hc0698a41, 32'hc2943294, 32'h429afc80, 32'hc2b965fe, 32'h41835e43, 32'h42af16e5};
test_output[4416:4423] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429afc80, 32'h0, 32'h41835e43, 32'h42af16e5};
test_input[4424:4431] = '{32'hc238931e, 32'h42013a16, 32'h419c0a19, 32'h423bc579, 32'hc2062508, 32'hc2104611, 32'hc2c0cd1d, 32'hc23e008b};
test_output[4424:4431] = '{32'h0, 32'h42013a16, 32'h419c0a19, 32'h423bc579, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4432:4439] = '{32'hc2a2f3cd, 32'hc281c2dd, 32'hc21d4e32, 32'h42bea7e5, 32'hc2b3b80e, 32'hc1546d8a, 32'h420ab173, 32'h4229e40a};
test_output[4432:4439] = '{32'h0, 32'h0, 32'h0, 32'h42bea7e5, 32'h0, 32'h0, 32'h420ab173, 32'h4229e40a};
test_input[4440:4447] = '{32'h42510494, 32'hc2523f44, 32'h41d44320, 32'h42a7bc8c, 32'h41cb02dd, 32'h420e53c5, 32'hc196796d, 32'h4240f0dd};
test_output[4440:4447] = '{32'h42510494, 32'h0, 32'h41d44320, 32'h42a7bc8c, 32'h41cb02dd, 32'h420e53c5, 32'h0, 32'h4240f0dd};
test_input[4448:4455] = '{32'hc268d7e0, 32'hc135275e, 32'h4217333d, 32'h4180b9ca, 32'h4295a8de, 32'hc2a7a6ba, 32'h42ab172d, 32'h42c26b38};
test_output[4448:4455] = '{32'h0, 32'h0, 32'h4217333d, 32'h4180b9ca, 32'h4295a8de, 32'h0, 32'h42ab172d, 32'h42c26b38};
test_input[4456:4463] = '{32'hc1a970d5, 32'hc23d2753, 32'hc2885900, 32'hc2b0c53c, 32'h4207dc73, 32'hc24bff62, 32'h42b01fd9, 32'hc226c073};
test_output[4456:4463] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4207dc73, 32'h0, 32'h42b01fd9, 32'h0};
test_input[4464:4471] = '{32'hc0c50030, 32'hc2bdebae, 32'h4103aa3f, 32'hc29e08e9, 32'h429070c0, 32'h424d5093, 32'h424251ff, 32'h41c50eee};
test_output[4464:4471] = '{32'h0, 32'h0, 32'h4103aa3f, 32'h0, 32'h429070c0, 32'h424d5093, 32'h424251ff, 32'h41c50eee};
test_input[4472:4479] = '{32'hc2746650, 32'h420ed568, 32'h42c401d1, 32'h422e570c, 32'h410f793e, 32'h4237f173, 32'h428daaba, 32'h4223577a};
test_output[4472:4479] = '{32'h0, 32'h420ed568, 32'h42c401d1, 32'h422e570c, 32'h410f793e, 32'h4237f173, 32'h428daaba, 32'h4223577a};
test_input[4480:4487] = '{32'hc0e873c6, 32'h42987401, 32'hc105c28c, 32'hc139337e, 32'hc22e5929, 32'h42442dd3, 32'h3ff7d6c5, 32'hc2961861};
test_output[4480:4487] = '{32'h0, 32'h42987401, 32'h0, 32'h0, 32'h0, 32'h42442dd3, 32'h3ff7d6c5, 32'h0};
test_input[4488:4495] = '{32'hc200977a, 32'h41b3c621, 32'h41a8c6bb, 32'hc21be1bd, 32'h42b34739, 32'hc29b2a40, 32'hc2369469, 32'hc01c88f8};
test_output[4488:4495] = '{32'h0, 32'h41b3c621, 32'h41a8c6bb, 32'h0, 32'h42b34739, 32'h0, 32'h0, 32'h0};
test_input[4496:4503] = '{32'hc22e6375, 32'hc2592f16, 32'hc2995a1f, 32'hc2b5e8e6, 32'hc2b1ba86, 32'hc2752871, 32'hc28c6fa4, 32'hc180e110};
test_output[4496:4503] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4504:4511] = '{32'h427d65d1, 32'h42a34086, 32'hc2b254d3, 32'hc283ea15, 32'h4232ddf5, 32'hc2b5cf88, 32'h42c32dc7, 32'h4143f8d8};
test_output[4504:4511] = '{32'h427d65d1, 32'h42a34086, 32'h0, 32'h0, 32'h4232ddf5, 32'h0, 32'h42c32dc7, 32'h4143f8d8};
test_input[4512:4519] = '{32'h428c4c2d, 32'hc1d79dce, 32'hc1a1709a, 32'h419cd221, 32'h42bbb108, 32'h405aba78, 32'hc122b39e, 32'h426903cb};
test_output[4512:4519] = '{32'h428c4c2d, 32'h0, 32'h0, 32'h419cd221, 32'h42bbb108, 32'h405aba78, 32'h0, 32'h426903cb};
test_input[4520:4527] = '{32'hc2a07dc3, 32'h422f6f59, 32'h42bcde40, 32'hc25b6983, 32'h4227ef75, 32'h418d9ea2, 32'hc22fcdd1, 32'hc27785be};
test_output[4520:4527] = '{32'h0, 32'h422f6f59, 32'h42bcde40, 32'h0, 32'h4227ef75, 32'h418d9ea2, 32'h0, 32'h0};
test_input[4528:4535] = '{32'h42950752, 32'h4260aa07, 32'h42504b69, 32'hc2597d66, 32'h42bb5108, 32'hc28cc7c6, 32'hc2b12557, 32'h42c51b3a};
test_output[4528:4535] = '{32'h42950752, 32'h4260aa07, 32'h42504b69, 32'h0, 32'h42bb5108, 32'h0, 32'h0, 32'h42c51b3a};
test_input[4536:4543] = '{32'hc23f33ac, 32'h427ecfb3, 32'hc2c4bd84, 32'h4297580c, 32'h42235485, 32'hc122e4df, 32'hc1b7400a, 32'hc226d55d};
test_output[4536:4543] = '{32'h0, 32'h427ecfb3, 32'h0, 32'h4297580c, 32'h42235485, 32'h0, 32'h0, 32'h0};
test_input[4544:4551] = '{32'hc202602a, 32'h42873e7d, 32'hc1c5ea69, 32'hc218dfd7, 32'h4227062d, 32'h40db04f6, 32'h41102a9a, 32'hbf22ff1c};
test_output[4544:4551] = '{32'h0, 32'h42873e7d, 32'h0, 32'h0, 32'h4227062d, 32'h40db04f6, 32'h41102a9a, 32'h0};
test_input[4552:4559] = '{32'hc23da72c, 32'h42b23a86, 32'h4284f5fa, 32'h42bcd020, 32'hc25b7f04, 32'hc248aed8, 32'hc119d174, 32'h42815beb};
test_output[4552:4559] = '{32'h0, 32'h42b23a86, 32'h4284f5fa, 32'h42bcd020, 32'h0, 32'h0, 32'h0, 32'h42815beb};
test_input[4560:4567] = '{32'hc1bdb5d0, 32'hc2a34599, 32'hc18eec1d, 32'h415bed29, 32'h429dad1b, 32'h41a3f0cd, 32'hc23b1e21, 32'h41e1fb11};
test_output[4560:4567] = '{32'h0, 32'h0, 32'h0, 32'h415bed29, 32'h429dad1b, 32'h41a3f0cd, 32'h0, 32'h41e1fb11};
test_input[4568:4575] = '{32'hc2a45b73, 32'hc231345a, 32'hc2125251, 32'hc218cd50, 32'h4259ba03, 32'hc1fc5610, 32'h42c1452e, 32'hc20cd762};
test_output[4568:4575] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4259ba03, 32'h0, 32'h42c1452e, 32'h0};
test_input[4576:4583] = '{32'hc20107fa, 32'h421d7eaf, 32'h429c09e2, 32'hc1bd4a6c, 32'hc2783817, 32'hc2af0f4f, 32'hc21ac227, 32'h412113f2};
test_output[4576:4583] = '{32'h0, 32'h421d7eaf, 32'h429c09e2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h412113f2};
test_input[4584:4591] = '{32'h4216f9e5, 32'hc177ec75, 32'h42a657b3, 32'h41f0b172, 32'hc2590f76, 32'h42c5d6e3, 32'h42bdc178, 32'h42a2a81e};
test_output[4584:4591] = '{32'h4216f9e5, 32'h0, 32'h42a657b3, 32'h41f0b172, 32'h0, 32'h42c5d6e3, 32'h42bdc178, 32'h42a2a81e};
test_input[4592:4599] = '{32'h42b98844, 32'hc29257e0, 32'hc215219c, 32'h42350bed, 32'hc285cdb1, 32'hc219524a, 32'hc2acc843, 32'h415c7d24};
test_output[4592:4599] = '{32'h42b98844, 32'h0, 32'h0, 32'h42350bed, 32'h0, 32'h0, 32'h0, 32'h415c7d24};
test_input[4600:4607] = '{32'hc2aaa49b, 32'hc2be8691, 32'hc05f0dcf, 32'h4208c555, 32'hc28adbbe, 32'hc2c70c74, 32'hc210ad7d, 32'hc1c9189e};
test_output[4600:4607] = '{32'h0, 32'h0, 32'h0, 32'h4208c555, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4608:4615] = '{32'h40ddd2bb, 32'hc2a4a580, 32'hc249afcd, 32'hc299dd18, 32'h41ca71e3, 32'h4164bcce, 32'h42bd6d16, 32'hc24b03b4};
test_output[4608:4615] = '{32'h40ddd2bb, 32'h0, 32'h0, 32'h0, 32'h41ca71e3, 32'h4164bcce, 32'h42bd6d16, 32'h0};
test_input[4616:4623] = '{32'h4283fa6a, 32'h42894bba, 32'hc283d028, 32'hc20825f6, 32'hc19d1bb9, 32'h422c18bc, 32'hc15b927a, 32'h3f45e759};
test_output[4616:4623] = '{32'h4283fa6a, 32'h42894bba, 32'h0, 32'h0, 32'h0, 32'h422c18bc, 32'h0, 32'h3f45e759};
test_input[4624:4631] = '{32'h424b828e, 32'hc26f9329, 32'h4208a2d6, 32'hc2c4ed19, 32'hc1ae743f, 32'hbf3d64f6, 32'h3fcbd8d5, 32'h4219a5db};
test_output[4624:4631] = '{32'h424b828e, 32'h0, 32'h4208a2d6, 32'h0, 32'h0, 32'h0, 32'h3fcbd8d5, 32'h4219a5db};
test_input[4632:4639] = '{32'h429d53b1, 32'h421d36a6, 32'h42b4606e, 32'hc25d0248, 32'hc29d392b, 32'hc24075b5, 32'h424a4ffd, 32'h425f6429};
test_output[4632:4639] = '{32'h429d53b1, 32'h421d36a6, 32'h42b4606e, 32'h0, 32'h0, 32'h0, 32'h424a4ffd, 32'h425f6429};
test_input[4640:4647] = '{32'h411c95da, 32'h426487ee, 32'h407ceadd, 32'hc263840e, 32'h41e11bf0, 32'h41d5fd51, 32'hc2213285, 32'hc2b85be6};
test_output[4640:4647] = '{32'h411c95da, 32'h426487ee, 32'h407ceadd, 32'h0, 32'h41e11bf0, 32'h41d5fd51, 32'h0, 32'h0};
test_input[4648:4655] = '{32'h41dc2c73, 32'hc29d6c27, 32'h41827374, 32'h4293a06a, 32'hc2bd47e5, 32'hc0df49a7, 32'h4251837c, 32'h428ae1ea};
test_output[4648:4655] = '{32'h41dc2c73, 32'h0, 32'h41827374, 32'h4293a06a, 32'h0, 32'h0, 32'h4251837c, 32'h428ae1ea};
test_input[4656:4663] = '{32'h428eb660, 32'hc2317dfd, 32'hc21226a9, 32'h424ca0c3, 32'hc2b53923, 32'hc1e455b2, 32'h42c7be53, 32'hbfc074a9};
test_output[4656:4663] = '{32'h428eb660, 32'h0, 32'h0, 32'h424ca0c3, 32'h0, 32'h0, 32'h42c7be53, 32'h0};
test_input[4664:4671] = '{32'h41c2832a, 32'h41f780cd, 32'hc15d5eb2, 32'hc207d597, 32'h42896609, 32'h4289180a, 32'h41c50bb2, 32'hc2c59ee8};
test_output[4664:4671] = '{32'h41c2832a, 32'h41f780cd, 32'h0, 32'h0, 32'h42896609, 32'h4289180a, 32'h41c50bb2, 32'h0};
test_input[4672:4679] = '{32'hc284676c, 32'hc23d8e62, 32'h41b3b15b, 32'hc07ba5bc, 32'hc2960b9b, 32'hc2334035, 32'h4297d426, 32'hc27de26f};
test_output[4672:4679] = '{32'h0, 32'h0, 32'h41b3b15b, 32'h0, 32'h0, 32'h0, 32'h4297d426, 32'h0};
test_input[4680:4687] = '{32'h4293d541, 32'hc264454a, 32'h42ab82b9, 32'h42457a5b, 32'h42b5c7b7, 32'hc1c6f6f9, 32'hc1831634, 32'h3f0001a4};
test_output[4680:4687] = '{32'h4293d541, 32'h0, 32'h42ab82b9, 32'h42457a5b, 32'h42b5c7b7, 32'h0, 32'h0, 32'h3f0001a4};
test_input[4688:4695] = '{32'h4295ace5, 32'h423bfdca, 32'h42a06bfd, 32'hc2327786, 32'h400b982d, 32'h42c03483, 32'hc20a4403, 32'hc2abfe77};
test_output[4688:4695] = '{32'h4295ace5, 32'h423bfdca, 32'h42a06bfd, 32'h0, 32'h400b982d, 32'h42c03483, 32'h0, 32'h0};
test_input[4696:4703] = '{32'hc19697aa, 32'hc2ba99e3, 32'hc18a2413, 32'h425416ae, 32'hc1a3f85f, 32'h425e9045, 32'h42bd4083, 32'h421f726a};
test_output[4696:4703] = '{32'h0, 32'h0, 32'h0, 32'h425416ae, 32'h0, 32'h425e9045, 32'h42bd4083, 32'h421f726a};
test_input[4704:4711] = '{32'h42217308, 32'hc1c4536a, 32'hc2709584, 32'h42bda1df, 32'h407d50d8, 32'hc2a15edf, 32'h42a50dde, 32'hc09b8e02};
test_output[4704:4711] = '{32'h42217308, 32'h0, 32'h0, 32'h42bda1df, 32'h407d50d8, 32'h0, 32'h42a50dde, 32'h0};
test_input[4712:4719] = '{32'h42b5fcec, 32'h42b2c836, 32'hc2918375, 32'hc210c0c6, 32'hbfdf1a32, 32'hc11a0e68, 32'hc09d4a3b, 32'h3eb1ca26};
test_output[4712:4719] = '{32'h42b5fcec, 32'h42b2c836, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3eb1ca26};
test_input[4720:4727] = '{32'hc040f5b5, 32'h4177e242, 32'h4261ce10, 32'h42c6e601, 32'hc12faf45, 32'h42042bb2, 32'hc1fc9454, 32'h41fb4e5f};
test_output[4720:4727] = '{32'h0, 32'h4177e242, 32'h4261ce10, 32'h42c6e601, 32'h0, 32'h42042bb2, 32'h0, 32'h41fb4e5f};
test_input[4728:4735] = '{32'h408d75ab, 32'h428d69c8, 32'h4293c92b, 32'hc0b07ba9, 32'hc1e4cb00, 32'hc2b1538f, 32'hc2ad156d, 32'h428a92db};
test_output[4728:4735] = '{32'h408d75ab, 32'h428d69c8, 32'h4293c92b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428a92db};
test_input[4736:4743] = '{32'h4262aa93, 32'hc18b01f5, 32'h42a15dd8, 32'h421be18e, 32'h40487be6, 32'h42bee9b6, 32'h415261cc, 32'hc2adcb05};
test_output[4736:4743] = '{32'h4262aa93, 32'h0, 32'h42a15dd8, 32'h421be18e, 32'h40487be6, 32'h42bee9b6, 32'h415261cc, 32'h0};
test_input[4744:4751] = '{32'h4290a2b9, 32'h41b6daeb, 32'hc235392b, 32'hc2a2cb38, 32'hc15be3df, 32'hc2bb0c27, 32'hc12967a5, 32'hc106f3e9};
test_output[4744:4751] = '{32'h4290a2b9, 32'h41b6daeb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4752:4759] = '{32'h42b71052, 32'hc2a395c9, 32'h426ab4f1, 32'h421011e5, 32'h421de407, 32'hc280da6e, 32'hc291e815, 32'h42bee394};
test_output[4752:4759] = '{32'h42b71052, 32'h0, 32'h426ab4f1, 32'h421011e5, 32'h421de407, 32'h0, 32'h0, 32'h42bee394};
test_input[4760:4767] = '{32'h42b5589d, 32'hc294d8fb, 32'h42a0bea9, 32'h41192555, 32'hc1c56b8c, 32'hc2402b4b, 32'hc232de11, 32'hc2a5ac2c};
test_output[4760:4767] = '{32'h42b5589d, 32'h0, 32'h42a0bea9, 32'h41192555, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[4768:4775] = '{32'hc2898c13, 32'h4289d6ff, 32'hc05cadda, 32'h429d15be, 32'hc13ef545, 32'h42553269, 32'h41071b6d, 32'hc291a92d};
test_output[4768:4775] = '{32'h0, 32'h4289d6ff, 32'h0, 32'h429d15be, 32'h0, 32'h42553269, 32'h41071b6d, 32'h0};
test_input[4776:4783] = '{32'hc2b7b5cc, 32'hc1cb86af, 32'hc267795a, 32'hc29d756b, 32'hc19f9cad, 32'h41ba4055, 32'hc251e5d3, 32'hc1a6e130};
test_output[4776:4783] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ba4055, 32'h0, 32'h0};
test_input[4784:4791] = '{32'hc2bb574f, 32'h4228280b, 32'hc2891a93, 32'h419d64f3, 32'hc16f5353, 32'hc1f9e9e2, 32'hc2ac6220, 32'h4225dab8};
test_output[4784:4791] = '{32'h0, 32'h4228280b, 32'h0, 32'h419d64f3, 32'h0, 32'h0, 32'h0, 32'h4225dab8};
test_input[4792:4799] = '{32'hc27051b0, 32'h423f8bc7, 32'h3f8a0bdc, 32'h424b1b39, 32'h42a12a93, 32'hc209988d, 32'h42a2762b, 32'hc2373877};
test_output[4792:4799] = '{32'h0, 32'h423f8bc7, 32'h3f8a0bdc, 32'h424b1b39, 32'h42a12a93, 32'h0, 32'h42a2762b, 32'h0};
test_input[4800:4807] = '{32'h42658664, 32'h40f1da72, 32'hc28d45eb, 32'h42b5d263, 32'h421ad9c1, 32'hc1b4a952, 32'hc2358c00, 32'hc28cea66};
test_output[4800:4807] = '{32'h42658664, 32'h40f1da72, 32'h0, 32'h42b5d263, 32'h421ad9c1, 32'h0, 32'h0, 32'h0};
test_input[4808:4815] = '{32'h428981d9, 32'hc108696f, 32'hc1c938cd, 32'h423c66b0, 32'hc2767a13, 32'h4208ab44, 32'hc2a4f234, 32'hc2a585e5};
test_output[4808:4815] = '{32'h428981d9, 32'h0, 32'h0, 32'h423c66b0, 32'h0, 32'h4208ab44, 32'h0, 32'h0};
test_input[4816:4823] = '{32'h42a042b8, 32'hc2854fec, 32'h42c7a6ae, 32'hc1c5a2ff, 32'hc19e6729, 32'hc1413487, 32'hbfb41243, 32'h428c69e6};
test_output[4816:4823] = '{32'h42a042b8, 32'h0, 32'h42c7a6ae, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428c69e6};
test_input[4824:4831] = '{32'hc210ec5e, 32'h42be5a67, 32'hc299e3db, 32'h4040fa96, 32'hc11b7520, 32'h42a01ad1, 32'hc24c74c8, 32'h42801f51};
test_output[4824:4831] = '{32'h0, 32'h42be5a67, 32'h0, 32'h4040fa96, 32'h0, 32'h42a01ad1, 32'h0, 32'h42801f51};
test_input[4832:4839] = '{32'hc20256d5, 32'hc293ba1a, 32'h42a6be35, 32'h42a27fde, 32'hc202d51d, 32'hc2c3af51, 32'hc2a93b20, 32'h41c95a6c};
test_output[4832:4839] = '{32'h0, 32'h0, 32'h42a6be35, 32'h42a27fde, 32'h0, 32'h0, 32'h0, 32'h41c95a6c};
test_input[4840:4847] = '{32'hc1f3c85f, 32'hc2470ca6, 32'hc29e1bb7, 32'hc29367d4, 32'hc2765314, 32'hc2c51154, 32'h414043a7, 32'h420fbb03};
test_output[4840:4847] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h414043a7, 32'h420fbb03};
test_input[4848:4855] = '{32'h428c9ead, 32'h400b796b, 32'h42a3538a, 32'h4210e8b7, 32'h4260a37d, 32'h41e9dab6, 32'hc1aaef3a, 32'hc05efee1};
test_output[4848:4855] = '{32'h428c9ead, 32'h400b796b, 32'h42a3538a, 32'h4210e8b7, 32'h4260a37d, 32'h41e9dab6, 32'h0, 32'h0};
test_input[4856:4863] = '{32'hc263c164, 32'hc29e1869, 32'hc2823462, 32'hc186043d, 32'hc23022c8, 32'hc2824344, 32'hc29806d3, 32'h41ab0731};
test_output[4856:4863] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ab0731};
test_input[4864:4871] = '{32'hc2a2f7dc, 32'hc2197430, 32'h429d8123, 32'hc1dac7fa, 32'hc23c6d05, 32'h41b82522, 32'h4146a5df, 32'hc2b67f29};
test_output[4864:4871] = '{32'h0, 32'h0, 32'h429d8123, 32'h0, 32'h0, 32'h41b82522, 32'h4146a5df, 32'h0};
test_input[4872:4879] = '{32'hc2bc3823, 32'h419c6777, 32'h4284e4a1, 32'h42a51f8e, 32'h42b91143, 32'hc20d98af, 32'hc2c2b6d2, 32'h42aa0334};
test_output[4872:4879] = '{32'h0, 32'h419c6777, 32'h4284e4a1, 32'h42a51f8e, 32'h42b91143, 32'h0, 32'h0, 32'h42aa0334};
test_input[4880:4887] = '{32'h424f5879, 32'h41d3c3da, 32'hc2c1b20c, 32'hbe8d4f0f, 32'h4215500a, 32'h42a4282f, 32'hc2b4be50, 32'h427ac177};
test_output[4880:4887] = '{32'h424f5879, 32'h41d3c3da, 32'h0, 32'h0, 32'h4215500a, 32'h42a4282f, 32'h0, 32'h427ac177};
test_input[4888:4895] = '{32'hc2aab029, 32'hc16e5df5, 32'h4165592d, 32'h42a13b33, 32'h42c49a76, 32'h42bc5267, 32'h428ec4c6, 32'h42c2d43e};
test_output[4888:4895] = '{32'h0, 32'h0, 32'h4165592d, 32'h42a13b33, 32'h42c49a76, 32'h42bc5267, 32'h428ec4c6, 32'h42c2d43e};
test_input[4896:4903] = '{32'h4281eab6, 32'hc2290bfb, 32'hc21e9745, 32'hc22b9c20, 32'hc2428891, 32'hc27520fe, 32'h4299892b, 32'h42b7466a};
test_output[4896:4903] = '{32'h4281eab6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4299892b, 32'h42b7466a};
test_input[4904:4911] = '{32'hc2172dbe, 32'hc293062b, 32'h4296554c, 32'hc2a3a49d, 32'h42c4acee, 32'h424517f2, 32'h42aba6ce, 32'h41b787e5};
test_output[4904:4911] = '{32'h0, 32'h0, 32'h4296554c, 32'h0, 32'h42c4acee, 32'h424517f2, 32'h42aba6ce, 32'h41b787e5};
test_input[4912:4919] = '{32'h42109f8e, 32'h42432c30, 32'h42667094, 32'hc2bc2c41, 32'hc271894d, 32'h409fc483, 32'h42828f4a, 32'hc2801794};
test_output[4912:4919] = '{32'h42109f8e, 32'h42432c30, 32'h42667094, 32'h0, 32'h0, 32'h409fc483, 32'h42828f4a, 32'h0};
test_input[4920:4927] = '{32'h42703b8c, 32'hc2336f23, 32'h408e2610, 32'h429a6d76, 32'hc15af629, 32'hc1c714fb, 32'hc2586a88, 32'h4207bcd2};
test_output[4920:4927] = '{32'h42703b8c, 32'h0, 32'h408e2610, 32'h429a6d76, 32'h0, 32'h0, 32'h0, 32'h4207bcd2};
test_input[4928:4935] = '{32'h42aebbd7, 32'hbf7135d6, 32'h4205b6f1, 32'h4243474d, 32'hc2c3db17, 32'hc238421d, 32'h42bc186d, 32'h424adb47};
test_output[4928:4935] = '{32'h42aebbd7, 32'h0, 32'h4205b6f1, 32'h4243474d, 32'h0, 32'h0, 32'h42bc186d, 32'h424adb47};
test_input[4936:4943] = '{32'h413d5a7c, 32'h420c2933, 32'h42b55411, 32'hc1f2b25e, 32'hc291a023, 32'hc2237172, 32'hbf90123a, 32'h423cc350};
test_output[4936:4943] = '{32'h413d5a7c, 32'h420c2933, 32'h42b55411, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423cc350};
test_input[4944:4951] = '{32'h422d3f4d, 32'h421950c8, 32'h3d4a3c7a, 32'hc2a0a3df, 32'h4133fef9, 32'h428d483d, 32'h4258303c, 32'hc2a906b4};
test_output[4944:4951] = '{32'h422d3f4d, 32'h421950c8, 32'h3d4a3c7a, 32'h0, 32'h4133fef9, 32'h428d483d, 32'h4258303c, 32'h0};
test_input[4952:4959] = '{32'hc193cd20, 32'h41c35a79, 32'h4205502c, 32'hc1cde7df, 32'hc285cfbf, 32'hc29e994c, 32'h424a99fe, 32'h40c5efe1};
test_output[4952:4959] = '{32'h0, 32'h41c35a79, 32'h4205502c, 32'h0, 32'h0, 32'h0, 32'h424a99fe, 32'h40c5efe1};
test_input[4960:4967] = '{32'h428b0d90, 32'h42558b59, 32'h4277dfe7, 32'hc1fda9fd, 32'h418ab609, 32'hc2ba156a, 32'hc1f5d5a3, 32'hc1a74b7c};
test_output[4960:4967] = '{32'h428b0d90, 32'h42558b59, 32'h4277dfe7, 32'h0, 32'h418ab609, 32'h0, 32'h0, 32'h0};
test_input[4968:4975] = '{32'h41991357, 32'hc0a68850, 32'hc249ab29, 32'h3ffa2bc1, 32'h42223ff5, 32'hc2bc2a5f, 32'h42a9b49f, 32'h422f578b};
test_output[4968:4975] = '{32'h41991357, 32'h0, 32'h0, 32'h3ffa2bc1, 32'h42223ff5, 32'h0, 32'h42a9b49f, 32'h422f578b};
test_input[4976:4983] = '{32'h41af7f3a, 32'h428a5c0e, 32'hc282dce1, 32'hbe91f8bd, 32'hc295f572, 32'h41773573, 32'h4290d0b5, 32'h4266b0a6};
test_output[4976:4983] = '{32'h41af7f3a, 32'h428a5c0e, 32'h0, 32'h0, 32'h0, 32'h41773573, 32'h4290d0b5, 32'h4266b0a6};
test_input[4984:4991] = '{32'h42966b97, 32'hc106835b, 32'hc171f049, 32'hc10554df, 32'hc0243d87, 32'hc0294ee6, 32'h40f3ffe7, 32'hc2b9e539};
test_output[4984:4991] = '{32'h42966b97, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40f3ffe7, 32'h0};
test_input[4992:4999] = '{32'hc1d146e4, 32'h410a5aef, 32'hc173c3a9, 32'hc2b8ef5d, 32'hc1c58c08, 32'hc2447b43, 32'hc29340cd, 32'hc0de0f8b};
test_output[4992:4999] = '{32'h0, 32'h410a5aef, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5000:5007] = '{32'hc1d202c7, 32'h428ac7fd, 32'hc2805b45, 32'hc1ab101f, 32'hc2be83ce, 32'h42abb035, 32'h41d63f30, 32'hc21e5c98};
test_output[5000:5007] = '{32'h0, 32'h428ac7fd, 32'h0, 32'h0, 32'h0, 32'h42abb035, 32'h41d63f30, 32'h0};
test_input[5008:5015] = '{32'hc282fc24, 32'hc2c78cbb, 32'h41a25c8b, 32'h42b645a8, 32'h426058fd, 32'hc293614b, 32'h40a00953, 32'hc21fec16};
test_output[5008:5015] = '{32'h0, 32'h0, 32'h41a25c8b, 32'h42b645a8, 32'h426058fd, 32'h0, 32'h40a00953, 32'h0};
test_input[5016:5023] = '{32'h417b84e5, 32'hc15b6ac0, 32'h42c7f74c, 32'h41c875aa, 32'hc2bb1c8a, 32'hc201ce78, 32'h4222ccce, 32'hc23c6570};
test_output[5016:5023] = '{32'h417b84e5, 32'h0, 32'h42c7f74c, 32'h41c875aa, 32'h0, 32'h0, 32'h4222ccce, 32'h0};
test_input[5024:5031] = '{32'hc2b6411c, 32'hc29d9c67, 32'h400c2398, 32'h42c3e81e, 32'hc221de24, 32'hc26db2cf, 32'h426f7e12, 32'hc2b3a5e3};
test_output[5024:5031] = '{32'h0, 32'h0, 32'h400c2398, 32'h42c3e81e, 32'h0, 32'h0, 32'h426f7e12, 32'h0};
test_input[5032:5039] = '{32'hc19f2eed, 32'h41681ac9, 32'h42a6fa88, 32'h4206f17a, 32'hc1356f7d, 32'hc2814f00, 32'hc2baaa8b, 32'hc1fc7356};
test_output[5032:5039] = '{32'h0, 32'h41681ac9, 32'h42a6fa88, 32'h4206f17a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5040:5047] = '{32'h405333f1, 32'h421b5e72, 32'hc2274a0c, 32'hc2844274, 32'hc174be49, 32'h42122f67, 32'hc2c1d06e, 32'h42693057};
test_output[5040:5047] = '{32'h405333f1, 32'h421b5e72, 32'h0, 32'h0, 32'h0, 32'h42122f67, 32'h0, 32'h42693057};
test_input[5048:5055] = '{32'hc29a6bb9, 32'h424ec4c0, 32'h42ac7ec3, 32'hc103afca, 32'h425cbe1b, 32'hc2a4d938, 32'h42a610ae, 32'h41de5dc9};
test_output[5048:5055] = '{32'h0, 32'h424ec4c0, 32'h42ac7ec3, 32'h0, 32'h425cbe1b, 32'h0, 32'h42a610ae, 32'h41de5dc9};
test_input[5056:5063] = '{32'h42845153, 32'hc29712f2, 32'hc28cf281, 32'h4285741a, 32'hc23472b0, 32'hc2830a1e, 32'h428e2125, 32'hc17c0ed1};
test_output[5056:5063] = '{32'h42845153, 32'h0, 32'h0, 32'h4285741a, 32'h0, 32'h0, 32'h428e2125, 32'h0};
test_input[5064:5071] = '{32'h41a8e0a2, 32'h420dc5d7, 32'hc24a72ad, 32'h4220d8d7, 32'h42859024, 32'h426e1a26, 32'h418c7dff, 32'hc1106597};
test_output[5064:5071] = '{32'h41a8e0a2, 32'h420dc5d7, 32'h0, 32'h4220d8d7, 32'h42859024, 32'h426e1a26, 32'h418c7dff, 32'h0};
test_input[5072:5079] = '{32'hc0b49bd0, 32'hc1d30697, 32'h42b20331, 32'hc20a2fb6, 32'hc23513cb, 32'hc24ec859, 32'h42bcf65c, 32'h415564c1};
test_output[5072:5079] = '{32'h0, 32'h0, 32'h42b20331, 32'h0, 32'h0, 32'h0, 32'h42bcf65c, 32'h415564c1};
test_input[5080:5087] = '{32'hc2a4d24f, 32'h41dea38c, 32'h411f706a, 32'hc2ac6f5e, 32'h4213d054, 32'hc137f883, 32'h427706fb, 32'hc18151fe};
test_output[5080:5087] = '{32'h0, 32'h41dea38c, 32'h411f706a, 32'h0, 32'h4213d054, 32'h0, 32'h427706fb, 32'h0};
test_input[5088:5095] = '{32'h42a206fb, 32'h42c30a1b, 32'h428c9f80, 32'hc20a7384, 32'hc2a92dfe, 32'h42c52a32, 32'hc1b9e777, 32'hc1c72b40};
test_output[5088:5095] = '{32'h42a206fb, 32'h42c30a1b, 32'h428c9f80, 32'h0, 32'h0, 32'h42c52a32, 32'h0, 32'h0};
test_input[5096:5103] = '{32'hc23c599f, 32'h4234ca86, 32'hc2c32420, 32'h42691354, 32'hc21ea448, 32'h428b6ef0, 32'h4181e9ad, 32'hc219b408};
test_output[5096:5103] = '{32'h0, 32'h4234ca86, 32'h0, 32'h42691354, 32'h0, 32'h428b6ef0, 32'h4181e9ad, 32'h0};
test_input[5104:5111] = '{32'h422d1e91, 32'hc28f5fa0, 32'h40b2d132, 32'hc285ee7d, 32'hc1af0025, 32'hc28e17ca, 32'h42996d36, 32'hc21e6d59};
test_output[5104:5111] = '{32'h422d1e91, 32'h0, 32'h40b2d132, 32'h0, 32'h0, 32'h0, 32'h42996d36, 32'h0};
test_input[5112:5119] = '{32'h427000e9, 32'h3e9635eb, 32'hc29f52f2, 32'h4180150f, 32'hc2a5de01, 32'h42513b91, 32'hc29995b2, 32'h4101546a};
test_output[5112:5119] = '{32'h427000e9, 32'h3e9635eb, 32'h0, 32'h4180150f, 32'h0, 32'h42513b91, 32'h0, 32'h4101546a};
test_input[5120:5127] = '{32'hc25ba2f8, 32'h4254ecdd, 32'h41a4078e, 32'h426cf5b6, 32'hc173e477, 32'hc043d85f, 32'h420f7929, 32'h42bce803};
test_output[5120:5127] = '{32'h0, 32'h4254ecdd, 32'h41a4078e, 32'h426cf5b6, 32'h0, 32'h0, 32'h420f7929, 32'h42bce803};
test_input[5128:5135] = '{32'hc27f7491, 32'h41bd91da, 32'hc28fcea1, 32'hc25272f8, 32'h41f1b13f, 32'hc1a0d3f1, 32'h4217c12a, 32'h42ba365d};
test_output[5128:5135] = '{32'h0, 32'h41bd91da, 32'h0, 32'h0, 32'h41f1b13f, 32'h0, 32'h4217c12a, 32'h42ba365d};
test_input[5136:5143] = '{32'hc27c7bda, 32'hc2887e78, 32'h4287fe09, 32'hc25b2ff4, 32'h411ba5fd, 32'hc295b04b, 32'h4286ba6e, 32'h41920b55};
test_output[5136:5143] = '{32'h0, 32'h0, 32'h4287fe09, 32'h0, 32'h411ba5fd, 32'h0, 32'h4286ba6e, 32'h41920b55};
test_input[5144:5151] = '{32'h424a4779, 32'h424163bd, 32'h413e2862, 32'hc29a3dfa, 32'hc0abc10d, 32'h42075bf2, 32'h417d6827, 32'h4217b84b};
test_output[5144:5151] = '{32'h424a4779, 32'h424163bd, 32'h413e2862, 32'h0, 32'h0, 32'h42075bf2, 32'h417d6827, 32'h4217b84b};
test_input[5152:5159] = '{32'h424e0dea, 32'h42162b3a, 32'h42320291, 32'hc2142f58, 32'hc2222f1c, 32'h40588b43, 32'h42c303f3, 32'hbfd84a3f};
test_output[5152:5159] = '{32'h424e0dea, 32'h42162b3a, 32'h42320291, 32'h0, 32'h0, 32'h40588b43, 32'h42c303f3, 32'h0};
test_input[5160:5167] = '{32'hc2bb4eff, 32'hc1589449, 32'h42b1dc95, 32'hc2b1cef5, 32'h4288098f, 32'hc26076cd, 32'h42a0b505, 32'h41e85f4c};
test_output[5160:5167] = '{32'h0, 32'h0, 32'h42b1dc95, 32'h0, 32'h4288098f, 32'h0, 32'h42a0b505, 32'h41e85f4c};
test_input[5168:5175] = '{32'h428ef687, 32'h4217fb4f, 32'h428e65f2, 32'h41712023, 32'hc2c0bc71, 32'h42553fb6, 32'h42b21f00, 32'h422387c0};
test_output[5168:5175] = '{32'h428ef687, 32'h4217fb4f, 32'h428e65f2, 32'h41712023, 32'h0, 32'h42553fb6, 32'h42b21f00, 32'h422387c0};
test_input[5176:5183] = '{32'hc1e36692, 32'hc24de9b0, 32'hc2b36375, 32'hc0ceb947, 32'h40b558bc, 32'hc25763c6, 32'hc2c0ce31, 32'h419aca43};
test_output[5176:5183] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40b558bc, 32'h0, 32'h0, 32'h419aca43};
test_input[5184:5191] = '{32'h41a86029, 32'h429b170c, 32'hc2ba317f, 32'hc137854a, 32'hc2ba15f1, 32'h41f3f613, 32'h4271e93f, 32'h425bca07};
test_output[5184:5191] = '{32'h41a86029, 32'h429b170c, 32'h0, 32'h0, 32'h0, 32'h41f3f613, 32'h4271e93f, 32'h425bca07};
test_input[5192:5199] = '{32'h422afb9f, 32'h42938c18, 32'h40fdc6e9, 32'h4188f8f7, 32'hc2139702, 32'hc21bc5be, 32'h4261b533, 32'h42c20ee8};
test_output[5192:5199] = '{32'h422afb9f, 32'h42938c18, 32'h40fdc6e9, 32'h4188f8f7, 32'h0, 32'h0, 32'h4261b533, 32'h42c20ee8};
test_input[5200:5207] = '{32'h4056c7c8, 32'h418f79e4, 32'hc20fe642, 32'h42015058, 32'hbfaa9b16, 32'hc1f3f3c0, 32'hc25a3eb1, 32'hc1ceca2a};
test_output[5200:5207] = '{32'h4056c7c8, 32'h418f79e4, 32'h0, 32'h42015058, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5208:5215] = '{32'hc11080cd, 32'h41c990e3, 32'h42ac5b15, 32'h427d1a94, 32'hc29f32c3, 32'hc28eb21e, 32'h42a5f025, 32'hc29f2da1};
test_output[5208:5215] = '{32'h0, 32'h41c990e3, 32'h42ac5b15, 32'h427d1a94, 32'h0, 32'h0, 32'h42a5f025, 32'h0};
test_input[5216:5223] = '{32'h40e2409b, 32'h42190342, 32'hc296a3ad, 32'h420e6d02, 32'h4190ae9b, 32'hbf51a2b0, 32'h41939845, 32'hc0702953};
test_output[5216:5223] = '{32'h40e2409b, 32'h42190342, 32'h0, 32'h420e6d02, 32'h4190ae9b, 32'h0, 32'h41939845, 32'h0};
test_input[5224:5231] = '{32'h427a1e88, 32'h428d0fc9, 32'hc286fb00, 32'h42b2feae, 32'hc26147e6, 32'hbfb06caa, 32'h418b1459, 32'h42950db8};
test_output[5224:5231] = '{32'h427a1e88, 32'h428d0fc9, 32'h0, 32'h42b2feae, 32'h0, 32'h0, 32'h418b1459, 32'h42950db8};
test_input[5232:5239] = '{32'h428bba92, 32'h40c1b7bc, 32'hc264e606, 32'hc2aa814b, 32'hc2464d25, 32'hc1ce3b2b, 32'h4259c6a8, 32'hc223daea};
test_output[5232:5239] = '{32'h428bba92, 32'h40c1b7bc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4259c6a8, 32'h0};
test_input[5240:5247] = '{32'hc1e8efcf, 32'hc234811f, 32'h42b23003, 32'h42396c6f, 32'hc2c68375, 32'h428f9b82, 32'h42a735e6, 32'h420a8a2f};
test_output[5240:5247] = '{32'h0, 32'h0, 32'h42b23003, 32'h42396c6f, 32'h0, 32'h428f9b82, 32'h42a735e6, 32'h420a8a2f};
test_input[5248:5255] = '{32'h421ebedd, 32'hc29db400, 32'hc1152562, 32'hc1c93a38, 32'h42900c44, 32'hc2186ff4, 32'h42ae8bde, 32'h423c5dba};
test_output[5248:5255] = '{32'h421ebedd, 32'h0, 32'h0, 32'h0, 32'h42900c44, 32'h0, 32'h42ae8bde, 32'h423c5dba};
test_input[5256:5263] = '{32'h41e9357a, 32'hc2a0ced9, 32'hc207bff8, 32'h421b3067, 32'hc27c9df7, 32'h4285acba, 32'h4214883e, 32'h403f3e4c};
test_output[5256:5263] = '{32'h41e9357a, 32'h0, 32'h0, 32'h421b3067, 32'h0, 32'h4285acba, 32'h4214883e, 32'h403f3e4c};
test_input[5264:5271] = '{32'hc2a125d7, 32'hc276e32e, 32'hc25fdeec, 32'h3ff0a096, 32'h40898008, 32'h429bbaa3, 32'hc2b67248, 32'h427393bd};
test_output[5264:5271] = '{32'h0, 32'h0, 32'h0, 32'h3ff0a096, 32'h40898008, 32'h429bbaa3, 32'h0, 32'h427393bd};
test_input[5272:5279] = '{32'h41b543e7, 32'hc13293e1, 32'hc28db7d7, 32'h423ffa6c, 32'hc1dc0290, 32'hc19d1182, 32'h4241e410, 32'h41e2c124};
test_output[5272:5279] = '{32'h41b543e7, 32'h0, 32'h0, 32'h423ffa6c, 32'h0, 32'h0, 32'h4241e410, 32'h41e2c124};
test_input[5280:5287] = '{32'hc26f9567, 32'h42a4beb6, 32'h405a0af5, 32'h42332286, 32'h41df7582, 32'hc184c1c9, 32'hc2b69258, 32'hc1dee1e5};
test_output[5280:5287] = '{32'h0, 32'h42a4beb6, 32'h405a0af5, 32'h42332286, 32'h41df7582, 32'h0, 32'h0, 32'h0};
test_input[5288:5295] = '{32'hc249ac11, 32'h426ce2f7, 32'h4290d8d4, 32'hc2b9e1c1, 32'hc2408b8b, 32'h42c3e075, 32'hc21f30ed, 32'hc2ada0fc};
test_output[5288:5295] = '{32'h0, 32'h426ce2f7, 32'h4290d8d4, 32'h0, 32'h0, 32'h42c3e075, 32'h0, 32'h0};
test_input[5296:5303] = '{32'h40446246, 32'hc25980ac, 32'hc24d2921, 32'hc2b3d39f, 32'h428226af, 32'h4280a1af, 32'h4281752c, 32'hc2543250};
test_output[5296:5303] = '{32'h40446246, 32'h0, 32'h0, 32'h0, 32'h428226af, 32'h4280a1af, 32'h4281752c, 32'h0};
test_input[5304:5311] = '{32'hc2bdb2cc, 32'hc242594f, 32'hc22ade71, 32'hc27565b8, 32'h42229ed3, 32'hc142c61a, 32'hc092fdf3, 32'h4284cee0};
test_output[5304:5311] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42229ed3, 32'h0, 32'h0, 32'h4284cee0};
test_input[5312:5319] = '{32'h423e3f0f, 32'h42bef1a8, 32'h42ad47dd, 32'hc1907610, 32'hc27e8c75, 32'h413ac0fe, 32'hc11b5f46, 32'hc230286f};
test_output[5312:5319] = '{32'h423e3f0f, 32'h42bef1a8, 32'h42ad47dd, 32'h0, 32'h0, 32'h413ac0fe, 32'h0, 32'h0};
test_input[5320:5327] = '{32'hc2226785, 32'hc2a52263, 32'hc25e6de7, 32'h3dd4d926, 32'h410c2838, 32'h4296081a, 32'hc24315eb, 32'h41fd2338};
test_output[5320:5327] = '{32'h0, 32'h0, 32'h0, 32'h3dd4d926, 32'h410c2838, 32'h4296081a, 32'h0, 32'h41fd2338};
test_input[5328:5335] = '{32'hc2896b63, 32'hc1d37aa9, 32'hc2a022f3, 32'hc22689b8, 32'h401bea30, 32'h428ab5d6, 32'h42befc61, 32'hc2c2b654};
test_output[5328:5335] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h401bea30, 32'h428ab5d6, 32'h42befc61, 32'h0};
test_input[5336:5343] = '{32'h42acdb03, 32'h42942746, 32'hc2b9884c, 32'h4265ea55, 32'hc1e7f3c8, 32'hc2b7fcb0, 32'hc238f2e9, 32'h429ab42b};
test_output[5336:5343] = '{32'h42acdb03, 32'h42942746, 32'h0, 32'h4265ea55, 32'h0, 32'h0, 32'h0, 32'h429ab42b};
test_input[5344:5351] = '{32'h413f50fe, 32'h41c9b343, 32'h42a3ec36, 32'hc2908da9, 32'h4284f794, 32'hc2001b2f, 32'h41bdfb4b, 32'h406397d0};
test_output[5344:5351] = '{32'h413f50fe, 32'h41c9b343, 32'h42a3ec36, 32'h0, 32'h4284f794, 32'h0, 32'h41bdfb4b, 32'h406397d0};
test_input[5352:5359] = '{32'hc2af6ba0, 32'hc2a07d97, 32'hc0e679ee, 32'hc20867b3, 32'h41f98593, 32'h418c9dc1, 32'hc2177661, 32'hc2c3465d};
test_output[5352:5359] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41f98593, 32'h418c9dc1, 32'h0, 32'h0};
test_input[5360:5367] = '{32'hc2a7cd8f, 32'h42ad7126, 32'h4014b8e0, 32'h42385a4f, 32'hc2a3c882, 32'h4246405e, 32'h42b9d22a, 32'hc1b9197b};
test_output[5360:5367] = '{32'h0, 32'h42ad7126, 32'h4014b8e0, 32'h42385a4f, 32'h0, 32'h4246405e, 32'h42b9d22a, 32'h0};
test_input[5368:5375] = '{32'h41c424f9, 32'h42a013e1, 32'h42a04369, 32'hc2a36ebd, 32'hc287765b, 32'h42a8c977, 32'hc1bdc878, 32'hc27cd6ea};
test_output[5368:5375] = '{32'h41c424f9, 32'h42a013e1, 32'h42a04369, 32'h0, 32'h0, 32'h42a8c977, 32'h0, 32'h0};
test_input[5376:5383] = '{32'hc2bd5bd4, 32'h42b99c8d, 32'h40eebdc1, 32'hc1efd12f, 32'hc2aa2eb7, 32'h4229bf78, 32'h41ec1307, 32'hc29a0532};
test_output[5376:5383] = '{32'h0, 32'h42b99c8d, 32'h40eebdc1, 32'h0, 32'h0, 32'h4229bf78, 32'h41ec1307, 32'h0};
test_input[5384:5391] = '{32'hc20cfbb3, 32'hc2c75bba, 32'h4209de84, 32'hc2ab2f39, 32'hc12f0833, 32'h4289c39f, 32'hc2986f0b, 32'hc1e8d322};
test_output[5384:5391] = '{32'h0, 32'h0, 32'h4209de84, 32'h0, 32'h0, 32'h4289c39f, 32'h0, 32'h0};
test_input[5392:5399] = '{32'hc1fd4854, 32'h42b48acb, 32'hc25bcffd, 32'hc1fca025, 32'hc1f62021, 32'h42c3fe06, 32'hc13d11f6, 32'hc118a796};
test_output[5392:5399] = '{32'h0, 32'h42b48acb, 32'h0, 32'h0, 32'h0, 32'h42c3fe06, 32'h0, 32'h0};
test_input[5400:5407] = '{32'h420dd15d, 32'h4292dcdf, 32'hc2c1f936, 32'hc2a11664, 32'h424c5e11, 32'h42506c7b, 32'h42c404bc, 32'h42a661c0};
test_output[5400:5407] = '{32'h420dd15d, 32'h4292dcdf, 32'h0, 32'h0, 32'h424c5e11, 32'h42506c7b, 32'h42c404bc, 32'h42a661c0};
test_input[5408:5415] = '{32'hc01ac833, 32'hc14be01b, 32'h3d949c4d, 32'h42ad5200, 32'hc1f254a2, 32'h426735f6, 32'h423972cd, 32'hc2977403};
test_output[5408:5415] = '{32'h0, 32'h0, 32'h3d949c4d, 32'h42ad5200, 32'h0, 32'h426735f6, 32'h423972cd, 32'h0};
test_input[5416:5423] = '{32'hc1f5bff3, 32'h4293213e, 32'hc1a8ca45, 32'hc29858ac, 32'hc2a5e043, 32'hc2638e21, 32'hc225097f, 32'h42701ed2};
test_output[5416:5423] = '{32'h0, 32'h4293213e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42701ed2};
test_input[5424:5431] = '{32'h42838f6e, 32'h42ac1b63, 32'hc1929d5f, 32'hc23110a2, 32'hc252ac62, 32'h42341fea, 32'h4289d2b9, 32'h428f99c4};
test_output[5424:5431] = '{32'h42838f6e, 32'h42ac1b63, 32'h0, 32'h0, 32'h0, 32'h42341fea, 32'h4289d2b9, 32'h428f99c4};
test_input[5432:5439] = '{32'hc1dffe4e, 32'hc095ae06, 32'hc1cf462c, 32'h42753997, 32'hc2649bc7, 32'hc2699f4e, 32'hc1082175, 32'h41b5a189};
test_output[5432:5439] = '{32'h0, 32'h0, 32'h0, 32'h42753997, 32'h0, 32'h0, 32'h0, 32'h41b5a189};
test_input[5440:5447] = '{32'h423dea49, 32'h429b43e5, 32'hc2634fe1, 32'hc2033586, 32'h4289a138, 32'h3f567a73, 32'hc2a2507d, 32'h4242e53b};
test_output[5440:5447] = '{32'h423dea49, 32'h429b43e5, 32'h0, 32'h0, 32'h4289a138, 32'h3f567a73, 32'h0, 32'h4242e53b};
test_input[5448:5455] = '{32'hc2b66714, 32'hc2130e75, 32'hc24f9b4e, 32'hc298b456, 32'h425d1f9d, 32'h42a32aba, 32'hc159f15d, 32'h42011dc3};
test_output[5448:5455] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h425d1f9d, 32'h42a32aba, 32'h0, 32'h42011dc3};
test_input[5456:5463] = '{32'hc2404338, 32'hc2b01803, 32'h42255837, 32'hc18154be, 32'hc2962c9b, 32'h42c28572, 32'hc1a6bea9, 32'hc271391f};
test_output[5456:5463] = '{32'h0, 32'h0, 32'h42255837, 32'h0, 32'h0, 32'h42c28572, 32'h0, 32'h0};
test_input[5464:5471] = '{32'hc1d9c2fe, 32'h42a52253, 32'hc2b74dec, 32'hc1214f0d, 32'hc25c1ff8, 32'h42132f1e, 32'hc284ba73, 32'h42994acf};
test_output[5464:5471] = '{32'h0, 32'h42a52253, 32'h0, 32'h0, 32'h0, 32'h42132f1e, 32'h0, 32'h42994acf};
test_input[5472:5479] = '{32'h4271e35e, 32'hc1bdd3d7, 32'h42b8c16d, 32'hc190a5a0, 32'hc2bb142b, 32'hc0bcb20e, 32'h42bb6005, 32'hc2074517};
test_output[5472:5479] = '{32'h4271e35e, 32'h0, 32'h42b8c16d, 32'h0, 32'h0, 32'h0, 32'h42bb6005, 32'h0};
test_input[5480:5487] = '{32'hc2118d2d, 32'hc29517e5, 32'h4207cc5b, 32'h42c28b96, 32'h41c514ef, 32'hc2847896, 32'hc2621189, 32'h42454f64};
test_output[5480:5487] = '{32'h0, 32'h0, 32'h4207cc5b, 32'h42c28b96, 32'h41c514ef, 32'h0, 32'h0, 32'h42454f64};
test_input[5488:5495] = '{32'hc270832f, 32'hc243f663, 32'hc24aac99, 32'hc28fe04f, 32'hc27bebd6, 32'hc27cd5b1, 32'hc18b42e5, 32'hc28eb3af};
test_output[5488:5495] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5496:5503] = '{32'hc24b2209, 32'h42b6d77d, 32'h419dffe8, 32'hc0d099d4, 32'hc2416333, 32'hc2a58959, 32'hc29a8158, 32'h4244292f};
test_output[5496:5503] = '{32'h0, 32'h42b6d77d, 32'h419dffe8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4244292f};
test_input[5504:5511] = '{32'h428221aa, 32'h41a04886, 32'hc1d13746, 32'hc231a6f9, 32'hc2792234, 32'hc29a3934, 32'h41a92640, 32'hc248d042};
test_output[5504:5511] = '{32'h428221aa, 32'h41a04886, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41a92640, 32'h0};
test_input[5512:5519] = '{32'h425b9138, 32'h42b668e3, 32'hc07ecbe0, 32'h4216c0e8, 32'h41f4b760, 32'hc25ba355, 32'h414e8f97, 32'h429522de};
test_output[5512:5519] = '{32'h425b9138, 32'h42b668e3, 32'h0, 32'h4216c0e8, 32'h41f4b760, 32'h0, 32'h414e8f97, 32'h429522de};
test_input[5520:5527] = '{32'h3fbfedee, 32'hc2438029, 32'hc26bdb9f, 32'hc1a79924, 32'hc27b5d65, 32'hc21b714e, 32'hc268ac8a, 32'h4242e417};
test_output[5520:5527] = '{32'h3fbfedee, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4242e417};
test_input[5528:5535] = '{32'h42c11ff2, 32'hc2b9f8f5, 32'hc0971c1c, 32'h42c52ba5, 32'hc217898f, 32'h42208920, 32'h428710e1, 32'h42514e8c};
test_output[5528:5535] = '{32'h42c11ff2, 32'h0, 32'h0, 32'h42c52ba5, 32'h0, 32'h42208920, 32'h428710e1, 32'h42514e8c};
test_input[5536:5543] = '{32'hc260908e, 32'hc20c8012, 32'hc0f46c17, 32'hc17d4da2, 32'hc1bf0d8d, 32'h4183b03e, 32'h42996200, 32'hc22c9d53};
test_output[5536:5543] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4183b03e, 32'h42996200, 32'h0};
test_input[5544:5551] = '{32'hc186afd2, 32'h41f1631e, 32'hc271f8e2, 32'h428c0389, 32'hc1d0c4f7, 32'hc29848bd, 32'hc10eb56b, 32'hc1cc5cb4};
test_output[5544:5551] = '{32'h0, 32'h41f1631e, 32'h0, 32'h428c0389, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5552:5559] = '{32'h41a2df3d, 32'hc19a5118, 32'hc1a3d50e, 32'h42a73acb, 32'hc111efe0, 32'hc26b0580, 32'h42998b89, 32'h42928a5d};
test_output[5552:5559] = '{32'h41a2df3d, 32'h0, 32'h0, 32'h42a73acb, 32'h0, 32'h0, 32'h42998b89, 32'h42928a5d};
test_input[5560:5567] = '{32'hc27f33c5, 32'hc28e964f, 32'hc2100601, 32'hc27c5c48, 32'h427a6beb, 32'h42139d78, 32'hc232fe44, 32'h4229f5af};
test_output[5560:5567] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h427a6beb, 32'h42139d78, 32'h0, 32'h4229f5af};
test_input[5568:5575] = '{32'h4271f81c, 32'hbe300891, 32'h425fd429, 32'hc2b36a62, 32'h423fa44b, 32'hc27ca315, 32'hc1b3328a, 32'h4268ba21};
test_output[5568:5575] = '{32'h4271f81c, 32'h0, 32'h425fd429, 32'h0, 32'h423fa44b, 32'h0, 32'h0, 32'h4268ba21};
test_input[5576:5583] = '{32'hc233a140, 32'hc1414201, 32'h418cbc30, 32'h42bc5be4, 32'h420ba480, 32'h4290b885, 32'h42bfd55f, 32'hc199a917};
test_output[5576:5583] = '{32'h0, 32'h0, 32'h418cbc30, 32'h42bc5be4, 32'h420ba480, 32'h4290b885, 32'h42bfd55f, 32'h0};
test_input[5584:5591] = '{32'h41f866ea, 32'h427ab6af, 32'hc21465b2, 32'hc21b638d, 32'h42827157, 32'hc2781bae, 32'h41a8fd2c, 32'h41e5d923};
test_output[5584:5591] = '{32'h41f866ea, 32'h427ab6af, 32'h0, 32'h0, 32'h42827157, 32'h0, 32'h41a8fd2c, 32'h41e5d923};
test_input[5592:5599] = '{32'h41609818, 32'h42962749, 32'hc29e4272, 32'hc26d13d7, 32'hc2a084ef, 32'h4299551a, 32'h4283a2d6, 32'h42630e40};
test_output[5592:5599] = '{32'h41609818, 32'h42962749, 32'h0, 32'h0, 32'h0, 32'h4299551a, 32'h4283a2d6, 32'h42630e40};
test_input[5600:5607] = '{32'hc25d7020, 32'hc29d9001, 32'hc16f0f90, 32'h4182e85b, 32'hc277ebb1, 32'hc21027f9, 32'h425afeee, 32'hc148affa};
test_output[5600:5607] = '{32'h0, 32'h0, 32'h0, 32'h4182e85b, 32'h0, 32'h0, 32'h425afeee, 32'h0};
test_input[5608:5615] = '{32'hc297709e, 32'h40e5a420, 32'h42876284, 32'h42905abc, 32'h42a17c3e, 32'h41b2dc04, 32'h429a3bda, 32'h42232975};
test_output[5608:5615] = '{32'h0, 32'h40e5a420, 32'h42876284, 32'h42905abc, 32'h42a17c3e, 32'h41b2dc04, 32'h429a3bda, 32'h42232975};
test_input[5616:5623] = '{32'h424e9efa, 32'h404e1371, 32'h427f31e2, 32'h424c787c, 32'hc2c39f5f, 32'h4189d4a6, 32'h41cbeb8a, 32'hc018f812};
test_output[5616:5623] = '{32'h424e9efa, 32'h404e1371, 32'h427f31e2, 32'h424c787c, 32'h0, 32'h4189d4a6, 32'h41cbeb8a, 32'h0};
test_input[5624:5631] = '{32'hc28b165a, 32'hc2433561, 32'hc1af5fa2, 32'h428371d9, 32'h422a2b18, 32'h42a40c54, 32'hc22fee8e, 32'hc1f8ed41};
test_output[5624:5631] = '{32'h0, 32'h0, 32'h0, 32'h428371d9, 32'h422a2b18, 32'h42a40c54, 32'h0, 32'h0};
test_input[5632:5639] = '{32'hc228a9d1, 32'h40b891b2, 32'h42a5e05b, 32'h42608256, 32'hbe1a1f16, 32'h41d6b034, 32'h420df820, 32'h419b1c3b};
test_output[5632:5639] = '{32'h0, 32'h40b891b2, 32'h42a5e05b, 32'h42608256, 32'h0, 32'h41d6b034, 32'h420df820, 32'h419b1c3b};
test_input[5640:5647] = '{32'hc2ad1963, 32'h429a039f, 32'h4228475c, 32'hc1f74a46, 32'hc28fc4d7, 32'h422c6bdb, 32'hc20db7ea, 32'h41a9c92a};
test_output[5640:5647] = '{32'h0, 32'h429a039f, 32'h4228475c, 32'h0, 32'h0, 32'h422c6bdb, 32'h0, 32'h41a9c92a};
test_input[5648:5655] = '{32'h429db4d3, 32'hc25a09e2, 32'hc1e0e0aa, 32'h41de770e, 32'hc1a97e90, 32'h421db11f, 32'h42573961, 32'h428b530e};
test_output[5648:5655] = '{32'h429db4d3, 32'h0, 32'h0, 32'h41de770e, 32'h0, 32'h421db11f, 32'h42573961, 32'h428b530e};
test_input[5656:5663] = '{32'h42c0d1a9, 32'hc2bd4a51, 32'h41414f0c, 32'h42366385, 32'h42c219ca, 32'h418dad44, 32'hc2c5751a, 32'h41a1c03d};
test_output[5656:5663] = '{32'h42c0d1a9, 32'h0, 32'h41414f0c, 32'h42366385, 32'h42c219ca, 32'h418dad44, 32'h0, 32'h41a1c03d};
test_input[5664:5671] = '{32'h412ed039, 32'h4180c43a, 32'h426fc069, 32'hc2b7cf4d, 32'hc19b35a8, 32'hc2588c97, 32'h421b9784, 32'hc2c5a149};
test_output[5664:5671] = '{32'h412ed039, 32'h4180c43a, 32'h426fc069, 32'h0, 32'h0, 32'h0, 32'h421b9784, 32'h0};
test_input[5672:5679] = '{32'h42165f94, 32'h42454abf, 32'hc135ec17, 32'h4267cf1e, 32'hc260fb67, 32'hc2099b27, 32'h40dd20c1, 32'hc1ae9f22};
test_output[5672:5679] = '{32'h42165f94, 32'h42454abf, 32'h0, 32'h4267cf1e, 32'h0, 32'h0, 32'h40dd20c1, 32'h0};
test_input[5680:5687] = '{32'h42a7dde7, 32'h42a1e603, 32'hc11773d5, 32'hc1b0c5e5, 32'h42a5cfe0, 32'h42b8124d, 32'h41e13253, 32'h41db5fc0};
test_output[5680:5687] = '{32'h42a7dde7, 32'h42a1e603, 32'h0, 32'h0, 32'h42a5cfe0, 32'h42b8124d, 32'h41e13253, 32'h41db5fc0};
test_input[5688:5695] = '{32'h41b31413, 32'hc235275f, 32'h41bd377f, 32'hc1b01f62, 32'h4104fa00, 32'hc02623d9, 32'hc2a954a6, 32'hc1be3d96};
test_output[5688:5695] = '{32'h41b31413, 32'h0, 32'h41bd377f, 32'h0, 32'h4104fa00, 32'h0, 32'h0, 32'h0};
test_input[5696:5703] = '{32'hc2ac409b, 32'hc2c50222, 32'hc2742763, 32'h429c05b8, 32'hc1e41385, 32'h42b203c0, 32'hc2c21653, 32'h4115366c};
test_output[5696:5703] = '{32'h0, 32'h0, 32'h0, 32'h429c05b8, 32'h0, 32'h42b203c0, 32'h0, 32'h4115366c};
test_input[5704:5711] = '{32'hc2a5180f, 32'hc044c8ac, 32'h4202ea64, 32'h41f111f5, 32'hc29f4611, 32'hc267e10d, 32'hc2b1c8f7, 32'hc2542567};
test_output[5704:5711] = '{32'h0, 32'h0, 32'h4202ea64, 32'h41f111f5, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5712:5719] = '{32'h4280a6df, 32'h42786190, 32'hc1c36d45, 32'h42ac0773, 32'hc23fce22, 32'hc2c1a831, 32'hc0603f81, 32'h428f3bf7};
test_output[5712:5719] = '{32'h4280a6df, 32'h42786190, 32'h0, 32'h42ac0773, 32'h0, 32'h0, 32'h0, 32'h428f3bf7};
test_input[5720:5727] = '{32'h42c55c91, 32'hc205e6d8, 32'h41ce7e35, 32'hc2a1cf65, 32'h42c4a93e, 32'h421b6fdb, 32'h429ab295, 32'h423f63f9};
test_output[5720:5727] = '{32'h42c55c91, 32'h0, 32'h41ce7e35, 32'h0, 32'h42c4a93e, 32'h421b6fdb, 32'h429ab295, 32'h423f63f9};
test_input[5728:5735] = '{32'h42355e4f, 32'hc2bf264d, 32'h41ea9bcc, 32'hc2b2498c, 32'hc12b7d96, 32'hc108df6b, 32'hc29fd9db, 32'hc296d4ae};
test_output[5728:5735] = '{32'h42355e4f, 32'h0, 32'h41ea9bcc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5736:5743] = '{32'hc260d28a, 32'hc2313777, 32'h419ccaa2, 32'h429ff784, 32'h41da6c00, 32'h42be1666, 32'h42bf3f2c, 32'hc263da7f};
test_output[5736:5743] = '{32'h0, 32'h0, 32'h419ccaa2, 32'h429ff784, 32'h41da6c00, 32'h42be1666, 32'h42bf3f2c, 32'h0};
test_input[5744:5751] = '{32'hc0f3b38b, 32'h42b3c5cc, 32'hc2473073, 32'hc2b628da, 32'hc27b39e8, 32'hc1e6e7e1, 32'hc29099ac, 32'h407d915b};
test_output[5744:5751] = '{32'h0, 32'h42b3c5cc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h407d915b};
test_input[5752:5759] = '{32'hc1f2eb31, 32'hc20d8b6f, 32'h427a341d, 32'h42ae1b05, 32'hc21aaff7, 32'h41caf232, 32'hc0604b77, 32'hc0185a1f};
test_output[5752:5759] = '{32'h0, 32'h0, 32'h427a341d, 32'h42ae1b05, 32'h0, 32'h41caf232, 32'h0, 32'h0};
test_input[5760:5767] = '{32'h42beffb3, 32'h3fc4f9c3, 32'hc28d1da7, 32'hc166dda4, 32'h4209a343, 32'hc10d2ff1, 32'hc1dec022, 32'h4194b73d};
test_output[5760:5767] = '{32'h42beffb3, 32'h3fc4f9c3, 32'h0, 32'h0, 32'h4209a343, 32'h0, 32'h0, 32'h4194b73d};
test_input[5768:5775] = '{32'hc2af76b7, 32'h4054d14b, 32'h408b27ba, 32'h42c3c03e, 32'hc141bab4, 32'h41babd94, 32'hc29a38d0, 32'hc2193d46};
test_output[5768:5775] = '{32'h0, 32'h4054d14b, 32'h408b27ba, 32'h42c3c03e, 32'h0, 32'h41babd94, 32'h0, 32'h0};
test_input[5776:5783] = '{32'hc22d13de, 32'hc2a2605e, 32'hc28f613c, 32'h3fe89fd9, 32'hc1a93676, 32'h41848531, 32'h428d940e, 32'hc1b73134};
test_output[5776:5783] = '{32'h0, 32'h0, 32'h0, 32'h3fe89fd9, 32'h0, 32'h41848531, 32'h428d940e, 32'h0};
test_input[5784:5791] = '{32'h412a8739, 32'hc2b08e40, 32'hc2acdcca, 32'h41f8004e, 32'h4276b1f8, 32'hc254198e, 32'hc29625e4, 32'h420ae9bc};
test_output[5784:5791] = '{32'h412a8739, 32'h0, 32'h0, 32'h41f8004e, 32'h4276b1f8, 32'h0, 32'h0, 32'h420ae9bc};
test_input[5792:5799] = '{32'hbdae87e9, 32'h40f863ce, 32'hc20f3b48, 32'h42b91cac, 32'hc282dad8, 32'hc23a5f24, 32'h426fd60c, 32'h4276d732};
test_output[5792:5799] = '{32'h0, 32'h40f863ce, 32'h0, 32'h42b91cac, 32'h0, 32'h0, 32'h426fd60c, 32'h4276d732};
test_input[5800:5807] = '{32'hc2996239, 32'hc283fe65, 32'h4234e4bc, 32'h42633b83, 32'h4265b219, 32'h41dc8021, 32'h41bd4483, 32'hc2b92595};
test_output[5800:5807] = '{32'h0, 32'h0, 32'h4234e4bc, 32'h42633b83, 32'h4265b219, 32'h41dc8021, 32'h41bd4483, 32'h0};
test_input[5808:5815] = '{32'h424d515c, 32'hc27a423e, 32'h41a9e50d, 32'hc2c2f55b, 32'hbfe5d3e8, 32'h41a18a24, 32'hc28ed70b, 32'h42b0d9a0};
test_output[5808:5815] = '{32'h424d515c, 32'h0, 32'h41a9e50d, 32'h0, 32'h0, 32'h41a18a24, 32'h0, 32'h42b0d9a0};
test_input[5816:5823] = '{32'hc2ae7715, 32'h42258a8f, 32'hc295bba5, 32'hc253f940, 32'h41e17504, 32'h40a93e5e, 32'h42c000fb, 32'h41af3a00};
test_output[5816:5823] = '{32'h0, 32'h42258a8f, 32'h0, 32'h0, 32'h41e17504, 32'h40a93e5e, 32'h42c000fb, 32'h41af3a00};
test_input[5824:5831] = '{32'hc2288cc9, 32'hc2b4d665, 32'hc2aa19b1, 32'hc131a615, 32'h42602a6f, 32'h42a168a1, 32'hc1d420ec, 32'hc20a50d1};
test_output[5824:5831] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42602a6f, 32'h42a168a1, 32'h0, 32'h0};
test_input[5832:5839] = '{32'hc276624c, 32'h42c561b9, 32'hc2be9731, 32'hc2977011, 32'hc2217863, 32'hc26d3044, 32'hc2c6a3a4, 32'hbf9d7fbe};
test_output[5832:5839] = '{32'h0, 32'h42c561b9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5840:5847] = '{32'h419ac5ae, 32'hbe8918a2, 32'h426cac96, 32'hc18555cf, 32'h4296e026, 32'hc25e5626, 32'h42219597, 32'hc12cb716};
test_output[5840:5847] = '{32'h419ac5ae, 32'h0, 32'h426cac96, 32'h0, 32'h4296e026, 32'h0, 32'h42219597, 32'h0};
test_input[5848:5855] = '{32'hc29b17dd, 32'hc1a282d5, 32'hc2a649b5, 32'h42425b5d, 32'hc2579052, 32'hc2c42075, 32'hc1871d33, 32'hc1233af8};
test_output[5848:5855] = '{32'h0, 32'h0, 32'h0, 32'h42425b5d, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5856:5863] = '{32'h42bbd933, 32'hc257409b, 32'h42a939e9, 32'h42931442, 32'hc245a47b, 32'h42442764, 32'hc2bb07fe, 32'h42ab8917};
test_output[5856:5863] = '{32'h42bbd933, 32'h0, 32'h42a939e9, 32'h42931442, 32'h0, 32'h42442764, 32'h0, 32'h42ab8917};
test_input[5864:5871] = '{32'hc29d5465, 32'hc120de8c, 32'hc1ea5c1e, 32'hc2457297, 32'h42422f2e, 32'h40efa243, 32'hc2848260, 32'hc23dbf1a};
test_output[5864:5871] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42422f2e, 32'h40efa243, 32'h0, 32'h0};
test_input[5872:5879] = '{32'hc2480144, 32'h42820d20, 32'h41e55bdb, 32'h42222699, 32'hc185ebc1, 32'hc2a71dc2, 32'hc24f209b, 32'hc2a4e79e};
test_output[5872:5879] = '{32'h0, 32'h42820d20, 32'h41e55bdb, 32'h42222699, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5880:5887] = '{32'hc20fcaf8, 32'hc19ba93a, 32'hc0e0444a, 32'hc28c570b, 32'hc2817458, 32'hc24edbd4, 32'h42a40a92, 32'hc090f305};
test_output[5880:5887] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a40a92, 32'h0};
test_input[5888:5895] = '{32'h41a431c6, 32'h4296f81d, 32'hc1ae46bc, 32'h4288cf06, 32'hc29abf12, 32'hc1f4e96c, 32'hc2414009, 32'h41ed8b4b};
test_output[5888:5895] = '{32'h41a431c6, 32'h4296f81d, 32'h0, 32'h4288cf06, 32'h0, 32'h0, 32'h0, 32'h41ed8b4b};
test_input[5896:5903] = '{32'h421da083, 32'hc1f07a1d, 32'hc147013d, 32'hc286f53f, 32'hc273a50d, 32'hc18d837b, 32'h41db8dbd, 32'hc1834b98};
test_output[5896:5903] = '{32'h421da083, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41db8dbd, 32'h0};
test_input[5904:5911] = '{32'h429a6388, 32'hc28fda34, 32'h426b2df2, 32'h41c61aee, 32'h4282f0ed, 32'hc256d872, 32'h42b3c9ab, 32'h425596e1};
test_output[5904:5911] = '{32'h429a6388, 32'h0, 32'h426b2df2, 32'h41c61aee, 32'h4282f0ed, 32'h0, 32'h42b3c9ab, 32'h425596e1};
test_input[5912:5919] = '{32'h3f9b5a9d, 32'hc21d7151, 32'h41a411cc, 32'h4210a494, 32'hc29f256b, 32'h424e7dea, 32'h414059b8, 32'hc24cadab};
test_output[5912:5919] = '{32'h3f9b5a9d, 32'h0, 32'h41a411cc, 32'h4210a494, 32'h0, 32'h424e7dea, 32'h414059b8, 32'h0};
test_input[5920:5927] = '{32'hc222f0f6, 32'hc1bf8826, 32'hc2abc8ab, 32'hc298c47f, 32'hc172c4c7, 32'hc268703a, 32'hc213efe2, 32'h4158ac90};
test_output[5920:5927] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4158ac90};
test_input[5928:5935] = '{32'hc24cd5b8, 32'h42139133, 32'h4256dc15, 32'h426b8919, 32'hc119ba59, 32'hc2a0c889, 32'hc2a57cac, 32'hc28f9986};
test_output[5928:5935] = '{32'h0, 32'h42139133, 32'h4256dc15, 32'h426b8919, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[5936:5943] = '{32'h3f746cb6, 32'h42165a31, 32'hc23f75d8, 32'h42b45b7d, 32'h42499726, 32'hc2bb650d, 32'h418c1937, 32'h428d6f17};
test_output[5936:5943] = '{32'h3f746cb6, 32'h42165a31, 32'h0, 32'h42b45b7d, 32'h42499726, 32'h0, 32'h418c1937, 32'h428d6f17};
test_input[5944:5951] = '{32'h422d935f, 32'h417f4365, 32'h41ac38fe, 32'h429c6c19, 32'h422f832c, 32'hc17d4ee9, 32'hc1081c0b, 32'hc19eeec1};
test_output[5944:5951] = '{32'h422d935f, 32'h417f4365, 32'h41ac38fe, 32'h429c6c19, 32'h422f832c, 32'h0, 32'h0, 32'h0};
test_input[5952:5959] = '{32'h423ed188, 32'hc2b9d3cf, 32'hc2646b8e, 32'hc29accc2, 32'h420b57c3, 32'h42a42528, 32'h4267d152, 32'h41bd6195};
test_output[5952:5959] = '{32'h423ed188, 32'h0, 32'h0, 32'h0, 32'h420b57c3, 32'h42a42528, 32'h4267d152, 32'h41bd6195};
test_input[5960:5967] = '{32'h4281ed45, 32'h4295357e, 32'hc299b711, 32'h405e004b, 32'hc2ac4005, 32'h40a637ea, 32'hc2a66b2e, 32'hc00d3b89};
test_output[5960:5967] = '{32'h4281ed45, 32'h4295357e, 32'h0, 32'h405e004b, 32'h0, 32'h40a637ea, 32'h0, 32'h0};
test_input[5968:5975] = '{32'hc2b89f61, 32'h4292d4d9, 32'h426aa80b, 32'hc2332ddb, 32'h41b5af89, 32'hc29e1325, 32'hc1b64cda, 32'h4232cb00};
test_output[5968:5975] = '{32'h0, 32'h4292d4d9, 32'h426aa80b, 32'h0, 32'h41b5af89, 32'h0, 32'h0, 32'h4232cb00};
test_input[5976:5983] = '{32'hc2bbba83, 32'h42a84b0a, 32'h42c54b58, 32'h42aa6a7b, 32'h42b5a04e, 32'h42bd4814, 32'h4205c39a, 32'h426b3542};
test_output[5976:5983] = '{32'h0, 32'h42a84b0a, 32'h42c54b58, 32'h42aa6a7b, 32'h42b5a04e, 32'h42bd4814, 32'h4205c39a, 32'h426b3542};
test_input[5984:5991] = '{32'hc0d46703, 32'h42994167, 32'h42bcc12b, 32'h424e6a3a, 32'hc2b4b400, 32'h4216440e, 32'hc25ec285, 32'hc2104ff6};
test_output[5984:5991] = '{32'h0, 32'h42994167, 32'h42bcc12b, 32'h424e6a3a, 32'h0, 32'h4216440e, 32'h0, 32'h0};
test_input[5992:5999] = '{32'h42b80a11, 32'h42b881fb, 32'h420a3db1, 32'h42948333, 32'hc1d5fb1d, 32'hc0d6868c, 32'hc01754b4, 32'hc19bfb63};
test_output[5992:5999] = '{32'h42b80a11, 32'h42b881fb, 32'h420a3db1, 32'h42948333, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6000:6007] = '{32'hc264ce65, 32'hc28adf4a, 32'hc19cb8f1, 32'h418da9ca, 32'h42a6b01a, 32'hc1def590, 32'h429b0787, 32'hc1349591};
test_output[6000:6007] = '{32'h0, 32'h0, 32'h0, 32'h418da9ca, 32'h42a6b01a, 32'h0, 32'h429b0787, 32'h0};
test_input[6008:6015] = '{32'h41de6883, 32'h428658cb, 32'h4130fb3a, 32'h42a7887f, 32'h42695c4c, 32'hc20ec019, 32'hc26dc63b, 32'h42bd395b};
test_output[6008:6015] = '{32'h41de6883, 32'h428658cb, 32'h4130fb3a, 32'h42a7887f, 32'h42695c4c, 32'h0, 32'h0, 32'h42bd395b};
test_input[6016:6023] = '{32'hc2b777c7, 32'hc1f98378, 32'hc2c60946, 32'h428f38f6, 32'hc26b690a, 32'hc2c2f79d, 32'hc28540be, 32'h41d0fb8b};
test_output[6016:6023] = '{32'h0, 32'h0, 32'h0, 32'h428f38f6, 32'h0, 32'h0, 32'h0, 32'h41d0fb8b};
test_input[6024:6031] = '{32'h42bbb8e6, 32'hc2b25a8e, 32'hc154b4b4, 32'h422e592b, 32'hc2637a66, 32'h400c6bb2, 32'h4026e7cd, 32'hc224380f};
test_output[6024:6031] = '{32'h42bbb8e6, 32'h0, 32'h0, 32'h422e592b, 32'h0, 32'h400c6bb2, 32'h4026e7cd, 32'h0};
test_input[6032:6039] = '{32'hc29570bb, 32'hc28aafea, 32'h4228e0e9, 32'h42a9900c, 32'h42085c0b, 32'hc1aee309, 32'h4282a693, 32'hc288fce8};
test_output[6032:6039] = '{32'h0, 32'h0, 32'h4228e0e9, 32'h42a9900c, 32'h42085c0b, 32'h0, 32'h4282a693, 32'h0};
test_input[6040:6047] = '{32'h426600a5, 32'hc29f94b3, 32'h42b138b4, 32'h429716e3, 32'hc2a32f19, 32'h422a0935, 32'h42226811, 32'hc13ebf7b};
test_output[6040:6047] = '{32'h426600a5, 32'h0, 32'h42b138b4, 32'h429716e3, 32'h0, 32'h422a0935, 32'h42226811, 32'h0};
test_input[6048:6055] = '{32'hc0aa58d7, 32'h42ad6851, 32'hc2b796c7, 32'hc29c0d1b, 32'hc24ddc0e, 32'h4233445e, 32'h42364d9a, 32'h42afc729};
test_output[6048:6055] = '{32'h0, 32'h42ad6851, 32'h0, 32'h0, 32'h0, 32'h4233445e, 32'h42364d9a, 32'h42afc729};
test_input[6056:6063] = '{32'hc28dab10, 32'h41e4bf6c, 32'h40a1854b, 32'hc28d9f9d, 32'hc171bbd3, 32'h42bdd9b8, 32'hc12a2ff8, 32'hc1d4f72e};
test_output[6056:6063] = '{32'h0, 32'h41e4bf6c, 32'h40a1854b, 32'h0, 32'h0, 32'h42bdd9b8, 32'h0, 32'h0};
test_input[6064:6071] = '{32'hc276c41f, 32'hbfd4c7d9, 32'hc2bab210, 32'hc20de3e7, 32'h4288191b, 32'h42186af9, 32'hc28672d0, 32'hc1db07b3};
test_output[6064:6071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4288191b, 32'h42186af9, 32'h0, 32'h0};
test_input[6072:6079] = '{32'hc12ee7cf, 32'hc1f73b40, 32'hc16960b7, 32'hc181e1fa, 32'hc1812304, 32'h422d8ee3, 32'hc246a1f7, 32'h4293f10c};
test_output[6072:6079] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422d8ee3, 32'h0, 32'h4293f10c};
test_input[6080:6087] = '{32'hc265c30d, 32'hc0487289, 32'hc2bf567d, 32'h4016e3a7, 32'hc279b0fd, 32'h4115f156, 32'h41b03cfb, 32'h422d7015};
test_output[6080:6087] = '{32'h0, 32'h0, 32'h0, 32'h4016e3a7, 32'h0, 32'h4115f156, 32'h41b03cfb, 32'h422d7015};
test_input[6088:6095] = '{32'hc20973d7, 32'h424c3144, 32'hc18441b1, 32'h4192f8da, 32'h4265bd52, 32'h428eed37, 32'h426d004a, 32'h4226cb8b};
test_output[6088:6095] = '{32'h0, 32'h424c3144, 32'h0, 32'h4192f8da, 32'h4265bd52, 32'h428eed37, 32'h426d004a, 32'h4226cb8b};
test_input[6096:6103] = '{32'hc2b85229, 32'hc2b311f7, 32'hc222de97, 32'h42c02d43, 32'h420c34a9, 32'h42639bec, 32'h428b414c, 32'hc1eb2ae0};
test_output[6096:6103] = '{32'h0, 32'h0, 32'h0, 32'h42c02d43, 32'h420c34a9, 32'h42639bec, 32'h428b414c, 32'h0};
test_input[6104:6111] = '{32'h42c132ef, 32'h4295a3c5, 32'hc1d70cbf, 32'hc297e044, 32'h4285cd21, 32'hc2201146, 32'hc1390a67, 32'hbfbe1632};
test_output[6104:6111] = '{32'h42c132ef, 32'h4295a3c5, 32'h0, 32'h0, 32'h4285cd21, 32'h0, 32'h0, 32'h0};
test_input[6112:6119] = '{32'hbf13a002, 32'hc229ccb7, 32'hc26c55bd, 32'h41b7395d, 32'hc2a6cb0a, 32'h420ed6dd, 32'h42bf6f33, 32'h4294554d};
test_output[6112:6119] = '{32'h0, 32'h0, 32'h0, 32'h41b7395d, 32'h0, 32'h420ed6dd, 32'h42bf6f33, 32'h4294554d};
test_input[6120:6127] = '{32'hc21e6a91, 32'h41da4bba, 32'h426f828c, 32'hc234e5fe, 32'hc15ddf92, 32'hc2b1e174, 32'hc29739de, 32'h42a3454f};
test_output[6120:6127] = '{32'h0, 32'h41da4bba, 32'h426f828c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a3454f};
test_input[6128:6135] = '{32'hc295ff72, 32'hc18f1969, 32'h4245e98f, 32'hc285870b, 32'h42c0613b, 32'hc24111c4, 32'h42a26a64, 32'h41fa858d};
test_output[6128:6135] = '{32'h0, 32'h0, 32'h4245e98f, 32'h0, 32'h42c0613b, 32'h0, 32'h42a26a64, 32'h41fa858d};
test_input[6136:6143] = '{32'h4236f6f9, 32'hc20c9b17, 32'h42bb02c1, 32'hc2bee6be, 32'h42a07d1f, 32'h4209e512, 32'hc28e7afd, 32'h4132ae25};
test_output[6136:6143] = '{32'h4236f6f9, 32'h0, 32'h42bb02c1, 32'h0, 32'h42a07d1f, 32'h4209e512, 32'h0, 32'h4132ae25};
test_input[6144:6151] = '{32'h4091f5f6, 32'h42aefd99, 32'h429a287f, 32'h420f6166, 32'hc01bdad5, 32'hc284c96c, 32'hc249efd1, 32'h4114a88b};
test_output[6144:6151] = '{32'h4091f5f6, 32'h42aefd99, 32'h429a287f, 32'h420f6166, 32'h0, 32'h0, 32'h0, 32'h4114a88b};
test_input[6152:6159] = '{32'h42485d35, 32'h42624402, 32'hc2a979bf, 32'hc23453ab, 32'h429d2e27, 32'h41c3dfc5, 32'hc0ea59f5, 32'h42b5d648};
test_output[6152:6159] = '{32'h42485d35, 32'h42624402, 32'h0, 32'h0, 32'h429d2e27, 32'h41c3dfc5, 32'h0, 32'h42b5d648};
test_input[6160:6167] = '{32'h41af7664, 32'h411a1232, 32'hc2ac934c, 32'hc251f310, 32'h42777136, 32'h42ae04cb, 32'hc2340d4a, 32'h427e2936};
test_output[6160:6167] = '{32'h41af7664, 32'h411a1232, 32'h0, 32'h0, 32'h42777136, 32'h42ae04cb, 32'h0, 32'h427e2936};
test_input[6168:6175] = '{32'hc2278e08, 32'h429781f1, 32'hc2a746f6, 32'hc1cd13da, 32'h4218cd26, 32'h429abf7a, 32'hbec200a2, 32'hc2598129};
test_output[6168:6175] = '{32'h0, 32'h429781f1, 32'h0, 32'h0, 32'h4218cd26, 32'h429abf7a, 32'h0, 32'h0};
test_input[6176:6183] = '{32'h412a8245, 32'hc2480766, 32'hc2c0ed23, 32'hc1de24c2, 32'hc1624a6a, 32'hc256688f, 32'hc2829674, 32'h42ad4d47};
test_output[6176:6183] = '{32'h412a8245, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ad4d47};
test_input[6184:6191] = '{32'h41368d36, 32'h4040c364, 32'hc2680490, 32'h4296d127, 32'h42b7f3f5, 32'hc2b60ffa, 32'h42a33b5d, 32'h4180f596};
test_output[6184:6191] = '{32'h41368d36, 32'h4040c364, 32'h0, 32'h4296d127, 32'h42b7f3f5, 32'h0, 32'h42a33b5d, 32'h4180f596};
test_input[6192:6199] = '{32'h42c355d2, 32'hc2bb94c8, 32'hc293ba36, 32'hc128ed2f, 32'hc21b4849, 32'h429166bb, 32'hc221094e, 32'hc2b73e63};
test_output[6192:6199] = '{32'h42c355d2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429166bb, 32'h0, 32'h0};
test_input[6200:6207] = '{32'hc2b3cb38, 32'hc281dec9, 32'h426ed669, 32'h42802f47, 32'hc275f243, 32'hc2a26346, 32'h420b3313, 32'hc1cfe78c};
test_output[6200:6207] = '{32'h0, 32'h0, 32'h426ed669, 32'h42802f47, 32'h0, 32'h0, 32'h420b3313, 32'h0};
test_input[6208:6215] = '{32'hc29d9b27, 32'h42251d69, 32'hc2b9b196, 32'h42465b52, 32'hc27e7576, 32'h4249d2f4, 32'h41cca67c, 32'hc2556440};
test_output[6208:6215] = '{32'h0, 32'h42251d69, 32'h0, 32'h42465b52, 32'h0, 32'h4249d2f4, 32'h41cca67c, 32'h0};
test_input[6216:6223] = '{32'h4203813a, 32'h4257658f, 32'h419b1fc0, 32'h4202aab8, 32'hc16cb302, 32'hc242e570, 32'hc09ae3ca, 32'hc2793699};
test_output[6216:6223] = '{32'h4203813a, 32'h4257658f, 32'h419b1fc0, 32'h4202aab8, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6224:6231] = '{32'hc2c40b90, 32'hc25e3886, 32'hc22fc00d, 32'hc0adfa0e, 32'hc1f79499, 32'hc2c2d3d7, 32'h42bd20ae, 32'h42b0b753};
test_output[6224:6231] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bd20ae, 32'h42b0b753};
test_input[6232:6239] = '{32'hc2a7b0f4, 32'h40fb668e, 32'hc2180605, 32'h41613d5a, 32'hc29d2787, 32'hc2bd8e21, 32'hc2a284fe, 32'hc29c0b9f};
test_output[6232:6239] = '{32'h0, 32'h40fb668e, 32'h0, 32'h41613d5a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6240:6247] = '{32'h41a1eddd, 32'hc2bd5bd3, 32'h4248cef0, 32'hc29b1cf7, 32'hc2c022aa, 32'h424c8637, 32'hc1c5a29f, 32'h42b88770};
test_output[6240:6247] = '{32'h41a1eddd, 32'h0, 32'h4248cef0, 32'h0, 32'h0, 32'h424c8637, 32'h0, 32'h42b88770};
test_input[6248:6255] = '{32'hc07225ee, 32'hc23d15c3, 32'hc29af294, 32'h42346838, 32'hc25db093, 32'h40242c32, 32'hc1ff3c33, 32'hc2900342};
test_output[6248:6255] = '{32'h0, 32'h0, 32'h0, 32'h42346838, 32'h0, 32'h40242c32, 32'h0, 32'h0};
test_input[6256:6263] = '{32'hc2b84471, 32'h41ff63c9, 32'h41859d91, 32'h41064f6d, 32'h428d00ce, 32'h40f6f32a, 32'h42957970, 32'h42965974};
test_output[6256:6263] = '{32'h0, 32'h41ff63c9, 32'h41859d91, 32'h41064f6d, 32'h428d00ce, 32'h40f6f32a, 32'h42957970, 32'h42965974};
test_input[6264:6271] = '{32'hc2191b08, 32'h424810b7, 32'h4222aac4, 32'h42b85d8e, 32'h42aa9806, 32'hc1c9ea03, 32'h428d9b86, 32'h42a7962a};
test_output[6264:6271] = '{32'h0, 32'h424810b7, 32'h4222aac4, 32'h42b85d8e, 32'h42aa9806, 32'h0, 32'h428d9b86, 32'h42a7962a};
test_input[6272:6279] = '{32'hc2bc1adb, 32'h420d8148, 32'h416e29f5, 32'h4157d80a, 32'h41c5ed35, 32'hc04c2cc1, 32'h4265be6f, 32'h41c5d901};
test_output[6272:6279] = '{32'h0, 32'h420d8148, 32'h416e29f5, 32'h4157d80a, 32'h41c5ed35, 32'h0, 32'h4265be6f, 32'h41c5d901};
test_input[6280:6287] = '{32'h422eb7ca, 32'h4266bad1, 32'h41280a1e, 32'h41a256d8, 32'hc2c203ab, 32'hc220127d, 32'hc0fdca9b, 32'h4211e457};
test_output[6280:6287] = '{32'h422eb7ca, 32'h4266bad1, 32'h41280a1e, 32'h41a256d8, 32'h0, 32'h0, 32'h0, 32'h4211e457};
test_input[6288:6295] = '{32'h412aaeb8, 32'h3f01a53c, 32'hc2790372, 32'hc14f908a, 32'hc2c6242e, 32'h41e45496, 32'hc02ca50a, 32'hc159e53d};
test_output[6288:6295] = '{32'h412aaeb8, 32'h3f01a53c, 32'h0, 32'h0, 32'h0, 32'h41e45496, 32'h0, 32'h0};
test_input[6296:6303] = '{32'hc1322072, 32'h422f6b4e, 32'hc265fe2d, 32'hc2b125a8, 32'hc1f19909, 32'hc2733e92, 32'h4295485a, 32'h427fb499};
test_output[6296:6303] = '{32'h0, 32'h422f6b4e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4295485a, 32'h427fb499};
test_input[6304:6311] = '{32'hc2a9f28c, 32'h41bd9c68, 32'hc27ed4d6, 32'h4217c116, 32'h41071c39, 32'h4270a668, 32'hc1a52d35, 32'h429fb9b9};
test_output[6304:6311] = '{32'h0, 32'h41bd9c68, 32'h0, 32'h4217c116, 32'h41071c39, 32'h4270a668, 32'h0, 32'h429fb9b9};
test_input[6312:6319] = '{32'hc21be500, 32'h42b32f68, 32'h413459ff, 32'hc2792c62, 32'hc2a58bff, 32'h4200d30e, 32'hc2bf4d7b, 32'h41888e02};
test_output[6312:6319] = '{32'h0, 32'h42b32f68, 32'h413459ff, 32'h0, 32'h0, 32'h4200d30e, 32'h0, 32'h41888e02};
test_input[6320:6327] = '{32'hc297a47e, 32'h3f913b99, 32'hc2c50171, 32'hc29813bd, 32'h42b86e06, 32'hc206e15a, 32'hc25a1b2f, 32'hc21f75aa};
test_output[6320:6327] = '{32'h0, 32'h3f913b99, 32'h0, 32'h0, 32'h42b86e06, 32'h0, 32'h0, 32'h0};
test_input[6328:6335] = '{32'h4275586c, 32'h41902510, 32'h41c98651, 32'h4219c906, 32'h4287f295, 32'hc2b86718, 32'hc267fe95, 32'h41fa6dc5};
test_output[6328:6335] = '{32'h4275586c, 32'h41902510, 32'h41c98651, 32'h4219c906, 32'h4287f295, 32'h0, 32'h0, 32'h41fa6dc5};
test_input[6336:6343] = '{32'hc1f79005, 32'h42b5b2d1, 32'hc2232fe9, 32'h42437cfd, 32'hc2b81555, 32'hc28d8d62, 32'h428b9428, 32'h41c519f3};
test_output[6336:6343] = '{32'h0, 32'h42b5b2d1, 32'h0, 32'h42437cfd, 32'h0, 32'h0, 32'h428b9428, 32'h41c519f3};
test_input[6344:6351] = '{32'hc22e3e87, 32'hc1da589a, 32'hc1e0f4f0, 32'h41a54bb6, 32'h42178677, 32'h42bfb42e, 32'hc279e3f6, 32'h417d8479};
test_output[6344:6351] = '{32'h0, 32'h0, 32'h0, 32'h41a54bb6, 32'h42178677, 32'h42bfb42e, 32'h0, 32'h417d8479};
test_input[6352:6359] = '{32'hc268d771, 32'h4287b989, 32'h4213ee76, 32'hc284655c, 32'hc2602bf3, 32'h3c5b32ba, 32'hc254108a, 32'h4245b04c};
test_output[6352:6359] = '{32'h0, 32'h4287b989, 32'h4213ee76, 32'h0, 32'h0, 32'h3c5b32ba, 32'h0, 32'h4245b04c};
test_input[6360:6367] = '{32'hc201dd01, 32'hc1df6987, 32'h418618e8, 32'hc2bff785, 32'hc0075c51, 32'h426cbd58, 32'hc2accde5, 32'hc2abccd5};
test_output[6360:6367] = '{32'h0, 32'h0, 32'h418618e8, 32'h0, 32'h0, 32'h426cbd58, 32'h0, 32'h0};
test_input[6368:6375] = '{32'h423d644d, 32'h4211b88a, 32'h40e474b1, 32'hc28b8e2d, 32'h424d4357, 32'h413c0c6f, 32'hc24a3ef1, 32'hc0b7ce18};
test_output[6368:6375] = '{32'h423d644d, 32'h4211b88a, 32'h40e474b1, 32'h0, 32'h424d4357, 32'h413c0c6f, 32'h0, 32'h0};
test_input[6376:6383] = '{32'h4091cb91, 32'hc16e9c6e, 32'hc2338d04, 32'hc2878a7b, 32'h41f23530, 32'h42c6a39f, 32'hc192c869, 32'h40816f44};
test_output[6376:6383] = '{32'h4091cb91, 32'h0, 32'h0, 32'h0, 32'h41f23530, 32'h42c6a39f, 32'h0, 32'h40816f44};
test_input[6384:6391] = '{32'h429a4c1a, 32'hc289ef94, 32'hc2965c56, 32'hc2749773, 32'h426f212d, 32'h429e0735, 32'hc23b00fb, 32'hc1bd52bf};
test_output[6384:6391] = '{32'h429a4c1a, 32'h0, 32'h0, 32'h0, 32'h426f212d, 32'h429e0735, 32'h0, 32'h0};
test_input[6392:6399] = '{32'hc22f443b, 32'h429c135b, 32'hc1a9716d, 32'h428ba47a, 32'h4174c918, 32'hc2aac94d, 32'h428a6a2d, 32'hc2a29ce7};
test_output[6392:6399] = '{32'h0, 32'h429c135b, 32'h0, 32'h428ba47a, 32'h4174c918, 32'h0, 32'h428a6a2d, 32'h0};
test_input[6400:6407] = '{32'hc13b2745, 32'h41602edc, 32'hc2c63e2c, 32'hc2bf5933, 32'h427542b9, 32'hc14340d5, 32'hc2ab8518, 32'hc28b46a3};
test_output[6400:6407] = '{32'h0, 32'h41602edc, 32'h0, 32'h0, 32'h427542b9, 32'h0, 32'h0, 32'h0};
test_input[6408:6415] = '{32'h42742e8b, 32'h42b27430, 32'hc1c2824a, 32'h42a71f25, 32'h416daf5a, 32'h423c9f98, 32'hc2079c1e, 32'hc2458b77};
test_output[6408:6415] = '{32'h42742e8b, 32'h42b27430, 32'h0, 32'h42a71f25, 32'h416daf5a, 32'h423c9f98, 32'h0, 32'h0};
test_input[6416:6423] = '{32'h426c8da3, 32'h41569ef6, 32'h420fef42, 32'h4267dab1, 32'h400f6884, 32'h42041aae, 32'h427d1b59, 32'h42611159};
test_output[6416:6423] = '{32'h426c8da3, 32'h41569ef6, 32'h420fef42, 32'h4267dab1, 32'h400f6884, 32'h42041aae, 32'h427d1b59, 32'h42611159};
test_input[6424:6431] = '{32'hc2b9cb16, 32'h42a32e6e, 32'h424d9122, 32'h42a2464f, 32'h42beebd5, 32'hc26ec057, 32'hc1094d49, 32'h42998b0b};
test_output[6424:6431] = '{32'h0, 32'h42a32e6e, 32'h424d9122, 32'h42a2464f, 32'h42beebd5, 32'h0, 32'h0, 32'h42998b0b};
test_input[6432:6439] = '{32'hc2a4baa2, 32'hc1b4d688, 32'h424a1e40, 32'hc22a0c0a, 32'h42474eac, 32'h41bdae0f, 32'h42b0aa73, 32'h42307874};
test_output[6432:6439] = '{32'h0, 32'h0, 32'h424a1e40, 32'h0, 32'h42474eac, 32'h41bdae0f, 32'h42b0aa73, 32'h42307874};
test_input[6440:6447] = '{32'h424604cb, 32'h42a2d917, 32'hc20ddd80, 32'h412de628, 32'h42c36b71, 32'h42143c79, 32'hc017da43, 32'hc20f2b24};
test_output[6440:6447] = '{32'h424604cb, 32'h42a2d917, 32'h0, 32'h412de628, 32'h42c36b71, 32'h42143c79, 32'h0, 32'h0};
test_input[6448:6455] = '{32'hc2acc86d, 32'h42a08669, 32'hc281a50f, 32'hc294c525, 32'hc2a3a95b, 32'h4124ff8d, 32'h4216b256, 32'hc22b2cfe};
test_output[6448:6455] = '{32'h0, 32'h42a08669, 32'h0, 32'h0, 32'h0, 32'h4124ff8d, 32'h4216b256, 32'h0};
test_input[6456:6463] = '{32'h40dacecf, 32'hc28b554a, 32'hc2b9d748, 32'h411daba4, 32'hc290ab7c, 32'hc2b5b632, 32'hc2c1fbe2, 32'h429ef4f2};
test_output[6456:6463] = '{32'h40dacecf, 32'h0, 32'h0, 32'h411daba4, 32'h0, 32'h0, 32'h0, 32'h429ef4f2};
test_input[6464:6471] = '{32'h42675fcd, 32'h4263edc7, 32'hc0877bbc, 32'h4274e2e6, 32'h41f099e6, 32'h42638731, 32'hc1913f54, 32'h422f3d4e};
test_output[6464:6471] = '{32'h42675fcd, 32'h4263edc7, 32'h0, 32'h4274e2e6, 32'h41f099e6, 32'h42638731, 32'h0, 32'h422f3d4e};
test_input[6472:6479] = '{32'h4294f55a, 32'hc2a9b654, 32'hc2c4412e, 32'h4218cfd3, 32'h42a047dd, 32'h4288a72d, 32'hc2948318, 32'h40f28242};
test_output[6472:6479] = '{32'h4294f55a, 32'h0, 32'h0, 32'h4218cfd3, 32'h42a047dd, 32'h4288a72d, 32'h0, 32'h40f28242};
test_input[6480:6487] = '{32'hc238f364, 32'hc2817884, 32'hc2b81ff6, 32'hc29234ed, 32'hc29d012c, 32'h426b7b1f, 32'hc23fe678, 32'h42942757};
test_output[6480:6487] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426b7b1f, 32'h0, 32'h42942757};
test_input[6488:6495] = '{32'h42b44b92, 32'hc2087802, 32'h428cae8c, 32'hc180f482, 32'h41d61c2d, 32'h41c50273, 32'h41796b4a, 32'h421999af};
test_output[6488:6495] = '{32'h42b44b92, 32'h0, 32'h428cae8c, 32'h0, 32'h41d61c2d, 32'h41c50273, 32'h41796b4a, 32'h421999af};
test_input[6496:6503] = '{32'h41a7cc95, 32'hc14d27e3, 32'h42818286, 32'hc2a02a41, 32'hc29691e8, 32'hc29473fc, 32'hc1cd7f91, 32'h4280a109};
test_output[6496:6503] = '{32'h41a7cc95, 32'h0, 32'h42818286, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4280a109};
test_input[6504:6511] = '{32'h42bebff5, 32'hc1d593ca, 32'hc02a4d6f, 32'h42b53ccd, 32'hc206f28f, 32'hc2adadc4, 32'hc0bb35ba, 32'hc2170a6d};
test_output[6504:6511] = '{32'h42bebff5, 32'h0, 32'h0, 32'h42b53ccd, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6512:6519] = '{32'h42494bbf, 32'hc2b6a988, 32'h40a4b307, 32'hc18184c9, 32'hc113c661, 32'h42755197, 32'hc0120528, 32'hc0a6a152};
test_output[6512:6519] = '{32'h42494bbf, 32'h0, 32'h40a4b307, 32'h0, 32'h0, 32'h42755197, 32'h0, 32'h0};
test_input[6520:6527] = '{32'h41c9c1e7, 32'h3f6a5a20, 32'h4169e22b, 32'hc2c49cce, 32'h40a5f03c, 32'hc191cc95, 32'hc273930f, 32'hc24c9964};
test_output[6520:6527] = '{32'h41c9c1e7, 32'h3f6a5a20, 32'h4169e22b, 32'h0, 32'h40a5f03c, 32'h0, 32'h0, 32'h0};
test_input[6528:6535] = '{32'h42c20011, 32'hc11f740c, 32'hc0f4bf68, 32'h420f0534, 32'hc2c7aa33, 32'h422d4e8a, 32'h42be91da, 32'h42bcb5fb};
test_output[6528:6535] = '{32'h42c20011, 32'h0, 32'h0, 32'h420f0534, 32'h0, 32'h422d4e8a, 32'h42be91da, 32'h42bcb5fb};
test_input[6536:6543] = '{32'hc2a8a58d, 32'h42429ff7, 32'hc18cd30d, 32'hc24b287d, 32'hc29baae0, 32'h425cfcaa, 32'h4277c305, 32'h4290152a};
test_output[6536:6543] = '{32'h0, 32'h42429ff7, 32'h0, 32'h0, 32'h0, 32'h425cfcaa, 32'h4277c305, 32'h4290152a};
test_input[6544:6551] = '{32'h41c1e395, 32'hc2a712a8, 32'h423ebf1a, 32'h422bc676, 32'h4291a64a, 32'h425a2252, 32'hc2b6688e, 32'hc0650226};
test_output[6544:6551] = '{32'h41c1e395, 32'h0, 32'h423ebf1a, 32'h422bc676, 32'h4291a64a, 32'h425a2252, 32'h0, 32'h0};
test_input[6552:6559] = '{32'h42834ee4, 32'h419e639f, 32'h40c02725, 32'h427eb696, 32'hc2a57951, 32'hc13a3b94, 32'hc1cf6726, 32'hc222a754};
test_output[6552:6559] = '{32'h42834ee4, 32'h419e639f, 32'h40c02725, 32'h427eb696, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6560:6567] = '{32'hc20eff77, 32'h426d544e, 32'h416b6bc6, 32'h42c62096, 32'h3f0942ed, 32'hc2153b5d, 32'h415416fb, 32'hc173fd51};
test_output[6560:6567] = '{32'h0, 32'h426d544e, 32'h416b6bc6, 32'h42c62096, 32'h3f0942ed, 32'h0, 32'h415416fb, 32'h0};
test_input[6568:6575] = '{32'hc1a58df9, 32'h428190d2, 32'hc233fcde, 32'hc15aa017, 32'hc26178f1, 32'hc22554af, 32'hc28f9579, 32'hc2a229cd};
test_output[6568:6575] = '{32'h0, 32'h428190d2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6576:6583] = '{32'hc20a356a, 32'h41eaef6b, 32'hc2c47543, 32'hc2395f9c, 32'hc1bb740f, 32'hc2a332be, 32'h41aaa4f4, 32'h420e584d};
test_output[6576:6583] = '{32'h0, 32'h41eaef6b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41aaa4f4, 32'h420e584d};
test_input[6584:6591] = '{32'h412ee041, 32'hc21f9264, 32'hc1cd4c9b, 32'hc24f612b, 32'hc209a92f, 32'hc27e8850, 32'h425e2d2c, 32'h42bf9a0c};
test_output[6584:6591] = '{32'h412ee041, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425e2d2c, 32'h42bf9a0c};
test_input[6592:6599] = '{32'h4225ee39, 32'h4212087d, 32'hc2acd4b2, 32'hc2907230, 32'hc2b0a9c3, 32'h4218bc0c, 32'hc293e0e6, 32'hc2c33c21};
test_output[6592:6599] = '{32'h4225ee39, 32'h4212087d, 32'h0, 32'h0, 32'h0, 32'h4218bc0c, 32'h0, 32'h0};
test_input[6600:6607] = '{32'hbe61af6a, 32'h421a16f7, 32'hc2b99c99, 32'h412bb593, 32'h4259ff93, 32'hc15ab691, 32'h429151a1, 32'h4246d938};
test_output[6600:6607] = '{32'h0, 32'h421a16f7, 32'h0, 32'h412bb593, 32'h4259ff93, 32'h0, 32'h429151a1, 32'h4246d938};
test_input[6608:6615] = '{32'hc243856b, 32'h4236ae7e, 32'hc2c24b8d, 32'hc0d0065e, 32'hc2ab3ad1, 32'h423d5cfe, 32'hc2bc249f, 32'h4213a5a2};
test_output[6608:6615] = '{32'h0, 32'h4236ae7e, 32'h0, 32'h0, 32'h0, 32'h423d5cfe, 32'h0, 32'h4213a5a2};
test_input[6616:6623] = '{32'h40be46e0, 32'h41b0aa24, 32'hc21f4f7b, 32'hc29c8427, 32'h4111903c, 32'h4190346e, 32'h420f8da1, 32'hc29212d5};
test_output[6616:6623] = '{32'h40be46e0, 32'h41b0aa24, 32'h0, 32'h0, 32'h4111903c, 32'h4190346e, 32'h420f8da1, 32'h0};
test_input[6624:6631] = '{32'hc27351ba, 32'h42adad3c, 32'hc2c4ce7e, 32'hbf10e76a, 32'h424a5ba1, 32'hc1e81aef, 32'h42ac1557, 32'hc213a98a};
test_output[6624:6631] = '{32'h0, 32'h42adad3c, 32'h0, 32'h0, 32'h424a5ba1, 32'h0, 32'h42ac1557, 32'h0};
test_input[6632:6639] = '{32'h429dd5ef, 32'h423d1dcc, 32'hc26e1d35, 32'hc294e9c4, 32'h42c61197, 32'h42bf4bd6, 32'h425cf32c, 32'h417ed0e8};
test_output[6632:6639] = '{32'h429dd5ef, 32'h423d1dcc, 32'h0, 32'h0, 32'h42c61197, 32'h42bf4bd6, 32'h425cf32c, 32'h417ed0e8};
test_input[6640:6647] = '{32'hc26c9597, 32'hc238267f, 32'hc18525db, 32'hc2c00821, 32'h42c11cd3, 32'h41b6cf75, 32'hc20792b5, 32'hc29ce34e};
test_output[6640:6647] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42c11cd3, 32'h41b6cf75, 32'h0, 32'h0};
test_input[6648:6655] = '{32'hc20a0207, 32'h42685379, 32'hc295f95c, 32'h410edef5, 32'h426569c1, 32'h420c728d, 32'hc2c76f99, 32'hc26ae957};
test_output[6648:6655] = '{32'h0, 32'h42685379, 32'h0, 32'h410edef5, 32'h426569c1, 32'h420c728d, 32'h0, 32'h0};
test_input[6656:6663] = '{32'h42aa9c3f, 32'hc2b3d610, 32'h423df5d5, 32'hbfcb9e77, 32'hc2c08499, 32'h41226d0f, 32'h42c2bb0c, 32'hc19889cb};
test_output[6656:6663] = '{32'h42aa9c3f, 32'h0, 32'h423df5d5, 32'h0, 32'h0, 32'h41226d0f, 32'h42c2bb0c, 32'h0};
test_input[6664:6671] = '{32'h41d24c9c, 32'hc2a12ee9, 32'h425ddd92, 32'h41a8647e, 32'h429946ce, 32'h3fda756b, 32'hc2870b58, 32'hc1db605a};
test_output[6664:6671] = '{32'h41d24c9c, 32'h0, 32'h425ddd92, 32'h41a8647e, 32'h429946ce, 32'h3fda756b, 32'h0, 32'h0};
test_input[6672:6679] = '{32'h429ab1f5, 32'hc20f9ce8, 32'hc2c255cf, 32'hc1e73992, 32'h41ea8bd1, 32'hc23fb9bd, 32'h42474384, 32'hc1c3581e};
test_output[6672:6679] = '{32'h429ab1f5, 32'h0, 32'h0, 32'h0, 32'h41ea8bd1, 32'h0, 32'h42474384, 32'h0};
test_input[6680:6687] = '{32'hc2b0de2c, 32'h3f5e94f9, 32'h4255888a, 32'hc1dde352, 32'h41157db1, 32'hc28d2b3c, 32'h42be8cd2, 32'h40adae87};
test_output[6680:6687] = '{32'h0, 32'h3f5e94f9, 32'h4255888a, 32'h0, 32'h41157db1, 32'h0, 32'h42be8cd2, 32'h40adae87};
test_input[6688:6695] = '{32'h429d61cd, 32'h4122c186, 32'h410ee74f, 32'h42bb1ab0, 32'hc24ed02d, 32'hc2c1ff1b, 32'hc16c81c0, 32'h40f02f60};
test_output[6688:6695] = '{32'h429d61cd, 32'h4122c186, 32'h410ee74f, 32'h42bb1ab0, 32'h0, 32'h0, 32'h0, 32'h40f02f60};
test_input[6696:6703] = '{32'h427b06ce, 32'h42b8a1ac, 32'hc2a20389, 32'hc2c0ff63, 32'hc25b76ee, 32'h42af499e, 32'h425579e5, 32'h423446e4};
test_output[6696:6703] = '{32'h427b06ce, 32'h42b8a1ac, 32'h0, 32'h0, 32'h0, 32'h42af499e, 32'h425579e5, 32'h423446e4};
test_input[6704:6711] = '{32'hc1664706, 32'hc11ff1f4, 32'hc193d186, 32'h428b0a7b, 32'h42060ede, 32'hc298205f, 32'h41826110, 32'h4215ca58};
test_output[6704:6711] = '{32'h0, 32'h0, 32'h0, 32'h428b0a7b, 32'h42060ede, 32'h0, 32'h41826110, 32'h4215ca58};
test_input[6712:6719] = '{32'hc1916f5f, 32'hc26be206, 32'hc29d51df, 32'h429e0916, 32'hc1002ad5, 32'h42a10ea7, 32'hc2c0d961, 32'h42abd7ed};
test_output[6712:6719] = '{32'h0, 32'h0, 32'h0, 32'h429e0916, 32'h0, 32'h42a10ea7, 32'h0, 32'h42abd7ed};
test_input[6720:6727] = '{32'hc2b94110, 32'hc2a63bc2, 32'hc2212752, 32'hc2343336, 32'hc1238879, 32'hc22f3d2d, 32'h40062180, 32'h41eea356};
test_output[6720:6727] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40062180, 32'h41eea356};
test_input[6728:6735] = '{32'h42ae18ac, 32'hc207ca8e, 32'h42169cba, 32'h421991b1, 32'hc248ed62, 32'hc2502906, 32'h424ddfce, 32'h42587e6b};
test_output[6728:6735] = '{32'h42ae18ac, 32'h0, 32'h42169cba, 32'h421991b1, 32'h0, 32'h0, 32'h424ddfce, 32'h42587e6b};
test_input[6736:6743] = '{32'hc1f1d0db, 32'h412358b9, 32'hc095cc06, 32'hc19f5bda, 32'h41717045, 32'hc1c0bab8, 32'h4097b9a4, 32'hc2a49296};
test_output[6736:6743] = '{32'h0, 32'h412358b9, 32'h0, 32'h0, 32'h41717045, 32'h0, 32'h4097b9a4, 32'h0};
test_input[6744:6751] = '{32'hc23bd3c6, 32'h423ce251, 32'h419575c6, 32'hc28c3e8e, 32'h42a65256, 32'hc22580a5, 32'hc1964598, 32'hc28b84be};
test_output[6744:6751] = '{32'h0, 32'h423ce251, 32'h419575c6, 32'h0, 32'h42a65256, 32'h0, 32'h0, 32'h0};
test_input[6752:6759] = '{32'hc28a3f6e, 32'hc273853c, 32'h41e42da8, 32'hc28b9a8b, 32'h41febc67, 32'h419f0cc6, 32'h428cf82c, 32'h4192ea0a};
test_output[6752:6759] = '{32'h0, 32'h0, 32'h41e42da8, 32'h0, 32'h41febc67, 32'h419f0cc6, 32'h428cf82c, 32'h4192ea0a};
test_input[6760:6767] = '{32'hc1ab4ce3, 32'hc1c74b05, 32'hbfc579bb, 32'h41990a85, 32'h40b33235, 32'hc26af2b5, 32'h42bca8db, 32'hc282f108};
test_output[6760:6767] = '{32'h0, 32'h0, 32'h0, 32'h41990a85, 32'h40b33235, 32'h0, 32'h42bca8db, 32'h0};
test_input[6768:6775] = '{32'h42294f24, 32'hc2408b5d, 32'hc185833e, 32'h42a7e987, 32'h42a5f6a6, 32'h42b09f0d, 32'h42023274, 32'h42906f25};
test_output[6768:6775] = '{32'h42294f24, 32'h0, 32'h0, 32'h42a7e987, 32'h42a5f6a6, 32'h42b09f0d, 32'h42023274, 32'h42906f25};
test_input[6776:6783] = '{32'hc2c2a32a, 32'h41dabf19, 32'hc269c2be, 32'hc231ceda, 32'hc1cdc80a, 32'h42761fca, 32'hc0f4f2c1, 32'hc234febc};
test_output[6776:6783] = '{32'h0, 32'h41dabf19, 32'h0, 32'h0, 32'h0, 32'h42761fca, 32'h0, 32'h0};
test_input[6784:6791] = '{32'hc2a54064, 32'hc2ab9e9b, 32'hc2bb3996, 32'h3ee19a7f, 32'hc24f62d8, 32'hc2767ec3, 32'hc2af61ac, 32'hc2ad0ad8};
test_output[6784:6791] = '{32'h0, 32'h0, 32'h0, 32'h3ee19a7f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6792:6799] = '{32'h4294bc31, 32'h42c358c5, 32'hc293cfb3, 32'hc29aa597, 32'h42074ca5, 32'h420e5099, 32'h42a5f19c, 32'h42a3e29b};
test_output[6792:6799] = '{32'h4294bc31, 32'h42c358c5, 32'h0, 32'h0, 32'h42074ca5, 32'h420e5099, 32'h42a5f19c, 32'h42a3e29b};
test_input[6800:6807] = '{32'hc227e180, 32'h426f77bd, 32'hc02471e3, 32'hc1e982e9, 32'hc219f0a6, 32'hc1a2cea6, 32'h425be4b1, 32'h41caba31};
test_output[6800:6807] = '{32'h0, 32'h426f77bd, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425be4b1, 32'h41caba31};
test_input[6808:6815] = '{32'hc011152b, 32'h425baa72, 32'hc1792f10, 32'hc2687efa, 32'hc2a2f659, 32'h41978c25, 32'hc2170fe0, 32'hc15fc257};
test_output[6808:6815] = '{32'h0, 32'h425baa72, 32'h0, 32'h0, 32'h0, 32'h41978c25, 32'h0, 32'h0};
test_input[6816:6823] = '{32'h41fc6919, 32'hc28ef12d, 32'h421d1498, 32'h3f89383d, 32'hc24b4091, 32'h4090a4e6, 32'h4259aa27, 32'hc2bd4b1c};
test_output[6816:6823] = '{32'h41fc6919, 32'h0, 32'h421d1498, 32'h3f89383d, 32'h0, 32'h4090a4e6, 32'h4259aa27, 32'h0};
test_input[6824:6831] = '{32'h423d3052, 32'h429d36a4, 32'h41974e3e, 32'h42a08170, 32'h421c0195, 32'hc18a14f2, 32'hc1ad60e7, 32'hc281864f};
test_output[6824:6831] = '{32'h423d3052, 32'h429d36a4, 32'h41974e3e, 32'h42a08170, 32'h421c0195, 32'h0, 32'h0, 32'h0};
test_input[6832:6839] = '{32'h41665b68, 32'h4195a3b8, 32'h41dd692e, 32'h42937afa, 32'hc223bd8a, 32'h41995b63, 32'h4106caa7, 32'h412d71b5};
test_output[6832:6839] = '{32'h41665b68, 32'h4195a3b8, 32'h41dd692e, 32'h42937afa, 32'h0, 32'h41995b63, 32'h4106caa7, 32'h412d71b5};
test_input[6840:6847] = '{32'hc0e0ae84, 32'h41e632e9, 32'hc1737384, 32'h427bf883, 32'h42971ca3, 32'h429ff9b1, 32'h426e573a, 32'h4294de9f};
test_output[6840:6847] = '{32'h0, 32'h41e632e9, 32'h0, 32'h427bf883, 32'h42971ca3, 32'h429ff9b1, 32'h426e573a, 32'h4294de9f};
test_input[6848:6855] = '{32'hc10a684d, 32'h3ff7da86, 32'hc2a05676, 32'hc28d5658, 32'hc2b0e0b8, 32'hc2393f21, 32'h427c0692, 32'hc2b8fc75};
test_output[6848:6855] = '{32'h0, 32'h3ff7da86, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427c0692, 32'h0};
test_input[6856:6863] = '{32'h42293b90, 32'hc2b4a2ed, 32'h41751e9e, 32'hc1ea73de, 32'h40473e8a, 32'h40682b9f, 32'hc29ec12e, 32'h42183ae1};
test_output[6856:6863] = '{32'h42293b90, 32'h0, 32'h41751e9e, 32'h0, 32'h40473e8a, 32'h40682b9f, 32'h0, 32'h42183ae1};
test_input[6864:6871] = '{32'hc2b66b33, 32'h41e33fcd, 32'hc1e3a404, 32'hc09d8009, 32'hc2be72fa, 32'hc2699f31, 32'hc0e0c142, 32'hc2ad17e8};
test_output[6864:6871] = '{32'h0, 32'h41e33fcd, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6872:6879] = '{32'h4221c76e, 32'hc28e6ace, 32'hc23d3e06, 32'h40d01736, 32'hc1a7ed76, 32'h4272e1aa, 32'h4246b1f0, 32'hc2bfd84f};
test_output[6872:6879] = '{32'h4221c76e, 32'h0, 32'h0, 32'h40d01736, 32'h0, 32'h4272e1aa, 32'h4246b1f0, 32'h0};
test_input[6880:6887] = '{32'hc18933bc, 32'h42b26c13, 32'hc2b0ee42, 32'hc2aab123, 32'h429a7344, 32'h41db5449, 32'hc03f464f, 32'hc2b6dee1};
test_output[6880:6887] = '{32'h0, 32'h42b26c13, 32'h0, 32'h0, 32'h429a7344, 32'h41db5449, 32'h0, 32'h0};
test_input[6888:6895] = '{32'hc1923a36, 32'hc1c7257a, 32'h41cc1989, 32'hc210360e, 32'h4297941c, 32'h4238f094, 32'hc128ec05, 32'h41139d33};
test_output[6888:6895] = '{32'h0, 32'h0, 32'h41cc1989, 32'h0, 32'h4297941c, 32'h4238f094, 32'h0, 32'h41139d33};
test_input[6896:6903] = '{32'h40ba98ff, 32'hc1f33e5f, 32'h41fedb6d, 32'hc1e83a6f, 32'h42b1bbdd, 32'hc2aeb586, 32'hc2add92c, 32'h4025cec2};
test_output[6896:6903] = '{32'h40ba98ff, 32'h0, 32'h41fedb6d, 32'h0, 32'h42b1bbdd, 32'h0, 32'h0, 32'h4025cec2};
test_input[6904:6911] = '{32'h42b877ba, 32'h420b2745, 32'hc2bc1cb3, 32'h425fc4fa, 32'h4284be6f, 32'h41b217dd, 32'h42316a48, 32'hc28faa71};
test_output[6904:6911] = '{32'h42b877ba, 32'h420b2745, 32'h0, 32'h425fc4fa, 32'h4284be6f, 32'h41b217dd, 32'h42316a48, 32'h0};
test_input[6912:6919] = '{32'hc05baae3, 32'hc2491f07, 32'h4181308f, 32'hc27105b3, 32'h425ecbc1, 32'h428d31fc, 32'hc2a45e2d, 32'hc13a0438};
test_output[6912:6919] = '{32'h0, 32'h0, 32'h4181308f, 32'h0, 32'h425ecbc1, 32'h428d31fc, 32'h0, 32'h0};
test_input[6920:6927] = '{32'hc1c0a520, 32'hc2bbc290, 32'hc147c355, 32'h42748f68, 32'h4298d836, 32'h42ac59eb, 32'hc2763ef0, 32'hc28f6de4};
test_output[6920:6927] = '{32'h0, 32'h0, 32'h0, 32'h42748f68, 32'h4298d836, 32'h42ac59eb, 32'h0, 32'h0};
test_input[6928:6935] = '{32'hc2261002, 32'hc25dcc15, 32'hc25e2309, 32'hc2620a9f, 32'h419af103, 32'h427d5d72, 32'hc1aa879a, 32'hc1453ed1};
test_output[6928:6935] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h419af103, 32'h427d5d72, 32'h0, 32'h0};
test_input[6936:6943] = '{32'hc28f174b, 32'h426ad29d, 32'hc25f12d3, 32'h42282821, 32'h42bdebfb, 32'h428b6d4c, 32'hc2b8738b, 32'h421f9e2d};
test_output[6936:6943] = '{32'h0, 32'h426ad29d, 32'h0, 32'h42282821, 32'h42bdebfb, 32'h428b6d4c, 32'h0, 32'h421f9e2d};
test_input[6944:6951] = '{32'h42583db0, 32'h42c738e1, 32'h4172b955, 32'hc246be9d, 32'h425ced21, 32'hc0575aaa, 32'h4205ae9a, 32'h42581792};
test_output[6944:6951] = '{32'h42583db0, 32'h42c738e1, 32'h4172b955, 32'h0, 32'h425ced21, 32'h0, 32'h4205ae9a, 32'h42581792};
test_input[6952:6959] = '{32'hc2ab7375, 32'hc290266f, 32'h42a3c4c3, 32'h4291f68a, 32'h41f63f66, 32'h41d1a48e, 32'h41228fa2, 32'hc2a78927};
test_output[6952:6959] = '{32'h0, 32'h0, 32'h42a3c4c3, 32'h4291f68a, 32'h41f63f66, 32'h41d1a48e, 32'h41228fa2, 32'h0};
test_input[6960:6967] = '{32'hc1fde18e, 32'hc00a7a9f, 32'hc2c7da16, 32'hc1c1cdd1, 32'h4195befb, 32'hc2887947, 32'hc2778393, 32'hc23bfe24};
test_output[6960:6967] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4195befb, 32'h0, 32'h0, 32'h0};
test_input[6968:6975] = '{32'h41d0c2da, 32'h429d31f9, 32'h42b8ceec, 32'h42c3ca2e, 32'h4290cdf6, 32'hc29d9722, 32'h41ee1d5b, 32'h429478a2};
test_output[6968:6975] = '{32'h41d0c2da, 32'h429d31f9, 32'h42b8ceec, 32'h42c3ca2e, 32'h4290cdf6, 32'h0, 32'h41ee1d5b, 32'h429478a2};
test_input[6976:6983] = '{32'hc267479a, 32'hc2255509, 32'hc28349b5, 32'h4092d736, 32'hc2648918, 32'hc23e059e, 32'hc0fa7993, 32'hc17b61f7};
test_output[6976:6983] = '{32'h0, 32'h0, 32'h0, 32'h4092d736, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[6984:6991] = '{32'hc29b7ca9, 32'hc223c9b5, 32'h41bc11bc, 32'h416ace6b, 32'hc2b84808, 32'h42ab7eff, 32'h427b2dcc, 32'hc2997473};
test_output[6984:6991] = '{32'h0, 32'h0, 32'h41bc11bc, 32'h416ace6b, 32'h0, 32'h42ab7eff, 32'h427b2dcc, 32'h0};
test_input[6992:6999] = '{32'hc15f9b01, 32'h427e0887, 32'hc25eed86, 32'hc16abbc0, 32'h42bdf72d, 32'h41b8d004, 32'hc273ebd5, 32'hc1c2675c};
test_output[6992:6999] = '{32'h0, 32'h427e0887, 32'h0, 32'h0, 32'h42bdf72d, 32'h41b8d004, 32'h0, 32'h0};
test_input[7000:7007] = '{32'h427aff3e, 32'h4173bc02, 32'h41f79667, 32'hc22e1e43, 32'hc151e459, 32'h427a68d1, 32'h42c2385b, 32'hc293e12c};
test_output[7000:7007] = '{32'h427aff3e, 32'h4173bc02, 32'h41f79667, 32'h0, 32'h0, 32'h427a68d1, 32'h42c2385b, 32'h0};
test_input[7008:7015] = '{32'h40ca472f, 32'hc273d046, 32'h42c21482, 32'h42a73f57, 32'h426ce9e1, 32'hc2ba435a, 32'h4223137c, 32'hc2585a2a};
test_output[7008:7015] = '{32'h40ca472f, 32'h0, 32'h42c21482, 32'h42a73f57, 32'h426ce9e1, 32'h0, 32'h4223137c, 32'h0};
test_input[7016:7023] = '{32'h41fc0fd8, 32'hc292debc, 32'h42658e7f, 32'h427cce59, 32'h4253ad22, 32'h4296326d, 32'h41d3b65d, 32'hc2999828};
test_output[7016:7023] = '{32'h41fc0fd8, 32'h0, 32'h42658e7f, 32'h427cce59, 32'h4253ad22, 32'h4296326d, 32'h41d3b65d, 32'h0};
test_input[7024:7031] = '{32'hc2a015dd, 32'h428dbcee, 32'h3db36e88, 32'hc28e169a, 32'hc2af47b1, 32'hc2ab1157, 32'h4227c465, 32'h428a68da};
test_output[7024:7031] = '{32'h0, 32'h428dbcee, 32'h3db36e88, 32'h0, 32'h0, 32'h0, 32'h4227c465, 32'h428a68da};
test_input[7032:7039] = '{32'hc10115d7, 32'h42a61f87, 32'h42aa2d77, 32'h42518f6b, 32'hc148dae0, 32'hc26264ea, 32'h409200f7, 32'hc1dd032d};
test_output[7032:7039] = '{32'h0, 32'h42a61f87, 32'h42aa2d77, 32'h42518f6b, 32'h0, 32'h0, 32'h409200f7, 32'h0};
test_input[7040:7047] = '{32'h429d4345, 32'h418a8208, 32'hc1f61971, 32'h424c20c2, 32'hc24e3532, 32'hc1be6ac5, 32'h42251f89, 32'h426a2f14};
test_output[7040:7047] = '{32'h429d4345, 32'h418a8208, 32'h0, 32'h424c20c2, 32'h0, 32'h0, 32'h42251f89, 32'h426a2f14};
test_input[7048:7055] = '{32'hc267a52b, 32'h42568f63, 32'h428d53d8, 32'hc0a00e31, 32'hc17dca11, 32'h425b1847, 32'h426ea2c9, 32'hc2891cfc};
test_output[7048:7055] = '{32'h0, 32'h42568f63, 32'h428d53d8, 32'h0, 32'h0, 32'h425b1847, 32'h426ea2c9, 32'h0};
test_input[7056:7063] = '{32'h4277359d, 32'h42a1017e, 32'hc1a662bd, 32'hc20cc624, 32'h42c35fef, 32'h404785b3, 32'h41748423, 32'hc2598caa};
test_output[7056:7063] = '{32'h4277359d, 32'h42a1017e, 32'h0, 32'h0, 32'h42c35fef, 32'h404785b3, 32'h41748423, 32'h0};
test_input[7064:7071] = '{32'hc2a3fb7a, 32'h40523901, 32'h425aa226, 32'h427818d8, 32'hc2be0959, 32'hc26b8aaa, 32'hc112a208, 32'h411019e1};
test_output[7064:7071] = '{32'h0, 32'h40523901, 32'h425aa226, 32'h427818d8, 32'h0, 32'h0, 32'h0, 32'h411019e1};
test_input[7072:7079] = '{32'hc2184896, 32'h41c7af30, 32'h4291db49, 32'hc2c14c9c, 32'hc20b372b, 32'h424ec968, 32'hc21bf1b3, 32'h42a277e5};
test_output[7072:7079] = '{32'h0, 32'h41c7af30, 32'h4291db49, 32'h0, 32'h0, 32'h424ec968, 32'h0, 32'h42a277e5};
test_input[7080:7087] = '{32'hc1b4141f, 32'h423ce862, 32'hc290d6d3, 32'h429759de, 32'h4240c293, 32'hc25004dc, 32'h41f1e15b, 32'h422e2cc2};
test_output[7080:7087] = '{32'h0, 32'h423ce862, 32'h0, 32'h429759de, 32'h4240c293, 32'h0, 32'h41f1e15b, 32'h422e2cc2};
test_input[7088:7095] = '{32'h4023dea4, 32'h40a68644, 32'hc210fd18, 32'h426d6eb5, 32'hc2a6d80e, 32'hc065f360, 32'hc2bf0b46, 32'hc291fbdf};
test_output[7088:7095] = '{32'h4023dea4, 32'h40a68644, 32'h0, 32'h426d6eb5, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7096:7103] = '{32'hc05edfc4, 32'h4273abca, 32'hc2936f1c, 32'hc2891144, 32'hc22c7f3d, 32'h419a9485, 32'hc241381c, 32'h41745dd2};
test_output[7096:7103] = '{32'h0, 32'h4273abca, 32'h0, 32'h0, 32'h0, 32'h419a9485, 32'h0, 32'h41745dd2};
test_input[7104:7111] = '{32'hc19a48ab, 32'hbfe6d334, 32'hc245a31a, 32'hc25c9d83, 32'h419ea4db, 32'h421c7419, 32'h42babd77, 32'hc2c21809};
test_output[7104:7111] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h419ea4db, 32'h421c7419, 32'h42babd77, 32'h0};
test_input[7112:7119] = '{32'h40e12a7f, 32'h42200b1f, 32'h41e26a6b, 32'hc29c0202, 32'hc276be51, 32'h41909c09, 32'h42a3d8be, 32'hc2b51304};
test_output[7112:7119] = '{32'h40e12a7f, 32'h42200b1f, 32'h41e26a6b, 32'h0, 32'h0, 32'h41909c09, 32'h42a3d8be, 32'h0};
test_input[7120:7127] = '{32'h40168bd1, 32'hc2213547, 32'h42a9341b, 32'h41471b1f, 32'hc294de4a, 32'h42a5a34a, 32'h42728833, 32'h41def56a};
test_output[7120:7127] = '{32'h40168bd1, 32'h0, 32'h42a9341b, 32'h41471b1f, 32'h0, 32'h42a5a34a, 32'h42728833, 32'h41def56a};
test_input[7128:7135] = '{32'hc2986a46, 32'hc0a9c132, 32'hc2c0178d, 32'h42aec3d7, 32'hc11f811d, 32'hc2b03b15, 32'h42566647, 32'hc0784400};
test_output[7128:7135] = '{32'h0, 32'h0, 32'h0, 32'h42aec3d7, 32'h0, 32'h0, 32'h42566647, 32'h0};
test_input[7136:7143] = '{32'h4222400a, 32'h422a32ea, 32'h42b01d9a, 32'h4293b064, 32'h42ace340, 32'hc234a17b, 32'h41d8ada1, 32'hc27cfda6};
test_output[7136:7143] = '{32'h4222400a, 32'h422a32ea, 32'h42b01d9a, 32'h4293b064, 32'h42ace340, 32'h0, 32'h41d8ada1, 32'h0};
test_input[7144:7151] = '{32'h41810b22, 32'h427d3689, 32'hc2b43946, 32'hc285d338, 32'h428c56ae, 32'h41ff7ae9, 32'h40f9e758, 32'h41b8571a};
test_output[7144:7151] = '{32'h41810b22, 32'h427d3689, 32'h0, 32'h0, 32'h428c56ae, 32'h41ff7ae9, 32'h40f9e758, 32'h41b8571a};
test_input[7152:7159] = '{32'hc16c90cf, 32'hc26bee96, 32'hc0806e7a, 32'hc2b390fc, 32'hc212d295, 32'h42273271, 32'h42c74b2e, 32'hc14fcd2e};
test_output[7152:7159] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42273271, 32'h42c74b2e, 32'h0};
test_input[7160:7167] = '{32'hc2846f95, 32'h421d356f, 32'hc2105d2e, 32'h421579c2, 32'hc0c152f7, 32'h428ccaad, 32'hc2a81eb3, 32'hc29f7f3b};
test_output[7160:7167] = '{32'h0, 32'h421d356f, 32'h0, 32'h421579c2, 32'h0, 32'h428ccaad, 32'h0, 32'h0};
test_input[7168:7175] = '{32'h41df74b8, 32'hc2476511, 32'hc1300415, 32'hc21c143e, 32'hc2959cc2, 32'h42860c5e, 32'hc2975882, 32'hc2674c2e};
test_output[7168:7175] = '{32'h41df74b8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42860c5e, 32'h0, 32'h0};
test_input[7176:7183] = '{32'hc21a6045, 32'h42bdacaa, 32'h403c0dc2, 32'hc28f26c4, 32'h4264d752, 32'hc2584ed0, 32'hc0193ee0, 32'hc2476b67};
test_output[7176:7183] = '{32'h0, 32'h42bdacaa, 32'h403c0dc2, 32'h0, 32'h4264d752, 32'h0, 32'h0, 32'h0};
test_input[7184:7191] = '{32'h4121e9e6, 32'h4293bc57, 32'h42c55671, 32'hc2a883dd, 32'h4286617d, 32'h4256aacc, 32'h42595957, 32'h429ea1b3};
test_output[7184:7191] = '{32'h4121e9e6, 32'h4293bc57, 32'h42c55671, 32'h0, 32'h4286617d, 32'h4256aacc, 32'h42595957, 32'h429ea1b3};
test_input[7192:7199] = '{32'h421af1eb, 32'hc24fed4a, 32'h42902307, 32'h419ec8ba, 32'h4258b8a3, 32'hc21aad6d, 32'h4100283c, 32'h41c4fcf0};
test_output[7192:7199] = '{32'h421af1eb, 32'h0, 32'h42902307, 32'h419ec8ba, 32'h4258b8a3, 32'h0, 32'h4100283c, 32'h41c4fcf0};
test_input[7200:7207] = '{32'hc248efb1, 32'h402c9761, 32'h429ae010, 32'h4297d356, 32'hc28d1d40, 32'hc247120d, 32'hc1483c4b, 32'h429a4aab};
test_output[7200:7207] = '{32'h0, 32'h402c9761, 32'h429ae010, 32'h4297d356, 32'h0, 32'h0, 32'h0, 32'h429a4aab};
test_input[7208:7215] = '{32'hc166ce8c, 32'hc1bbdd89, 32'hc145dd8f, 32'hc2274cff, 32'h42ba16f8, 32'h41ded503, 32'h42705d10, 32'hc286937a};
test_output[7208:7215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42ba16f8, 32'h41ded503, 32'h42705d10, 32'h0};
test_input[7216:7223] = '{32'hc2408a8d, 32'hc12ecbbd, 32'h41c929b2, 32'h418c0f77, 32'h3fd298fb, 32'h4286c65f, 32'hc0f9233c, 32'h4295115a};
test_output[7216:7223] = '{32'h0, 32'h0, 32'h41c929b2, 32'h418c0f77, 32'h3fd298fb, 32'h4286c65f, 32'h0, 32'h4295115a};
test_input[7224:7231] = '{32'h42b9597a, 32'hc0c7397d, 32'h3f482543, 32'h42b9dff7, 32'hc259bc24, 32'hc22aa45c, 32'hc2a77d90, 32'hc29921c4};
test_output[7224:7231] = '{32'h42b9597a, 32'h0, 32'h3f482543, 32'h42b9dff7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7232:7239] = '{32'h4211dd70, 32'h4211b614, 32'h422287ce, 32'h42561ab2, 32'h42bcd147, 32'hc2b845a9, 32'h40a080ef, 32'h41590c7f};
test_output[7232:7239] = '{32'h4211dd70, 32'h4211b614, 32'h422287ce, 32'h42561ab2, 32'h42bcd147, 32'h0, 32'h40a080ef, 32'h41590c7f};
test_input[7240:7247] = '{32'h3f1031da, 32'hc1dd6f40, 32'hc2b6ce39, 32'hc136b5f7, 32'hc1c23864, 32'hc2be5047, 32'hc1668e1c, 32'hc20b46e0};
test_output[7240:7247] = '{32'h3f1031da, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7248:7255] = '{32'h42b04c20, 32'h3d562c59, 32'h4296628f, 32'hc295a28a, 32'h42780895, 32'h42627923, 32'h42128a22, 32'h42680d9c};
test_output[7248:7255] = '{32'h42b04c20, 32'h3d562c59, 32'h4296628f, 32'h0, 32'h42780895, 32'h42627923, 32'h42128a22, 32'h42680d9c};
test_input[7256:7263] = '{32'h428b4ed8, 32'hc29418fe, 32'h423823db, 32'h425e40fd, 32'hc0b85e2e, 32'h4241c6c8, 32'h42866202, 32'hc16601f3};
test_output[7256:7263] = '{32'h428b4ed8, 32'h0, 32'h423823db, 32'h425e40fd, 32'h0, 32'h4241c6c8, 32'h42866202, 32'h0};
test_input[7264:7271] = '{32'h4299edbe, 32'hc22292c8, 32'h4237b533, 32'hc236e91d, 32'h42b0d3dd, 32'h41ac4e28, 32'hc2bd8265, 32'hc1a1c7eb};
test_output[7264:7271] = '{32'h4299edbe, 32'h0, 32'h4237b533, 32'h0, 32'h42b0d3dd, 32'h41ac4e28, 32'h0, 32'h0};
test_input[7272:7279] = '{32'hc1f30d80, 32'hc2c3e515, 32'hc2b4f4d0, 32'h421b7547, 32'hc2893a24, 32'hc2c2ae10, 32'hc143a40e, 32'hc1fad3f8};
test_output[7272:7279] = '{32'h0, 32'h0, 32'h0, 32'h421b7547, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7280:7287] = '{32'hc28d4238, 32'hc2bcb5ac, 32'hc20a4997, 32'h42b7034a, 32'h42b61923, 32'hc2aaea67, 32'h424b903f, 32'hc28931ea};
test_output[7280:7287] = '{32'h0, 32'h0, 32'h0, 32'h42b7034a, 32'h42b61923, 32'h0, 32'h424b903f, 32'h0};
test_input[7288:7295] = '{32'h423352f1, 32'hc2a77d9f, 32'h42649830, 32'hc165afa3, 32'hc0152f72, 32'h42a3d42b, 32'h426ccf71, 32'hc0671d83};
test_output[7288:7295] = '{32'h423352f1, 32'h0, 32'h42649830, 32'h0, 32'h0, 32'h42a3d42b, 32'h426ccf71, 32'h0};
test_input[7296:7303] = '{32'hc2c68b08, 32'hc2c4cc81, 32'hc2c13dcb, 32'hc2039868, 32'hc1c99f68, 32'hc26f7d6c, 32'h415f5714, 32'hbf0c2ae7};
test_output[7296:7303] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h415f5714, 32'h0};
test_input[7304:7311] = '{32'h426f4c4c, 32'h429de646, 32'h41009b06, 32'hc2baf782, 32'h4232b378, 32'h422338c2, 32'hc21ff9b9, 32'h42abdadb};
test_output[7304:7311] = '{32'h426f4c4c, 32'h429de646, 32'h41009b06, 32'h0, 32'h4232b378, 32'h422338c2, 32'h0, 32'h42abdadb};
test_input[7312:7319] = '{32'hc26686ba, 32'h4228a72f, 32'h42b8cff4, 32'hc2bd8646, 32'hc19323be, 32'hc281be57, 32'hc0da14f4, 32'h428b276b};
test_output[7312:7319] = '{32'h0, 32'h4228a72f, 32'h42b8cff4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428b276b};
test_input[7320:7327] = '{32'h42402478, 32'hc1a37eb1, 32'h418f9b8b, 32'h420e03ad, 32'h428e6792, 32'hc2a97280, 32'hc19b1ee0, 32'h4285d883};
test_output[7320:7327] = '{32'h42402478, 32'h0, 32'h418f9b8b, 32'h420e03ad, 32'h428e6792, 32'h0, 32'h0, 32'h4285d883};
test_input[7328:7335] = '{32'h41d923a8, 32'hc2bc24fe, 32'hbfc81685, 32'hc29d8096, 32'h41a7ddd5, 32'hc219edfd, 32'h419b744a, 32'h4226f949};
test_output[7328:7335] = '{32'h41d923a8, 32'h0, 32'h0, 32'h0, 32'h41a7ddd5, 32'h0, 32'h419b744a, 32'h4226f949};
test_input[7336:7343] = '{32'h42b2894d, 32'hc2a3dc95, 32'h42b02933, 32'h40d0260a, 32'h424dfd76, 32'hc238dd20, 32'h42b9a111, 32'hc170ade5};
test_output[7336:7343] = '{32'h42b2894d, 32'h0, 32'h42b02933, 32'h40d0260a, 32'h424dfd76, 32'h0, 32'h42b9a111, 32'h0};
test_input[7344:7351] = '{32'h423bdfef, 32'hc2c3480b, 32'h41a4817d, 32'hc23f8256, 32'h427c388a, 32'h42947a16, 32'hc2c1b8a8, 32'h42a689da};
test_output[7344:7351] = '{32'h423bdfef, 32'h0, 32'h41a4817d, 32'h0, 32'h427c388a, 32'h42947a16, 32'h0, 32'h42a689da};
test_input[7352:7359] = '{32'h4221fefa, 32'h42b3ccca, 32'hc271d066, 32'h4210f487, 32'h42a5a6f1, 32'hc267956f, 32'h422545ce, 32'hc260e1fc};
test_output[7352:7359] = '{32'h4221fefa, 32'h42b3ccca, 32'h0, 32'h4210f487, 32'h42a5a6f1, 32'h0, 32'h422545ce, 32'h0};
test_input[7360:7367] = '{32'h404e49fb, 32'hc282ded7, 32'hc19e3b90, 32'hc215eb79, 32'hc1c4a54d, 32'h41bbe1e9, 32'hc29f5db5, 32'h42598073};
test_output[7360:7367] = '{32'h404e49fb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41bbe1e9, 32'h0, 32'h42598073};
test_input[7368:7375] = '{32'h41b91d4e, 32'hc2634173, 32'h3eac0583, 32'hc28d0a4d, 32'h41d86c7b, 32'h3f4c0359, 32'h42535225, 32'h4298ea80};
test_output[7368:7375] = '{32'h41b91d4e, 32'h0, 32'h3eac0583, 32'h0, 32'h41d86c7b, 32'h3f4c0359, 32'h42535225, 32'h4298ea80};
test_input[7376:7383] = '{32'h42c0ef1f, 32'hc2846433, 32'h4188703e, 32'h42b663cc, 32'hc1b84b74, 32'hc29a87bb, 32'hc242596b, 32'h429bcc88};
test_output[7376:7383] = '{32'h42c0ef1f, 32'h0, 32'h4188703e, 32'h42b663cc, 32'h0, 32'h0, 32'h0, 32'h429bcc88};
test_input[7384:7391] = '{32'hc1738c96, 32'hc28aa842, 32'hc20f7c05, 32'hc2432b05, 32'h411b34b1, 32'h42972932, 32'hc1a1d8ce, 32'h41a3c547};
test_output[7384:7391] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h411b34b1, 32'h42972932, 32'h0, 32'h41a3c547};
test_input[7392:7399] = '{32'h427ed562, 32'hc166ef20, 32'hc2535b3a, 32'hc1a8dc68, 32'hc26a4bd0, 32'h42a52275, 32'hc23ac2de, 32'hc28f5e5d};
test_output[7392:7399] = '{32'h427ed562, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a52275, 32'h0, 32'h0};
test_input[7400:7407] = '{32'h42b530e4, 32'hc2b89c0b, 32'h42a9973d, 32'h4089f5a0, 32'h42a702d0, 32'h42c4b116, 32'h41c32fda, 32'h41cd05a3};
test_output[7400:7407] = '{32'h42b530e4, 32'h0, 32'h42a9973d, 32'h4089f5a0, 32'h42a702d0, 32'h42c4b116, 32'h41c32fda, 32'h41cd05a3};
test_input[7408:7415] = '{32'hc1989e92, 32'hc24dc33b, 32'h3fb1ba27, 32'h418d4e0c, 32'h411b8841, 32'hbe1fb095, 32'h42413803, 32'hbec8699e};
test_output[7408:7415] = '{32'h0, 32'h0, 32'h3fb1ba27, 32'h418d4e0c, 32'h411b8841, 32'h0, 32'h42413803, 32'h0};
test_input[7416:7423] = '{32'hc266d175, 32'hc127b341, 32'hc20082b0, 32'h42b3b290, 32'h4265c06f, 32'h42c77dea, 32'h428a63ba, 32'hc1b30175};
test_output[7416:7423] = '{32'h0, 32'h0, 32'h0, 32'h42b3b290, 32'h4265c06f, 32'h42c77dea, 32'h428a63ba, 32'h0};
test_input[7424:7431] = '{32'hbfe7ca39, 32'hc2963705, 32'hc2b91a3d, 32'hc23b620e, 32'hc28c6bef, 32'h429e5213, 32'hc2b890cd, 32'hc23371ff};
test_output[7424:7431] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429e5213, 32'h0, 32'h0};
test_input[7432:7439] = '{32'h40a5a161, 32'h41de7a44, 32'h42389e96, 32'hc296e3f3, 32'h4297e6ec, 32'hc29fa139, 32'hc0e1e27b, 32'h42c604bc};
test_output[7432:7439] = '{32'h40a5a161, 32'h41de7a44, 32'h42389e96, 32'h0, 32'h4297e6ec, 32'h0, 32'h0, 32'h42c604bc};
test_input[7440:7447] = '{32'hc1357b1a, 32'h419bf259, 32'hc232529c, 32'h3fc7d9da, 32'hc2a0ca4c, 32'hc2c34553, 32'hc1aca3a0, 32'h421144b3};
test_output[7440:7447] = '{32'h0, 32'h419bf259, 32'h0, 32'h3fc7d9da, 32'h0, 32'h0, 32'h0, 32'h421144b3};
test_input[7448:7455] = '{32'hc2c55af1, 32'h429f021d, 32'hc210e61b, 32'hc2b06d35, 32'h42aefa8e, 32'hc2c1a049, 32'hc1288e6d, 32'hc279731f};
test_output[7448:7455] = '{32'h0, 32'h429f021d, 32'h0, 32'h0, 32'h42aefa8e, 32'h0, 32'h0, 32'h0};
test_input[7456:7463] = '{32'h42a79cde, 32'h4260833b, 32'h427998ae, 32'h421d6368, 32'h4209eef7, 32'hc0d3609a, 32'hc25ac6a8, 32'h4007c388};
test_output[7456:7463] = '{32'h42a79cde, 32'h4260833b, 32'h427998ae, 32'h421d6368, 32'h4209eef7, 32'h0, 32'h0, 32'h4007c388};
test_input[7464:7471] = '{32'h4002bb30, 32'hc25be239, 32'h412742af, 32'h4298ce60, 32'hc28eab4b, 32'hc1be09f5, 32'hc297fcae, 32'h421088da};
test_output[7464:7471] = '{32'h4002bb30, 32'h0, 32'h412742af, 32'h4298ce60, 32'h0, 32'h0, 32'h0, 32'h421088da};
test_input[7472:7479] = '{32'hc08c03f5, 32'h428d05be, 32'hc161d2e6, 32'hc29bd0c7, 32'hc271e06f, 32'h41a68d4a, 32'h42bd2023, 32'h4211ca11};
test_output[7472:7479] = '{32'h0, 32'h428d05be, 32'h0, 32'h0, 32'h0, 32'h41a68d4a, 32'h42bd2023, 32'h4211ca11};
test_input[7480:7487] = '{32'hc209034f, 32'hc2a14235, 32'hc13eb182, 32'h3fadeac9, 32'hc158a5e6, 32'h42bb8b87, 32'hc2b386f8, 32'h42981dd0};
test_output[7480:7487] = '{32'h0, 32'h0, 32'h0, 32'h3fadeac9, 32'h0, 32'h42bb8b87, 32'h0, 32'h42981dd0};
test_input[7488:7495] = '{32'hc1e5e9b6, 32'hc2138a27, 32'hc28773e9, 32'h40e904b7, 32'h420152c0, 32'hc217a746, 32'h42282bf1, 32'hc235a8f2};
test_output[7488:7495] = '{32'h0, 32'h0, 32'h0, 32'h40e904b7, 32'h420152c0, 32'h0, 32'h42282bf1, 32'h0};
test_input[7496:7503] = '{32'hc22dc07b, 32'h418c6427, 32'hc2289a1c, 32'hc29b43bd, 32'h4299bd2d, 32'h42c290eb, 32'h418e1b48, 32'h425ed17e};
test_output[7496:7503] = '{32'h0, 32'h418c6427, 32'h0, 32'h0, 32'h4299bd2d, 32'h42c290eb, 32'h418e1b48, 32'h425ed17e};
test_input[7504:7511] = '{32'h42c6a49b, 32'h42aea902, 32'h425b6a68, 32'hc26589d7, 32'h418e4a95, 32'h40810d51, 32'h42937233, 32'h3faaec40};
test_output[7504:7511] = '{32'h42c6a49b, 32'h42aea902, 32'h425b6a68, 32'h0, 32'h418e4a95, 32'h40810d51, 32'h42937233, 32'h3faaec40};
test_input[7512:7519] = '{32'h42bb23b5, 32'hc23f88f5, 32'h40dd652b, 32'hc2c7fa9d, 32'hc228361f, 32'h42619f52, 32'hc0cca74f, 32'h4191dc52};
test_output[7512:7519] = '{32'h42bb23b5, 32'h0, 32'h40dd652b, 32'h0, 32'h0, 32'h42619f52, 32'h0, 32'h4191dc52};
test_input[7520:7527] = '{32'h4207cd23, 32'hc29648f5, 32'h4274414f, 32'hc2c1f965, 32'hc261977d, 32'h428bb68f, 32'h420aa269, 32'hc2a6d1c1};
test_output[7520:7527] = '{32'h4207cd23, 32'h0, 32'h4274414f, 32'h0, 32'h0, 32'h428bb68f, 32'h420aa269, 32'h0};
test_input[7528:7535] = '{32'hc1d5a193, 32'hc146c961, 32'h42a64bda, 32'hc289d641, 32'hc1c0cc12, 32'hc1460afa, 32'hbfac5055, 32'hc2032c5c};
test_output[7528:7535] = '{32'h0, 32'h0, 32'h42a64bda, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[7536:7543] = '{32'h41e2dee6, 32'h41b6217e, 32'h424372d4, 32'hc08fbe5c, 32'h429513c2, 32'h426efa74, 32'hc28cfd94, 32'h41f52777};
test_output[7536:7543] = '{32'h41e2dee6, 32'h41b6217e, 32'h424372d4, 32'h0, 32'h429513c2, 32'h426efa74, 32'h0, 32'h41f52777};
test_input[7544:7551] = '{32'h42114e41, 32'h3ef49bd4, 32'hc18df92f, 32'h419c4fc9, 32'h40c61355, 32'h42a58844, 32'h41b3d043, 32'hc1d08dbb};
test_output[7544:7551] = '{32'h42114e41, 32'h3ef49bd4, 32'h0, 32'h419c4fc9, 32'h40c61355, 32'h42a58844, 32'h41b3d043, 32'h0};
test_input[7552:7559] = '{32'hc0644089, 32'h42b9e1fd, 32'h42bfa427, 32'h4268f75c, 32'hc28c54f6, 32'h4205b330, 32'hc1c9f86c, 32'h42801233};
test_output[7552:7559] = '{32'h0, 32'h42b9e1fd, 32'h42bfa427, 32'h4268f75c, 32'h0, 32'h4205b330, 32'h0, 32'h42801233};
test_input[7560:7567] = '{32'h42a844b2, 32'h4250facc, 32'hc1f10cfd, 32'hc1861588, 32'h42a6c4e6, 32'h42b6bbff, 32'hc2b6edb9, 32'h41ccf2d6};
test_output[7560:7567] = '{32'h42a844b2, 32'h4250facc, 32'h0, 32'h0, 32'h42a6c4e6, 32'h42b6bbff, 32'h0, 32'h41ccf2d6};
test_input[7568:7575] = '{32'hc24ccc10, 32'hc2b711b4, 32'h429a80b7, 32'h3f99f9cb, 32'h42694fbf, 32'hc2416db1, 32'h42a38798, 32'h42648701};
test_output[7568:7575] = '{32'h0, 32'h0, 32'h429a80b7, 32'h3f99f9cb, 32'h42694fbf, 32'h0, 32'h42a38798, 32'h42648701};
test_input[7576:7583] = '{32'h428bd724, 32'hc1ae7c9a, 32'h422e616f, 32'h4201aee8, 32'hc1bfed29, 32'hc1d15cd2, 32'hc2136f2c, 32'h42aac074};
test_output[7576:7583] = '{32'h428bd724, 32'h0, 32'h422e616f, 32'h4201aee8, 32'h0, 32'h0, 32'h0, 32'h42aac074};
test_input[7584:7591] = '{32'hc238d5cd, 32'h4268b7a4, 32'h413b74cf, 32'hc1bfe6f2, 32'h3f5f1f15, 32'h4244a4d0, 32'hc1352869, 32'h4249ddd9};
test_output[7584:7591] = '{32'h0, 32'h4268b7a4, 32'h413b74cf, 32'h0, 32'h3f5f1f15, 32'h4244a4d0, 32'h0, 32'h4249ddd9};
test_input[7592:7599] = '{32'hc1a157d7, 32'h429f08c5, 32'hc28e8570, 32'h420b603f, 32'hc2a6549f, 32'h4253ae0b, 32'h42b8be6d, 32'hc2c71e64};
test_output[7592:7599] = '{32'h0, 32'h429f08c5, 32'h0, 32'h420b603f, 32'h0, 32'h4253ae0b, 32'h42b8be6d, 32'h0};
test_input[7600:7607] = '{32'h42c1dcef, 32'h42b381aa, 32'h4295a5b6, 32'h425350ed, 32'h428e73ae, 32'h42827ae3, 32'hc23066ed, 32'h41c0d6e7};
test_output[7600:7607] = '{32'h42c1dcef, 32'h42b381aa, 32'h4295a5b6, 32'h425350ed, 32'h428e73ae, 32'h42827ae3, 32'h0, 32'h41c0d6e7};
test_input[7608:7615] = '{32'hc0fcc804, 32'hc2ba599c, 32'hc2214733, 32'h42a90430, 32'h42130e8c, 32'h42855f67, 32'h428b93cc, 32'hc2739e18};
test_output[7608:7615] = '{32'h0, 32'h0, 32'h0, 32'h42a90430, 32'h42130e8c, 32'h42855f67, 32'h428b93cc, 32'h0};
test_input[7616:7623] = '{32'h424e91bb, 32'h4246b4fb, 32'hc2af4c26, 32'h4208de8d, 32'h40c417f9, 32'h42b0ae62, 32'h422eb178, 32'hc2b83f00};
test_output[7616:7623] = '{32'h424e91bb, 32'h4246b4fb, 32'h0, 32'h4208de8d, 32'h40c417f9, 32'h42b0ae62, 32'h422eb178, 32'h0};
test_input[7624:7631] = '{32'hc1c0898e, 32'h42a379cf, 32'h424617f1, 32'hc284b18e, 32'hc25931df, 32'h428bccc4, 32'h4284b7ac, 32'hc1764e70};
test_output[7624:7631] = '{32'h0, 32'h42a379cf, 32'h424617f1, 32'h0, 32'h0, 32'h428bccc4, 32'h4284b7ac, 32'h0};
test_input[7632:7639] = '{32'hc1690ed0, 32'hc215b9e3, 32'h42a960b1, 32'hc2b07ad8, 32'h42b442d5, 32'hc24b7127, 32'h4102fee6, 32'hc2a9fced};
test_output[7632:7639] = '{32'h0, 32'h0, 32'h42a960b1, 32'h0, 32'h42b442d5, 32'h0, 32'h4102fee6, 32'h0};
test_input[7640:7647] = '{32'hc2445b0a, 32'h42287430, 32'hc2653f54, 32'h4131e518, 32'hc2243caa, 32'h41b3bbdd, 32'hc2a66213, 32'hc2491763};
test_output[7640:7647] = '{32'h0, 32'h42287430, 32'h0, 32'h4131e518, 32'h0, 32'h41b3bbdd, 32'h0, 32'h0};
test_input[7648:7655] = '{32'h425b00a8, 32'hc26dd009, 32'h42013331, 32'h41f453aa, 32'hc265a8c3, 32'h4168e7dd, 32'hc2c113a2, 32'h417ce341};
test_output[7648:7655] = '{32'h425b00a8, 32'h0, 32'h42013331, 32'h41f453aa, 32'h0, 32'h4168e7dd, 32'h0, 32'h417ce341};
test_input[7656:7663] = '{32'h422b93af, 32'hc0ca8bbb, 32'h421dc345, 32'h422aa168, 32'hc1875a72, 32'hc187815e, 32'hc29e2502, 32'h429e3ac9};
test_output[7656:7663] = '{32'h422b93af, 32'h0, 32'h421dc345, 32'h422aa168, 32'h0, 32'h0, 32'h0, 32'h429e3ac9};
test_input[7664:7671] = '{32'h421bfbd7, 32'hc0ceb9ec, 32'hc112218c, 32'h42869ada, 32'hc1bbbe11, 32'h42801c40, 32'hc2591708, 32'h417b30ee};
test_output[7664:7671] = '{32'h421bfbd7, 32'h0, 32'h0, 32'h42869ada, 32'h0, 32'h42801c40, 32'h0, 32'h417b30ee};
test_input[7672:7679] = '{32'h42383e7e, 32'h424b33ac, 32'hc28a602c, 32'hc2863a6f, 32'h422d77c9, 32'h42814ee2, 32'h42aff51e, 32'hc286fd84};
test_output[7672:7679] = '{32'h42383e7e, 32'h424b33ac, 32'h0, 32'h0, 32'h422d77c9, 32'h42814ee2, 32'h42aff51e, 32'h0};
test_input[7680:7687] = '{32'h3ffc038e, 32'hbf4250ca, 32'h424d1ccd, 32'h42357372, 32'h4253b6fa, 32'h426980c6, 32'hc2a756d5, 32'h419a1bae};
test_output[7680:7687] = '{32'h3ffc038e, 32'h0, 32'h424d1ccd, 32'h42357372, 32'h4253b6fa, 32'h426980c6, 32'h0, 32'h419a1bae};
test_input[7688:7695] = '{32'h42796a55, 32'h4217aa31, 32'h424c87c0, 32'hc02051bc, 32'hc23b1434, 32'h421f632e, 32'h41908cbf, 32'hc2bf1617};
test_output[7688:7695] = '{32'h42796a55, 32'h4217aa31, 32'h424c87c0, 32'h0, 32'h0, 32'h421f632e, 32'h41908cbf, 32'h0};
test_input[7696:7703] = '{32'h4001f50d, 32'h41e21b20, 32'h42ba4757, 32'h423499c4, 32'h4263d1df, 32'hc05ed143, 32'h4188f12a, 32'hc0bfb872};
test_output[7696:7703] = '{32'h4001f50d, 32'h41e21b20, 32'h42ba4757, 32'h423499c4, 32'h4263d1df, 32'h0, 32'h4188f12a, 32'h0};
test_input[7704:7711] = '{32'hc28c39de, 32'hc2752b46, 32'h423cab73, 32'hc2c558a0, 32'hc0e6b2d6, 32'h3fc01475, 32'hc2721560, 32'h42460d67};
test_output[7704:7711] = '{32'h0, 32'h0, 32'h423cab73, 32'h0, 32'h0, 32'h3fc01475, 32'h0, 32'h42460d67};
test_input[7712:7719] = '{32'hc1fa1117, 32'h4198c0fe, 32'h420943ff, 32'h42bc9362, 32'h42ad1c23, 32'h42156950, 32'hc1fd42c8, 32'h41c7e57e};
test_output[7712:7719] = '{32'h0, 32'h4198c0fe, 32'h420943ff, 32'h42bc9362, 32'h42ad1c23, 32'h42156950, 32'h0, 32'h41c7e57e};
test_input[7720:7727] = '{32'hc29f6afc, 32'h425ae670, 32'h4282b5ef, 32'h4221397e, 32'h42b88b60, 32'hc262bf5b, 32'hc275d864, 32'h423f2334};
test_output[7720:7727] = '{32'h0, 32'h425ae670, 32'h4282b5ef, 32'h4221397e, 32'h42b88b60, 32'h0, 32'h0, 32'h423f2334};
test_input[7728:7735] = '{32'h422b9bdd, 32'hc293b1e2, 32'hbf3eaff9, 32'hc24f4fab, 32'hc29e76ca, 32'hc29938ac, 32'h422245e4, 32'hc21809ce};
test_output[7728:7735] = '{32'h422b9bdd, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422245e4, 32'h0};
test_input[7736:7743] = '{32'hc28943e2, 32'h423d7b80, 32'hc19397e5, 32'h423b1f50, 32'h42b23ee8, 32'h422ff4fb, 32'h4297f6f0, 32'hc2ad7065};
test_output[7736:7743] = '{32'h0, 32'h423d7b80, 32'h0, 32'h423b1f50, 32'h42b23ee8, 32'h422ff4fb, 32'h4297f6f0, 32'h0};
test_input[7744:7751] = '{32'h42963864, 32'hc2a5bf10, 32'hc1fa5af8, 32'hc2ad5325, 32'hc2c15c9d, 32'hc0faed7e, 32'h429402d6, 32'h42c705d5};
test_output[7744:7751] = '{32'h42963864, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429402d6, 32'h42c705d5};
test_input[7752:7759] = '{32'hc28003ba, 32'hc2b0cd84, 32'h42402722, 32'hc2ab563c, 32'hc1bf9ca3, 32'hc275800b, 32'h42794d28, 32'h42878132};
test_output[7752:7759] = '{32'h0, 32'h0, 32'h42402722, 32'h0, 32'h0, 32'h0, 32'h42794d28, 32'h42878132};
test_input[7760:7767] = '{32'hc2b0b790, 32'hc28766c6, 32'h41c0c8b7, 32'h42977f87, 32'hc1e24610, 32'hc175997d, 32'h42c43762, 32'h41b8aa65};
test_output[7760:7767] = '{32'h0, 32'h0, 32'h41c0c8b7, 32'h42977f87, 32'h0, 32'h0, 32'h42c43762, 32'h41b8aa65};
test_input[7768:7775] = '{32'hc290eb45, 32'hc2ab3b5c, 32'h422d8dbb, 32'h4189c61b, 32'hc24ebe23, 32'hc2a93395, 32'hc119c735, 32'h423ff2a1};
test_output[7768:7775] = '{32'h0, 32'h0, 32'h422d8dbb, 32'h4189c61b, 32'h0, 32'h0, 32'h0, 32'h423ff2a1};
test_input[7776:7783] = '{32'h42418756, 32'hc248e2e0, 32'h42afe8b7, 32'hbf40ebd8, 32'h422b91cb, 32'hc29f3a5d, 32'h40a3d9c9, 32'h425c0214};
test_output[7776:7783] = '{32'h42418756, 32'h0, 32'h42afe8b7, 32'h0, 32'h422b91cb, 32'h0, 32'h40a3d9c9, 32'h425c0214};
test_input[7784:7791] = '{32'h4218c25f, 32'hc0861668, 32'h42ac38df, 32'h417e48ec, 32'hc1b62319, 32'h42a13bfa, 32'h41ae5fa9, 32'hc22e6eda};
test_output[7784:7791] = '{32'h4218c25f, 32'h0, 32'h42ac38df, 32'h417e48ec, 32'h0, 32'h42a13bfa, 32'h41ae5fa9, 32'h0};
test_input[7792:7799] = '{32'h42bb49cf, 32'hc26ea09d, 32'h41b5e24c, 32'hc2bc5e44, 32'h428a676b, 32'h42ac360b, 32'h42a07f5b, 32'hc1ac0d7c};
test_output[7792:7799] = '{32'h42bb49cf, 32'h0, 32'h41b5e24c, 32'h0, 32'h428a676b, 32'h42ac360b, 32'h42a07f5b, 32'h0};
test_input[7800:7807] = '{32'hc1940b5a, 32'h4130b27e, 32'h3f822aa3, 32'hc26faabf, 32'h42ae2fca, 32'h423e4c7d, 32'h424b243e, 32'hc29d7604};
test_output[7800:7807] = '{32'h0, 32'h4130b27e, 32'h3f822aa3, 32'h0, 32'h42ae2fca, 32'h423e4c7d, 32'h424b243e, 32'h0};
test_input[7808:7815] = '{32'hc200ed21, 32'h42b41757, 32'h4267ceea, 32'h42978eed, 32'h42bebe15, 32'hc28ef50a, 32'h426315e3, 32'hc22fb220};
test_output[7808:7815] = '{32'h0, 32'h42b41757, 32'h4267ceea, 32'h42978eed, 32'h42bebe15, 32'h0, 32'h426315e3, 32'h0};
test_input[7816:7823] = '{32'hc21f620d, 32'h425245d9, 32'h429f8d79, 32'h429495be, 32'hc292494a, 32'hc051263d, 32'h403dc519, 32'h42049a3e};
test_output[7816:7823] = '{32'h0, 32'h425245d9, 32'h429f8d79, 32'h429495be, 32'h0, 32'h0, 32'h403dc519, 32'h42049a3e};
test_input[7824:7831] = '{32'hc0c1338a, 32'hc2c3dbe3, 32'hc291d5a6, 32'h42b1ab74, 32'hc2c2d5cf, 32'h42a52936, 32'hbfcac309, 32'hc17ab013};
test_output[7824:7831] = '{32'h0, 32'h0, 32'h0, 32'h42b1ab74, 32'h0, 32'h42a52936, 32'h0, 32'h0};
test_input[7832:7839] = '{32'h4039e490, 32'hbf457526, 32'hc200c9c1, 32'h4107fd4e, 32'hc29d295f, 32'hc0a5254f, 32'hc1ac65a4, 32'h429a46c8};
test_output[7832:7839] = '{32'h4039e490, 32'h0, 32'h0, 32'h4107fd4e, 32'h0, 32'h0, 32'h0, 32'h429a46c8};
test_input[7840:7847] = '{32'hc2568264, 32'hc2bbb5c0, 32'h413fcf95, 32'hc2925b20, 32'hc1ddf8b6, 32'hc28084e4, 32'h41327847, 32'hc2c0b40f};
test_output[7840:7847] = '{32'h0, 32'h0, 32'h413fcf95, 32'h0, 32'h0, 32'h0, 32'h41327847, 32'h0};
test_input[7848:7855] = '{32'hc26f6791, 32'hc1351499, 32'h42b6988e, 32'h42078b9b, 32'hc29081a0, 32'h422c9f75, 32'h41676430, 32'h4104e129};
test_output[7848:7855] = '{32'h0, 32'h0, 32'h42b6988e, 32'h42078b9b, 32'h0, 32'h422c9f75, 32'h41676430, 32'h4104e129};
test_input[7856:7863] = '{32'hc153d933, 32'h428af7c1, 32'hc232abf6, 32'h42423024, 32'hc27b842a, 32'hc258b42d, 32'h4286f201, 32'h40e898c6};
test_output[7856:7863] = '{32'h0, 32'h428af7c1, 32'h0, 32'h42423024, 32'h0, 32'h0, 32'h4286f201, 32'h40e898c6};
test_input[7864:7871] = '{32'h421a48ae, 32'h42ad5e20, 32'h42aa6fa9, 32'h41de5247, 32'h42057977, 32'h4234829e, 32'h41fa8557, 32'hc1717394};
test_output[7864:7871] = '{32'h421a48ae, 32'h42ad5e20, 32'h42aa6fa9, 32'h41de5247, 32'h42057977, 32'h4234829e, 32'h41fa8557, 32'h0};
test_input[7872:7879] = '{32'hc249deba, 32'h4210ff4a, 32'hc074d71b, 32'h427db7b8, 32'h427f2a7a, 32'hc108460e, 32'hc18171b0, 32'hc1d16947};
test_output[7872:7879] = '{32'h0, 32'h4210ff4a, 32'h0, 32'h427db7b8, 32'h427f2a7a, 32'h0, 32'h0, 32'h0};
test_input[7880:7887] = '{32'hc28c213d, 32'hbf438f22, 32'hc275e370, 32'hc0fe6dcb, 32'h42127cef, 32'h40e75dbc, 32'h42a4fc12, 32'hc21f5d63};
test_output[7880:7887] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42127cef, 32'h40e75dbc, 32'h42a4fc12, 32'h0};
test_input[7888:7895] = '{32'h42b57770, 32'hc290b391, 32'h412551a9, 32'h424242fb, 32'h402cac1f, 32'h42b265ce, 32'h40f3e31a, 32'hc180c5c8};
test_output[7888:7895] = '{32'h42b57770, 32'h0, 32'h412551a9, 32'h424242fb, 32'h402cac1f, 32'h42b265ce, 32'h40f3e31a, 32'h0};
test_input[7896:7903] = '{32'hc231dbdc, 32'hc02d5c6f, 32'h429f309e, 32'hc2538c26, 32'hc2b2bc8a, 32'h4299fbde, 32'hc2950076, 32'h41b59771};
test_output[7896:7903] = '{32'h0, 32'h0, 32'h429f309e, 32'h0, 32'h0, 32'h4299fbde, 32'h0, 32'h41b59771};
test_input[7904:7911] = '{32'h40d3be28, 32'hc19dd57f, 32'h423b9f23, 32'h42648ff3, 32'hc1c28ae2, 32'h4277a3e9, 32'hc23a7850, 32'h42a3a1a8};
test_output[7904:7911] = '{32'h40d3be28, 32'h0, 32'h423b9f23, 32'h42648ff3, 32'h0, 32'h4277a3e9, 32'h0, 32'h42a3a1a8};
test_input[7912:7919] = '{32'h41bb4b00, 32'hc298f579, 32'hc2b92cd1, 32'hc1f43f19, 32'h42b14c63, 32'h4288d149, 32'hc2bf8407, 32'hc2c2e41d};
test_output[7912:7919] = '{32'h41bb4b00, 32'h0, 32'h0, 32'h0, 32'h42b14c63, 32'h4288d149, 32'h0, 32'h0};
test_input[7920:7927] = '{32'hc299000d, 32'hc09f9395, 32'h42b1414f, 32'hc28b1ef6, 32'h428ed199, 32'hc26b4f76, 32'hc087959f, 32'hc2880c59};
test_output[7920:7927] = '{32'h0, 32'h0, 32'h42b1414f, 32'h0, 32'h428ed199, 32'h0, 32'h0, 32'h0};
test_input[7928:7935] = '{32'hc241bdaf, 32'h429e7e52, 32'hc1b055a4, 32'hc1adc0fc, 32'h41c15849, 32'h425240a8, 32'hc15022b2, 32'h42b14dfa};
test_output[7928:7935] = '{32'h0, 32'h429e7e52, 32'h0, 32'h0, 32'h41c15849, 32'h425240a8, 32'h0, 32'h42b14dfa};
test_input[7936:7943] = '{32'hc2804c67, 32'hc1104cbc, 32'hc2231a73, 32'h42aa6ad7, 32'hc26f9924, 32'hc213e95d, 32'h42a367ad, 32'h42b068f6};
test_output[7936:7943] = '{32'h0, 32'h0, 32'h0, 32'h42aa6ad7, 32'h0, 32'h0, 32'h42a367ad, 32'h42b068f6};
test_input[7944:7951] = '{32'h428ee82a, 32'h41df6b81, 32'hc224ce7e, 32'hc1bfd4b5, 32'hc21011c0, 32'h42b3ab27, 32'h42bf7acf, 32'h41a4a9de};
test_output[7944:7951] = '{32'h428ee82a, 32'h41df6b81, 32'h0, 32'h0, 32'h0, 32'h42b3ab27, 32'h42bf7acf, 32'h41a4a9de};
test_input[7952:7959] = '{32'hc296f60f, 32'hc2162766, 32'hc157433b, 32'hc2b25e99, 32'hc191fe10, 32'h41b65991, 32'h41318395, 32'h42134577};
test_output[7952:7959] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b65991, 32'h41318395, 32'h42134577};
test_input[7960:7967] = '{32'h42bbd37c, 32'h42823135, 32'hc1fb3666, 32'hc259850f, 32'hc2264f15, 32'hc2562e6d, 32'h428c643b, 32'h420f4c52};
test_output[7960:7967] = '{32'h42bbd37c, 32'h42823135, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428c643b, 32'h420f4c52};
test_input[7968:7975] = '{32'hc12afb8b, 32'hc296695e, 32'hc25b0197, 32'h428d5395, 32'h41c3d913, 32'h429482ba, 32'h429f679f, 32'hc1124452};
test_output[7968:7975] = '{32'h0, 32'h0, 32'h0, 32'h428d5395, 32'h41c3d913, 32'h429482ba, 32'h429f679f, 32'h0};
test_input[7976:7983] = '{32'hc13f8d67, 32'h3f88ed5f, 32'hc2bda934, 32'hc2bfe306, 32'h413b8bc1, 32'h42a382fa, 32'hc19b5e50, 32'h42c15c3c};
test_output[7976:7983] = '{32'h0, 32'h3f88ed5f, 32'h0, 32'h0, 32'h413b8bc1, 32'h42a382fa, 32'h0, 32'h42c15c3c};
test_input[7984:7991] = '{32'hc297daa9, 32'h427a1ee4, 32'h41025ec7, 32'h41f72655, 32'hc25ed49b, 32'h422112f4, 32'h41b24966, 32'hc03970e9};
test_output[7984:7991] = '{32'h0, 32'h427a1ee4, 32'h41025ec7, 32'h41f72655, 32'h0, 32'h422112f4, 32'h41b24966, 32'h0};
test_input[7992:7999] = '{32'h4245ab9e, 32'h426b0e8b, 32'hc257bc69, 32'h428e4436, 32'hc1982aaf, 32'hc29f3329, 32'h420302a0, 32'h4274fa4d};
test_output[7992:7999] = '{32'h4245ab9e, 32'h426b0e8b, 32'h0, 32'h428e4436, 32'h0, 32'h0, 32'h420302a0, 32'h4274fa4d};
test_input[8000:8007] = '{32'hc274bd60, 32'h41ed7ce3, 32'h417bc4ec, 32'hc1ccf014, 32'hc0c286dd, 32'h426ad249, 32'hc282ab13, 32'hc2971f50};
test_output[8000:8007] = '{32'h0, 32'h41ed7ce3, 32'h417bc4ec, 32'h0, 32'h0, 32'h426ad249, 32'h0, 32'h0};
test_input[8008:8015] = '{32'h42ab4f10, 32'h42446f26, 32'hc13041bf, 32'hc23c3dcd, 32'h42c276e2, 32'h41f68d63, 32'hc2a458d0, 32'h42823394};
test_output[8008:8015] = '{32'h42ab4f10, 32'h42446f26, 32'h0, 32'h0, 32'h42c276e2, 32'h41f68d63, 32'h0, 32'h42823394};
test_input[8016:8023] = '{32'h42312d99, 32'hc2c1b804, 32'h3efb4d6d, 32'hc16c7995, 32'h42360893, 32'hc121de83, 32'hc22ea738, 32'h42bfe06b};
test_output[8016:8023] = '{32'h42312d99, 32'h0, 32'h3efb4d6d, 32'h0, 32'h42360893, 32'h0, 32'h0, 32'h42bfe06b};
test_input[8024:8031] = '{32'hc17d4a9b, 32'h4255c8f7, 32'h41407740, 32'hc196cc46, 32'h4299538e, 32'h4017de55, 32'hc2a89a55, 32'h41b2f997};
test_output[8024:8031] = '{32'h0, 32'h4255c8f7, 32'h41407740, 32'h0, 32'h4299538e, 32'h4017de55, 32'h0, 32'h41b2f997};
test_input[8032:8039] = '{32'h4134fa23, 32'h42bccef7, 32'hc202b8f1, 32'h41d6862a, 32'hc1996e57, 32'h41900dfa, 32'h42bd5e54, 32'hc2b9df5f};
test_output[8032:8039] = '{32'h4134fa23, 32'h42bccef7, 32'h0, 32'h41d6862a, 32'h0, 32'h41900dfa, 32'h42bd5e54, 32'h0};
test_input[8040:8047] = '{32'h428cb3b1, 32'h41e59bd7, 32'h3f2b16e0, 32'hc205684e, 32'hc258bf20, 32'hbe303301, 32'hc1bc6c32, 32'hc1703451};
test_output[8040:8047] = '{32'h428cb3b1, 32'h41e59bd7, 32'h3f2b16e0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8048:8055] = '{32'hc2b324e6, 32'hc1d0b07e, 32'h4284cece, 32'h41a92e48, 32'h429bcff8, 32'hc282e5f9, 32'hc216a065, 32'hc2247f37};
test_output[8048:8055] = '{32'h0, 32'h0, 32'h4284cece, 32'h41a92e48, 32'h429bcff8, 32'h0, 32'h0, 32'h0};
test_input[8056:8063] = '{32'h424fb014, 32'hc2030707, 32'hc18047d4, 32'hc22faab5, 32'hc047ed5f, 32'hc2ad7b89, 32'hc28c99ca, 32'h42187109};
test_output[8056:8063] = '{32'h424fb014, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42187109};
test_input[8064:8071] = '{32'hc29cd38d, 32'hc1ad5784, 32'hc2a5457a, 32'hc1874fc3, 32'hc2b94642, 32'h4158fd52, 32'hc29ed609, 32'hc26604ce};
test_output[8064:8071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4158fd52, 32'h0, 32'h0};
test_input[8072:8079] = '{32'h42b72bb2, 32'hc2adadf5, 32'h423e26ff, 32'hc28c416a, 32'hc1e3b4e7, 32'hc2ae901f, 32'hc1848b90, 32'h42beae82};
test_output[8072:8079] = '{32'h42b72bb2, 32'h0, 32'h423e26ff, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42beae82};
test_input[8080:8087] = '{32'hc2b56923, 32'hc1349240, 32'hc1c27771, 32'h4069692f, 32'h42c06f84, 32'h42119639, 32'hc2c075c3, 32'hc186ead5};
test_output[8080:8087] = '{32'h0, 32'h0, 32'h0, 32'h4069692f, 32'h42c06f84, 32'h42119639, 32'h0, 32'h0};
test_input[8088:8095] = '{32'h4286323a, 32'hc1d382a0, 32'h413c97bf, 32'h41f72c25, 32'h40c44680, 32'h425f78ef, 32'h41e1e918, 32'h426519b6};
test_output[8088:8095] = '{32'h4286323a, 32'h0, 32'h413c97bf, 32'h41f72c25, 32'h40c44680, 32'h425f78ef, 32'h41e1e918, 32'h426519b6};
test_input[8096:8103] = '{32'h428f2d06, 32'h42a3c2b1, 32'hc2beb74d, 32'h420c1583, 32'h4286205b, 32'hc2bd4745, 32'hc27a6cf7, 32'h42aad302};
test_output[8096:8103] = '{32'h428f2d06, 32'h42a3c2b1, 32'h0, 32'h420c1583, 32'h4286205b, 32'h0, 32'h0, 32'h42aad302};
test_input[8104:8111] = '{32'hc1ce059c, 32'hc2c5f552, 32'hc2abd674, 32'hc226042d, 32'h40f8a26a, 32'hc11dde22, 32'hc1e3a5b6, 32'hc1b94e9e};
test_output[8104:8111] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40f8a26a, 32'h0, 32'h0, 32'h0};
test_input[8112:8119] = '{32'h3f141e32, 32'hc29b6799, 32'h424f6983, 32'h41b61bea, 32'hc1f4cbb5, 32'h4285208f, 32'hc280b5e2, 32'hc117ac8f};
test_output[8112:8119] = '{32'h3f141e32, 32'h0, 32'h424f6983, 32'h41b61bea, 32'h0, 32'h4285208f, 32'h0, 32'h0};
test_input[8120:8127] = '{32'hc18a53e7, 32'h4143ee0a, 32'hc1c5c652, 32'h42458a9f, 32'h42366bc7, 32'hc1158316, 32'hc167162e, 32'hc18b93f8};
test_output[8120:8127] = '{32'h0, 32'h4143ee0a, 32'h0, 32'h42458a9f, 32'h42366bc7, 32'h0, 32'h0, 32'h0};
test_input[8128:8135] = '{32'h420a01a5, 32'hc252556e, 32'h4290853d, 32'h3fbf121c, 32'hc22193e7, 32'h42c32db4, 32'h42b339ea, 32'hc2439fec};
test_output[8128:8135] = '{32'h420a01a5, 32'h0, 32'h4290853d, 32'h3fbf121c, 32'h0, 32'h42c32db4, 32'h42b339ea, 32'h0};
test_input[8136:8143] = '{32'h404a779d, 32'h425cfbe1, 32'h429300a6, 32'hc2b84518, 32'h412fcabd, 32'hc2900471, 32'h42c77c1c, 32'hc2b8cda5};
test_output[8136:8143] = '{32'h404a779d, 32'h425cfbe1, 32'h429300a6, 32'h0, 32'h412fcabd, 32'h0, 32'h42c77c1c, 32'h0};
test_input[8144:8151] = '{32'hc2c10b5b, 32'hc1b35d00, 32'h41dbcb08, 32'h41da5d82, 32'hc00b7d4d, 32'h414999e6, 32'hc2c04657, 32'h404603ce};
test_output[8144:8151] = '{32'h0, 32'h0, 32'h41dbcb08, 32'h41da5d82, 32'h0, 32'h414999e6, 32'h0, 32'h404603ce};
test_input[8152:8159] = '{32'hc260a000, 32'hc27e2e8d, 32'h426a4328, 32'hc205a899, 32'h42271ee4, 32'h428c7e0a, 32'hc1c96f03, 32'hc1b10704};
test_output[8152:8159] = '{32'h0, 32'h0, 32'h426a4328, 32'h0, 32'h42271ee4, 32'h428c7e0a, 32'h0, 32'h0};
test_input[8160:8167] = '{32'hc277857d, 32'h4232a1e1, 32'h424fe38e, 32'h4295e585, 32'h4285bacf, 32'h420bd597, 32'h4191c868, 32'h429a3149};
test_output[8160:8167] = '{32'h0, 32'h4232a1e1, 32'h424fe38e, 32'h4295e585, 32'h4285bacf, 32'h420bd597, 32'h4191c868, 32'h429a3149};
test_input[8168:8175] = '{32'hc255d428, 32'hc29f58d5, 32'hc11119b0, 32'h42a718ad, 32'h419a7a26, 32'h4114c3fa, 32'hc23c3275, 32'h41a358f3};
test_output[8168:8175] = '{32'h0, 32'h0, 32'h0, 32'h42a718ad, 32'h419a7a26, 32'h4114c3fa, 32'h0, 32'h41a358f3};
test_input[8176:8183] = '{32'hc1ff6e52, 32'h42c0e3d3, 32'hc0676517, 32'h428762f2, 32'h4101b810, 32'h403ea234, 32'hc2248547, 32'hc1b42463};
test_output[8176:8183] = '{32'h0, 32'h42c0e3d3, 32'h0, 32'h428762f2, 32'h4101b810, 32'h403ea234, 32'h0, 32'h0};
test_input[8184:8191] = '{32'hbfbb6554, 32'h403c0c6c, 32'hc2c49890, 32'hc25e223d, 32'hc2967bb0, 32'hc2b19b46, 32'hc1969174, 32'hc25e4ffe};
test_output[8184:8191] = '{32'h0, 32'h403c0c6c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8192:8199] = '{32'hc27d9f6f, 32'h4174f69d, 32'h408b087a, 32'h41df0dce, 32'hc2b417de, 32'hc2a88bd1, 32'h41f7e0d5, 32'hc22943a7};
test_output[8192:8199] = '{32'h0, 32'h4174f69d, 32'h408b087a, 32'h41df0dce, 32'h0, 32'h0, 32'h41f7e0d5, 32'h0};
test_input[8200:8207] = '{32'hc26c9bdc, 32'hc1455faa, 32'h41abf846, 32'hc2ab4dad, 32'h414ad3b0, 32'h4292888e, 32'hc26e8047, 32'hc272adb8};
test_output[8200:8207] = '{32'h0, 32'h0, 32'h41abf846, 32'h0, 32'h414ad3b0, 32'h4292888e, 32'h0, 32'h0};
test_input[8208:8215] = '{32'hc2b04cb6, 32'hc212645a, 32'hc2c5a545, 32'hc2805d3d, 32'h42a5a8d6, 32'h428fe8a8, 32'h41e454d7, 32'hc21115bb};
test_output[8208:8215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a5a8d6, 32'h428fe8a8, 32'h41e454d7, 32'h0};
test_input[8216:8223] = '{32'h40bd715e, 32'hc1c4a1c6, 32'h42351380, 32'h4207b9fe, 32'h42797d6f, 32'h41688f94, 32'hc2769986, 32'h42ab2891};
test_output[8216:8223] = '{32'h40bd715e, 32'h0, 32'h42351380, 32'h4207b9fe, 32'h42797d6f, 32'h41688f94, 32'h0, 32'h42ab2891};
test_input[8224:8231] = '{32'h40d5b27b, 32'h41814fe7, 32'hc1e61dda, 32'hc2bcf959, 32'hc14f7a2d, 32'hc28d1d5f, 32'h42b5d701, 32'hc2a89db1};
test_output[8224:8231] = '{32'h40d5b27b, 32'h41814fe7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b5d701, 32'h0};
test_input[8232:8239] = '{32'hc27d6741, 32'h42b12c2a, 32'h41e2b162, 32'h3f7ff071, 32'hc0fec3d5, 32'hc215fca7, 32'h4268f73e, 32'hc298cdb0};
test_output[8232:8239] = '{32'h0, 32'h42b12c2a, 32'h41e2b162, 32'h3f7ff071, 32'h0, 32'h0, 32'h4268f73e, 32'h0};
test_input[8240:8247] = '{32'hc26d634d, 32'h42803d04, 32'hc2b8d054, 32'h42aa39e7, 32'h428b525b, 32'hc210f7a8, 32'h41ad1a78, 32'hc280bd96};
test_output[8240:8247] = '{32'h0, 32'h42803d04, 32'h0, 32'h42aa39e7, 32'h428b525b, 32'h0, 32'h41ad1a78, 32'h0};
test_input[8248:8255] = '{32'hc29aa2ff, 32'h41b18344, 32'h3f03a9cf, 32'hc17e6711, 32'hc2307227, 32'hc217daf5, 32'h41c19336, 32'h42b5fec2};
test_output[8248:8255] = '{32'h0, 32'h41b18344, 32'h3f03a9cf, 32'h0, 32'h0, 32'h0, 32'h41c19336, 32'h42b5fec2};
test_input[8256:8263] = '{32'h412ca902, 32'hc24a0aeb, 32'hc286ed58, 32'hc0ce4866, 32'hc21634f4, 32'h4222862d, 32'hc2c7d1bc, 32'h42a1e2d4};
test_output[8256:8263] = '{32'h412ca902, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4222862d, 32'h0, 32'h42a1e2d4};
test_input[8264:8271] = '{32'hc22b592a, 32'h42bd7ee9, 32'hc0c832dc, 32'h4173a272, 32'hc1af31d3, 32'h4291f62e, 32'h427f6df3, 32'h42b87f07};
test_output[8264:8271] = '{32'h0, 32'h42bd7ee9, 32'h0, 32'h4173a272, 32'h0, 32'h4291f62e, 32'h427f6df3, 32'h42b87f07};
test_input[8272:8279] = '{32'h42a30f4c, 32'h40a92b42, 32'hc2090ebd, 32'h419bacd7, 32'h41d33cf0, 32'hc28ea89b, 32'h42a69796, 32'h42426f8b};
test_output[8272:8279] = '{32'h42a30f4c, 32'h40a92b42, 32'h0, 32'h419bacd7, 32'h41d33cf0, 32'h0, 32'h42a69796, 32'h42426f8b};
test_input[8280:8287] = '{32'hc29d03c0, 32'h42c6c2cc, 32'hc23ae499, 32'h4220b079, 32'hbfcb7c26, 32'h42a2d04e, 32'hc1d2deba, 32'h428769de};
test_output[8280:8287] = '{32'h0, 32'h42c6c2cc, 32'h0, 32'h4220b079, 32'h0, 32'h42a2d04e, 32'h0, 32'h428769de};
test_input[8288:8295] = '{32'h4297cbb3, 32'hc2a1e5cb, 32'h42825074, 32'h429e3e7a, 32'hc2920d66, 32'hbf9ac6e7, 32'hc2162a64, 32'hbed56b93};
test_output[8288:8295] = '{32'h4297cbb3, 32'h0, 32'h42825074, 32'h429e3e7a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8296:8303] = '{32'hc2b055ff, 32'hc2a4f067, 32'hc25010a4, 32'h42b8a12e, 32'h41aa80fe, 32'h428b167e, 32'hc0e70065, 32'h4257459d};
test_output[8296:8303] = '{32'h0, 32'h0, 32'h0, 32'h42b8a12e, 32'h41aa80fe, 32'h428b167e, 32'h0, 32'h4257459d};
test_input[8304:8311] = '{32'h40535b0c, 32'h42badbe3, 32'hc2481604, 32'h4278ee5c, 32'hc1dd5fb4, 32'h421b3dba, 32'h41ccb857, 32'h424500cb};
test_output[8304:8311] = '{32'h40535b0c, 32'h42badbe3, 32'h0, 32'h4278ee5c, 32'h0, 32'h421b3dba, 32'h41ccb857, 32'h424500cb};
test_input[8312:8319] = '{32'hc2278b46, 32'hc2b4ca3b, 32'h4253b8b9, 32'hc240812b, 32'hc202565e, 32'hbfe4d46d, 32'h42becda7, 32'hc241e332};
test_output[8312:8319] = '{32'h0, 32'h0, 32'h4253b8b9, 32'h0, 32'h0, 32'h0, 32'h42becda7, 32'h0};
test_input[8320:8327] = '{32'hc1fb16cc, 32'h4224c2cc, 32'h421b80a1, 32'hc1b18eb3, 32'hc2326ca2, 32'hc0a7b15a, 32'h42b3db85, 32'h41014654};
test_output[8320:8327] = '{32'h0, 32'h4224c2cc, 32'h421b80a1, 32'h0, 32'h0, 32'h0, 32'h42b3db85, 32'h41014654};
test_input[8328:8335] = '{32'h423fc196, 32'hc29fe75f, 32'hc1ea9dc8, 32'h4283760d, 32'hc260584e, 32'hc0abcf64, 32'hc292c64c, 32'hc299987c};
test_output[8328:8335] = '{32'h423fc196, 32'h0, 32'h0, 32'h4283760d, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8336:8343] = '{32'h41ba0ad4, 32'hc23c5ad3, 32'hc0c2f228, 32'hc2bff3e2, 32'hc298397c, 32'hc2845487, 32'h42009213, 32'hc0316b50};
test_output[8336:8343] = '{32'h41ba0ad4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42009213, 32'h0};
test_input[8344:8351] = '{32'hc275d82f, 32'h42613096, 32'h42c30c05, 32'hc07d785e, 32'h421d21ea, 32'hc2090648, 32'hc110353a, 32'h4272c206};
test_output[8344:8351] = '{32'h0, 32'h42613096, 32'h42c30c05, 32'h0, 32'h421d21ea, 32'h0, 32'h0, 32'h4272c206};
test_input[8352:8359] = '{32'hc28a4f05, 32'h42c28439, 32'hc2867738, 32'h42c0ce24, 32'hc0eccaec, 32'h40b40c50, 32'h429be289, 32'h3f6c7d45};
test_output[8352:8359] = '{32'h0, 32'h42c28439, 32'h0, 32'h42c0ce24, 32'h0, 32'h40b40c50, 32'h429be289, 32'h3f6c7d45};
test_input[8360:8367] = '{32'h4266cf1b, 32'h42a9479c, 32'h427a3e02, 32'hc2931872, 32'hc2b4e20c, 32'h4284005c, 32'hc27530b7, 32'hc1a74425};
test_output[8360:8367] = '{32'h4266cf1b, 32'h42a9479c, 32'h427a3e02, 32'h0, 32'h0, 32'h4284005c, 32'h0, 32'h0};
test_input[8368:8375] = '{32'hc1f683d8, 32'h42117757, 32'hc21c421a, 32'hc29f2bd0, 32'hc249c9e8, 32'h42556632, 32'hc1926fb5, 32'hc249d94f};
test_output[8368:8375] = '{32'h0, 32'h42117757, 32'h0, 32'h0, 32'h0, 32'h42556632, 32'h0, 32'h0};
test_input[8376:8383] = '{32'h42b5a96c, 32'h405b57b1, 32'h428b421d, 32'hc28c8093, 32'h429f77c9, 32'h42bdd71b, 32'h418ea27d, 32'h41b54a64};
test_output[8376:8383] = '{32'h42b5a96c, 32'h405b57b1, 32'h428b421d, 32'h0, 32'h429f77c9, 32'h42bdd71b, 32'h418ea27d, 32'h41b54a64};
test_input[8384:8391] = '{32'hc29b5ed9, 32'hc27f588c, 32'h413bc205, 32'h4299220c, 32'h42a7214b, 32'h40336593, 32'h41f8633c, 32'hc1c65a8f};
test_output[8384:8391] = '{32'h0, 32'h0, 32'h413bc205, 32'h4299220c, 32'h42a7214b, 32'h40336593, 32'h41f8633c, 32'h0};
test_input[8392:8399] = '{32'hbf8d7b93, 32'hc266d892, 32'hc28bf733, 32'h42bb8d31, 32'h420d83c2, 32'h4237c653, 32'h4224b8c7, 32'h4211c229};
test_output[8392:8399] = '{32'h0, 32'h0, 32'h0, 32'h42bb8d31, 32'h420d83c2, 32'h4237c653, 32'h4224b8c7, 32'h4211c229};
test_input[8400:8407] = '{32'hc113bf73, 32'h42972787, 32'h42949ed1, 32'hc24c49b8, 32'h42a4f95f, 32'hc27cc978, 32'h4295f2a3, 32'h425ebcc3};
test_output[8400:8407] = '{32'h0, 32'h42972787, 32'h42949ed1, 32'h0, 32'h42a4f95f, 32'h0, 32'h4295f2a3, 32'h425ebcc3};
test_input[8408:8415] = '{32'hc288c28a, 32'hc2b315a6, 32'h423960a5, 32'hc2c1a7e3, 32'h42237ea6, 32'h42a255eb, 32'hc09c25fb, 32'hc2a0a7a6};
test_output[8408:8415] = '{32'h0, 32'h0, 32'h423960a5, 32'h0, 32'h42237ea6, 32'h42a255eb, 32'h0, 32'h0};
test_input[8416:8423] = '{32'hc2541ae1, 32'hc254fcab, 32'h42350ea0, 32'hc2946ca3, 32'hc2923998, 32'h400e6831, 32'hc2919d9a, 32'hc2a7cf9c};
test_output[8416:8423] = '{32'h0, 32'h0, 32'h42350ea0, 32'h0, 32'h0, 32'h400e6831, 32'h0, 32'h0};
test_input[8424:8431] = '{32'h4255054c, 32'h421e4577, 32'hc2757b66, 32'hc12160a5, 32'h42c6f261, 32'hc24bd2ab, 32'h41c1eb02, 32'hc20c4611};
test_output[8424:8431] = '{32'h4255054c, 32'h421e4577, 32'h0, 32'h0, 32'h42c6f261, 32'h0, 32'h41c1eb02, 32'h0};
test_input[8432:8439] = '{32'h41fc56e0, 32'h42445336, 32'h4126d791, 32'hc20afc2d, 32'hc297e47e, 32'h4228f1d5, 32'h420832b9, 32'h42a8108f};
test_output[8432:8439] = '{32'h41fc56e0, 32'h42445336, 32'h4126d791, 32'h0, 32'h0, 32'h4228f1d5, 32'h420832b9, 32'h42a8108f};
test_input[8440:8447] = '{32'hc264526d, 32'h42a8a563, 32'hc256ca2a, 32'hc14b8909, 32'hc2b0e5a8, 32'h4228da7a, 32'h4223ba32, 32'hc1244270};
test_output[8440:8447] = '{32'h0, 32'h42a8a563, 32'h0, 32'h0, 32'h0, 32'h4228da7a, 32'h4223ba32, 32'h0};
test_input[8448:8455] = '{32'h42c32ce5, 32'h4151bd68, 32'h42acd886, 32'h4110240c, 32'hc205d8c6, 32'h42528d58, 32'hc1b3f0f3, 32'h41545da9};
test_output[8448:8455] = '{32'h42c32ce5, 32'h4151bd68, 32'h42acd886, 32'h4110240c, 32'h0, 32'h42528d58, 32'h0, 32'h41545da9};
test_input[8456:8463] = '{32'hc2819c77, 32'h411d4a66, 32'hc14ddd56, 32'h42276980, 32'hc1920eb1, 32'hc27bdc8f, 32'h429e5b54, 32'hc1fca4db};
test_output[8456:8463] = '{32'h0, 32'h411d4a66, 32'h0, 32'h42276980, 32'h0, 32'h0, 32'h429e5b54, 32'h0};
test_input[8464:8471] = '{32'h422b3519, 32'hc273d7c0, 32'hc0c39c99, 32'hc25a6247, 32'h429505b8, 32'hc1b76a2b, 32'hc267a1d0, 32'h42b29361};
test_output[8464:8471] = '{32'h422b3519, 32'h0, 32'h0, 32'h0, 32'h429505b8, 32'h0, 32'h0, 32'h42b29361};
test_input[8472:8479] = '{32'h413ffad3, 32'hc298b41e, 32'h4281091c, 32'hc2c04ec1, 32'hc2740313, 32'hc2bda14a, 32'h42bf1b01, 32'hbf601fb4};
test_output[8472:8479] = '{32'h413ffad3, 32'h0, 32'h4281091c, 32'h0, 32'h0, 32'h0, 32'h42bf1b01, 32'h0};
test_input[8480:8487] = '{32'hc1c9fb48, 32'hc270ed6e, 32'h42a56d7d, 32'h429a478d, 32'hc2c4f385, 32'h42a23a62, 32'h42ab2344, 32'h41a86a2a};
test_output[8480:8487] = '{32'h0, 32'h0, 32'h42a56d7d, 32'h429a478d, 32'h0, 32'h42a23a62, 32'h42ab2344, 32'h41a86a2a};
test_input[8488:8495] = '{32'hc1cd18cd, 32'h403117dc, 32'h429be048, 32'h4198ecd0, 32'h42a3fe64, 32'h425c5a8a, 32'hc1ad0e6a, 32'h429d3a16};
test_output[8488:8495] = '{32'h0, 32'h403117dc, 32'h429be048, 32'h4198ecd0, 32'h42a3fe64, 32'h425c5a8a, 32'h0, 32'h429d3a16};
test_input[8496:8503] = '{32'hc1db89fb, 32'h4266cedc, 32'hc290c65d, 32'hc28a633d, 32'hc284c0e1, 32'hc1d3566e, 32'hc2296dc1, 32'hc0f7137b};
test_output[8496:8503] = '{32'h0, 32'h4266cedc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8504:8511] = '{32'hc28aa011, 32'h404cd596, 32'hc2360b76, 32'h4286138c, 32'h42b09cdc, 32'h41566c25, 32'hbea1ba35, 32'h40c47aea};
test_output[8504:8511] = '{32'h0, 32'h404cd596, 32'h0, 32'h4286138c, 32'h42b09cdc, 32'h41566c25, 32'h0, 32'h40c47aea};
test_input[8512:8519] = '{32'h4076eb62, 32'h425b8034, 32'h418ac85c, 32'hc288bd70, 32'h427cd3ec, 32'h41b07b21, 32'h41ee01aa, 32'hc2c6012b};
test_output[8512:8519] = '{32'h4076eb62, 32'h425b8034, 32'h418ac85c, 32'h0, 32'h427cd3ec, 32'h41b07b21, 32'h41ee01aa, 32'h0};
test_input[8520:8527] = '{32'hc1bdde24, 32'hc2a1757c, 32'h40d7ff1d, 32'h42a2efc2, 32'hc2805a97, 32'h42b2b86b, 32'hc282ba15, 32'h42bd435a};
test_output[8520:8527] = '{32'h0, 32'h0, 32'h40d7ff1d, 32'h42a2efc2, 32'h0, 32'h42b2b86b, 32'h0, 32'h42bd435a};
test_input[8528:8535] = '{32'hc199bf1c, 32'hc152b506, 32'h4218cd21, 32'h4218e24e, 32'hc03a0a8c, 32'h425a6e39, 32'h41954443, 32'hc205060b};
test_output[8528:8535] = '{32'h0, 32'h0, 32'h4218cd21, 32'h4218e24e, 32'h0, 32'h425a6e39, 32'h41954443, 32'h0};
test_input[8536:8543] = '{32'hc2046b58, 32'hc2b38a50, 32'hc29c6b6d, 32'h425d4022, 32'hc22974e6, 32'h42960188, 32'hc19a5b3f, 32'h42152f05};
test_output[8536:8543] = '{32'h0, 32'h0, 32'h0, 32'h425d4022, 32'h0, 32'h42960188, 32'h0, 32'h42152f05};
test_input[8544:8551] = '{32'hc299b32c, 32'h42612ad0, 32'h42ad6b04, 32'h41d15ed2, 32'hc142cfae, 32'h4109bcfd, 32'h41edbe35, 32'hc0ec8fb8};
test_output[8544:8551] = '{32'h0, 32'h42612ad0, 32'h42ad6b04, 32'h41d15ed2, 32'h0, 32'h4109bcfd, 32'h41edbe35, 32'h0};
test_input[8552:8559] = '{32'h42714a82, 32'h41cbf816, 32'h42ab86b1, 32'hc290b5a8, 32'h40653738, 32'h426e0bac, 32'hc1f5c806, 32'h4255a10c};
test_output[8552:8559] = '{32'h42714a82, 32'h41cbf816, 32'h42ab86b1, 32'h0, 32'h40653738, 32'h426e0bac, 32'h0, 32'h4255a10c};
test_input[8560:8567] = '{32'h40dcfdb7, 32'hc263e17c, 32'hc1c5a831, 32'h42a7b2ed, 32'h41a2c38f, 32'h41620875, 32'h429f5c2f, 32'h425f9ca1};
test_output[8560:8567] = '{32'h40dcfdb7, 32'h0, 32'h0, 32'h42a7b2ed, 32'h41a2c38f, 32'h41620875, 32'h429f5c2f, 32'h425f9ca1};
test_input[8568:8575] = '{32'hc1a7054c, 32'hc22ed873, 32'h418c72f4, 32'hc2526ba3, 32'hc2ac9c83, 32'h42348781, 32'h426888d4, 32'h420cd674};
test_output[8568:8575] = '{32'h0, 32'h0, 32'h418c72f4, 32'h0, 32'h0, 32'h42348781, 32'h426888d4, 32'h420cd674};
test_input[8576:8583] = '{32'hc29527ae, 32'h42210027, 32'hc16bde51, 32'h420a32cf, 32'h42c18535, 32'hc2345c3e, 32'hc288ec34, 32'hc26a08a5};
test_output[8576:8583] = '{32'h0, 32'h42210027, 32'h0, 32'h420a32cf, 32'h42c18535, 32'h0, 32'h0, 32'h0};
test_input[8584:8591] = '{32'h4106e9bf, 32'h421f82df, 32'hc29c8bd1, 32'h4276c90c, 32'h402d5b56, 32'h42854e76, 32'hc21d9207, 32'hc1eb93f1};
test_output[8584:8591] = '{32'h4106e9bf, 32'h421f82df, 32'h0, 32'h4276c90c, 32'h402d5b56, 32'h42854e76, 32'h0, 32'h0};
test_input[8592:8599] = '{32'h41e1aa4c, 32'h42b1db17, 32'hc18bb45c, 32'h421c2600, 32'hc213b3b5, 32'hc2be7e95, 32'h41a3cb72, 32'hc21df024};
test_output[8592:8599] = '{32'h41e1aa4c, 32'h42b1db17, 32'h0, 32'h421c2600, 32'h0, 32'h0, 32'h41a3cb72, 32'h0};
test_input[8600:8607] = '{32'h41ff3e87, 32'h419ca4e0, 32'hc14080d2, 32'hc2bb5f98, 32'hc26ec568, 32'h42bc4549, 32'hc1e8d5d9, 32'h42c797a0};
test_output[8600:8607] = '{32'h41ff3e87, 32'h419ca4e0, 32'h0, 32'h0, 32'h0, 32'h42bc4549, 32'h0, 32'h42c797a0};
test_input[8608:8615] = '{32'h40a287dd, 32'hc2854e25, 32'h4205f021, 32'h4282d3e6, 32'h414e64d6, 32'hc2c5e3f9, 32'h42a14a9f, 32'h42b6ea3b};
test_output[8608:8615] = '{32'h40a287dd, 32'h0, 32'h4205f021, 32'h4282d3e6, 32'h414e64d6, 32'h0, 32'h42a14a9f, 32'h42b6ea3b};
test_input[8616:8623] = '{32'h429c0174, 32'h425becf7, 32'h4249337d, 32'h42750b20, 32'h4227af62, 32'hc2b0b881, 32'hc17993a4, 32'h427a820a};
test_output[8616:8623] = '{32'h429c0174, 32'h425becf7, 32'h4249337d, 32'h42750b20, 32'h4227af62, 32'h0, 32'h0, 32'h427a820a};
test_input[8624:8631] = '{32'hc11c2383, 32'hc1987754, 32'h4252698b, 32'hc1099f21, 32'hc1052c17, 32'hc14c288c, 32'hc21e672b, 32'h42a10d75};
test_output[8624:8631] = '{32'h0, 32'h0, 32'h4252698b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a10d75};
test_input[8632:8639] = '{32'h4290cd10, 32'h4280461e, 32'hc2019b7f, 32'h42af523c, 32'h4232c5dc, 32'h427d9660, 32'hc2685192, 32'hc28827be};
test_output[8632:8639] = '{32'h4290cd10, 32'h4280461e, 32'h0, 32'h42af523c, 32'h4232c5dc, 32'h427d9660, 32'h0, 32'h0};
test_input[8640:8647] = '{32'h4282909d, 32'hc1fd66b4, 32'h42c18bcf, 32'h42901126, 32'hc2aeaf2d, 32'hc1e84da8, 32'h4088a0a5, 32'hc25f4e1d};
test_output[8640:8647] = '{32'h4282909d, 32'h0, 32'h42c18bcf, 32'h42901126, 32'h0, 32'h0, 32'h4088a0a5, 32'h0};
test_input[8648:8655] = '{32'hc0c17d48, 32'hc2119b3b, 32'h419dc367, 32'h42b39845, 32'h4087a83f, 32'h428ddf1a, 32'h41d39a1b, 32'h41e108a4};
test_output[8648:8655] = '{32'h0, 32'h0, 32'h419dc367, 32'h42b39845, 32'h4087a83f, 32'h428ddf1a, 32'h41d39a1b, 32'h41e108a4};
test_input[8656:8663] = '{32'hc2831e55, 32'hc1555cd6, 32'h426c32ca, 32'hc11fae3c, 32'h3f9a64ec, 32'hc1ab3a17, 32'h429e3942, 32'hc186d49f};
test_output[8656:8663] = '{32'h0, 32'h0, 32'h426c32ca, 32'h0, 32'h3f9a64ec, 32'h0, 32'h429e3942, 32'h0};
test_input[8664:8671] = '{32'hc2806d74, 32'h426e3395, 32'h4263101c, 32'hc22a404e, 32'h428c5e62, 32'hc2822603, 32'hc292c69d, 32'h426eb27b};
test_output[8664:8671] = '{32'h0, 32'h426e3395, 32'h4263101c, 32'h0, 32'h428c5e62, 32'h0, 32'h0, 32'h426eb27b};
test_input[8672:8679] = '{32'hc28a7931, 32'h42af0721, 32'hc294dce3, 32'hc2b9f1ba, 32'hc242f8af, 32'h40cda6eb, 32'hc2ae0d7b, 32'h429ae225};
test_output[8672:8679] = '{32'h0, 32'h42af0721, 32'h0, 32'h0, 32'h0, 32'h40cda6eb, 32'h0, 32'h429ae225};
test_input[8680:8687] = '{32'h41df084b, 32'hc29b255a, 32'hc2a0dd00, 32'hc282b5b0, 32'hc1e1dd23, 32'hc262107d, 32'h42001977, 32'hc176b392};
test_output[8680:8687] = '{32'h41df084b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42001977, 32'h0};
test_input[8688:8695] = '{32'hc2822b93, 32'hc24ab616, 32'hc26a534a, 32'h4270f5de, 32'h42041461, 32'hc2349c3b, 32'hc24446d9, 32'h42768ad3};
test_output[8688:8695] = '{32'h0, 32'h0, 32'h0, 32'h4270f5de, 32'h42041461, 32'h0, 32'h0, 32'h42768ad3};
test_input[8696:8703] = '{32'hc2734485, 32'hbeaf7654, 32'h42bf4e30, 32'hc14e54f0, 32'h429e4fc4, 32'h429c12bd, 32'h42386e79, 32'h42abadc3};
test_output[8696:8703] = '{32'h0, 32'h0, 32'h42bf4e30, 32'h0, 32'h429e4fc4, 32'h429c12bd, 32'h42386e79, 32'h42abadc3};
test_input[8704:8711] = '{32'hc1d3a5c7, 32'h42097b50, 32'h42490fa0, 32'hc2903e9a, 32'hc20d811d, 32'hc234d8ad, 32'h404481a7, 32'hc2826298};
test_output[8704:8711] = '{32'h0, 32'h42097b50, 32'h42490fa0, 32'h0, 32'h0, 32'h0, 32'h404481a7, 32'h0};
test_input[8712:8719] = '{32'h419d49d8, 32'hc2c16dee, 32'hc2893821, 32'h42a3edeb, 32'hc1259497, 32'hc2b56c59, 32'h42a49c29, 32'hc2993195};
test_output[8712:8719] = '{32'h419d49d8, 32'h0, 32'h0, 32'h42a3edeb, 32'h0, 32'h0, 32'h42a49c29, 32'h0};
test_input[8720:8727] = '{32'h40f74346, 32'h42c4472e, 32'h42c5eb30, 32'hc26abb6c, 32'h428f15e9, 32'h411ea11a, 32'hc2aab429, 32'h419a07ac};
test_output[8720:8727] = '{32'h40f74346, 32'h42c4472e, 32'h42c5eb30, 32'h0, 32'h428f15e9, 32'h411ea11a, 32'h0, 32'h419a07ac};
test_input[8728:8735] = '{32'hc1ed63ef, 32'hc2c52924, 32'h42592f11, 32'hc061e16a, 32'h429bb8c3, 32'hc153e07d, 32'hc2bf152d, 32'h4291b089};
test_output[8728:8735] = '{32'h0, 32'h0, 32'h42592f11, 32'h0, 32'h429bb8c3, 32'h0, 32'h0, 32'h4291b089};
test_input[8736:8743] = '{32'hc2bbd166, 32'hc261c158, 32'hc21ed731, 32'hc1eb1e0c, 32'h42501394, 32'h41330dcf, 32'h41ef889f, 32'hc1822691};
test_output[8736:8743] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42501394, 32'h41330dcf, 32'h41ef889f, 32'h0};
test_input[8744:8751] = '{32'hc27c1731, 32'hc2b76898, 32'hc17b6327, 32'h42bf650d, 32'hc1d3d5ef, 32'hc1915085, 32'h42b870a3, 32'h41d2b799};
test_output[8744:8751] = '{32'h0, 32'h0, 32'h0, 32'h42bf650d, 32'h0, 32'h0, 32'h42b870a3, 32'h41d2b799};
test_input[8752:8759] = '{32'hc249e53f, 32'hc28ff142, 32'h42491bb6, 32'hc200c1dd, 32'h42a58ed0, 32'hc2a26a12, 32'hc2c0c5af, 32'hc1a2dd96};
test_output[8752:8759] = '{32'h0, 32'h0, 32'h42491bb6, 32'h0, 32'h42a58ed0, 32'h0, 32'h0, 32'h0};
test_input[8760:8767] = '{32'hbea3bd06, 32'h4243b113, 32'h425fa091, 32'h422ba196, 32'h42578935, 32'hc0d01f6e, 32'hc2c7f4e0, 32'h427e28fa};
test_output[8760:8767] = '{32'h0, 32'h4243b113, 32'h425fa091, 32'h422ba196, 32'h42578935, 32'h0, 32'h0, 32'h427e28fa};
test_input[8768:8775] = '{32'hc1e48861, 32'hc218b302, 32'h4202a60c, 32'hbf990c8b, 32'h42115fad, 32'hc2738f3e, 32'h41d77577, 32'hc2648d83};
test_output[8768:8775] = '{32'h0, 32'h0, 32'h4202a60c, 32'h0, 32'h42115fad, 32'h0, 32'h41d77577, 32'h0};
test_input[8776:8783] = '{32'h41e13c72, 32'hc2911b59, 32'h429ca4da, 32'hc2081231, 32'h410df821, 32'h4208bf3e, 32'hc2c390f2, 32'hc1c32167};
test_output[8776:8783] = '{32'h41e13c72, 32'h0, 32'h429ca4da, 32'h0, 32'h410df821, 32'h4208bf3e, 32'h0, 32'h0};
test_input[8784:8791] = '{32'h4205fabe, 32'h4127f03c, 32'h425af5c1, 32'h42b54708, 32'h4262eff9, 32'h42695e4d, 32'hc2a9258b, 32'hc110b46f};
test_output[8784:8791] = '{32'h4205fabe, 32'h4127f03c, 32'h425af5c1, 32'h42b54708, 32'h4262eff9, 32'h42695e4d, 32'h0, 32'h0};
test_input[8792:8799] = '{32'hc286acc1, 32'hc067c04f, 32'h41a14785, 32'h42834812, 32'hc2b9aa59, 32'hc22324d0, 32'hc29bdb40, 32'hc2a2d7a2};
test_output[8792:8799] = '{32'h0, 32'h0, 32'h41a14785, 32'h42834812, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8800:8807] = '{32'h42c0b2ac, 32'h421c409b, 32'hc2c3dd26, 32'h41de01d7, 32'h428005a5, 32'h421220c9, 32'h420fc7c4, 32'hc1b7ed14};
test_output[8800:8807] = '{32'h42c0b2ac, 32'h421c409b, 32'h0, 32'h41de01d7, 32'h428005a5, 32'h421220c9, 32'h420fc7c4, 32'h0};
test_input[8808:8815] = '{32'hc1337165, 32'hc2ad5b05, 32'hc2132934, 32'h42937bdb, 32'hc21abca7, 32'hc26fb2f4, 32'h42350b56, 32'h429279ad};
test_output[8808:8815] = '{32'h0, 32'h0, 32'h0, 32'h42937bdb, 32'h0, 32'h0, 32'h42350b56, 32'h429279ad};
test_input[8816:8823] = '{32'h427fb5c8, 32'h414be66a, 32'hc10337a5, 32'hc0221e8e, 32'h42801f8f, 32'h4115c596, 32'h429c078a, 32'hc27c1325};
test_output[8816:8823] = '{32'h427fb5c8, 32'h414be66a, 32'h0, 32'h0, 32'h42801f8f, 32'h4115c596, 32'h429c078a, 32'h0};
test_input[8824:8831] = '{32'h429f7127, 32'h421594d3, 32'h41e08896, 32'hc137d1f9, 32'h421d1ea6, 32'h412d1f96, 32'hc2545c8f, 32'hc248fd9e};
test_output[8824:8831] = '{32'h429f7127, 32'h421594d3, 32'h41e08896, 32'h0, 32'h421d1ea6, 32'h412d1f96, 32'h0, 32'h0};
test_input[8832:8839] = '{32'h421f663e, 32'hc29f6865, 32'h4291bb0e, 32'h3ff58031, 32'h42c5b00d, 32'h419b8ed9, 32'h42310e39, 32'hc29c81d1};
test_output[8832:8839] = '{32'h421f663e, 32'h0, 32'h4291bb0e, 32'h3ff58031, 32'h42c5b00d, 32'h419b8ed9, 32'h42310e39, 32'h0};
test_input[8840:8847] = '{32'hc2b5a7a4, 32'h42a85ade, 32'h42b31aac, 32'h421785c4, 32'h42420bba, 32'hc14df2c4, 32'h41a878e5, 32'h42a0f783};
test_output[8840:8847] = '{32'h0, 32'h42a85ade, 32'h42b31aac, 32'h421785c4, 32'h42420bba, 32'h0, 32'h41a878e5, 32'h42a0f783};
test_input[8848:8855] = '{32'hc29f17cb, 32'h42c61323, 32'h42604e04, 32'h4155d85c, 32'h42860f76, 32'h4280eeaa, 32'h42392cf2, 32'h42880353};
test_output[8848:8855] = '{32'h0, 32'h42c61323, 32'h42604e04, 32'h4155d85c, 32'h42860f76, 32'h4280eeaa, 32'h42392cf2, 32'h42880353};
test_input[8856:8863] = '{32'h42b28b2f, 32'h411bbd82, 32'hc1d44df8, 32'h4242088d, 32'hc28c1234, 32'hc296a3b2, 32'h40be1084, 32'h42035e9c};
test_output[8856:8863] = '{32'h42b28b2f, 32'h411bbd82, 32'h0, 32'h4242088d, 32'h0, 32'h0, 32'h40be1084, 32'h42035e9c};
test_input[8864:8871] = '{32'h41f4e484, 32'hc1a894e0, 32'h42b0870e, 32'hc1f002ae, 32'h4238296a, 32'h42af15ed, 32'hbf874f4c, 32'h425e8bea};
test_output[8864:8871] = '{32'h41f4e484, 32'h0, 32'h42b0870e, 32'h0, 32'h4238296a, 32'h42af15ed, 32'h0, 32'h425e8bea};
test_input[8872:8879] = '{32'hc2af7234, 32'hc2acdea7, 32'hc11a6ee0, 32'hc2c094ba, 32'h4184535f, 32'hc2a19c75, 32'h42a4a118, 32'h42c796c2};
test_output[8872:8879] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4184535f, 32'h0, 32'h42a4a118, 32'h42c796c2};
test_input[8880:8887] = '{32'h422d7426, 32'h415b75fe, 32'h41d2ca81, 32'hc249a102, 32'h42c18ae8, 32'hc1d57085, 32'hc202ad5e, 32'h4188453c};
test_output[8880:8887] = '{32'h422d7426, 32'h415b75fe, 32'h41d2ca81, 32'h0, 32'h42c18ae8, 32'h0, 32'h0, 32'h4188453c};
test_input[8888:8895] = '{32'h4270f96e, 32'h429c6377, 32'hc2ad4528, 32'h412b82e6, 32'hc2b2c072, 32'hc28e3ee6, 32'hc1bb5319, 32'hc23800a2};
test_output[8888:8895] = '{32'h4270f96e, 32'h429c6377, 32'h0, 32'h412b82e6, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[8896:8903] = '{32'hc0d454e0, 32'h4215ad7a, 32'hc2a52250, 32'h429a9d8a, 32'hc2637bbf, 32'h4086db52, 32'hc0c0b3d4, 32'h424121f4};
test_output[8896:8903] = '{32'h0, 32'h4215ad7a, 32'h0, 32'h429a9d8a, 32'h0, 32'h4086db52, 32'h0, 32'h424121f4};
test_input[8904:8911] = '{32'h428d3b32, 32'h42898957, 32'hc28c7477, 32'h42b8b245, 32'hc20f7395, 32'h428f020e, 32'h4123d3e3, 32'h4264ad2c};
test_output[8904:8911] = '{32'h428d3b32, 32'h42898957, 32'h0, 32'h42b8b245, 32'h0, 32'h428f020e, 32'h4123d3e3, 32'h4264ad2c};
test_input[8912:8919] = '{32'hc1063810, 32'hc0f2ae33, 32'hc2a18817, 32'h4243cd9b, 32'h42a4c51c, 32'hc10c481d, 32'h42059a31, 32'hc1e59244};
test_output[8912:8919] = '{32'h0, 32'h0, 32'h0, 32'h4243cd9b, 32'h42a4c51c, 32'h0, 32'h42059a31, 32'h0};
test_input[8920:8927] = '{32'h4138934a, 32'hbf4a10e6, 32'hc2102352, 32'h40dcf440, 32'h427cb1d8, 32'h4291cdcb, 32'hc2065ee5, 32'hc264ece1};
test_output[8920:8927] = '{32'h4138934a, 32'h0, 32'h0, 32'h40dcf440, 32'h427cb1d8, 32'h4291cdcb, 32'h0, 32'h0};
test_input[8928:8935] = '{32'h41dc02c9, 32'hc1ef50a2, 32'h40058f8b, 32'hc264f820, 32'hc18d0bff, 32'h42203e5c, 32'h42ae40a7, 32'h42bc5aab};
test_output[8928:8935] = '{32'h41dc02c9, 32'h0, 32'h40058f8b, 32'h0, 32'h0, 32'h42203e5c, 32'h42ae40a7, 32'h42bc5aab};
test_input[8936:8943] = '{32'h418b5be8, 32'h40ca53a1, 32'h42b816f9, 32'hc2bd8645, 32'h41f56b8d, 32'h429d7a35, 32'hc1aa6490, 32'hc119f2e6};
test_output[8936:8943] = '{32'h418b5be8, 32'h40ca53a1, 32'h42b816f9, 32'h0, 32'h41f56b8d, 32'h429d7a35, 32'h0, 32'h0};
test_input[8944:8951] = '{32'h4201efe3, 32'hc28ed8ef, 32'h42be5016, 32'h428c467b, 32'hc224ab9d, 32'hc2bd0ef0, 32'h42bbcec2, 32'hc2b39e0b};
test_output[8944:8951] = '{32'h4201efe3, 32'h0, 32'h42be5016, 32'h428c467b, 32'h0, 32'h0, 32'h42bbcec2, 32'h0};
test_input[8952:8959] = '{32'h42b48970, 32'hc2b4fc26, 32'hc143ac85, 32'h429365eb, 32'h42ae5c2c, 32'hc2a2aaf8, 32'hc1fd9fa2, 32'hc25a1657};
test_output[8952:8959] = '{32'h42b48970, 32'h0, 32'h0, 32'h429365eb, 32'h42ae5c2c, 32'h0, 32'h0, 32'h0};
test_input[8960:8967] = '{32'h42240b90, 32'hc24207e8, 32'hc2adff23, 32'h42be241d, 32'h428ca401, 32'h4299865f, 32'hc2c501b5, 32'hc289ab9c};
test_output[8960:8967] = '{32'h42240b90, 32'h0, 32'h0, 32'h42be241d, 32'h428ca401, 32'h4299865f, 32'h0, 32'h0};
test_input[8968:8975] = '{32'h42a52418, 32'h4214cc45, 32'hc28b0a09, 32'h4139f75f, 32'h4285cffd, 32'hc283124c, 32'hc1d56237, 32'hc2713466};
test_output[8968:8975] = '{32'h42a52418, 32'h4214cc45, 32'h0, 32'h4139f75f, 32'h4285cffd, 32'h0, 32'h0, 32'h0};
test_input[8976:8983] = '{32'h426625cb, 32'hc23ad188, 32'hc2c7ef8f, 32'hc13cb320, 32'h42543269, 32'hc12d1f3e, 32'h4269e85a, 32'hc220b14e};
test_output[8976:8983] = '{32'h426625cb, 32'h0, 32'h0, 32'h0, 32'h42543269, 32'h0, 32'h4269e85a, 32'h0};
test_input[8984:8991] = '{32'hc285cb47, 32'hc2494ae2, 32'h42bd415c, 32'h428cd0f6, 32'hc2b7e13d, 32'hc2b8eb8f, 32'h42965974, 32'h42938b19};
test_output[8984:8991] = '{32'h0, 32'h0, 32'h42bd415c, 32'h428cd0f6, 32'h0, 32'h0, 32'h42965974, 32'h42938b19};
test_input[8992:8999] = '{32'hc0d4ccfb, 32'hc0562fda, 32'h42947aff, 32'hc259970f, 32'hc112ec3a, 32'h41ad49b6, 32'h41a10eb2, 32'h40fbc510};
test_output[8992:8999] = '{32'h0, 32'h0, 32'h42947aff, 32'h0, 32'h0, 32'h41ad49b6, 32'h41a10eb2, 32'h40fbc510};
test_input[9000:9007] = '{32'hc2bd0f0a, 32'h42309781, 32'h422366b4, 32'hc284535d, 32'h42acee74, 32'h4289262d, 32'hc2a870c9, 32'hc2a22778};
test_output[9000:9007] = '{32'h0, 32'h42309781, 32'h422366b4, 32'h0, 32'h42acee74, 32'h4289262d, 32'h0, 32'h0};
test_input[9008:9015] = '{32'hc0c5a884, 32'h42bdefe4, 32'h408b8260, 32'hc244fee8, 32'hc27ab349, 32'h424866bc, 32'h4295a150, 32'h4228b390};
test_output[9008:9015] = '{32'h0, 32'h42bdefe4, 32'h408b8260, 32'h0, 32'h0, 32'h424866bc, 32'h4295a150, 32'h4228b390};
test_input[9016:9023] = '{32'h42a3fe8b, 32'h4232d107, 32'hc242402d, 32'h4201ec99, 32'h4039c969, 32'h41932ff3, 32'h41eecb5e, 32'hc252454e};
test_output[9016:9023] = '{32'h42a3fe8b, 32'h4232d107, 32'h0, 32'h4201ec99, 32'h4039c969, 32'h41932ff3, 32'h41eecb5e, 32'h0};
test_input[9024:9031] = '{32'h42b70f8b, 32'h4293131a, 32'h42635af1, 32'h42c299e9, 32'h4254d88b, 32'hc257096d, 32'h42c085b7, 32'h42880e75};
test_output[9024:9031] = '{32'h42b70f8b, 32'h4293131a, 32'h42635af1, 32'h42c299e9, 32'h4254d88b, 32'h0, 32'h42c085b7, 32'h42880e75};
test_input[9032:9039] = '{32'hc0f1bef0, 32'h41b5a671, 32'hc2361eb3, 32'hc2244659, 32'h428a22f9, 32'h412c3388, 32'h41d6a46a, 32'h418f5c32};
test_output[9032:9039] = '{32'h0, 32'h41b5a671, 32'h0, 32'h0, 32'h428a22f9, 32'h412c3388, 32'h41d6a46a, 32'h418f5c32};
test_input[9040:9047] = '{32'hc29df9b6, 32'hc25253ba, 32'h42991fce, 32'h4249a39c, 32'hbf30ff85, 32'h421556db, 32'hc243c274, 32'h42bce6be};
test_output[9040:9047] = '{32'h0, 32'h0, 32'h42991fce, 32'h4249a39c, 32'h0, 32'h421556db, 32'h0, 32'h42bce6be};
test_input[9048:9055] = '{32'hc2c2c805, 32'h421c4d9b, 32'h41b93d01, 32'h41bafe2e, 32'hc16ed224, 32'hc2181aa6, 32'hc2b679b9, 32'hc2938e4e};
test_output[9048:9055] = '{32'h0, 32'h421c4d9b, 32'h41b93d01, 32'h41bafe2e, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9056:9063] = '{32'h42b78000, 32'hc2bd1c84, 32'hc0d92146, 32'hc2666652, 32'h40c3a751, 32'h426efe1d, 32'hc2b3e71b, 32'hc18b5cac};
test_output[9056:9063] = '{32'h42b78000, 32'h0, 32'h0, 32'h0, 32'h40c3a751, 32'h426efe1d, 32'h0, 32'h0};
test_input[9064:9071] = '{32'h42568d47, 32'hc2529865, 32'hc2b8ea8d, 32'h42860a25, 32'h420ac210, 32'h4246d816, 32'hc2377e7f, 32'h41a14490};
test_output[9064:9071] = '{32'h42568d47, 32'h0, 32'h0, 32'h42860a25, 32'h420ac210, 32'h4246d816, 32'h0, 32'h41a14490};
test_input[9072:9079] = '{32'hc2429872, 32'h42b947c3, 32'hc274e456, 32'hc19af6ff, 32'hc22077b1, 32'h42c1d61d, 32'hc2be1631, 32'hc1783ee7};
test_output[9072:9079] = '{32'h0, 32'h42b947c3, 32'h0, 32'h0, 32'h0, 32'h42c1d61d, 32'h0, 32'h0};
test_input[9080:9087] = '{32'hc21a0c47, 32'hc26bd85c, 32'hc2bc7da1, 32'hc21e7c02, 32'hc1f6991a, 32'hc29d4591, 32'h418c1bd5, 32'h428734bc};
test_output[9080:9087] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h418c1bd5, 32'h428734bc};
test_input[9088:9095] = '{32'h42022233, 32'h421536d6, 32'hc2a16319, 32'hc282bc33, 32'hc2232690, 32'hc283769e, 32'hc2b3a9b9, 32'hc2717903};
test_output[9088:9095] = '{32'h42022233, 32'h421536d6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9096:9103] = '{32'h4286a9d7, 32'hc2a1e09a, 32'h41c06cf2, 32'hc235bcb7, 32'h41bf7bce, 32'h422700ce, 32'h420830cb, 32'hc28c8bf7};
test_output[9096:9103] = '{32'h4286a9d7, 32'h0, 32'h41c06cf2, 32'h0, 32'h41bf7bce, 32'h422700ce, 32'h420830cb, 32'h0};
test_input[9104:9111] = '{32'hc26af21d, 32'hc2a07d88, 32'hc1fc6877, 32'hc1c28017, 32'h42a67830, 32'h42119768, 32'hc2b0a191, 32'hc23a2bbe};
test_output[9104:9111] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a67830, 32'h42119768, 32'h0, 32'h0};
test_input[9112:9119] = '{32'hc22c74bc, 32'h42c71b50, 32'h4196bdaf, 32'hc27db9ce, 32'h41ffa624, 32'h4155316e, 32'hc225d574, 32'h4282bc28};
test_output[9112:9119] = '{32'h0, 32'h42c71b50, 32'h4196bdaf, 32'h0, 32'h41ffa624, 32'h4155316e, 32'h0, 32'h4282bc28};
test_input[9120:9127] = '{32'hc244f9aa, 32'hc1a4ecd2, 32'hc253d927, 32'hc25dcf8c, 32'h42750f12, 32'h42c5b41f, 32'hc2535fd0, 32'hc1001e3e};
test_output[9120:9127] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42750f12, 32'h42c5b41f, 32'h0, 32'h0};
test_input[9128:9135] = '{32'hc290b5de, 32'hc1eb9e6a, 32'h42c3fbc6, 32'h4208b1eb, 32'h4286c0bc, 32'h429eccb0, 32'hc0d528db, 32'h42c3c363};
test_output[9128:9135] = '{32'h0, 32'h0, 32'h42c3fbc6, 32'h4208b1eb, 32'h4286c0bc, 32'h429eccb0, 32'h0, 32'h42c3c363};
test_input[9136:9143] = '{32'hc2a5dd76, 32'hc28edf29, 32'hc13ff935, 32'hc21b838e, 32'hc1d98ebe, 32'hc213670a, 32'h42748c14, 32'hc17ea5dd};
test_output[9136:9143] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42748c14, 32'h0};
test_input[9144:9151] = '{32'h42b9629c, 32'hc208d055, 32'hc1dbbbcf, 32'h4281f57a, 32'h42a93988, 32'hc2491212, 32'hc1fc9340, 32'h428e5ad8};
test_output[9144:9151] = '{32'h42b9629c, 32'h0, 32'h0, 32'h4281f57a, 32'h42a93988, 32'h0, 32'h0, 32'h428e5ad8};
test_input[9152:9159] = '{32'h426ff982, 32'hc273caa7, 32'hc29eca0b, 32'hc28e50a4, 32'h42407b86, 32'hc2b4ab6e, 32'h40a167af, 32'h42c7d0e7};
test_output[9152:9159] = '{32'h426ff982, 32'h0, 32'h0, 32'h0, 32'h42407b86, 32'h0, 32'h40a167af, 32'h42c7d0e7};
test_input[9160:9167] = '{32'hc29fc756, 32'h4284cfaa, 32'hc29cc74f, 32'hc2a7e63c, 32'h42b62ee5, 32'h4154fecd, 32'hc0963532, 32'hc21d9d90};
test_output[9160:9167] = '{32'h0, 32'h4284cfaa, 32'h0, 32'h0, 32'h42b62ee5, 32'h4154fecd, 32'h0, 32'h0};
test_input[9168:9175] = '{32'h40f65c3e, 32'hc1f5ae98, 32'h42bdef42, 32'hc28c5427, 32'h4273d35d, 32'h42a038cb, 32'h41dc51aa, 32'hc0be9d6d};
test_output[9168:9175] = '{32'h40f65c3e, 32'h0, 32'h42bdef42, 32'h0, 32'h4273d35d, 32'h42a038cb, 32'h41dc51aa, 32'h0};
test_input[9176:9183] = '{32'h42900a06, 32'h41af57fc, 32'h42aa7562, 32'hc2c3050d, 32'h42912f79, 32'hc24e2bb7, 32'hc1bb69fa, 32'hc283d8c4};
test_output[9176:9183] = '{32'h42900a06, 32'h41af57fc, 32'h42aa7562, 32'h0, 32'h42912f79, 32'h0, 32'h0, 32'h0};
test_input[9184:9191] = '{32'hc20735d5, 32'hc2042ffc, 32'hc1e25b58, 32'hc25aad19, 32'h41029b83, 32'h41ec7790, 32'h42c14f7f, 32'hc1c9ad8e};
test_output[9184:9191] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41029b83, 32'h41ec7790, 32'h42c14f7f, 32'h0};
test_input[9192:9199] = '{32'hc29eabc4, 32'hc149c14f, 32'h4197d76a, 32'h41f0e304, 32'h42a44f16, 32'h418fe047, 32'hc1d1bb04, 32'h42aea37b};
test_output[9192:9199] = '{32'h0, 32'h0, 32'h4197d76a, 32'h41f0e304, 32'h42a44f16, 32'h418fe047, 32'h0, 32'h42aea37b};
test_input[9200:9207] = '{32'hc2a54395, 32'h422aa66f, 32'hc2a911e6, 32'h42a7f083, 32'h415ed20b, 32'hc2c6da6c, 32'hbf09a931, 32'hc1e3a103};
test_output[9200:9207] = '{32'h0, 32'h422aa66f, 32'h0, 32'h42a7f083, 32'h415ed20b, 32'h0, 32'h0, 32'h0};
test_input[9208:9215] = '{32'h4053232c, 32'hc19d8150, 32'hc267e9ae, 32'hc0053e1d, 32'hc15516b8, 32'h426a3b46, 32'h42a5f269, 32'h41e7e186};
test_output[9208:9215] = '{32'h4053232c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426a3b46, 32'h42a5f269, 32'h41e7e186};
test_input[9216:9223] = '{32'h428c9224, 32'h423f01e9, 32'hc299c018, 32'h429911b5, 32'h41339c56, 32'hc21bac5a, 32'h427352fd, 32'h4202ce28};
test_output[9216:9223] = '{32'h428c9224, 32'h423f01e9, 32'h0, 32'h429911b5, 32'h41339c56, 32'h0, 32'h427352fd, 32'h4202ce28};
test_input[9224:9231] = '{32'h425113ad, 32'hc2b76b99, 32'h413df6aa, 32'h42aa3646, 32'h41ba64af, 32'hc241951a, 32'hc1507ad0, 32'hc204d28a};
test_output[9224:9231] = '{32'h425113ad, 32'h0, 32'h413df6aa, 32'h42aa3646, 32'h41ba64af, 32'h0, 32'h0, 32'h0};
test_input[9232:9239] = '{32'h41fc8122, 32'hc2084962, 32'hc2072177, 32'hc2904fa9, 32'h42bbe6f3, 32'hc2904dbf, 32'hc2af9b99, 32'h4205cc0a};
test_output[9232:9239] = '{32'h41fc8122, 32'h0, 32'h0, 32'h0, 32'h42bbe6f3, 32'h0, 32'h0, 32'h4205cc0a};
test_input[9240:9247] = '{32'hc2b83701, 32'hc2b3a94a, 32'hc28d6d48, 32'hc249603a, 32'h42923917, 32'h42a75a92, 32'hc1cd9f15, 32'hc2b4af77};
test_output[9240:9247] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42923917, 32'h42a75a92, 32'h0, 32'h0};
test_input[9248:9255] = '{32'hc2a04922, 32'h427eab23, 32'h42931b26, 32'h41a5079d, 32'hc28a0fdc, 32'hc0f5074b, 32'h42058d5c, 32'h42c651ed};
test_output[9248:9255] = '{32'h0, 32'h427eab23, 32'h42931b26, 32'h41a5079d, 32'h0, 32'h0, 32'h42058d5c, 32'h42c651ed};
test_input[9256:9263] = '{32'hc2112a17, 32'hc21748ad, 32'hc2b51edf, 32'hc276b416, 32'hc12871f9, 32'h4237e014, 32'hc205ce51, 32'hc2b9466c};
test_output[9256:9263] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4237e014, 32'h0, 32'h0};
test_input[9264:9271] = '{32'hc059d3cb, 32'h420f8f9a, 32'hc28263a2, 32'hc2a54644, 32'hc1eb32f5, 32'hc2a28f5b, 32'h41fd4576, 32'h42668691};
test_output[9264:9271] = '{32'h0, 32'h420f8f9a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41fd4576, 32'h42668691};
test_input[9272:9279] = '{32'h42b4db82, 32'h427b253f, 32'h429c8af3, 32'hc21bd4b5, 32'hc1c8f8b9, 32'hc06119fe, 32'hc23dba36, 32'hc2c18df0};
test_output[9272:9279] = '{32'h42b4db82, 32'h427b253f, 32'h429c8af3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9280:9287] = '{32'hc1c8b2e8, 32'hc2a5351c, 32'hc2c6016b, 32'h42a0834c, 32'h4269e09e, 32'h41f1ca4e, 32'h428ab4fd, 32'h42378d85};
test_output[9280:9287] = '{32'h0, 32'h0, 32'h0, 32'h42a0834c, 32'h4269e09e, 32'h41f1ca4e, 32'h428ab4fd, 32'h42378d85};
test_input[9288:9295] = '{32'h425dacc6, 32'h42a59292, 32'hc1898b3c, 32'h40a6201e, 32'hc2935aee, 32'h42c6eff4, 32'h420fa59a, 32'h42708f66};
test_output[9288:9295] = '{32'h425dacc6, 32'h42a59292, 32'h0, 32'h40a6201e, 32'h0, 32'h42c6eff4, 32'h420fa59a, 32'h42708f66};
test_input[9296:9303] = '{32'h4279e2cc, 32'hc290c64c, 32'hc2be11ab, 32'h429d8b75, 32'h4240f8c2, 32'hc2a0015f, 32'hc1a265e9, 32'hc02f828e};
test_output[9296:9303] = '{32'h4279e2cc, 32'h0, 32'h0, 32'h429d8b75, 32'h4240f8c2, 32'h0, 32'h0, 32'h0};
test_input[9304:9311] = '{32'h42a04ed1, 32'hc1196c09, 32'h41c4cd3f, 32'hbf7bb38b, 32'hc2c45af9, 32'hc27c1de5, 32'h4233a503, 32'hc2a6c7de};
test_output[9304:9311] = '{32'h42a04ed1, 32'h0, 32'h41c4cd3f, 32'h0, 32'h0, 32'h0, 32'h4233a503, 32'h0};
test_input[9312:9319] = '{32'h413a1f6c, 32'h42473c19, 32'hc2a59248, 32'h40e72ca8, 32'h42c21c0d, 32'h4267966c, 32'h4269cad0, 32'h42b6808f};
test_output[9312:9319] = '{32'h413a1f6c, 32'h42473c19, 32'h0, 32'h40e72ca8, 32'h42c21c0d, 32'h4267966c, 32'h4269cad0, 32'h42b6808f};
test_input[9320:9327] = '{32'h426f1001, 32'h42c449fc, 32'hc212b8d3, 32'hc2aa04d5, 32'h414ce111, 32'hc2905251, 32'hc2777d32, 32'h428d8054};
test_output[9320:9327] = '{32'h426f1001, 32'h42c449fc, 32'h0, 32'h0, 32'h414ce111, 32'h0, 32'h0, 32'h428d8054};
test_input[9328:9335] = '{32'hc28b347f, 32'hc1ede13a, 32'h40659aac, 32'hc2502b45, 32'h41523616, 32'hc2a74173, 32'h4158888f, 32'hc2277866};
test_output[9328:9335] = '{32'h0, 32'h0, 32'h40659aac, 32'h0, 32'h41523616, 32'h0, 32'h4158888f, 32'h0};
test_input[9336:9343] = '{32'h418ccd2a, 32'hc298dd51, 32'h42c26475, 32'hc1719c92, 32'h4245d30c, 32'hc1e73906, 32'h4292c523, 32'hc160a259};
test_output[9336:9343] = '{32'h418ccd2a, 32'h0, 32'h42c26475, 32'h0, 32'h4245d30c, 32'h0, 32'h4292c523, 32'h0};
test_input[9344:9351] = '{32'hc1905bc1, 32'hc27ccce4, 32'h4284bcb4, 32'h41210f35, 32'h410b2bc2, 32'hc0fcedd5, 32'hc2366c6c, 32'h428716ad};
test_output[9344:9351] = '{32'h0, 32'h0, 32'h4284bcb4, 32'h41210f35, 32'h410b2bc2, 32'h0, 32'h0, 32'h428716ad};
test_input[9352:9359] = '{32'hc26fdb46, 32'h424388ad, 32'hc1542cb4, 32'h42153b47, 32'hc1a3ec83, 32'h42585059, 32'h4246c99d, 32'hc05291d9};
test_output[9352:9359] = '{32'h0, 32'h424388ad, 32'h0, 32'h42153b47, 32'h0, 32'h42585059, 32'h4246c99d, 32'h0};
test_input[9360:9367] = '{32'h40be09b4, 32'h42a7c82b, 32'h42a11fa6, 32'h42b150f0, 32'hc2a76141, 32'hc02c45ca, 32'hc2713424, 32'h42bbeb26};
test_output[9360:9367] = '{32'h40be09b4, 32'h42a7c82b, 32'h42a11fa6, 32'h42b150f0, 32'h0, 32'h0, 32'h0, 32'h42bbeb26};
test_input[9368:9375] = '{32'hc19e2216, 32'h426d6770, 32'h41dfafc8, 32'h42c4470e, 32'h4294f572, 32'h418b9aa1, 32'h42978074, 32'h42acf727};
test_output[9368:9375] = '{32'h0, 32'h426d6770, 32'h41dfafc8, 32'h42c4470e, 32'h4294f572, 32'h418b9aa1, 32'h42978074, 32'h42acf727};
test_input[9376:9383] = '{32'hc288bd72, 32'hc05f2565, 32'hc27cdd3b, 32'hc1926ba1, 32'h4094acb8, 32'h42401b07, 32'h429e90d2, 32'h42909a51};
test_output[9376:9383] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4094acb8, 32'h42401b07, 32'h429e90d2, 32'h42909a51};
test_input[9384:9391] = '{32'h42877550, 32'h428c52e2, 32'hc292764c, 32'h41c194f9, 32'hc2c43b01, 32'hc21eda81, 32'h422b9f5b, 32'h4226ad4d};
test_output[9384:9391] = '{32'h42877550, 32'h428c52e2, 32'h0, 32'h41c194f9, 32'h0, 32'h0, 32'h422b9f5b, 32'h4226ad4d};
test_input[9392:9399] = '{32'hc1a27522, 32'hc2c0cf0f, 32'h41f375bd, 32'hc21c1a32, 32'hc200ed91, 32'h426a9d6f, 32'h4131fe1d, 32'h42c5348d};
test_output[9392:9399] = '{32'h0, 32'h0, 32'h41f375bd, 32'h0, 32'h0, 32'h426a9d6f, 32'h4131fe1d, 32'h42c5348d};
test_input[9400:9407] = '{32'hc281db07, 32'hc22fe8ac, 32'h4295b0fb, 32'h42b6587d, 32'h42b4bf2d, 32'h427986e3, 32'h427ddec8, 32'hc25bf8de};
test_output[9400:9407] = '{32'h0, 32'h0, 32'h4295b0fb, 32'h42b6587d, 32'h42b4bf2d, 32'h427986e3, 32'h427ddec8, 32'h0};
test_input[9408:9415] = '{32'h426f2b92, 32'hc228623a, 32'h408e5d24, 32'h42c773e7, 32'hc254b65f, 32'hc2ad0d2d, 32'h42966448, 32'h42424496};
test_output[9408:9415] = '{32'h426f2b92, 32'h0, 32'h408e5d24, 32'h42c773e7, 32'h0, 32'h0, 32'h42966448, 32'h42424496};
test_input[9416:9423] = '{32'h412b5fc8, 32'h42866c5f, 32'hc28df0a6, 32'h42254e25, 32'hc296dd6a, 32'h415259f3, 32'h428df0c3, 32'h42691eea};
test_output[9416:9423] = '{32'h412b5fc8, 32'h42866c5f, 32'h0, 32'h42254e25, 32'h0, 32'h415259f3, 32'h428df0c3, 32'h42691eea};
test_input[9424:9431] = '{32'hc11391fc, 32'hc1539497, 32'hc1e109d8, 32'hc2c38fd7, 32'h42747ef0, 32'h423b2a08, 32'hc28a251b, 32'h419c0c84};
test_output[9424:9431] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42747ef0, 32'h423b2a08, 32'h0, 32'h419c0c84};
test_input[9432:9439] = '{32'hc25fb285, 32'hc2a9f9d1, 32'hc27984d6, 32'hc0df5b46, 32'h421ef398, 32'h41cc844f, 32'hc2a84880, 32'h3f522011};
test_output[9432:9439] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h421ef398, 32'h41cc844f, 32'h0, 32'h3f522011};
test_input[9440:9447] = '{32'h417edbea, 32'h412dcaf2, 32'hc22501ee, 32'h41d1a1e9, 32'h426995b2, 32'h423adfdf, 32'h42a85648, 32'hc1cadba3};
test_output[9440:9447] = '{32'h417edbea, 32'h412dcaf2, 32'h0, 32'h41d1a1e9, 32'h426995b2, 32'h423adfdf, 32'h42a85648, 32'h0};
test_input[9448:9455] = '{32'h42b4aca0, 32'hc2221278, 32'hc14f95f0, 32'hc088957f, 32'h4232df18, 32'hc2972087, 32'hc1bb67cc, 32'h428a1c61};
test_output[9448:9455] = '{32'h42b4aca0, 32'h0, 32'h0, 32'h0, 32'h4232df18, 32'h0, 32'h0, 32'h428a1c61};
test_input[9456:9463] = '{32'hc04358fd, 32'hc137e770, 32'h423b99ed, 32'h42a4c42a, 32'hc1991021, 32'h42abeadd, 32'h427db343, 32'hc1eaf197};
test_output[9456:9463] = '{32'h0, 32'h0, 32'h423b99ed, 32'h42a4c42a, 32'h0, 32'h42abeadd, 32'h427db343, 32'h0};
test_input[9464:9471] = '{32'hc1edecac, 32'hc2a4198c, 32'h42c4e475, 32'hc0fe790a, 32'h3fe2a831, 32'hc014f996, 32'h40a2d7c5, 32'h42478862};
test_output[9464:9471] = '{32'h0, 32'h0, 32'h42c4e475, 32'h0, 32'h3fe2a831, 32'h0, 32'h40a2d7c5, 32'h42478862};
test_input[9472:9479] = '{32'h4276a583, 32'hbfb2c20e, 32'h428f4d54, 32'hc22d6e27, 32'h429581cd, 32'h4274d7a5, 32'h42257941, 32'hc1bac106};
test_output[9472:9479] = '{32'h4276a583, 32'h0, 32'h428f4d54, 32'h0, 32'h429581cd, 32'h4274d7a5, 32'h42257941, 32'h0};
test_input[9480:9487] = '{32'h41e0fae1, 32'h41806815, 32'h41cbfea5, 32'h42381d4e, 32'hc2346f50, 32'h413e5c46, 32'hc1fd45c9, 32'h409bd913};
test_output[9480:9487] = '{32'h41e0fae1, 32'h41806815, 32'h41cbfea5, 32'h42381d4e, 32'h0, 32'h413e5c46, 32'h0, 32'h409bd913};
test_input[9488:9495] = '{32'h41e03611, 32'h42c16c46, 32'hc2b0ab4c, 32'h427ede0a, 32'hc27a3468, 32'hc23b18e7, 32'h420eb514, 32'h42a3cbe0};
test_output[9488:9495] = '{32'h41e03611, 32'h42c16c46, 32'h0, 32'h427ede0a, 32'h0, 32'h0, 32'h420eb514, 32'h42a3cbe0};
test_input[9496:9503] = '{32'hc082597a, 32'hc274093a, 32'hc117e793, 32'hc281420f, 32'h425d013a, 32'h41b4a71b, 32'h3cb155fb, 32'hc1e014ae};
test_output[9496:9503] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h425d013a, 32'h41b4a71b, 32'h3cb155fb, 32'h0};
test_input[9504:9511] = '{32'h42a69729, 32'h42a1e912, 32'hc29d662f, 32'h42c479c6, 32'hc249f785, 32'hc2be5bc2, 32'hc135ccaa, 32'hc25a0400};
test_output[9504:9511] = '{32'h42a69729, 32'h42a1e912, 32'h0, 32'h42c479c6, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9512:9519] = '{32'h412f0360, 32'h426a7189, 32'h41c8cb46, 32'h421279f1, 32'hc2c0135c, 32'h42b4a6ff, 32'hc19be01d, 32'hc1d7cacb};
test_output[9512:9519] = '{32'h412f0360, 32'h426a7189, 32'h41c8cb46, 32'h421279f1, 32'h0, 32'h42b4a6ff, 32'h0, 32'h0};
test_input[9520:9527] = '{32'h42c2ee07, 32'hc2614e5c, 32'h42a2be73, 32'h4283c87a, 32'hc240b6eb, 32'h428ebc09, 32'hc2845210, 32'h424abbcc};
test_output[9520:9527] = '{32'h42c2ee07, 32'h0, 32'h42a2be73, 32'h4283c87a, 32'h0, 32'h428ebc09, 32'h0, 32'h424abbcc};
test_input[9528:9535] = '{32'hc197366f, 32'hc2246a88, 32'hbfb68267, 32'hc29a38f0, 32'hc22e9781, 32'h42c4097c, 32'h425a046d, 32'h41d2656f};
test_output[9528:9535] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c4097c, 32'h425a046d, 32'h41d2656f};
test_input[9536:9543] = '{32'hc2864977, 32'hc272e868, 32'hc033a752, 32'h41d0211f, 32'h428892f3, 32'hc29852f9, 32'hc18d6a50, 32'h4296023c};
test_output[9536:9543] = '{32'h0, 32'h0, 32'h0, 32'h41d0211f, 32'h428892f3, 32'h0, 32'h0, 32'h4296023c};
test_input[9544:9551] = '{32'h4008155e, 32'hc2955e4e, 32'hc29d7f9e, 32'hc287e5c7, 32'h41ccd321, 32'h429211b9, 32'h42280783, 32'h42a3b334};
test_output[9544:9551] = '{32'h4008155e, 32'h0, 32'h0, 32'h0, 32'h41ccd321, 32'h429211b9, 32'h42280783, 32'h42a3b334};
test_input[9552:9559] = '{32'hc29408ec, 32'h42800552, 32'h42bdd269, 32'hc243d30f, 32'h426375db, 32'h42573f86, 32'h415e48aa, 32'h4285bd67};
test_output[9552:9559] = '{32'h0, 32'h42800552, 32'h42bdd269, 32'h0, 32'h426375db, 32'h42573f86, 32'h415e48aa, 32'h4285bd67};
test_input[9560:9567] = '{32'hc226a083, 32'h424e0a7c, 32'hc2b3cb38, 32'h4150a797, 32'hc2889ba6, 32'h415ce8ee, 32'h3fb4b8c0, 32'hc1c09937};
test_output[9560:9567] = '{32'h0, 32'h424e0a7c, 32'h0, 32'h4150a797, 32'h0, 32'h415ce8ee, 32'h3fb4b8c0, 32'h0};
test_input[9568:9575] = '{32'h429011d5, 32'hc1d98544, 32'h40926d0f, 32'h424c84aa, 32'h42318e3f, 32'h41553d2e, 32'h42492681, 32'hc1d634cd};
test_output[9568:9575] = '{32'h429011d5, 32'h0, 32'h40926d0f, 32'h424c84aa, 32'h42318e3f, 32'h41553d2e, 32'h42492681, 32'h0};
test_input[9576:9583] = '{32'hc170dda1, 32'hc2ba2f16, 32'h4195f063, 32'hc2c36b24, 32'hc10be5c1, 32'h41a5fa5b, 32'hc241923d, 32'h42403ba6};
test_output[9576:9583] = '{32'h0, 32'h0, 32'h4195f063, 32'h0, 32'h0, 32'h41a5fa5b, 32'h0, 32'h42403ba6};
test_input[9584:9591] = '{32'hc171a9cd, 32'h4211f7ce, 32'hc1868b92, 32'h414391e8, 32'hc1decdb8, 32'h42b1e61f, 32'hc10bf6f5, 32'h42be1268};
test_output[9584:9591] = '{32'h0, 32'h4211f7ce, 32'h0, 32'h414391e8, 32'h0, 32'h42b1e61f, 32'h0, 32'h42be1268};
test_input[9592:9599] = '{32'hc29daad5, 32'h42158978, 32'h4260f01a, 32'h4218a954, 32'hc1408360, 32'hc27ff384, 32'hc0ae435a, 32'h426a57ab};
test_output[9592:9599] = '{32'h0, 32'h42158978, 32'h4260f01a, 32'h4218a954, 32'h0, 32'h0, 32'h0, 32'h426a57ab};
test_input[9600:9607] = '{32'h426dab1d, 32'hc20309d6, 32'h421658db, 32'h42b7af58, 32'h42b9d1f8, 32'hc1c4d3a9, 32'h429bbbe1, 32'h42bec7bb};
test_output[9600:9607] = '{32'h426dab1d, 32'h0, 32'h421658db, 32'h42b7af58, 32'h42b9d1f8, 32'h0, 32'h429bbbe1, 32'h42bec7bb};
test_input[9608:9615] = '{32'h40395175, 32'h41f6458e, 32'h42541bd2, 32'hc18eae1d, 32'hc22a9b05, 32'hc293ab26, 32'h42980779, 32'h4256c19f};
test_output[9608:9615] = '{32'h40395175, 32'h41f6458e, 32'h42541bd2, 32'h0, 32'h0, 32'h0, 32'h42980779, 32'h4256c19f};
test_input[9616:9623] = '{32'h428f89b5, 32'hc238a8bb, 32'h424cb22f, 32'hc2b65f9c, 32'hc2aea2fa, 32'hc23498ce, 32'h420eb8a2, 32'hc139f85e};
test_output[9616:9623] = '{32'h428f89b5, 32'h0, 32'h424cb22f, 32'h0, 32'h0, 32'h0, 32'h420eb8a2, 32'h0};
test_input[9624:9631] = '{32'h42324e18, 32'h41cd4eda, 32'hc1751091, 32'hc2b87650, 32'hc20c4d8e, 32'h41131031, 32'h41800fcd, 32'h41292a40};
test_output[9624:9631] = '{32'h42324e18, 32'h41cd4eda, 32'h0, 32'h0, 32'h0, 32'h41131031, 32'h41800fcd, 32'h41292a40};
test_input[9632:9639] = '{32'hc2557e72, 32'h426fe9cc, 32'hc0d009af, 32'hc1aea3b6, 32'h42a3081d, 32'h4122e192, 32'h422ab40a, 32'h41760298};
test_output[9632:9639] = '{32'h0, 32'h426fe9cc, 32'h0, 32'h0, 32'h42a3081d, 32'h4122e192, 32'h422ab40a, 32'h41760298};
test_input[9640:9647] = '{32'hc20b64d9, 32'hc1f41ade, 32'hc24e694b, 32'hc209cebc, 32'h42a18d75, 32'h41c8c46e, 32'h4013afe5, 32'h41454154};
test_output[9640:9647] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a18d75, 32'h41c8c46e, 32'h4013afe5, 32'h41454154};
test_input[9648:9655] = '{32'hc23ec9ae, 32'hc267e317, 32'hc2ae153d, 32'hc2141a80, 32'h41a75a16, 32'hc20370e5, 32'hc21fb143, 32'hc0f15eb7};
test_output[9648:9655] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41a75a16, 32'h0, 32'h0, 32'h0};
test_input[9656:9663] = '{32'hc27eafe4, 32'h4265cdc8, 32'hc299ee8c, 32'h419132e6, 32'hc2c5bef7, 32'hc23944d8, 32'hc12a5249, 32'hc2934f81};
test_output[9656:9663] = '{32'h0, 32'h4265cdc8, 32'h0, 32'h419132e6, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9664:9671] = '{32'hc2281e67, 32'hc1cac6ac, 32'h429ceaa0, 32'h3ec4eb51, 32'hc207dbac, 32'h418e3f9b, 32'hc26172c0, 32'h42c0dfca};
test_output[9664:9671] = '{32'h0, 32'h0, 32'h429ceaa0, 32'h3ec4eb51, 32'h0, 32'h418e3f9b, 32'h0, 32'h42c0dfca};
test_input[9672:9679] = '{32'h4209e296, 32'h42710021, 32'hc2bb971a, 32'h41dc2ca1, 32'h4293e501, 32'h4295d63b, 32'hc28e1a99, 32'h412c59ff};
test_output[9672:9679] = '{32'h4209e296, 32'h42710021, 32'h0, 32'h41dc2ca1, 32'h4293e501, 32'h4295d63b, 32'h0, 32'h412c59ff};
test_input[9680:9687] = '{32'hc28c3ede, 32'hc2a6d978, 32'h42b54df3, 32'h41cffd43, 32'h42aefced, 32'h41bacef7, 32'h42b9485d, 32'hc1a606c9};
test_output[9680:9687] = '{32'h0, 32'h0, 32'h42b54df3, 32'h41cffd43, 32'h42aefced, 32'h41bacef7, 32'h42b9485d, 32'h0};
test_input[9688:9695] = '{32'h41156c87, 32'h41ce7e98, 32'hbe46b199, 32'h429e4a8b, 32'hc2543c30, 32'hc23d2a24, 32'hc2905a8c, 32'hc016a71d};
test_output[9688:9695] = '{32'h41156c87, 32'h41ce7e98, 32'h0, 32'h429e4a8b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9696:9703] = '{32'h417430b6, 32'h425fbbf8, 32'hc2a51ff8, 32'h41c6a0ed, 32'h42bf8046, 32'h4298fc7b, 32'hc2604d77, 32'hc1ef8fb8};
test_output[9696:9703] = '{32'h417430b6, 32'h425fbbf8, 32'h0, 32'h41c6a0ed, 32'h42bf8046, 32'h4298fc7b, 32'h0, 32'h0};
test_input[9704:9711] = '{32'h424c8917, 32'h4230b5f9, 32'h426e7037, 32'h41f5c637, 32'h42187674, 32'hc1d31519, 32'hc20421c2, 32'h42404551};
test_output[9704:9711] = '{32'h424c8917, 32'h4230b5f9, 32'h426e7037, 32'h41f5c637, 32'h42187674, 32'h0, 32'h0, 32'h42404551};
test_input[9712:9719] = '{32'hc1717a96, 32'h42258425, 32'h41fc5141, 32'h41eafb47, 32'h4297c835, 32'h40158b3a, 32'h420f8027, 32'hbfc6d8d0};
test_output[9712:9719] = '{32'h0, 32'h42258425, 32'h41fc5141, 32'h41eafb47, 32'h4297c835, 32'h40158b3a, 32'h420f8027, 32'h0};
test_input[9720:9727] = '{32'hc2b9fe3d, 32'hc2c174ee, 32'hc28c8b35, 32'hc1c8659a, 32'hc1455801, 32'hc1352639, 32'hc0f5c8e7, 32'hc29f3542};
test_output[9720:9727] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9728:9735] = '{32'h426503ab, 32'hc0420e9a, 32'hc25038db, 32'h4150d8e0, 32'hc2b206a7, 32'h426ed520, 32'h40bc3513, 32'hc2b06d89};
test_output[9728:9735] = '{32'h426503ab, 32'h0, 32'h0, 32'h4150d8e0, 32'h0, 32'h426ed520, 32'h40bc3513, 32'h0};
test_input[9736:9743] = '{32'h429b0ec4, 32'h42bfddb6, 32'h42374049, 32'h42575a86, 32'h42a2b657, 32'h41a264c0, 32'h423ef37b, 32'hbfd3f2ce};
test_output[9736:9743] = '{32'h429b0ec4, 32'h42bfddb6, 32'h42374049, 32'h42575a86, 32'h42a2b657, 32'h41a264c0, 32'h423ef37b, 32'h0};
test_input[9744:9751] = '{32'hc2a40688, 32'h424e14c4, 32'h4152417b, 32'h4183bf2e, 32'hc205c904, 32'h423d667c, 32'h428a462f, 32'h422d3824};
test_output[9744:9751] = '{32'h0, 32'h424e14c4, 32'h4152417b, 32'h4183bf2e, 32'h0, 32'h423d667c, 32'h428a462f, 32'h422d3824};
test_input[9752:9759] = '{32'hc2a6279f, 32'h42629e3b, 32'h42815553, 32'hc1ff6a16, 32'h41f3e192, 32'hc253d3c3, 32'h42987094, 32'h420230cb};
test_output[9752:9759] = '{32'h0, 32'h42629e3b, 32'h42815553, 32'h0, 32'h41f3e192, 32'h0, 32'h42987094, 32'h420230cb};
test_input[9760:9767] = '{32'h42925b9d, 32'h421ee6c3, 32'hc17bb580, 32'h4274271d, 32'h4185a8ff, 32'h41a2d017, 32'hc2189dc4, 32'h421d6a6a};
test_output[9760:9767] = '{32'h42925b9d, 32'h421ee6c3, 32'h0, 32'h4274271d, 32'h4185a8ff, 32'h41a2d017, 32'h0, 32'h421d6a6a};
test_input[9768:9775] = '{32'hc203b6e5, 32'h40045f69, 32'h42b98d1e, 32'hc18e70c9, 32'h423ea7e7, 32'h41c1b805, 32'hc2a2bc83, 32'hc1ce4955};
test_output[9768:9775] = '{32'h0, 32'h40045f69, 32'h42b98d1e, 32'h0, 32'h423ea7e7, 32'h41c1b805, 32'h0, 32'h0};
test_input[9776:9783] = '{32'hc203c046, 32'hc2b8fd6e, 32'h426408cc, 32'h42577556, 32'hc13df735, 32'h423dc645, 32'h4293980b, 32'hc289b56c};
test_output[9776:9783] = '{32'h0, 32'h0, 32'h426408cc, 32'h42577556, 32'h0, 32'h423dc645, 32'h4293980b, 32'h0};
test_input[9784:9791] = '{32'h41b5bdb3, 32'hc25d8573, 32'h41eecdf8, 32'h4259bc9e, 32'h40cd08ec, 32'hc2222bbf, 32'hc2c48b14, 32'h42a52f05};
test_output[9784:9791] = '{32'h41b5bdb3, 32'h0, 32'h41eecdf8, 32'h4259bc9e, 32'h40cd08ec, 32'h0, 32'h0, 32'h42a52f05};
test_input[9792:9799] = '{32'hc2b12628, 32'hc23888c0, 32'hc2688cb1, 32'hc2635537, 32'hc0de4cab, 32'hc21f2d0c, 32'hc18be907, 32'hc24b2b15};
test_output[9792:9799] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[9800:9807] = '{32'h41a958bc, 32'hc1697f41, 32'h42758223, 32'hc0912fe2, 32'h402ccefd, 32'hc273b358, 32'h4297ecbd, 32'h428decc3};
test_output[9800:9807] = '{32'h41a958bc, 32'h0, 32'h42758223, 32'h0, 32'h402ccefd, 32'h0, 32'h4297ecbd, 32'h428decc3};
test_input[9808:9815] = '{32'h42b8e31c, 32'h4263a7b3, 32'h42641338, 32'hc20d6a52, 32'hc2a5de89, 32'hc27f720e, 32'h429a14a5, 32'h42bac256};
test_output[9808:9815] = '{32'h42b8e31c, 32'h4263a7b3, 32'h42641338, 32'h0, 32'h0, 32'h0, 32'h429a14a5, 32'h42bac256};
test_input[9816:9823] = '{32'h422c030f, 32'h42accaae, 32'h41ae0808, 32'hc1a38995, 32'hc271a84a, 32'hc29a9f89, 32'h425f3cea, 32'h42010adb};
test_output[9816:9823] = '{32'h422c030f, 32'h42accaae, 32'h41ae0808, 32'h0, 32'h0, 32'h0, 32'h425f3cea, 32'h42010adb};
test_input[9824:9831] = '{32'hc2b856d3, 32'hc25537c2, 32'h424ed640, 32'hc24f65c4, 32'h420e43a7, 32'hc28dc123, 32'hc178f616, 32'h41b76fe5};
test_output[9824:9831] = '{32'h0, 32'h0, 32'h424ed640, 32'h0, 32'h420e43a7, 32'h0, 32'h0, 32'h41b76fe5};
test_input[9832:9839] = '{32'hc28ab97b, 32'h42b72ca7, 32'h421785e7, 32'hc28ec57f, 32'hc1173243, 32'hc29af924, 32'hc24ac18a, 32'h42109c92};
test_output[9832:9839] = '{32'h0, 32'h42b72ca7, 32'h421785e7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42109c92};
test_input[9840:9847] = '{32'h42b06b09, 32'hc27c2197, 32'h42ab3d6b, 32'hc29da7f4, 32'h4298ff54, 32'hc237803b, 32'h42b23109, 32'h4218a95a};
test_output[9840:9847] = '{32'h42b06b09, 32'h0, 32'h42ab3d6b, 32'h0, 32'h4298ff54, 32'h0, 32'h42b23109, 32'h4218a95a};
test_input[9848:9855] = '{32'hc1fe0b35, 32'hc2028b74, 32'hc068b086, 32'hc14224d9, 32'hc1179cc6, 32'h425b4977, 32'hc1f80010, 32'h42a59694};
test_output[9848:9855] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425b4977, 32'h0, 32'h42a59694};
test_input[9856:9863] = '{32'h3fb5c19e, 32'hc29227f3, 32'h4206a31e, 32'hc2b3832a, 32'h40a92170, 32'h4215e330, 32'hc2938621, 32'hc1c3c8e2};
test_output[9856:9863] = '{32'h3fb5c19e, 32'h0, 32'h4206a31e, 32'h0, 32'h40a92170, 32'h4215e330, 32'h0, 32'h0};
test_input[9864:9871] = '{32'h42b7f05c, 32'hc1d39d28, 32'hc2a4278f, 32'h420b067c, 32'h42bb3576, 32'h4131fa9a, 32'hc2b8c40d, 32'hc1c09533};
test_output[9864:9871] = '{32'h42b7f05c, 32'h0, 32'h0, 32'h420b067c, 32'h42bb3576, 32'h4131fa9a, 32'h0, 32'h0};
test_input[9872:9879] = '{32'hc0b483e8, 32'h428619df, 32'h429aa6e4, 32'hc2ae207f, 32'h42755040, 32'h42a81ee3, 32'hc22ea8a6, 32'h4006bf92};
test_output[9872:9879] = '{32'h0, 32'h428619df, 32'h429aa6e4, 32'h0, 32'h42755040, 32'h42a81ee3, 32'h0, 32'h4006bf92};
test_input[9880:9887] = '{32'hc21a950a, 32'h41b1a195, 32'hc27fa083, 32'h42a29eb2, 32'h41eddde4, 32'h4174703f, 32'h40326686, 32'hc290461a};
test_output[9880:9887] = '{32'h0, 32'h41b1a195, 32'h0, 32'h42a29eb2, 32'h41eddde4, 32'h4174703f, 32'h40326686, 32'h0};
test_input[9888:9895] = '{32'hc258880b, 32'h42831687, 32'hc2941321, 32'h415e7464, 32'hc2a20605, 32'h41080106, 32'hc208cf6e, 32'h41fd492b};
test_output[9888:9895] = '{32'h0, 32'h42831687, 32'h0, 32'h415e7464, 32'h0, 32'h41080106, 32'h0, 32'h41fd492b};
test_input[9896:9903] = '{32'h42ae918c, 32'h421c6d7a, 32'hc1fc21c3, 32'h41f88332, 32'hc2bd7a41, 32'h42c32c44, 32'h416367a4, 32'h42b31114};
test_output[9896:9903] = '{32'h42ae918c, 32'h421c6d7a, 32'h0, 32'h41f88332, 32'h0, 32'h42c32c44, 32'h416367a4, 32'h42b31114};
test_input[9904:9911] = '{32'hc1f09d6a, 32'h428fe967, 32'h41a64f7a, 32'h4114a848, 32'h42b9c810, 32'h42be9ab7, 32'h428b7dc4, 32'hc2ba5e75};
test_output[9904:9911] = '{32'h0, 32'h428fe967, 32'h41a64f7a, 32'h4114a848, 32'h42b9c810, 32'h42be9ab7, 32'h428b7dc4, 32'h0};
test_input[9912:9919] = '{32'hc1c70d13, 32'hc267eeae, 32'h422566d9, 32'h42c0c6b8, 32'h41c7427b, 32'h42b48648, 32'h418112c6, 32'h4248e012};
test_output[9912:9919] = '{32'h0, 32'h0, 32'h422566d9, 32'h42c0c6b8, 32'h41c7427b, 32'h42b48648, 32'h418112c6, 32'h4248e012};
test_input[9920:9927] = '{32'hc03d1069, 32'hc246716b, 32'hc2775b9b, 32'hc17ca427, 32'hc2b14919, 32'h41bcf170, 32'h42346a2c, 32'h429ddd8f};
test_output[9920:9927] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41bcf170, 32'h42346a2c, 32'h429ddd8f};
test_input[9928:9935] = '{32'h429f47ab, 32'hc2c15558, 32'h42859932, 32'h4187e8e1, 32'h42738e0d, 32'hc1828814, 32'hc2a21aa2, 32'hc18da3fe};
test_output[9928:9935] = '{32'h429f47ab, 32'h0, 32'h42859932, 32'h4187e8e1, 32'h42738e0d, 32'h0, 32'h0, 32'h0};
test_input[9936:9943] = '{32'hc127615f, 32'hc2475821, 32'hc296eec4, 32'h41ff14b0, 32'hc2c07130, 32'hc24cd249, 32'h42a61e2f, 32'h422e453a};
test_output[9936:9943] = '{32'h0, 32'h0, 32'h0, 32'h41ff14b0, 32'h0, 32'h0, 32'h42a61e2f, 32'h422e453a};
test_input[9944:9951] = '{32'hc28ef41d, 32'hc02dece4, 32'h4288e698, 32'hc28aa5aa, 32'h4272e1eb, 32'hc2253877, 32'h42c706a7, 32'h4280c973};
test_output[9944:9951] = '{32'h0, 32'h0, 32'h4288e698, 32'h0, 32'h4272e1eb, 32'h0, 32'h42c706a7, 32'h4280c973};
test_input[9952:9959] = '{32'hc28dca09, 32'hc12eadd9, 32'h42b8c305, 32'h4281c993, 32'h42811ab1, 32'h41014836, 32'hc1e89841, 32'hc1a89ae2};
test_output[9952:9959] = '{32'h0, 32'h0, 32'h42b8c305, 32'h4281c993, 32'h42811ab1, 32'h41014836, 32'h0, 32'h0};
test_input[9960:9967] = '{32'hc1e6149f, 32'hc280a902, 32'h417b465f, 32'h429c76dd, 32'hc231df5e, 32'hc2547f79, 32'hc2a182e4, 32'h41429e43};
test_output[9960:9967] = '{32'h0, 32'h0, 32'h417b465f, 32'h429c76dd, 32'h0, 32'h0, 32'h0, 32'h41429e43};
test_input[9968:9975] = '{32'hc23c13f7, 32'h42b873af, 32'h4260ee2b, 32'h4232be88, 32'hc1932588, 32'h41116dfb, 32'h42b9798a, 32'hc1ac82f4};
test_output[9968:9975] = '{32'h0, 32'h42b873af, 32'h4260ee2b, 32'h4232be88, 32'h0, 32'h41116dfb, 32'h42b9798a, 32'h0};
test_input[9976:9983] = '{32'h42788c98, 32'hc20b9277, 32'hc227ede4, 32'hc192a8b8, 32'h4148ce60, 32'h42253ac0, 32'h421ed00e, 32'hc2b7437c};
test_output[9976:9983] = '{32'h42788c98, 32'h0, 32'h0, 32'h0, 32'h4148ce60, 32'h42253ac0, 32'h421ed00e, 32'h0};
test_input[9984:9991] = '{32'h42657cd9, 32'hc14e328b, 32'h42652895, 32'hc10240ba, 32'hc22880bc, 32'h3fc27c05, 32'hc1cfe1dc, 32'h42123370};
test_output[9984:9991] = '{32'h42657cd9, 32'h0, 32'h42652895, 32'h0, 32'h0, 32'h3fc27c05, 32'h0, 32'h42123370};
test_input[9992:9999] = '{32'hc25c89fb, 32'hc2715ebd, 32'h4244b99b, 32'hc28271e8, 32'h427f42b2, 32'hc2be0fca, 32'hc1ac2951, 32'hc27fa2ae};
test_output[9992:9999] = '{32'h0, 32'h0, 32'h4244b99b, 32'h0, 32'h427f42b2, 32'h0, 32'h0, 32'h0};
test_input[10000:10007] = '{32'h41a85b86, 32'hc1ad636e, 32'hc269b82b, 32'hc28be09c, 32'hc298e769, 32'h408b8d5e, 32'h420a5066, 32'hc2a106dd};
test_output[10000:10007] = '{32'h41a85b86, 32'h0, 32'h0, 32'h0, 32'h0, 32'h408b8d5e, 32'h420a5066, 32'h0};
test_input[10008:10015] = '{32'hc1881ca9, 32'hc13bb1cc, 32'h429d6878, 32'h41ea995b, 32'h428384ba, 32'h413cf086, 32'hc2350169, 32'h42b3fbb8};
test_output[10008:10015] = '{32'h0, 32'h0, 32'h429d6878, 32'h41ea995b, 32'h428384ba, 32'h413cf086, 32'h0, 32'h42b3fbb8};
test_input[10016:10023] = '{32'hc20da047, 32'h42892159, 32'h42701279, 32'h42893139, 32'hc2c07a98, 32'hc268eb22, 32'h41c8a5c2, 32'h42b74bfe};
test_output[10016:10023] = '{32'h0, 32'h42892159, 32'h42701279, 32'h42893139, 32'h0, 32'h0, 32'h41c8a5c2, 32'h42b74bfe};
test_input[10024:10031] = '{32'hc2ab4512, 32'hc250ba40, 32'hc1aa8fb2, 32'hc1e3fc98, 32'hc1f3e2a5, 32'h4181431b, 32'hc15ed16b, 32'hc16ba4b1};
test_output[10024:10031] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4181431b, 32'h0, 32'h0};
test_input[10032:10039] = '{32'h4212d9a2, 32'hc2a3efc9, 32'hc0792813, 32'hc23ab478, 32'h420e6b63, 32'h42c3537c, 32'hc2b6aad5, 32'h3e86937b};
test_output[10032:10039] = '{32'h4212d9a2, 32'h0, 32'h0, 32'h0, 32'h420e6b63, 32'h42c3537c, 32'h0, 32'h3e86937b};
test_input[10040:10047] = '{32'hc29814c5, 32'h4254e957, 32'hc26075ac, 32'hc247d032, 32'hc0e3d0a3, 32'hc29b4eed, 32'h42984b57, 32'hc24db7e4};
test_output[10040:10047] = '{32'h0, 32'h4254e957, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42984b57, 32'h0};
test_input[10048:10055] = '{32'h42524219, 32'hc26905ca, 32'h4286ba1c, 32'hc1d1f5e8, 32'h42847b08, 32'h42746c0c, 32'h41a846f3, 32'hc2815de6};
test_output[10048:10055] = '{32'h42524219, 32'h0, 32'h4286ba1c, 32'h0, 32'h42847b08, 32'h42746c0c, 32'h41a846f3, 32'h0};
test_input[10056:10063] = '{32'h421015f2, 32'h41b19017, 32'hc267ae1f, 32'hc2a33126, 32'h42b00f32, 32'h40c11de2, 32'hc2735530, 32'hc16014d3};
test_output[10056:10063] = '{32'h421015f2, 32'h41b19017, 32'h0, 32'h0, 32'h42b00f32, 32'h40c11de2, 32'h0, 32'h0};
test_input[10064:10071] = '{32'h429d188e, 32'h42bccc43, 32'hc2989603, 32'hc0cccf87, 32'h42c6e703, 32'h42969586, 32'hc206ab8d, 32'hc217107e};
test_output[10064:10071] = '{32'h429d188e, 32'h42bccc43, 32'h0, 32'h0, 32'h42c6e703, 32'h42969586, 32'h0, 32'h0};
test_input[10072:10079] = '{32'hc2268340, 32'h422fec3d, 32'hc0c61ad3, 32'hc24ded99, 32'hc28c0b69, 32'h42258e93, 32'h41a9ba2e, 32'h428281bb};
test_output[10072:10079] = '{32'h0, 32'h422fec3d, 32'h0, 32'h0, 32'h0, 32'h42258e93, 32'h41a9ba2e, 32'h428281bb};
test_input[10080:10087] = '{32'h41fca544, 32'h41a66a35, 32'h42bceff0, 32'h429ea857, 32'hc0f38a89, 32'hc1dae248, 32'h429fc8e3, 32'h42b57676};
test_output[10080:10087] = '{32'h41fca544, 32'h41a66a35, 32'h42bceff0, 32'h429ea857, 32'h0, 32'h0, 32'h429fc8e3, 32'h42b57676};
test_input[10088:10095] = '{32'h42c1b88e, 32'h4194a46e, 32'hc28caa50, 32'hc2b9e8a5, 32'h420b4b54, 32'h41e003de, 32'hc1b0197d, 32'hc22276fd};
test_output[10088:10095] = '{32'h42c1b88e, 32'h4194a46e, 32'h0, 32'h0, 32'h420b4b54, 32'h41e003de, 32'h0, 32'h0};
test_input[10096:10103] = '{32'hc2475a75, 32'hc203e644, 32'h425b9f04, 32'hc2c073e3, 32'h423d1bfe, 32'h42b4ec81, 32'hc2829375, 32'h4267f270};
test_output[10096:10103] = '{32'h0, 32'h0, 32'h425b9f04, 32'h0, 32'h423d1bfe, 32'h42b4ec81, 32'h0, 32'h4267f270};
test_input[10104:10111] = '{32'h42a29c8b, 32'h42be4eff, 32'hc280be02, 32'h428ac476, 32'hc2c4881a, 32'hc25ec1e5, 32'h4292a770, 32'hc2c7adda};
test_output[10104:10111] = '{32'h42a29c8b, 32'h42be4eff, 32'h0, 32'h428ac476, 32'h0, 32'h0, 32'h4292a770, 32'h0};
test_input[10112:10119] = '{32'h42922d88, 32'h41c149e3, 32'hc0994388, 32'h42a11021, 32'hc0767c49, 32'h41f6196b, 32'h425391d3, 32'h4081a20c};
test_output[10112:10119] = '{32'h42922d88, 32'h41c149e3, 32'h0, 32'h42a11021, 32'h0, 32'h41f6196b, 32'h425391d3, 32'h4081a20c};
test_input[10120:10127] = '{32'hc2955866, 32'h42b168d7, 32'hc28090f2, 32'hc28e5d86, 32'h3fcd8f95, 32'h41517439, 32'h41d89b3d, 32'hc2038b63};
test_output[10120:10127] = '{32'h0, 32'h42b168d7, 32'h0, 32'h0, 32'h3fcd8f95, 32'h41517439, 32'h41d89b3d, 32'h0};
test_input[10128:10135] = '{32'hc22d7ead, 32'h42a9357d, 32'hc27f28f2, 32'h42a2e377, 32'hc23c8046, 32'h42a4db1b, 32'hc29a524b, 32'hc252fc2f};
test_output[10128:10135] = '{32'h0, 32'h42a9357d, 32'h0, 32'h42a2e377, 32'h0, 32'h42a4db1b, 32'h0, 32'h0};
test_input[10136:10143] = '{32'h3f07462c, 32'hbf5281f7, 32'hc213ccaa, 32'hc1779e41, 32'hc0e487ac, 32'h4282d030, 32'hc29a70a0, 32'hc11f106d};
test_output[10136:10143] = '{32'h3f07462c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4282d030, 32'h0, 32'h0};
test_input[10144:10151] = '{32'h40199e2c, 32'hc2081642, 32'h42b60f58, 32'h4269f6ee, 32'hc27d0273, 32'hc2a755b4, 32'hc1cdfc14, 32'h42930755};
test_output[10144:10151] = '{32'h40199e2c, 32'h0, 32'h42b60f58, 32'h4269f6ee, 32'h0, 32'h0, 32'h0, 32'h42930755};
test_input[10152:10159] = '{32'h42b1fc11, 32'h41a1bd90, 32'h421a0556, 32'h422e77b0, 32'hc171efef, 32'h42587dc4, 32'hc23cde72, 32'hc11399aa};
test_output[10152:10159] = '{32'h42b1fc11, 32'h41a1bd90, 32'h421a0556, 32'h422e77b0, 32'h0, 32'h42587dc4, 32'h0, 32'h0};
test_input[10160:10167] = '{32'hc1f92e5e, 32'h41ccdc0e, 32'h421c104f, 32'hc21c2128, 32'h42b23a41, 32'hc13c8ef8, 32'hc203585b, 32'hc29d037b};
test_output[10160:10167] = '{32'h0, 32'h41ccdc0e, 32'h421c104f, 32'h0, 32'h42b23a41, 32'h0, 32'h0, 32'h0};
test_input[10168:10175] = '{32'h42578c2e, 32'h41e13a6d, 32'hc2bf4cb5, 32'hc2aa2686, 32'hc28a4f21, 32'h42b7ad72, 32'h4130a0d2, 32'h42a080cf};
test_output[10168:10175] = '{32'h42578c2e, 32'h41e13a6d, 32'h0, 32'h0, 32'h0, 32'h42b7ad72, 32'h4130a0d2, 32'h42a080cf};
test_input[10176:10183] = '{32'h41f867ba, 32'hc14ebec6, 32'h41385f27, 32'hc29b2799, 32'h42300ed7, 32'h420b89e8, 32'h41082a93, 32'hc1bcec3a};
test_output[10176:10183] = '{32'h41f867ba, 32'h0, 32'h41385f27, 32'h0, 32'h42300ed7, 32'h420b89e8, 32'h41082a93, 32'h0};
test_input[10184:10191] = '{32'h421a6a94, 32'h4191da7e, 32'h41b9ea7a, 32'hc21ec942, 32'h4251af98, 32'hc29f517b, 32'h429b2dd4, 32'h41ed4001};
test_output[10184:10191] = '{32'h421a6a94, 32'h4191da7e, 32'h41b9ea7a, 32'h0, 32'h4251af98, 32'h0, 32'h429b2dd4, 32'h41ed4001};
test_input[10192:10199] = '{32'h419457bc, 32'h41f77ce8, 32'h420c920d, 32'h41043e03, 32'h42b52536, 32'h41cd20fb, 32'h428fbd9b, 32'h4280d76f};
test_output[10192:10199] = '{32'h419457bc, 32'h41f77ce8, 32'h420c920d, 32'h41043e03, 32'h42b52536, 32'h41cd20fb, 32'h428fbd9b, 32'h4280d76f};
test_input[10200:10207] = '{32'h42c3c110, 32'h42c6489d, 32'h42b63a99, 32'hc13194e0, 32'h40654af0, 32'hc2abf187, 32'hc2832472, 32'hc29de752};
test_output[10200:10207] = '{32'h42c3c110, 32'h42c6489d, 32'h42b63a99, 32'h0, 32'h40654af0, 32'h0, 32'h0, 32'h0};
test_input[10208:10215] = '{32'h42873588, 32'hc1c915c2, 32'h41f566e5, 32'hc04057b6, 32'h42b899de, 32'h42783250, 32'hc225b79c, 32'hc2ae6400};
test_output[10208:10215] = '{32'h42873588, 32'h0, 32'h41f566e5, 32'h0, 32'h42b899de, 32'h42783250, 32'h0, 32'h0};
test_input[10216:10223] = '{32'hc2a886da, 32'hc24c60bb, 32'h425cbfc2, 32'h42821dc9, 32'h428edd1b, 32'hc2829b37, 32'h42c2c30c, 32'h408366c7};
test_output[10216:10223] = '{32'h0, 32'h0, 32'h425cbfc2, 32'h42821dc9, 32'h428edd1b, 32'h0, 32'h42c2c30c, 32'h408366c7};
test_input[10224:10231] = '{32'hc28c721d, 32'h42599ba7, 32'hc0ae2bd1, 32'hc278aab2, 32'h428774f9, 32'hc04e9102, 32'hc2314e18, 32'h42693ec5};
test_output[10224:10231] = '{32'h0, 32'h42599ba7, 32'h0, 32'h0, 32'h428774f9, 32'h0, 32'h0, 32'h42693ec5};
test_input[10232:10239] = '{32'h41d0d6e9, 32'hc2851c52, 32'hc0ebe44b, 32'h422951a5, 32'h41973112, 32'hc104302c, 32'h4148b5de, 32'h41f6e45e};
test_output[10232:10239] = '{32'h41d0d6e9, 32'h0, 32'h0, 32'h422951a5, 32'h41973112, 32'h0, 32'h4148b5de, 32'h41f6e45e};
test_input[10240:10247] = '{32'h42bfe7dd, 32'hc1acc7f8, 32'h42c31e19, 32'hc0ec21a4, 32'h4295be2a, 32'hc2c6137d, 32'h42972826, 32'hc25181a4};
test_output[10240:10247] = '{32'h42bfe7dd, 32'h0, 32'h42c31e19, 32'h0, 32'h4295be2a, 32'h0, 32'h42972826, 32'h0};
test_input[10248:10255] = '{32'hc2b69e3f, 32'h421c41dd, 32'h427a647a, 32'hc28603dc, 32'hc2ab4811, 32'hc235a478, 32'h41c75334, 32'h42527522};
test_output[10248:10255] = '{32'h0, 32'h421c41dd, 32'h427a647a, 32'h0, 32'h0, 32'h0, 32'h41c75334, 32'h42527522};
test_input[10256:10263] = '{32'hc294c4b7, 32'hc2980376, 32'hc2adf79b, 32'h422e066c, 32'h415a02e6, 32'h410f9931, 32'h4259c2e5, 32'h4240dbc3};
test_output[10256:10263] = '{32'h0, 32'h0, 32'h0, 32'h422e066c, 32'h415a02e6, 32'h410f9931, 32'h4259c2e5, 32'h4240dbc3};
test_input[10264:10271] = '{32'h4133fd5e, 32'h42b7b1d8, 32'h41608d28, 32'h42c6fb9c, 32'hc18a3189, 32'h42b65def, 32'h42c4a132, 32'hc1d65dda};
test_output[10264:10271] = '{32'h4133fd5e, 32'h42b7b1d8, 32'h41608d28, 32'h42c6fb9c, 32'h0, 32'h42b65def, 32'h42c4a132, 32'h0};
test_input[10272:10279] = '{32'h4187b4b1, 32'h418562c6, 32'hc0c06000, 32'hc2a0ff22, 32'h42419024, 32'hc2023a4a, 32'hc2979237, 32'hc24488b4};
test_output[10272:10279] = '{32'h4187b4b1, 32'h418562c6, 32'h0, 32'h0, 32'h42419024, 32'h0, 32'h0, 32'h0};
test_input[10280:10287] = '{32'hc25a0762, 32'h427c2f8e, 32'h428319f9, 32'hc2408c84, 32'h421092f9, 32'hc0fc0257, 32'hc2bae5d9, 32'h4293ffbe};
test_output[10280:10287] = '{32'h0, 32'h427c2f8e, 32'h428319f9, 32'h0, 32'h421092f9, 32'h0, 32'h0, 32'h4293ffbe};
test_input[10288:10295] = '{32'hc2b5a343, 32'hc289c1c4, 32'hc2a7c1aa, 32'hc27b2e50, 32'hc167f42c, 32'h411f90a2, 32'hc27aba60, 32'h42a55f43};
test_output[10288:10295] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h411f90a2, 32'h0, 32'h42a55f43};
test_input[10296:10303] = '{32'hc1a20091, 32'h42a2548f, 32'hc2bd70bb, 32'h41c26e9e, 32'hc21033c6, 32'hc2c424bf, 32'h428f1633, 32'hc2acd203};
test_output[10296:10303] = '{32'h0, 32'h42a2548f, 32'h0, 32'h41c26e9e, 32'h0, 32'h0, 32'h428f1633, 32'h0};
test_input[10304:10311] = '{32'hc2823058, 32'h41e11d53, 32'hc27dcbd9, 32'hc2a12b86, 32'h42aa5de5, 32'h42660255, 32'hc1260bbb, 32'h428fafbd};
test_output[10304:10311] = '{32'h0, 32'h41e11d53, 32'h0, 32'h0, 32'h42aa5de5, 32'h42660255, 32'h0, 32'h428fafbd};
test_input[10312:10319] = '{32'hc26f97df, 32'h428689cb, 32'hc21cfeb4, 32'h41992898, 32'hc1d9413f, 32'h428e50dc, 32'hc22a521d, 32'hc101a24c};
test_output[10312:10319] = '{32'h0, 32'h428689cb, 32'h0, 32'h41992898, 32'h0, 32'h428e50dc, 32'h0, 32'h0};
test_input[10320:10327] = '{32'h422b0f1b, 32'hc1cb09a9, 32'h40a45fab, 32'hc28e29bb, 32'hc19fa5c6, 32'hc2ba1283, 32'hc296f180, 32'h41738d4a};
test_output[10320:10327] = '{32'h422b0f1b, 32'h0, 32'h40a45fab, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41738d4a};
test_input[10328:10335] = '{32'h42bfadb0, 32'h42aacaf7, 32'h42931f1b, 32'hc295d9ff, 32'hc2252f43, 32'h427865a1, 32'h424e6e73, 32'h40a93eb3};
test_output[10328:10335] = '{32'h42bfadb0, 32'h42aacaf7, 32'h42931f1b, 32'h0, 32'h0, 32'h427865a1, 32'h424e6e73, 32'h40a93eb3};
test_input[10336:10343] = '{32'h423a7e34, 32'hc1342c51, 32'h41aa38c4, 32'h42bc790f, 32'hc22fcdf0, 32'hc20b8c60, 32'hc2b4b986, 32'h42bc10d4};
test_output[10336:10343] = '{32'h423a7e34, 32'h0, 32'h41aa38c4, 32'h42bc790f, 32'h0, 32'h0, 32'h0, 32'h42bc10d4};
test_input[10344:10351] = '{32'hc201a366, 32'h42886730, 32'h42c1ef5e, 32'hc29538b1, 32'hc1cfb579, 32'hc218462a, 32'h42c59aa2, 32'hc1189767};
test_output[10344:10351] = '{32'h0, 32'h42886730, 32'h42c1ef5e, 32'h0, 32'h0, 32'h0, 32'h42c59aa2, 32'h0};
test_input[10352:10359] = '{32'h42c7d141, 32'hc220072f, 32'h4100177e, 32'hc0369b66, 32'hc22574a9, 32'hc1ba9e53, 32'h428c6dda, 32'h41ed5e6f};
test_output[10352:10359] = '{32'h42c7d141, 32'h0, 32'h4100177e, 32'h0, 32'h0, 32'h0, 32'h428c6dda, 32'h41ed5e6f};
test_input[10360:10367] = '{32'hc1fe711b, 32'hc2c58088, 32'h42854114, 32'hc1a35199, 32'h42b0ccf1, 32'h426c3813, 32'hc111faea, 32'h425598e3};
test_output[10360:10367] = '{32'h0, 32'h0, 32'h42854114, 32'h0, 32'h42b0ccf1, 32'h426c3813, 32'h0, 32'h425598e3};
test_input[10368:10375] = '{32'h42601ca4, 32'hc1a2deef, 32'h426aad48, 32'h4261d73b, 32'h424d8621, 32'hc225a110, 32'h410d00b4, 32'hc22c2e5e};
test_output[10368:10375] = '{32'h42601ca4, 32'h0, 32'h426aad48, 32'h4261d73b, 32'h424d8621, 32'h0, 32'h410d00b4, 32'h0};
test_input[10376:10383] = '{32'hc1e6119d, 32'h41cdf39e, 32'hc269d32a, 32'h4282404d, 32'h409c4b83, 32'hc1b9890d, 32'hc2c1b051, 32'hc2bce8f2};
test_output[10376:10383] = '{32'h0, 32'h41cdf39e, 32'h0, 32'h4282404d, 32'h409c4b83, 32'h0, 32'h0, 32'h0};
test_input[10384:10391] = '{32'hc1e8b99c, 32'h40a52498, 32'hc0b445a7, 32'hc27b13d2, 32'h42c07fab, 32'hc25b5921, 32'h4297077d, 32'h41b18e35};
test_output[10384:10391] = '{32'h0, 32'h40a52498, 32'h0, 32'h0, 32'h42c07fab, 32'h0, 32'h4297077d, 32'h41b18e35};
test_input[10392:10399] = '{32'hc255571f, 32'h421142ad, 32'hc2aa18dd, 32'hc239eea9, 32'h41a70856, 32'hc1dc244d, 32'h42b1a4f5, 32'hc2b15264};
test_output[10392:10399] = '{32'h0, 32'h421142ad, 32'h0, 32'h0, 32'h41a70856, 32'h0, 32'h42b1a4f5, 32'h0};
test_input[10400:10407] = '{32'hc2292860, 32'hc1afcf62, 32'hc146fa1f, 32'hc29cabfa, 32'hc200982b, 32'hc1bb1c96, 32'hc20994ce, 32'hc1d007fb};
test_output[10400:10407] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10408:10415] = '{32'h4121ba45, 32'hc0ca24a4, 32'hc208b097, 32'hc22be179, 32'h408ee7e7, 32'hc1f3517c, 32'hc1e3d954, 32'hc288a9ff};
test_output[10408:10415] = '{32'h4121ba45, 32'h0, 32'h0, 32'h0, 32'h408ee7e7, 32'h0, 32'h0, 32'h0};
test_input[10416:10423] = '{32'h41652b18, 32'h42561929, 32'h4266071f, 32'h42039bf0, 32'hc24ef97e, 32'h3eb87fd4, 32'h41f5b8df, 32'h42c37101};
test_output[10416:10423] = '{32'h41652b18, 32'h42561929, 32'h4266071f, 32'h42039bf0, 32'h0, 32'h3eb87fd4, 32'h41f5b8df, 32'h42c37101};
test_input[10424:10431] = '{32'h4022c920, 32'hc1fe5c95, 32'h428477f3, 32'hc127cded, 32'h42ba01b2, 32'hc208b9fb, 32'h4232055c, 32'hc267947d};
test_output[10424:10431] = '{32'h4022c920, 32'h0, 32'h428477f3, 32'h0, 32'h42ba01b2, 32'h0, 32'h4232055c, 32'h0};
test_input[10432:10439] = '{32'h42c2ba6a, 32'hc2bf52e0, 32'hc2aef545, 32'h4118c8ab, 32'h428d48c2, 32'hc19722a7, 32'h429f2e37, 32'h42c0c7af};
test_output[10432:10439] = '{32'h42c2ba6a, 32'h0, 32'h0, 32'h4118c8ab, 32'h428d48c2, 32'h0, 32'h429f2e37, 32'h42c0c7af};
test_input[10440:10447] = '{32'hc28ac532, 32'hc2254e14, 32'h4269a4dc, 32'h42c238ff, 32'hc288ead3, 32'h423397a5, 32'hc2212e8b, 32'h4215bcb7};
test_output[10440:10447] = '{32'h0, 32'h0, 32'h4269a4dc, 32'h42c238ff, 32'h0, 32'h423397a5, 32'h0, 32'h4215bcb7};
test_input[10448:10455] = '{32'hc2c18979, 32'h414c46d0, 32'h411e1ce0, 32'h42afe0de, 32'h40c396a3, 32'h41ff5120, 32'h420c0d1e, 32'h42aeb7d2};
test_output[10448:10455] = '{32'h0, 32'h414c46d0, 32'h411e1ce0, 32'h42afe0de, 32'h40c396a3, 32'h41ff5120, 32'h420c0d1e, 32'h42aeb7d2};
test_input[10456:10463] = '{32'h4277abfe, 32'hc2bcb998, 32'h3fe65745, 32'hc2047a32, 32'hc14fb428, 32'hc23460ca, 32'h4104eb8e, 32'hc2c7d461};
test_output[10456:10463] = '{32'h4277abfe, 32'h0, 32'h3fe65745, 32'h0, 32'h0, 32'h0, 32'h4104eb8e, 32'h0};
test_input[10464:10471] = '{32'hc299b51f, 32'hc252ecb1, 32'hc2af0fc3, 32'hc274fe54, 32'h420c5981, 32'hc1448532, 32'h42974cc2, 32'hc1ac74a0};
test_output[10464:10471] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h420c5981, 32'h0, 32'h42974cc2, 32'h0};
test_input[10472:10479] = '{32'h428e404a, 32'hc29bbe8c, 32'hc2737cc9, 32'h4222bc7d, 32'h423a474f, 32'h4178ee7f, 32'hc24b05f2, 32'hc223c54d};
test_output[10472:10479] = '{32'h428e404a, 32'h0, 32'h0, 32'h4222bc7d, 32'h423a474f, 32'h4178ee7f, 32'h0, 32'h0};
test_input[10480:10487] = '{32'hc2882f4d, 32'hc1e37bfb, 32'h405924ff, 32'hc1693509, 32'hc1d226f8, 32'hc2335d10, 32'h42a128a8, 32'hc2b48033};
test_output[10480:10487] = '{32'h0, 32'h0, 32'h405924ff, 32'h0, 32'h0, 32'h0, 32'h42a128a8, 32'h0};
test_input[10488:10495] = '{32'h42917194, 32'h42809186, 32'h42bd47ec, 32'hc0d9a616, 32'hc194d596, 32'h421f58b3, 32'h41acfa85, 32'hc06e93d9};
test_output[10488:10495] = '{32'h42917194, 32'h42809186, 32'h42bd47ec, 32'h0, 32'h0, 32'h421f58b3, 32'h41acfa85, 32'h0};
test_input[10496:10503] = '{32'hc26cc205, 32'hc233bd54, 32'h429e4146, 32'hc2bb878a, 32'hc145cb3e, 32'hc2c00907, 32'hc1dba7e1, 32'hc2bf2988};
test_output[10496:10503] = '{32'h0, 32'h0, 32'h429e4146, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10504:10511] = '{32'hc29853ee, 32'h3d8f1296, 32'h41dd2ab2, 32'h42016660, 32'h42ad7193, 32'h400c3a9c, 32'h42386fd6, 32'h4296aa8f};
test_output[10504:10511] = '{32'h0, 32'h3d8f1296, 32'h41dd2ab2, 32'h42016660, 32'h42ad7193, 32'h400c3a9c, 32'h42386fd6, 32'h4296aa8f};
test_input[10512:10519] = '{32'h4063266a, 32'h423837b9, 32'hc25accb4, 32'h420537f1, 32'hc23ff195, 32'h4149a040, 32'h428ecf68, 32'hbfaae4b7};
test_output[10512:10519] = '{32'h4063266a, 32'h423837b9, 32'h0, 32'h420537f1, 32'h0, 32'h4149a040, 32'h428ecf68, 32'h0};
test_input[10520:10527] = '{32'h424c1627, 32'hbd58f03d, 32'hc25731df, 32'h421f3261, 32'h41cee725, 32'hc2701bb4, 32'h413d5df5, 32'hc2156994};
test_output[10520:10527] = '{32'h424c1627, 32'h0, 32'h0, 32'h421f3261, 32'h41cee725, 32'h0, 32'h413d5df5, 32'h0};
test_input[10528:10535] = '{32'hc2888062, 32'h42abc8c1, 32'hc24ac3d3, 32'h429f64ff, 32'hc2206b3f, 32'hc109c3ee, 32'hc23581b8, 32'h4247fb7b};
test_output[10528:10535] = '{32'h0, 32'h42abc8c1, 32'h0, 32'h429f64ff, 32'h0, 32'h0, 32'h0, 32'h4247fb7b};
test_input[10536:10543] = '{32'hc201d667, 32'h3fc9befc, 32'hc0b1c955, 32'hc2acef36, 32'h4217a284, 32'hc1ec5b4b, 32'hc2aabc7f, 32'hc02825c1};
test_output[10536:10543] = '{32'h0, 32'h3fc9befc, 32'h0, 32'h0, 32'h4217a284, 32'h0, 32'h0, 32'h0};
test_input[10544:10551] = '{32'h4165d876, 32'h41ac43d3, 32'hc211b52a, 32'h42c4bd5f, 32'h419a481c, 32'hc296cc75, 32'hc26303c3, 32'hc1e76890};
test_output[10544:10551] = '{32'h4165d876, 32'h41ac43d3, 32'h0, 32'h42c4bd5f, 32'h419a481c, 32'h0, 32'h0, 32'h0};
test_input[10552:10559] = '{32'h426c62e7, 32'hc29f8b58, 32'hc29f1c13, 32'hc2311aa0, 32'hc22e480f, 32'hc24698aa, 32'hc23bc5f9, 32'h42bfed17};
test_output[10552:10559] = '{32'h426c62e7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bfed17};
test_input[10560:10567] = '{32'hc2261642, 32'h42344fab, 32'hc21cfbdf, 32'h40d87b54, 32'hc042e790, 32'h42b9e942, 32'h41a83616, 32'hc28a44d5};
test_output[10560:10567] = '{32'h0, 32'h42344fab, 32'h0, 32'h40d87b54, 32'h0, 32'h42b9e942, 32'h41a83616, 32'h0};
test_input[10568:10575] = '{32'h42ad2ace, 32'h42c7b779, 32'h42609af6, 32'h429ae66a, 32'hc2c2da28, 32'hc2c48ef2, 32'hc251c15c, 32'h4203efeb};
test_output[10568:10575] = '{32'h42ad2ace, 32'h42c7b779, 32'h42609af6, 32'h429ae66a, 32'h0, 32'h0, 32'h0, 32'h4203efeb};
test_input[10576:10583] = '{32'hc26803bf, 32'h42b27fed, 32'h426c92a7, 32'hc2bc8c26, 32'hc24f44ff, 32'hc18fee55, 32'hc2c00e8b, 32'hc1793ef7};
test_output[10576:10583] = '{32'h0, 32'h42b27fed, 32'h426c92a7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10584:10591] = '{32'h4254cafd, 32'h420394ed, 32'h42c15089, 32'hc24bf254, 32'hc21b9d7f, 32'h42319340, 32'hc248fb45, 32'hc1043094};
test_output[10584:10591] = '{32'h4254cafd, 32'h420394ed, 32'h42c15089, 32'h0, 32'h0, 32'h42319340, 32'h0, 32'h0};
test_input[10592:10599] = '{32'h42048102, 32'h422a9218, 32'h41142b6c, 32'hc2bfc0ce, 32'hc19b8db3, 32'h42650239, 32'h429861ab, 32'h42c731d5};
test_output[10592:10599] = '{32'h42048102, 32'h422a9218, 32'h41142b6c, 32'h0, 32'h0, 32'h42650239, 32'h429861ab, 32'h42c731d5};
test_input[10600:10607] = '{32'h401f0108, 32'hc027926b, 32'h41fab996, 32'h4243ebf0, 32'hc19a680b, 32'h41e32c8e, 32'hc0c0b3bb, 32'hc2088c93};
test_output[10600:10607] = '{32'h401f0108, 32'h0, 32'h41fab996, 32'h4243ebf0, 32'h0, 32'h41e32c8e, 32'h0, 32'h0};
test_input[10608:10615] = '{32'hc21f674b, 32'h411a65aa, 32'hc28e5155, 32'h415a1f39, 32'hc027a701, 32'h42202563, 32'hc264e30f, 32'h425fcce4};
test_output[10608:10615] = '{32'h0, 32'h411a65aa, 32'h0, 32'h415a1f39, 32'h0, 32'h42202563, 32'h0, 32'h425fcce4};
test_input[10616:10623] = '{32'h4299ec42, 32'hc2af5678, 32'hc13536f6, 32'hc2c635c6, 32'hc2a3739f, 32'hc1f827d4, 32'hc1795b03, 32'hc1dbdc75};
test_output[10616:10623] = '{32'h4299ec42, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10624:10631] = '{32'hc2b06341, 32'hc289635c, 32'hc295e761, 32'h42ac0e13, 32'hc1f1409d, 32'hc284dde1, 32'hc29f766a, 32'h4063121c};
test_output[10624:10631] = '{32'h0, 32'h0, 32'h0, 32'h42ac0e13, 32'h0, 32'h0, 32'h0, 32'h4063121c};
test_input[10632:10639] = '{32'hc1c2aa9c, 32'h4244bd28, 32'hc1bacb88, 32'hbffddaed, 32'h429d434d, 32'hc2168c48, 32'hc0459912, 32'hc094d962};
test_output[10632:10639] = '{32'h0, 32'h4244bd28, 32'h0, 32'h0, 32'h429d434d, 32'h0, 32'h0, 32'h0};
test_input[10640:10647] = '{32'h42b9047e, 32'hc1192658, 32'hc29c7190, 32'hc23fd1b2, 32'h428a1e10, 32'h40fa5de9, 32'h41eebcab, 32'hc28d9ed2};
test_output[10640:10647] = '{32'h42b9047e, 32'h0, 32'h0, 32'h0, 32'h428a1e10, 32'h40fa5de9, 32'h41eebcab, 32'h0};
test_input[10648:10655] = '{32'hc28ba1d3, 32'h425b3bec, 32'hc1b11ab8, 32'h424ff84a, 32'hc1c70fd8, 32'hc258a2de, 32'h42c46615, 32'hc17c5d0d};
test_output[10648:10655] = '{32'h0, 32'h425b3bec, 32'h0, 32'h424ff84a, 32'h0, 32'h0, 32'h42c46615, 32'h0};
test_input[10656:10663] = '{32'h41ec9de8, 32'hc2b4f8d7, 32'h42664c9f, 32'h41b13309, 32'hc091ad76, 32'hc1b11fd7, 32'h42aca5d3, 32'hc2984479};
test_output[10656:10663] = '{32'h41ec9de8, 32'h0, 32'h42664c9f, 32'h41b13309, 32'h0, 32'h0, 32'h42aca5d3, 32'h0};
test_input[10664:10671] = '{32'hc29b6fb8, 32'h42b504f4, 32'h415c05a0, 32'hc2aa5a33, 32'h422d2ac8, 32'h42b5ad35, 32'hc24d2bc8, 32'h4299f8d3};
test_output[10664:10671] = '{32'h0, 32'h42b504f4, 32'h415c05a0, 32'h0, 32'h422d2ac8, 32'h42b5ad35, 32'h0, 32'h4299f8d3};
test_input[10672:10679] = '{32'hc24e2106, 32'h413f4dee, 32'hc26b2f8e, 32'h423affc2, 32'hc290f0b8, 32'h420adbff, 32'h42a5784a, 32'h4213a55e};
test_output[10672:10679] = '{32'h0, 32'h413f4dee, 32'h0, 32'h423affc2, 32'h0, 32'h420adbff, 32'h42a5784a, 32'h4213a55e};
test_input[10680:10687] = '{32'h42815fce, 32'hc2b24a53, 32'h42b6733c, 32'h42c5a411, 32'h42c7135d, 32'hc1f6a478, 32'h407037fa, 32'h4290a5ff};
test_output[10680:10687] = '{32'h42815fce, 32'h0, 32'h42b6733c, 32'h42c5a411, 32'h42c7135d, 32'h0, 32'h407037fa, 32'h4290a5ff};
test_input[10688:10695] = '{32'h4110174d, 32'h3f909a44, 32'hc29be9a2, 32'h4255bc31, 32'h403e93a5, 32'hc1126b6c, 32'h42079d03, 32'hc1b8992b};
test_output[10688:10695] = '{32'h4110174d, 32'h3f909a44, 32'h0, 32'h4255bc31, 32'h403e93a5, 32'h0, 32'h42079d03, 32'h0};
test_input[10696:10703] = '{32'hc2260397, 32'hc2913a63, 32'h42b2139a, 32'h4279f1e1, 32'h421d6174, 32'hc2a9c98c, 32'h4253afa3, 32'h413c283e};
test_output[10696:10703] = '{32'h0, 32'h0, 32'h42b2139a, 32'h4279f1e1, 32'h421d6174, 32'h0, 32'h4253afa3, 32'h413c283e};
test_input[10704:10711] = '{32'h42892055, 32'hc21331f4, 32'h425fc7a7, 32'h413bb5d9, 32'h42b58433, 32'hc29391e1, 32'hc2512ffe, 32'h42b3f398};
test_output[10704:10711] = '{32'h42892055, 32'h0, 32'h425fc7a7, 32'h413bb5d9, 32'h42b58433, 32'h0, 32'h0, 32'h42b3f398};
test_input[10712:10719] = '{32'h4292e6e0, 32'h41cedfa3, 32'h420fb54b, 32'h428d3797, 32'hc21b5048, 32'hc19a97fc, 32'h41a62b64, 32'h424b0388};
test_output[10712:10719] = '{32'h4292e6e0, 32'h41cedfa3, 32'h420fb54b, 32'h428d3797, 32'h0, 32'h0, 32'h41a62b64, 32'h424b0388};
test_input[10720:10727] = '{32'h42079baa, 32'h41afdebe, 32'hc2282759, 32'h40aff643, 32'hc02ae219, 32'hc10701e7, 32'h4197de7a, 32'h42a5418d};
test_output[10720:10727] = '{32'h42079baa, 32'h41afdebe, 32'h0, 32'h40aff643, 32'h0, 32'h0, 32'h4197de7a, 32'h42a5418d};
test_input[10728:10735] = '{32'hc21583e2, 32'hc29849c7, 32'hc25d2cbc, 32'h4295a230, 32'h429e9ad5, 32'h41ddfc22, 32'h420b7407, 32'hc2142014};
test_output[10728:10735] = '{32'h0, 32'h0, 32'h0, 32'h4295a230, 32'h429e9ad5, 32'h41ddfc22, 32'h420b7407, 32'h0};
test_input[10736:10743] = '{32'h42c08d58, 32'hc2b5d84d, 32'hc287d8ba, 32'hc1fbcc50, 32'h4021ecfa, 32'h4115f677, 32'h42749890, 32'h41b9d74a};
test_output[10736:10743] = '{32'h42c08d58, 32'h0, 32'h0, 32'h0, 32'h4021ecfa, 32'h4115f677, 32'h42749890, 32'h41b9d74a};
test_input[10744:10751] = '{32'hc29fbf40, 32'hc27a6ac8, 32'hc2814d9e, 32'hc1fc073d, 32'hc195b04a, 32'hc25d3d9c, 32'h4245bfc0, 32'h424af58f};
test_output[10744:10751] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4245bfc0, 32'h424af58f};
test_input[10752:10759] = '{32'h41d203af, 32'h42a52aa2, 32'hc0ac2356, 32'h413a3fa8, 32'hc2c7195e, 32'hc281b0ba, 32'h42696357, 32'hc26c0d3a};
test_output[10752:10759] = '{32'h41d203af, 32'h42a52aa2, 32'h0, 32'h413a3fa8, 32'h0, 32'h0, 32'h42696357, 32'h0};
test_input[10760:10767] = '{32'hc2107bd2, 32'hc15172d8, 32'hc25aa6f5, 32'hc23ee6ee, 32'h41ac8fcd, 32'h4000f161, 32'h4225a0f1, 32'h42a3fdaf};
test_output[10760:10767] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41ac8fcd, 32'h4000f161, 32'h4225a0f1, 32'h42a3fdaf};
test_input[10768:10775] = '{32'hc2bd4872, 32'h40d479f4, 32'h42238fb8, 32'h41fef2f2, 32'h4224c31f, 32'h42b11c2a, 32'h421437f9, 32'hc2057b05};
test_output[10768:10775] = '{32'h0, 32'h40d479f4, 32'h42238fb8, 32'h41fef2f2, 32'h4224c31f, 32'h42b11c2a, 32'h421437f9, 32'h0};
test_input[10776:10783] = '{32'h42869828, 32'hc2333747, 32'h42984a2c, 32'hc15e7d08, 32'hc262bb15, 32'hc2ba4dfa, 32'hc188c052, 32'hc2bd41b4};
test_output[10776:10783] = '{32'h42869828, 32'h0, 32'h42984a2c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10784:10791] = '{32'hc2236483, 32'h42a98a7b, 32'h4126e846, 32'hc27bc593, 32'h4284991a, 32'hc29e8ea6, 32'h415236c2, 32'hc178893a};
test_output[10784:10791] = '{32'h0, 32'h42a98a7b, 32'h4126e846, 32'h0, 32'h4284991a, 32'h0, 32'h415236c2, 32'h0};
test_input[10792:10799] = '{32'hc28d83aa, 32'hc29757b5, 32'h429daaa4, 32'h426a67ac, 32'h42ae14b7, 32'h42c45e82, 32'h41ace29c, 32'hc29cbecb};
test_output[10792:10799] = '{32'h0, 32'h0, 32'h429daaa4, 32'h426a67ac, 32'h42ae14b7, 32'h42c45e82, 32'h41ace29c, 32'h0};
test_input[10800:10807] = '{32'hc28c694a, 32'hc229187f, 32'h41b43394, 32'h4211c0aa, 32'hc1afbb59, 32'hc14fe54e, 32'h423fa4a9, 32'h41a2ebbb};
test_output[10800:10807] = '{32'h0, 32'h0, 32'h41b43394, 32'h4211c0aa, 32'h0, 32'h0, 32'h423fa4a9, 32'h41a2ebbb};
test_input[10808:10815] = '{32'hc12a337c, 32'h4232259a, 32'hc1c5e419, 32'h42bf77fd, 32'hc1fdd326, 32'h42aafb41, 32'h429d07d9, 32'h41ae0c03};
test_output[10808:10815] = '{32'h0, 32'h4232259a, 32'h0, 32'h42bf77fd, 32'h0, 32'h42aafb41, 32'h429d07d9, 32'h41ae0c03};
test_input[10816:10823] = '{32'h412302f5, 32'hbf34b204, 32'h416f4a4c, 32'h429de00d, 32'h419cab0b, 32'h412a1e5a, 32'hc2a61fc9, 32'h41d0c345};
test_output[10816:10823] = '{32'h412302f5, 32'h0, 32'h416f4a4c, 32'h429de00d, 32'h419cab0b, 32'h412a1e5a, 32'h0, 32'h41d0c345};
test_input[10824:10831] = '{32'hc2ad30e7, 32'hc28e62b0, 32'h42b1e7df, 32'hc1af9a10, 32'h40c8b0e6, 32'h420cc1eb, 32'hc24d2f4e, 32'hc24bb31f};
test_output[10824:10831] = '{32'h0, 32'h0, 32'h42b1e7df, 32'h0, 32'h40c8b0e6, 32'h420cc1eb, 32'h0, 32'h0};
test_input[10832:10839] = '{32'hc2a5b1c7, 32'hc21df78f, 32'hc2868b61, 32'h41da7d44, 32'hc2132748, 32'hc2413fe1, 32'hc24e76b8, 32'hc2a4ab94};
test_output[10832:10839] = '{32'h0, 32'h0, 32'h0, 32'h41da7d44, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10840:10847] = '{32'h4151ef5d, 32'hc2070203, 32'hc0ad8e9f, 32'h4299bfe2, 32'hc2c465ed, 32'h4246da20, 32'h42916d7a, 32'h425cabcc};
test_output[10840:10847] = '{32'h4151ef5d, 32'h0, 32'h0, 32'h4299bfe2, 32'h0, 32'h4246da20, 32'h42916d7a, 32'h425cabcc};
test_input[10848:10855] = '{32'hc2c1628b, 32'hc24ac952, 32'h42c139bf, 32'h41c65786, 32'h4268f6c3, 32'hc2aecc06, 32'h42561461, 32'hc205cd1f};
test_output[10848:10855] = '{32'h0, 32'h0, 32'h42c139bf, 32'h41c65786, 32'h4268f6c3, 32'h0, 32'h42561461, 32'h0};
test_input[10856:10863] = '{32'h418bcb11, 32'hc2b471dd, 32'h41149528, 32'h42b945e8, 32'hc296f3b7, 32'h4294d7aa, 32'h41e62c6b, 32'h4206610b};
test_output[10856:10863] = '{32'h418bcb11, 32'h0, 32'h41149528, 32'h42b945e8, 32'h0, 32'h4294d7aa, 32'h41e62c6b, 32'h4206610b};
test_input[10864:10871] = '{32'hc2b75622, 32'hc262df76, 32'hc2b3c31d, 32'h40aa4f8f, 32'hc2922f92, 32'h40fc8c6b, 32'h429ab9e0, 32'hc1f2d735};
test_output[10864:10871] = '{32'h0, 32'h0, 32'h0, 32'h40aa4f8f, 32'h0, 32'h40fc8c6b, 32'h429ab9e0, 32'h0};
test_input[10872:10879] = '{32'hc20d648d, 32'h405a196d, 32'h427a7b43, 32'h4222fad0, 32'hc2adbfb8, 32'h428d2bc3, 32'h418e7ca7, 32'h42b4a34d};
test_output[10872:10879] = '{32'h0, 32'h405a196d, 32'h427a7b43, 32'h4222fad0, 32'h0, 32'h428d2bc3, 32'h418e7ca7, 32'h42b4a34d};
test_input[10880:10887] = '{32'h3f25ab89, 32'hc29ca88a, 32'h4286a57e, 32'hc2788a2d, 32'hc0db5e45, 32'h4243926e, 32'h4195afdf, 32'h426e75cf};
test_output[10880:10887] = '{32'h3f25ab89, 32'h0, 32'h4286a57e, 32'h0, 32'h0, 32'h4243926e, 32'h4195afdf, 32'h426e75cf};
test_input[10888:10895] = '{32'h42a605cc, 32'hc1eaba78, 32'h42070433, 32'h42089782, 32'hc22b2e28, 32'h42ab0274, 32'hc23cb206, 32'h42209b52};
test_output[10888:10895] = '{32'h42a605cc, 32'h0, 32'h42070433, 32'h42089782, 32'h0, 32'h42ab0274, 32'h0, 32'h42209b52};
test_input[10896:10903] = '{32'hc22eab62, 32'hc2aa8ee5, 32'h41ad6ec3, 32'hc1bd7b8a, 32'h42ab2486, 32'h42a87456, 32'hc1954c5a, 32'hc23a8a2a};
test_output[10896:10903] = '{32'h0, 32'h0, 32'h41ad6ec3, 32'h0, 32'h42ab2486, 32'h42a87456, 32'h0, 32'h0};
test_input[10904:10911] = '{32'h423423b7, 32'hc24a49b4, 32'h42038635, 32'hc2af8e34, 32'hc26f487a, 32'h42a72c9e, 32'h42983d5f, 32'h41da8065};
test_output[10904:10911] = '{32'h423423b7, 32'h0, 32'h42038635, 32'h0, 32'h0, 32'h42a72c9e, 32'h42983d5f, 32'h41da8065};
test_input[10912:10919] = '{32'hc2a7f250, 32'h414b43d1, 32'hc1d848bd, 32'hc05c09ef, 32'hc2586380, 32'hc20e3f94, 32'hc2657bcc, 32'h40a10ad9};
test_output[10912:10919] = '{32'h0, 32'h414b43d1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40a10ad9};
test_input[10920:10927] = '{32'h3f773b4d, 32'h42b405e4, 32'hc206114d, 32'h4222170a, 32'hc2b25ab8, 32'h4298b4b5, 32'h42b99e38, 32'h42a4f44c};
test_output[10920:10927] = '{32'h3f773b4d, 32'h42b405e4, 32'h0, 32'h4222170a, 32'h0, 32'h4298b4b5, 32'h42b99e38, 32'h42a4f44c};
test_input[10928:10935] = '{32'hc2039ea8, 32'hc0cd28cd, 32'hc242fc91, 32'hc20d3028, 32'h3fcad3e8, 32'h401c69ea, 32'hc22fcec8, 32'hc2a92875};
test_output[10928:10935] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h3fcad3e8, 32'h401c69ea, 32'h0, 32'h0};
test_input[10936:10943] = '{32'hc2b05f8b, 32'hc1965aeb, 32'h4291113c, 32'h429b9d78, 32'hc1c886a7, 32'hc28b9165, 32'hc2096e39, 32'hc250418a};
test_output[10936:10943] = '{32'h0, 32'h0, 32'h4291113c, 32'h429b9d78, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10944:10951] = '{32'hc22fc208, 32'hc22c6035, 32'hc16dc776, 32'hc2124da7, 32'h423cd430, 32'hc115ca01, 32'hc257aeb2, 32'h4125d5e8};
test_output[10944:10951] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h423cd430, 32'h0, 32'h0, 32'h4125d5e8};
test_input[10952:10959] = '{32'hc26b5fa1, 32'h4079aa82, 32'hc284abce, 32'hc0d12a53, 32'hc2aede7f, 32'hc2c01d01, 32'hc26c0f11, 32'hc194fab4};
test_output[10952:10959] = '{32'h0, 32'h4079aa82, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[10960:10967] = '{32'h418c7051, 32'hc2c7b3e9, 32'hc2001296, 32'h425ac90e, 32'h4189b60f, 32'h423e4252, 32'h416a670e, 32'hc1cba357};
test_output[10960:10967] = '{32'h418c7051, 32'h0, 32'h0, 32'h425ac90e, 32'h4189b60f, 32'h423e4252, 32'h416a670e, 32'h0};
test_input[10968:10975] = '{32'hc2a36fd0, 32'h41d737a9, 32'h428b1430, 32'hc28437e7, 32'hc2a97c4e, 32'hc234a000, 32'hc298ddf0, 32'h42c7659b};
test_output[10968:10975] = '{32'h0, 32'h41d737a9, 32'h428b1430, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c7659b};
test_input[10976:10983] = '{32'h42ab31a3, 32'h4277b404, 32'h421392d2, 32'h42b5d113, 32'h42965a9a, 32'hc2194cea, 32'hc200de45, 32'hc2c578b7};
test_output[10976:10983] = '{32'h42ab31a3, 32'h4277b404, 32'h421392d2, 32'h42b5d113, 32'h42965a9a, 32'h0, 32'h0, 32'h0};
test_input[10984:10991] = '{32'hc2477bb2, 32'h4103c58a, 32'hc2b5ec03, 32'h3f867b89, 32'hc292a017, 32'hc1ecd1d0, 32'hc23c3564, 32'h42b32ef9};
test_output[10984:10991] = '{32'h0, 32'h4103c58a, 32'h0, 32'h3f867b89, 32'h0, 32'h0, 32'h0, 32'h42b32ef9};
test_input[10992:10999] = '{32'hc2bd98cc, 32'h42b54766, 32'hc24ae92c, 32'h42081849, 32'h4228675a, 32'hc291526f, 32'hc2aabcbf, 32'hc2a6b134};
test_output[10992:10999] = '{32'h0, 32'h42b54766, 32'h0, 32'h42081849, 32'h4228675a, 32'h0, 32'h0, 32'h0};
test_input[11000:11007] = '{32'h41dfd0f8, 32'hc0afaab2, 32'h419cdc26, 32'hc2459cdf, 32'hc1391f19, 32'hc1907ffe, 32'hc0ed7ff7, 32'hc2789877};
test_output[11000:11007] = '{32'h41dfd0f8, 32'h0, 32'h419cdc26, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11008:11015] = '{32'h403ac241, 32'h4216444c, 32'h41d5c4e5, 32'hc1bb1a67, 32'hc263b805, 32'h422e9813, 32'hc2991413, 32'h42b03d38};
test_output[11008:11015] = '{32'h403ac241, 32'h4216444c, 32'h41d5c4e5, 32'h0, 32'h0, 32'h422e9813, 32'h0, 32'h42b03d38};
test_input[11016:11023] = '{32'h4248cd63, 32'h4241d584, 32'h424d4564, 32'hc1db9fa6, 32'h42011016, 32'hc23bea52, 32'h41a11aed, 32'hc26c1d98};
test_output[11016:11023] = '{32'h4248cd63, 32'h4241d584, 32'h424d4564, 32'h0, 32'h42011016, 32'h0, 32'h41a11aed, 32'h0};
test_input[11024:11031] = '{32'hc2bf618d, 32'hc1cff7b4, 32'h40459ca4, 32'hc25034d9, 32'h422c6c3e, 32'hc2910fa4, 32'h419d32a7, 32'hc27f3eca};
test_output[11024:11031] = '{32'h0, 32'h0, 32'h40459ca4, 32'h0, 32'h422c6c3e, 32'h0, 32'h419d32a7, 32'h0};
test_input[11032:11039] = '{32'h4219140a, 32'hc29833a3, 32'h4167b3c8, 32'h42432b22, 32'h42aed66c, 32'h40ba0505, 32'h42af64f7, 32'hc216653c};
test_output[11032:11039] = '{32'h4219140a, 32'h0, 32'h4167b3c8, 32'h42432b22, 32'h42aed66c, 32'h40ba0505, 32'h42af64f7, 32'h0};
test_input[11040:11047] = '{32'h4179df71, 32'h3fd1c70d, 32'h429ae12c, 32'h42808728, 32'h41144834, 32'h42c4f071, 32'h428b4afd, 32'hc2a06c48};
test_output[11040:11047] = '{32'h4179df71, 32'h3fd1c70d, 32'h429ae12c, 32'h42808728, 32'h41144834, 32'h42c4f071, 32'h428b4afd, 32'h0};
test_input[11048:11055] = '{32'hc28df659, 32'hc1a8b16b, 32'hc2bfa4ef, 32'h4065459a, 32'h429e4d34, 32'hc2bcfcf4, 32'hc1cc9f23, 32'h4280cd0d};
test_output[11048:11055] = '{32'h0, 32'h0, 32'h0, 32'h4065459a, 32'h429e4d34, 32'h0, 32'h0, 32'h4280cd0d};
test_input[11056:11063] = '{32'h41858b10, 32'h4129be43, 32'hc247ed69, 32'hc2b317e4, 32'hc1bde723, 32'h422eb858, 32'hc29052ee, 32'h421975af};
test_output[11056:11063] = '{32'h41858b10, 32'h4129be43, 32'h0, 32'h0, 32'h0, 32'h422eb858, 32'h0, 32'h421975af};
test_input[11064:11071] = '{32'hc1110ec9, 32'hc14fce4b, 32'hc10e13f0, 32'hc2899483, 32'hc24f3cb9, 32'h41ef8891, 32'h42b7830f, 32'h42bd8e0b};
test_output[11064:11071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ef8891, 32'h42b7830f, 32'h42bd8e0b};
test_input[11072:11079] = '{32'h428beed0, 32'h424c70f8, 32'hc2bfebc4, 32'h41f1ed97, 32'h423ffab8, 32'h42398594, 32'h421bbbc0, 32'h41f5064d};
test_output[11072:11079] = '{32'h428beed0, 32'h424c70f8, 32'h0, 32'h41f1ed97, 32'h423ffab8, 32'h42398594, 32'h421bbbc0, 32'h41f5064d};
test_input[11080:11087] = '{32'h429117a1, 32'h415ccdf5, 32'hc28661db, 32'hc2a1677c, 32'h423ff4fe, 32'h413c2154, 32'h41ff87da, 32'h427117cf};
test_output[11080:11087] = '{32'h429117a1, 32'h415ccdf5, 32'h0, 32'h0, 32'h423ff4fe, 32'h413c2154, 32'h41ff87da, 32'h427117cf};
test_input[11088:11095] = '{32'hc089d19b, 32'h4263e8c5, 32'h411448aa, 32'h3fcb5d96, 32'hc2c0d97d, 32'h4200868d, 32'h41e0c15d, 32'h400db841};
test_output[11088:11095] = '{32'h0, 32'h4263e8c5, 32'h411448aa, 32'h3fcb5d96, 32'h0, 32'h4200868d, 32'h41e0c15d, 32'h400db841};
test_input[11096:11103] = '{32'hc2595d03, 32'h42afbe2c, 32'h411ed4b5, 32'hc21d9ecf, 32'hc2bbeb4e, 32'hc2925146, 32'h4011e335, 32'h42a47b31};
test_output[11096:11103] = '{32'h0, 32'h42afbe2c, 32'h411ed4b5, 32'h0, 32'h0, 32'h0, 32'h4011e335, 32'h42a47b31};
test_input[11104:11111] = '{32'h420d67d4, 32'hc1e2ed0a, 32'hc2166833, 32'h428be1ef, 32'hc2119818, 32'hc2beb809, 32'h423be76b, 32'h42a047d1};
test_output[11104:11111] = '{32'h420d67d4, 32'h0, 32'h0, 32'h428be1ef, 32'h0, 32'h0, 32'h423be76b, 32'h42a047d1};
test_input[11112:11119] = '{32'h3fca1fc4, 32'hc184ded7, 32'h42ba61e7, 32'hc185c253, 32'hc14fbd5b, 32'hc2a847b8, 32'h42a16fd5, 32'hc20ca518};
test_output[11112:11119] = '{32'h3fca1fc4, 32'h0, 32'h42ba61e7, 32'h0, 32'h0, 32'h0, 32'h42a16fd5, 32'h0};
test_input[11120:11127] = '{32'h42c0eba6, 32'h42be9185, 32'h42408d87, 32'h427eec97, 32'h404c6c5c, 32'h4266bc7c, 32'hc25c5c95, 32'h419ead7a};
test_output[11120:11127] = '{32'h42c0eba6, 32'h42be9185, 32'h42408d87, 32'h427eec97, 32'h404c6c5c, 32'h4266bc7c, 32'h0, 32'h419ead7a};
test_input[11128:11135] = '{32'h41dbf6db, 32'h42b2e6c9, 32'hc2848eca, 32'h42543f52, 32'h40d4f9bc, 32'hc253fd76, 32'h40808645, 32'h421cb3fa};
test_output[11128:11135] = '{32'h41dbf6db, 32'h42b2e6c9, 32'h0, 32'h42543f52, 32'h40d4f9bc, 32'h0, 32'h40808645, 32'h421cb3fa};
test_input[11136:11143] = '{32'hc2b4da29, 32'h4211c4a0, 32'hbfedd52b, 32'h4235e4ad, 32'h402966a3, 32'h428e023d, 32'h4273c949, 32'h424bc1b0};
test_output[11136:11143] = '{32'h0, 32'h4211c4a0, 32'h0, 32'h4235e4ad, 32'h402966a3, 32'h428e023d, 32'h4273c949, 32'h424bc1b0};
test_input[11144:11151] = '{32'h422d8839, 32'hc263576e, 32'h4108db80, 32'h41c9953d, 32'h4159e1da, 32'hc039cda9, 32'h42bb3660, 32'h42bd7d3a};
test_output[11144:11151] = '{32'h422d8839, 32'h0, 32'h4108db80, 32'h41c9953d, 32'h4159e1da, 32'h0, 32'h42bb3660, 32'h42bd7d3a};
test_input[11152:11159] = '{32'h416c1fe1, 32'h421e7232, 32'hc20ddcc4, 32'h41760268, 32'hc00d0d57, 32'hc2b2dce8, 32'hc2b446e2, 32'h42ad9cb3};
test_output[11152:11159] = '{32'h416c1fe1, 32'h421e7232, 32'h0, 32'h41760268, 32'h0, 32'h0, 32'h0, 32'h42ad9cb3};
test_input[11160:11167] = '{32'hc2a85003, 32'hc14b676c, 32'hc210f57e, 32'h426ce23b, 32'hc29a484e, 32'hc20e7615, 32'h4294c648, 32'h4195f419};
test_output[11160:11167] = '{32'h0, 32'h0, 32'h0, 32'h426ce23b, 32'h0, 32'h0, 32'h4294c648, 32'h4195f419};
test_input[11168:11175] = '{32'h41d33bdb, 32'h42b99862, 32'hc1cfa248, 32'hc0961aa3, 32'h41e12f4a, 32'h42283d02, 32'h412e6d74, 32'hc115348a};
test_output[11168:11175] = '{32'h41d33bdb, 32'h42b99862, 32'h0, 32'h0, 32'h41e12f4a, 32'h42283d02, 32'h412e6d74, 32'h0};
test_input[11176:11183] = '{32'hc2075f1c, 32'hc25684d8, 32'h4290c1cb, 32'hc2544062, 32'h429bcc3f, 32'hc1f32e14, 32'h429ff287, 32'h42b5c62b};
test_output[11176:11183] = '{32'h0, 32'h0, 32'h4290c1cb, 32'h0, 32'h429bcc3f, 32'h0, 32'h429ff287, 32'h42b5c62b};
test_input[11184:11191] = '{32'h42c4f7f8, 32'h4019853d, 32'h421c9704, 32'h42b32a99, 32'h4048adbf, 32'hc2c4fc3d, 32'hc2b465dd, 32'h411308bd};
test_output[11184:11191] = '{32'h42c4f7f8, 32'h4019853d, 32'h421c9704, 32'h42b32a99, 32'h4048adbf, 32'h0, 32'h0, 32'h411308bd};
test_input[11192:11199] = '{32'h428cedef, 32'h41d4cde1, 32'hc10ab210, 32'hc19e5b04, 32'h4230e688, 32'hc2b74a51, 32'h428de741, 32'hc2b8f417};
test_output[11192:11199] = '{32'h428cedef, 32'h41d4cde1, 32'h0, 32'h0, 32'h4230e688, 32'h0, 32'h428de741, 32'h0};
test_input[11200:11207] = '{32'hc01f0c76, 32'hc194fd92, 32'hc26f0cbe, 32'hc2817d80, 32'h41adf7b5, 32'h4281208d, 32'hc1382bb2, 32'hc291845e};
test_output[11200:11207] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41adf7b5, 32'h4281208d, 32'h0, 32'h0};
test_input[11208:11215] = '{32'hc28f8e73, 32'hc2c09c01, 32'hc2aa391a, 32'h411dc53f, 32'hc2ab7819, 32'h42c5e48a, 32'hc1d800c6, 32'h42a7d70a};
test_output[11208:11215] = '{32'h0, 32'h0, 32'h0, 32'h411dc53f, 32'h0, 32'h42c5e48a, 32'h0, 32'h42a7d70a};
test_input[11216:11223] = '{32'hc2409eaf, 32'h428dfb9d, 32'hc217ff82, 32'h42931bb3, 32'h42b5ba40, 32'h411b2308, 32'h41cdaaf2, 32'hc1d2f408};
test_output[11216:11223] = '{32'h0, 32'h428dfb9d, 32'h0, 32'h42931bb3, 32'h42b5ba40, 32'h411b2308, 32'h41cdaaf2, 32'h0};
test_input[11224:11231] = '{32'h3fc8cf39, 32'hc26e8bd4, 32'hc29edcfa, 32'h427cf404, 32'hc196cccd, 32'hc187a3b0, 32'h428d6674, 32'h426823c4};
test_output[11224:11231] = '{32'h3fc8cf39, 32'h0, 32'h0, 32'h427cf404, 32'h0, 32'h0, 32'h428d6674, 32'h426823c4};
test_input[11232:11239] = '{32'hc20deb16, 32'hc1034792, 32'hc269beba, 32'h4295fb63, 32'h42adccb8, 32'h42abd7d2, 32'h421af762, 32'hc1749f0e};
test_output[11232:11239] = '{32'h0, 32'h0, 32'h0, 32'h4295fb63, 32'h42adccb8, 32'h42abd7d2, 32'h421af762, 32'h0};
test_input[11240:11247] = '{32'hc21bb29e, 32'h4282588e, 32'hc2b8a993, 32'h41ce56c3, 32'hc14c91f7, 32'hc2a0d9c1, 32'hc270df5c, 32'h427bc7ee};
test_output[11240:11247] = '{32'h0, 32'h4282588e, 32'h0, 32'h41ce56c3, 32'h0, 32'h0, 32'h0, 32'h427bc7ee};
test_input[11248:11255] = '{32'h42b13169, 32'h429cb37d, 32'h42773484, 32'hc2ac3c96, 32'h422f0681, 32'hc1fbe907, 32'h41237ffc, 32'hc2093c02};
test_output[11248:11255] = '{32'h42b13169, 32'h429cb37d, 32'h42773484, 32'h0, 32'h422f0681, 32'h0, 32'h41237ffc, 32'h0};
test_input[11256:11263] = '{32'h40ae82c0, 32'hc2305f4d, 32'hc24e19a1, 32'hc2983b20, 32'hc2279955, 32'h42a16efe, 32'h421710b7, 32'h428bff6a};
test_output[11256:11263] = '{32'h40ae82c0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a16efe, 32'h421710b7, 32'h428bff6a};
test_input[11264:11271] = '{32'h4241f22f, 32'hc25755c9, 32'h428adc5c, 32'h401a5446, 32'hc1be1b0b, 32'hc121de29, 32'h42a60f50, 32'hc25334ba};
test_output[11264:11271] = '{32'h4241f22f, 32'h0, 32'h428adc5c, 32'h401a5446, 32'h0, 32'h0, 32'h42a60f50, 32'h0};
test_input[11272:11279] = '{32'hc244ffb7, 32'h41919d99, 32'hc247f6c4, 32'hc21c1d11, 32'h4276f992, 32'h41f2494e, 32'h40d99272, 32'hc2927320};
test_output[11272:11279] = '{32'h0, 32'h41919d99, 32'h0, 32'h0, 32'h4276f992, 32'h41f2494e, 32'h40d99272, 32'h0};
test_input[11280:11287] = '{32'h42a53ac1, 32'h4294d5f5, 32'h421c6cb9, 32'hc27fe83f, 32'hc29f837c, 32'hc1eb8edb, 32'h428f6ac0, 32'h41513fa1};
test_output[11280:11287] = '{32'h42a53ac1, 32'h4294d5f5, 32'h421c6cb9, 32'h0, 32'h0, 32'h0, 32'h428f6ac0, 32'h41513fa1};
test_input[11288:11295] = '{32'h4259781f, 32'hc2bc0b1c, 32'h42abf7a3, 32'h429e3135, 32'hc281001b, 32'h410b268f, 32'h3fb24443, 32'hc23fc499};
test_output[11288:11295] = '{32'h4259781f, 32'h0, 32'h42abf7a3, 32'h429e3135, 32'h0, 32'h410b268f, 32'h3fb24443, 32'h0};
test_input[11296:11303] = '{32'h42c58317, 32'hc29708a7, 32'h413aa983, 32'hc24f18fb, 32'hc1821d8a, 32'hc285f60b, 32'h42a56a18, 32'h408265a4};
test_output[11296:11303] = '{32'h42c58317, 32'h0, 32'h413aa983, 32'h0, 32'h0, 32'h0, 32'h42a56a18, 32'h408265a4};
test_input[11304:11311] = '{32'h41158a39, 32'h429c75b4, 32'hc2aa39ac, 32'hc220727c, 32'hc252584f, 32'hc1cbf7fb, 32'hc2b51ff7, 32'hc2b66146};
test_output[11304:11311] = '{32'h41158a39, 32'h429c75b4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11312:11319] = '{32'hc20cc47e, 32'hc276a744, 32'hc2a392c1, 32'h418c1996, 32'hc15d0eb8, 32'h4278de5e, 32'hc2897c0e, 32'hc24560b7};
test_output[11312:11319] = '{32'h0, 32'h0, 32'h0, 32'h418c1996, 32'h0, 32'h4278de5e, 32'h0, 32'h0};
test_input[11320:11327] = '{32'hc2b34d14, 32'h4286718d, 32'hc1d6857d, 32'h424305f9, 32'h41ea1b00, 32'hc1fdd0fc, 32'hc2b6645e, 32'hc1ebe860};
test_output[11320:11327] = '{32'h0, 32'h4286718d, 32'h0, 32'h424305f9, 32'h41ea1b00, 32'h0, 32'h0, 32'h0};
test_input[11328:11335] = '{32'hc1a8275f, 32'h415fb162, 32'hc08bb529, 32'h40c879a1, 32'h42b6cb39, 32'hc19d2df5, 32'hc29791be, 32'h423b5305};
test_output[11328:11335] = '{32'h0, 32'h415fb162, 32'h0, 32'h40c879a1, 32'h42b6cb39, 32'h0, 32'h0, 32'h423b5305};
test_input[11336:11343] = '{32'h421dde5f, 32'h4296dbda, 32'h40ad9221, 32'hc21e5380, 32'h41863ce3, 32'h41bc42b0, 32'hc194cba1, 32'h4267eb36};
test_output[11336:11343] = '{32'h421dde5f, 32'h4296dbda, 32'h40ad9221, 32'h0, 32'h41863ce3, 32'h41bc42b0, 32'h0, 32'h4267eb36};
test_input[11344:11351] = '{32'hc28c8cc8, 32'h42bed431, 32'hc1b33ff7, 32'hc1c353b1, 32'hc12b0b3f, 32'hc29b56d6, 32'h42aae3bd, 32'h41e0dddf};
test_output[11344:11351] = '{32'h0, 32'h42bed431, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42aae3bd, 32'h41e0dddf};
test_input[11352:11359] = '{32'h41e0812a, 32'hc245b7d0, 32'hc1efa629, 32'h42b57f78, 32'hc21f2b23, 32'hc1cf0897, 32'hc1ac5c3c, 32'h4215748f};
test_output[11352:11359] = '{32'h41e0812a, 32'h0, 32'h0, 32'h42b57f78, 32'h0, 32'h0, 32'h0, 32'h4215748f};
test_input[11360:11367] = '{32'h424c1f7b, 32'hc10b76bd, 32'hc1027b38, 32'hc2bb7525, 32'h42b8bd5d, 32'h42806081, 32'hc22fb6b9, 32'hc2ae84b4};
test_output[11360:11367] = '{32'h424c1f7b, 32'h0, 32'h0, 32'h0, 32'h42b8bd5d, 32'h42806081, 32'h0, 32'h0};
test_input[11368:11375] = '{32'h425167e6, 32'hc27bbfa9, 32'h427fc885, 32'hc27cffe7, 32'h4236712e, 32'h419d3967, 32'h41a7d794, 32'hc28be4d4};
test_output[11368:11375] = '{32'h425167e6, 32'h0, 32'h427fc885, 32'h0, 32'h4236712e, 32'h419d3967, 32'h41a7d794, 32'h0};
test_input[11376:11383] = '{32'h4288031f, 32'hc278a672, 32'h42078e23, 32'hc1d7af8e, 32'h422365e5, 32'h41dd1536, 32'h4286b760, 32'h3fed1e43};
test_output[11376:11383] = '{32'h4288031f, 32'h0, 32'h42078e23, 32'h0, 32'h422365e5, 32'h41dd1536, 32'h4286b760, 32'h3fed1e43};
test_input[11384:11391] = '{32'h42a93d34, 32'hc295ada8, 32'h4235f1ac, 32'h41e3a96e, 32'hc2b73c0a, 32'hc1dd5562, 32'hc1ef440a, 32'h4143ba6a};
test_output[11384:11391] = '{32'h42a93d34, 32'h0, 32'h4235f1ac, 32'h41e3a96e, 32'h0, 32'h0, 32'h0, 32'h4143ba6a};
test_input[11392:11399] = '{32'hc212d773, 32'h426430a0, 32'hc2b7fefd, 32'h428943ac, 32'h426a88cf, 32'h425a0cb7, 32'hc26c311e, 32'hc15e429e};
test_output[11392:11399] = '{32'h0, 32'h426430a0, 32'h0, 32'h428943ac, 32'h426a88cf, 32'h425a0cb7, 32'h0, 32'h0};
test_input[11400:11407] = '{32'hc28d4dc8, 32'h41905c69, 32'h40f9ac13, 32'h423044b5, 32'hc23aa577, 32'hc2b8725d, 32'hc21beff8, 32'hc1ec9011};
test_output[11400:11407] = '{32'h0, 32'h41905c69, 32'h40f9ac13, 32'h423044b5, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11408:11415] = '{32'hc18d4dfb, 32'h4212eb1a, 32'hc1517b20, 32'h428ddf03, 32'hc20b1257, 32'hc2ba48bc, 32'h424e2c27, 32'h429476e8};
test_output[11408:11415] = '{32'h0, 32'h4212eb1a, 32'h0, 32'h428ddf03, 32'h0, 32'h0, 32'h424e2c27, 32'h429476e8};
test_input[11416:11423] = '{32'h41fbf928, 32'hc2bb2be7, 32'hc214fa96, 32'hc00f49f7, 32'hc2929175, 32'h42537bcd, 32'hc2a37516, 32'h4203bd66};
test_output[11416:11423] = '{32'h41fbf928, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42537bcd, 32'h0, 32'h4203bd66};
test_input[11424:11431] = '{32'h42c1edb0, 32'h40301bdc, 32'hc229ece7, 32'h4206e439, 32'hc1f16c0e, 32'hc1912c0e, 32'h42a4adcc, 32'hc2912bfb};
test_output[11424:11431] = '{32'h42c1edb0, 32'h40301bdc, 32'h0, 32'h4206e439, 32'h0, 32'h0, 32'h42a4adcc, 32'h0};
test_input[11432:11439] = '{32'hc1c52347, 32'h429981bf, 32'hc20637b3, 32'hc24e2a3b, 32'h4286d1e9, 32'h42843351, 32'h42a50187, 32'h42a06195};
test_output[11432:11439] = '{32'h0, 32'h429981bf, 32'h0, 32'h0, 32'h4286d1e9, 32'h42843351, 32'h42a50187, 32'h42a06195};
test_input[11440:11447] = '{32'h418ca212, 32'h4251d3c7, 32'h42967cf2, 32'h428a29c6, 32'h4184f6a7, 32'h42866b25, 32'h42ad3afb, 32'h4280bc99};
test_output[11440:11447] = '{32'h418ca212, 32'h4251d3c7, 32'h42967cf2, 32'h428a29c6, 32'h4184f6a7, 32'h42866b25, 32'h42ad3afb, 32'h4280bc99};
test_input[11448:11455] = '{32'hc2c40ba1, 32'h4290045b, 32'hc1576a8d, 32'hc2accaf4, 32'h42b07ab4, 32'h42bad337, 32'h4149d319, 32'hc2ab20da};
test_output[11448:11455] = '{32'h0, 32'h4290045b, 32'h0, 32'h0, 32'h42b07ab4, 32'h42bad337, 32'h4149d319, 32'h0};
test_input[11456:11463] = '{32'h42a9f766, 32'hc24cedc7, 32'hc2999960, 32'h42a282bb, 32'h423a0ff2, 32'h426b6f07, 32'hc2a6e8ad, 32'hc2a56a1b};
test_output[11456:11463] = '{32'h42a9f766, 32'h0, 32'h0, 32'h42a282bb, 32'h423a0ff2, 32'h426b6f07, 32'h0, 32'h0};
test_input[11464:11471] = '{32'hc220ffa2, 32'hc28f4d6d, 32'hc23f4676, 32'h4114f383, 32'hc2c2334d, 32'hc08d20a5, 32'h42446a98, 32'h42833d86};
test_output[11464:11471] = '{32'h0, 32'h0, 32'h0, 32'h4114f383, 32'h0, 32'h0, 32'h42446a98, 32'h42833d86};
test_input[11472:11479] = '{32'h42133bee, 32'hc2a80129, 32'hc1786ca8, 32'hc2a69436, 32'hc1f0fa55, 32'h4288f6ab, 32'hc2747d3d, 32'h428f0802};
test_output[11472:11479] = '{32'h42133bee, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4288f6ab, 32'h0, 32'h428f0802};
test_input[11480:11487] = '{32'hc27fc4bc, 32'hc24ec379, 32'hc2c2e3bb, 32'hc202a5b5, 32'h41664b73, 32'h40e94710, 32'hc221945b, 32'h41725e9e};
test_output[11480:11487] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41664b73, 32'h40e94710, 32'h0, 32'h41725e9e};
test_input[11488:11495] = '{32'hc25e0e11, 32'h3f290e1d, 32'h419f458d, 32'hc28b1638, 32'hc1c4b7b9, 32'h427fba3b, 32'h42938405, 32'h421cdf57};
test_output[11488:11495] = '{32'h0, 32'h3f290e1d, 32'h419f458d, 32'h0, 32'h0, 32'h427fba3b, 32'h42938405, 32'h421cdf57};
test_input[11496:11503] = '{32'hc20c928a, 32'h42af5b42, 32'h40d6e908, 32'h41c73efc, 32'h421866cf, 32'h42bc9eba, 32'hc14b6a95, 32'h428b5237};
test_output[11496:11503] = '{32'h0, 32'h42af5b42, 32'h40d6e908, 32'h41c73efc, 32'h421866cf, 32'h42bc9eba, 32'h0, 32'h428b5237};
test_input[11504:11511] = '{32'hc1c9d209, 32'hc28b0ae4, 32'hc22b156f, 32'h4275e180, 32'hc0834158, 32'h42713eb9, 32'h42a25911, 32'hc29be816};
test_output[11504:11511] = '{32'h0, 32'h0, 32'h0, 32'h4275e180, 32'h0, 32'h42713eb9, 32'h42a25911, 32'h0};
test_input[11512:11519] = '{32'h4244e0f0, 32'h429733f7, 32'hc2b5b1be, 32'hc2b4a86d, 32'h42957e69, 32'h425a5722, 32'hc18dc33d, 32'hc1cd98bc};
test_output[11512:11519] = '{32'h4244e0f0, 32'h429733f7, 32'h0, 32'h0, 32'h42957e69, 32'h425a5722, 32'h0, 32'h0};
test_input[11520:11527] = '{32'h40215d0a, 32'hc0bc64ad, 32'h427875b1, 32'hc28c5860, 32'hc2041275, 32'hc2998a90, 32'hc2ab1127, 32'hc2396164};
test_output[11520:11527] = '{32'h40215d0a, 32'h0, 32'h427875b1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11528:11535] = '{32'hc226e76c, 32'hc25db5e0, 32'hc2681cb4, 32'hc14ca5ab, 32'h4237ac01, 32'hc1be0290, 32'hc2777841, 32'hc145daa0};
test_output[11528:11535] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4237ac01, 32'h0, 32'h0, 32'h0};
test_input[11536:11543] = '{32'hc2c6c1e4, 32'hc29c11c4, 32'hc2c28286, 32'hc2575195, 32'h42972714, 32'hc29e4afe, 32'h40ec465d, 32'h42c0f47f};
test_output[11536:11543] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42972714, 32'h0, 32'h40ec465d, 32'h42c0f47f};
test_input[11544:11551] = '{32'h42b971c9, 32'h425ddc98, 32'h42bd98f5, 32'h421b9b14, 32'h40f166eb, 32'h42c404b2, 32'h427b325a, 32'hc0faa494};
test_output[11544:11551] = '{32'h42b971c9, 32'h425ddc98, 32'h42bd98f5, 32'h421b9b14, 32'h40f166eb, 32'h42c404b2, 32'h427b325a, 32'h0};
test_input[11552:11559] = '{32'h4296b9b7, 32'hc2b1e151, 32'hc1c7396e, 32'hc28be8e1, 32'hc092e12e, 32'h42c23cf2, 32'hc2b55971, 32'hc27f08f6};
test_output[11552:11559] = '{32'h4296b9b7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c23cf2, 32'h0, 32'h0};
test_input[11560:11567] = '{32'h42c6f795, 32'h42640a86, 32'hc2bb969b, 32'h42647eea, 32'hc2347ac9, 32'hc20e331a, 32'hc1bec9bb, 32'h423dea3d};
test_output[11560:11567] = '{32'h42c6f795, 32'h42640a86, 32'h0, 32'h42647eea, 32'h0, 32'h0, 32'h0, 32'h423dea3d};
test_input[11568:11575] = '{32'h42b8619a, 32'hc19d39a2, 32'hc290b165, 32'h407e8aca, 32'hc2853cf7, 32'hc2c028ac, 32'hc298d57b, 32'hc1ff54fc};
test_output[11568:11575] = '{32'h42b8619a, 32'h0, 32'h0, 32'h407e8aca, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11576:11583] = '{32'h42625f15, 32'h42bb791c, 32'h414a1ce2, 32'hc1064d02, 32'hc21b7450, 32'h42419c3f, 32'hc2aab7d7, 32'hc20cf938};
test_output[11576:11583] = '{32'h42625f15, 32'h42bb791c, 32'h414a1ce2, 32'h0, 32'h0, 32'h42419c3f, 32'h0, 32'h0};
test_input[11584:11591] = '{32'hc1bced77, 32'h429f3299, 32'h415c6d24, 32'hc119a1eb, 32'hc2771e60, 32'h42bcf7b4, 32'hc1a8d29e, 32'h41d80523};
test_output[11584:11591] = '{32'h0, 32'h429f3299, 32'h415c6d24, 32'h0, 32'h0, 32'h42bcf7b4, 32'h0, 32'h41d80523};
test_input[11592:11599] = '{32'hc297f29e, 32'h424d1c1f, 32'hc23ebb80, 32'h4294cc3b, 32'h42043d2a, 32'h42b345c6, 32'h41d9691a, 32'h4241326c};
test_output[11592:11599] = '{32'h0, 32'h424d1c1f, 32'h0, 32'h4294cc3b, 32'h42043d2a, 32'h42b345c6, 32'h41d9691a, 32'h4241326c};
test_input[11600:11607] = '{32'hc2861900, 32'hc2903408, 32'h4086d973, 32'hc24b59e7, 32'h41dbb902, 32'h41856713, 32'h428de6d0, 32'hc1c54472};
test_output[11600:11607] = '{32'h0, 32'h0, 32'h4086d973, 32'h0, 32'h41dbb902, 32'h41856713, 32'h428de6d0, 32'h0};
test_input[11608:11615] = '{32'h424510e4, 32'h42143034, 32'h42ba7879, 32'hc212ef16, 32'hc2c4e172, 32'hc2857d41, 32'hc1c6a442, 32'h42af35cd};
test_output[11608:11615] = '{32'h424510e4, 32'h42143034, 32'h42ba7879, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42af35cd};
test_input[11616:11623] = '{32'h3e7bf543, 32'hc20c054f, 32'hc2ba9d54, 32'h425227db, 32'hc2506584, 32'h3fa35a3a, 32'hc221fc7d, 32'h408a02ad};
test_output[11616:11623] = '{32'h3e7bf543, 32'h0, 32'h0, 32'h425227db, 32'h0, 32'h3fa35a3a, 32'h0, 32'h408a02ad};
test_input[11624:11631] = '{32'hc2985724, 32'hc253708e, 32'h41350c29, 32'hc2262a6c, 32'h422a8180, 32'h42c390d3, 32'hc27d23de, 32'h4229ab57};
test_output[11624:11631] = '{32'h0, 32'h0, 32'h41350c29, 32'h0, 32'h422a8180, 32'h42c390d3, 32'h0, 32'h4229ab57};
test_input[11632:11639] = '{32'hc1e721be, 32'h4254b47b, 32'h42a1893f, 32'hc1a1a5b2, 32'hc2bda19e, 32'hc25ba447, 32'hc2846dc9, 32'hc20730bc};
test_output[11632:11639] = '{32'h0, 32'h4254b47b, 32'h42a1893f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11640:11647] = '{32'h42c380c6, 32'hc12f22e2, 32'h41929322, 32'h42c2319c, 32'h42966ad4, 32'hc2428e21, 32'h4035e140, 32'hc274a61b};
test_output[11640:11647] = '{32'h42c380c6, 32'h0, 32'h41929322, 32'h42c2319c, 32'h42966ad4, 32'h0, 32'h4035e140, 32'h0};
test_input[11648:11655] = '{32'hc201ed11, 32'h40f31a95, 32'hc2051511, 32'hc27c4f85, 32'h423e529b, 32'hc219ee25, 32'h42982b18, 32'hc278a02c};
test_output[11648:11655] = '{32'h0, 32'h40f31a95, 32'h0, 32'h0, 32'h423e529b, 32'h0, 32'h42982b18, 32'h0};
test_input[11656:11663] = '{32'h4052300b, 32'h429ca013, 32'h4289dee1, 32'hc1aa1643, 32'hc20815eb, 32'hc15462be, 32'h42b502ab, 32'hc27c8296};
test_output[11656:11663] = '{32'h4052300b, 32'h429ca013, 32'h4289dee1, 32'h0, 32'h0, 32'h0, 32'h42b502ab, 32'h0};
test_input[11664:11671] = '{32'hc29a9b2b, 32'h42bfe015, 32'hc0481ba8, 32'h4295f6f9, 32'hc20efeca, 32'hc112a616, 32'h41d2a318, 32'hc258c6af};
test_output[11664:11671] = '{32'h0, 32'h42bfe015, 32'h0, 32'h4295f6f9, 32'h0, 32'h0, 32'h41d2a318, 32'h0};
test_input[11672:11679] = '{32'h42b01805, 32'hc18024c0, 32'h42696fab, 32'h412f171e, 32'hc2810dbf, 32'h426a0597, 32'hc250ad9b, 32'h429471f3};
test_output[11672:11679] = '{32'h42b01805, 32'h0, 32'h42696fab, 32'h412f171e, 32'h0, 32'h426a0597, 32'h0, 32'h429471f3};
test_input[11680:11687] = '{32'h428a2b58, 32'h41dc5f88, 32'hc289c431, 32'hc1382df8, 32'h418a49ab, 32'hc26ce4d9, 32'h4265f7b2, 32'hc2c4dae5};
test_output[11680:11687] = '{32'h428a2b58, 32'h41dc5f88, 32'h0, 32'h0, 32'h418a49ab, 32'h0, 32'h4265f7b2, 32'h0};
test_input[11688:11695] = '{32'h420ad912, 32'h423990eb, 32'h4232251c, 32'h42108f37, 32'hc1e95c41, 32'h42a01842, 32'h41df96c2, 32'hc2ba4a32};
test_output[11688:11695] = '{32'h420ad912, 32'h423990eb, 32'h4232251c, 32'h42108f37, 32'h0, 32'h42a01842, 32'h41df96c2, 32'h0};
test_input[11696:11703] = '{32'h4280973e, 32'h41f8c509, 32'hc21fe325, 32'hc23e4b08, 32'hc18cc6a0, 32'h426e202d, 32'h416b6712, 32'hc28356cc};
test_output[11696:11703] = '{32'h4280973e, 32'h41f8c509, 32'h0, 32'h0, 32'h0, 32'h426e202d, 32'h416b6712, 32'h0};
test_input[11704:11711] = '{32'h429ce872, 32'h42b7eea9, 32'h41b3f013, 32'hc2a22d46, 32'h42293c31, 32'hc2b1b951, 32'h42bd83e7, 32'h42bfa009};
test_output[11704:11711] = '{32'h429ce872, 32'h42b7eea9, 32'h41b3f013, 32'h0, 32'h42293c31, 32'h0, 32'h42bd83e7, 32'h42bfa009};
test_input[11712:11719] = '{32'hc2a2a0fb, 32'hc2b53cb0, 32'hc2870ace, 32'h429f33de, 32'h42012041, 32'h422a4752, 32'hc2b9787f, 32'h4213a87e};
test_output[11712:11719] = '{32'h0, 32'h0, 32'h0, 32'h429f33de, 32'h42012041, 32'h422a4752, 32'h0, 32'h4213a87e};
test_input[11720:11727] = '{32'hc2ae8cd5, 32'hbeb36580, 32'h42a3c4c6, 32'h42ba33f4, 32'hc0da98d4, 32'h40fc8b75, 32'h419a4d51, 32'h41a05f4b};
test_output[11720:11727] = '{32'h0, 32'h0, 32'h42a3c4c6, 32'h42ba33f4, 32'h0, 32'h40fc8b75, 32'h419a4d51, 32'h41a05f4b};
test_input[11728:11735] = '{32'h42c7b715, 32'hc2abc76c, 32'h427b08ba, 32'hc11c399a, 32'hc25f2556, 32'h42772858, 32'hc2844ced, 32'h4202aec2};
test_output[11728:11735] = '{32'h42c7b715, 32'h0, 32'h427b08ba, 32'h0, 32'h0, 32'h42772858, 32'h0, 32'h4202aec2};
test_input[11736:11743] = '{32'h423f1cea, 32'h41f22afb, 32'h428ffa2c, 32'h42aad1db, 32'hc25a1023, 32'hc2af4b62, 32'hc19d4001, 32'hc1f8a578};
test_output[11736:11743] = '{32'h423f1cea, 32'h41f22afb, 32'h428ffa2c, 32'h42aad1db, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11744:11751] = '{32'hc1c1a5a0, 32'h428918d2, 32'h3f0774a0, 32'hc1b95ed2, 32'h4238520e, 32'hc1412f29, 32'h4285417e, 32'hc274134d};
test_output[11744:11751] = '{32'h0, 32'h428918d2, 32'h3f0774a0, 32'h0, 32'h4238520e, 32'h0, 32'h4285417e, 32'h0};
test_input[11752:11759] = '{32'h42257331, 32'hc2c7df79, 32'h419738fc, 32'hc2c66305, 32'h42243b74, 32'h4222d036, 32'h429237e0, 32'h421569ae};
test_output[11752:11759] = '{32'h42257331, 32'h0, 32'h419738fc, 32'h0, 32'h42243b74, 32'h4222d036, 32'h429237e0, 32'h421569ae};
test_input[11760:11767] = '{32'h4294c35d, 32'hc26a8094, 32'hc1eb2306, 32'hc21ab6c4, 32'hc1d71a30, 32'hc26779d8, 32'h42c7bb0c, 32'h41046b31};
test_output[11760:11767] = '{32'h4294c35d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c7bb0c, 32'h41046b31};
test_input[11768:11775] = '{32'hc2a64bbd, 32'h41a0bcc2, 32'h40c14c6a, 32'h42377887, 32'h420a3ef9, 32'h42bbed29, 32'h4143f3c0, 32'hc1d105ad};
test_output[11768:11775] = '{32'h0, 32'h41a0bcc2, 32'h40c14c6a, 32'h42377887, 32'h420a3ef9, 32'h42bbed29, 32'h4143f3c0, 32'h0};
test_input[11776:11783] = '{32'h42667910, 32'h42bc476f, 32'h421b057d, 32'hc1e79d9c, 32'h4215447e, 32'h42b10eeb, 32'hc2863ec7, 32'h42a75877};
test_output[11776:11783] = '{32'h42667910, 32'h42bc476f, 32'h421b057d, 32'h0, 32'h4215447e, 32'h42b10eeb, 32'h0, 32'h42a75877};
test_input[11784:11791] = '{32'h42926601, 32'h4285bbe5, 32'hc25a320a, 32'h40af1bac, 32'hc1aa4ef2, 32'h4204f7bf, 32'h4217b5d2, 32'hc1effd1a};
test_output[11784:11791] = '{32'h42926601, 32'h4285bbe5, 32'h0, 32'h40af1bac, 32'h0, 32'h4204f7bf, 32'h4217b5d2, 32'h0};
test_input[11792:11799] = '{32'hc17d90e0, 32'hc1cf9db0, 32'h42c416a7, 32'h41609dc5, 32'h427c5b05, 32'hbffe7412, 32'h425c800b, 32'hc2c39fed};
test_output[11792:11799] = '{32'h0, 32'h0, 32'h42c416a7, 32'h41609dc5, 32'h427c5b05, 32'h0, 32'h425c800b, 32'h0};
test_input[11800:11807] = '{32'hc240f8a4, 32'h410bcdf9, 32'h417995a0, 32'h41fbb6e2, 32'h42762dfc, 32'h429354aa, 32'hc25ca71a, 32'hc1efffa5};
test_output[11800:11807] = '{32'h0, 32'h410bcdf9, 32'h417995a0, 32'h41fbb6e2, 32'h42762dfc, 32'h429354aa, 32'h0, 32'h0};
test_input[11808:11815] = '{32'h426e2370, 32'hc295f0cb, 32'h40cbdadc, 32'hc189c778, 32'hc25c656b, 32'hc209d2cf, 32'hc28d4bca, 32'h427fa6ef};
test_output[11808:11815] = '{32'h426e2370, 32'h0, 32'h40cbdadc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427fa6ef};
test_input[11816:11823] = '{32'h4235bdb3, 32'h42a12be8, 32'h42c027ec, 32'h42bf8cb2, 32'hc27d470c, 32'h4296241f, 32'hc1a87056, 32'hc2a31857};
test_output[11816:11823] = '{32'h4235bdb3, 32'h42a12be8, 32'h42c027ec, 32'h42bf8cb2, 32'h0, 32'h4296241f, 32'h0, 32'h0};
test_input[11824:11831] = '{32'hc25ae2b7, 32'h42c06d9d, 32'h42304731, 32'h4032a43d, 32'hc296b240, 32'hc236fe1c, 32'hc2bc3377, 32'h42a292ad};
test_output[11824:11831] = '{32'h0, 32'h42c06d9d, 32'h42304731, 32'h4032a43d, 32'h0, 32'h0, 32'h0, 32'h42a292ad};
test_input[11832:11839] = '{32'hc2067f89, 32'hc24de751, 32'hc1ed8d36, 32'hc10b9c4d, 32'h408ab5d7, 32'h4205b98c, 32'h4274d54e, 32'hc10fe5d9};
test_output[11832:11839] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h408ab5d7, 32'h4205b98c, 32'h4274d54e, 32'h0};
test_input[11840:11847] = '{32'h42bec76b, 32'h42a615c6, 32'h417d22d1, 32'hc1dd5600, 32'h4277d39e, 32'h42ad85b9, 32'h41b4b5d4, 32'hc0ff7265};
test_output[11840:11847] = '{32'h42bec76b, 32'h42a615c6, 32'h417d22d1, 32'h0, 32'h4277d39e, 32'h42ad85b9, 32'h41b4b5d4, 32'h0};
test_input[11848:11855] = '{32'h420d8896, 32'hc2a9d23f, 32'h42aaaa66, 32'hc2070c63, 32'hc29781e8, 32'h42976186, 32'hc24406cf, 32'h42621717};
test_output[11848:11855] = '{32'h420d8896, 32'h0, 32'h42aaaa66, 32'h0, 32'h0, 32'h42976186, 32'h0, 32'h42621717};
test_input[11856:11863] = '{32'h428285fd, 32'h428c3faf, 32'h423f0049, 32'h42abc93c, 32'h428bd146, 32'hc212ed3b, 32'h429a3834, 32'h40d709a8};
test_output[11856:11863] = '{32'h428285fd, 32'h428c3faf, 32'h423f0049, 32'h42abc93c, 32'h428bd146, 32'h0, 32'h429a3834, 32'h40d709a8};
test_input[11864:11871] = '{32'h4250c774, 32'hc2c62884, 32'hc2621eb5, 32'hc23632c1, 32'h42395586, 32'hc2992dc2, 32'h42b87fcd, 32'hc2874760};
test_output[11864:11871] = '{32'h4250c774, 32'h0, 32'h0, 32'h0, 32'h42395586, 32'h0, 32'h42b87fcd, 32'h0};
test_input[11872:11879] = '{32'h429da8a3, 32'h424651f6, 32'h4153ed29, 32'hc2b087fb, 32'hc28021b3, 32'hc2a2a78f, 32'h429dc818, 32'hc1becbfe};
test_output[11872:11879] = '{32'h429da8a3, 32'h424651f6, 32'h4153ed29, 32'h0, 32'h0, 32'h0, 32'h429dc818, 32'h0};
test_input[11880:11887] = '{32'h4286dbf4, 32'h4251c020, 32'hc2b085c8, 32'h42c1027e, 32'h426a4850, 32'h420161b1, 32'h40b37962, 32'hc2124ffc};
test_output[11880:11887] = '{32'h4286dbf4, 32'h4251c020, 32'h0, 32'h42c1027e, 32'h426a4850, 32'h420161b1, 32'h40b37962, 32'h0};
test_input[11888:11895] = '{32'h40bf0026, 32'h42455dd8, 32'h428f7cb3, 32'h42a878c1, 32'hc28df158, 32'h42c35a3b, 32'hc2861e43, 32'hc2789839};
test_output[11888:11895] = '{32'h40bf0026, 32'h42455dd8, 32'h428f7cb3, 32'h42a878c1, 32'h0, 32'h42c35a3b, 32'h0, 32'h0};
test_input[11896:11903] = '{32'h429cb5ac, 32'h41ffb076, 32'hc22cdad9, 32'h4288e9f6, 32'hc2a113f5, 32'hc2843f11, 32'hc2646a9f, 32'hc29fa177};
test_output[11896:11903] = '{32'h429cb5ac, 32'h41ffb076, 32'h0, 32'h4288e9f6, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11904:11911] = '{32'hc1920a86, 32'h4296e47d, 32'h428b9077, 32'hc2608f3a, 32'hc225c8d6, 32'hc2a42443, 32'hc2825d60, 32'hc2377423};
test_output[11904:11911] = '{32'h0, 32'h4296e47d, 32'h428b9077, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11912:11919] = '{32'h42b499d6, 32'h41dd7d57, 32'hc26f3cef, 32'hc2babb2c, 32'hc244a83e, 32'h426f2056, 32'h41f2f1ea, 32'h41d7ccf7};
test_output[11912:11919] = '{32'h42b499d6, 32'h41dd7d57, 32'h0, 32'h0, 32'h0, 32'h426f2056, 32'h41f2f1ea, 32'h41d7ccf7};
test_input[11920:11927] = '{32'hc2553e2d, 32'h41c79faf, 32'h42a2244a, 32'hc2a7400f, 32'h403b1939, 32'h419de7d6, 32'hc0e4222a, 32'h427ae43d};
test_output[11920:11927] = '{32'h0, 32'h41c79faf, 32'h42a2244a, 32'h0, 32'h403b1939, 32'h419de7d6, 32'h0, 32'h427ae43d};
test_input[11928:11935] = '{32'hc20bf76b, 32'hc1abe3b5, 32'h4232bab4, 32'hc10e76fb, 32'hc2b50687, 32'h42258a9e, 32'hc298c65f, 32'hc2045dc1};
test_output[11928:11935] = '{32'h0, 32'h0, 32'h4232bab4, 32'h0, 32'h0, 32'h42258a9e, 32'h0, 32'h0};
test_input[11936:11943] = '{32'h4240ddaa, 32'hc2053fac, 32'h427e9ef8, 32'hc2ad870c, 32'hc2bcbef8, 32'h3da3b323, 32'hc29b4cfd, 32'hc050b565};
test_output[11936:11943] = '{32'h4240ddaa, 32'h0, 32'h427e9ef8, 32'h0, 32'h0, 32'h3da3b323, 32'h0, 32'h0};
test_input[11944:11951] = '{32'hc2770f65, 32'hc19df2ba, 32'h42816049, 32'hc2b69b17, 32'hc24fa683, 32'h41ec8563, 32'h41c6d6f0, 32'hc2957e2a};
test_output[11944:11951] = '{32'h0, 32'h0, 32'h42816049, 32'h0, 32'h0, 32'h41ec8563, 32'h41c6d6f0, 32'h0};
test_input[11952:11959] = '{32'h42927a82, 32'hc1020a43, 32'hc24c8f08, 32'h422e95b3, 32'h42b49f54, 32'hc1e28858, 32'hc2b75160, 32'hc2612702};
test_output[11952:11959] = '{32'h42927a82, 32'h0, 32'h0, 32'h422e95b3, 32'h42b49f54, 32'h0, 32'h0, 32'h0};
test_input[11960:11967] = '{32'h4266e8b7, 32'hc23f4756, 32'h423b53f8, 32'h42559d1b, 32'hc28cd61d, 32'h42b2cc2b, 32'hc1a1859b, 32'h42c42726};
test_output[11960:11967] = '{32'h4266e8b7, 32'h0, 32'h423b53f8, 32'h42559d1b, 32'h0, 32'h42b2cc2b, 32'h0, 32'h42c42726};
test_input[11968:11975] = '{32'hc2ae62db, 32'hc1cb6e89, 32'hc243c00f, 32'h428398db, 32'hc2a83f11, 32'h42ab5da9, 32'h420b0c7e, 32'h42991622};
test_output[11968:11975] = '{32'h0, 32'h0, 32'h0, 32'h428398db, 32'h0, 32'h42ab5da9, 32'h420b0c7e, 32'h42991622};
test_input[11976:11983] = '{32'h42b711c6, 32'hc2812256, 32'h3fc7b879, 32'hbec42e3d, 32'h428ab3f8, 32'h42b2a1bc, 32'hc1a9d700, 32'h420467ab};
test_output[11976:11983] = '{32'h42b711c6, 32'h0, 32'h3fc7b879, 32'h0, 32'h428ab3f8, 32'h42b2a1bc, 32'h0, 32'h420467ab};
test_input[11984:11991] = '{32'hc20636c9, 32'h42a82bb1, 32'h4211dc1d, 32'h421cfa77, 32'hc1ffd73f, 32'hc2843690, 32'hc2bdcabc, 32'hc2c08131};
test_output[11984:11991] = '{32'h0, 32'h42a82bb1, 32'h4211dc1d, 32'h421cfa77, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[11992:11999] = '{32'hc2c06d4c, 32'h405b2ba2, 32'h424b5f10, 32'h42040214, 32'h420dab27, 32'h4246fce2, 32'hc17cbd4b, 32'h411ef663};
test_output[11992:11999] = '{32'h0, 32'h405b2ba2, 32'h424b5f10, 32'h42040214, 32'h420dab27, 32'h4246fce2, 32'h0, 32'h411ef663};
test_input[12000:12007] = '{32'hc226e31c, 32'h3e14d671, 32'hc12f506f, 32'hc1a888ea, 32'hc28e7348, 32'hc1fd6bff, 32'hc1c6dbc3, 32'h429e1ad6};
test_output[12000:12007] = '{32'h0, 32'h3e14d671, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429e1ad6};
test_input[12008:12015] = '{32'h4246ca3b, 32'hc2644c22, 32'hc2a5dd87, 32'h40c24c70, 32'h40c7e5e4, 32'h42b187a7, 32'hc2b867b2, 32'hc04a242d};
test_output[12008:12015] = '{32'h4246ca3b, 32'h0, 32'h0, 32'h40c24c70, 32'h40c7e5e4, 32'h42b187a7, 32'h0, 32'h0};
test_input[12016:12023] = '{32'h41ceb2e0, 32'hc27bb1b3, 32'hc2825d5a, 32'h400ff2b8, 32'hc1a857a0, 32'hc2b1d921, 32'h4207e00b, 32'hc261cf11};
test_output[12016:12023] = '{32'h41ceb2e0, 32'h0, 32'h0, 32'h400ff2b8, 32'h0, 32'h0, 32'h4207e00b, 32'h0};
test_input[12024:12031] = '{32'h4206bdbd, 32'h42332584, 32'hc2820940, 32'hc246d4d5, 32'hc25393ad, 32'h414dfbbf, 32'h42b78fa3, 32'h41cdade6};
test_output[12024:12031] = '{32'h4206bdbd, 32'h42332584, 32'h0, 32'h0, 32'h0, 32'h414dfbbf, 32'h42b78fa3, 32'h41cdade6};
test_input[12032:12039] = '{32'h4286d610, 32'h422d289c, 32'hc2abab44, 32'h41c6f530, 32'h42aec3a6, 32'h42290a59, 32'hc249bac5, 32'h3fded7df};
test_output[12032:12039] = '{32'h4286d610, 32'h422d289c, 32'h0, 32'h41c6f530, 32'h42aec3a6, 32'h42290a59, 32'h0, 32'h3fded7df};
test_input[12040:12047] = '{32'h42039abc, 32'h423625c4, 32'hc2c582fe, 32'h42c474ee, 32'hc22d1159, 32'h41d0d9cd, 32'hc2b1d742, 32'h41c2ce0e};
test_output[12040:12047] = '{32'h42039abc, 32'h423625c4, 32'h0, 32'h42c474ee, 32'h0, 32'h41d0d9cd, 32'h0, 32'h41c2ce0e};
test_input[12048:12055] = '{32'h403b009f, 32'h4224e678, 32'h4261a94c, 32'h419b529b, 32'hc0f04a54, 32'hc2a84f84, 32'hc23e75cf, 32'hc129d6fe};
test_output[12048:12055] = '{32'h403b009f, 32'h4224e678, 32'h4261a94c, 32'h419b529b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12056:12063] = '{32'h42abfb8f, 32'hc289d443, 32'hc1d1c291, 32'h42bad1fd, 32'h4282195b, 32'h42c0a6ae, 32'h42b10629, 32'h41cd9cf0};
test_output[12056:12063] = '{32'h42abfb8f, 32'h0, 32'h0, 32'h42bad1fd, 32'h4282195b, 32'h42c0a6ae, 32'h42b10629, 32'h41cd9cf0};
test_input[12064:12071] = '{32'h42820c16, 32'h41d155bb, 32'hc1dceebc, 32'hc288f07c, 32'hc1df57c3, 32'hc29c964c, 32'h400af323, 32'hc2631068};
test_output[12064:12071] = '{32'h42820c16, 32'h41d155bb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h400af323, 32'h0};
test_input[12072:12079] = '{32'h42b9aa8e, 32'hc2275c7a, 32'hc1edad3e, 32'hc1b997ca, 32'hc2a330c2, 32'h42640e52, 32'h42083852, 32'h4141ac9a};
test_output[12072:12079] = '{32'h42b9aa8e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42640e52, 32'h42083852, 32'h4141ac9a};
test_input[12080:12087] = '{32'hc12f8cc0, 32'hc28f120a, 32'h40725da9, 32'h4167105c, 32'h4180bd41, 32'hc1dfcc05, 32'h41fffc0a, 32'hc1f627f9};
test_output[12080:12087] = '{32'h0, 32'h0, 32'h40725da9, 32'h4167105c, 32'h4180bd41, 32'h0, 32'h41fffc0a, 32'h0};
test_input[12088:12095] = '{32'hc29931d2, 32'hc2507eec, 32'hc2986b46, 32'hc21bf281, 32'hc29c91ff, 32'h4256b8aa, 32'hc1b94b9a, 32'hc260c0dc};
test_output[12088:12095] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4256b8aa, 32'h0, 32'h0};
test_input[12096:12103] = '{32'hc1710e22, 32'hc29b7810, 32'h4220190f, 32'hc126d55d, 32'hc25503e3, 32'hc19b7239, 32'h4271f59f, 32'hc0c72622};
test_output[12096:12103] = '{32'h0, 32'h0, 32'h4220190f, 32'h0, 32'h0, 32'h0, 32'h4271f59f, 32'h0};
test_input[12104:12111] = '{32'h42489772, 32'hc2897558, 32'hc20ab4dc, 32'h426d576c, 32'h42af2e72, 32'hc2c032a8, 32'h423bfc80, 32'hc1d20e4f};
test_output[12104:12111] = '{32'h42489772, 32'h0, 32'h0, 32'h426d576c, 32'h42af2e72, 32'h0, 32'h423bfc80, 32'h0};
test_input[12112:12119] = '{32'h42864c58, 32'h40cd434c, 32'hc2743673, 32'h421c811a, 32'hc20bff39, 32'hc29d3e7b, 32'hc282f6c0, 32'h4136a00d};
test_output[12112:12119] = '{32'h42864c58, 32'h40cd434c, 32'h0, 32'h421c811a, 32'h0, 32'h0, 32'h0, 32'h4136a00d};
test_input[12120:12127] = '{32'hc296729f, 32'h4216a143, 32'h42ab57cc, 32'h426b8eeb, 32'hc235e47a, 32'hc14321ca, 32'hc2a51fcf, 32'hc2b8533f};
test_output[12120:12127] = '{32'h0, 32'h4216a143, 32'h42ab57cc, 32'h426b8eeb, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12128:12135] = '{32'hc1375f38, 32'hc1b42d77, 32'hc233216c, 32'h42992119, 32'h428b1aaa, 32'h4268376e, 32'h42b6c693, 32'h42b69cfe};
test_output[12128:12135] = '{32'h0, 32'h0, 32'h0, 32'h42992119, 32'h428b1aaa, 32'h4268376e, 32'h42b6c693, 32'h42b69cfe};
test_input[12136:12143] = '{32'hc1cc138a, 32'h423346ee, 32'h429361e1, 32'hc2265505, 32'hc2b9b60b, 32'hc2b7cd0c, 32'h429e765b, 32'h426a171d};
test_output[12136:12143] = '{32'h0, 32'h423346ee, 32'h429361e1, 32'h0, 32'h0, 32'h0, 32'h429e765b, 32'h426a171d};
test_input[12144:12151] = '{32'h42208f73, 32'hc28971e6, 32'h42a320f4, 32'h411add8b, 32'hc23f4ba4, 32'h42318efa, 32'h42b5fb72, 32'h4249dc86};
test_output[12144:12151] = '{32'h42208f73, 32'h0, 32'h42a320f4, 32'h411add8b, 32'h0, 32'h42318efa, 32'h42b5fb72, 32'h4249dc86};
test_input[12152:12159] = '{32'h40930888, 32'hbf05a8cf, 32'hc2b07e4d, 32'h428f80db, 32'h42c4de8e, 32'h42bde5b0, 32'h42866dcc, 32'hc20223bd};
test_output[12152:12159] = '{32'h40930888, 32'h0, 32'h0, 32'h428f80db, 32'h42c4de8e, 32'h42bde5b0, 32'h42866dcc, 32'h0};
test_input[12160:12167] = '{32'hc29c6a52, 32'hc25b90a8, 32'hc106c2aa, 32'h4238f4f5, 32'h424296d1, 32'hc25fbfc7, 32'hc1c9bd6d, 32'h41b5205c};
test_output[12160:12167] = '{32'h0, 32'h0, 32'h0, 32'h4238f4f5, 32'h424296d1, 32'h0, 32'h0, 32'h41b5205c};
test_input[12168:12175] = '{32'h4280d492, 32'hc132268f, 32'hc262bfad, 32'hc1ca4d3b, 32'hc28bf6ad, 32'h428340fb, 32'hc26b8af3, 32'hc292d4d9};
test_output[12168:12175] = '{32'h4280d492, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428340fb, 32'h0, 32'h0};
test_input[12176:12183] = '{32'h4006ff70, 32'hc29cd2a8, 32'hc2735414, 32'hc1ae620e, 32'h42bb1c7a, 32'hc29d24ea, 32'hc23f037a, 32'h426f5b31};
test_output[12176:12183] = '{32'h4006ff70, 32'h0, 32'h0, 32'h0, 32'h42bb1c7a, 32'h0, 32'h0, 32'h426f5b31};
test_input[12184:12191] = '{32'hc2942452, 32'hc29159a2, 32'hc1fbb7e0, 32'hbf93c107, 32'h422297a8, 32'h41c8a276, 32'hc2a6f88d, 32'hc2720cd7};
test_output[12184:12191] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h422297a8, 32'h41c8a276, 32'h0, 32'h0};
test_input[12192:12199] = '{32'hc1b8a00b, 32'hc2410b9a, 32'hc242431f, 32'h40dc4d84, 32'hc126f0ae, 32'hc1c2a243, 32'h420f1344, 32'h428ca636};
test_output[12192:12199] = '{32'h0, 32'h0, 32'h0, 32'h40dc4d84, 32'h0, 32'h0, 32'h420f1344, 32'h428ca636};
test_input[12200:12207] = '{32'hc18b629d, 32'h42bcd42b, 32'h41dbc09b, 32'h428921e3, 32'h42206c7b, 32'hc03f8d06, 32'hc212f53b, 32'h41cfe20f};
test_output[12200:12207] = '{32'h0, 32'h42bcd42b, 32'h41dbc09b, 32'h428921e3, 32'h42206c7b, 32'h0, 32'h0, 32'h41cfe20f};
test_input[12208:12215] = '{32'h4292d5b8, 32'h42c394fb, 32'hc2aa669d, 32'hc29756a2, 32'hc29dae95, 32'hc18e57cd, 32'hc26139c2, 32'h40cc4188};
test_output[12208:12215] = '{32'h4292d5b8, 32'h42c394fb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40cc4188};
test_input[12216:12223] = '{32'hc2742a03, 32'hc136860c, 32'h41c02dff, 32'hc29b29c6, 32'h4006829f, 32'hc10a65fa, 32'h41997872, 32'h41f42a0f};
test_output[12216:12223] = '{32'h0, 32'h0, 32'h41c02dff, 32'h0, 32'h4006829f, 32'h0, 32'h41997872, 32'h41f42a0f};
test_input[12224:12231] = '{32'hc1a94f40, 32'hc245583f, 32'h4205a27b, 32'hc26cc243, 32'h42949637, 32'hc1c3ad82, 32'hc032a000, 32'h42714404};
test_output[12224:12231] = '{32'h0, 32'h0, 32'h4205a27b, 32'h0, 32'h42949637, 32'h0, 32'h0, 32'h42714404};
test_input[12232:12239] = '{32'hc2494393, 32'hc28d9aff, 32'h4223ce19, 32'hc2b8c866, 32'h40c58392, 32'hc217a388, 32'h419412d2, 32'hc29b0357};
test_output[12232:12239] = '{32'h0, 32'h0, 32'h4223ce19, 32'h0, 32'h40c58392, 32'h0, 32'h419412d2, 32'h0};
test_input[12240:12247] = '{32'hc1a5a6c2, 32'hc28acdef, 32'h42a6bed5, 32'hc2bacc29, 32'hc0d9e1d6, 32'hc0943b60, 32'h423143bd, 32'hc21c98d0};
test_output[12240:12247] = '{32'h0, 32'h0, 32'h42a6bed5, 32'h0, 32'h0, 32'h0, 32'h423143bd, 32'h0};
test_input[12248:12255] = '{32'hc1dd1a0b, 32'hc225a05b, 32'hc2264e03, 32'h42acdcca, 32'h42c58467, 32'h42948d82, 32'hc2633d9b, 32'hc2336ea9};
test_output[12248:12255] = '{32'h0, 32'h0, 32'h0, 32'h42acdcca, 32'h42c58467, 32'h42948d82, 32'h0, 32'h0};
test_input[12256:12263] = '{32'h42826835, 32'hc1db8e22, 32'h422139f6, 32'h42847926, 32'hc2c291d4, 32'h41d060ed, 32'hc295f71d, 32'h42a67ce1};
test_output[12256:12263] = '{32'h42826835, 32'h0, 32'h422139f6, 32'h42847926, 32'h0, 32'h41d060ed, 32'h0, 32'h42a67ce1};
test_input[12264:12271] = '{32'h417446b9, 32'hc1a4c88c, 32'h42204b79, 32'hc2817632, 32'hc25bea02, 32'h42577f86, 32'hc25aa87b, 32'h429118df};
test_output[12264:12271] = '{32'h417446b9, 32'h0, 32'h42204b79, 32'h0, 32'h0, 32'h42577f86, 32'h0, 32'h429118df};
test_input[12272:12279] = '{32'hc108e0d2, 32'hc22b112e, 32'hc28c8e38, 32'h429922f1, 32'hc07a90ce, 32'hc2af92cb, 32'hc20ca92c, 32'hc268a7ad};
test_output[12272:12279] = '{32'h0, 32'h0, 32'h0, 32'h429922f1, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12280:12287] = '{32'hc2ae094c, 32'hc11573c3, 32'hc2a86f3b, 32'hc1680271, 32'hc21566ce, 32'h42a01a88, 32'h41e76b83, 32'h41fe9ecf};
test_output[12280:12287] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a01a88, 32'h41e76b83, 32'h41fe9ecf};
test_input[12288:12295] = '{32'hc1bcb422, 32'h40a494c7, 32'hc2983a33, 32'h41a3552d, 32'h4205d626, 32'h41521ff2, 32'h41bf9c3c, 32'h41746689};
test_output[12288:12295] = '{32'h0, 32'h40a494c7, 32'h0, 32'h41a3552d, 32'h4205d626, 32'h41521ff2, 32'h41bf9c3c, 32'h41746689};
test_input[12296:12303] = '{32'h41fcc811, 32'h42824e84, 32'hc0f228a1, 32'h421e646b, 32'h42847e3b, 32'hc06c9202, 32'h419753e8, 32'h418e4267};
test_output[12296:12303] = '{32'h41fcc811, 32'h42824e84, 32'h0, 32'h421e646b, 32'h42847e3b, 32'h0, 32'h419753e8, 32'h418e4267};
test_input[12304:12311] = '{32'h41e885af, 32'h4211cb19, 32'hc2a51b87, 32'h42881672, 32'h42636a36, 32'hc2c18f9c, 32'h42b346bb, 32'hc23fb2d0};
test_output[12304:12311] = '{32'h41e885af, 32'h4211cb19, 32'h0, 32'h42881672, 32'h42636a36, 32'h0, 32'h42b346bb, 32'h0};
test_input[12312:12319] = '{32'hc0f110e5, 32'h4243c0e1, 32'h41100e5c, 32'h418d8f38, 32'h41dbe48a, 32'h41e4d58b, 32'hc216ec97, 32'hc2acbdc1};
test_output[12312:12319] = '{32'h0, 32'h4243c0e1, 32'h41100e5c, 32'h418d8f38, 32'h41dbe48a, 32'h41e4d58b, 32'h0, 32'h0};
test_input[12320:12327] = '{32'h42a3c75f, 32'hc2ab8740, 32'h42038fb2, 32'hc2123e1a, 32'h428f5a2b, 32'hc1b63f83, 32'hc1b4d0e3, 32'hc280784d};
test_output[12320:12327] = '{32'h42a3c75f, 32'h0, 32'h42038fb2, 32'h0, 32'h428f5a2b, 32'h0, 32'h0, 32'h0};
test_input[12328:12335] = '{32'h4019a05a, 32'h42ad18a6, 32'h40f42f62, 32'h42bccaa7, 32'h3fc1f31e, 32'hc2286101, 32'hc2b9e116, 32'h42566acf};
test_output[12328:12335] = '{32'h4019a05a, 32'h42ad18a6, 32'h40f42f62, 32'h42bccaa7, 32'h3fc1f31e, 32'h0, 32'h0, 32'h42566acf};
test_input[12336:12343] = '{32'h42969124, 32'hc242eb2c, 32'h418d82d4, 32'h42262e17, 32'hc23a73ae, 32'hc19d1128, 32'h42b4b763, 32'h419b08f4};
test_output[12336:12343] = '{32'h42969124, 32'h0, 32'h418d82d4, 32'h42262e17, 32'h0, 32'h0, 32'h42b4b763, 32'h419b08f4};
test_input[12344:12351] = '{32'hc27aad8d, 32'h42652585, 32'hc2ab276f, 32'h412a8a7c, 32'h42b68eec, 32'hc235a9d1, 32'h42941c6c, 32'hc2b242b1};
test_output[12344:12351] = '{32'h0, 32'h42652585, 32'h0, 32'h412a8a7c, 32'h42b68eec, 32'h0, 32'h42941c6c, 32'h0};
test_input[12352:12359] = '{32'hc23aef5f, 32'h423d8fa9, 32'hc2a75c1d, 32'h42a1260e, 32'h4182cf80, 32'hc2803a7a, 32'hc2bfd2b1, 32'hc1f9524a};
test_output[12352:12359] = '{32'h0, 32'h423d8fa9, 32'h0, 32'h42a1260e, 32'h4182cf80, 32'h0, 32'h0, 32'h0};
test_input[12360:12367] = '{32'hc2a46ae6, 32'h429759b2, 32'h41ca8d3e, 32'hc12b0a93, 32'hc068a37b, 32'hc2bf1bf1, 32'h4299aa16, 32'hc2863d15};
test_output[12360:12367] = '{32'h0, 32'h429759b2, 32'h41ca8d3e, 32'h0, 32'h0, 32'h0, 32'h4299aa16, 32'h0};
test_input[12368:12375] = '{32'h413080e5, 32'h415e90b2, 32'hc2418e8a, 32'hc1efb8a2, 32'h42b80e12, 32'h42b08b4a, 32'h429342b4, 32'h425a9141};
test_output[12368:12375] = '{32'h413080e5, 32'h415e90b2, 32'h0, 32'h0, 32'h42b80e12, 32'h42b08b4a, 32'h429342b4, 32'h425a9141};
test_input[12376:12383] = '{32'h4295f4a0, 32'hc22e98b9, 32'hc243c699, 32'h3f240792, 32'h419f6772, 32'hc29d2d50, 32'hc2c2c3bb, 32'hc2a60295};
test_output[12376:12383] = '{32'h4295f4a0, 32'h0, 32'h0, 32'h3f240792, 32'h419f6772, 32'h0, 32'h0, 32'h0};
test_input[12384:12391] = '{32'h424c5767, 32'h42613a8d, 32'h41e8bcd3, 32'h419f9e94, 32'h4282a6ff, 32'hc22cc45e, 32'hc25c4b8b, 32'h42b1dd79};
test_output[12384:12391] = '{32'h424c5767, 32'h42613a8d, 32'h41e8bcd3, 32'h419f9e94, 32'h4282a6ff, 32'h0, 32'h0, 32'h42b1dd79};
test_input[12392:12399] = '{32'h412d9e61, 32'hc13ae52e, 32'hc24aa3e0, 32'hc1dbbf12, 32'hc2314c09, 32'hc2c60f87, 32'h41f9112a, 32'hc1f7bc3e};
test_output[12392:12399] = '{32'h412d9e61, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f9112a, 32'h0};
test_input[12400:12407] = '{32'h424d7784, 32'h41c42dc6, 32'hc08736ce, 32'hc2bfeb6b, 32'hc192e3ce, 32'h41f3b50e, 32'hc29bdc12, 32'hc2792b23};
test_output[12400:12407] = '{32'h424d7784, 32'h41c42dc6, 32'h0, 32'h0, 32'h0, 32'h41f3b50e, 32'h0, 32'h0};
test_input[12408:12415] = '{32'h4277b2d5, 32'hc19b9465, 32'hc2c6f1c7, 32'hc1c7a73c, 32'hc1ac956b, 32'hc2243df0, 32'h428eca07, 32'h41d45ebf};
test_output[12408:12415] = '{32'h4277b2d5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428eca07, 32'h41d45ebf};
test_input[12416:12423] = '{32'hc0957537, 32'h42456080, 32'h412cd00a, 32'h420fd634, 32'hc28a42c3, 32'hc29dfc12, 32'hc1e41bd5, 32'h42b9cb01};
test_output[12416:12423] = '{32'h0, 32'h42456080, 32'h412cd00a, 32'h420fd634, 32'h0, 32'h0, 32'h0, 32'h42b9cb01};
test_input[12424:12431] = '{32'hc29c3612, 32'h4155e037, 32'hc27ce77a, 32'h4122665f, 32'hc27cd375, 32'h42a50aeb, 32'h42c380c1, 32'hc1d0640f};
test_output[12424:12431] = '{32'h0, 32'h4155e037, 32'h0, 32'h4122665f, 32'h0, 32'h42a50aeb, 32'h42c380c1, 32'h0};
test_input[12432:12439] = '{32'hc2ad8e26, 32'hc29293d4, 32'h41f9113c, 32'h4085966f, 32'h4272617c, 32'hc29fd77f, 32'hbec7a268, 32'h418d332a};
test_output[12432:12439] = '{32'h0, 32'h0, 32'h41f9113c, 32'h4085966f, 32'h4272617c, 32'h0, 32'h0, 32'h418d332a};
test_input[12440:12447] = '{32'h41d6809a, 32'hc13d7aa0, 32'hc21fc8ec, 32'h42bc61cc, 32'h420fd3cf, 32'h42a2827c, 32'h424ebb7e, 32'hc28c94d8};
test_output[12440:12447] = '{32'h41d6809a, 32'h0, 32'h0, 32'h42bc61cc, 32'h420fd3cf, 32'h42a2827c, 32'h424ebb7e, 32'h0};
test_input[12448:12455] = '{32'h426c019d, 32'h418d7ad0, 32'h41d5dcfd, 32'hc2a5cb20, 32'hc2539a3d, 32'h42ad119f, 32'h41df7ded, 32'hc28a63ea};
test_output[12448:12455] = '{32'h426c019d, 32'h418d7ad0, 32'h41d5dcfd, 32'h0, 32'h0, 32'h42ad119f, 32'h41df7ded, 32'h0};
test_input[12456:12463] = '{32'h428d037b, 32'h41212140, 32'hc25ceac8, 32'hc2b26845, 32'h421945b4, 32'h4120ea15, 32'hc20164fa, 32'hc0fb0955};
test_output[12456:12463] = '{32'h428d037b, 32'h41212140, 32'h0, 32'h0, 32'h421945b4, 32'h4120ea15, 32'h0, 32'h0};
test_input[12464:12471] = '{32'h421e0dfe, 32'h420a5ee1, 32'h42b3d014, 32'hc25eef17, 32'hc2c3eb7f, 32'h40b877fb, 32'hc2b33caa, 32'h41ba2884};
test_output[12464:12471] = '{32'h421e0dfe, 32'h420a5ee1, 32'h42b3d014, 32'h0, 32'h0, 32'h40b877fb, 32'h0, 32'h41ba2884};
test_input[12472:12479] = '{32'h426de0af, 32'hc2b2819b, 32'h41b7db72, 32'hc0e07cc3, 32'hc254c903, 32'hbfdc8559, 32'hc1c447a6, 32'hc1c46ffb};
test_output[12472:12479] = '{32'h426de0af, 32'h0, 32'h41b7db72, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12480:12487] = '{32'h41aabd4a, 32'hc0094b2a, 32'h42ba9e52, 32'hc2573097, 32'hc2505660, 32'hc004c307, 32'h42860dc6, 32'h422e167e};
test_output[12480:12487] = '{32'h41aabd4a, 32'h0, 32'h42ba9e52, 32'h0, 32'h0, 32'h0, 32'h42860dc6, 32'h422e167e};
test_input[12488:12495] = '{32'hc286c275, 32'h42b46eca, 32'hc2c6e093, 32'h42538bfa, 32'hc203eaac, 32'hc2a1d88c, 32'hc1505efa, 32'h42860a71};
test_output[12488:12495] = '{32'h0, 32'h42b46eca, 32'h0, 32'h42538bfa, 32'h0, 32'h0, 32'h0, 32'h42860a71};
test_input[12496:12503] = '{32'hc271013d, 32'hc2a2b23b, 32'hc25aea0f, 32'hc26ac7c3, 32'h422fed6a, 32'h42571637, 32'hc1acb002, 32'h424c5b88};
test_output[12496:12503] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h422fed6a, 32'h42571637, 32'h0, 32'h424c5b88};
test_input[12504:12511] = '{32'h42b27c56, 32'h3f9459ab, 32'h42a80fb2, 32'hc2972461, 32'hc2212f08, 32'hc2b04b74, 32'hc1ec23dc, 32'hc2954b8d};
test_output[12504:12511] = '{32'h42b27c56, 32'h3f9459ab, 32'h42a80fb2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12512:12519] = '{32'hc246bb92, 32'hc20a9010, 32'hc2a5486f, 32'hc28e07ee, 32'h429ed140, 32'hc2757f9b, 32'hc2ad2c2b, 32'h41c88f6d};
test_output[12512:12519] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429ed140, 32'h0, 32'h0, 32'h41c88f6d};
test_input[12520:12527] = '{32'hc13da921, 32'h41c439c1, 32'hc1e7600b, 32'h4204c5f6, 32'h422258f1, 32'h42832187, 32'hc22a5abd, 32'h41f6ddb7};
test_output[12520:12527] = '{32'h0, 32'h41c439c1, 32'h0, 32'h4204c5f6, 32'h422258f1, 32'h42832187, 32'h0, 32'h41f6ddb7};
test_input[12528:12535] = '{32'hc2b31ee2, 32'h42c39bfb, 32'hc24181fe, 32'h42c45213, 32'h42b430bd, 32'hc2c085ec, 32'h42c36265, 32'h42999c10};
test_output[12528:12535] = '{32'h0, 32'h42c39bfb, 32'h0, 32'h42c45213, 32'h42b430bd, 32'h0, 32'h42c36265, 32'h42999c10};
test_input[12536:12543] = '{32'h40376716, 32'h42333bc2, 32'h42ab44ff, 32'h417054da, 32'hc12e2275, 32'hc2babcc9, 32'hc29c590a, 32'h42a5d90b};
test_output[12536:12543] = '{32'h40376716, 32'h42333bc2, 32'h42ab44ff, 32'h417054da, 32'h0, 32'h0, 32'h0, 32'h42a5d90b};
test_input[12544:12551] = '{32'hc23044d4, 32'hc287e166, 32'hc2c527f0, 32'hc29dd17b, 32'hc2b53906, 32'hc23ba309, 32'hc29b2dac, 32'h42accbe3};
test_output[12544:12551] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42accbe3};
test_input[12552:12559] = '{32'hc06da3cf, 32'hc207ca9e, 32'h42aa05d9, 32'hc2c6daa1, 32'h421ccdb8, 32'h41d85e93, 32'h422d21db, 32'hc28b669f};
test_output[12552:12559] = '{32'h0, 32'h0, 32'h42aa05d9, 32'h0, 32'h421ccdb8, 32'h41d85e93, 32'h422d21db, 32'h0};
test_input[12560:12567] = '{32'hc2bda554, 32'hc2a7d8d0, 32'hc257f794, 32'hc285c940, 32'hc19538e9, 32'h42b06dff, 32'hc0eb40ac, 32'h42a3fc29};
test_output[12560:12567] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b06dff, 32'h0, 32'h42a3fc29};
test_input[12568:12575] = '{32'hc170d10e, 32'h422a121a, 32'h4212a3d9, 32'h420f3873, 32'hc0e12d11, 32'hc2832f24, 32'hc1123737, 32'hc1afd1f8};
test_output[12568:12575] = '{32'h0, 32'h422a121a, 32'h4212a3d9, 32'h420f3873, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12576:12583] = '{32'h42c65cd5, 32'hc293995f, 32'hc1157dd2, 32'h42c00add, 32'h4289fba1, 32'h4297c6a8, 32'hc1ddcb2d, 32'hc2a24fb7};
test_output[12576:12583] = '{32'h42c65cd5, 32'h0, 32'h0, 32'h42c00add, 32'h4289fba1, 32'h4297c6a8, 32'h0, 32'h0};
test_input[12584:12591] = '{32'h421bca8a, 32'hc23e1a13, 32'hc203e974, 32'hc228528b, 32'hc1e9da97, 32'hc246331b, 32'h4241360b, 32'h42274af6};
test_output[12584:12591] = '{32'h421bca8a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4241360b, 32'h42274af6};
test_input[12592:12599] = '{32'h42775625, 32'hbff6c319, 32'hc1aafdef, 32'h41958dca, 32'h418ab2a7, 32'hc285c817, 32'h4248ca8b, 32'h4299a422};
test_output[12592:12599] = '{32'h42775625, 32'h0, 32'h0, 32'h41958dca, 32'h418ab2a7, 32'h0, 32'h4248ca8b, 32'h4299a422};
test_input[12600:12607] = '{32'hc10da79b, 32'h42ba2a17, 32'h42b6e71e, 32'h428f24c4, 32'h425c1696, 32'h40f2b283, 32'h42bacd2a, 32'h419e9f19};
test_output[12600:12607] = '{32'h0, 32'h42ba2a17, 32'h42b6e71e, 32'h428f24c4, 32'h425c1696, 32'h40f2b283, 32'h42bacd2a, 32'h419e9f19};
test_input[12608:12615] = '{32'h42b2f475, 32'h427413f2, 32'h418d195a, 32'hc2b8d165, 32'hc1218295, 32'hc214e695, 32'hc2b9179a, 32'h42c0ffce};
test_output[12608:12615] = '{32'h42b2f475, 32'h427413f2, 32'h418d195a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c0ffce};
test_input[12616:12623] = '{32'hbf01f0ff, 32'h42aedc7f, 32'h4240f0ba, 32'hc27fe553, 32'h41b0beed, 32'h42352638, 32'hc1f0d1f1, 32'h42a361e5};
test_output[12616:12623] = '{32'h0, 32'h42aedc7f, 32'h4240f0ba, 32'h0, 32'h41b0beed, 32'h42352638, 32'h0, 32'h42a361e5};
test_input[12624:12631] = '{32'h42c42a2a, 32'h4252b7c0, 32'h42c7e1ff, 32'hc1a7d1e8, 32'hc29a15cb, 32'hc2b9508c, 32'h421cee12, 32'h41ca4961};
test_output[12624:12631] = '{32'h42c42a2a, 32'h4252b7c0, 32'h42c7e1ff, 32'h0, 32'h0, 32'h0, 32'h421cee12, 32'h41ca4961};
test_input[12632:12639] = '{32'hc2aef0e4, 32'hc288caa6, 32'h4239d3f2, 32'hc208c61c, 32'h419762b1, 32'h413dedf8, 32'hc230f816, 32'h429815c4};
test_output[12632:12639] = '{32'h0, 32'h0, 32'h4239d3f2, 32'h0, 32'h419762b1, 32'h413dedf8, 32'h0, 32'h429815c4};
test_input[12640:12647] = '{32'hc23d9720, 32'h421588b2, 32'hc20d1f2b, 32'h42139732, 32'hc2121dbe, 32'hc038932f, 32'hc2701f85, 32'hc2c12f39};
test_output[12640:12647] = '{32'h0, 32'h421588b2, 32'h0, 32'h42139732, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[12648:12655] = '{32'hc2940af4, 32'hc2bc61af, 32'hc2bec896, 32'hc0a631e3, 32'h42776103, 32'hc23a1e3f, 32'h42a838f3, 32'hc18900d1};
test_output[12648:12655] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42776103, 32'h0, 32'h42a838f3, 32'h0};
test_input[12656:12663] = '{32'hc2814d2e, 32'h40c28991, 32'hc217dac8, 32'h42b015df, 32'hc21d73c3, 32'hc29f0d42, 32'h41b9f10e, 32'h423f445d};
test_output[12656:12663] = '{32'h0, 32'h40c28991, 32'h0, 32'h42b015df, 32'h0, 32'h0, 32'h41b9f10e, 32'h423f445d};
test_input[12664:12671] = '{32'hc251b253, 32'h42c5da9f, 32'h4280ff7f, 32'h4245717d, 32'hc27a8f9b, 32'hc290aa40, 32'h4281eb74, 32'hc0dbe255};
test_output[12664:12671] = '{32'h0, 32'h42c5da9f, 32'h4280ff7f, 32'h4245717d, 32'h0, 32'h0, 32'h4281eb74, 32'h0};
test_input[12672:12679] = '{32'hc22bf196, 32'hbe029585, 32'h429daa97, 32'h42a97e0f, 32'h42699000, 32'h42149d2a, 32'hc2520b0c, 32'hc1b5c8ac};
test_output[12672:12679] = '{32'h0, 32'h0, 32'h429daa97, 32'h42a97e0f, 32'h42699000, 32'h42149d2a, 32'h0, 32'h0};
test_input[12680:12687] = '{32'hc2a812aa, 32'h42aee734, 32'h4250cd9e, 32'h408d487c, 32'hc186c329, 32'hc271ba76, 32'h40ba0e8e, 32'hc17bcaec};
test_output[12680:12687] = '{32'h0, 32'h42aee734, 32'h4250cd9e, 32'h408d487c, 32'h0, 32'h0, 32'h40ba0e8e, 32'h0};
test_input[12688:12695] = '{32'hc1a44b9e, 32'hc216b3e0, 32'hc2c43f47, 32'hc24a4fd4, 32'hc28a7f4e, 32'h423318ac, 32'hc28b0efa, 32'hc1173703};
test_output[12688:12695] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423318ac, 32'h0, 32'h0};
test_input[12696:12703] = '{32'h429c1509, 32'h42916845, 32'h426d7213, 32'h42249048, 32'hc28c6fe1, 32'h428f2701, 32'h42afd48c, 32'hc0a3a319};
test_output[12696:12703] = '{32'h429c1509, 32'h42916845, 32'h426d7213, 32'h42249048, 32'h0, 32'h428f2701, 32'h42afd48c, 32'h0};
test_input[12704:12711] = '{32'h4213a293, 32'h41d9f7d7, 32'hc0b0fcff, 32'h41919437, 32'hc26af51a, 32'h425c35c8, 32'hc1e0e43e, 32'hc296ff6d};
test_output[12704:12711] = '{32'h4213a293, 32'h41d9f7d7, 32'h0, 32'h41919437, 32'h0, 32'h425c35c8, 32'h0, 32'h0};
test_input[12712:12719] = '{32'hc2a7c7d0, 32'h4286d4c2, 32'h4041bfd2, 32'h4286e398, 32'hc24d629e, 32'hc1b2e0e9, 32'h42535f6a, 32'h4119b975};
test_output[12712:12719] = '{32'h0, 32'h4286d4c2, 32'h4041bfd2, 32'h4286e398, 32'h0, 32'h0, 32'h42535f6a, 32'h4119b975};
test_input[12720:12727] = '{32'hc229e631, 32'h42ac89c6, 32'h42ada436, 32'h428c0d5e, 32'h426d60fc, 32'h4207be8c, 32'hc1648783, 32'h4286159d};
test_output[12720:12727] = '{32'h0, 32'h42ac89c6, 32'h42ada436, 32'h428c0d5e, 32'h426d60fc, 32'h4207be8c, 32'h0, 32'h4286159d};
test_input[12728:12735] = '{32'hc24135bc, 32'hc283cb11, 32'hc2a16c10, 32'h424ac794, 32'hc1c4457c, 32'hc22b48c1, 32'h423be80c, 32'h42a5d307};
test_output[12728:12735] = '{32'h0, 32'h0, 32'h0, 32'h424ac794, 32'h0, 32'h0, 32'h423be80c, 32'h42a5d307};
test_input[12736:12743] = '{32'h4241cedc, 32'hc23a79ad, 32'h42bbaf76, 32'hc2a9aa55, 32'h410c493d, 32'h42a33682, 32'h42a93746, 32'hc27b4e7b};
test_output[12736:12743] = '{32'h4241cedc, 32'h0, 32'h42bbaf76, 32'h0, 32'h410c493d, 32'h42a33682, 32'h42a93746, 32'h0};
test_input[12744:12751] = '{32'hc1f2814a, 32'h4292e440, 32'h42a4dd9e, 32'hc2219a63, 32'h3f05cd98, 32'h42bdf1aa, 32'h419a52ca, 32'h42bd4183};
test_output[12744:12751] = '{32'h0, 32'h4292e440, 32'h42a4dd9e, 32'h0, 32'h3f05cd98, 32'h42bdf1aa, 32'h419a52ca, 32'h42bd4183};
test_input[12752:12759] = '{32'h41cc63d6, 32'h41bf5aaa, 32'hc2935f12, 32'h428db3e2, 32'h424bffe1, 32'hc115458c, 32'h3ffedaac, 32'h41c36d94};
test_output[12752:12759] = '{32'h41cc63d6, 32'h41bf5aaa, 32'h0, 32'h428db3e2, 32'h424bffe1, 32'h0, 32'h3ffedaac, 32'h41c36d94};
test_input[12760:12767] = '{32'hc2aaca80, 32'hc18e0183, 32'h420274c3, 32'h41b0677a, 32'h4290716d, 32'hc28011f9, 32'h4269bfe1, 32'h40846cc2};
test_output[12760:12767] = '{32'h0, 32'h0, 32'h420274c3, 32'h41b0677a, 32'h4290716d, 32'h0, 32'h4269bfe1, 32'h40846cc2};
test_input[12768:12775] = '{32'hc155eb65, 32'h42976cf5, 32'h422c2c80, 32'hc2abbd36, 32'h42056b7d, 32'h42a13265, 32'hc284503b, 32'h4052e9e1};
test_output[12768:12775] = '{32'h0, 32'h42976cf5, 32'h422c2c80, 32'h0, 32'h42056b7d, 32'h42a13265, 32'h0, 32'h4052e9e1};
test_input[12776:12783] = '{32'h4295cafe, 32'hc29fe1fb, 32'hc2c600c2, 32'hbf862c84, 32'h41b2fa56, 32'h42a77c05, 32'hc1bc8cf3, 32'h427ec1e1};
test_output[12776:12783] = '{32'h4295cafe, 32'h0, 32'h0, 32'h0, 32'h41b2fa56, 32'h42a77c05, 32'h0, 32'h427ec1e1};
test_input[12784:12791] = '{32'hc1632815, 32'h428688e2, 32'h4230a545, 32'hc101f729, 32'h424b3c40, 32'hc197dd69, 32'hc21bbe2b, 32'hc0c569fd};
test_output[12784:12791] = '{32'h0, 32'h428688e2, 32'h4230a545, 32'h0, 32'h424b3c40, 32'h0, 32'h0, 32'h0};
test_input[12792:12799] = '{32'h42be1917, 32'h419f10cf, 32'hc265351e, 32'h420dd861, 32'hc2ad95f8, 32'hc29b2423, 32'h41b014a2, 32'hc2635da8};
test_output[12792:12799] = '{32'h42be1917, 32'h419f10cf, 32'h0, 32'h420dd861, 32'h0, 32'h0, 32'h41b014a2, 32'h0};
test_input[12800:12807] = '{32'hc2af6328, 32'h4287755f, 32'h41f26bac, 32'h41dc4321, 32'hc269ec22, 32'hc28a4224, 32'h42b49732, 32'h428c5b4d};
test_output[12800:12807] = '{32'h0, 32'h4287755f, 32'h41f26bac, 32'h41dc4321, 32'h0, 32'h0, 32'h42b49732, 32'h428c5b4d};
test_input[12808:12815] = '{32'h42ab9142, 32'h42461337, 32'h3fde3eed, 32'h429ab7d9, 32'hc2bbe4dc, 32'h41956e15, 32'h3ed26a69, 32'hc28aac27};
test_output[12808:12815] = '{32'h42ab9142, 32'h42461337, 32'h3fde3eed, 32'h429ab7d9, 32'h0, 32'h41956e15, 32'h3ed26a69, 32'h0};
test_input[12816:12823] = '{32'hc2aed2fc, 32'hc2479b5d, 32'hc2866008, 32'h41da4b4d, 32'hc15e03cb, 32'hc2a70562, 32'h42363af7, 32'hc2aeeb95};
test_output[12816:12823] = '{32'h0, 32'h0, 32'h0, 32'h41da4b4d, 32'h0, 32'h0, 32'h42363af7, 32'h0};
test_input[12824:12831] = '{32'h42ae8f04, 32'hc18a46ca, 32'hc1b1b6c8, 32'h4211041e, 32'hc1f5d2d6, 32'h41743813, 32'h40cbc4d8, 32'h42c3ce1a};
test_output[12824:12831] = '{32'h42ae8f04, 32'h0, 32'h0, 32'h4211041e, 32'h0, 32'h41743813, 32'h40cbc4d8, 32'h42c3ce1a};
test_input[12832:12839] = '{32'hc1247f3e, 32'h423004e0, 32'h4034ec61, 32'h42ba063c, 32'hc2c577d1, 32'h4277e43f, 32'h426ee5d0, 32'h41583bed};
test_output[12832:12839] = '{32'h0, 32'h423004e0, 32'h4034ec61, 32'h42ba063c, 32'h0, 32'h4277e43f, 32'h426ee5d0, 32'h41583bed};
test_input[12840:12847] = '{32'hc290d715, 32'hc17089ed, 32'h428f5c4d, 32'h41d0e8a9, 32'h42089ba7, 32'hc19b4911, 32'hc0e88045, 32'hc2294444};
test_output[12840:12847] = '{32'h0, 32'h0, 32'h428f5c4d, 32'h41d0e8a9, 32'h42089ba7, 32'h0, 32'h0, 32'h0};
test_input[12848:12855] = '{32'h404e5e5e, 32'hc1f36cb9, 32'hc0e225b1, 32'hc1e7f967, 32'h42a8a11f, 32'h427ed01f, 32'hc29ecf78, 32'h4131d67c};
test_output[12848:12855] = '{32'h404e5e5e, 32'h0, 32'h0, 32'h0, 32'h42a8a11f, 32'h427ed01f, 32'h0, 32'h4131d67c};
test_input[12856:12863] = '{32'hc2891f7b, 32'h42a0caa1, 32'h429f50ab, 32'hc0ec2d18, 32'hc1bdc40f, 32'hc2c592ee, 32'h42aa510f, 32'h42c5a8c8};
test_output[12856:12863] = '{32'h0, 32'h42a0caa1, 32'h429f50ab, 32'h0, 32'h0, 32'h0, 32'h42aa510f, 32'h42c5a8c8};
test_input[12864:12871] = '{32'hc1c4f80d, 32'h428d5519, 32'hc248a46e, 32'h420ce4db, 32'h4220dca2, 32'h3c83d042, 32'hc1e858b3, 32'hc0fe573a};
test_output[12864:12871] = '{32'h0, 32'h428d5519, 32'h0, 32'h420ce4db, 32'h4220dca2, 32'h3c83d042, 32'h0, 32'h0};
test_input[12872:12879] = '{32'h42567169, 32'h429dd673, 32'hc277887a, 32'hc2ab8e87, 32'hc2c7cd5d, 32'hc1f5bff5, 32'hc1ce63d5, 32'h426f9b8c};
test_output[12872:12879] = '{32'h42567169, 32'h429dd673, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426f9b8c};
test_input[12880:12887] = '{32'h42067a13, 32'h41cd903f, 32'h412d0da9, 32'hc2325a75, 32'h41c1ef93, 32'h42b4edb0, 32'h4259b062, 32'h427a73a1};
test_output[12880:12887] = '{32'h42067a13, 32'h41cd903f, 32'h412d0da9, 32'h0, 32'h41c1ef93, 32'h42b4edb0, 32'h4259b062, 32'h427a73a1};
test_input[12888:12895] = '{32'h42ac2863, 32'h42b9095b, 32'hc2981f9e, 32'h42a25b3b, 32'hc1626ec9, 32'h42a5436b, 32'h42b7c468, 32'hc26b2e88};
test_output[12888:12895] = '{32'h42ac2863, 32'h42b9095b, 32'h0, 32'h42a25b3b, 32'h0, 32'h42a5436b, 32'h42b7c468, 32'h0};
test_input[12896:12903] = '{32'hc0feff12, 32'hc2806c2e, 32'h421e50e5, 32'h4271cfdf, 32'h41a96bf6, 32'h428001aa, 32'h42bf4b37, 32'h42b0d99e};
test_output[12896:12903] = '{32'h0, 32'h0, 32'h421e50e5, 32'h4271cfdf, 32'h41a96bf6, 32'h428001aa, 32'h42bf4b37, 32'h42b0d99e};
test_input[12904:12911] = '{32'hc2345a4a, 32'h40fadd44, 32'hc28da005, 32'hc1c0b596, 32'h4285957a, 32'h422747a2, 32'h41ae8119, 32'h420accad};
test_output[12904:12911] = '{32'h0, 32'h40fadd44, 32'h0, 32'h0, 32'h4285957a, 32'h422747a2, 32'h41ae8119, 32'h420accad};
test_input[12912:12919] = '{32'h4296d90c, 32'h42ade3d9, 32'hc043323b, 32'h4241971d, 32'hc020ce64, 32'h41da0d32, 32'h42b75da6, 32'h42815e0b};
test_output[12912:12919] = '{32'h4296d90c, 32'h42ade3d9, 32'h0, 32'h4241971d, 32'h0, 32'h41da0d32, 32'h42b75da6, 32'h42815e0b};
test_input[12920:12927] = '{32'h429ff53c, 32'hc2317926, 32'h40be6c5d, 32'h429e790e, 32'h42477bac, 32'h42331e09, 32'hc292a4e5, 32'hc2976e3e};
test_output[12920:12927] = '{32'h429ff53c, 32'h0, 32'h40be6c5d, 32'h429e790e, 32'h42477bac, 32'h42331e09, 32'h0, 32'h0};
test_input[12928:12935] = '{32'hc25b1e90, 32'h4263ba4b, 32'hc2afa0a6, 32'hc11905c0, 32'h41a9ca50, 32'hc09d8a44, 32'h42039271, 32'hc24eb1b0};
test_output[12928:12935] = '{32'h0, 32'h4263ba4b, 32'h0, 32'h0, 32'h41a9ca50, 32'h0, 32'h42039271, 32'h0};
test_input[12936:12943] = '{32'h42adf22c, 32'h4213cdb0, 32'hc2a43f3b, 32'hc2c1ab6c, 32'h41b7b049, 32'h416e6030, 32'h40824a35, 32'hc26869cd};
test_output[12936:12943] = '{32'h42adf22c, 32'h4213cdb0, 32'h0, 32'h0, 32'h41b7b049, 32'h416e6030, 32'h40824a35, 32'h0};
test_input[12944:12951] = '{32'h42b84434, 32'hc295e665, 32'h429a6f78, 32'hc21350d1, 32'hc24608b4, 32'h4252f696, 32'h426f0cb9, 32'hc28cfe7f};
test_output[12944:12951] = '{32'h42b84434, 32'h0, 32'h429a6f78, 32'h0, 32'h0, 32'h4252f696, 32'h426f0cb9, 32'h0};
test_input[12952:12959] = '{32'hc218f0e2, 32'hc1c1b39a, 32'h428e82d6, 32'h42c703f2, 32'hc20043f4, 32'hc2babdfe, 32'h42471020, 32'hc290da40};
test_output[12952:12959] = '{32'h0, 32'h0, 32'h428e82d6, 32'h42c703f2, 32'h0, 32'h0, 32'h42471020, 32'h0};
test_input[12960:12967] = '{32'h420575fb, 32'h429bd57a, 32'hc282e8bb, 32'hc26f97e0, 32'h42c413a7, 32'hc268dc13, 32'h41b773f6, 32'h41fd2fa9};
test_output[12960:12967] = '{32'h420575fb, 32'h429bd57a, 32'h0, 32'h0, 32'h42c413a7, 32'h0, 32'h41b773f6, 32'h41fd2fa9};
test_input[12968:12975] = '{32'hc2bd9c99, 32'hc1c9fbdd, 32'h40878580, 32'h42bf723f, 32'h41389442, 32'hc001c2c8, 32'hc2649d9b, 32'h41ecffef};
test_output[12968:12975] = '{32'h0, 32'h0, 32'h40878580, 32'h42bf723f, 32'h41389442, 32'h0, 32'h0, 32'h41ecffef};
test_input[12976:12983] = '{32'h424b6368, 32'hc28eb44f, 32'h40d26f60, 32'h420f635a, 32'h423dec82, 32'h4235f3ad, 32'h42a7b9ce, 32'h424d2d21};
test_output[12976:12983] = '{32'h424b6368, 32'h0, 32'h40d26f60, 32'h420f635a, 32'h423dec82, 32'h4235f3ad, 32'h42a7b9ce, 32'h424d2d21};
test_input[12984:12991] = '{32'h42492532, 32'hc292f41c, 32'h42722bde, 32'hc1b1fdc7, 32'hc2840655, 32'hc20e9646, 32'hc14986eb, 32'h428c5e51};
test_output[12984:12991] = '{32'h42492532, 32'h0, 32'h42722bde, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428c5e51};
test_input[12992:12999] = '{32'h428da9ac, 32'h424e1b43, 32'h413ffaf7, 32'h41061084, 32'h427c3591, 32'h414976a2, 32'h42ab5799, 32'hc151bfe8};
test_output[12992:12999] = '{32'h428da9ac, 32'h424e1b43, 32'h413ffaf7, 32'h41061084, 32'h427c3591, 32'h414976a2, 32'h42ab5799, 32'h0};
test_input[13000:13007] = '{32'h41f32af7, 32'h42740617, 32'hc236d685, 32'hc2345415, 32'hc21ed6ff, 32'h42acd2ef, 32'h414c65ab, 32'h42b50b73};
test_output[13000:13007] = '{32'h41f32af7, 32'h42740617, 32'h0, 32'h0, 32'h0, 32'h42acd2ef, 32'h414c65ab, 32'h42b50b73};
test_input[13008:13015] = '{32'hc203fef0, 32'h40bf2f83, 32'hc220a5c6, 32'hc1d0d797, 32'hc2540c6e, 32'hc2626f66, 32'h410c441a, 32'hc1b2bb8c};
test_output[13008:13015] = '{32'h0, 32'h40bf2f83, 32'h0, 32'h0, 32'h0, 32'h0, 32'h410c441a, 32'h0};
test_input[13016:13023] = '{32'h418fc280, 32'h426671d9, 32'hc1a40bc5, 32'h41fb27a2, 32'hc1820081, 32'hc22f8739, 32'hc1fe4942, 32'hc28bc256};
test_output[13016:13023] = '{32'h418fc280, 32'h426671d9, 32'h0, 32'h41fb27a2, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13024:13031] = '{32'h41666886, 32'h41d98387, 32'h42972471, 32'h429cbc09, 32'hc2c04a46, 32'h42999372, 32'h42c113f4, 32'h4290b8b6};
test_output[13024:13031] = '{32'h41666886, 32'h41d98387, 32'h42972471, 32'h429cbc09, 32'h0, 32'h42999372, 32'h42c113f4, 32'h4290b8b6};
test_input[13032:13039] = '{32'h40ea74cb, 32'h41f08ef1, 32'h423171cb, 32'h418b1d83, 32'hc2c42f8e, 32'h41bf7967, 32'hc1b95caf, 32'h41569291};
test_output[13032:13039] = '{32'h40ea74cb, 32'h41f08ef1, 32'h423171cb, 32'h418b1d83, 32'h0, 32'h41bf7967, 32'h0, 32'h41569291};
test_input[13040:13047] = '{32'h4286ea9d, 32'hc2659b86, 32'hc0af2c0d, 32'h42b5d88c, 32'h42b38a07, 32'hc2c1133e, 32'h429cc744, 32'h4187287b};
test_output[13040:13047] = '{32'h4286ea9d, 32'h0, 32'h0, 32'h42b5d88c, 32'h42b38a07, 32'h0, 32'h429cc744, 32'h4187287b};
test_input[13048:13055] = '{32'h429bd0a1, 32'h41579174, 32'h429c1f51, 32'h41c98fb1, 32'hc23986f1, 32'hc2accf08, 32'hc2b9446a, 32'h402767c2};
test_output[13048:13055] = '{32'h429bd0a1, 32'h41579174, 32'h429c1f51, 32'h41c98fb1, 32'h0, 32'h0, 32'h0, 32'h402767c2};
test_input[13056:13063] = '{32'hc28b806c, 32'hc2b25e55, 32'hc108cbcb, 32'h412d79af, 32'h42556c4a, 32'h4289349e, 32'h428354da, 32'h417a11e6};
test_output[13056:13063] = '{32'h0, 32'h0, 32'h0, 32'h412d79af, 32'h42556c4a, 32'h4289349e, 32'h428354da, 32'h417a11e6};
test_input[13064:13071] = '{32'h421dad05, 32'h4252b3be, 32'h424a4093, 32'hc1b88be9, 32'h4280bf22, 32'h42c58434, 32'hc20d0fa6, 32'h425d2b18};
test_output[13064:13071] = '{32'h421dad05, 32'h4252b3be, 32'h424a4093, 32'h0, 32'h4280bf22, 32'h42c58434, 32'h0, 32'h425d2b18};
test_input[13072:13079] = '{32'h4150788d, 32'hc0f2a40b, 32'hc2958446, 32'hc0155b5c, 32'hc24cb9bb, 32'hc17a4cdf, 32'h419dc907, 32'h412f0971};
test_output[13072:13079] = '{32'h4150788d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h419dc907, 32'h412f0971};
test_input[13080:13087] = '{32'hc28af80d, 32'hc2994ed6, 32'h42be29fe, 32'hc194d998, 32'hc2892e5b, 32'h429c293d, 32'hc21e1f51, 32'hc1f9bc6f};
test_output[13080:13087] = '{32'h0, 32'h0, 32'h42be29fe, 32'h0, 32'h0, 32'h429c293d, 32'h0, 32'h0};
test_input[13088:13095] = '{32'h4271d8e4, 32'hc2b8a725, 32'hc297f75c, 32'h42c3eb85, 32'hc0a9b576, 32'hc233e1e7, 32'hc27a2a92, 32'hc2a1e973};
test_output[13088:13095] = '{32'h4271d8e4, 32'h0, 32'h0, 32'h42c3eb85, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13096:13103] = '{32'h4170edd6, 32'h42bd3d7f, 32'hc118d79c, 32'hc29a520d, 32'h423ec318, 32'hc2454b7f, 32'hc288bd54, 32'hc2588360};
test_output[13096:13103] = '{32'h4170edd6, 32'h42bd3d7f, 32'h0, 32'h0, 32'h423ec318, 32'h0, 32'h0, 32'h0};
test_input[13104:13111] = '{32'hc28258bf, 32'h4156f7ad, 32'h422d70fb, 32'h422a64bb, 32'h41d3a052, 32'h42b32fbf, 32'h412dae4b, 32'h42aeea5f};
test_output[13104:13111] = '{32'h0, 32'h4156f7ad, 32'h422d70fb, 32'h422a64bb, 32'h41d3a052, 32'h42b32fbf, 32'h412dae4b, 32'h42aeea5f};
test_input[13112:13119] = '{32'h409852d2, 32'hc28a0326, 32'hc2720282, 32'h42c7129f, 32'hc1e6c8f0, 32'hc2c5a0ff, 32'h42c11fbf, 32'hc29805f6};
test_output[13112:13119] = '{32'h409852d2, 32'h0, 32'h0, 32'h42c7129f, 32'h0, 32'h0, 32'h42c11fbf, 32'h0};
test_input[13120:13127] = '{32'h42449239, 32'hc10773ff, 32'h4293c25e, 32'h42ba42fc, 32'h4207feb0, 32'hc24c9b45, 32'hc246fa62, 32'h41c954ce};
test_output[13120:13127] = '{32'h42449239, 32'h0, 32'h4293c25e, 32'h42ba42fc, 32'h4207feb0, 32'h0, 32'h0, 32'h41c954ce};
test_input[13128:13135] = '{32'hc2c24596, 32'h42307afc, 32'hc2b25762, 32'h42a6855f, 32'hc16fda19, 32'hc2ad114e, 32'h422d4b63, 32'hc27249cf};
test_output[13128:13135] = '{32'h0, 32'h42307afc, 32'h0, 32'h42a6855f, 32'h0, 32'h0, 32'h422d4b63, 32'h0};
test_input[13136:13143] = '{32'hc29537f1, 32'h42878220, 32'h415024c2, 32'hc2a763b3, 32'h41ed97e4, 32'h41c59337, 32'h427433ac, 32'hc282226d};
test_output[13136:13143] = '{32'h0, 32'h42878220, 32'h415024c2, 32'h0, 32'h41ed97e4, 32'h41c59337, 32'h427433ac, 32'h0};
test_input[13144:13151] = '{32'hc269d649, 32'h4210883f, 32'hc2823375, 32'h422b97f1, 32'hc209e5d3, 32'hc2172b8f, 32'hc1545864, 32'h42119371};
test_output[13144:13151] = '{32'h0, 32'h4210883f, 32'h0, 32'h422b97f1, 32'h0, 32'h0, 32'h0, 32'h42119371};
test_input[13152:13159] = '{32'h3fc4d3c1, 32'h42b12fe6, 32'h42b8531c, 32'hc2c36d74, 32'hc297c88d, 32'hc2abb5a7, 32'h4283629f, 32'h429d63d4};
test_output[13152:13159] = '{32'h3fc4d3c1, 32'h42b12fe6, 32'h42b8531c, 32'h0, 32'h0, 32'h0, 32'h4283629f, 32'h429d63d4};
test_input[13160:13167] = '{32'h409e8191, 32'h426020f3, 32'h42037a17, 32'hc25e143e, 32'h42b84d33, 32'hc288c5cb, 32'hc2368575, 32'hbdad46d4};
test_output[13160:13167] = '{32'h409e8191, 32'h426020f3, 32'h42037a17, 32'h0, 32'h42b84d33, 32'h0, 32'h0, 32'h0};
test_input[13168:13175] = '{32'h427a7a60, 32'h42a73409, 32'h41f8ad1d, 32'h42b0355c, 32'hc201dec4, 32'h422a8dfc, 32'h4200dfef, 32'hc0c75b52};
test_output[13168:13175] = '{32'h427a7a60, 32'h42a73409, 32'h41f8ad1d, 32'h42b0355c, 32'h0, 32'h422a8dfc, 32'h4200dfef, 32'h0};
test_input[13176:13183] = '{32'hc19a4d2a, 32'hc28a8632, 32'h40ad641e, 32'hc28e80d9, 32'h4186d242, 32'hc2712317, 32'h423314b9, 32'hc1ad8db1};
test_output[13176:13183] = '{32'h0, 32'h0, 32'h40ad641e, 32'h0, 32'h4186d242, 32'h0, 32'h423314b9, 32'h0};
test_input[13184:13191] = '{32'hc2c43d5e, 32'hc0e51018, 32'h41db2519, 32'hc22332a0, 32'hc2677ec1, 32'hc219044b, 32'h41f342f7, 32'h42ac8e97};
test_output[13184:13191] = '{32'h0, 32'h0, 32'h41db2519, 32'h0, 32'h0, 32'h0, 32'h41f342f7, 32'h42ac8e97};
test_input[13192:13199] = '{32'h41a21c51, 32'hc254186a, 32'h42bf1d55, 32'hc15dc29a, 32'hc0dd8d2f, 32'h42bc8687, 32'hc163298a, 32'h40df958b};
test_output[13192:13199] = '{32'h41a21c51, 32'h0, 32'h42bf1d55, 32'h0, 32'h0, 32'h42bc8687, 32'h0, 32'h40df958b};
test_input[13200:13207] = '{32'hc2709bd7, 32'hc24730f6, 32'hc26679e1, 32'h421aa917, 32'h42431347, 32'hc22af128, 32'hc18d1b26, 32'hc239846b};
test_output[13200:13207] = '{32'h0, 32'h0, 32'h0, 32'h421aa917, 32'h42431347, 32'h0, 32'h0, 32'h0};
test_input[13208:13215] = '{32'h429ae4be, 32'hc19f1827, 32'hc22b8576, 32'hc2624b84, 32'hc2aede73, 32'hc130fa69, 32'h420cd06b, 32'h427e1e22};
test_output[13208:13215] = '{32'h429ae4be, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420cd06b, 32'h427e1e22};
test_input[13216:13223] = '{32'h4206bca0, 32'hc279f085, 32'hc26b0db1, 32'h408f4c07, 32'hbf64b000, 32'hc28adbfc, 32'hc1c38a11, 32'hc0f236f3};
test_output[13216:13223] = '{32'h4206bca0, 32'h0, 32'h0, 32'h408f4c07, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13224:13231] = '{32'hc1bfd97a, 32'h42205409, 32'h42464494, 32'h41be50af, 32'h42586a57, 32'h429c1f24, 32'h42939a05, 32'h42aacea8};
test_output[13224:13231] = '{32'h0, 32'h42205409, 32'h42464494, 32'h41be50af, 32'h42586a57, 32'h429c1f24, 32'h42939a05, 32'h42aacea8};
test_input[13232:13239] = '{32'hc2956003, 32'hc2a51326, 32'h424dbd97, 32'h42a0ee7b, 32'hc2936bc6, 32'h426db818, 32'hc29389b0, 32'hc0dcb8ae};
test_output[13232:13239] = '{32'h0, 32'h0, 32'h424dbd97, 32'h42a0ee7b, 32'h0, 32'h426db818, 32'h0, 32'h0};
test_input[13240:13247] = '{32'h42591a50, 32'hc20e3042, 32'hc287e317, 32'hc2bc01d9, 32'hc217c682, 32'hc2999549, 32'h42077aa3, 32'hc238eb37};
test_output[13240:13247] = '{32'h42591a50, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42077aa3, 32'h0};
test_input[13248:13255] = '{32'hc2bee574, 32'h4290e4eb, 32'hc2b5fb67, 32'h428224b8, 32'hbfb4e666, 32'h4189112e, 32'hc233b4e0, 32'h424abca7};
test_output[13248:13255] = '{32'h0, 32'h4290e4eb, 32'h0, 32'h428224b8, 32'h0, 32'h4189112e, 32'h0, 32'h424abca7};
test_input[13256:13263] = '{32'hc29a43b6, 32'h42163d7e, 32'hbe72dfe6, 32'hc2a14185, 32'h412c2356, 32'hc29475d9, 32'hc21366a7, 32'h42213eda};
test_output[13256:13263] = '{32'h0, 32'h42163d7e, 32'h0, 32'h0, 32'h412c2356, 32'h0, 32'h0, 32'h42213eda};
test_input[13264:13271] = '{32'h424fd134, 32'h42b9e5b9, 32'h41bd64c6, 32'h42a08aa3, 32'h42a17a6a, 32'h42884850, 32'h3fa78588, 32'hc2829643};
test_output[13264:13271] = '{32'h424fd134, 32'h42b9e5b9, 32'h41bd64c6, 32'h42a08aa3, 32'h42a17a6a, 32'h42884850, 32'h3fa78588, 32'h0};
test_input[13272:13279] = '{32'h41a79fa3, 32'hc2806d85, 32'hc1d37cbe, 32'hc28f6ca7, 32'hc132a46b, 32'h42968b0c, 32'hc1bf0a07, 32'h42b596b2};
test_output[13272:13279] = '{32'h41a79fa3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42968b0c, 32'h0, 32'h42b596b2};
test_input[13280:13287] = '{32'h42260aae, 32'hc0f792ff, 32'h4157d3b9, 32'hc253a237, 32'h425e732b, 32'h42af9ec5, 32'hc2a911df, 32'h4288a976};
test_output[13280:13287] = '{32'h42260aae, 32'h0, 32'h4157d3b9, 32'h0, 32'h425e732b, 32'h42af9ec5, 32'h0, 32'h4288a976};
test_input[13288:13295] = '{32'hc28da513, 32'hc2707e02, 32'hc282099a, 32'h41bb20e7, 32'hc2ada8f6, 32'hc27826cf, 32'h42ad2f9c, 32'h426d1543};
test_output[13288:13295] = '{32'h0, 32'h0, 32'h0, 32'h41bb20e7, 32'h0, 32'h0, 32'h42ad2f9c, 32'h426d1543};
test_input[13296:13303] = '{32'hc207e398, 32'h41806c2b, 32'h4289c887, 32'hc2101284, 32'hc2a2c8e6, 32'h424dce26, 32'h40d12d82, 32'h42c37cc2};
test_output[13296:13303] = '{32'h0, 32'h41806c2b, 32'h4289c887, 32'h0, 32'h0, 32'h424dce26, 32'h40d12d82, 32'h42c37cc2};
test_input[13304:13311] = '{32'hc1b4bf1e, 32'hc067a334, 32'h42165a50, 32'h42991d1c, 32'hc27b4494, 32'h41b795e2, 32'h42af7444, 32'hc1fedec4};
test_output[13304:13311] = '{32'h0, 32'h0, 32'h42165a50, 32'h42991d1c, 32'h0, 32'h41b795e2, 32'h42af7444, 32'h0};
test_input[13312:13319] = '{32'hc1f1e038, 32'h4180d0af, 32'h4159bdb2, 32'hc279f7fb, 32'h42b15072, 32'h42761dd2, 32'hc10b0e02, 32'hc2bb1a3f};
test_output[13312:13319] = '{32'h0, 32'h4180d0af, 32'h4159bdb2, 32'h0, 32'h42b15072, 32'h42761dd2, 32'h0, 32'h0};
test_input[13320:13327] = '{32'h420662b9, 32'hc27dae05, 32'h42a0d66f, 32'h42a76ee7, 32'h41a9375c, 32'h42c38e60, 32'hc1babce1, 32'hc2747152};
test_output[13320:13327] = '{32'h420662b9, 32'h0, 32'h42a0d66f, 32'h42a76ee7, 32'h41a9375c, 32'h42c38e60, 32'h0, 32'h0};
test_input[13328:13335] = '{32'hc2586ffb, 32'hc0086ded, 32'h42bff690, 32'hc2b3408b, 32'hc2be7474, 32'hc28bc8f5, 32'hc075de11, 32'hc23622b4};
test_output[13328:13335] = '{32'h0, 32'h0, 32'h42bff690, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13336:13343] = '{32'hc228d3b3, 32'h42beb3a6, 32'hc2b9d29a, 32'h421679a1, 32'hc2c6aa33, 32'h429da5e2, 32'h422eef16, 32'hc223099e};
test_output[13336:13343] = '{32'h0, 32'h42beb3a6, 32'h0, 32'h421679a1, 32'h0, 32'h429da5e2, 32'h422eef16, 32'h0};
test_input[13344:13351] = '{32'h425281a0, 32'hc2a24ba0, 32'hc288b855, 32'hc2b5c411, 32'h42b02183, 32'hc2820272, 32'h42c67517, 32'hc28d1ae7};
test_output[13344:13351] = '{32'h425281a0, 32'h0, 32'h0, 32'h0, 32'h42b02183, 32'h0, 32'h42c67517, 32'h0};
test_input[13352:13359] = '{32'hc24c5608, 32'h4260d8ee, 32'h419d3e28, 32'hc217e79d, 32'h4189e328, 32'hc198a0e9, 32'hc2442817, 32'hc2c187c8};
test_output[13352:13359] = '{32'h0, 32'h4260d8ee, 32'h419d3e28, 32'h0, 32'h4189e328, 32'h0, 32'h0, 32'h0};
test_input[13360:13367] = '{32'h4295e262, 32'hc2b0fdd9, 32'h41e4b044, 32'hc251d5eb, 32'hc2b7d7d5, 32'h4130eef7, 32'h42a7b760, 32'h4299ba7f};
test_output[13360:13367] = '{32'h4295e262, 32'h0, 32'h41e4b044, 32'h0, 32'h0, 32'h4130eef7, 32'h42a7b760, 32'h4299ba7f};
test_input[13368:13375] = '{32'hc249a3b6, 32'h41110791, 32'h42967207, 32'h42a55dd5, 32'hc21bee58, 32'h4251a53b, 32'hc2c2f6f8, 32'hc29c1b41};
test_output[13368:13375] = '{32'h0, 32'h41110791, 32'h42967207, 32'h42a55dd5, 32'h0, 32'h4251a53b, 32'h0, 32'h0};
test_input[13376:13383] = '{32'hc13d951e, 32'hc2b80470, 32'h422c0457, 32'hc287236a, 32'h429e30d2, 32'hc252849c, 32'h425f1c12, 32'hc20f40de};
test_output[13376:13383] = '{32'h0, 32'h0, 32'h422c0457, 32'h0, 32'h429e30d2, 32'h0, 32'h425f1c12, 32'h0};
test_input[13384:13391] = '{32'hc29e39b7, 32'hc2a623c3, 32'h41c96a7f, 32'hc2b858e5, 32'hbf49c0f9, 32'h422485be, 32'hc29a69a0, 32'hc1af8513};
test_output[13384:13391] = '{32'h0, 32'h0, 32'h41c96a7f, 32'h0, 32'h0, 32'h422485be, 32'h0, 32'h0};
test_input[13392:13399] = '{32'hc1426e30, 32'h428f7fdc, 32'hc2a9f0ad, 32'hc1ce279a, 32'hc159dbfe, 32'hc2be47ad, 32'h42966f20, 32'hc16d07e5};
test_output[13392:13399] = '{32'h0, 32'h428f7fdc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42966f20, 32'h0};
test_input[13400:13407] = '{32'h4101c278, 32'hc1bcfcbe, 32'hc2995ea9, 32'hc1c5a401, 32'h42af017e, 32'h42a54df4, 32'hc02b7141, 32'hc1e78160};
test_output[13400:13407] = '{32'h4101c278, 32'h0, 32'h0, 32'h0, 32'h42af017e, 32'h42a54df4, 32'h0, 32'h0};
test_input[13408:13415] = '{32'hc1edf016, 32'h42b98cc6, 32'h420e2921, 32'hc11c0d9e, 32'hc1c9cfff, 32'hc2578a7d, 32'hc2603fbd, 32'hc2ac4891};
test_output[13408:13415] = '{32'h0, 32'h42b98cc6, 32'h420e2921, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13416:13423] = '{32'hc250ce91, 32'hc03442d1, 32'hc1258874, 32'hc29e1243, 32'h422e0e38, 32'hc2c59aaa, 32'hc276cf45, 32'h41e7581f};
test_output[13416:13423] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h422e0e38, 32'h0, 32'h0, 32'h41e7581f};
test_input[13424:13431] = '{32'hc24aa2ff, 32'hc2aead2e, 32'h40e14e2b, 32'h421cee10, 32'h42826a5c, 32'hc20c8f96, 32'h42c35bdb, 32'h42792cc9};
test_output[13424:13431] = '{32'h0, 32'h0, 32'h40e14e2b, 32'h421cee10, 32'h42826a5c, 32'h0, 32'h42c35bdb, 32'h42792cc9};
test_input[13432:13439] = '{32'h404e9aaf, 32'hc29ae0f0, 32'h41e34d26, 32'hc2c2a4fd, 32'hc2bc65a6, 32'hc29edf17, 32'hc2c5364a, 32'hc1ed39aa};
test_output[13432:13439] = '{32'h404e9aaf, 32'h0, 32'h41e34d26, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13440:13447] = '{32'h428e4334, 32'hc0a0bf94, 32'h4192ff75, 32'hc28fca6c, 32'h42a1284e, 32'hc27abca4, 32'hc2862b09, 32'h42c4eb84};
test_output[13440:13447] = '{32'h428e4334, 32'h0, 32'h4192ff75, 32'h0, 32'h42a1284e, 32'h0, 32'h0, 32'h42c4eb84};
test_input[13448:13455] = '{32'h4251f68f, 32'hc1869505, 32'h42c6209f, 32'h4157e40f, 32'hc1520e47, 32'h415387ed, 32'h425465db, 32'hc2630414};
test_output[13448:13455] = '{32'h4251f68f, 32'h0, 32'h42c6209f, 32'h4157e40f, 32'h0, 32'h415387ed, 32'h425465db, 32'h0};
test_input[13456:13463] = '{32'hc2b6fe04, 32'hc1f97a32, 32'h41adbd45, 32'hc204bb5b, 32'h4001bdd2, 32'h42757ee1, 32'hc1ea19b9, 32'h42a21b8c};
test_output[13456:13463] = '{32'h0, 32'h0, 32'h41adbd45, 32'h0, 32'h4001bdd2, 32'h42757ee1, 32'h0, 32'h42a21b8c};
test_input[13464:13471] = '{32'hc2864f5b, 32'hc2b304b4, 32'h41d42928, 32'h42a06afe, 32'h42606139, 32'h41e5dcb2, 32'hc21f7292, 32'hc2c07a3b};
test_output[13464:13471] = '{32'h0, 32'h0, 32'h41d42928, 32'h42a06afe, 32'h42606139, 32'h41e5dcb2, 32'h0, 32'h0};
test_input[13472:13479] = '{32'h42913ed2, 32'hc2a23547, 32'hc298b058, 32'h41c9d46a, 32'hc2bf1d97, 32'h4294e303, 32'h418081aa, 32'h41cc9e88};
test_output[13472:13479] = '{32'h42913ed2, 32'h0, 32'h0, 32'h41c9d46a, 32'h0, 32'h4294e303, 32'h418081aa, 32'h41cc9e88};
test_input[13480:13487] = '{32'h4255a2a7, 32'hc218c631, 32'h3ec0bdc1, 32'hc23000ab, 32'hc2560112, 32'hc1bafa2b, 32'h420ae811, 32'hc22ec79f};
test_output[13480:13487] = '{32'h4255a2a7, 32'h0, 32'h3ec0bdc1, 32'h0, 32'h0, 32'h0, 32'h420ae811, 32'h0};
test_input[13488:13495] = '{32'h426d947e, 32'hc28a07fd, 32'h42b573e7, 32'hc25ab2e8, 32'hc183d58d, 32'hc2aa5661, 32'hc1315e9b, 32'h42a4197d};
test_output[13488:13495] = '{32'h426d947e, 32'h0, 32'h42b573e7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a4197d};
test_input[13496:13503] = '{32'hc0d98374, 32'hc2ae4d46, 32'h42b639b9, 32'h41c4b815, 32'hc2108aa3, 32'hc2ad70ea, 32'h42c039cc, 32'hc2b4e050};
test_output[13496:13503] = '{32'h0, 32'h0, 32'h42b639b9, 32'h41c4b815, 32'h0, 32'h0, 32'h42c039cc, 32'h0};
test_input[13504:13511] = '{32'h42b03647, 32'h42b8d8e8, 32'hc27d7ff7, 32'hc202d06d, 32'hc25c62a5, 32'h426b1838, 32'h422ce3ad, 32'hc28ac0d1};
test_output[13504:13511] = '{32'h42b03647, 32'h42b8d8e8, 32'h0, 32'h0, 32'h0, 32'h426b1838, 32'h422ce3ad, 32'h0};
test_input[13512:13519] = '{32'hc0e4f720, 32'hc1c2faf8, 32'h41918335, 32'hc2bbcc79, 32'hc1558eb2, 32'hc2b16107, 32'h42bb14d4, 32'h4226316b};
test_output[13512:13519] = '{32'h0, 32'h0, 32'h41918335, 32'h0, 32'h0, 32'h0, 32'h42bb14d4, 32'h4226316b};
test_input[13520:13527] = '{32'h425c581f, 32'hc211e4a6, 32'hc2254a20, 32'hc203f2af, 32'hc277eda3, 32'hc20726a5, 32'hc28a227f, 32'h41e35597};
test_output[13520:13527] = '{32'h425c581f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41e35597};
test_input[13528:13535] = '{32'h42c3baea, 32'h423acb34, 32'h41492067, 32'hc0ee5805, 32'h3f22b7a7, 32'hc2887eb8, 32'h42434b4c, 32'h41ee2bab};
test_output[13528:13535] = '{32'h42c3baea, 32'h423acb34, 32'h41492067, 32'h0, 32'h3f22b7a7, 32'h0, 32'h42434b4c, 32'h41ee2bab};
test_input[13536:13543] = '{32'hc1a2bb37, 32'hc12db5ee, 32'h42746f3e, 32'h428dfd4f, 32'h40ea5550, 32'h408b734e, 32'h4244b9ee, 32'hc2a8871c};
test_output[13536:13543] = '{32'h0, 32'h0, 32'h42746f3e, 32'h428dfd4f, 32'h40ea5550, 32'h408b734e, 32'h4244b9ee, 32'h0};
test_input[13544:13551] = '{32'h42bf6d3f, 32'hc28e7c29, 32'hc2847f62, 32'h42236579, 32'h428495a6, 32'hc204d1c4, 32'h421aa32a, 32'hc18ea1db};
test_output[13544:13551] = '{32'h42bf6d3f, 32'h0, 32'h0, 32'h42236579, 32'h428495a6, 32'h0, 32'h421aa32a, 32'h0};
test_input[13552:13559] = '{32'h427e3ffe, 32'h40825f9d, 32'hc2496e22, 32'h41cfd0d3, 32'hc1ac7751, 32'h42bd781b, 32'h427cca26, 32'hc29c75ba};
test_output[13552:13559] = '{32'h427e3ffe, 32'h40825f9d, 32'h0, 32'h41cfd0d3, 32'h0, 32'h42bd781b, 32'h427cca26, 32'h0};
test_input[13560:13567] = '{32'hc272c482, 32'hc280faba, 32'h4297db14, 32'hc2063a5f, 32'h4227e8e1, 32'h415f9b7b, 32'hc1faeac0, 32'hc2b868fb};
test_output[13560:13567] = '{32'h0, 32'h0, 32'h4297db14, 32'h0, 32'h4227e8e1, 32'h415f9b7b, 32'h0, 32'h0};
test_input[13568:13575] = '{32'h42374339, 32'hc2c40260, 32'hc2a81928, 32'h3f152aaa, 32'h42c09c2a, 32'h41aed5d6, 32'hc1f022f2, 32'h42a1d68d};
test_output[13568:13575] = '{32'h42374339, 32'h0, 32'h0, 32'h3f152aaa, 32'h42c09c2a, 32'h41aed5d6, 32'h0, 32'h42a1d68d};
test_input[13576:13583] = '{32'hc25c01d2, 32'h42c06ddc, 32'h41fc1b49, 32'hc29c8254, 32'h41ba3a91, 32'h3f541166, 32'hc2bbacad, 32'hc2a93543};
test_output[13576:13583] = '{32'h0, 32'h42c06ddc, 32'h41fc1b49, 32'h0, 32'h41ba3a91, 32'h3f541166, 32'h0, 32'h0};
test_input[13584:13591] = '{32'hc29e4362, 32'h41173f1a, 32'h4205b0d7, 32'hc25b25e1, 32'hc2147a4b, 32'hc1cef5f4, 32'hc1db499d, 32'h41b6a497};
test_output[13584:13591] = '{32'h0, 32'h41173f1a, 32'h4205b0d7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b6a497};
test_input[13592:13599] = '{32'h409dda12, 32'hc2a91422, 32'hc24e8523, 32'hc00afcdf, 32'h428f6190, 32'h4295b1a9, 32'h40aa5f36, 32'hc2046966};
test_output[13592:13599] = '{32'h409dda12, 32'h0, 32'h0, 32'h0, 32'h428f6190, 32'h4295b1a9, 32'h40aa5f36, 32'h0};
test_input[13600:13607] = '{32'hc1bb223f, 32'hc14a7fae, 32'h41bb87ad, 32'h405be4f2, 32'hc29c96ff, 32'h40d5edd9, 32'hc2a296b0, 32'hc27fc735};
test_output[13600:13607] = '{32'h0, 32'h0, 32'h41bb87ad, 32'h405be4f2, 32'h0, 32'h40d5edd9, 32'h0, 32'h0};
test_input[13608:13615] = '{32'hc1a2fe38, 32'h423c845b, 32'h4283c344, 32'h4292b7bb, 32'h42c1833a, 32'hc2153084, 32'h42009586, 32'hc266b7ec};
test_output[13608:13615] = '{32'h0, 32'h423c845b, 32'h4283c344, 32'h4292b7bb, 32'h42c1833a, 32'h0, 32'h42009586, 32'h0};
test_input[13616:13623] = '{32'h42955f64, 32'h4297bc9d, 32'h42684f8c, 32'h40ebcb9e, 32'hc245e551, 32'hc1e382ce, 32'hc2a12b13, 32'h42a9c117};
test_output[13616:13623] = '{32'h42955f64, 32'h4297bc9d, 32'h42684f8c, 32'h40ebcb9e, 32'h0, 32'h0, 32'h0, 32'h42a9c117};
test_input[13624:13631] = '{32'h4220cf26, 32'h3d472214, 32'hc286b762, 32'hc19100b1, 32'hc23f0eed, 32'hc2ae337d, 32'h414c5325, 32'h42a0f793};
test_output[13624:13631] = '{32'h4220cf26, 32'h3d472214, 32'h0, 32'h0, 32'h0, 32'h0, 32'h414c5325, 32'h42a0f793};
test_input[13632:13639] = '{32'h41181de6, 32'hc219f5c2, 32'hc2c46b42, 32'hc1dc935b, 32'h41c42a1d, 32'h42892e34, 32'hc29ad444, 32'h42a1fcfc};
test_output[13632:13639] = '{32'h41181de6, 32'h0, 32'h0, 32'h0, 32'h41c42a1d, 32'h42892e34, 32'h0, 32'h42a1fcfc};
test_input[13640:13647] = '{32'h42c2c186, 32'h428244de, 32'hc2082a72, 32'h429c4254, 32'hc272b686, 32'hc182a0ff, 32'h428d730b, 32'h4286ee98};
test_output[13640:13647] = '{32'h42c2c186, 32'h428244de, 32'h0, 32'h429c4254, 32'h0, 32'h0, 32'h428d730b, 32'h4286ee98};
test_input[13648:13655] = '{32'hc11fb61c, 32'hc2079c49, 32'h42506c55, 32'hc2898a11, 32'h4268c151, 32'h42433bda, 32'h42b6cacb, 32'hc2bed436};
test_output[13648:13655] = '{32'h0, 32'h0, 32'h42506c55, 32'h0, 32'h4268c151, 32'h42433bda, 32'h42b6cacb, 32'h0};
test_input[13656:13663] = '{32'hc0b519a7, 32'h41bd8d93, 32'hc2a62522, 32'h429666ba, 32'h42a70548, 32'h428506f2, 32'h4234bcd0, 32'hc1d589f5};
test_output[13656:13663] = '{32'h0, 32'h41bd8d93, 32'h0, 32'h429666ba, 32'h42a70548, 32'h428506f2, 32'h4234bcd0, 32'h0};
test_input[13664:13671] = '{32'h429c9bd9, 32'h42207458, 32'h41a72a45, 32'hc25f3b92, 32'h423bc462, 32'h42527a6c, 32'hc2c046de, 32'hc1b7bcb9};
test_output[13664:13671] = '{32'h429c9bd9, 32'h42207458, 32'h41a72a45, 32'h0, 32'h423bc462, 32'h42527a6c, 32'h0, 32'h0};
test_input[13672:13679] = '{32'hc29a6b94, 32'h42ab355b, 32'h41563a98, 32'hc28aebbd, 32'hc20eeb42, 32'h428780d2, 32'hc0a07799, 32'hc2951853};
test_output[13672:13679] = '{32'h0, 32'h42ab355b, 32'h41563a98, 32'h0, 32'h0, 32'h428780d2, 32'h0, 32'h0};
test_input[13680:13687] = '{32'h42c506f3, 32'h40bc58dc, 32'hc2bb784f, 32'h41e32611, 32'h4272e819, 32'h422c17a9, 32'hc2210277, 32'hc27997f5};
test_output[13680:13687] = '{32'h42c506f3, 32'h40bc58dc, 32'h0, 32'h41e32611, 32'h4272e819, 32'h422c17a9, 32'h0, 32'h0};
test_input[13688:13695] = '{32'h41ff9b7c, 32'hc1d9e9b2, 32'hc28a15b3, 32'h42757e0f, 32'hc2203245, 32'hc1c2e7b2, 32'h420e8506, 32'hc283b3d8};
test_output[13688:13695] = '{32'h41ff9b7c, 32'h0, 32'h0, 32'h42757e0f, 32'h0, 32'h0, 32'h420e8506, 32'h0};
test_input[13696:13703] = '{32'h42147d33, 32'h40abad40, 32'h429c0f3d, 32'h41f111c5, 32'hc0306ffe, 32'h4204eca0, 32'hc2365c66, 32'hc160e898};
test_output[13696:13703] = '{32'h42147d33, 32'h40abad40, 32'h429c0f3d, 32'h41f111c5, 32'h0, 32'h4204eca0, 32'h0, 32'h0};
test_input[13704:13711] = '{32'h4240c1a0, 32'h41eb0410, 32'hc2293cb4, 32'h4080b26e, 32'h424d022b, 32'hc29d04b1, 32'h428b37ec, 32'h412c4f1d};
test_output[13704:13711] = '{32'h4240c1a0, 32'h41eb0410, 32'h0, 32'h4080b26e, 32'h424d022b, 32'h0, 32'h428b37ec, 32'h412c4f1d};
test_input[13712:13719] = '{32'h428b14c3, 32'h41171ab5, 32'h428f9c3b, 32'hc2b070eb, 32'hc25fd9b6, 32'hc2afeaba, 32'hc14ad32a, 32'hc21c1fe8};
test_output[13712:13719] = '{32'h428b14c3, 32'h41171ab5, 32'h428f9c3b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13720:13727] = '{32'h42b4e8e7, 32'hc1c2c960, 32'h421239ac, 32'h42c0308c, 32'hc2654cae, 32'h42837cea, 32'hc2887ea7, 32'hc215d9e3};
test_output[13720:13727] = '{32'h42b4e8e7, 32'h0, 32'h421239ac, 32'h42c0308c, 32'h0, 32'h42837cea, 32'h0, 32'h0};
test_input[13728:13735] = '{32'hc2a805ef, 32'h4244ca5b, 32'hc040f7bf, 32'h428c168d, 32'hc106cda0, 32'hc176736a, 32'hc27b0206, 32'hc2c7bc2c};
test_output[13728:13735] = '{32'h0, 32'h4244ca5b, 32'h0, 32'h428c168d, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13736:13743] = '{32'hc29a4096, 32'hc23a4e4b, 32'hc21a0e92, 32'h423d218d, 32'hc18dbf5f, 32'hc1ffdb84, 32'h4289e158, 32'h42586be2};
test_output[13736:13743] = '{32'h0, 32'h0, 32'h0, 32'h423d218d, 32'h0, 32'h0, 32'h4289e158, 32'h42586be2};
test_input[13744:13751] = '{32'h4283ccd8, 32'hc1c3a1bd, 32'h42081976, 32'h42aff2e5, 32'hc25f121c, 32'hc19e7b51, 32'h41cc5da4, 32'h422c501e};
test_output[13744:13751] = '{32'h4283ccd8, 32'h0, 32'h42081976, 32'h42aff2e5, 32'h0, 32'h0, 32'h41cc5da4, 32'h422c501e};
test_input[13752:13759] = '{32'hc2afc5c7, 32'hc29b0f81, 32'hc2125557, 32'h415936bd, 32'h428e3ef1, 32'h4198c7ae, 32'hc181b3b9, 32'hc26f4894};
test_output[13752:13759] = '{32'h0, 32'h0, 32'h0, 32'h415936bd, 32'h428e3ef1, 32'h4198c7ae, 32'h0, 32'h0};
test_input[13760:13767] = '{32'hbfde7084, 32'h40b8b241, 32'hc26575b9, 32'hc18ceb2a, 32'h41a1fada, 32'h42a22116, 32'hc2aed031, 32'hc22143a1};
test_output[13760:13767] = '{32'h0, 32'h40b8b241, 32'h0, 32'h0, 32'h41a1fada, 32'h42a22116, 32'h0, 32'h0};
test_input[13768:13775] = '{32'hc1d0be74, 32'h429684b8, 32'hc2971c44, 32'hc1b23b01, 32'h41a30412, 32'h41b4a93a, 32'hc195bbbb, 32'hc1228a8e};
test_output[13768:13775] = '{32'h0, 32'h429684b8, 32'h0, 32'h0, 32'h41a30412, 32'h41b4a93a, 32'h0, 32'h0};
test_input[13776:13783] = '{32'hc235210b, 32'hc184eadb, 32'h42776d62, 32'hc20d770e, 32'hc20430b8, 32'hc23b9d64, 32'hc2483d02, 32'hc0dfd194};
test_output[13776:13783] = '{32'h0, 32'h0, 32'h42776d62, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13784:13791] = '{32'h42b123b4, 32'hc17520c7, 32'hc1fbbe6e, 32'h4202bfac, 32'h42098b6e, 32'hc29adc11, 32'h423fd12e, 32'hc1816f6c};
test_output[13784:13791] = '{32'h42b123b4, 32'h0, 32'h0, 32'h4202bfac, 32'h42098b6e, 32'h0, 32'h423fd12e, 32'h0};
test_input[13792:13799] = '{32'hc2449869, 32'hc25681d7, 32'hc28e6336, 32'h42871b30, 32'hc20d3004, 32'hc20f131e, 32'h421a1964, 32'hc2325f50};
test_output[13792:13799] = '{32'h0, 32'h0, 32'h0, 32'h42871b30, 32'h0, 32'h0, 32'h421a1964, 32'h0};
test_input[13800:13807] = '{32'hc2a1e2b0, 32'hc22d903b, 32'hc24eb6c1, 32'h423dd563, 32'hc2132a3e, 32'h420235ac, 32'h42a47b3f, 32'hc29fe643};
test_output[13800:13807] = '{32'h0, 32'h0, 32'h0, 32'h423dd563, 32'h0, 32'h420235ac, 32'h42a47b3f, 32'h0};
test_input[13808:13815] = '{32'hc2750c9f, 32'hc21fbb7f, 32'hc212a47b, 32'h4295a5b5, 32'h421405b8, 32'hc2433a4e, 32'hc278ea70, 32'hc1a5bcb1};
test_output[13808:13815] = '{32'h0, 32'h0, 32'h0, 32'h4295a5b5, 32'h421405b8, 32'h0, 32'h0, 32'h0};
test_input[13816:13823] = '{32'h40bf2b4a, 32'hc2487244, 32'hc286b54f, 32'h41d5a078, 32'h42910372, 32'h429808f0, 32'h42b811cd, 32'hc177424f};
test_output[13816:13823] = '{32'h40bf2b4a, 32'h0, 32'h0, 32'h41d5a078, 32'h42910372, 32'h429808f0, 32'h42b811cd, 32'h0};
test_input[13824:13831] = '{32'h42b5c6e5, 32'hc2b25b66, 32'h42bd5599, 32'h42858ff6, 32'h42ade395, 32'hc204b23d, 32'hc259b7f9, 32'h427bf5c4};
test_output[13824:13831] = '{32'h42b5c6e5, 32'h0, 32'h42bd5599, 32'h42858ff6, 32'h42ade395, 32'h0, 32'h0, 32'h427bf5c4};
test_input[13832:13839] = '{32'hc0fc3e6f, 32'h42c35177, 32'h4291a4bc, 32'hc15ae82f, 32'h41655272, 32'hc2b76f28, 32'hc186ec1f, 32'h42a50e99};
test_output[13832:13839] = '{32'h0, 32'h42c35177, 32'h4291a4bc, 32'h0, 32'h41655272, 32'h0, 32'h0, 32'h42a50e99};
test_input[13840:13847] = '{32'hc0eb6bfc, 32'hc2c404e0, 32'h42783e7d, 32'h41e5ae1a, 32'hc227a8ae, 32'h42893a43, 32'h429ab180, 32'hc1cadb3c};
test_output[13840:13847] = '{32'h0, 32'h0, 32'h42783e7d, 32'h41e5ae1a, 32'h0, 32'h42893a43, 32'h429ab180, 32'h0};
test_input[13848:13855] = '{32'h41a04156, 32'hc26c648b, 32'hc1fca074, 32'h4174b14d, 32'hc19c756c, 32'hc1f934d6, 32'hc28b69a3, 32'hc2a6e8e7};
test_output[13848:13855] = '{32'h41a04156, 32'h0, 32'h0, 32'h4174b14d, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13856:13863] = '{32'h4194c31a, 32'h42abb577, 32'h410067ee, 32'h42a0fcca, 32'h42b7d244, 32'hc0c42063, 32'hc28116bd, 32'h428dff1f};
test_output[13856:13863] = '{32'h4194c31a, 32'h42abb577, 32'h410067ee, 32'h42a0fcca, 32'h42b7d244, 32'h0, 32'h0, 32'h428dff1f};
test_input[13864:13871] = '{32'hc23d0799, 32'h42920005, 32'hc23d6f8b, 32'hc23f9098, 32'hc085c181, 32'h4254dc30, 32'h42995457, 32'h41c73dd4};
test_output[13864:13871] = '{32'h0, 32'h42920005, 32'h0, 32'h0, 32'h0, 32'h4254dc30, 32'h42995457, 32'h41c73dd4};
test_input[13872:13879] = '{32'h41bb5afd, 32'hc0be3247, 32'h42c33315, 32'hc2baf184, 32'hc278d88c, 32'hc1938f66, 32'hc2a356d4, 32'hc271a9d4};
test_output[13872:13879] = '{32'h41bb5afd, 32'h0, 32'h42c33315, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13880:13887] = '{32'h41ee475f, 32'hc28a47d2, 32'h41ff7a4b, 32'h42a27d80, 32'h4203ca59, 32'hc2493674, 32'hc20614b3, 32'h427e3372};
test_output[13880:13887] = '{32'h41ee475f, 32'h0, 32'h41ff7a4b, 32'h42a27d80, 32'h4203ca59, 32'h0, 32'h0, 32'h427e3372};
test_input[13888:13895] = '{32'hc2afc5fb, 32'h41c261cd, 32'h42bd53a6, 32'h428bbf59, 32'hbfe9876c, 32'hc2886520, 32'hc299ac5f, 32'h42a849af};
test_output[13888:13895] = '{32'h0, 32'h41c261cd, 32'h42bd53a6, 32'h428bbf59, 32'h0, 32'h0, 32'h0, 32'h42a849af};
test_input[13896:13903] = '{32'hc21bf96f, 32'h428d39c7, 32'h428cd178, 32'h411a67f7, 32'hc2576f4d, 32'hc2a645e2, 32'hc20e8610, 32'h41c9813e};
test_output[13896:13903] = '{32'h0, 32'h428d39c7, 32'h428cd178, 32'h411a67f7, 32'h0, 32'h0, 32'h0, 32'h41c9813e};
test_input[13904:13911] = '{32'hc2778ee2, 32'h4295f8da, 32'h427ff91b, 32'hc2722fb9, 32'hc2034cd6, 32'h41951bbc, 32'h414adff1, 32'h42a99889};
test_output[13904:13911] = '{32'h0, 32'h4295f8da, 32'h427ff91b, 32'h0, 32'h0, 32'h41951bbc, 32'h414adff1, 32'h42a99889};
test_input[13912:13919] = '{32'h42b7a8b4, 32'hc26c580d, 32'h4295c3e4, 32'h428f7326, 32'hc297a1cf, 32'hc13be037, 32'h425e2905, 32'h42ab4013};
test_output[13912:13919] = '{32'h42b7a8b4, 32'h0, 32'h4295c3e4, 32'h428f7326, 32'h0, 32'h0, 32'h425e2905, 32'h42ab4013};
test_input[13920:13927] = '{32'h4292b27a, 32'hc16c6662, 32'hc0f9010e, 32'h4286e01d, 32'h4283301a, 32'h421e411e, 32'h4279ed87, 32'h42801c55};
test_output[13920:13927] = '{32'h4292b27a, 32'h0, 32'h0, 32'h4286e01d, 32'h4283301a, 32'h421e411e, 32'h4279ed87, 32'h42801c55};
test_input[13928:13935] = '{32'h42876789, 32'hc24af4e6, 32'hc2ba0194, 32'h41308dc6, 32'hc1a03547, 32'hc16fef75, 32'h41190fb1, 32'hc18f67e5};
test_output[13928:13935] = '{32'h42876789, 32'h0, 32'h0, 32'h41308dc6, 32'h0, 32'h0, 32'h41190fb1, 32'h0};
test_input[13936:13943] = '{32'h42b62f70, 32'hc2701d10, 32'hc2c6be26, 32'hc10c4974, 32'h42c1dc72, 32'h42c3a14e, 32'h42ad370b, 32'h42337c70};
test_output[13936:13943] = '{32'h42b62f70, 32'h0, 32'h0, 32'h0, 32'h42c1dc72, 32'h42c3a14e, 32'h42ad370b, 32'h42337c70};
test_input[13944:13951] = '{32'hc2af0389, 32'hc0d670ff, 32'h42bdbf45, 32'h40d36dab, 32'hc205eb1d, 32'hc2a05d90, 32'hc21fd0c7, 32'hc1f5b400};
test_output[13944:13951] = '{32'h0, 32'h0, 32'h42bdbf45, 32'h40d36dab, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[13952:13959] = '{32'hc1965265, 32'hc1061322, 32'hc293a7aa, 32'h422ce9da, 32'hc276f985, 32'hc1e38fc7, 32'hc2adb1ae, 32'h40ee91ee};
test_output[13952:13959] = '{32'h0, 32'h0, 32'h0, 32'h422ce9da, 32'h0, 32'h0, 32'h0, 32'h40ee91ee};
test_input[13960:13967] = '{32'h4190120c, 32'hc11ceb4a, 32'h42468e15, 32'h42490b45, 32'h42710b00, 32'hc2b65c37, 32'hc280d1b6, 32'hc17f7332};
test_output[13960:13967] = '{32'h4190120c, 32'h0, 32'h42468e15, 32'h42490b45, 32'h42710b00, 32'h0, 32'h0, 32'h0};
test_input[13968:13975] = '{32'hc1864782, 32'h423da031, 32'hc2967964, 32'hc2859dd1, 32'h41a71c64, 32'hc2b92ae1, 32'hc01239f3, 32'h418a081d};
test_output[13968:13975] = '{32'h0, 32'h423da031, 32'h0, 32'h0, 32'h41a71c64, 32'h0, 32'h0, 32'h418a081d};
test_input[13976:13983] = '{32'hc2c510a6, 32'h422e94c5, 32'h42719bec, 32'hc2a4bbcc, 32'h421d2814, 32'h4269dcde, 32'h41c8f61f, 32'hc26a6123};
test_output[13976:13983] = '{32'h0, 32'h422e94c5, 32'h42719bec, 32'h0, 32'h421d2814, 32'h4269dcde, 32'h41c8f61f, 32'h0};
test_input[13984:13991] = '{32'hbf8d8e4f, 32'hc21aa6da, 32'hc1739211, 32'h42bfdf0d, 32'hc298c85b, 32'h4247da6b, 32'h42bf41b3, 32'h41a32a8b};
test_output[13984:13991] = '{32'h0, 32'h0, 32'h0, 32'h42bfdf0d, 32'h0, 32'h4247da6b, 32'h42bf41b3, 32'h41a32a8b};
test_input[13992:13999] = '{32'hc2b4824c, 32'h428505ec, 32'hc1fcd196, 32'hc0b9eee5, 32'hc26d4091, 32'h42aa91b1, 32'hc1863e9c, 32'h41bfb0c4};
test_output[13992:13999] = '{32'h0, 32'h428505ec, 32'h0, 32'h0, 32'h0, 32'h42aa91b1, 32'h0, 32'h41bfb0c4};
test_input[14000:14007] = '{32'h42253523, 32'h4257036f, 32'hc1c005cc, 32'h42b68fe9, 32'h41f90f63, 32'hbfd06511, 32'h426fe828, 32'h4227d51a};
test_output[14000:14007] = '{32'h42253523, 32'h4257036f, 32'h0, 32'h42b68fe9, 32'h41f90f63, 32'h0, 32'h426fe828, 32'h4227d51a};
test_input[14008:14015] = '{32'h41168121, 32'hc1b911bd, 32'hc287ce84, 32'h42aad90a, 32'h41e8d4ff, 32'h41db79d5, 32'h41eaf946, 32'hc20a1f16};
test_output[14008:14015] = '{32'h41168121, 32'h0, 32'h0, 32'h42aad90a, 32'h41e8d4ff, 32'h41db79d5, 32'h41eaf946, 32'h0};
test_input[14016:14023] = '{32'hc255dfe9, 32'h4148d9d0, 32'h41ce1e4f, 32'h416dc2f2, 32'h42458468, 32'hc29f689c, 32'h42a71b92, 32'h42ae4dab};
test_output[14016:14023] = '{32'h0, 32'h4148d9d0, 32'h41ce1e4f, 32'h416dc2f2, 32'h42458468, 32'h0, 32'h42a71b92, 32'h42ae4dab};
test_input[14024:14031] = '{32'h429e08e7, 32'h42a71d22, 32'h4257de29, 32'h427b5d00, 32'hc195ba69, 32'h415586b5, 32'h422cab2b, 32'h4147995e};
test_output[14024:14031] = '{32'h429e08e7, 32'h42a71d22, 32'h4257de29, 32'h427b5d00, 32'h0, 32'h415586b5, 32'h422cab2b, 32'h4147995e};
test_input[14032:14039] = '{32'h42a1553d, 32'h429a600c, 32'h4294bbb1, 32'hc21aaacd, 32'hc1e74611, 32'h42160fdd, 32'h4227d620, 32'h403a9777};
test_output[14032:14039] = '{32'h42a1553d, 32'h429a600c, 32'h4294bbb1, 32'h0, 32'h0, 32'h42160fdd, 32'h4227d620, 32'h403a9777};
test_input[14040:14047] = '{32'h40bb3dc8, 32'h42202851, 32'h42416376, 32'h41d14afb, 32'hc26869a1, 32'h424d2165, 32'hc10eb4b9, 32'h426911fe};
test_output[14040:14047] = '{32'h40bb3dc8, 32'h42202851, 32'h42416376, 32'h41d14afb, 32'h0, 32'h424d2165, 32'h0, 32'h426911fe};
test_input[14048:14055] = '{32'hc24aeb75, 32'hc22c510a, 32'h421c283a, 32'h40eed189, 32'hc25320d2, 32'h41561873, 32'h424fa9c9, 32'hc10eef11};
test_output[14048:14055] = '{32'h0, 32'h0, 32'h421c283a, 32'h40eed189, 32'h0, 32'h41561873, 32'h424fa9c9, 32'h0};
test_input[14056:14063] = '{32'h4280c743, 32'hc10084f2, 32'hc19dcd26, 32'h41d26df9, 32'h4244efc4, 32'hc28bc636, 32'hc29ce77e, 32'hc2bb6dab};
test_output[14056:14063] = '{32'h4280c743, 32'h0, 32'h0, 32'h41d26df9, 32'h4244efc4, 32'h0, 32'h0, 32'h0};
test_input[14064:14071] = '{32'hc226aafe, 32'hc1db4be5, 32'hc0ed7d52, 32'hc2c7cd9b, 32'h426a2ab6, 32'h3f15d8c9, 32'h42aec982, 32'h4281f0f8};
test_output[14064:14071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h426a2ab6, 32'h3f15d8c9, 32'h42aec982, 32'h4281f0f8};
test_input[14072:14079] = '{32'h42bf8207, 32'h429fbfe8, 32'hc26a6a26, 32'hc2ad9081, 32'hc1d81ed1, 32'hc2bf0fb7, 32'hc159486b, 32'h419026fd};
test_output[14072:14079] = '{32'h42bf8207, 32'h429fbfe8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h419026fd};
test_input[14080:14087] = '{32'hbdbc70d0, 32'hc2917f00, 32'h42574b09, 32'hc1e2cd3a, 32'h41fd6e81, 32'hc2877fb1, 32'h423d821b, 32'hc2b07ff2};
test_output[14080:14087] = '{32'h0, 32'h0, 32'h42574b09, 32'h0, 32'h41fd6e81, 32'h0, 32'h423d821b, 32'h0};
test_input[14088:14095] = '{32'h429bc80f, 32'hc26ee708, 32'hbf373f70, 32'h42bf25a4, 32'h4204802f, 32'h4126d353, 32'h4288e53f, 32'h428118b4};
test_output[14088:14095] = '{32'h429bc80f, 32'h0, 32'h0, 32'h42bf25a4, 32'h4204802f, 32'h4126d353, 32'h4288e53f, 32'h428118b4};
test_input[14096:14103] = '{32'h423ad069, 32'h4281f74f, 32'h4285aa03, 32'hc0c4f6db, 32'h42941e93, 32'hc2aafb2f, 32'h42a45971, 32'hc2c641b7};
test_output[14096:14103] = '{32'h423ad069, 32'h4281f74f, 32'h4285aa03, 32'h0, 32'h42941e93, 32'h0, 32'h42a45971, 32'h0};
test_input[14104:14111] = '{32'h42954969, 32'hc2adaa04, 32'hc29a5df2, 32'h4218832f, 32'hc2b4c6d9, 32'h4283af81, 32'h3fc730bf, 32'hc216be8d};
test_output[14104:14111] = '{32'h42954969, 32'h0, 32'h0, 32'h4218832f, 32'h0, 32'h4283af81, 32'h3fc730bf, 32'h0};
test_input[14112:14119] = '{32'h422ca58f, 32'h42c593ea, 32'h41cbf5e3, 32'h42936070, 32'h4211a851, 32'hc2a78eff, 32'hc21bd4b7, 32'hc0fbc161};
test_output[14112:14119] = '{32'h422ca58f, 32'h42c593ea, 32'h41cbf5e3, 32'h42936070, 32'h4211a851, 32'h0, 32'h0, 32'h0};
test_input[14120:14127] = '{32'hc2853ed1, 32'h422bf120, 32'h429edcfa, 32'hc2aa6daf, 32'hc2934a90, 32'h42c3567a, 32'h41c572c4, 32'h420fbc61};
test_output[14120:14127] = '{32'h0, 32'h422bf120, 32'h429edcfa, 32'h0, 32'h0, 32'h42c3567a, 32'h41c572c4, 32'h420fbc61};
test_input[14128:14135] = '{32'h42b394f0, 32'h40073a5e, 32'h429230b1, 32'h423503aa, 32'h41998953, 32'h429fe2ea, 32'hbfb91a2e, 32'h41aae351};
test_output[14128:14135] = '{32'h42b394f0, 32'h40073a5e, 32'h429230b1, 32'h423503aa, 32'h41998953, 32'h429fe2ea, 32'h0, 32'h41aae351};
test_input[14136:14143] = '{32'h42ad9b01, 32'h42153f83, 32'hc2497e3c, 32'hc17ad30b, 32'h418723c5, 32'h4232ec04, 32'h42c63cb1, 32'hc29c1aa7};
test_output[14136:14143] = '{32'h42ad9b01, 32'h42153f83, 32'h0, 32'h0, 32'h418723c5, 32'h4232ec04, 32'h42c63cb1, 32'h0};
test_input[14144:14151] = '{32'hc2bcf67c, 32'h40e2796d, 32'hc28f26e2, 32'h41c2fcc9, 32'h423582d1, 32'h421a1a00, 32'hc295ff47, 32'h42c5399c};
test_output[14144:14151] = '{32'h0, 32'h40e2796d, 32'h0, 32'h41c2fcc9, 32'h423582d1, 32'h421a1a00, 32'h0, 32'h42c5399c};
test_input[14152:14159] = '{32'hc2bd4c0c, 32'h4209cc92, 32'hc199cbda, 32'hbfff09f4, 32'hc25f3195, 32'h41df696b, 32'hc2c09f7d, 32'hc265e978};
test_output[14152:14159] = '{32'h0, 32'h4209cc92, 32'h0, 32'h0, 32'h0, 32'h41df696b, 32'h0, 32'h0};
test_input[14160:14167] = '{32'hc25c5d41, 32'hc251dcd4, 32'h42a83134, 32'h4257dd06, 32'hc2b2ca23, 32'hc288e8b8, 32'hc2a340c2, 32'h429aae4e};
test_output[14160:14167] = '{32'h0, 32'h0, 32'h42a83134, 32'h4257dd06, 32'h0, 32'h0, 32'h0, 32'h429aae4e};
test_input[14168:14175] = '{32'hc29876eb, 32'h40865985, 32'h42b92e8c, 32'h41a2665f, 32'hc2646786, 32'h425b7948, 32'h418323ba, 32'h4212630e};
test_output[14168:14175] = '{32'h0, 32'h40865985, 32'h42b92e8c, 32'h41a2665f, 32'h0, 32'h425b7948, 32'h418323ba, 32'h4212630e};
test_input[14176:14183] = '{32'hc2127aae, 32'hbf75d8f2, 32'hc24d757a, 32'h4221d05b, 32'h4241e2fb, 32'h42bb02d4, 32'hc24ef102, 32'hc2c75532};
test_output[14176:14183] = '{32'h0, 32'h0, 32'h0, 32'h4221d05b, 32'h4241e2fb, 32'h42bb02d4, 32'h0, 32'h0};
test_input[14184:14191] = '{32'h42b50cca, 32'h3f209b70, 32'hc08edec1, 32'h416bb0fd, 32'h41de536a, 32'hc1c2da6c, 32'h42a8017c, 32'h42930c55};
test_output[14184:14191] = '{32'h42b50cca, 32'h3f209b70, 32'h0, 32'h416bb0fd, 32'h41de536a, 32'h0, 32'h42a8017c, 32'h42930c55};
test_input[14192:14199] = '{32'h417201fb, 32'h42c42b2c, 32'hc2932cca, 32'h4281baaa, 32'hc2572f60, 32'h423b5817, 32'h421c1c39, 32'h41d4f248};
test_output[14192:14199] = '{32'h417201fb, 32'h42c42b2c, 32'h0, 32'h4281baaa, 32'h0, 32'h423b5817, 32'h421c1c39, 32'h41d4f248};
test_input[14200:14207] = '{32'h42bbf891, 32'h42221988, 32'h4082252d, 32'h4239d81e, 32'h4128c5df, 32'h40f9594c, 32'h41ea4d66, 32'h429e3e9a};
test_output[14200:14207] = '{32'h42bbf891, 32'h42221988, 32'h4082252d, 32'h4239d81e, 32'h4128c5df, 32'h40f9594c, 32'h41ea4d66, 32'h429e3e9a};
test_input[14208:14215] = '{32'h42425b73, 32'hc2348fa3, 32'hc2c1a8af, 32'h42c37e3b, 32'hc28a8868, 32'hc20a15b4, 32'hc2655a9c, 32'hc28c96fa};
test_output[14208:14215] = '{32'h42425b73, 32'h0, 32'h0, 32'h42c37e3b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14216:14223] = '{32'h4282b7f0, 32'hc167e2be, 32'h42a5aa9a, 32'hc212bbfa, 32'h41eabbdc, 32'hc2999222, 32'hc22ba8ba, 32'hc29c5558};
test_output[14216:14223] = '{32'h4282b7f0, 32'h0, 32'h42a5aa9a, 32'h0, 32'h41eabbdc, 32'h0, 32'h0, 32'h0};
test_input[14224:14231] = '{32'hc1618ea6, 32'hc1607940, 32'h42ae7c8d, 32'hc1815be7, 32'hc23fcabc, 32'h4225ba3b, 32'hc291d14c, 32'h4292a731};
test_output[14224:14231] = '{32'h0, 32'h0, 32'h42ae7c8d, 32'h0, 32'h0, 32'h4225ba3b, 32'h0, 32'h4292a731};
test_input[14232:14239] = '{32'h42aadd9f, 32'hc019655e, 32'h42277da9, 32'hc2aec186, 32'hc26b2183, 32'hc1b57674, 32'h42bd8798, 32'hc28b6f7f};
test_output[14232:14239] = '{32'h42aadd9f, 32'h0, 32'h42277da9, 32'h0, 32'h0, 32'h0, 32'h42bd8798, 32'h0};
test_input[14240:14247] = '{32'h41f318d6, 32'h4278116f, 32'hc292a6a2, 32'hc27e9bc7, 32'hc27fd4ec, 32'h4268d1dd, 32'hc1c45ab5, 32'h4289c215};
test_output[14240:14247] = '{32'h41f318d6, 32'h4278116f, 32'h0, 32'h0, 32'h0, 32'h4268d1dd, 32'h0, 32'h4289c215};
test_input[14248:14255] = '{32'h42827e7f, 32'hc1fa3f9e, 32'hc140fa92, 32'h4247e63d, 32'hc1e861d2, 32'h42c514e9, 32'hc27f5f4e, 32'hc1ab1893};
test_output[14248:14255] = '{32'h42827e7f, 32'h0, 32'h0, 32'h4247e63d, 32'h0, 32'h42c514e9, 32'h0, 32'h0};
test_input[14256:14263] = '{32'hc28079c6, 32'h4107813a, 32'hc225cbef, 32'hc19a663d, 32'h40ad615d, 32'hc1a3f0fb, 32'hc2671084, 32'hc2a7665e};
test_output[14256:14263] = '{32'h0, 32'h4107813a, 32'h0, 32'h0, 32'h40ad615d, 32'h0, 32'h0, 32'h0};
test_input[14264:14271] = '{32'hc25e5403, 32'h41f070b6, 32'hc271a817, 32'hc1e43527, 32'hc27b15af, 32'h426bb5fb, 32'hc1099772, 32'h414dc4ca};
test_output[14264:14271] = '{32'h0, 32'h41f070b6, 32'h0, 32'h0, 32'h0, 32'h426bb5fb, 32'h0, 32'h414dc4ca};
test_input[14272:14279] = '{32'h424ac089, 32'hc2b8c080, 32'h425130d9, 32'h41e9dc1c, 32'hc045c495, 32'hbfb4e0e6, 32'hc283643b, 32'hc2bbe7da};
test_output[14272:14279] = '{32'h424ac089, 32'h0, 32'h425130d9, 32'h41e9dc1c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14280:14287] = '{32'h40b90792, 32'hc27ef9f3, 32'hc2c414d5, 32'hc23abec4, 32'hc283d4f5, 32'hc2c3b6be, 32'hc19fd185, 32'h41c4dc54};
test_output[14280:14287] = '{32'h40b90792, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41c4dc54};
test_input[14288:14295] = '{32'hc26da33b, 32'h42005bd0, 32'h413dd9ed, 32'h428a4174, 32'h421b6bf6, 32'hc1d0e5bb, 32'hc04dbd47, 32'hc26484f5};
test_output[14288:14295] = '{32'h0, 32'h42005bd0, 32'h413dd9ed, 32'h428a4174, 32'h421b6bf6, 32'h0, 32'h0, 32'h0};
test_input[14296:14303] = '{32'hc1e05d5e, 32'hc21796b6, 32'h427db603, 32'hc22d8992, 32'h4084fe4f, 32'h42973f2e, 32'h421f507e, 32'h420513cb};
test_output[14296:14303] = '{32'h0, 32'h0, 32'h427db603, 32'h0, 32'h4084fe4f, 32'h42973f2e, 32'h421f507e, 32'h420513cb};
test_input[14304:14311] = '{32'hc101f931, 32'hc29be9bf, 32'hc1931fb1, 32'hc2849856, 32'h428adebb, 32'h4291dc55, 32'h429f878d, 32'h42bf1d35};
test_output[14304:14311] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h428adebb, 32'h4291dc55, 32'h429f878d, 32'h42bf1d35};
test_input[14312:14319] = '{32'h42887fd1, 32'hc280c4fc, 32'h4180b6a6, 32'h4285e762, 32'h42bfaae8, 32'h41eec8bf, 32'h41a463df, 32'h40c568a0};
test_output[14312:14319] = '{32'h42887fd1, 32'h0, 32'h4180b6a6, 32'h4285e762, 32'h42bfaae8, 32'h41eec8bf, 32'h41a463df, 32'h40c568a0};
test_input[14320:14327] = '{32'h42983775, 32'h41c8352d, 32'hc22a00da, 32'h42828e39, 32'hc21cfe42, 32'h4188f4b8, 32'h41c9f4b2, 32'hc115b82f};
test_output[14320:14327] = '{32'h42983775, 32'h41c8352d, 32'h0, 32'h42828e39, 32'h0, 32'h4188f4b8, 32'h41c9f4b2, 32'h0};
test_input[14328:14335] = '{32'hc1d1acf0, 32'hc296e8e6, 32'hc2a8082f, 32'hc0ce68e9, 32'h42a82b02, 32'h42b34c26, 32'hc189cc79, 32'hc236ff9e};
test_output[14328:14335] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a82b02, 32'h42b34c26, 32'h0, 32'h0};
test_input[14336:14343] = '{32'hc287a222, 32'hc0dadf07, 32'h41b2495d, 32'hc263900c, 32'hc2b6a5fb, 32'hc29a3b21, 32'h3f8f854c, 32'hc06c7124};
test_output[14336:14343] = '{32'h0, 32'h0, 32'h41b2495d, 32'h0, 32'h0, 32'h0, 32'h3f8f854c, 32'h0};
test_input[14344:14351] = '{32'hc0be166a, 32'hc27482ce, 32'hc0ce8a3e, 32'h41edf5c3, 32'h425fe0c6, 32'hc2a9948d, 32'hc1b4f62f, 32'hc2adb9ba};
test_output[14344:14351] = '{32'h0, 32'h0, 32'h0, 32'h41edf5c3, 32'h425fe0c6, 32'h0, 32'h0, 32'h0};
test_input[14352:14359] = '{32'hc0b0696b, 32'hc1ca038b, 32'hc2114537, 32'h4141d23a, 32'hc2b9f879, 32'hc2b2fa07, 32'h42724036, 32'hc2bd3aa7};
test_output[14352:14359] = '{32'h0, 32'h0, 32'h0, 32'h4141d23a, 32'h0, 32'h0, 32'h42724036, 32'h0};
test_input[14360:14367] = '{32'h42c3215f, 32'hc20f7426, 32'h41dd0e03, 32'h4112f60c, 32'hc03fbd2c, 32'h419ee832, 32'h4291fa8a, 32'h41a9ba8a};
test_output[14360:14367] = '{32'h42c3215f, 32'h0, 32'h41dd0e03, 32'h4112f60c, 32'h0, 32'h419ee832, 32'h4291fa8a, 32'h41a9ba8a};
test_input[14368:14375] = '{32'hc291e198, 32'hc24aee89, 32'h4155ad44, 32'hc2c2819f, 32'h429de67b, 32'hc28abb12, 32'hc287531f, 32'h42b1fe44};
test_output[14368:14375] = '{32'h0, 32'h0, 32'h4155ad44, 32'h0, 32'h429de67b, 32'h0, 32'h0, 32'h42b1fe44};
test_input[14376:14383] = '{32'h42501469, 32'hc1b05232, 32'h4299663f, 32'h413597ef, 32'hc2a72d96, 32'hc27caaa6, 32'hc2041016, 32'h41c95dbe};
test_output[14376:14383] = '{32'h42501469, 32'h0, 32'h4299663f, 32'h413597ef, 32'h0, 32'h0, 32'h0, 32'h41c95dbe};
test_input[14384:14391] = '{32'h40d7b1e4, 32'h42889b11, 32'h423e5154, 32'h42b3befa, 32'hc1979920, 32'hc2ae9f82, 32'h40661738, 32'hc225b47b};
test_output[14384:14391] = '{32'h40d7b1e4, 32'h42889b11, 32'h423e5154, 32'h42b3befa, 32'h0, 32'h0, 32'h40661738, 32'h0};
test_input[14392:14399] = '{32'hc2bd916d, 32'h42921623, 32'hc2077fc0, 32'hc2845bca, 32'h4064cf1f, 32'hc24168a0, 32'hc2272897, 32'hc2a3d1fc};
test_output[14392:14399] = '{32'h0, 32'h42921623, 32'h0, 32'h0, 32'h4064cf1f, 32'h0, 32'h0, 32'h0};
test_input[14400:14407] = '{32'hc2ac30d6, 32'h40981935, 32'h41fe8fab, 32'hc22ace2f, 32'h426f93a2, 32'hc14a2827, 32'h429d9716, 32'hc2c0809b};
test_output[14400:14407] = '{32'h0, 32'h40981935, 32'h41fe8fab, 32'h0, 32'h426f93a2, 32'h0, 32'h429d9716, 32'h0};
test_input[14408:14415] = '{32'hc2a67557, 32'hc2b3ce81, 32'h42b7b93e, 32'hc2332f2d, 32'hc29f00a9, 32'hc25c0462, 32'hc1f1854f, 32'hc22a8a11};
test_output[14408:14415] = '{32'h0, 32'h0, 32'h42b7b93e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14416:14423] = '{32'hc2609d16, 32'hc2af0a4d, 32'hc29f1214, 32'h42392a2b, 32'h41aff919, 32'h418949af, 32'hc0bc0668, 32'hc1c1d940};
test_output[14416:14423] = '{32'h0, 32'h0, 32'h0, 32'h42392a2b, 32'h41aff919, 32'h418949af, 32'h0, 32'h0};
test_input[14424:14431] = '{32'h41125e03, 32'h41f3167c, 32'h421ead45, 32'h4182728d, 32'hc29b5b7e, 32'h419242b3, 32'hc2727fd7, 32'h42c63342};
test_output[14424:14431] = '{32'h41125e03, 32'h41f3167c, 32'h421ead45, 32'h4182728d, 32'h0, 32'h419242b3, 32'h0, 32'h42c63342};
test_input[14432:14439] = '{32'h427597c1, 32'hc15f6a7a, 32'hc0c9a3b6, 32'hc1da7730, 32'h40ada5cc, 32'hc2b68e9b, 32'hc2b349da, 32'h429dff65};
test_output[14432:14439] = '{32'h427597c1, 32'h0, 32'h0, 32'h0, 32'h40ada5cc, 32'h0, 32'h0, 32'h429dff65};
test_input[14440:14447] = '{32'h42b80752, 32'h4193f5bb, 32'hc1cb8fe9, 32'hc1b84090, 32'hc15ed521, 32'h416c82dd, 32'h415ddcab, 32'h4221f716};
test_output[14440:14447] = '{32'h42b80752, 32'h4193f5bb, 32'h0, 32'h0, 32'h0, 32'h416c82dd, 32'h415ddcab, 32'h4221f716};
test_input[14448:14455] = '{32'hc1f35bf9, 32'h4195b326, 32'h40f312e9, 32'h41ba3834, 32'h428468a6, 32'hc0ec5cc4, 32'h42a3c03d, 32'hc2a64cb2};
test_output[14448:14455] = '{32'h0, 32'h4195b326, 32'h40f312e9, 32'h41ba3834, 32'h428468a6, 32'h0, 32'h42a3c03d, 32'h0};
test_input[14456:14463] = '{32'h42b9def7, 32'hc2076f4e, 32'h42b0e7e5, 32'h42352725, 32'hc097f805, 32'hc1fb8dcd, 32'h41eb25ec, 32'hc24afe52};
test_output[14456:14463] = '{32'h42b9def7, 32'h0, 32'h42b0e7e5, 32'h42352725, 32'h0, 32'h0, 32'h41eb25ec, 32'h0};
test_input[14464:14471] = '{32'h42af4d48, 32'h41bebaa1, 32'hc03f89d0, 32'h42a46fb5, 32'h42545658, 32'h41d75a94, 32'hc25b0d6c, 32'hc1c1f793};
test_output[14464:14471] = '{32'h42af4d48, 32'h41bebaa1, 32'h0, 32'h42a46fb5, 32'h42545658, 32'h41d75a94, 32'h0, 32'h0};
test_input[14472:14479] = '{32'hbf05e9ed, 32'hc1d43817, 32'hc248b0d2, 32'h410b7f80, 32'hc2a2878e, 32'hc2191c72, 32'hc2738e73, 32'hc25ad615};
test_output[14472:14479] = '{32'h0, 32'h0, 32'h0, 32'h410b7f80, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14480:14487] = '{32'h426e2d4d, 32'hc169b389, 32'h41ee78e6, 32'h417c160e, 32'hc2984adf, 32'hc25e8137, 32'hc2aa06f9, 32'h42c5365d};
test_output[14480:14487] = '{32'h426e2d4d, 32'h0, 32'h41ee78e6, 32'h417c160e, 32'h0, 32'h0, 32'h0, 32'h42c5365d};
test_input[14488:14495] = '{32'hc28417e0, 32'h412b1898, 32'h429dfabd, 32'h4146d11f, 32'h429b7640, 32'h4261f741, 32'hc28f294f, 32'h41a6992b};
test_output[14488:14495] = '{32'h0, 32'h412b1898, 32'h429dfabd, 32'h4146d11f, 32'h429b7640, 32'h4261f741, 32'h0, 32'h41a6992b};
test_input[14496:14503] = '{32'h3f641c0c, 32'h41a9fe7f, 32'h42311330, 32'hc2a8983e, 32'h428808f1, 32'hc2820415, 32'h42269eb5, 32'h41c711e2};
test_output[14496:14503] = '{32'h3f641c0c, 32'h41a9fe7f, 32'h42311330, 32'h0, 32'h428808f1, 32'h0, 32'h42269eb5, 32'h41c711e2};
test_input[14504:14511] = '{32'h42b8572b, 32'hc249a510, 32'hc225d0ea, 32'h4135e251, 32'h423c1bbd, 32'h42866d47, 32'h418e98a2, 32'h42a4d812};
test_output[14504:14511] = '{32'h42b8572b, 32'h0, 32'h0, 32'h4135e251, 32'h423c1bbd, 32'h42866d47, 32'h418e98a2, 32'h42a4d812};
test_input[14512:14519] = '{32'h40773dea, 32'hc2aaf832, 32'h42a598f1, 32'hc22a52a0, 32'h425b19a1, 32'h419a6318, 32'h4285b6f7, 32'h41e3defa};
test_output[14512:14519] = '{32'h40773dea, 32'h0, 32'h42a598f1, 32'h0, 32'h425b19a1, 32'h419a6318, 32'h4285b6f7, 32'h41e3defa};
test_input[14520:14527] = '{32'hc2c02875, 32'hc1e95d33, 32'h42525fb6, 32'h41c443fc, 32'h41cd0193, 32'hc2900603, 32'h42c1d536, 32'hc25617e5};
test_output[14520:14527] = '{32'h0, 32'h0, 32'h42525fb6, 32'h41c443fc, 32'h41cd0193, 32'h0, 32'h42c1d536, 32'h0};
test_input[14528:14535] = '{32'hc28b63b1, 32'h3faed1fc, 32'h416710d4, 32'hc2c5e737, 32'hc2563801, 32'hc245e488, 32'hc20e2011, 32'hc276bf4e};
test_output[14528:14535] = '{32'h0, 32'h3faed1fc, 32'h416710d4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14536:14543] = '{32'h42c654ff, 32'h41e7b1ea, 32'hc0da826f, 32'h41d809e2, 32'h42ab610e, 32'h41daad9f, 32'h3ead6cd8, 32'h422a25ae};
test_output[14536:14543] = '{32'h42c654ff, 32'h41e7b1ea, 32'h0, 32'h41d809e2, 32'h42ab610e, 32'h41daad9f, 32'h3ead6cd8, 32'h422a25ae};
test_input[14544:14551] = '{32'h40fc94cb, 32'hc2b41ffe, 32'hc286a2e9, 32'hc291b297, 32'h4291bf54, 32'hc185d653, 32'h423af5f1, 32'hc2c2636e};
test_output[14544:14551] = '{32'h40fc94cb, 32'h0, 32'h0, 32'h0, 32'h4291bf54, 32'h0, 32'h423af5f1, 32'h0};
test_input[14552:14559] = '{32'hc1d1558b, 32'hc2868507, 32'hc23e1354, 32'hc081c1f1, 32'hc27ed1c1, 32'h420d8a46, 32'h42938ffb, 32'hc286f842};
test_output[14552:14559] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420d8a46, 32'h42938ffb, 32'h0};
test_input[14560:14567] = '{32'h42304252, 32'hc2c5c95a, 32'hc243368d, 32'h42806ebd, 32'h412bd37c, 32'hc2ae3278, 32'h4282d2e0, 32'h42b52563};
test_output[14560:14567] = '{32'h42304252, 32'h0, 32'h0, 32'h42806ebd, 32'h412bd37c, 32'h0, 32'h4282d2e0, 32'h42b52563};
test_input[14568:14575] = '{32'h423e26df, 32'h415abee1, 32'hc29c9b95, 32'h42b9b417, 32'hc2733581, 32'h4267628f, 32'hc291ec5f, 32'hc1f92c6b};
test_output[14568:14575] = '{32'h423e26df, 32'h415abee1, 32'h0, 32'h42b9b417, 32'h0, 32'h4267628f, 32'h0, 32'h0};
test_input[14576:14583] = '{32'hc11f51c5, 32'hc2852e6c, 32'hc23bd99b, 32'hc1de9a1c, 32'hc29940a1, 32'h42b19799, 32'hc2c3f998, 32'h40a639ba};
test_output[14576:14583] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b19799, 32'h0, 32'h40a639ba};
test_input[14584:14591] = '{32'h4287417c, 32'h41c7e16c, 32'hc1c4b2af, 32'h42a70422, 32'hc1373398, 32'h4269d492, 32'hc2b7cfa1, 32'hc2478325};
test_output[14584:14591] = '{32'h4287417c, 32'h41c7e16c, 32'h0, 32'h42a70422, 32'h0, 32'h4269d492, 32'h0, 32'h0};
test_input[14592:14599] = '{32'h42baba18, 32'hc05e8d37, 32'h429d0c09, 32'h41b129a2, 32'hc29d691f, 32'hc1d703e1, 32'hc1ee8f0e, 32'hc2b0fd2e};
test_output[14592:14599] = '{32'h42baba18, 32'h0, 32'h429d0c09, 32'h41b129a2, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14600:14607] = '{32'h41bf3058, 32'hc20a7799, 32'hc272edcc, 32'hc2809b52, 32'h416a9c42, 32'hc28eab6a, 32'h4210014d, 32'hc26448d6};
test_output[14600:14607] = '{32'h41bf3058, 32'h0, 32'h0, 32'h0, 32'h416a9c42, 32'h0, 32'h4210014d, 32'h0};
test_input[14608:14615] = '{32'h414f41ae, 32'h41fbf521, 32'hc23a89dc, 32'h426165f7, 32'h41c5fa01, 32'hc2b643e3, 32'h426923a0, 32'hc18f80c7};
test_output[14608:14615] = '{32'h414f41ae, 32'h41fbf521, 32'h0, 32'h426165f7, 32'h41c5fa01, 32'h0, 32'h426923a0, 32'h0};
test_input[14616:14623] = '{32'hc1213c8a, 32'h42149f7b, 32'hc21d01d5, 32'hc1589170, 32'hc24fbfbd, 32'h4219cc0c, 32'h40ae50fb, 32'h4268070c};
test_output[14616:14623] = '{32'h0, 32'h42149f7b, 32'h0, 32'h0, 32'h0, 32'h4219cc0c, 32'h40ae50fb, 32'h4268070c};
test_input[14624:14631] = '{32'hc27b19b7, 32'h4250aae3, 32'h420c6b8c, 32'h4152c164, 32'hbf00f330, 32'hc2c406fa, 32'hc2924b58, 32'hc12791b0};
test_output[14624:14631] = '{32'h0, 32'h4250aae3, 32'h420c6b8c, 32'h4152c164, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14632:14639] = '{32'hc088df08, 32'hc212af1d, 32'h426c0be6, 32'hc2995da1, 32'h42920153, 32'hc27a766f, 32'hc068c5ab, 32'h427ab778};
test_output[14632:14639] = '{32'h0, 32'h0, 32'h426c0be6, 32'h0, 32'h42920153, 32'h0, 32'h0, 32'h427ab778};
test_input[14640:14647] = '{32'h42a2a6d5, 32'h4234863f, 32'h4101cd11, 32'hc23de547, 32'h42a18ead, 32'h41705ee1, 32'h41a477a4, 32'hc23025e4};
test_output[14640:14647] = '{32'h42a2a6d5, 32'h4234863f, 32'h4101cd11, 32'h0, 32'h42a18ead, 32'h41705ee1, 32'h41a477a4, 32'h0};
test_input[14648:14655] = '{32'hc2c7c7f5, 32'hc278d1de, 32'hc2ba4519, 32'h42a5ab7b, 32'hc254a007, 32'h4263ea3e, 32'hc1e488c1, 32'h4190eed9};
test_output[14648:14655] = '{32'h0, 32'h0, 32'h0, 32'h42a5ab7b, 32'h0, 32'h4263ea3e, 32'h0, 32'h4190eed9};
test_input[14656:14663] = '{32'hc2bc1f4e, 32'h41158cfd, 32'hc2223884, 32'h41c62a97, 32'h422cbd54, 32'h422db0f3, 32'h42a2f55b, 32'hc2738c64};
test_output[14656:14663] = '{32'h0, 32'h41158cfd, 32'h0, 32'h41c62a97, 32'h422cbd54, 32'h422db0f3, 32'h42a2f55b, 32'h0};
test_input[14664:14671] = '{32'h42576c30, 32'hc2c14ebd, 32'h42a18656, 32'hc21e2794, 32'hc1f956f0, 32'hc290d4cf, 32'h420b00e9, 32'hc27eda97};
test_output[14664:14671] = '{32'h42576c30, 32'h0, 32'h42a18656, 32'h0, 32'h0, 32'h0, 32'h420b00e9, 32'h0};
test_input[14672:14679] = '{32'hc2659f1f, 32'hc23bc899, 32'hc156fb9f, 32'h3f945052, 32'hc1943f97, 32'h4249986d, 32'hc2c72a34, 32'h3ef99ce0};
test_output[14672:14679] = '{32'h0, 32'h0, 32'h0, 32'h3f945052, 32'h0, 32'h4249986d, 32'h0, 32'h3ef99ce0};
test_input[14680:14687] = '{32'h42a69b0b, 32'hc22f6307, 32'h421cc133, 32'hc23c30d5, 32'h42c22814, 32'h42c26774, 32'h42377233, 32'h424b1143};
test_output[14680:14687] = '{32'h42a69b0b, 32'h0, 32'h421cc133, 32'h0, 32'h42c22814, 32'h42c26774, 32'h42377233, 32'h424b1143};
test_input[14688:14695] = '{32'hc28e56b0, 32'hc1bfdd26, 32'hc1cef328, 32'h41a115bf, 32'hc29e6204, 32'h41c63890, 32'h42c1bf6c, 32'hc2aa9e2a};
test_output[14688:14695] = '{32'h0, 32'h0, 32'h0, 32'h41a115bf, 32'h0, 32'h41c63890, 32'h42c1bf6c, 32'h0};
test_input[14696:14703] = '{32'hc2a6fc65, 32'hc25bee47, 32'h40b7e000, 32'h4031fd48, 32'h4249e21a, 32'hc287cd03, 32'h415bcc5e, 32'hc22c616f};
test_output[14696:14703] = '{32'h0, 32'h0, 32'h40b7e000, 32'h4031fd48, 32'h4249e21a, 32'h0, 32'h415bcc5e, 32'h0};
test_input[14704:14711] = '{32'hc0ce1952, 32'hc2400dfd, 32'hc2a5f0f9, 32'hc29ef766, 32'h420bd2bf, 32'h4249d786, 32'hc1360fe9, 32'hc205f2d5};
test_output[14704:14711] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h420bd2bf, 32'h4249d786, 32'h0, 32'h0};
test_input[14712:14719] = '{32'hc281826e, 32'h4289b4e4, 32'h417e5222, 32'h4106a194, 32'h4049ee2e, 32'h4242fd29, 32'hc20867a7, 32'h41383e43};
test_output[14712:14719] = '{32'h0, 32'h4289b4e4, 32'h417e5222, 32'h4106a194, 32'h4049ee2e, 32'h4242fd29, 32'h0, 32'h41383e43};
test_input[14720:14727] = '{32'hc15a5246, 32'h4222eafb, 32'hbf67d622, 32'h4164a117, 32'hc1866309, 32'h427e58e6, 32'h40d8d217, 32'hc264bf49};
test_output[14720:14727] = '{32'h0, 32'h4222eafb, 32'h0, 32'h4164a117, 32'h0, 32'h427e58e6, 32'h40d8d217, 32'h0};
test_input[14728:14735] = '{32'hc2a7ca44, 32'h42a3f5ba, 32'h40337f69, 32'h42a0bba7, 32'hc2939845, 32'hc10c7bc8, 32'h41dea667, 32'hc2b1e2b1};
test_output[14728:14735] = '{32'h0, 32'h42a3f5ba, 32'h40337f69, 32'h42a0bba7, 32'h0, 32'h0, 32'h41dea667, 32'h0};
test_input[14736:14743] = '{32'h42b401e4, 32'h41f26634, 32'h41b0b931, 32'hc22ebd5f, 32'hc2bd1569, 32'hc211f3d5, 32'h419d4d62, 32'hc2a6be9b};
test_output[14736:14743] = '{32'h42b401e4, 32'h41f26634, 32'h41b0b931, 32'h0, 32'h0, 32'h0, 32'h419d4d62, 32'h0};
test_input[14744:14751] = '{32'hc2bc82d7, 32'h42c4aa24, 32'h4131552f, 32'h42545f55, 32'h429ce5a4, 32'h42931613, 32'hc2634cb0, 32'h42a14ae8};
test_output[14744:14751] = '{32'h0, 32'h42c4aa24, 32'h4131552f, 32'h42545f55, 32'h429ce5a4, 32'h42931613, 32'h0, 32'h42a14ae8};
test_input[14752:14759] = '{32'hc2bd1e8d, 32'h40a540b5, 32'h4202993d, 32'h423cdffe, 32'h4283b00e, 32'hc295910f, 32'hc2172494, 32'hc2ba4a33};
test_output[14752:14759] = '{32'h0, 32'h40a540b5, 32'h4202993d, 32'h423cdffe, 32'h4283b00e, 32'h0, 32'h0, 32'h0};
test_input[14760:14767] = '{32'h428e119f, 32'hc2a76c54, 32'h41da7bad, 32'hc20fedcc, 32'hc20a2546, 32'hc2208780, 32'h42b7ee6e, 32'h42b33826};
test_output[14760:14767] = '{32'h428e119f, 32'h0, 32'h41da7bad, 32'h0, 32'h0, 32'h0, 32'h42b7ee6e, 32'h42b33826};
test_input[14768:14775] = '{32'h42a969fd, 32'hc2a34df2, 32'h411033b6, 32'h42b4c679, 32'h41494788, 32'hc281150b, 32'h41a46ae8, 32'h42220d21};
test_output[14768:14775] = '{32'h42a969fd, 32'h0, 32'h411033b6, 32'h42b4c679, 32'h41494788, 32'h0, 32'h41a46ae8, 32'h42220d21};
test_input[14776:14783] = '{32'h42ae4311, 32'hc2bb48cb, 32'h429dd07f, 32'h428a3387, 32'hc219ea71, 32'h4294068a, 32'hc2ab6f2f, 32'h42460e53};
test_output[14776:14783] = '{32'h42ae4311, 32'h0, 32'h429dd07f, 32'h428a3387, 32'h0, 32'h4294068a, 32'h0, 32'h42460e53};
test_input[14784:14791] = '{32'h42aa3cdb, 32'hc284fc54, 32'h427af7de, 32'h42b10e16, 32'hc261d35d, 32'h40177317, 32'h42a2daaa, 32'h42945e08};
test_output[14784:14791] = '{32'h42aa3cdb, 32'h0, 32'h427af7de, 32'h42b10e16, 32'h0, 32'h40177317, 32'h42a2daaa, 32'h42945e08};
test_input[14792:14799] = '{32'hc1d7dbe1, 32'hc2bd5bbe, 32'hc2bef341, 32'h425027fe, 32'hc246fc71, 32'hc26fe0c8, 32'h41c6f94e, 32'h428b6ccb};
test_output[14792:14799] = '{32'h0, 32'h0, 32'h0, 32'h425027fe, 32'h0, 32'h0, 32'h41c6f94e, 32'h428b6ccb};
test_input[14800:14807] = '{32'hc25d99c5, 32'hc29904e2, 32'h41ce4891, 32'h427a56f9, 32'hc200bb8a, 32'h414f6e1e, 32'hc0fd7a12, 32'hc19c26f5};
test_output[14800:14807] = '{32'h0, 32'h0, 32'h41ce4891, 32'h427a56f9, 32'h0, 32'h414f6e1e, 32'h0, 32'h0};
test_input[14808:14815] = '{32'hbfbf3df7, 32'h42696bbc, 32'h42c2af2f, 32'h42b6a76d, 32'hc2136bc4, 32'h42928fcd, 32'hc27199f5, 32'h4233591e};
test_output[14808:14815] = '{32'h0, 32'h42696bbc, 32'h42c2af2f, 32'h42b6a76d, 32'h0, 32'h42928fcd, 32'h0, 32'h4233591e};
test_input[14816:14823] = '{32'hc2583e68, 32'hc250043b, 32'h4243345b, 32'h414af860, 32'hc20704a4, 32'h4190716b, 32'h4124d210, 32'h4269d3fb};
test_output[14816:14823] = '{32'h0, 32'h0, 32'h4243345b, 32'h414af860, 32'h0, 32'h4190716b, 32'h4124d210, 32'h4269d3fb};
test_input[14824:14831] = '{32'hc28cd2e3, 32'hc250a695, 32'h429df59c, 32'h428adb72, 32'hc19d10ff, 32'hc28d105f, 32'hc2b8c080, 32'h42009ffe};
test_output[14824:14831] = '{32'h0, 32'h0, 32'h429df59c, 32'h428adb72, 32'h0, 32'h0, 32'h0, 32'h42009ffe};
test_input[14832:14839] = '{32'hc16ce06e, 32'h4278c717, 32'hc2162aa4, 32'h4291d0c5, 32'hc2b7cf4a, 32'hc21d46f2, 32'hc1e695d1, 32'h41e57a80};
test_output[14832:14839] = '{32'h0, 32'h4278c717, 32'h0, 32'h4291d0c5, 32'h0, 32'h0, 32'h0, 32'h41e57a80};
test_input[14840:14847] = '{32'h427d55c5, 32'h425540a2, 32'h42c6dea7, 32'hc2a6bde1, 32'h42ab5a21, 32'h4184aa53, 32'hc269584c, 32'hc2b83427};
test_output[14840:14847] = '{32'h427d55c5, 32'h425540a2, 32'h42c6dea7, 32'h0, 32'h42ab5a21, 32'h4184aa53, 32'h0, 32'h0};
test_input[14848:14855] = '{32'h424df668, 32'h41baa76b, 32'h424ef1cb, 32'hc1bf9aee, 32'hc1242cfa, 32'h42556167, 32'hc138cf48, 32'h408591b2};
test_output[14848:14855] = '{32'h424df668, 32'h41baa76b, 32'h424ef1cb, 32'h0, 32'h0, 32'h42556167, 32'h0, 32'h408591b2};
test_input[14856:14863] = '{32'h421d4fde, 32'h41cb60f6, 32'hc1ed7783, 32'hc284a0c3, 32'h42927d5c, 32'hc2878e89, 32'hc1b19ef3, 32'hc2a240a0};
test_output[14856:14863] = '{32'h421d4fde, 32'h41cb60f6, 32'h0, 32'h0, 32'h42927d5c, 32'h0, 32'h0, 32'h0};
test_input[14864:14871] = '{32'hc2aaad02, 32'h42bb8b9a, 32'h428d52c4, 32'h425f5756, 32'hc2aea8be, 32'hc25c8155, 32'hc1a98c27, 32'hc154bbf9};
test_output[14864:14871] = '{32'h0, 32'h42bb8b9a, 32'h428d52c4, 32'h425f5756, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14872:14879] = '{32'h42b11dfe, 32'h426685ff, 32'h423d7c41, 32'h4037035c, 32'h42171092, 32'hc2aadf05, 32'hbe9faf45, 32'hc2244229};
test_output[14872:14879] = '{32'h42b11dfe, 32'h426685ff, 32'h423d7c41, 32'h4037035c, 32'h42171092, 32'h0, 32'h0, 32'h0};
test_input[14880:14887] = '{32'h42b46108, 32'h4291fa39, 32'hc1ab85f0, 32'hc23fe1ac, 32'h42188cfb, 32'h40b826ed, 32'h42a19d66, 32'h42b3759f};
test_output[14880:14887] = '{32'h42b46108, 32'h4291fa39, 32'h0, 32'h0, 32'h42188cfb, 32'h40b826ed, 32'h42a19d66, 32'h42b3759f};
test_input[14888:14895] = '{32'hc295693d, 32'h4293fb00, 32'h4269feba, 32'h42403920, 32'hc29834ea, 32'hc166ea8c, 32'hc2a803c2, 32'hc18b4e07};
test_output[14888:14895] = '{32'h0, 32'h4293fb00, 32'h4269feba, 32'h42403920, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14896:14903] = '{32'h425a17a7, 32'h42052f61, 32'hc119cc17, 32'h429cbde7, 32'h425d1223, 32'hc19f294e, 32'hc12969e5, 32'h4283bf49};
test_output[14896:14903] = '{32'h425a17a7, 32'h42052f61, 32'h0, 32'h429cbde7, 32'h425d1223, 32'h0, 32'h0, 32'h4283bf49};
test_input[14904:14911] = '{32'h424b685f, 32'h422a13b7, 32'h4140a623, 32'h428d9001, 32'h426cef5a, 32'hc16050b4, 32'h4284d8b2, 32'h427c7c81};
test_output[14904:14911] = '{32'h424b685f, 32'h422a13b7, 32'h4140a623, 32'h428d9001, 32'h426cef5a, 32'h0, 32'h4284d8b2, 32'h427c7c81};
test_input[14912:14919] = '{32'h42b89390, 32'hc191af2d, 32'hc2520ecd, 32'hc03f36aa, 32'hc2ab38f3, 32'h4216e6c0, 32'hc293fe26, 32'hc2abeea8};
test_output[14912:14919] = '{32'h42b89390, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4216e6c0, 32'h0, 32'h0};
test_input[14920:14927] = '{32'hc279dcf9, 32'h42920be0, 32'hc1477006, 32'h42beb9f3, 32'hc2a21b2b, 32'h4297398a, 32'hc286f1f4, 32'hc107707c};
test_output[14920:14927] = '{32'h0, 32'h42920be0, 32'h0, 32'h42beb9f3, 32'h0, 32'h4297398a, 32'h0, 32'h0};
test_input[14928:14935] = '{32'h41d7be77, 32'hc2c15901, 32'hc248a746, 32'h405b54e5, 32'h4247d690, 32'h42811173, 32'h41df0765, 32'hc25b8fea};
test_output[14928:14935] = '{32'h41d7be77, 32'h0, 32'h0, 32'h405b54e5, 32'h4247d690, 32'h42811173, 32'h41df0765, 32'h0};
test_input[14936:14943] = '{32'h4243a755, 32'h42c1bec1, 32'h42aa08d4, 32'hc2491e74, 32'h42a6eef9, 32'hc299a917, 32'h4248fa91, 32'h427b24b9};
test_output[14936:14943] = '{32'h4243a755, 32'h42c1bec1, 32'h42aa08d4, 32'h0, 32'h42a6eef9, 32'h0, 32'h4248fa91, 32'h427b24b9};
test_input[14944:14951] = '{32'h42bd679a, 32'hc0df4d85, 32'hc2056c76, 32'h422a8724, 32'h42c40555, 32'h425e7d41, 32'h429fdf2c, 32'hc22bf53b};
test_output[14944:14951] = '{32'h42bd679a, 32'h0, 32'h0, 32'h422a8724, 32'h42c40555, 32'h425e7d41, 32'h429fdf2c, 32'h0};
test_input[14952:14959] = '{32'h4281f33c, 32'h42aceba9, 32'h42843283, 32'hc1ff675a, 32'hc239e742, 32'hc2b70aee, 32'hc16babf2, 32'h3fc3d610};
test_output[14952:14959] = '{32'h4281f33c, 32'h42aceba9, 32'h42843283, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3fc3d610};
test_input[14960:14967] = '{32'h42a0ad79, 32'hc20944de, 32'hc26f4df6, 32'hc210b8a9, 32'h422d3982, 32'h412afd3c, 32'hc28ce6ed, 32'hc2817eee};
test_output[14960:14967] = '{32'h42a0ad79, 32'h0, 32'h0, 32'h0, 32'h422d3982, 32'h412afd3c, 32'h0, 32'h0};
test_input[14968:14975] = '{32'hc22ee1d9, 32'hc286db36, 32'h426add02, 32'h3fac88d4, 32'hc2b9cd83, 32'h4248e7cb, 32'hc0859b31, 32'hbe9137e6};
test_output[14968:14975] = '{32'h0, 32'h0, 32'h426add02, 32'h3fac88d4, 32'h0, 32'h4248e7cb, 32'h0, 32'h0};
test_input[14976:14983] = '{32'h41cfb7cc, 32'hc2341092, 32'h425f4a2b, 32'h42881e10, 32'hc202196c, 32'h41db6e53, 32'h42ab97c2, 32'hc2bc8d7e};
test_output[14976:14983] = '{32'h41cfb7cc, 32'h0, 32'h425f4a2b, 32'h42881e10, 32'h0, 32'h41db6e53, 32'h42ab97c2, 32'h0};
test_input[14984:14991] = '{32'h425e5368, 32'hc2baf306, 32'hc20d70dd, 32'h42a532c5, 32'hc0016f2d, 32'hbf781ad3, 32'hc28f65f7, 32'hc2a5df00};
test_output[14984:14991] = '{32'h425e5368, 32'h0, 32'h0, 32'h42a532c5, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[14992:14999] = '{32'h4223539f, 32'h421a89bf, 32'hc2bf769d, 32'hc27bb277, 32'h42248a0c, 32'h3f4eb79a, 32'hc1a70cea, 32'h4276ed81};
test_output[14992:14999] = '{32'h4223539f, 32'h421a89bf, 32'h0, 32'h0, 32'h42248a0c, 32'h3f4eb79a, 32'h0, 32'h4276ed81};
test_input[15000:15007] = '{32'h42a9b71e, 32'h413e80ab, 32'h4223a974, 32'h42c74ee8, 32'hc244d536, 32'h4284a6af, 32'h42c0d6f3, 32'hc1dfd364};
test_output[15000:15007] = '{32'h42a9b71e, 32'h413e80ab, 32'h4223a974, 32'h42c74ee8, 32'h0, 32'h4284a6af, 32'h42c0d6f3, 32'h0};
test_input[15008:15015] = '{32'hc2857366, 32'hc2054cf6, 32'hc1bb3cf8, 32'h415dd77c, 32'h421e1d49, 32'hc0d68258, 32'h42694f0f, 32'hc20a04a5};
test_output[15008:15015] = '{32'h0, 32'h0, 32'h0, 32'h415dd77c, 32'h421e1d49, 32'h0, 32'h42694f0f, 32'h0};
test_input[15016:15023] = '{32'h4264bf96, 32'h42ad610f, 32'hc10b6980, 32'h40b677ae, 32'hc2b558b1, 32'h429566fe, 32'hc1a1c4f0, 32'hc246de90};
test_output[15016:15023] = '{32'h4264bf96, 32'h42ad610f, 32'h0, 32'h40b677ae, 32'h0, 32'h429566fe, 32'h0, 32'h0};
test_input[15024:15031] = '{32'h41e945ca, 32'h42115722, 32'h42400da3, 32'hc259c0c9, 32'hc187a857, 32'hc22e9425, 32'h428d4885, 32'h425480cb};
test_output[15024:15031] = '{32'h41e945ca, 32'h42115722, 32'h42400da3, 32'h0, 32'h0, 32'h0, 32'h428d4885, 32'h425480cb};
test_input[15032:15039] = '{32'h423b3707, 32'h425ae8d0, 32'hc2747dbf, 32'h3fbcc613, 32'hc24bb96b, 32'h4156b8f1, 32'hc2568082, 32'h42325a13};
test_output[15032:15039] = '{32'h423b3707, 32'h425ae8d0, 32'h0, 32'h3fbcc613, 32'h0, 32'h4156b8f1, 32'h0, 32'h42325a13};
test_input[15040:15047] = '{32'hc22716b4, 32'h41f78488, 32'h41bff7ef, 32'h427489e2, 32'h419b9229, 32'h4232f324, 32'hc298377f, 32'hc24adb81};
test_output[15040:15047] = '{32'h0, 32'h41f78488, 32'h41bff7ef, 32'h427489e2, 32'h419b9229, 32'h4232f324, 32'h0, 32'h0};
test_input[15048:15055] = '{32'h41b6cf24, 32'hc29739ec, 32'hc21e5bbb, 32'hc2ab8658, 32'hc277de10, 32'hc2bd354d, 32'h423fd98c, 32'hc2121f0c};
test_output[15048:15055] = '{32'h41b6cf24, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423fd98c, 32'h0};
test_input[15056:15063] = '{32'h40f39f91, 32'h428378a4, 32'h424bcb5a, 32'h41db7b2c, 32'hc1dbc784, 32'hc14614bf, 32'h42409921, 32'h4286f201};
test_output[15056:15063] = '{32'h40f39f91, 32'h428378a4, 32'h424bcb5a, 32'h41db7b2c, 32'h0, 32'h0, 32'h42409921, 32'h4286f201};
test_input[15064:15071] = '{32'hc03f946c, 32'hc2c3ab32, 32'h40b31873, 32'hc28646df, 32'h40a4a6a6, 32'h406ab36e, 32'hc0f81cf5, 32'hc2a38366};
test_output[15064:15071] = '{32'h0, 32'h0, 32'h40b31873, 32'h0, 32'h40a4a6a6, 32'h406ab36e, 32'h0, 32'h0};
test_input[15072:15079] = '{32'hc2bbe4f4, 32'h424fb0d2, 32'hc2371d8c, 32'hc2a696f4, 32'h428ab497, 32'h417886ed, 32'hc1bddc42, 32'h41a32613};
test_output[15072:15079] = '{32'h0, 32'h424fb0d2, 32'h0, 32'h0, 32'h428ab497, 32'h417886ed, 32'h0, 32'h41a32613};
test_input[15080:15087] = '{32'hc2be59a2, 32'h40c530cd, 32'hc0e376d0, 32'hc11bc0ef, 32'h417f7044, 32'h4280948c, 32'h42c1d3e8, 32'h41f25f1d};
test_output[15080:15087] = '{32'h0, 32'h40c530cd, 32'h0, 32'h0, 32'h417f7044, 32'h4280948c, 32'h42c1d3e8, 32'h41f25f1d};
test_input[15088:15095] = '{32'h42af6a45, 32'h42379509, 32'hc1ffe4e0, 32'h417f12c8, 32'h41d96b9b, 32'h42b0ece6, 32'hc22fa05d, 32'h4035fd9d};
test_output[15088:15095] = '{32'h42af6a45, 32'h42379509, 32'h0, 32'h417f12c8, 32'h41d96b9b, 32'h42b0ece6, 32'h0, 32'h4035fd9d};
test_input[15096:15103] = '{32'h42b4546d, 32'h429be230, 32'hc243fc8e, 32'h42611981, 32'h42a477d1, 32'h41bb4ea8, 32'hc18c65f4, 32'h429b9c93};
test_output[15096:15103] = '{32'h42b4546d, 32'h429be230, 32'h0, 32'h42611981, 32'h42a477d1, 32'h41bb4ea8, 32'h0, 32'h429b9c93};
test_input[15104:15111] = '{32'h41e287b6, 32'hc26da4c9, 32'h41ce0abc, 32'hc2177fb8, 32'h428ced38, 32'hc27fe23a, 32'hc1e9fb8a, 32'hc29f43a7};
test_output[15104:15111] = '{32'h41e287b6, 32'h0, 32'h41ce0abc, 32'h0, 32'h428ced38, 32'h0, 32'h0, 32'h0};
test_input[15112:15119] = '{32'hc29bd15d, 32'h4282c871, 32'h4269fde2, 32'h4121a44a, 32'h42243fee, 32'h426a9319, 32'h413d7b7b, 32'h42c1d9b9};
test_output[15112:15119] = '{32'h0, 32'h4282c871, 32'h4269fde2, 32'h4121a44a, 32'h42243fee, 32'h426a9319, 32'h413d7b7b, 32'h42c1d9b9};
test_input[15120:15127] = '{32'hc2b40e56, 32'hc266c09b, 32'hc259ae88, 32'hc03808d6, 32'hc26566a3, 32'h426dcd53, 32'hc29a9e04, 32'hc28ec499};
test_output[15120:15127] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426dcd53, 32'h0, 32'h0};
test_input[15128:15135] = '{32'h41a98f90, 32'hc19bcb74, 32'h4284cc2e, 32'h428892ad, 32'hc2c43605, 32'hc296b49f, 32'hc28d0ea2, 32'hc2914bc8};
test_output[15128:15135] = '{32'h41a98f90, 32'h0, 32'h4284cc2e, 32'h428892ad, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15136:15143] = '{32'hc2c42eda, 32'h41d36555, 32'hc1d66a09, 32'h4122046f, 32'h427cc28a, 32'h42092a52, 32'hc21e5a12, 32'hc267e61d};
test_output[15136:15143] = '{32'h0, 32'h41d36555, 32'h0, 32'h4122046f, 32'h427cc28a, 32'h42092a52, 32'h0, 32'h0};
test_input[15144:15151] = '{32'hbfa34a56, 32'h42989d4a, 32'h3ee9085b, 32'hc111a80c, 32'hc28f67b3, 32'h42959fb1, 32'hc29ff2f7, 32'h42b44e96};
test_output[15144:15151] = '{32'h0, 32'h42989d4a, 32'h3ee9085b, 32'h0, 32'h0, 32'h42959fb1, 32'h0, 32'h42b44e96};
test_input[15152:15159] = '{32'hc23533cb, 32'hc1fd5175, 32'h41ee9934, 32'h425f565c, 32'hc2493f28, 32'hc2526910, 32'h422b127f, 32'h42b2720b};
test_output[15152:15159] = '{32'h0, 32'h0, 32'h41ee9934, 32'h425f565c, 32'h0, 32'h0, 32'h422b127f, 32'h42b2720b};
test_input[15160:15167] = '{32'h42850d7d, 32'hc27b1363, 32'h420df201, 32'h42489c73, 32'hc2abe426, 32'h41ff2ee4, 32'h426bc19f, 32'hc2b18ea3};
test_output[15160:15167] = '{32'h42850d7d, 32'h0, 32'h420df201, 32'h42489c73, 32'h0, 32'h41ff2ee4, 32'h426bc19f, 32'h0};
test_input[15168:15175] = '{32'hc2b37301, 32'h40cdc83d, 32'hc20e07b5, 32'hc2701d8e, 32'hc2516e20, 32'hc23d2403, 32'h415a040d, 32'hc2ba3513};
test_output[15168:15175] = '{32'h0, 32'h40cdc83d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h415a040d, 32'h0};
test_input[15176:15183] = '{32'h42b32838, 32'hc19eaf6a, 32'hc1df6a4b, 32'h41d912d8, 32'hc2070e06, 32'h418d2e8d, 32'h4294da1f, 32'hc2526be9};
test_output[15176:15183] = '{32'h42b32838, 32'h0, 32'h0, 32'h41d912d8, 32'h0, 32'h418d2e8d, 32'h4294da1f, 32'h0};
test_input[15184:15191] = '{32'hc217a9ef, 32'hc052ce5e, 32'hc1cad0cb, 32'h42a89722, 32'h42aea03d, 32'hc277770d, 32'h4180773b, 32'hc0ae51d8};
test_output[15184:15191] = '{32'h0, 32'h0, 32'h0, 32'h42a89722, 32'h42aea03d, 32'h0, 32'h4180773b, 32'h0};
test_input[15192:15199] = '{32'hc25cfe1b, 32'hc1f3ab4a, 32'h42ada56d, 32'hc269849b, 32'h41c249af, 32'h4134d16f, 32'h422fd40a, 32'h4236368f};
test_output[15192:15199] = '{32'h0, 32'h0, 32'h42ada56d, 32'h0, 32'h41c249af, 32'h4134d16f, 32'h422fd40a, 32'h4236368f};
test_input[15200:15207] = '{32'hc2b3c981, 32'hc2a802c8, 32'hc2bd57c9, 32'h421091d4, 32'hc1df1748, 32'hc1e57db5, 32'h4256d4b5, 32'h4274eee2};
test_output[15200:15207] = '{32'h0, 32'h0, 32'h0, 32'h421091d4, 32'h0, 32'h0, 32'h4256d4b5, 32'h4274eee2};
test_input[15208:15215] = '{32'h423ac12c, 32'h406aa275, 32'hc2be093c, 32'h42240041, 32'h40ecd982, 32'h40ef049f, 32'hc18d7bef, 32'hc23edd96};
test_output[15208:15215] = '{32'h423ac12c, 32'h406aa275, 32'h0, 32'h42240041, 32'h40ecd982, 32'h40ef049f, 32'h0, 32'h0};
test_input[15216:15223] = '{32'h425b8bbe, 32'hc2c28310, 32'h42a794b5, 32'h4074d370, 32'h429b40be, 32'hc1bdfa24, 32'h40a2869c, 32'h41edc84a};
test_output[15216:15223] = '{32'h425b8bbe, 32'h0, 32'h42a794b5, 32'h4074d370, 32'h429b40be, 32'h0, 32'h40a2869c, 32'h41edc84a};
test_input[15224:15231] = '{32'hc2a44127, 32'h42b04cad, 32'h422a77fc, 32'hc200070d, 32'hc2c2a08d, 32'h40ef6969, 32'hc20a42c2, 32'hc120e311};
test_output[15224:15231] = '{32'h0, 32'h42b04cad, 32'h422a77fc, 32'h0, 32'h0, 32'h40ef6969, 32'h0, 32'h0};
test_input[15232:15239] = '{32'hc219cb6d, 32'hc29384b8, 32'hc13e2ab3, 32'h422a702b, 32'hc095bd06, 32'hc241f593, 32'h4192f64f, 32'hc2841bfe};
test_output[15232:15239] = '{32'h0, 32'h0, 32'h0, 32'h422a702b, 32'h0, 32'h0, 32'h4192f64f, 32'h0};
test_input[15240:15247] = '{32'hc2abaff7, 32'h42794800, 32'hc293cf76, 32'hc28a48c8, 32'h3f57d1c2, 32'hc0919184, 32'hc0ed1e3b, 32'hc1e0f7b6};
test_output[15240:15247] = '{32'h0, 32'h42794800, 32'h0, 32'h0, 32'h3f57d1c2, 32'h0, 32'h0, 32'h0};
test_input[15248:15255] = '{32'hc2070b62, 32'hc2ac5f13, 32'hc279bca1, 32'h3e67c729, 32'h42155c79, 32'h426c6bba, 32'hc1fb0bb4, 32'h426e179d};
test_output[15248:15255] = '{32'h0, 32'h0, 32'h0, 32'h3e67c729, 32'h42155c79, 32'h426c6bba, 32'h0, 32'h426e179d};
test_input[15256:15263] = '{32'hc24a4727, 32'h42336fd1, 32'hc2a5f3d9, 32'hbf5ce19f, 32'hc229c8e3, 32'hc1ce21fc, 32'hc28cfdf3, 32'hc20c7108};
test_output[15256:15263] = '{32'h0, 32'h42336fd1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15264:15271] = '{32'hbef284fd, 32'hc2aa4b79, 32'h42b4c095, 32'hc01d3bde, 32'h41f2e3ad, 32'hc248f9af, 32'h401541d3, 32'hc217cb72};
test_output[15264:15271] = '{32'h0, 32'h0, 32'h42b4c095, 32'h0, 32'h41f2e3ad, 32'h0, 32'h401541d3, 32'h0};
test_input[15272:15279] = '{32'h42970a56, 32'hc2c693b0, 32'hc2c03bb9, 32'hc215c6e3, 32'h42976e7c, 32'hc15e0e00, 32'hc2c040ec, 32'h42a15fbe};
test_output[15272:15279] = '{32'h42970a56, 32'h0, 32'h0, 32'h0, 32'h42976e7c, 32'h0, 32'h0, 32'h42a15fbe};
test_input[15280:15287] = '{32'h426cf000, 32'h427fd3e3, 32'hc2341d00, 32'h42a7fae5, 32'h422784ec, 32'hc2696a21, 32'h41711ac0, 32'h42914699};
test_output[15280:15287] = '{32'h426cf000, 32'h427fd3e3, 32'h0, 32'h42a7fae5, 32'h422784ec, 32'h0, 32'h41711ac0, 32'h42914699};
test_input[15288:15295] = '{32'h42389436, 32'h42372676, 32'hc10366ea, 32'h3f47fe56, 32'h425b80a2, 32'hc212aaa2, 32'h42974ba0, 32'hc225470c};
test_output[15288:15295] = '{32'h42389436, 32'h42372676, 32'h0, 32'h3f47fe56, 32'h425b80a2, 32'h0, 32'h42974ba0, 32'h0};
test_input[15296:15303] = '{32'hc1d745e1, 32'h41fcdab4, 32'h42c12f61, 32'hc2b98d75, 32'hc220e022, 32'h40e9b50a, 32'h424b4df1, 32'h4298f8b6};
test_output[15296:15303] = '{32'h0, 32'h41fcdab4, 32'h42c12f61, 32'h0, 32'h0, 32'h40e9b50a, 32'h424b4df1, 32'h4298f8b6};
test_input[15304:15311] = '{32'hc1a7abd3, 32'h41bf1523, 32'hc29fcc3c, 32'hc1823b49, 32'h42aeab8a, 32'hc1a13e9d, 32'hc27a7934, 32'hc11ad43e};
test_output[15304:15311] = '{32'h0, 32'h41bf1523, 32'h0, 32'h0, 32'h42aeab8a, 32'h0, 32'h0, 32'h0};
test_input[15312:15319] = '{32'h428db261, 32'h4220c25f, 32'h4299ed43, 32'hc2b42b5f, 32'hc29baed1, 32'hc1903bf9, 32'hc22c517c, 32'h41f3de16};
test_output[15312:15319] = '{32'h428db261, 32'h4220c25f, 32'h4299ed43, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f3de16};
test_input[15320:15327] = '{32'hc2bda57a, 32'hc113ec2a, 32'h4293301a, 32'hc173e22f, 32'hc1eeeb8e, 32'hc0f929e0, 32'h42350a63, 32'hc2936945};
test_output[15320:15327] = '{32'h0, 32'h0, 32'h4293301a, 32'h0, 32'h0, 32'h0, 32'h42350a63, 32'h0};
test_input[15328:15335] = '{32'hc05631b9, 32'h41de5847, 32'h42baa0fa, 32'hc216f6d3, 32'hc2124760, 32'h42a45d51, 32'hc21e21ae, 32'hc241668f};
test_output[15328:15335] = '{32'h0, 32'h41de5847, 32'h42baa0fa, 32'h0, 32'h0, 32'h42a45d51, 32'h0, 32'h0};
test_input[15336:15343] = '{32'h42353520, 32'h42c2ac3a, 32'hc234d6e8, 32'hc1ddbfa7, 32'h4203fe94, 32'h415ba404, 32'h42b5fc29, 32'h42be1f55};
test_output[15336:15343] = '{32'h42353520, 32'h42c2ac3a, 32'h0, 32'h0, 32'h4203fe94, 32'h415ba404, 32'h42b5fc29, 32'h42be1f55};
test_input[15344:15351] = '{32'h4215c11b, 32'h4283a53e, 32'hc1eb78e3, 32'hc23c27f0, 32'h42c4070b, 32'h420b4f32, 32'hc25a39f8, 32'hc298b3d9};
test_output[15344:15351] = '{32'h4215c11b, 32'h4283a53e, 32'h0, 32'h0, 32'h42c4070b, 32'h420b4f32, 32'h0, 32'h0};
test_input[15352:15359] = '{32'hc1a433ca, 32'hc2b39ae2, 32'h4180cf5f, 32'h411d6244, 32'hc2c05431, 32'hc24b8639, 32'h41c830fa, 32'h419e045d};
test_output[15352:15359] = '{32'h0, 32'h0, 32'h4180cf5f, 32'h411d6244, 32'h0, 32'h0, 32'h41c830fa, 32'h419e045d};
test_input[15360:15367] = '{32'h3fe2cee7, 32'hc29dfadc, 32'hc21d9c90, 32'h40dc0e1d, 32'h41e87644, 32'h42c40a33, 32'hc1adf2a8, 32'hc2972ed2};
test_output[15360:15367] = '{32'h3fe2cee7, 32'h0, 32'h0, 32'h40dc0e1d, 32'h41e87644, 32'h42c40a33, 32'h0, 32'h0};
test_input[15368:15375] = '{32'h426224c4, 32'h41d7d27a, 32'hbf1b8da9, 32'hc08c23cc, 32'hc224f3ca, 32'h41e9ab26, 32'hc21d2079, 32'h42729724};
test_output[15368:15375] = '{32'h426224c4, 32'h41d7d27a, 32'h0, 32'h0, 32'h0, 32'h41e9ab26, 32'h0, 32'h42729724};
test_input[15376:15383] = '{32'hc2b56d7d, 32'h426609b0, 32'hc0b77492, 32'hc21986ed, 32'h42395a94, 32'hc23ceeeb, 32'h41e4a568, 32'hc26e3f6a};
test_output[15376:15383] = '{32'h0, 32'h426609b0, 32'h0, 32'h0, 32'h42395a94, 32'h0, 32'h41e4a568, 32'h0};
test_input[15384:15391] = '{32'hc213ae56, 32'hc23bbb5e, 32'hc2bcb88a, 32'h429b57fa, 32'h421b63bf, 32'hc242dab7, 32'hc175a1d9, 32'h4278a3c8};
test_output[15384:15391] = '{32'h0, 32'h0, 32'h0, 32'h429b57fa, 32'h421b63bf, 32'h0, 32'h0, 32'h4278a3c8};
test_input[15392:15399] = '{32'hc2c4017b, 32'hc1177f69, 32'h428e0cb3, 32'h412d74b8, 32'h41f35ea9, 32'hc2111e84, 32'hc13744cb, 32'hbe8f8bb0};
test_output[15392:15399] = '{32'h0, 32'h0, 32'h428e0cb3, 32'h412d74b8, 32'h41f35ea9, 32'h0, 32'h0, 32'h0};
test_input[15400:15407] = '{32'h42b14511, 32'hc2a9e362, 32'h421990bc, 32'h42a62f1c, 32'hc2972325, 32'hc1962f8b, 32'h4264079b, 32'hc1bde082};
test_output[15400:15407] = '{32'h42b14511, 32'h0, 32'h421990bc, 32'h42a62f1c, 32'h0, 32'h0, 32'h4264079b, 32'h0};
test_input[15408:15415] = '{32'h42377a3e, 32'hc176308e, 32'hc2c37082, 32'h423ea4fe, 32'h427ef1a3, 32'hc27b3ec2, 32'h41dfd959, 32'h42200163};
test_output[15408:15415] = '{32'h42377a3e, 32'h0, 32'h0, 32'h423ea4fe, 32'h427ef1a3, 32'h0, 32'h41dfd959, 32'h42200163};
test_input[15416:15423] = '{32'h429d74d6, 32'hc2255f85, 32'h411641c2, 32'hc2b531ce, 32'h428252df, 32'hc28f4010, 32'h42ac06ae, 32'h428c6f5c};
test_output[15416:15423] = '{32'h429d74d6, 32'h0, 32'h411641c2, 32'h0, 32'h428252df, 32'h0, 32'h42ac06ae, 32'h428c6f5c};
test_input[15424:15431] = '{32'h42bbdc68, 32'h41b35111, 32'h42aeb0bd, 32'hc1b92d02, 32'hc0d5d7af, 32'h426ef05f, 32'h4271b9d2, 32'h3faf87be};
test_output[15424:15431] = '{32'h42bbdc68, 32'h41b35111, 32'h42aeb0bd, 32'h0, 32'h0, 32'h426ef05f, 32'h4271b9d2, 32'h3faf87be};
test_input[15432:15439] = '{32'hc2c77d46, 32'hc1edb689, 32'hc28ebee4, 32'hc27d6aca, 32'hc2ba3bbf, 32'h42972ba7, 32'h42b357b1, 32'h425fc3d9};
test_output[15432:15439] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42972ba7, 32'h42b357b1, 32'h425fc3d9};
test_input[15440:15447] = '{32'hc21533b3, 32'hc29d66bb, 32'hc2101301, 32'h42b4e2f9, 32'h426d5949, 32'hc2aabbf5, 32'hc10df905, 32'hc2c66d81};
test_output[15440:15447] = '{32'h0, 32'h0, 32'h0, 32'h42b4e2f9, 32'h426d5949, 32'h0, 32'h0, 32'h0};
test_input[15448:15455] = '{32'hc2958533, 32'h4113583d, 32'h429ca98f, 32'h4058b4f1, 32'hc2050bee, 32'h413d01d3, 32'hc2c1f9ae, 32'hc2421ec6};
test_output[15448:15455] = '{32'h0, 32'h4113583d, 32'h429ca98f, 32'h4058b4f1, 32'h0, 32'h413d01d3, 32'h0, 32'h0};
test_input[15456:15463] = '{32'h429ea010, 32'hc156c915, 32'hc1f3344b, 32'hc111d01c, 32'h428f3e55, 32'hc293f4b7, 32'h4214eebf, 32'h428caa35};
test_output[15456:15463] = '{32'h429ea010, 32'h0, 32'h0, 32'h0, 32'h428f3e55, 32'h0, 32'h4214eebf, 32'h428caa35};
test_input[15464:15471] = '{32'h42433ed2, 32'h41bae369, 32'hc2314f9f, 32'hc1fc2177, 32'h4258a56d, 32'h42809d28, 32'hc116b923, 32'hc2a1425c};
test_output[15464:15471] = '{32'h42433ed2, 32'h41bae369, 32'h0, 32'h0, 32'h4258a56d, 32'h42809d28, 32'h0, 32'h0};
test_input[15472:15479] = '{32'h3f58a9fb, 32'hc2101cc8, 32'hc2419ebe, 32'h41f78262, 32'hc2679d09, 32'h425c72e5, 32'h4296674b, 32'h42440a16};
test_output[15472:15479] = '{32'h3f58a9fb, 32'h0, 32'h0, 32'h41f78262, 32'h0, 32'h425c72e5, 32'h4296674b, 32'h42440a16};
test_input[15480:15487] = '{32'h3eab3ece, 32'hc277c751, 32'hc0be5b7c, 32'h42231675, 32'h429fd262, 32'hc297249a, 32'h4233d74f, 32'h4243cf76};
test_output[15480:15487] = '{32'h3eab3ece, 32'h0, 32'h0, 32'h42231675, 32'h429fd262, 32'h0, 32'h4233d74f, 32'h4243cf76};
test_input[15488:15495] = '{32'h42735636, 32'hc19cb4a3, 32'h428d81c0, 32'h42868cf0, 32'hc070bda0, 32'hc0c3c66f, 32'h40a1a68c, 32'h429800a9};
test_output[15488:15495] = '{32'h42735636, 32'h0, 32'h428d81c0, 32'h42868cf0, 32'h0, 32'h0, 32'h40a1a68c, 32'h429800a9};
test_input[15496:15503] = '{32'hc29fcc6d, 32'hc2c4dc1b, 32'hc23a7a49, 32'h42a7c76d, 32'hc238a6a7, 32'hc151bd7e, 32'hc28d4d2b, 32'hc182659e};
test_output[15496:15503] = '{32'h0, 32'h0, 32'h0, 32'h42a7c76d, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15504:15511] = '{32'h428d6186, 32'hc26fad3a, 32'h42384502, 32'hc18f8517, 32'h42075630, 32'h42be8d54, 32'hc29cb7d7, 32'hc25da783};
test_output[15504:15511] = '{32'h428d6186, 32'h0, 32'h42384502, 32'h0, 32'h42075630, 32'h42be8d54, 32'h0, 32'h0};
test_input[15512:15519] = '{32'h40ce27f9, 32'h42168199, 32'hc286be51, 32'h429677ca, 32'hc18574ca, 32'h411e7082, 32'hc0a3d77a, 32'h4287e809};
test_output[15512:15519] = '{32'h40ce27f9, 32'h42168199, 32'h0, 32'h429677ca, 32'h0, 32'h411e7082, 32'h0, 32'h4287e809};
test_input[15520:15527] = '{32'h418f4af8, 32'hc25940d9, 32'hc2be1b2b, 32'h41ad7b39, 32'hc12c1e99, 32'hc1208dd1, 32'h42a26566, 32'h4209fdb1};
test_output[15520:15527] = '{32'h418f4af8, 32'h0, 32'h0, 32'h41ad7b39, 32'h0, 32'h0, 32'h42a26566, 32'h4209fdb1};
test_input[15528:15535] = '{32'h413f27a0, 32'hc240f2ed, 32'h42312d7d, 32'hc2837a1c, 32'hc252eb35, 32'hc2b96284, 32'hc1937125, 32'hc1f6fe66};
test_output[15528:15535] = '{32'h413f27a0, 32'h0, 32'h42312d7d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15536:15543] = '{32'hc1f4a4ed, 32'hc22e706c, 32'hc0937792, 32'h4193a7a4, 32'h42732f9d, 32'hc22fc98f, 32'h42ad5f49, 32'h4238918c};
test_output[15536:15543] = '{32'h0, 32'h0, 32'h0, 32'h4193a7a4, 32'h42732f9d, 32'h0, 32'h42ad5f49, 32'h4238918c};
test_input[15544:15551] = '{32'hc1a1cb65, 32'h40dad5f0, 32'h41bec9b7, 32'h422fa2cd, 32'hc248c202, 32'h428ce515, 32'hc00f4d23, 32'h41d3386a};
test_output[15544:15551] = '{32'h0, 32'h40dad5f0, 32'h41bec9b7, 32'h422fa2cd, 32'h0, 32'h428ce515, 32'h0, 32'h41d3386a};
test_input[15552:15559] = '{32'hc2840f0c, 32'h42bdc62a, 32'hc20cda8f, 32'h412467c9, 32'hc1943eb7, 32'h41fcd6c0, 32'h42764858, 32'h424c6628};
test_output[15552:15559] = '{32'h0, 32'h42bdc62a, 32'h0, 32'h412467c9, 32'h0, 32'h41fcd6c0, 32'h42764858, 32'h424c6628};
test_input[15560:15567] = '{32'hc2416167, 32'h42aca592, 32'h423bbcb5, 32'h427de2bd, 32'h4112c59e, 32'hc02a5f7a, 32'h4214f7b7, 32'h425a95c1};
test_output[15560:15567] = '{32'h0, 32'h42aca592, 32'h423bbcb5, 32'h427de2bd, 32'h4112c59e, 32'h0, 32'h4214f7b7, 32'h425a95c1};
test_input[15568:15575] = '{32'h423f3ab0, 32'hc23674f7, 32'h42509b42, 32'h424815ee, 32'h41abcd48, 32'h427427bc, 32'hc232da9e, 32'h42a1f615};
test_output[15568:15575] = '{32'h423f3ab0, 32'h0, 32'h42509b42, 32'h424815ee, 32'h41abcd48, 32'h427427bc, 32'h0, 32'h42a1f615};
test_input[15576:15583] = '{32'hc292b6f4, 32'hc253ed83, 32'h41c5f3d4, 32'h41e342c2, 32'hc2acb588, 32'hc2312de4, 32'hc1ba7a48, 32'hc2369c5d};
test_output[15576:15583] = '{32'h0, 32'h0, 32'h41c5f3d4, 32'h41e342c2, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15584:15591] = '{32'hc2ba94a3, 32'h42a29145, 32'h41de5342, 32'h4288d385, 32'h41871f29, 32'hc1a06cab, 32'h42b8c744, 32'hc2bc48d4};
test_output[15584:15591] = '{32'h0, 32'h42a29145, 32'h41de5342, 32'h4288d385, 32'h41871f29, 32'h0, 32'h42b8c744, 32'h0};
test_input[15592:15599] = '{32'h42b6c313, 32'h416d8be7, 32'h4290a420, 32'h42b8d838, 32'hc2aa07eb, 32'h42bd149e, 32'hc2516c1b, 32'hc22afb15};
test_output[15592:15599] = '{32'h42b6c313, 32'h416d8be7, 32'h4290a420, 32'h42b8d838, 32'h0, 32'h42bd149e, 32'h0, 32'h0};
test_input[15600:15607] = '{32'hc2133094, 32'h41715493, 32'hc27d5df9, 32'hc2170390, 32'hc1ab2b65, 32'hc2967698, 32'h420e2f6c, 32'h42c21a04};
test_output[15600:15607] = '{32'h0, 32'h41715493, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420e2f6c, 32'h42c21a04};
test_input[15608:15615] = '{32'h42726c0c, 32'h42104687, 32'h42a24952, 32'h4207dfb7, 32'hc0ce9aa9, 32'hc199de57, 32'hc1b5200e, 32'hc1fb8afb};
test_output[15608:15615] = '{32'h42726c0c, 32'h42104687, 32'h42a24952, 32'h4207dfb7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15616:15623] = '{32'hc2b491f8, 32'hc1be49c0, 32'hc15f4a3d, 32'h41fb2455, 32'h422d1e38, 32'hbede4f3c, 32'h423cb612, 32'h427c5abc};
test_output[15616:15623] = '{32'h0, 32'h0, 32'h0, 32'h41fb2455, 32'h422d1e38, 32'h0, 32'h423cb612, 32'h427c5abc};
test_input[15624:15631] = '{32'h42b5241a, 32'h40ec6d17, 32'h412252bc, 32'hc2521b4c, 32'h4192ed0e, 32'hc2624975, 32'h41d71b4f, 32'hc1b455e7};
test_output[15624:15631] = '{32'h42b5241a, 32'h40ec6d17, 32'h412252bc, 32'h0, 32'h4192ed0e, 32'h0, 32'h41d71b4f, 32'h0};
test_input[15632:15639] = '{32'h41e09c28, 32'hc228a5ab, 32'hc2170e71, 32'hc288dbf8, 32'h42a6258f, 32'h41016cdf, 32'hc2823cf0, 32'h417b659a};
test_output[15632:15639] = '{32'h41e09c28, 32'h0, 32'h0, 32'h0, 32'h42a6258f, 32'h41016cdf, 32'h0, 32'h417b659a};
test_input[15640:15647] = '{32'hc2b7b6a5, 32'hc21732ad, 32'hc1cc5b39, 32'hc2bc3b52, 32'h4241a3e3, 32'h429307b4, 32'h41425a2e, 32'h41f03c66};
test_output[15640:15647] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4241a3e3, 32'h429307b4, 32'h41425a2e, 32'h41f03c66};
test_input[15648:15655] = '{32'hc0052888, 32'h42227e81, 32'h4132ea3c, 32'h4282f609, 32'hc28a0824, 32'hc2b3a543, 32'hc2a99ec8, 32'hc24f86c2};
test_output[15648:15655] = '{32'h0, 32'h42227e81, 32'h4132ea3c, 32'h4282f609, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15656:15663] = '{32'hc1028476, 32'hc29262e4, 32'hc2b6430d, 32'h41b8db4e, 32'h4218d6da, 32'hc2a96293, 32'hc1d4c219, 32'h41f76620};
test_output[15656:15663] = '{32'h0, 32'h0, 32'h0, 32'h41b8db4e, 32'h4218d6da, 32'h0, 32'h0, 32'h41f76620};
test_input[15664:15671] = '{32'h4280eff2, 32'h40c247ed, 32'h41007f55, 32'hc0f23e76, 32'h42966e49, 32'h4274e592, 32'hc28fd45c, 32'h42bd619a};
test_output[15664:15671] = '{32'h4280eff2, 32'h40c247ed, 32'h41007f55, 32'h0, 32'h42966e49, 32'h4274e592, 32'h0, 32'h42bd619a};
test_input[15672:15679] = '{32'h419d3916, 32'h426349fd, 32'h42982a3b, 32'hc25fd12c, 32'hc29061b8, 32'hc15a5031, 32'h42aff0ef, 32'hc2888de4};
test_output[15672:15679] = '{32'h419d3916, 32'h426349fd, 32'h42982a3b, 32'h0, 32'h0, 32'h0, 32'h42aff0ef, 32'h0};
test_input[15680:15687] = '{32'hc27fa409, 32'h426a6bf0, 32'h42c032aa, 32'h421eb743, 32'h42bfd90c, 32'hc1de9103, 32'hc260cea0, 32'hc2c4ad05};
test_output[15680:15687] = '{32'h0, 32'h426a6bf0, 32'h42c032aa, 32'h421eb743, 32'h42bfd90c, 32'h0, 32'h0, 32'h0};
test_input[15688:15695] = '{32'h41fa8aa7, 32'h403522d4, 32'hc2b0fd68, 32'hc25fea0c, 32'hc255a827, 32'h42947780, 32'h4224a083, 32'hc11fb0de};
test_output[15688:15695] = '{32'h41fa8aa7, 32'h403522d4, 32'h0, 32'h0, 32'h0, 32'h42947780, 32'h4224a083, 32'h0};
test_input[15696:15703] = '{32'hc2329d0b, 32'hc2b6cf65, 32'hc297bfd9, 32'hc1681279, 32'h42b9a386, 32'hc284ce9d, 32'hc245b419, 32'h3de4a78f};
test_output[15696:15703] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42b9a386, 32'h0, 32'h0, 32'h3de4a78f};
test_input[15704:15711] = '{32'hc11a34e0, 32'hc2aa5b25, 32'h4293ecc2, 32'hc1aefd32, 32'h42c2ce1e, 32'hc24c6a32, 32'h4206aca3, 32'h42bbc0b4};
test_output[15704:15711] = '{32'h0, 32'h0, 32'h4293ecc2, 32'h0, 32'h42c2ce1e, 32'h0, 32'h4206aca3, 32'h42bbc0b4};
test_input[15712:15719] = '{32'h41d1c14b, 32'h429c9947, 32'hc1f8214b, 32'h42a6cecd, 32'hc28a2e34, 32'h421d98ca, 32'h4286895d, 32'h42a45b8a};
test_output[15712:15719] = '{32'h41d1c14b, 32'h429c9947, 32'h0, 32'h42a6cecd, 32'h0, 32'h421d98ca, 32'h4286895d, 32'h42a45b8a};
test_input[15720:15727] = '{32'h428b9b9e, 32'h42b60275, 32'h41f9465d, 32'hc24dc8ee, 32'h428c2c71, 32'hc12506f6, 32'hc2c0b39d, 32'hc2c44e8b};
test_output[15720:15727] = '{32'h428b9b9e, 32'h42b60275, 32'h41f9465d, 32'h0, 32'h428c2c71, 32'h0, 32'h0, 32'h0};
test_input[15728:15735] = '{32'h4222bf3f, 32'hc26f6e12, 32'h42717630, 32'hc1207a8f, 32'hc1a671c7, 32'hc1d00857, 32'hbfaae984, 32'h420c0384};
test_output[15728:15735] = '{32'h4222bf3f, 32'h0, 32'h42717630, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420c0384};
test_input[15736:15743] = '{32'h409d5fca, 32'hc126b396, 32'h412d3456, 32'hc1e7fa66, 32'h42adc6b0, 32'h42705420, 32'hc2b46518, 32'hc14c3c14};
test_output[15736:15743] = '{32'h409d5fca, 32'h0, 32'h412d3456, 32'h0, 32'h42adc6b0, 32'h42705420, 32'h0, 32'h0};
test_input[15744:15751] = '{32'h428159e7, 32'h4288b167, 32'h4291ce92, 32'hc27d7e97, 32'hc2194ee2, 32'h40d80ce9, 32'hc258fd35, 32'hc0596557};
test_output[15744:15751] = '{32'h428159e7, 32'h4288b167, 32'h4291ce92, 32'h0, 32'h0, 32'h40d80ce9, 32'h0, 32'h0};
test_input[15752:15759] = '{32'h409bd26d, 32'hc1948c9c, 32'h42bf3709, 32'hc1b2f76e, 32'hc1ef57d8, 32'hc1fbaa53, 32'hc22e6bac, 32'hc25fb22b};
test_output[15752:15759] = '{32'h409bd26d, 32'h0, 32'h42bf3709, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15760:15767] = '{32'h4265d5bc, 32'hc2719879, 32'hc1d16242, 32'h426ddff2, 32'hc22a1210, 32'h42b38baa, 32'h4291e347, 32'hc2acb325};
test_output[15760:15767] = '{32'h4265d5bc, 32'h0, 32'h0, 32'h426ddff2, 32'h0, 32'h42b38baa, 32'h4291e347, 32'h0};
test_input[15768:15775] = '{32'hc12fdfce, 32'h42914061, 32'hc2365fea, 32'h429f7501, 32'h4221949a, 32'h42a3e83c, 32'hc24a4ea4, 32'h42c2eddd};
test_output[15768:15775] = '{32'h0, 32'h42914061, 32'h0, 32'h429f7501, 32'h4221949a, 32'h42a3e83c, 32'h0, 32'h42c2eddd};
test_input[15776:15783] = '{32'hc289e71a, 32'h429f677c, 32'hc27606c6, 32'hc2b47204, 32'hc21a4205, 32'hc2585c23, 32'hc2a917d0, 32'hc261da55};
test_output[15776:15783] = '{32'h0, 32'h429f677c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15784:15791] = '{32'hc29c9f98, 32'hc21f2451, 32'hc2b8a549, 32'hc28c3eb2, 32'hc152d9a8, 32'hc1c0299a, 32'h41ae5f9f, 32'hc1ac7142};
test_output[15784:15791] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ae5f9f, 32'h0};
test_input[15792:15799] = '{32'h41a6495b, 32'h41ad869a, 32'hc2b2ecda, 32'hc22d5d29, 32'hc17e1fce, 32'h42abf9fa, 32'h4062c981, 32'h42350d61};
test_output[15792:15799] = '{32'h41a6495b, 32'h41ad869a, 32'h0, 32'h0, 32'h0, 32'h42abf9fa, 32'h4062c981, 32'h42350d61};
test_input[15800:15807] = '{32'h42b03e43, 32'h42c70100, 32'h4220cd95, 32'hc19d363f, 32'hc2b07ad1, 32'hc256d2ba, 32'hc25b3b85, 32'h426c0af3};
test_output[15800:15807] = '{32'h42b03e43, 32'h42c70100, 32'h4220cd95, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426c0af3};
test_input[15808:15815] = '{32'h4299dbc3, 32'hc2ba54eb, 32'hc29f3848, 32'hc24177e7, 32'h42ae2bd1, 32'hc29d2c15, 32'h4286d763, 32'hc234664c};
test_output[15808:15815] = '{32'h4299dbc3, 32'h0, 32'h0, 32'h0, 32'h42ae2bd1, 32'h0, 32'h4286d763, 32'h0};
test_input[15816:15823] = '{32'hc2b08d39, 32'h42c5dc7e, 32'h4297a5a4, 32'hc217665a, 32'h3fa48087, 32'hc1068ee2, 32'hc282cff5, 32'hc29f60bb};
test_output[15816:15823] = '{32'h0, 32'h42c5dc7e, 32'h4297a5a4, 32'h0, 32'h3fa48087, 32'h0, 32'h0, 32'h0};
test_input[15824:15831] = '{32'hc1a82f97, 32'hc286c6cf, 32'hc2c33df7, 32'h42327866, 32'hc2bc0a42, 32'h416ff2a6, 32'hc04038e8, 32'h429489bd};
test_output[15824:15831] = '{32'h0, 32'h0, 32'h0, 32'h42327866, 32'h0, 32'h416ff2a6, 32'h0, 32'h429489bd};
test_input[15832:15839] = '{32'hc0449ba7, 32'h42a4313b, 32'hc2328c3a, 32'h42b205d0, 32'hc1b1bbee, 32'hc2935ed9, 32'hc29f65e0, 32'hc249ccc0};
test_output[15832:15839] = '{32'h0, 32'h42a4313b, 32'h0, 32'h42b205d0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[15840:15847] = '{32'hc2b9fba5, 32'h4296ba38, 32'hc283d6f7, 32'h42bc766f, 32'hc1f52e01, 32'hc256d012, 32'h3faf92ef, 32'h422314db};
test_output[15840:15847] = '{32'h0, 32'h4296ba38, 32'h0, 32'h42bc766f, 32'h0, 32'h0, 32'h3faf92ef, 32'h422314db};
test_input[15848:15855] = '{32'h4269c771, 32'hc1f7d0c2, 32'h4284ac9c, 32'h42aa47ac, 32'h4159db42, 32'hc1bdafc9, 32'h429ea349, 32'hc2a3a1ea};
test_output[15848:15855] = '{32'h4269c771, 32'h0, 32'h4284ac9c, 32'h42aa47ac, 32'h4159db42, 32'h0, 32'h429ea349, 32'h0};
test_input[15856:15863] = '{32'hc2537441, 32'hc2a051f8, 32'h428134b7, 32'h42914bff, 32'h400725de, 32'h4274b10a, 32'h41c66a4f, 32'h41852944};
test_output[15856:15863] = '{32'h0, 32'h0, 32'h428134b7, 32'h42914bff, 32'h400725de, 32'h4274b10a, 32'h41c66a4f, 32'h41852944};
test_input[15864:15871] = '{32'hc2779417, 32'h429298f3, 32'hc1fd96f3, 32'hc27aab28, 32'hc2662126, 32'h414d46ec, 32'hc13024d0, 32'h4245fe3c};
test_output[15864:15871] = '{32'h0, 32'h429298f3, 32'h0, 32'h0, 32'h0, 32'h414d46ec, 32'h0, 32'h4245fe3c};
test_input[15872:15879] = '{32'h424d143a, 32'h41a0ec80, 32'h41d29acb, 32'hc2392c61, 32'h427d79b4, 32'hc185227e, 32'h42539286, 32'hc0c1b281};
test_output[15872:15879] = '{32'h424d143a, 32'h41a0ec80, 32'h41d29acb, 32'h0, 32'h427d79b4, 32'h0, 32'h42539286, 32'h0};
test_input[15880:15887] = '{32'h4216cc69, 32'hc057eff9, 32'h41d1d42f, 32'hc2633ac4, 32'h41165b39, 32'hc0c122c7, 32'hc29a8730, 32'hc2819b3e};
test_output[15880:15887] = '{32'h4216cc69, 32'h0, 32'h41d1d42f, 32'h0, 32'h41165b39, 32'h0, 32'h0, 32'h0};
test_input[15888:15895] = '{32'h42b49aa4, 32'h42935869, 32'hc1d7a321, 32'h42b17c28, 32'h424c314c, 32'h42317fab, 32'h41cda7ce, 32'h42552c0f};
test_output[15888:15895] = '{32'h42b49aa4, 32'h42935869, 32'h0, 32'h42b17c28, 32'h424c314c, 32'h42317fab, 32'h41cda7ce, 32'h42552c0f};
test_input[15896:15903] = '{32'hc29e450c, 32'h42601e6f, 32'hc25c12da, 32'hc11ba5b0, 32'h417cd20f, 32'hc25690ad, 32'hbf97a383, 32'h425f47f8};
test_output[15896:15903] = '{32'h0, 32'h42601e6f, 32'h0, 32'h0, 32'h417cd20f, 32'h0, 32'h0, 32'h425f47f8};
test_input[15904:15911] = '{32'hc15eb545, 32'h3f84e64a, 32'h424e3127, 32'h420b2923, 32'hc28100ed, 32'h4286be4b, 32'hc21bf984, 32'hc296342c};
test_output[15904:15911] = '{32'h0, 32'h3f84e64a, 32'h424e3127, 32'h420b2923, 32'h0, 32'h4286be4b, 32'h0, 32'h0};
test_input[15912:15919] = '{32'h42777e95, 32'hc2972d59, 32'hc186a650, 32'hc2013590, 32'hc1229aec, 32'h41af610f, 32'h4192ffce, 32'hc25fcd04};
test_output[15912:15919] = '{32'h42777e95, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41af610f, 32'h4192ffce, 32'h0};
test_input[15920:15927] = '{32'h42a8e453, 32'h4205a5cf, 32'hc10d1f11, 32'h416b2caf, 32'h42290fda, 32'hc24faed2, 32'h4272204c, 32'hc1c68f83};
test_output[15920:15927] = '{32'h42a8e453, 32'h4205a5cf, 32'h0, 32'h416b2caf, 32'h42290fda, 32'h0, 32'h4272204c, 32'h0};
test_input[15928:15935] = '{32'hc2ad8613, 32'h42ba3b47, 32'h4225856a, 32'hc25bbcb1, 32'h42b44fb6, 32'hc2333d69, 32'h4247caf7, 32'hc1d9c4b3};
test_output[15928:15935] = '{32'h0, 32'h42ba3b47, 32'h4225856a, 32'h0, 32'h42b44fb6, 32'h0, 32'h4247caf7, 32'h0};
test_input[15936:15943] = '{32'h42b5f789, 32'h410cf89c, 32'h417cf332, 32'hbf1a759e, 32'h425ed04f, 32'hc21b6e08, 32'h4215e132, 32'h42b9b68d};
test_output[15936:15943] = '{32'h42b5f789, 32'h410cf89c, 32'h417cf332, 32'h0, 32'h425ed04f, 32'h0, 32'h4215e132, 32'h42b9b68d};
test_input[15944:15951] = '{32'h42a4b076, 32'hc29f4eae, 32'hc280120f, 32'hc285451b, 32'h42883800, 32'hc1b0bcbf, 32'h40ec1fed, 32'h4116b91e};
test_output[15944:15951] = '{32'h42a4b076, 32'h0, 32'h0, 32'h0, 32'h42883800, 32'h0, 32'h40ec1fed, 32'h4116b91e};
test_input[15952:15959] = '{32'h42225131, 32'hc2848ac0, 32'h42596d81, 32'h409abca4, 32'h40925ec7, 32'hc29f55c5, 32'h421b9646, 32'h42113eb7};
test_output[15952:15959] = '{32'h42225131, 32'h0, 32'h42596d81, 32'h409abca4, 32'h40925ec7, 32'h0, 32'h421b9646, 32'h42113eb7};
test_input[15960:15967] = '{32'h42ab87e0, 32'h42723dff, 32'h414f84c4, 32'h41fdf8d4, 32'hc02fd63b, 32'hc18c40aa, 32'h4210c496, 32'hc1296634};
test_output[15960:15967] = '{32'h42ab87e0, 32'h42723dff, 32'h414f84c4, 32'h41fdf8d4, 32'h0, 32'h0, 32'h4210c496, 32'h0};
test_input[15968:15975] = '{32'hc24e21a7, 32'h4140ed84, 32'hc1f5d910, 32'h42852fa7, 32'hc2ab48e8, 32'h4264a16c, 32'hc21f52ea, 32'h42acaa0c};
test_output[15968:15975] = '{32'h0, 32'h4140ed84, 32'h0, 32'h42852fa7, 32'h0, 32'h4264a16c, 32'h0, 32'h42acaa0c};
test_input[15976:15983] = '{32'hc261c966, 32'h426590a2, 32'hc272c15e, 32'h41adb16c, 32'h42c29809, 32'h424ec40d, 32'h428ed533, 32'h41f3ed93};
test_output[15976:15983] = '{32'h0, 32'h426590a2, 32'h0, 32'h41adb16c, 32'h42c29809, 32'h424ec40d, 32'h428ed533, 32'h41f3ed93};
test_input[15984:15991] = '{32'h41720833, 32'hc28dd5e0, 32'h42b39fd3, 32'h41bb4d7c, 32'h40869e98, 32'h4179a318, 32'h428702d5, 32'h4276ba06};
test_output[15984:15991] = '{32'h41720833, 32'h0, 32'h42b39fd3, 32'h41bb4d7c, 32'h40869e98, 32'h4179a318, 32'h428702d5, 32'h4276ba06};
test_input[15992:15999] = '{32'hc1c67e0d, 32'hc2a96983, 32'hc25fe92e, 32'h42244043, 32'hc0ee42fb, 32'hc28f5613, 32'hc2363dbc, 32'hbec243c1};
test_output[15992:15999] = '{32'h0, 32'h0, 32'h0, 32'h42244043, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16000:16007] = '{32'h42887193, 32'hc29fd4e1, 32'hc0e45553, 32'h42c566ab, 32'hc1e2c1d6, 32'h424e11c3, 32'hc2b16239, 32'hc2b9b7bd};
test_output[16000:16007] = '{32'h42887193, 32'h0, 32'h0, 32'h42c566ab, 32'h0, 32'h424e11c3, 32'h0, 32'h0};
test_input[16008:16015] = '{32'h4266eeb9, 32'hc1ac491b, 32'h42b3b95b, 32'hc2331cb2, 32'h429d7da7, 32'h4276fdd9, 32'hc263d53f, 32'h4279b9a3};
test_output[16008:16015] = '{32'h4266eeb9, 32'h0, 32'h42b3b95b, 32'h0, 32'h429d7da7, 32'h4276fdd9, 32'h0, 32'h4279b9a3};
test_input[16016:16023] = '{32'hc26c037d, 32'hc0a8a3dc, 32'hc0b38193, 32'h4233c2c1, 32'h41293ed6, 32'hc1451b4d, 32'h410ae908, 32'hc2083bf2};
test_output[16016:16023] = '{32'h0, 32'h0, 32'h0, 32'h4233c2c1, 32'h41293ed6, 32'h0, 32'h410ae908, 32'h0};
test_input[16024:16031] = '{32'hc23512f2, 32'hc28a5075, 32'h41cc149c, 32'hc05bbb76, 32'hc26375e5, 32'hc0a221fe, 32'hc2550106, 32'hc29dae5e};
test_output[16024:16031] = '{32'h0, 32'h0, 32'h41cc149c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16032:16039] = '{32'h42bb244e, 32'h426d65c9, 32'h416f27f5, 32'h42aeaf73, 32'hc28947f4, 32'hc1e86d14, 32'h42c4dd0f, 32'h40e878ba};
test_output[16032:16039] = '{32'h42bb244e, 32'h426d65c9, 32'h416f27f5, 32'h42aeaf73, 32'h0, 32'h0, 32'h42c4dd0f, 32'h40e878ba};
test_input[16040:16047] = '{32'hc0d4e107, 32'h422ec383, 32'hc21df682, 32'h42649c1f, 32'h42a368a7, 32'hc241defe, 32'hc2c1d4cf, 32'hc29debfb};
test_output[16040:16047] = '{32'h0, 32'h422ec383, 32'h0, 32'h42649c1f, 32'h42a368a7, 32'h0, 32'h0, 32'h0};
test_input[16048:16055] = '{32'hc2928c3a, 32'h4216205c, 32'hc286228a, 32'hc231b737, 32'hc29712d1, 32'h42bdf3b6, 32'h41b76c70, 32'hc2a25aa2};
test_output[16048:16055] = '{32'h0, 32'h4216205c, 32'h0, 32'h0, 32'h0, 32'h42bdf3b6, 32'h41b76c70, 32'h0};
test_input[16056:16063] = '{32'h428d0fb2, 32'hc220280c, 32'hc24b6de3, 32'h426ddf5e, 32'h41f3b93f, 32'h4201f95f, 32'h4120292a, 32'hc294ae7f};
test_output[16056:16063] = '{32'h428d0fb2, 32'h0, 32'h0, 32'h426ddf5e, 32'h41f3b93f, 32'h4201f95f, 32'h4120292a, 32'h0};
test_input[16064:16071] = '{32'hc1a576bc, 32'h42791d81, 32'h420c326c, 32'hc1deea21, 32'hc27d8343, 32'hc166dc5c, 32'h424dfdf5, 32'hc183683f};
test_output[16064:16071] = '{32'h0, 32'h42791d81, 32'h420c326c, 32'h0, 32'h0, 32'h0, 32'h424dfdf5, 32'h0};
test_input[16072:16079] = '{32'hc2a86a81, 32'hc2c3c794, 32'h41de3001, 32'h423a0f92, 32'h422b9279, 32'h4055f019, 32'h42b5e286, 32'h42bcbde8};
test_output[16072:16079] = '{32'h0, 32'h0, 32'h41de3001, 32'h423a0f92, 32'h422b9279, 32'h4055f019, 32'h42b5e286, 32'h42bcbde8};
test_input[16080:16087] = '{32'hc1cde925, 32'hc2aefbf8, 32'hc29c949f, 32'hc290b517, 32'h41c643c6, 32'h41846a48, 32'h42b25dca, 32'hc289a982};
test_output[16080:16087] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41c643c6, 32'h41846a48, 32'h42b25dca, 32'h0};
test_input[16088:16095] = '{32'h4183f09e, 32'hc20702e9, 32'h42bec0be, 32'hc2751f02, 32'h41d3df40, 32'hc2c33086, 32'hc26d3b7e, 32'h4140b596};
test_output[16088:16095] = '{32'h4183f09e, 32'h0, 32'h42bec0be, 32'h0, 32'h41d3df40, 32'h0, 32'h0, 32'h4140b596};
test_input[16096:16103] = '{32'h418db81a, 32'h42b6b088, 32'hc1d8d65d, 32'h4201caef, 32'h42713db9, 32'hc293f376, 32'h4155069c, 32'hc28f3f1e};
test_output[16096:16103] = '{32'h418db81a, 32'h42b6b088, 32'h0, 32'h4201caef, 32'h42713db9, 32'h0, 32'h4155069c, 32'h0};
test_input[16104:16111] = '{32'hc195a460, 32'h4299e97f, 32'h42615ccd, 32'h42b6ca57, 32'hbf26e5d9, 32'hc22373b7, 32'hc29ad6cf, 32'hc1941771};
test_output[16104:16111] = '{32'h0, 32'h4299e97f, 32'h42615ccd, 32'h42b6ca57, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16112:16119] = '{32'h429d448b, 32'h429496ec, 32'hbf0b459d, 32'h40938064, 32'hc1810756, 32'h4296a3b7, 32'hc298c530, 32'hc197d04d};
test_output[16112:16119] = '{32'h429d448b, 32'h429496ec, 32'h0, 32'h40938064, 32'h0, 32'h4296a3b7, 32'h0, 32'h0};
test_input[16120:16127] = '{32'h426d3bfc, 32'h41b84f2a, 32'h4281ba87, 32'h42307dce, 32'hc2924600, 32'h4221af51, 32'h423b916b, 32'hc2c6aaf5};
test_output[16120:16127] = '{32'h426d3bfc, 32'h41b84f2a, 32'h4281ba87, 32'h42307dce, 32'h0, 32'h4221af51, 32'h423b916b, 32'h0};
test_input[16128:16135] = '{32'h424dd52d, 32'h42b78db1, 32'h426e9853, 32'hc22d7076, 32'hc2a29ed4, 32'h422d57bf, 32'h41d9477e, 32'hc27df062};
test_output[16128:16135] = '{32'h424dd52d, 32'h42b78db1, 32'h426e9853, 32'h0, 32'h0, 32'h422d57bf, 32'h41d9477e, 32'h0};
test_input[16136:16143] = '{32'h411eddec, 32'hc2c4b768, 32'h41c961c2, 32'hc2909ac1, 32'h425125de, 32'hc220e347, 32'h404e8903, 32'h422d08b2};
test_output[16136:16143] = '{32'h411eddec, 32'h0, 32'h41c961c2, 32'h0, 32'h425125de, 32'h0, 32'h404e8903, 32'h422d08b2};
test_input[16144:16151] = '{32'h4197318a, 32'hc27916b9, 32'h428ff37c, 32'hc2af4b04, 32'hc25cbbfc, 32'h4243f848, 32'h41e1162d, 32'hc2002c72};
test_output[16144:16151] = '{32'h4197318a, 32'h0, 32'h428ff37c, 32'h0, 32'h0, 32'h4243f848, 32'h41e1162d, 32'h0};
test_input[16152:16159] = '{32'h41ca21ea, 32'hc2576f3a, 32'h428c6619, 32'h42a0f323, 32'h41eb0f60, 32'h42bf511f, 32'hc22e2ecd, 32'hc147c08c};
test_output[16152:16159] = '{32'h41ca21ea, 32'h0, 32'h428c6619, 32'h42a0f323, 32'h41eb0f60, 32'h42bf511f, 32'h0, 32'h0};
test_input[16160:16167] = '{32'h41e042dc, 32'hc1f6ef1e, 32'h40d82039, 32'h41c5d8a2, 32'hc28daa62, 32'h42a1be19, 32'h429a1261, 32'hc190f29d};
test_output[16160:16167] = '{32'h41e042dc, 32'h0, 32'h40d82039, 32'h41c5d8a2, 32'h0, 32'h42a1be19, 32'h429a1261, 32'h0};
test_input[16168:16175] = '{32'hc2a4af36, 32'h429964c2, 32'hc17555f8, 32'hc2c0f7c7, 32'hc0724867, 32'hc24da0da, 32'hc2864d48, 32'h4213d0d1};
test_output[16168:16175] = '{32'h0, 32'h429964c2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4213d0d1};
test_input[16176:16183] = '{32'h4242e44e, 32'h4246545d, 32'hc28a1f0e, 32'h42a1063c, 32'h412a0168, 32'hc2b9ee0c, 32'hc1fa51b4, 32'h4241699c};
test_output[16176:16183] = '{32'h4242e44e, 32'h4246545d, 32'h0, 32'h42a1063c, 32'h412a0168, 32'h0, 32'h0, 32'h4241699c};
test_input[16184:16191] = '{32'hc190124f, 32'hc24e7269, 32'h41867bdd, 32'h423fe5bf, 32'h4270e28c, 32'hc2a72a57, 32'hc2bd8511, 32'h42a1a165};
test_output[16184:16191] = '{32'h0, 32'h0, 32'h41867bdd, 32'h423fe5bf, 32'h4270e28c, 32'h0, 32'h0, 32'h42a1a165};
test_input[16192:16199] = '{32'h42993f26, 32'hc28a3782, 32'h42be118d, 32'hc159148f, 32'hc1a45131, 32'h42206e20, 32'hc272df5c, 32'hc1f3bd74};
test_output[16192:16199] = '{32'h42993f26, 32'h0, 32'h42be118d, 32'h0, 32'h0, 32'h42206e20, 32'h0, 32'h0};
test_input[16200:16207] = '{32'h4041ea7c, 32'hc25a3a92, 32'h4283ebd2, 32'h42b8df31, 32'h42234fa4, 32'h417c0f54, 32'h41965e3b, 32'hc2c1a03c};
test_output[16200:16207] = '{32'h4041ea7c, 32'h0, 32'h4283ebd2, 32'h42b8df31, 32'h42234fa4, 32'h417c0f54, 32'h41965e3b, 32'h0};
test_input[16208:16215] = '{32'hc11dfc8c, 32'hc25442e0, 32'hc2985839, 32'h429b67ed, 32'h41d41a94, 32'h42ad04d3, 32'h42281fa6, 32'h41e8b56d};
test_output[16208:16215] = '{32'h0, 32'h0, 32'h0, 32'h429b67ed, 32'h41d41a94, 32'h42ad04d3, 32'h42281fa6, 32'h41e8b56d};
test_input[16216:16223] = '{32'hc2833672, 32'hc267ec11, 32'h428f63b7, 32'hc2894606, 32'hc2b0c489, 32'h423b9de8, 32'hc1a23c96, 32'hc0e28650};
test_output[16216:16223] = '{32'h0, 32'h0, 32'h428f63b7, 32'h0, 32'h0, 32'h423b9de8, 32'h0, 32'h0};
test_input[16224:16231] = '{32'h41e9df3b, 32'h3f456fd3, 32'hc1b32673, 32'hc29645a4, 32'h4090c1f3, 32'h4080b7e1, 32'h424eea76, 32'hc28c01cb};
test_output[16224:16231] = '{32'h41e9df3b, 32'h3f456fd3, 32'h0, 32'h0, 32'h4090c1f3, 32'h4080b7e1, 32'h424eea76, 32'h0};
test_input[16232:16239] = '{32'h429374a8, 32'hc1a453ed, 32'hc2b83579, 32'hc1f7bd28, 32'h423a65c6, 32'h424104eb, 32'h428d300c, 32'h40b68d48};
test_output[16232:16239] = '{32'h429374a8, 32'h0, 32'h0, 32'h0, 32'h423a65c6, 32'h424104eb, 32'h428d300c, 32'h40b68d48};
test_input[16240:16247] = '{32'h428e7ebe, 32'h429f0ec5, 32'h420aa6df, 32'h423d5405, 32'h426669ea, 32'h41aa7bba, 32'h425770d5, 32'hc2ba03e9};
test_output[16240:16247] = '{32'h428e7ebe, 32'h429f0ec5, 32'h420aa6df, 32'h423d5405, 32'h426669ea, 32'h41aa7bba, 32'h425770d5, 32'h0};
test_input[16248:16255] = '{32'hc2b05158, 32'hc1807d4a, 32'h42c67e7e, 32'h419c1fed, 32'hc29217a0, 32'h4277ae67, 32'h4291f953, 32'hc16f9723};
test_output[16248:16255] = '{32'h0, 32'h0, 32'h42c67e7e, 32'h419c1fed, 32'h0, 32'h4277ae67, 32'h4291f953, 32'h0};
test_input[16256:16263] = '{32'hc2ba7da9, 32'hc2037ace, 32'h41f4f3d8, 32'h417b7b46, 32'hc2a5fd2c, 32'hc1a78f62, 32'h42b76176, 32'h41e88dde};
test_output[16256:16263] = '{32'h0, 32'h0, 32'h41f4f3d8, 32'h417b7b46, 32'h0, 32'h0, 32'h42b76176, 32'h41e88dde};
test_input[16264:16271] = '{32'hc2410b8f, 32'hc2a06abb, 32'hc1b006e2, 32'h42bf33fe, 32'h4209d128, 32'h4067b36f, 32'hc2894f01, 32'hc258a7e3};
test_output[16264:16271] = '{32'h0, 32'h0, 32'h0, 32'h42bf33fe, 32'h4209d128, 32'h4067b36f, 32'h0, 32'h0};
test_input[16272:16279] = '{32'hc1c71a79, 32'h42aeac7c, 32'h427bd5dc, 32'h41c232d7, 32'h42096b8a, 32'hbfe0ffe2, 32'h4279b0b7, 32'hc2b75ae0};
test_output[16272:16279] = '{32'h0, 32'h42aeac7c, 32'h427bd5dc, 32'h41c232d7, 32'h42096b8a, 32'h0, 32'h4279b0b7, 32'h0};
test_input[16280:16287] = '{32'hc2833678, 32'h428599b6, 32'hc1e15d89, 32'h429f647b, 32'hc24d90f1, 32'hc2a64c25, 32'h426e4b2f, 32'hc2b75fb1};
test_output[16280:16287] = '{32'h0, 32'h428599b6, 32'h0, 32'h429f647b, 32'h0, 32'h0, 32'h426e4b2f, 32'h0};
test_input[16288:16295] = '{32'hc2b60b6e, 32'hc049819b, 32'hc1561f9f, 32'hc2acb5c9, 32'hc28566b3, 32'hc2534582, 32'h4224af97, 32'hc203adc6};
test_output[16288:16295] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4224af97, 32'h0};
test_input[16296:16303] = '{32'hc1b4cdd8, 32'h42af55cb, 32'hc2938502, 32'hbf48d3e3, 32'hc299ca48, 32'hc2bf3665, 32'hc2a12622, 32'h41c2ac07};
test_output[16296:16303] = '{32'h0, 32'h42af55cb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41c2ac07};
test_input[16304:16311] = '{32'h41046291, 32'hc16363aa, 32'hc17a9b3c, 32'h41aa2a8c, 32'hc2abcdd3, 32'h41954677, 32'h41919178, 32'hc199f279};
test_output[16304:16311] = '{32'h41046291, 32'h0, 32'h0, 32'h41aa2a8c, 32'h0, 32'h41954677, 32'h41919178, 32'h0};
test_input[16312:16319] = '{32'h42a039d9, 32'hc1b9136b, 32'h42ba125b, 32'h42b8626c, 32'hc250535a, 32'h422eeec1, 32'h42055d4e, 32'hc207c656};
test_output[16312:16319] = '{32'h42a039d9, 32'h0, 32'h42ba125b, 32'h42b8626c, 32'h0, 32'h422eeec1, 32'h42055d4e, 32'h0};
test_input[16320:16327] = '{32'hc1cd3d3d, 32'h40eb3c4a, 32'hc1b8c698, 32'h422dc2f6, 32'h411ccbb7, 32'hc2b01d73, 32'hc242ff53, 32'hbfb579ff};
test_output[16320:16327] = '{32'h0, 32'h40eb3c4a, 32'h0, 32'h422dc2f6, 32'h411ccbb7, 32'h0, 32'h0, 32'h0};
test_input[16328:16335] = '{32'h429b263b, 32'h429dd02a, 32'h41eb5edf, 32'h4253e785, 32'hc29bc546, 32'h41f12d2d, 32'h40304d55, 32'hc2929696};
test_output[16328:16335] = '{32'h429b263b, 32'h429dd02a, 32'h41eb5edf, 32'h4253e785, 32'h0, 32'h41f12d2d, 32'h40304d55, 32'h0};
test_input[16336:16343] = '{32'h4205a81e, 32'h42092a0f, 32'hc28e27ae, 32'h42099db1, 32'hc2c22975, 32'hc1bbad9a, 32'h41d507ae, 32'hc0ace749};
test_output[16336:16343] = '{32'h4205a81e, 32'h42092a0f, 32'h0, 32'h42099db1, 32'h0, 32'h0, 32'h41d507ae, 32'h0};
test_input[16344:16351] = '{32'h424679b6, 32'h4282c73a, 32'hc274065c, 32'h42436fe8, 32'hc2b028ee, 32'h425bece4, 32'hc2be6689, 32'hc12abfb6};
test_output[16344:16351] = '{32'h424679b6, 32'h4282c73a, 32'h0, 32'h42436fe8, 32'h0, 32'h425bece4, 32'h0, 32'h0};
test_input[16352:16359] = '{32'h42aa0b07, 32'h424ee08e, 32'h428ef3eb, 32'h41cc28a9, 32'hc2514a42, 32'h428133b2, 32'h42a9cc0b, 32'hc29c72da};
test_output[16352:16359] = '{32'h42aa0b07, 32'h424ee08e, 32'h428ef3eb, 32'h41cc28a9, 32'h0, 32'h428133b2, 32'h42a9cc0b, 32'h0};
test_input[16360:16367] = '{32'h41e92042, 32'hc2ad2c6f, 32'h419e6bb4, 32'h425b001a, 32'h40e4e143, 32'h428ea6c2, 32'h42b574c4, 32'h426c9444};
test_output[16360:16367] = '{32'h41e92042, 32'h0, 32'h419e6bb4, 32'h425b001a, 32'h40e4e143, 32'h428ea6c2, 32'h42b574c4, 32'h426c9444};
test_input[16368:16375] = '{32'hc2654cf0, 32'hc2537b98, 32'hc1d7a010, 32'hc2a8dfb3, 32'hc1fd1757, 32'h40af3799, 32'h4151ec70, 32'h4154da5a};
test_output[16368:16375] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40af3799, 32'h4151ec70, 32'h4154da5a};
test_input[16376:16383] = '{32'h429f8346, 32'hc1669963, 32'h42c37aa1, 32'h41cd2ce9, 32'h42891a33, 32'h41afbffa, 32'h4177f4ce, 32'hc26f8651};
test_output[16376:16383] = '{32'h429f8346, 32'h0, 32'h42c37aa1, 32'h41cd2ce9, 32'h42891a33, 32'h41afbffa, 32'h4177f4ce, 32'h0};
test_input[16384:16391] = '{32'hc29fe088, 32'hc2abc630, 32'hc250a3ce, 32'hc2adede2, 32'h423b32b3, 32'hc1f3b63c, 32'h408ed1b6, 32'hc28dc211};
test_output[16384:16391] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h423b32b3, 32'h0, 32'h408ed1b6, 32'h0};
test_input[16392:16399] = '{32'h418f3935, 32'hc29e907b, 32'hc290504f, 32'h4152f147, 32'hc25eebf0, 32'hc2b1aebf, 32'h41f08aa7, 32'h4199d7a0};
test_output[16392:16399] = '{32'h418f3935, 32'h0, 32'h0, 32'h4152f147, 32'h0, 32'h0, 32'h41f08aa7, 32'h4199d7a0};
test_input[16400:16407] = '{32'hc209405f, 32'h4285d147, 32'h42252ff2, 32'h42914c1c, 32'hc0d91861, 32'h4287dc0a, 32'h41eaf547, 32'h422d83ae};
test_output[16400:16407] = '{32'h0, 32'h4285d147, 32'h42252ff2, 32'h42914c1c, 32'h0, 32'h4287dc0a, 32'h41eaf547, 32'h422d83ae};
test_input[16408:16415] = '{32'h400e83c5, 32'h41ae5a15, 32'hc2797604, 32'h42606d42, 32'h42aa4759, 32'hc2aef180, 32'hc27221f8, 32'hc1ee67fc};
test_output[16408:16415] = '{32'h400e83c5, 32'h41ae5a15, 32'h0, 32'h42606d42, 32'h42aa4759, 32'h0, 32'h0, 32'h0};
test_input[16416:16423] = '{32'h42b0f5fc, 32'h3f24a93d, 32'h4267accb, 32'hbfbe4862, 32'h422922b6, 32'h42c2fbc2, 32'h4289a043, 32'hc2b13882};
test_output[16416:16423] = '{32'h42b0f5fc, 32'h3f24a93d, 32'h4267accb, 32'h0, 32'h422922b6, 32'h42c2fbc2, 32'h4289a043, 32'h0};
test_input[16424:16431] = '{32'h419a8964, 32'hc288de9f, 32'hc2adc11b, 32'hc29e6db7, 32'hc2958e8e, 32'hc2041911, 32'hc27cb5e3, 32'h424c9d37};
test_output[16424:16431] = '{32'h419a8964, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h424c9d37};
test_input[16432:16439] = '{32'hc25c137d, 32'h429c8ca8, 32'hc254b8b7, 32'h41f3f43d, 32'h4268a927, 32'hc1ce9a74, 32'h40f3da4b, 32'hc28f4d25};
test_output[16432:16439] = '{32'h0, 32'h429c8ca8, 32'h0, 32'h41f3f43d, 32'h4268a927, 32'h0, 32'h40f3da4b, 32'h0};
test_input[16440:16447] = '{32'h426ded99, 32'hc24b595c, 32'hc1d79c23, 32'hc25dd4bd, 32'hc23e52f9, 32'hc2b896cb, 32'hbec18ad4, 32'h4274f257};
test_output[16440:16447] = '{32'h426ded99, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4274f257};
test_input[16448:16455] = '{32'hc253cca0, 32'hc275fdb7, 32'hc1e057e8, 32'h429204dc, 32'h416bb478, 32'h424e5f6a, 32'h429c19de, 32'hc2a710c1};
test_output[16448:16455] = '{32'h0, 32'h0, 32'h0, 32'h429204dc, 32'h416bb478, 32'h424e5f6a, 32'h429c19de, 32'h0};
test_input[16456:16463] = '{32'hc01a05a1, 32'hc2af92ac, 32'hc2b4023a, 32'hc1147b60, 32'hc184eda2, 32'hc268c88e, 32'h40a18792, 32'h42655d3c};
test_output[16456:16463] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40a18792, 32'h42655d3c};
test_input[16464:16471] = '{32'h40ca5e00, 32'h42a3b8c4, 32'h41f43ad7, 32'hc196a0c3, 32'h42910409, 32'h427f1b22, 32'hc222de3f, 32'h417aad86};
test_output[16464:16471] = '{32'h40ca5e00, 32'h42a3b8c4, 32'h41f43ad7, 32'h0, 32'h42910409, 32'h427f1b22, 32'h0, 32'h417aad86};
test_input[16472:16479] = '{32'hc285f607, 32'h41ae7300, 32'hc2a64c0e, 32'hc28ae4bd, 32'hc2731d2a, 32'hc20dc5df, 32'h428e1e98, 32'h428d40cc};
test_output[16472:16479] = '{32'h0, 32'h41ae7300, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428e1e98, 32'h428d40cc};
test_input[16480:16487] = '{32'h42c1d1a7, 32'hc23a0636, 32'h421f7397, 32'hc26640c4, 32'hc210bbe2, 32'hc28b4ab5, 32'h42b3a63f, 32'hc285bc42};
test_output[16480:16487] = '{32'h42c1d1a7, 32'h0, 32'h421f7397, 32'h0, 32'h0, 32'h0, 32'h42b3a63f, 32'h0};
test_input[16488:16495] = '{32'hc2474a75, 32'hc29064d3, 32'h4292a166, 32'hc1e12653, 32'h423c1e78, 32'hc1d97457, 32'hc2a3f410, 32'h42ba5c11};
test_output[16488:16495] = '{32'h0, 32'h0, 32'h4292a166, 32'h0, 32'h423c1e78, 32'h0, 32'h0, 32'h42ba5c11};
test_input[16496:16503] = '{32'hc25f885b, 32'h42b10ff7, 32'h42a53db6, 32'h4115d5d8, 32'h4204c67a, 32'hc247b050, 32'h4299dee2, 32'hc24d4b1d};
test_output[16496:16503] = '{32'h0, 32'h42b10ff7, 32'h42a53db6, 32'h4115d5d8, 32'h4204c67a, 32'h0, 32'h4299dee2, 32'h0};
test_input[16504:16511] = '{32'h418f4d58, 32'h416cb607, 32'h41cf288f, 32'hc1ab5972, 32'hc2c0ab89, 32'hc26a9e33, 32'h42a5a602, 32'hc280e579};
test_output[16504:16511] = '{32'h418f4d58, 32'h416cb607, 32'h41cf288f, 32'h0, 32'h0, 32'h0, 32'h42a5a602, 32'h0};
test_input[16512:16519] = '{32'hc2b2a44f, 32'h423426c8, 32'h4299868c, 32'hc27974d0, 32'hc24aa59d, 32'h42b0ddcd, 32'h41f9e789, 32'h41c229a2};
test_output[16512:16519] = '{32'h0, 32'h423426c8, 32'h4299868c, 32'h0, 32'h0, 32'h42b0ddcd, 32'h41f9e789, 32'h41c229a2};
test_input[16520:16527] = '{32'hc19e1dbe, 32'h418cbb9a, 32'h414be06e, 32'h400d38d6, 32'h4258d0e6, 32'h41d65d7c, 32'h420385a8, 32'hc283f17b};
test_output[16520:16527] = '{32'h0, 32'h418cbb9a, 32'h414be06e, 32'h400d38d6, 32'h4258d0e6, 32'h41d65d7c, 32'h420385a8, 32'h0};
test_input[16528:16535] = '{32'hc29d0633, 32'h4219af69, 32'h41ac76ba, 32'hc24768e4, 32'hc227089b, 32'hc0dc9021, 32'h42056f1f, 32'hc28df562};
test_output[16528:16535] = '{32'h0, 32'h4219af69, 32'h41ac76ba, 32'h0, 32'h0, 32'h0, 32'h42056f1f, 32'h0};
test_input[16536:16543] = '{32'hc2969b84, 32'h42953f9a, 32'h42beb230, 32'h421a928b, 32'h41d4ccb1, 32'hc2a2f6b0, 32'hc283c2e8, 32'h42c18faa};
test_output[16536:16543] = '{32'h0, 32'h42953f9a, 32'h42beb230, 32'h421a928b, 32'h41d4ccb1, 32'h0, 32'h0, 32'h42c18faa};
test_input[16544:16551] = '{32'h41a09c72, 32'hc23e8a47, 32'hc258833a, 32'hc2732e62, 32'h42ab0321, 32'hc25fdd66, 32'h416f8f1e, 32'hc2649ae4};
test_output[16544:16551] = '{32'h41a09c72, 32'h0, 32'h0, 32'h0, 32'h42ab0321, 32'h0, 32'h416f8f1e, 32'h0};
test_input[16552:16559] = '{32'h3fd98942, 32'h41f23d63, 32'h409a02e6, 32'hc283bd9f, 32'hc038065d, 32'h424c1b1d, 32'hc2772b78, 32'h3fb43e04};
test_output[16552:16559] = '{32'h3fd98942, 32'h41f23d63, 32'h409a02e6, 32'h0, 32'h0, 32'h424c1b1d, 32'h0, 32'h3fb43e04};
test_input[16560:16567] = '{32'h42a34b3b, 32'hc285cdb7, 32'h418640f2, 32'hc1f74dce, 32'hc2c706c0, 32'hc06b6fc8, 32'h42b0f852, 32'hc1c19e51};
test_output[16560:16567] = '{32'h42a34b3b, 32'h0, 32'h418640f2, 32'h0, 32'h0, 32'h0, 32'h42b0f852, 32'h0};
test_input[16568:16575] = '{32'h42bb7c9c, 32'hc232c9e3, 32'hc146ac38, 32'h4249155d, 32'hc22437f8, 32'h423a3e0a, 32'hc22da885, 32'h424b25bd};
test_output[16568:16575] = '{32'h42bb7c9c, 32'h0, 32'h0, 32'h4249155d, 32'h0, 32'h423a3e0a, 32'h0, 32'h424b25bd};
test_input[16576:16583] = '{32'hc25c4956, 32'h428eb217, 32'h40ea6934, 32'hc244b32a, 32'hc00e7e65, 32'h42415c47, 32'h425fa6b3, 32'h4113b0bf};
test_output[16576:16583] = '{32'h0, 32'h428eb217, 32'h40ea6934, 32'h0, 32'h0, 32'h42415c47, 32'h425fa6b3, 32'h4113b0bf};
test_input[16584:16591] = '{32'h42956dda, 32'h41cd189b, 32'h42c04518, 32'h41acad9a, 32'hc125c960, 32'h422772f0, 32'h420a99de, 32'hc0dfdc83};
test_output[16584:16591] = '{32'h42956dda, 32'h41cd189b, 32'h42c04518, 32'h41acad9a, 32'h0, 32'h422772f0, 32'h420a99de, 32'h0};
test_input[16592:16599] = '{32'hc22f2a5b, 32'hc2859940, 32'hc275aac4, 32'hc286c313, 32'hc217fee0, 32'hc25c6909, 32'hc10ce87f, 32'hc2b1ab97};
test_output[16592:16599] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[16600:16607] = '{32'hc2a84fad, 32'hc1498ca4, 32'h423ab7f8, 32'hc16c898f, 32'h42b8e888, 32'hc24cb914, 32'h42a00728, 32'h42616dc4};
test_output[16600:16607] = '{32'h0, 32'h0, 32'h423ab7f8, 32'h0, 32'h42b8e888, 32'h0, 32'h42a00728, 32'h42616dc4};
test_input[16608:16615] = '{32'h42764262, 32'hc2b9d27b, 32'h42a17789, 32'h42c388fa, 32'h42469111, 32'h419a4c3a, 32'h40426e95, 32'h41866c79};
test_output[16608:16615] = '{32'h42764262, 32'h0, 32'h42a17789, 32'h42c388fa, 32'h42469111, 32'h419a4c3a, 32'h40426e95, 32'h41866c79};
test_input[16616:16623] = '{32'h41b33200, 32'h42697b16, 32'hc227004f, 32'hc2aa2ebd, 32'hc1190104, 32'h3e55100d, 32'hc2859607, 32'h41212c19};
test_output[16616:16623] = '{32'h41b33200, 32'h42697b16, 32'h0, 32'h0, 32'h0, 32'h3e55100d, 32'h0, 32'h41212c19};
test_input[16624:16631] = '{32'h4229666c, 32'h42b73829, 32'h42aecea6, 32'h427e4950, 32'h425878d2, 32'hc182e6d9, 32'hc25bac14, 32'h41889b26};
test_output[16624:16631] = '{32'h4229666c, 32'h42b73829, 32'h42aecea6, 32'h427e4950, 32'h425878d2, 32'h0, 32'h0, 32'h41889b26};
test_input[16632:16639] = '{32'hc29f3796, 32'hc269cfaa, 32'h4293c76c, 32'h426411cf, 32'h417ca313, 32'hc15744cb, 32'h42b50378, 32'hc265b5be};
test_output[16632:16639] = '{32'h0, 32'h0, 32'h4293c76c, 32'h426411cf, 32'h417ca313, 32'h0, 32'h42b50378, 32'h0};
test_input[16640:16647] = '{32'h4231644a, 32'hc229dd1a, 32'hc2a1e3dd, 32'hc26a59cd, 32'h4223b343, 32'hc1309830, 32'hc2b66f6f, 32'hc2a38f87};
test_output[16640:16647] = '{32'h4231644a, 32'h0, 32'h0, 32'h0, 32'h4223b343, 32'h0, 32'h0, 32'h0};
test_input[16648:16655] = '{32'h411c1d42, 32'hc188aabb, 32'h42b50d32, 32'hbf548c07, 32'h41abbe10, 32'hc2c3c749, 32'h4253ce3a, 32'h4204d794};
test_output[16648:16655] = '{32'h411c1d42, 32'h0, 32'h42b50d32, 32'h0, 32'h41abbe10, 32'h0, 32'h4253ce3a, 32'h4204d794};
test_input[16656:16663] = '{32'h420c0885, 32'h425a4382, 32'hc1e680ea, 32'hc214a0c4, 32'hc0fb87a3, 32'hc1ffe9d5, 32'hc19cab7c, 32'h4256cd2c};
test_output[16656:16663] = '{32'h420c0885, 32'h425a4382, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4256cd2c};
test_input[16664:16671] = '{32'hc2165c94, 32'hc2968edd, 32'hc25b476b, 32'hc16b179e, 32'h42bc55ce, 32'hc221fdd4, 32'h42b9b80b, 32'h4273ab9b};
test_output[16664:16671] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42bc55ce, 32'h0, 32'h42b9b80b, 32'h4273ab9b};
test_input[16672:16679] = '{32'h42618774, 32'hbe61145d, 32'h41887a4b, 32'h4214cea6, 32'hc18fa4aa, 32'h425bffe5, 32'hc22d1e65, 32'hc23b2941};
test_output[16672:16679] = '{32'h42618774, 32'h0, 32'h41887a4b, 32'h4214cea6, 32'h0, 32'h425bffe5, 32'h0, 32'h0};
test_input[16680:16687] = '{32'hc2a16763, 32'hc14ad287, 32'h40edaa1a, 32'h420e7f9d, 32'h41ec2bd1, 32'h41f1631e, 32'hc274cd4c, 32'hc25d64ea};
test_output[16680:16687] = '{32'h0, 32'h0, 32'h40edaa1a, 32'h420e7f9d, 32'h41ec2bd1, 32'h41f1631e, 32'h0, 32'h0};
test_input[16688:16695] = '{32'h4282b421, 32'h42326257, 32'hc2b020b3, 32'h415405cb, 32'hc2b093a8, 32'h429fe483, 32'h429056cd, 32'h429a0e4d};
test_output[16688:16695] = '{32'h4282b421, 32'h42326257, 32'h0, 32'h415405cb, 32'h0, 32'h429fe483, 32'h429056cd, 32'h429a0e4d};
test_input[16696:16703] = '{32'h425b411f, 32'hc2504a2d, 32'hc2315d23, 32'h4127fd7a, 32'h41885fd0, 32'hc2b2bb38, 32'hc260a687, 32'hc206d2e3};
test_output[16696:16703] = '{32'h425b411f, 32'h0, 32'h0, 32'h4127fd7a, 32'h41885fd0, 32'h0, 32'h0, 32'h0};
test_input[16704:16711] = '{32'hc233aa5f, 32'hc29cecf4, 32'h420c1c7c, 32'hc2b8ebaa, 32'hc241038e, 32'hc12f8564, 32'h42ae5b2d, 32'hc2c4989d};
test_output[16704:16711] = '{32'h0, 32'h0, 32'h420c1c7c, 32'h0, 32'h0, 32'h0, 32'h42ae5b2d, 32'h0};
test_input[16712:16719] = '{32'h41f10e44, 32'h4281e450, 32'h422cb173, 32'hc2a304ce, 32'h424fb51a, 32'h42a96d95, 32'hc2377218, 32'hc21e39b6};
test_output[16712:16719] = '{32'h41f10e44, 32'h4281e450, 32'h422cb173, 32'h0, 32'h424fb51a, 32'h42a96d95, 32'h0, 32'h0};
test_input[16720:16727] = '{32'hc1dff07c, 32'h418d32fb, 32'h40a77646, 32'hc2adfbe7, 32'h42967297, 32'hc210a3d7, 32'h41f2add9, 32'hc2010a82};
test_output[16720:16727] = '{32'h0, 32'h418d32fb, 32'h40a77646, 32'h0, 32'h42967297, 32'h0, 32'h41f2add9, 32'h0};
test_input[16728:16735] = '{32'hc0b9255c, 32'h42322409, 32'hc1ad22af, 32'h429c3de4, 32'h42726304, 32'hc0e9f4b3, 32'hc2c44851, 32'hc2be643b};
test_output[16728:16735] = '{32'h0, 32'h42322409, 32'h0, 32'h429c3de4, 32'h42726304, 32'h0, 32'h0, 32'h0};
test_input[16736:16743] = '{32'h4242d73e, 32'h42955279, 32'hc1a4161f, 32'hc2c7875f, 32'hc272cb5c, 32'h4256df6f, 32'h428842d1, 32'hc29ad4c0};
test_output[16736:16743] = '{32'h4242d73e, 32'h42955279, 32'h0, 32'h0, 32'h0, 32'h4256df6f, 32'h428842d1, 32'h0};
test_input[16744:16751] = '{32'hc271850a, 32'h4247a1f9, 32'h40c40acd, 32'hbff38e10, 32'hc1929c65, 32'hc2085b29, 32'h428b45f8, 32'hc0e2da58};
test_output[16744:16751] = '{32'h0, 32'h4247a1f9, 32'h40c40acd, 32'h0, 32'h0, 32'h0, 32'h428b45f8, 32'h0};
test_input[16752:16759] = '{32'hc2b6fe66, 32'hc2a95442, 32'h4291561e, 32'h42acbd35, 32'hc296582e, 32'h42205f3e, 32'h413e9bd9, 32'hc23d216b};
test_output[16752:16759] = '{32'h0, 32'h0, 32'h4291561e, 32'h42acbd35, 32'h0, 32'h42205f3e, 32'h413e9bd9, 32'h0};
test_input[16760:16767] = '{32'h4256e6d5, 32'h420a020f, 32'h4212e0d6, 32'hc0ad44ea, 32'hc22e11cc, 32'hc191ccde, 32'h427a1741, 32'h42c7ea16};
test_output[16760:16767] = '{32'h4256e6d5, 32'h420a020f, 32'h4212e0d6, 32'h0, 32'h0, 32'h0, 32'h427a1741, 32'h42c7ea16};
test_input[16768:16775] = '{32'hc24f0806, 32'h4283f4c0, 32'hc1dddf3e, 32'hc2984d5b, 32'hc284f057, 32'hc20c41d4, 32'hc295861b, 32'h42a21916};
test_output[16768:16775] = '{32'h0, 32'h4283f4c0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a21916};
test_input[16776:16783] = '{32'h42938c9f, 32'h42654115, 32'h420fa8c7, 32'hc2bde60b, 32'h42bdbd46, 32'h41569f3e, 32'h418730a5, 32'hc0b4b82b};
test_output[16776:16783] = '{32'h42938c9f, 32'h42654115, 32'h420fa8c7, 32'h0, 32'h42bdbd46, 32'h41569f3e, 32'h418730a5, 32'h0};
test_input[16784:16791] = '{32'hc29d59a3, 32'h41713555, 32'hc198120f, 32'hc2645827, 32'hc291f16a, 32'h42604eeb, 32'h428dbbeb, 32'hc1f68099};
test_output[16784:16791] = '{32'h0, 32'h41713555, 32'h0, 32'h0, 32'h0, 32'h42604eeb, 32'h428dbbeb, 32'h0};
test_input[16792:16799] = '{32'h4295bfd5, 32'hc1f21e49, 32'hc249f5d1, 32'h4239e99c, 32'hc263d745, 32'h42779c43, 32'h429f9f4b, 32'h4094e3ab};
test_output[16792:16799] = '{32'h4295bfd5, 32'h0, 32'h0, 32'h4239e99c, 32'h0, 32'h42779c43, 32'h429f9f4b, 32'h4094e3ab};
test_input[16800:16807] = '{32'h4294ab95, 32'hc2c251c6, 32'h4213b1b2, 32'hc26f1155, 32'hc1f8be82, 32'h4280b143, 32'hc2093d57, 32'hc1c33fc2};
test_output[16800:16807] = '{32'h4294ab95, 32'h0, 32'h4213b1b2, 32'h0, 32'h0, 32'h4280b143, 32'h0, 32'h0};
test_input[16808:16815] = '{32'h4212b377, 32'hc1903a60, 32'h428209bd, 32'hc2695a3a, 32'hc29a7322, 32'hc0d8ab45, 32'h429d1627, 32'h42c59cfa};
test_output[16808:16815] = '{32'h4212b377, 32'h0, 32'h428209bd, 32'h0, 32'h0, 32'h0, 32'h429d1627, 32'h42c59cfa};
test_input[16816:16823] = '{32'h40aa2b7e, 32'hc1d5bc53, 32'hc25caf79, 32'h427e5224, 32'hc0c90919, 32'h40ce9adf, 32'h42583dd0, 32'h4264e205};
test_output[16816:16823] = '{32'h40aa2b7e, 32'h0, 32'h0, 32'h427e5224, 32'h0, 32'h40ce9adf, 32'h42583dd0, 32'h4264e205};
test_input[16824:16831] = '{32'hc233ca62, 32'hc1bacbe6, 32'h427d39b2, 32'h424cf2b7, 32'h40c6c758, 32'h40558dbc, 32'h42b8990f, 32'h415035c4};
test_output[16824:16831] = '{32'h0, 32'h0, 32'h427d39b2, 32'h424cf2b7, 32'h40c6c758, 32'h40558dbc, 32'h42b8990f, 32'h415035c4};
test_input[16832:16839] = '{32'hc28b829f, 32'h41e8fbf3, 32'hc2b00f93, 32'hc28663e0, 32'hc15a0f39, 32'hc2b39008, 32'hc21ac7c1, 32'h4211e96e};
test_output[16832:16839] = '{32'h0, 32'h41e8fbf3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4211e96e};
test_input[16840:16847] = '{32'hc2ba4edd, 32'h41932fbd, 32'hc28814b2, 32'h4111a8fe, 32'h4232ef33, 32'hc2b10c3d, 32'h428ba279, 32'h41c2967f};
test_output[16840:16847] = '{32'h0, 32'h41932fbd, 32'h0, 32'h4111a8fe, 32'h4232ef33, 32'h0, 32'h428ba279, 32'h41c2967f};
test_input[16848:16855] = '{32'hc2b7091d, 32'h41812c6d, 32'hc119b0ee, 32'h4279b61f, 32'h42aef4f3, 32'hc29dcc28, 32'h426f731b, 32'hc25f3560};
test_output[16848:16855] = '{32'h0, 32'h41812c6d, 32'h0, 32'h4279b61f, 32'h42aef4f3, 32'h0, 32'h426f731b, 32'h0};
test_input[16856:16863] = '{32'hc18b2b8a, 32'h4165cc66, 32'hc0c833eb, 32'h429a9c23, 32'h422276cc, 32'hc2ae5897, 32'h421124bd, 32'h42bf6ea9};
test_output[16856:16863] = '{32'h0, 32'h4165cc66, 32'h0, 32'h429a9c23, 32'h422276cc, 32'h0, 32'h421124bd, 32'h42bf6ea9};
test_input[16864:16871] = '{32'hc2791160, 32'h4295fd5b, 32'hc1813f66, 32'h41d5c1ad, 32'h4220759c, 32'hc125f760, 32'hc156811f, 32'h421d7b1f};
test_output[16864:16871] = '{32'h0, 32'h4295fd5b, 32'h0, 32'h41d5c1ad, 32'h4220759c, 32'h0, 32'h0, 32'h421d7b1f};
test_input[16872:16879] = '{32'h3fbd065d, 32'h4262a9b6, 32'h428f5f66, 32'hc1927e98, 32'hc26561aa, 32'hc289faa3, 32'h42199220, 32'h4202b204};
test_output[16872:16879] = '{32'h3fbd065d, 32'h4262a9b6, 32'h428f5f66, 32'h0, 32'h0, 32'h0, 32'h42199220, 32'h4202b204};
test_input[16880:16887] = '{32'hc0d91dc0, 32'h429ebf32, 32'h42c5e01f, 32'hc2b9122b, 32'h4205df6e, 32'hc197be3c, 32'hc242e8e8, 32'h42bc1bef};
test_output[16880:16887] = '{32'h0, 32'h429ebf32, 32'h42c5e01f, 32'h0, 32'h4205df6e, 32'h0, 32'h0, 32'h42bc1bef};
test_input[16888:16895] = '{32'hc262dc88, 32'hc1f2b4f2, 32'hc256a41a, 32'hc19dcfd3, 32'hc222bb52, 32'h4246ec73, 32'h426c773b, 32'h41c3ea2a};
test_output[16888:16895] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4246ec73, 32'h426c773b, 32'h41c3ea2a};
test_input[16896:16903] = '{32'hc14319fd, 32'h428b483b, 32'hc280e9c6, 32'hc165bdd0, 32'hc20ea92d, 32'h4248c089, 32'h42bd6784, 32'h42228560};
test_output[16896:16903] = '{32'h0, 32'h428b483b, 32'h0, 32'h0, 32'h0, 32'h4248c089, 32'h42bd6784, 32'h42228560};
test_input[16904:16911] = '{32'h421df59b, 32'h41e8384d, 32'h4273a3e2, 32'hc2bf0af8, 32'h41cdecba, 32'h422335a8, 32'h42b09954, 32'hc27cbe2c};
test_output[16904:16911] = '{32'h421df59b, 32'h41e8384d, 32'h4273a3e2, 32'h0, 32'h41cdecba, 32'h422335a8, 32'h42b09954, 32'h0};
test_input[16912:16919] = '{32'h42b90dbb, 32'hc299834a, 32'h41b98194, 32'h42a731b0, 32'h41326944, 32'h41de1873, 32'hc1115788, 32'hc1acd78a};
test_output[16912:16919] = '{32'h42b90dbb, 32'h0, 32'h41b98194, 32'h42a731b0, 32'h41326944, 32'h41de1873, 32'h0, 32'h0};
test_input[16920:16927] = '{32'hc18ca17b, 32'hc16e3082, 32'hc28a06a9, 32'h426d0fbc, 32'hc28e4c81, 32'h420b2e61, 32'hc238bf6d, 32'h409481fc};
test_output[16920:16927] = '{32'h0, 32'h0, 32'h0, 32'h426d0fbc, 32'h0, 32'h420b2e61, 32'h0, 32'h409481fc};
test_input[16928:16935] = '{32'h421b66f3, 32'h412ac62d, 32'hc28f04a3, 32'h41b5375e, 32'hc1a60711, 32'h407084b7, 32'h4186906b, 32'hc28672a8};
test_output[16928:16935] = '{32'h421b66f3, 32'h412ac62d, 32'h0, 32'h41b5375e, 32'h0, 32'h407084b7, 32'h4186906b, 32'h0};
test_input[16936:16943] = '{32'h423fa4ac, 32'hc2a833ae, 32'h42bd7583, 32'hc2c57306, 32'hc11faa86, 32'hc1afd4a6, 32'h413ac3a7, 32'hc0860237};
test_output[16936:16943] = '{32'h423fa4ac, 32'h0, 32'h42bd7583, 32'h0, 32'h0, 32'h0, 32'h413ac3a7, 32'h0};
test_input[16944:16951] = '{32'hc20872fa, 32'h4224ae46, 32'h40717b2d, 32'h41861583, 32'hc1e0e3ec, 32'h42546239, 32'hc2b84b03, 32'hc2931c00};
test_output[16944:16951] = '{32'h0, 32'h4224ae46, 32'h40717b2d, 32'h41861583, 32'h0, 32'h42546239, 32'h0, 32'h0};
test_input[16952:16959] = '{32'h4284a2ed, 32'hc1b5a617, 32'h42c7a30f, 32'hc2a158ca, 32'hbffb8578, 32'h42476a10, 32'hc288f770, 32'hc12438a9};
test_output[16952:16959] = '{32'h4284a2ed, 32'h0, 32'h42c7a30f, 32'h0, 32'h0, 32'h42476a10, 32'h0, 32'h0};
test_input[16960:16967] = '{32'h42a5b183, 32'hc2b01cba, 32'hc22250b0, 32'h42bb2c68, 32'h4125f25f, 32'h42ae9627, 32'hc29dc3ef, 32'h4286881c};
test_output[16960:16967] = '{32'h42a5b183, 32'h0, 32'h0, 32'h42bb2c68, 32'h4125f25f, 32'h42ae9627, 32'h0, 32'h4286881c};
test_input[16968:16975] = '{32'h4239e632, 32'hc232bbd4, 32'hc1ef66ad, 32'h41c132ed, 32'hc13f5141, 32'hc1e02a6f, 32'hc19f7481, 32'h42af6f03};
test_output[16968:16975] = '{32'h4239e632, 32'h0, 32'h0, 32'h41c132ed, 32'h0, 32'h0, 32'h0, 32'h42af6f03};
test_input[16976:16983] = '{32'hc2a21b9e, 32'hc250d606, 32'h4250d4d6, 32'h42255d2b, 32'hc29c1557, 32'h4118e501, 32'hc0727dfb, 32'h42a879cb};
test_output[16976:16983] = '{32'h0, 32'h0, 32'h4250d4d6, 32'h42255d2b, 32'h0, 32'h4118e501, 32'h0, 32'h42a879cb};
test_input[16984:16991] = '{32'hc14c677e, 32'h42b1643b, 32'h418df890, 32'h42934048, 32'hc291f875, 32'h41f3faae, 32'hc121eeb4, 32'hc284a4ef};
test_output[16984:16991] = '{32'h0, 32'h42b1643b, 32'h418df890, 32'h42934048, 32'h0, 32'h41f3faae, 32'h0, 32'h0};
test_input[16992:16999] = '{32'h41b477be, 32'h42a1c815, 32'hc22d70fd, 32'hc2ab9bcd, 32'hc2c48d1f, 32'h429d02d0, 32'hc24e1d89, 32'h42a92358};
test_output[16992:16999] = '{32'h41b477be, 32'h42a1c815, 32'h0, 32'h0, 32'h0, 32'h429d02d0, 32'h0, 32'h42a92358};
test_input[17000:17007] = '{32'hc202b60e, 32'hc29e8c3d, 32'h4298c641, 32'h425b0fcf, 32'hc28ad86c, 32'h42b95e16, 32'hc1113c9e, 32'hc2b07edf};
test_output[17000:17007] = '{32'h0, 32'h0, 32'h4298c641, 32'h425b0fcf, 32'h0, 32'h42b95e16, 32'h0, 32'h0};
test_input[17008:17015] = '{32'h42bd4011, 32'h42417bbc, 32'h41f90fad, 32'h426d6d33, 32'h4157fb24, 32'h41e03bce, 32'hc20c6cfd, 32'h42266503};
test_output[17008:17015] = '{32'h42bd4011, 32'h42417bbc, 32'h41f90fad, 32'h426d6d33, 32'h4157fb24, 32'h41e03bce, 32'h0, 32'h42266503};
test_input[17016:17023] = '{32'hc116fbec, 32'hc176dcf6, 32'h41e4b89c, 32'h42a989d3, 32'h40de682b, 32'h40f4158c, 32'hc29d7e3c, 32'h42b56db0};
test_output[17016:17023] = '{32'h0, 32'h0, 32'h41e4b89c, 32'h42a989d3, 32'h40de682b, 32'h40f4158c, 32'h0, 32'h42b56db0};
test_input[17024:17031] = '{32'hc26c5107, 32'hc256d4f1, 32'hc0dbd954, 32'h4042e4e8, 32'hc0d710a3, 32'hc2ae5b1c, 32'h42728900, 32'hc26fc053};
test_output[17024:17031] = '{32'h0, 32'h0, 32'h0, 32'h4042e4e8, 32'h0, 32'h0, 32'h42728900, 32'h0};
test_input[17032:17039] = '{32'hc2369239, 32'hc1c57717, 32'h3f6228a6, 32'h41d2dd21, 32'hc2744f17, 32'hc2b50e54, 32'h426947a1, 32'h4238a9ba};
test_output[17032:17039] = '{32'h0, 32'h0, 32'h3f6228a6, 32'h41d2dd21, 32'h0, 32'h0, 32'h426947a1, 32'h4238a9ba};
test_input[17040:17047] = '{32'hc2506dd8, 32'h42b831e3, 32'hc2a61088, 32'hc2b23998, 32'h420e6252, 32'h41c39443, 32'hc298c307, 32'h41a7ff0f};
test_output[17040:17047] = '{32'h0, 32'h42b831e3, 32'h0, 32'h0, 32'h420e6252, 32'h41c39443, 32'h0, 32'h41a7ff0f};
test_input[17048:17055] = '{32'h421be5e7, 32'h42987b07, 32'h42791424, 32'h4294f29d, 32'h42bc5ad0, 32'hc2386100, 32'h419f8847, 32'h42779cad};
test_output[17048:17055] = '{32'h421be5e7, 32'h42987b07, 32'h42791424, 32'h4294f29d, 32'h42bc5ad0, 32'h0, 32'h419f8847, 32'h42779cad};
test_input[17056:17063] = '{32'h41adbc5c, 32'hc1d0fec2, 32'h4299b450, 32'h4092739d, 32'h42af4940, 32'hc2c050d7, 32'h42848c94, 32'hc2a32a78};
test_output[17056:17063] = '{32'h41adbc5c, 32'h0, 32'h4299b450, 32'h4092739d, 32'h42af4940, 32'h0, 32'h42848c94, 32'h0};
test_input[17064:17071] = '{32'hc0220af8, 32'h42720fa2, 32'hc2ae82e2, 32'h40a4a6aa, 32'h427d9be2, 32'h42973547, 32'hc1d50578, 32'h41ea7e2a};
test_output[17064:17071] = '{32'h0, 32'h42720fa2, 32'h0, 32'h40a4a6aa, 32'h427d9be2, 32'h42973547, 32'h0, 32'h41ea7e2a};
test_input[17072:17079] = '{32'h41e4057e, 32'hc28bf244, 32'h41b6ecfd, 32'hc216f657, 32'hc23d6e70, 32'h4207cf1d, 32'hc1b22aeb, 32'h4292af6a};
test_output[17072:17079] = '{32'h41e4057e, 32'h0, 32'h41b6ecfd, 32'h0, 32'h0, 32'h4207cf1d, 32'h0, 32'h4292af6a};
test_input[17080:17087] = '{32'h424c8843, 32'h42976be6, 32'hc0c4bfff, 32'hc2a48afd, 32'h425e2e45, 32'hc081ef77, 32'hc17b1220, 32'hc24fb576};
test_output[17080:17087] = '{32'h424c8843, 32'h42976be6, 32'h0, 32'h0, 32'h425e2e45, 32'h0, 32'h0, 32'h0};
test_input[17088:17095] = '{32'h41871d73, 32'h41a1f556, 32'hc20e797b, 32'hc26c4271, 32'h4087c55f, 32'h4247270f, 32'hc2374639, 32'hc263ff03};
test_output[17088:17095] = '{32'h41871d73, 32'h41a1f556, 32'h0, 32'h0, 32'h4087c55f, 32'h4247270f, 32'h0, 32'h0};
test_input[17096:17103] = '{32'h412427f7, 32'hc1807851, 32'h40eba908, 32'hc26491ea, 32'h418ad4ab, 32'hc283c0a5, 32'h41f68281, 32'h42befc0b};
test_output[17096:17103] = '{32'h412427f7, 32'h0, 32'h40eba908, 32'h0, 32'h418ad4ab, 32'h0, 32'h41f68281, 32'h42befc0b};
test_input[17104:17111] = '{32'h429b3750, 32'hc0b7c55e, 32'hc17fe7f1, 32'hc1309d7e, 32'hc1e8f31b, 32'h41ce5cbf, 32'hc1b2c846, 32'h42bbdde1};
test_output[17104:17111] = '{32'h429b3750, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ce5cbf, 32'h0, 32'h42bbdde1};
test_input[17112:17119] = '{32'h42afc99c, 32'hc29a633f, 32'hc22b14b0, 32'h41f10ad9, 32'h42ac8798, 32'hc257440c, 32'hc12c4d1e, 32'h42a06dc0};
test_output[17112:17119] = '{32'h42afc99c, 32'h0, 32'h0, 32'h41f10ad9, 32'h42ac8798, 32'h0, 32'h0, 32'h42a06dc0};
test_input[17120:17127] = '{32'h429af45c, 32'h3f7a03db, 32'h41fff3de, 32'h42b65a99, 32'h411fd9b6, 32'h411b6d62, 32'h40c0a241, 32'h4295a5bb};
test_output[17120:17127] = '{32'h429af45c, 32'h3f7a03db, 32'h41fff3de, 32'h42b65a99, 32'h411fd9b6, 32'h411b6d62, 32'h40c0a241, 32'h4295a5bb};
test_input[17128:17135] = '{32'h42303ce0, 32'h418f6599, 32'h42b0ae3d, 32'h428a759f, 32'hc22aebdd, 32'hc21a9519, 32'h3f046ebe, 32'hc20fe30d};
test_output[17128:17135] = '{32'h42303ce0, 32'h418f6599, 32'h42b0ae3d, 32'h428a759f, 32'h0, 32'h0, 32'h3f046ebe, 32'h0};
test_input[17136:17143] = '{32'hc1b02ffb, 32'hc192db73, 32'h421e1805, 32'hc1bf8373, 32'hc1aa4f67, 32'h417a35b8, 32'hc273dffb, 32'h426a5d5b};
test_output[17136:17143] = '{32'h0, 32'h0, 32'h421e1805, 32'h0, 32'h0, 32'h417a35b8, 32'h0, 32'h426a5d5b};
test_input[17144:17151] = '{32'h424069f2, 32'h42adb20d, 32'hc257776d, 32'h41d28447, 32'h419af38a, 32'hc0b512aa, 32'hc2a51aed, 32'h42139518};
test_output[17144:17151] = '{32'h424069f2, 32'h42adb20d, 32'h0, 32'h41d28447, 32'h419af38a, 32'h0, 32'h0, 32'h42139518};
test_input[17152:17159] = '{32'h42a5cfcd, 32'hc293992f, 32'h42957eae, 32'hc1a81090, 32'hc25b8867, 32'hc2153550, 32'hc22e7d4c, 32'hc20cd8fb};
test_output[17152:17159] = '{32'h42a5cfcd, 32'h0, 32'h42957eae, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[17160:17167] = '{32'hc1a3f404, 32'h422381e4, 32'h427b0ffe, 32'hc20f035b, 32'hbf269077, 32'h427c7d7c, 32'h4153f80a, 32'h42246571};
test_output[17160:17167] = '{32'h0, 32'h422381e4, 32'h427b0ffe, 32'h0, 32'h0, 32'h427c7d7c, 32'h4153f80a, 32'h42246571};
test_input[17168:17175] = '{32'h40917a99, 32'hc26d1d7e, 32'hc2c5647d, 32'hc2b9ce68, 32'hc29737e3, 32'h4230bc69, 32'hc1f41223, 32'h3ee98ba5};
test_output[17168:17175] = '{32'h40917a99, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4230bc69, 32'h0, 32'h3ee98ba5};
test_input[17176:17183] = '{32'h42b039a5, 32'h40979290, 32'h402fb2ee, 32'h4163d921, 32'h428194c3, 32'hc2697ecf, 32'hc28c5566, 32'h4295713a};
test_output[17176:17183] = '{32'h42b039a5, 32'h40979290, 32'h402fb2ee, 32'h4163d921, 32'h428194c3, 32'h0, 32'h0, 32'h4295713a};
test_input[17184:17191] = '{32'hc2c71515, 32'h4221705c, 32'h41215a99, 32'hc23fe5f1, 32'h4242d8d9, 32'hc28409d5, 32'h42814931, 32'h40b088ad};
test_output[17184:17191] = '{32'h0, 32'h4221705c, 32'h41215a99, 32'h0, 32'h4242d8d9, 32'h0, 32'h42814931, 32'h40b088ad};
test_input[17192:17199] = '{32'h42a221bd, 32'h41633297, 32'hc2bf4419, 32'h4209d4bf, 32'hc26d2613, 32'h42b57b33, 32'h424aa0f3, 32'h4275af2f};
test_output[17192:17199] = '{32'h42a221bd, 32'h41633297, 32'h0, 32'h4209d4bf, 32'h0, 32'h42b57b33, 32'h424aa0f3, 32'h4275af2f};
test_input[17200:17207] = '{32'h421ed2e7, 32'hc26692dd, 32'hc286a094, 32'h41c6d95d, 32'h40d995b0, 32'hc1d129a5, 32'h3f8b3e1e, 32'h422952bd};
test_output[17200:17207] = '{32'h421ed2e7, 32'h0, 32'h0, 32'h41c6d95d, 32'h40d995b0, 32'h0, 32'h3f8b3e1e, 32'h422952bd};
test_input[17208:17215] = '{32'hc2c460a6, 32'h4212086c, 32'h4241b666, 32'h417ddcd3, 32'hc15daf55, 32'h41837c9d, 32'h4289bf82, 32'h4276e659};
test_output[17208:17215] = '{32'h0, 32'h4212086c, 32'h4241b666, 32'h417ddcd3, 32'h0, 32'h41837c9d, 32'h4289bf82, 32'h4276e659};
test_input[17216:17223] = '{32'h424c9df1, 32'h429b3475, 32'hc27e850d, 32'hc2c1dc27, 32'h4097a71e, 32'hc23b9902, 32'h424f1687, 32'h4238d6d0};
test_output[17216:17223] = '{32'h424c9df1, 32'h429b3475, 32'h0, 32'h0, 32'h4097a71e, 32'h0, 32'h424f1687, 32'h4238d6d0};
test_input[17224:17231] = '{32'hc286d1e0, 32'hc2ae54a1, 32'hc24ce832, 32'h420106a3, 32'h42c34370, 32'hc27f5efc, 32'h4213c5fd, 32'hc258d733};
test_output[17224:17231] = '{32'h0, 32'h0, 32'h0, 32'h420106a3, 32'h42c34370, 32'h0, 32'h4213c5fd, 32'h0};
test_input[17232:17239] = '{32'hc2b80983, 32'h426837ad, 32'h42b262e4, 32'hc2a0221f, 32'hc2bb80a5, 32'h4274ff93, 32'h40e3d60d, 32'hc1828596};
test_output[17232:17239] = '{32'h0, 32'h426837ad, 32'h42b262e4, 32'h0, 32'h0, 32'h4274ff93, 32'h40e3d60d, 32'h0};
test_input[17240:17247] = '{32'hc28fdf7c, 32'h42b0e4b5, 32'hc28c8278, 32'h4200f428, 32'hc29312e5, 32'h4023ff4e, 32'hc05e07c9, 32'hc27e68dc};
test_output[17240:17247] = '{32'h0, 32'h42b0e4b5, 32'h0, 32'h4200f428, 32'h0, 32'h4023ff4e, 32'h0, 32'h0};
test_input[17248:17255] = '{32'hc1c0b6cf, 32'hc236f798, 32'hc2290b78, 32'hc2c5cba0, 32'hc10f1ed3, 32'h4276d872, 32'h42a2def9, 32'hc2b8c656};
test_output[17248:17255] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4276d872, 32'h42a2def9, 32'h0};
test_input[17256:17263] = '{32'h426a1a40, 32'h40f2b6c4, 32'hc21adc24, 32'h42a60f91, 32'hc1d9c6d8, 32'h429b00d8, 32'hc1dfb293, 32'hc08cb6a9};
test_output[17256:17263] = '{32'h426a1a40, 32'h40f2b6c4, 32'h0, 32'h42a60f91, 32'h0, 32'h429b00d8, 32'h0, 32'h0};
test_input[17264:17271] = '{32'hc228daa4, 32'h42bedcd0, 32'h420fe94b, 32'hc1aaf44f, 32'h42baafad, 32'hc1d75fd9, 32'h42a45881, 32'hc21950b5};
test_output[17264:17271] = '{32'h0, 32'h42bedcd0, 32'h420fe94b, 32'h0, 32'h42baafad, 32'h0, 32'h42a45881, 32'h0};
test_input[17272:17279] = '{32'h4269dd57, 32'h42b8f4d1, 32'hc2c21996, 32'hc2506012, 32'hc2af1abc, 32'hc2911d47, 32'hc238dd0f, 32'h42bd0a16};
test_output[17272:17279] = '{32'h4269dd57, 32'h42b8f4d1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bd0a16};
test_input[17280:17287] = '{32'h41f92d79, 32'h42602c6d, 32'h423a8c06, 32'hc213e317, 32'h420dee94, 32'h42bfe7c1, 32'h42a95fd5, 32'h423c47eb};
test_output[17280:17287] = '{32'h41f92d79, 32'h42602c6d, 32'h423a8c06, 32'h0, 32'h420dee94, 32'h42bfe7c1, 32'h42a95fd5, 32'h423c47eb};
test_input[17288:17295] = '{32'hc2afcfc7, 32'hc1dd7258, 32'hc1dd69ba, 32'h4063ef79, 32'h4292704d, 32'h4270f1ca, 32'hc2b829d1, 32'hc29abd43};
test_output[17288:17295] = '{32'h0, 32'h0, 32'h0, 32'h4063ef79, 32'h4292704d, 32'h4270f1ca, 32'h0, 32'h0};
test_input[17296:17303] = '{32'hc18577d4, 32'hc28262f8, 32'hbfcea4c4, 32'hc2524f24, 32'hc2c5c942, 32'hc1fbb011, 32'hc23321b2, 32'h41fd1bdd};
test_output[17296:17303] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41fd1bdd};
test_input[17304:17311] = '{32'h41f780eb, 32'hc2787745, 32'hc1fc0ccf, 32'hc2138a46, 32'hc2393bf6, 32'h4243fc0a, 32'hc189c2cc, 32'h423a084e};
test_output[17304:17311] = '{32'h41f780eb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4243fc0a, 32'h0, 32'h423a084e};
test_input[17312:17319] = '{32'h429d124f, 32'h422b4de2, 32'h4125ac80, 32'h426f3928, 32'hc24ec55a, 32'h41b215d9, 32'h42804150, 32'h42231489};
test_output[17312:17319] = '{32'h429d124f, 32'h422b4de2, 32'h4125ac80, 32'h426f3928, 32'h0, 32'h41b215d9, 32'h42804150, 32'h42231489};
test_input[17320:17327] = '{32'hc2048573, 32'hc295af43, 32'hc2b5a88d, 32'hc273c5d2, 32'hc2b76e51, 32'hc29d4d39, 32'h421c9d7a, 32'h42a6aca0};
test_output[17320:17327] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h421c9d7a, 32'h42a6aca0};
test_input[17328:17335] = '{32'hc1b960d2, 32'h42b522a4, 32'h429de023, 32'h42a4b80c, 32'hc093aaa2, 32'h41e1456a, 32'hc26e15a9, 32'h421db54d};
test_output[17328:17335] = '{32'h0, 32'h42b522a4, 32'h429de023, 32'h42a4b80c, 32'h0, 32'h41e1456a, 32'h0, 32'h421db54d};
test_input[17336:17343] = '{32'hc130612e, 32'h407eac8d, 32'hc1c0944f, 32'hc25f9b1c, 32'h3fe0c586, 32'h417e3eea, 32'h42244642, 32'hc22f03ef};
test_output[17336:17343] = '{32'h0, 32'h407eac8d, 32'h0, 32'h0, 32'h3fe0c586, 32'h417e3eea, 32'h42244642, 32'h0};
test_input[17344:17351] = '{32'h42376828, 32'hc17b1068, 32'h42bffd2c, 32'hc1add3c1, 32'hc0cccbfe, 32'hc275b66f, 32'hc26a839f, 32'h4208fad4};
test_output[17344:17351] = '{32'h42376828, 32'h0, 32'h42bffd2c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4208fad4};
test_input[17352:17359] = '{32'h42785d1c, 32'h42105e0a, 32'hc1bf5593, 32'hc28c71d0, 32'hc223b3f8, 32'hc127e343, 32'h428d99e1, 32'hc2abac0a};
test_output[17352:17359] = '{32'h42785d1c, 32'h42105e0a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428d99e1, 32'h0};
test_input[17360:17367] = '{32'h41c103a7, 32'hc2688b96, 32'hc29df70f, 32'hc22f0e80, 32'hc23a6211, 32'h42ade151, 32'hc0279d8f, 32'h42b239e7};
test_output[17360:17367] = '{32'h41c103a7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ade151, 32'h0, 32'h42b239e7};
test_input[17368:17375] = '{32'h42c7d7c2, 32'h3f14c977, 32'h42ae9f10, 32'hc282fe42, 32'hc29f159a, 32'hc28b8246, 32'h410e4f43, 32'hc140887a};
test_output[17368:17375] = '{32'h42c7d7c2, 32'h3f14c977, 32'h42ae9f10, 32'h0, 32'h0, 32'h0, 32'h410e4f43, 32'h0};
test_input[17376:17383] = '{32'h4275668d, 32'h4293193a, 32'hc1c9f936, 32'hc299c068, 32'hc2ac7c3c, 32'hc29c621b, 32'hc25a599c, 32'hc25a16a7};
test_output[17376:17383] = '{32'h4275668d, 32'h4293193a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[17384:17391] = '{32'hc298dae7, 32'hc1be5151, 32'hc285ba11, 32'hc198dd5c, 32'hc2692c67, 32'hc2830976, 32'h40a2c501, 32'hc2bda546};
test_output[17384:17391] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40a2c501, 32'h0};
test_input[17392:17399] = '{32'h42a5cdd6, 32'hc10e8ebf, 32'h427fb4ba, 32'h41350cb2, 32'hc29ba859, 32'h42b628de, 32'hc22bd835, 32'hc25ed8be};
test_output[17392:17399] = '{32'h42a5cdd6, 32'h0, 32'h427fb4ba, 32'h41350cb2, 32'h0, 32'h42b628de, 32'h0, 32'h0};
test_input[17400:17407] = '{32'hc265d9a6, 32'h426d3ad1, 32'h428ab146, 32'hc2a0b279, 32'h429cff92, 32'hc2c3e0b1, 32'hc2338217, 32'hc2812332};
test_output[17400:17407] = '{32'h0, 32'h426d3ad1, 32'h428ab146, 32'h0, 32'h429cff92, 32'h0, 32'h0, 32'h0};
test_input[17408:17415] = '{32'h4235e75f, 32'hc28ddbac, 32'hc2b043bf, 32'hc09352d2, 32'h4271428c, 32'hc256ae3f, 32'hc1d6ae89, 32'hc20a181a};
test_output[17408:17415] = '{32'h4235e75f, 32'h0, 32'h0, 32'h0, 32'h4271428c, 32'h0, 32'h0, 32'h0};
test_input[17416:17423] = '{32'hc1ef50ac, 32'h424df0bd, 32'hc24dbb65, 32'h42ae1208, 32'hc29d4c8b, 32'h42b03f0f, 32'h42a3395b, 32'hc2309499};
test_output[17416:17423] = '{32'h0, 32'h424df0bd, 32'h0, 32'h42ae1208, 32'h0, 32'h42b03f0f, 32'h42a3395b, 32'h0};
test_input[17424:17431] = '{32'h41f65700, 32'hc2459a2c, 32'hc29acd72, 32'h429bd647, 32'h42b3a428, 32'h425cb836, 32'h42984710, 32'hc202f281};
test_output[17424:17431] = '{32'h41f65700, 32'h0, 32'h0, 32'h429bd647, 32'h42b3a428, 32'h425cb836, 32'h42984710, 32'h0};
test_input[17432:17439] = '{32'hc22e5a87, 32'h41873f16, 32'hc1f35fc9, 32'hc06c257e, 32'h42041d18, 32'hc2a90ad2, 32'hc2b8c058, 32'hc257932e};
test_output[17432:17439] = '{32'h0, 32'h41873f16, 32'h0, 32'h0, 32'h42041d18, 32'h0, 32'h0, 32'h0};
test_input[17440:17447] = '{32'hc08de943, 32'h4265a804, 32'hc27c56f2, 32'h427daed8, 32'hc22324ce, 32'hc2b5ce53, 32'h42613b8f, 32'hc29b6a6d};
test_output[17440:17447] = '{32'h0, 32'h4265a804, 32'h0, 32'h427daed8, 32'h0, 32'h0, 32'h42613b8f, 32'h0};
test_input[17448:17455] = '{32'h426a4831, 32'h42c2e047, 32'h42b29df2, 32'hc21b4503, 32'hc24159f5, 32'h42c2e645, 32'h42921b91, 32'hc2a02050};
test_output[17448:17455] = '{32'h426a4831, 32'h42c2e047, 32'h42b29df2, 32'h0, 32'h0, 32'h42c2e645, 32'h42921b91, 32'h0};
test_input[17456:17463] = '{32'h429e176d, 32'hc285503e, 32'h420b17b8, 32'hc1962988, 32'hc0a75e6d, 32'h42638c79, 32'hc224e135, 32'hc1cd485f};
test_output[17456:17463] = '{32'h429e176d, 32'h0, 32'h420b17b8, 32'h0, 32'h0, 32'h42638c79, 32'h0, 32'h0};
test_input[17464:17471] = '{32'h42a53e56, 32'hc2aac7cb, 32'hc1f87aad, 32'hc19eb718, 32'h42712a3e, 32'h4267b84e, 32'h42ad77b2, 32'hc27bedc1};
test_output[17464:17471] = '{32'h42a53e56, 32'h0, 32'h0, 32'h0, 32'h42712a3e, 32'h4267b84e, 32'h42ad77b2, 32'h0};
test_input[17472:17479] = '{32'h424ae18a, 32'h41a3f177, 32'hc28ebf9a, 32'h42be74e0, 32'hc2a518a7, 32'h41bdf8d8, 32'h420c6b7b, 32'hc2756663};
test_output[17472:17479] = '{32'h424ae18a, 32'h41a3f177, 32'h0, 32'h42be74e0, 32'h0, 32'h41bdf8d8, 32'h420c6b7b, 32'h0};
test_input[17480:17487] = '{32'hc22d34b4, 32'h429fbe07, 32'hc1c77484, 32'h4186c381, 32'h41a3d703, 32'hc2054fd9, 32'h42345ee4, 32'hc24f79f2};
test_output[17480:17487] = '{32'h0, 32'h429fbe07, 32'h0, 32'h4186c381, 32'h41a3d703, 32'h0, 32'h42345ee4, 32'h0};
test_input[17488:17495] = '{32'h4281774d, 32'hc1cead1e, 32'hc1eb8e69, 32'hc0fae092, 32'hc2b73bc9, 32'hc20d490a, 32'hc27bdb97, 32'h4150da26};
test_output[17488:17495] = '{32'h4281774d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4150da26};
test_input[17496:17503] = '{32'hc2c7a176, 32'hc28dde50, 32'hc288d53a, 32'h42bdef04, 32'h418b5691, 32'hc26a7725, 32'h411080b2, 32'hc1dba4ea};
test_output[17496:17503] = '{32'h0, 32'h0, 32'h0, 32'h42bdef04, 32'h418b5691, 32'h0, 32'h411080b2, 32'h0};
test_input[17504:17511] = '{32'hc1bc5198, 32'hc2677e6a, 32'hc21bdeac, 32'h425566e2, 32'h42420c7a, 32'h428def4a, 32'hc2a7a09a, 32'h39ccc7bb};
test_output[17504:17511] = '{32'h0, 32'h0, 32'h0, 32'h425566e2, 32'h42420c7a, 32'h428def4a, 32'h0, 32'h39ccc7bb};
test_input[17512:17519] = '{32'h428567e9, 32'hc24785c3, 32'hc223e970, 32'hc18f15a9, 32'hc25afd09, 32'h40d63d6f, 32'hc2b2cc79, 32'h41ff7864};
test_output[17512:17519] = '{32'h428567e9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40d63d6f, 32'h0, 32'h41ff7864};
test_input[17520:17527] = '{32'h41f984b1, 32'hc1c86092, 32'h424dae0d, 32'h427183b2, 32'hc27621fb, 32'h42659d9b, 32'h4228b37c, 32'hc0210219};
test_output[17520:17527] = '{32'h41f984b1, 32'h0, 32'h424dae0d, 32'h427183b2, 32'h0, 32'h42659d9b, 32'h4228b37c, 32'h0};
test_input[17528:17535] = '{32'hc28eb099, 32'hc2a94f4e, 32'h429d45f9, 32'h4113d6ed, 32'h41c3b7d9, 32'hc24250d6, 32'h423b34a9, 32'h4268032b};
test_output[17528:17535] = '{32'h0, 32'h0, 32'h429d45f9, 32'h4113d6ed, 32'h41c3b7d9, 32'h0, 32'h423b34a9, 32'h4268032b};
test_input[17536:17543] = '{32'h42843f86, 32'hc2c1aaba, 32'hc2bf989d, 32'hc01eac60, 32'h41a0d060, 32'hc2a97121, 32'hc2c43abd, 32'h411667a7};
test_output[17536:17543] = '{32'h42843f86, 32'h0, 32'h0, 32'h0, 32'h41a0d060, 32'h0, 32'h0, 32'h411667a7};
test_input[17544:17551] = '{32'h42aaf479, 32'h41fb4e2e, 32'hc2c4fe45, 32'h42445550, 32'hc1aaf1ee, 32'h42365c03, 32'h42744a3b, 32'hc2155a3e};
test_output[17544:17551] = '{32'h42aaf479, 32'h41fb4e2e, 32'h0, 32'h42445550, 32'h0, 32'h42365c03, 32'h42744a3b, 32'h0};
test_input[17552:17559] = '{32'hc2531d87, 32'h41645953, 32'h416cfae0, 32'h4220a570, 32'h424328af, 32'h4247f8bd, 32'h421ebcf7, 32'h4180d449};
test_output[17552:17559] = '{32'h0, 32'h41645953, 32'h416cfae0, 32'h4220a570, 32'h424328af, 32'h4247f8bd, 32'h421ebcf7, 32'h4180d449};
test_input[17560:17567] = '{32'hc26152a8, 32'hc11c11b0, 32'h427d75fc, 32'hc2467d60, 32'h41b28977, 32'hc1a0cd4c, 32'h42066317, 32'hc258449a};
test_output[17560:17567] = '{32'h0, 32'h0, 32'h427d75fc, 32'h0, 32'h41b28977, 32'h0, 32'h42066317, 32'h0};
test_input[17568:17575] = '{32'h412599f5, 32'hc091c31e, 32'h41494b81, 32'h41d4c7c5, 32'h41ebdd8d, 32'hc1e9a3c4, 32'h42c08f09, 32'h425682e7};
test_output[17568:17575] = '{32'h412599f5, 32'h0, 32'h41494b81, 32'h41d4c7c5, 32'h41ebdd8d, 32'h0, 32'h42c08f09, 32'h425682e7};
test_input[17576:17583] = '{32'h42bacb72, 32'hc2b93c69, 32'hc2006d63, 32'hc2328d1a, 32'hc11df65b, 32'hc1a37a8c, 32'h42b4b712, 32'h42a92557};
test_output[17576:17583] = '{32'h42bacb72, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b4b712, 32'h42a92557};
test_input[17584:17591] = '{32'hc1849dc8, 32'hc23af0f9, 32'h42868040, 32'h4290d169, 32'hc2345518, 32'hc26c5a48, 32'h41c78e04, 32'hc17ac484};
test_output[17584:17591] = '{32'h0, 32'h0, 32'h42868040, 32'h4290d169, 32'h0, 32'h0, 32'h41c78e04, 32'h0};
test_input[17592:17599] = '{32'h4293e1fd, 32'hc1cfa27f, 32'hc194548b, 32'hc23bd7b4, 32'hc1d125c0, 32'hc2b5ec67, 32'h42c4ddf5, 32'hc0b0d3c2};
test_output[17592:17599] = '{32'h4293e1fd, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c4ddf5, 32'h0};
test_input[17600:17607] = '{32'h42ba2511, 32'h4284cab6, 32'h4130222f, 32'hc276e552, 32'h422afeed, 32'hc2bff4c6, 32'h40a55977, 32'h428cf0e5};
test_output[17600:17607] = '{32'h42ba2511, 32'h4284cab6, 32'h4130222f, 32'h0, 32'h422afeed, 32'h0, 32'h40a55977, 32'h428cf0e5};
test_input[17608:17615] = '{32'h42432a29, 32'hc28dd42d, 32'h42b7a906, 32'h42aa6a9e, 32'h4263dd63, 32'h421d20c4, 32'h427f0cc7, 32'h4240ee93};
test_output[17608:17615] = '{32'h42432a29, 32'h0, 32'h42b7a906, 32'h42aa6a9e, 32'h4263dd63, 32'h421d20c4, 32'h427f0cc7, 32'h4240ee93};
test_input[17616:17623] = '{32'h4192fdbb, 32'h42c475fa, 32'hc0c24768, 32'h42613e96, 32'hc29ae620, 32'hc2b4e804, 32'h4202a3e5, 32'h42122dc7};
test_output[17616:17623] = '{32'h4192fdbb, 32'h42c475fa, 32'h0, 32'h42613e96, 32'h0, 32'h0, 32'h4202a3e5, 32'h42122dc7};
test_input[17624:17631] = '{32'h421306be, 32'hc1e6c79b, 32'hc294cd9a, 32'h42b83752, 32'h41918c31, 32'h42480edc, 32'h40f0f693, 32'h42927224};
test_output[17624:17631] = '{32'h421306be, 32'h0, 32'h0, 32'h42b83752, 32'h41918c31, 32'h42480edc, 32'h40f0f693, 32'h42927224};
test_input[17632:17639] = '{32'h423fe91c, 32'h429b657a, 32'h42bfbbac, 32'h41c64c3b, 32'h4275387b, 32'h428a6790, 32'hc285517a, 32'h429fbc7a};
test_output[17632:17639] = '{32'h423fe91c, 32'h429b657a, 32'h42bfbbac, 32'h41c64c3b, 32'h4275387b, 32'h428a6790, 32'h0, 32'h429fbc7a};
test_input[17640:17647] = '{32'hc1da1e7e, 32'h41cb3a93, 32'hc2c79df0, 32'hc28c67d9, 32'h41f0f56f, 32'hc194eb8d, 32'h42ad8d86, 32'hc1a05ea8};
test_output[17640:17647] = '{32'h0, 32'h41cb3a93, 32'h0, 32'h0, 32'h41f0f56f, 32'h0, 32'h42ad8d86, 32'h0};
test_input[17648:17655] = '{32'hc29f896f, 32'h42a5e91e, 32'hc29e3036, 32'hc28e0618, 32'hc28218fd, 32'hc235ab19, 32'h427a20a5, 32'h4231e420};
test_output[17648:17655] = '{32'h0, 32'h42a5e91e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427a20a5, 32'h4231e420};
test_input[17656:17663] = '{32'h4270ae8c, 32'h4291bb48, 32'h421f08a9, 32'h428ece9d, 32'h42b5aa45, 32'h4201b59d, 32'h420b5530, 32'h4126f53e};
test_output[17656:17663] = '{32'h4270ae8c, 32'h4291bb48, 32'h421f08a9, 32'h428ece9d, 32'h42b5aa45, 32'h4201b59d, 32'h420b5530, 32'h4126f53e};
test_input[17664:17671] = '{32'h4276d647, 32'h4266790f, 32'hc191cd92, 32'hc0cf1424, 32'hc18a7786, 32'hc208608a, 32'h42baf334, 32'hc2798d04};
test_output[17664:17671] = '{32'h4276d647, 32'h4266790f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42baf334, 32'h0};
test_input[17672:17679] = '{32'h420d562e, 32'hc2933d98, 32'h421836fe, 32'h407216df, 32'hc2b422a0, 32'h40079240, 32'h428a4216, 32'h4287cfb1};
test_output[17672:17679] = '{32'h420d562e, 32'h0, 32'h421836fe, 32'h407216df, 32'h0, 32'h40079240, 32'h428a4216, 32'h4287cfb1};
test_input[17680:17687] = '{32'h42a25a0a, 32'hc284736a, 32'h425390e7, 32'h42189d09, 32'h423ba2c7, 32'h42560795, 32'h42916794, 32'hc2bf5e63};
test_output[17680:17687] = '{32'h42a25a0a, 32'h0, 32'h425390e7, 32'h42189d09, 32'h423ba2c7, 32'h42560795, 32'h42916794, 32'h0};
test_input[17688:17695] = '{32'h41ee897d, 32'hc2b76e80, 32'h429a4989, 32'hc2aaead0, 32'h423e0dea, 32'hc1af9b13, 32'hc029b042, 32'h414bc3e8};
test_output[17688:17695] = '{32'h41ee897d, 32'h0, 32'h429a4989, 32'h0, 32'h423e0dea, 32'h0, 32'h0, 32'h414bc3e8};
test_input[17696:17703] = '{32'h4054baa1, 32'h4223a54d, 32'h417fef43, 32'hc2bc3f59, 32'h42aeddc4, 32'h41639200, 32'h42687e0c, 32'h42551b56};
test_output[17696:17703] = '{32'h4054baa1, 32'h4223a54d, 32'h417fef43, 32'h0, 32'h42aeddc4, 32'h41639200, 32'h42687e0c, 32'h42551b56};
test_input[17704:17711] = '{32'hc23b0e77, 32'h41810411, 32'h4210f434, 32'h40637313, 32'hc2892fe3, 32'hc18ce58c, 32'h41be33bf, 32'hc28eb775};
test_output[17704:17711] = '{32'h0, 32'h41810411, 32'h4210f434, 32'h40637313, 32'h0, 32'h0, 32'h41be33bf, 32'h0};
test_input[17712:17719] = '{32'h429850a6, 32'h40752481, 32'h4299e49f, 32'h42441c90, 32'h4149b8b2, 32'h41ea3bd0, 32'hc2adc915, 32'hc298cfb3};
test_output[17712:17719] = '{32'h429850a6, 32'h40752481, 32'h4299e49f, 32'h42441c90, 32'h4149b8b2, 32'h41ea3bd0, 32'h0, 32'h0};
test_input[17720:17727] = '{32'h4261293d, 32'h42afeb5a, 32'hc2a8b0fa, 32'hc2804bcd, 32'hc285a116, 32'hc16dbb24, 32'h4291a5be, 32'hc08f08a6};
test_output[17720:17727] = '{32'h4261293d, 32'h42afeb5a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4291a5be, 32'h0};
test_input[17728:17735] = '{32'h427ad5b2, 32'hc2c3793d, 32'hc2a4de65, 32'hc2705398, 32'hc1f76554, 32'hc11175b1, 32'h420ea823, 32'hc211029d};
test_output[17728:17735] = '{32'h427ad5b2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420ea823, 32'h0};
test_input[17736:17743] = '{32'h41c7277e, 32'h40607b78, 32'h429a4039, 32'hc2098631, 32'hc2730cd6, 32'hc2a36715, 32'hc206d177, 32'hc1aadf6b};
test_output[17736:17743] = '{32'h41c7277e, 32'h40607b78, 32'h429a4039, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[17744:17751] = '{32'h4265357c, 32'hc14c30d7, 32'h4274c7ed, 32'h413fa35a, 32'hc2b971d0, 32'h42a1e5a2, 32'hc1700202, 32'h428036e4};
test_output[17744:17751] = '{32'h4265357c, 32'h0, 32'h4274c7ed, 32'h413fa35a, 32'h0, 32'h42a1e5a2, 32'h0, 32'h428036e4};
test_input[17752:17759] = '{32'h42286df6, 32'h424fd562, 32'hc1b23ca2, 32'hc29fcabb, 32'hc239d570, 32'hc29c1c77, 32'hc28c67b0, 32'h4246877e};
test_output[17752:17759] = '{32'h42286df6, 32'h424fd562, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4246877e};
test_input[17760:17767] = '{32'hc0901d75, 32'hc2a7e024, 32'h4132bca8, 32'h40850291, 32'h42af0931, 32'h42547e11, 32'h42a52866, 32'h421c3c33};
test_output[17760:17767] = '{32'h0, 32'h0, 32'h4132bca8, 32'h40850291, 32'h42af0931, 32'h42547e11, 32'h42a52866, 32'h421c3c33};
test_input[17768:17775] = '{32'h41e6f9ed, 32'h420ab649, 32'hc2a1043a, 32'hc28c7307, 32'h4297b094, 32'h429cb6f2, 32'h4279bf08, 32'hc2110cfa};
test_output[17768:17775] = '{32'h41e6f9ed, 32'h420ab649, 32'h0, 32'h0, 32'h4297b094, 32'h429cb6f2, 32'h4279bf08, 32'h0};
test_input[17776:17783] = '{32'h42bed695, 32'hc2848618, 32'hc0bedd30, 32'hc1c5ca0e, 32'hc24530e8, 32'hc1acf121, 32'h429b20aa, 32'hc14c262c};
test_output[17776:17783] = '{32'h42bed695, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429b20aa, 32'h0};
test_input[17784:17791] = '{32'hc1d9a5d6, 32'h4286081d, 32'hc2a4178c, 32'h424e33e2, 32'h41f23db7, 32'h42c5879b, 32'h41c8f267, 32'h4290b846};
test_output[17784:17791] = '{32'h0, 32'h4286081d, 32'h0, 32'h424e33e2, 32'h41f23db7, 32'h42c5879b, 32'h41c8f267, 32'h4290b846};
test_input[17792:17799] = '{32'hc283c237, 32'hc2ad1103, 32'h423eaf8d, 32'hc115cc42, 32'hc249b0d7, 32'hc2743025, 32'h414ebe91, 32'h42876915};
test_output[17792:17799] = '{32'h0, 32'h0, 32'h423eaf8d, 32'h0, 32'h0, 32'h0, 32'h414ebe91, 32'h42876915};
test_input[17800:17807] = '{32'h41c6e19a, 32'hc1fe5b50, 32'h41f00b91, 32'h421fe75b, 32'hc24e202d, 32'hc2871d0d, 32'h42b8e092, 32'h42b959c1};
test_output[17800:17807] = '{32'h41c6e19a, 32'h0, 32'h41f00b91, 32'h421fe75b, 32'h0, 32'h0, 32'h42b8e092, 32'h42b959c1};
test_input[17808:17815] = '{32'hc1ea6641, 32'hc24ec1a0, 32'hc24b58a8, 32'hc286397c, 32'hbf9cf4dd, 32'hc24972ec, 32'hc230ab95, 32'hc1606568};
test_output[17808:17815] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[17816:17823] = '{32'hc294d6e0, 32'h410b5dac, 32'hc263e22f, 32'h41b6ab6f, 32'hc0d102d0, 32'h423694bf, 32'hc27d9716, 32'hc2c70244};
test_output[17816:17823] = '{32'h0, 32'h410b5dac, 32'h0, 32'h41b6ab6f, 32'h0, 32'h423694bf, 32'h0, 32'h0};
test_input[17824:17831] = '{32'hc2804b66, 32'h42810962, 32'h42ad23e0, 32'h412a457d, 32'h3e8ce89d, 32'h40174ba8, 32'h41b119f9, 32'hc2ac17fe};
test_output[17824:17831] = '{32'h0, 32'h42810962, 32'h42ad23e0, 32'h412a457d, 32'h3e8ce89d, 32'h40174ba8, 32'h41b119f9, 32'h0};
test_input[17832:17839] = '{32'h42311be1, 32'hc1b840c1, 32'hc266aa42, 32'hc1273db5, 32'h428138eb, 32'h403be4db, 32'h42bf5567, 32'h4259010b};
test_output[17832:17839] = '{32'h42311be1, 32'h0, 32'h0, 32'h0, 32'h428138eb, 32'h403be4db, 32'h42bf5567, 32'h4259010b};
test_input[17840:17847] = '{32'hc1a2dcdc, 32'hc2a8223c, 32'hc1cf3f36, 32'h421a7553, 32'h424d9bfe, 32'hc1973a3e, 32'h41d926fe, 32'h4286ebcd};
test_output[17840:17847] = '{32'h0, 32'h0, 32'h0, 32'h421a7553, 32'h424d9bfe, 32'h0, 32'h41d926fe, 32'h4286ebcd};
test_input[17848:17855] = '{32'h404e418a, 32'hc22c0c16, 32'hc28d84f1, 32'h428805f2, 32'h42a67607, 32'h40982909, 32'h42962c00, 32'h405d2bb9};
test_output[17848:17855] = '{32'h404e418a, 32'h0, 32'h0, 32'h428805f2, 32'h42a67607, 32'h40982909, 32'h42962c00, 32'h405d2bb9};
test_input[17856:17863] = '{32'h42b714ef, 32'hc23d69f9, 32'hc251d243, 32'h429038a8, 32'h42b6cc13, 32'h41fccacf, 32'hc251b1e5, 32'h4237599e};
test_output[17856:17863] = '{32'h42b714ef, 32'h0, 32'h0, 32'h429038a8, 32'h42b6cc13, 32'h41fccacf, 32'h0, 32'h4237599e};
test_input[17864:17871] = '{32'hc21af0af, 32'hc2641109, 32'h427359d1, 32'h4127e144, 32'hc253ce96, 32'h41b2d487, 32'hc284f3e8, 32'hc2c4e7b6};
test_output[17864:17871] = '{32'h0, 32'h0, 32'h427359d1, 32'h4127e144, 32'h0, 32'h41b2d487, 32'h0, 32'h0};
test_input[17872:17879] = '{32'h42a79482, 32'hc2c60120, 32'h42961ed0, 32'hc2998aff, 32'h4242f2e3, 32'hc2b900eb, 32'hc2add9a2, 32'hc29c4bdf};
test_output[17872:17879] = '{32'h42a79482, 32'h0, 32'h42961ed0, 32'h0, 32'h4242f2e3, 32'h0, 32'h0, 32'h0};
test_input[17880:17887] = '{32'hc2a34e60, 32'h42c4aa37, 32'h422bed94, 32'hc2a835d3, 32'h423fab3f, 32'hc044a299, 32'hc29dd6b9, 32'hc2955632};
test_output[17880:17887] = '{32'h0, 32'h42c4aa37, 32'h422bed94, 32'h0, 32'h423fab3f, 32'h0, 32'h0, 32'h0};
test_input[17888:17895] = '{32'hc2b526da, 32'h416bb9b6, 32'h422fd1e6, 32'hc0fa1421, 32'hc290f695, 32'hc29050fa, 32'h423627d1, 32'hc270379d};
test_output[17888:17895] = '{32'h0, 32'h416bb9b6, 32'h422fd1e6, 32'h0, 32'h0, 32'h0, 32'h423627d1, 32'h0};
test_input[17896:17903] = '{32'hc0687a46, 32'hc2b6aef0, 32'hc2b461bf, 32'hc1deed9a, 32'h42c70e2e, 32'hc206d268, 32'h4283d96e, 32'h42104389};
test_output[17896:17903] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42c70e2e, 32'h0, 32'h4283d96e, 32'h42104389};
test_input[17904:17911] = '{32'h423a82eb, 32'hc1aaa4bf, 32'hc03d37b7, 32'h42c26151, 32'h428fd8bd, 32'hc2100ed0, 32'h42b866a1, 32'h40fa995a};
test_output[17904:17911] = '{32'h423a82eb, 32'h0, 32'h0, 32'h42c26151, 32'h428fd8bd, 32'h0, 32'h42b866a1, 32'h40fa995a};
test_input[17912:17919] = '{32'h42a60e6f, 32'h41b714a5, 32'hc2a1936b, 32'h4266bb81, 32'hc2b70246, 32'h42c5eadf, 32'hc2498a82, 32'h425bc37a};
test_output[17912:17919] = '{32'h42a60e6f, 32'h41b714a5, 32'h0, 32'h4266bb81, 32'h0, 32'h42c5eadf, 32'h0, 32'h425bc37a};
test_input[17920:17927] = '{32'hc189581f, 32'hc1e2fb30, 32'h429e6500, 32'h40f2f82a, 32'hc2648a1d, 32'h42b36d8f, 32'h417ffd10, 32'h422120f6};
test_output[17920:17927] = '{32'h0, 32'h0, 32'h429e6500, 32'h40f2f82a, 32'h0, 32'h42b36d8f, 32'h417ffd10, 32'h422120f6};
test_input[17928:17935] = '{32'h4282dd40, 32'h4132c673, 32'h42a2baff, 32'h426d55f7, 32'h40545802, 32'hc265314c, 32'hc2ab8e3b, 32'h4214fe32};
test_output[17928:17935] = '{32'h4282dd40, 32'h4132c673, 32'h42a2baff, 32'h426d55f7, 32'h40545802, 32'h0, 32'h0, 32'h4214fe32};
test_input[17936:17943] = '{32'h424b5e80, 32'hc2943fd6, 32'h41090187, 32'h429a8dae, 32'h42a25b83, 32'h41ea129a, 32'hc15e1fa8, 32'h419758b1};
test_output[17936:17943] = '{32'h424b5e80, 32'h0, 32'h41090187, 32'h429a8dae, 32'h42a25b83, 32'h41ea129a, 32'h0, 32'h419758b1};
test_input[17944:17951] = '{32'hc256a547, 32'hc2963411, 32'hc0b5096d, 32'hc2ae1b96, 32'hc2962678, 32'hc295e1fe, 32'h423fb081, 32'hc21dab12};
test_output[17944:17951] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423fb081, 32'h0};
test_input[17952:17959] = '{32'h4292c4f3, 32'h42214f83, 32'hc280eb93, 32'h424e0eca, 32'h4219b83e, 32'hc2a82957, 32'hc2b1f14a, 32'hc2c01c61};
test_output[17952:17959] = '{32'h4292c4f3, 32'h42214f83, 32'h0, 32'h424e0eca, 32'h4219b83e, 32'h0, 32'h0, 32'h0};
test_input[17960:17967] = '{32'hc202ed1f, 32'hc2192ff1, 32'hc230e5e1, 32'h42ac4275, 32'h4211626b, 32'hc295865c, 32'hc2a28465, 32'hc24666b1};
test_output[17960:17967] = '{32'h0, 32'h0, 32'h0, 32'h42ac4275, 32'h4211626b, 32'h0, 32'h0, 32'h0};
test_input[17968:17975] = '{32'h421cf1e8, 32'h41a0222a, 32'h4148e8f8, 32'hc0fb2346, 32'hc2bf26f3, 32'h429b32f2, 32'hc2b2a5fb, 32'hc2a5fd6b};
test_output[17968:17975] = '{32'h421cf1e8, 32'h41a0222a, 32'h4148e8f8, 32'h0, 32'h0, 32'h429b32f2, 32'h0, 32'h0};
test_input[17976:17983] = '{32'hc208a486, 32'h424a0041, 32'hc2826bac, 32'hc2b9d5c7, 32'hc1f074a3, 32'h42bed6a5, 32'h40497c9a, 32'h409d008e};
test_output[17976:17983] = '{32'h0, 32'h424a0041, 32'h0, 32'h0, 32'h0, 32'h42bed6a5, 32'h40497c9a, 32'h409d008e};
test_input[17984:17991] = '{32'hc2500e34, 32'hc23f647e, 32'h4266e0cd, 32'hc1940048, 32'h42662ade, 32'hc10be788, 32'hc255b2bc, 32'h41dfd86e};
test_output[17984:17991] = '{32'h0, 32'h0, 32'h4266e0cd, 32'h0, 32'h42662ade, 32'h0, 32'h0, 32'h41dfd86e};
test_input[17992:17999] = '{32'hc29a3746, 32'hc29980fd, 32'hc1e39b9a, 32'hc0c4a04b, 32'hc13e3128, 32'hc139291b, 32'hc1ac5b84, 32'hc27e8ac1};
test_output[17992:17999] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18000:18007] = '{32'hc29399e5, 32'h4234414a, 32'hc29a7320, 32'h42c61f80, 32'hc250dd33, 32'h4282a3d8, 32'hc2b2eb7f, 32'hc1155028};
test_output[18000:18007] = '{32'h0, 32'h4234414a, 32'h0, 32'h42c61f80, 32'h0, 32'h4282a3d8, 32'h0, 32'h0};
test_input[18008:18015] = '{32'h414eff28, 32'h41ad9fa4, 32'h41921e9f, 32'hc280c43e, 32'hc1d67b45, 32'hc2c45157, 32'h429424ab, 32'h42b0bc02};
test_output[18008:18015] = '{32'h414eff28, 32'h41ad9fa4, 32'h41921e9f, 32'h0, 32'h0, 32'h0, 32'h429424ab, 32'h42b0bc02};
test_input[18016:18023] = '{32'hc1d578cf, 32'h4250b3b7, 32'h422e5681, 32'h429bcae8, 32'h42bcc928, 32'hc21833b3, 32'hc2538c7f, 32'h4105913a};
test_output[18016:18023] = '{32'h0, 32'h4250b3b7, 32'h422e5681, 32'h429bcae8, 32'h42bcc928, 32'h0, 32'h0, 32'h4105913a};
test_input[18024:18031] = '{32'hc19c9fdc, 32'h428e4e4d, 32'h4205d729, 32'h4260e8e8, 32'hc2a52e23, 32'hc1a60ce1, 32'h40d21cff, 32'hc232d605};
test_output[18024:18031] = '{32'h0, 32'h428e4e4d, 32'h4205d729, 32'h4260e8e8, 32'h0, 32'h0, 32'h40d21cff, 32'h0};
test_input[18032:18039] = '{32'hc2914a24, 32'hc225f2a3, 32'h425ccea6, 32'h419a58fe, 32'hc22217c1, 32'hc28c4336, 32'h41958214, 32'h424c881e};
test_output[18032:18039] = '{32'h0, 32'h0, 32'h425ccea6, 32'h419a58fe, 32'h0, 32'h0, 32'h41958214, 32'h424c881e};
test_input[18040:18047] = '{32'h42069181, 32'h41e5492e, 32'hc257cfaa, 32'h41dff0ad, 32'hc1b4ff91, 32'h3f8268a9, 32'hbfc0b81b, 32'h418955e5};
test_output[18040:18047] = '{32'h42069181, 32'h41e5492e, 32'h0, 32'h41dff0ad, 32'h0, 32'h3f8268a9, 32'h0, 32'h418955e5};
test_input[18048:18055] = '{32'hc1c5a84a, 32'hc2691b2a, 32'h42b62c09, 32'h4262c577, 32'hc255f962, 32'hc2173cbf, 32'h42a56062, 32'h42681f8d};
test_output[18048:18055] = '{32'h0, 32'h0, 32'h42b62c09, 32'h4262c577, 32'h0, 32'h0, 32'h42a56062, 32'h42681f8d};
test_input[18056:18063] = '{32'hc21863eb, 32'h4291e169, 32'h41a6ff24, 32'h4299eaad, 32'h424b3c5d, 32'h41a6522a, 32'h427a0982, 32'hc1d01bef};
test_output[18056:18063] = '{32'h0, 32'h4291e169, 32'h41a6ff24, 32'h4299eaad, 32'h424b3c5d, 32'h41a6522a, 32'h427a0982, 32'h0};
test_input[18064:18071] = '{32'hc2a09a76, 32'hc2833327, 32'hc28a1bf9, 32'hc262bc90, 32'h425f85a6, 32'h419ceaf8, 32'hc29ed626, 32'h428c5c91};
test_output[18064:18071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h425f85a6, 32'h419ceaf8, 32'h0, 32'h428c5c91};
test_input[18072:18079] = '{32'h425caaef, 32'h4238fced, 32'hc28edce2, 32'h428a1596, 32'hc29f233a, 32'hc287f721, 32'h428cc5ba, 32'hc26ea450};
test_output[18072:18079] = '{32'h425caaef, 32'h4238fced, 32'h0, 32'h428a1596, 32'h0, 32'h0, 32'h428cc5ba, 32'h0};
test_input[18080:18087] = '{32'hc2b3bd19, 32'hc2b546d6, 32'hc1fe1d15, 32'hc275c4a6, 32'h420d56c8, 32'hc199958d, 32'hc156f18f, 32'hc2952907};
test_output[18080:18087] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h420d56c8, 32'h0, 32'h0, 32'h0};
test_input[18088:18095] = '{32'h41a6dbc7, 32'h4255f2be, 32'hc0ec7566, 32'h41bd4957, 32'h429051aa, 32'h42b88f8f, 32'hc28dc9c4, 32'hc2c6feed};
test_output[18088:18095] = '{32'h41a6dbc7, 32'h4255f2be, 32'h0, 32'h41bd4957, 32'h429051aa, 32'h42b88f8f, 32'h0, 32'h0};
test_input[18096:18103] = '{32'h41d01724, 32'h41b2abed, 32'h4197f55b, 32'h421366e3, 32'h3ff3485c, 32'hc0871298, 32'hc221a6f7, 32'hc22ecf93};
test_output[18096:18103] = '{32'h41d01724, 32'h41b2abed, 32'h4197f55b, 32'h421366e3, 32'h3ff3485c, 32'h0, 32'h0, 32'h0};
test_input[18104:18111] = '{32'hc28f073a, 32'h41c0b231, 32'h416c470d, 32'h42803df0, 32'h429cb97d, 32'h42849ad4, 32'hc211e98a, 32'h4142fa7e};
test_output[18104:18111] = '{32'h0, 32'h41c0b231, 32'h416c470d, 32'h42803df0, 32'h429cb97d, 32'h42849ad4, 32'h0, 32'h4142fa7e};
test_input[18112:18119] = '{32'h41e79c25, 32'hc21efdfa, 32'h41721a6c, 32'hc21278a1, 32'h41f83954, 32'hc1384e8f, 32'h42ad3fa7, 32'hc265ce44};
test_output[18112:18119] = '{32'h41e79c25, 32'h0, 32'h41721a6c, 32'h0, 32'h41f83954, 32'h0, 32'h42ad3fa7, 32'h0};
test_input[18120:18127] = '{32'h41cd65f1, 32'hc270e234, 32'hc1ce0dc5, 32'h42051b4f, 32'h423d2fa8, 32'h42b36ceb, 32'h419a6776, 32'h420bc5d7};
test_output[18120:18127] = '{32'h41cd65f1, 32'h0, 32'h0, 32'h42051b4f, 32'h423d2fa8, 32'h42b36ceb, 32'h419a6776, 32'h420bc5d7};
test_input[18128:18135] = '{32'hc1e37f79, 32'hc2b4afcd, 32'hc2a579f9, 32'h42c4009d, 32'h41c47881, 32'h42983e33, 32'h4283fa47, 32'h42c76c68};
test_output[18128:18135] = '{32'h0, 32'h0, 32'h0, 32'h42c4009d, 32'h41c47881, 32'h42983e33, 32'h4283fa47, 32'h42c76c68};
test_input[18136:18143] = '{32'hc19e608c, 32'h4165d20a, 32'h42903fab, 32'h423eddb4, 32'h42736e31, 32'h420bce41, 32'h41da73de, 32'h42807dba};
test_output[18136:18143] = '{32'h0, 32'h4165d20a, 32'h42903fab, 32'h423eddb4, 32'h42736e31, 32'h420bce41, 32'h41da73de, 32'h42807dba};
test_input[18144:18151] = '{32'h428eced0, 32'hc20d7e6f, 32'hc219d7ff, 32'hc1d7bd7e, 32'hc2816753, 32'hc2c18b3c, 32'hc23b1d5a, 32'h425d9b96};
test_output[18144:18151] = '{32'h428eced0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425d9b96};
test_input[18152:18159] = '{32'hc248a0a1, 32'hc25a7b94, 32'hc2a257d2, 32'hc283842b, 32'hc2beaeab, 32'h41b5c28e, 32'hc22228a7, 32'hc2800f3f};
test_output[18152:18159] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b5c28e, 32'h0, 32'h0};
test_input[18160:18167] = '{32'h4291d921, 32'hc218fec2, 32'h416308ef, 32'hc22a4860, 32'h41b55983, 32'h424265ad, 32'h403e999c, 32'hc2bb1216};
test_output[18160:18167] = '{32'h4291d921, 32'h0, 32'h416308ef, 32'h0, 32'h41b55983, 32'h424265ad, 32'h403e999c, 32'h0};
test_input[18168:18175] = '{32'h4188325c, 32'hc2b83f08, 32'hc2b9b707, 32'hc21ffd4e, 32'hc2a0841e, 32'hc1817086, 32'h42a5a20a, 32'hc2ac67ab};
test_output[18168:18175] = '{32'h4188325c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a5a20a, 32'h0};
test_input[18176:18183] = '{32'h427b0ba4, 32'hc2b3c364, 32'h42999716, 32'hc1835f3d, 32'h4090f65e, 32'hc29d8f0e, 32'hc2c54cd4, 32'h42c0ef16};
test_output[18176:18183] = '{32'h427b0ba4, 32'h0, 32'h42999716, 32'h0, 32'h4090f65e, 32'h0, 32'h0, 32'h42c0ef16};
test_input[18184:18191] = '{32'hc29c9c20, 32'h42071b4e, 32'h417d4f9d, 32'hc1d06173, 32'hc1bb13f2, 32'hc2937ad4, 32'h426eb0bd, 32'h41870635};
test_output[18184:18191] = '{32'h0, 32'h42071b4e, 32'h417d4f9d, 32'h0, 32'h0, 32'h0, 32'h426eb0bd, 32'h41870635};
test_input[18192:18199] = '{32'hc28ae883, 32'hc158f107, 32'h41b2687a, 32'h41b1d4c8, 32'h42ad60ea, 32'hc27e6300, 32'h41bac080, 32'hc21ca0f3};
test_output[18192:18199] = '{32'h0, 32'h0, 32'h41b2687a, 32'h41b1d4c8, 32'h42ad60ea, 32'h0, 32'h41bac080, 32'h0};
test_input[18200:18207] = '{32'h429aa2a8, 32'h42af57c5, 32'hc27f41b3, 32'h42428a4e, 32'hc2c7776b, 32'h42058d58, 32'hc10b104b, 32'hc1ac9743};
test_output[18200:18207] = '{32'h429aa2a8, 32'h42af57c5, 32'h0, 32'h42428a4e, 32'h0, 32'h42058d58, 32'h0, 32'h0};
test_input[18208:18215] = '{32'hc0002e0a, 32'hbff2f091, 32'hc27f8aca, 32'h41cafb83, 32'hc20738be, 32'hc285ebe1, 32'hc27e1f38, 32'h4239aad3};
test_output[18208:18215] = '{32'h0, 32'h0, 32'h0, 32'h41cafb83, 32'h0, 32'h0, 32'h0, 32'h4239aad3};
test_input[18216:18223] = '{32'h4293c15e, 32'hc2957939, 32'h409c39ed, 32'h42c06ff9, 32'h42725ab8, 32'h409b9081, 32'hc2c08ce7, 32'hc1adb067};
test_output[18216:18223] = '{32'h4293c15e, 32'h0, 32'h409c39ed, 32'h42c06ff9, 32'h42725ab8, 32'h409b9081, 32'h0, 32'h0};
test_input[18224:18231] = '{32'h423215d1, 32'h426ab268, 32'hc23082ee, 32'hc27b7fbf, 32'h429d5f2d, 32'h41527dbc, 32'h426767fa, 32'h4185ead4};
test_output[18224:18231] = '{32'h423215d1, 32'h426ab268, 32'h0, 32'h0, 32'h429d5f2d, 32'h41527dbc, 32'h426767fa, 32'h4185ead4};
test_input[18232:18239] = '{32'hc1d61266, 32'hc281d96e, 32'hc2b6000c, 32'h42466f2d, 32'hc27ee070, 32'hc2363c01, 32'h42b33f6f, 32'h42bdde48};
test_output[18232:18239] = '{32'h0, 32'h0, 32'h0, 32'h42466f2d, 32'h0, 32'h0, 32'h42b33f6f, 32'h42bdde48};
test_input[18240:18247] = '{32'hc154f2a9, 32'h4241a136, 32'hc27bde09, 32'h42a4d049, 32'h42747648, 32'h42c41c0e, 32'h428a9802, 32'h42a42304};
test_output[18240:18247] = '{32'h0, 32'h4241a136, 32'h0, 32'h42a4d049, 32'h42747648, 32'h42c41c0e, 32'h428a9802, 32'h42a42304};
test_input[18248:18255] = '{32'hc25fd151, 32'h42b45290, 32'h4242ccf3, 32'h411e2d96, 32'hc2b66e77, 32'hc10794b4, 32'h4267a9f0, 32'h418d43dd};
test_output[18248:18255] = '{32'h0, 32'h42b45290, 32'h4242ccf3, 32'h411e2d96, 32'h0, 32'h0, 32'h4267a9f0, 32'h418d43dd};
test_input[18256:18263] = '{32'hc207979b, 32'h4207c8e5, 32'h423275c7, 32'h42728142, 32'hc0c7a64d, 32'hc1a06262, 32'h4225909f, 32'hc28976b8};
test_output[18256:18263] = '{32'h0, 32'h4207c8e5, 32'h423275c7, 32'h42728142, 32'h0, 32'h0, 32'h4225909f, 32'h0};
test_input[18264:18271] = '{32'hbe795d50, 32'hc2960613, 32'hc29b1a5f, 32'hc13cf023, 32'h426b8f30, 32'hc29f56da, 32'hc23c813b, 32'hc221bb98};
test_output[18264:18271] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h426b8f30, 32'h0, 32'h0, 32'h0};
test_input[18272:18279] = '{32'hc2577d66, 32'h428d5610, 32'hc238b11a, 32'hc2b0d321, 32'h426fa74d, 32'h428e6f50, 32'hc2c5296d, 32'h413bd93e};
test_output[18272:18279] = '{32'h0, 32'h428d5610, 32'h0, 32'h0, 32'h426fa74d, 32'h428e6f50, 32'h0, 32'h413bd93e};
test_input[18280:18287] = '{32'h40356d06, 32'hc237c0c6, 32'h424240aa, 32'h429482f1, 32'h4278113c, 32'h42a7dedb, 32'hc21c4554, 32'h428b3191};
test_output[18280:18287] = '{32'h40356d06, 32'h0, 32'h424240aa, 32'h429482f1, 32'h4278113c, 32'h42a7dedb, 32'h0, 32'h428b3191};
test_input[18288:18295] = '{32'h4036eaaa, 32'h425ca8e7, 32'h4292f598, 32'h41748f00, 32'hc1e66382, 32'h4231af4f, 32'h40698822, 32'hc2380ffd};
test_output[18288:18295] = '{32'h4036eaaa, 32'h425ca8e7, 32'h4292f598, 32'h41748f00, 32'h0, 32'h4231af4f, 32'h40698822, 32'h0};
test_input[18296:18303] = '{32'h41081fe3, 32'h423f7efd, 32'hc2bdf439, 32'hc213aca7, 32'h41b91190, 32'hc2b0e0d5, 32'hc22bfffc, 32'hc28e1d76};
test_output[18296:18303] = '{32'h41081fe3, 32'h423f7efd, 32'h0, 32'h0, 32'h41b91190, 32'h0, 32'h0, 32'h0};
test_input[18304:18311] = '{32'h41b18f14, 32'h40847808, 32'h4275bc09, 32'h428d68af, 32'hc1d0a575, 32'h429c5a8b, 32'hc1e630af, 32'hc2909929};
test_output[18304:18311] = '{32'h41b18f14, 32'h40847808, 32'h4275bc09, 32'h428d68af, 32'h0, 32'h429c5a8b, 32'h0, 32'h0};
test_input[18312:18319] = '{32'h428f1585, 32'hc1947a27, 32'hc20ce9b3, 32'hc2aa35d6, 32'hc21fef85, 32'hc2ba773e, 32'h428f5f60, 32'h42befafe};
test_output[18312:18319] = '{32'h428f1585, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428f5f60, 32'h42befafe};
test_input[18320:18327] = '{32'h428d66ec, 32'hc2679e58, 32'hc1c4103b, 32'h42a41c67, 32'hc1c01a75, 32'hc1ab02dd, 32'hc0d81285, 32'hc2a62ea4};
test_output[18320:18327] = '{32'h428d66ec, 32'h0, 32'h0, 32'h42a41c67, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18328:18335] = '{32'h42c37ac7, 32'hc1b46df4, 32'h41492111, 32'h42790d06, 32'hc223f86c, 32'h42a55775, 32'h424b2b87, 32'hc2af7e95};
test_output[18328:18335] = '{32'h42c37ac7, 32'h0, 32'h41492111, 32'h42790d06, 32'h0, 32'h42a55775, 32'h424b2b87, 32'h0};
test_input[18336:18343] = '{32'hc0cb8386, 32'hc077c297, 32'hc28c0d1f, 32'hc269ecd5, 32'hc29189ca, 32'hc2ba4b4e, 32'h42ba6a24, 32'h42aff0c5};
test_output[18336:18343] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ba6a24, 32'h42aff0c5};
test_input[18344:18351] = '{32'h4211c384, 32'h4174a9fb, 32'h428b0dcc, 32'hc1ee6c49, 32'h421aaa47, 32'hc0ef0ccd, 32'hc20bedf2, 32'hbfed19a2};
test_output[18344:18351] = '{32'h4211c384, 32'h4174a9fb, 32'h428b0dcc, 32'h0, 32'h421aaa47, 32'h0, 32'h0, 32'h0};
test_input[18352:18359] = '{32'h429161e5, 32'hc25a0632, 32'hc25794f5, 32'hc0369be3, 32'h42492b62, 32'h41e5dd17, 32'hc2969c11, 32'hc24f59d2};
test_output[18352:18359] = '{32'h429161e5, 32'h0, 32'h0, 32'h0, 32'h42492b62, 32'h41e5dd17, 32'h0, 32'h0};
test_input[18360:18367] = '{32'hc1121a3f, 32'h42870aae, 32'h42756ebb, 32'h42b5ce82, 32'h423b54e5, 32'h42a22327, 32'hc1f6db39, 32'h42addd4a};
test_output[18360:18367] = '{32'h0, 32'h42870aae, 32'h42756ebb, 32'h42b5ce82, 32'h423b54e5, 32'h42a22327, 32'h0, 32'h42addd4a};
test_input[18368:18375] = '{32'hc2c677b7, 32'h427ac455, 32'h40fe7f68, 32'hc2909564, 32'h4288fcbb, 32'h417f2d39, 32'hc2b00367, 32'hc12804aa};
test_output[18368:18375] = '{32'h0, 32'h427ac455, 32'h40fe7f68, 32'h0, 32'h4288fcbb, 32'h417f2d39, 32'h0, 32'h0};
test_input[18376:18383] = '{32'hc2236c49, 32'h41124276, 32'h4287fba1, 32'h41183245, 32'h4242d6bb, 32'h42a53fa0, 32'hc20410df, 32'h41b2b11a};
test_output[18376:18383] = '{32'h0, 32'h41124276, 32'h4287fba1, 32'h41183245, 32'h4242d6bb, 32'h42a53fa0, 32'h0, 32'h41b2b11a};
test_input[18384:18391] = '{32'h422e4da9, 32'h42ad62a4, 32'hc2a4ac63, 32'h42a54040, 32'h42a765fa, 32'hc2890eef, 32'hc226061e, 32'hc18db6f2};
test_output[18384:18391] = '{32'h422e4da9, 32'h42ad62a4, 32'h0, 32'h42a54040, 32'h42a765fa, 32'h0, 32'h0, 32'h0};
test_input[18392:18399] = '{32'h42a32b8f, 32'hc2bbe29a, 32'hc2070f31, 32'hc2c47e57, 32'hc17011e6, 32'hc250df52, 32'h415d7c6f, 32'h40e6ac42};
test_output[18392:18399] = '{32'h42a32b8f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h415d7c6f, 32'h40e6ac42};
test_input[18400:18407] = '{32'hc23892f9, 32'hc2369f4b, 32'h425fb966, 32'h425134ef, 32'hbfe87dde, 32'hc26c0af7, 32'h42add44e, 32'h42576c15};
test_output[18400:18407] = '{32'h0, 32'h0, 32'h425fb966, 32'h425134ef, 32'h0, 32'h0, 32'h42add44e, 32'h42576c15};
test_input[18408:18415] = '{32'hbfaeb97c, 32'hc2220386, 32'hc069828a, 32'h4208edd8, 32'h4168b97b, 32'hbf554712, 32'h42048bc0, 32'h427d3227};
test_output[18408:18415] = '{32'h0, 32'h0, 32'h0, 32'h4208edd8, 32'h4168b97b, 32'h0, 32'h42048bc0, 32'h427d3227};
test_input[18416:18423] = '{32'hc28da154, 32'hc2543a22, 32'hc29d0eb4, 32'hc2535acc, 32'h4280cbd3, 32'hc20283bd, 32'hc28ef5d0, 32'hc293f6ec};
test_output[18416:18423] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4280cbd3, 32'h0, 32'h0, 32'h0};
test_input[18424:18431] = '{32'hc22d25a4, 32'h429e3acd, 32'hc0d47a05, 32'h3de05523, 32'h42167104, 32'hc2190029, 32'hc29605a4, 32'h42bb93dc};
test_output[18424:18431] = '{32'h0, 32'h429e3acd, 32'h0, 32'h3de05523, 32'h42167104, 32'h0, 32'h0, 32'h42bb93dc};
test_input[18432:18439] = '{32'h42a6d024, 32'h42c2df14, 32'hc2c25c8a, 32'h425894a9, 32'hc1e5a315, 32'h3fb1eeba, 32'h41ed929f, 32'h423bb84c};
test_output[18432:18439] = '{32'h42a6d024, 32'h42c2df14, 32'h0, 32'h425894a9, 32'h0, 32'h3fb1eeba, 32'h41ed929f, 32'h423bb84c};
test_input[18440:18447] = '{32'hc2704c58, 32'h426c2860, 32'hc2283cd5, 32'h41ad8fef, 32'hc1fab4e9, 32'hc2a2e0b0, 32'h420c6dbe, 32'h420c8146};
test_output[18440:18447] = '{32'h0, 32'h426c2860, 32'h0, 32'h41ad8fef, 32'h0, 32'h0, 32'h420c6dbe, 32'h420c8146};
test_input[18448:18455] = '{32'h426aed60, 32'hc2c2d219, 32'hc22b522c, 32'hc2bacd70, 32'hc1239ef0, 32'hc10efb5e, 32'hc2c3337d, 32'h425299b5};
test_output[18448:18455] = '{32'h426aed60, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425299b5};
test_input[18456:18463] = '{32'hc198eaab, 32'hc28afc69, 32'hc21f5371, 32'hc2892b54, 32'hc240a2e8, 32'hc2bfb8ce, 32'hc26b7a42, 32'hc2c33556};
test_output[18456:18463] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18464:18471] = '{32'hc289537a, 32'hc219ceb6, 32'h42aa137f, 32'h429d7004, 32'h42bce573, 32'hc1e930f8, 32'h4249bce3, 32'h423c18a3};
test_output[18464:18471] = '{32'h0, 32'h0, 32'h42aa137f, 32'h429d7004, 32'h42bce573, 32'h0, 32'h4249bce3, 32'h423c18a3};
test_input[18472:18479] = '{32'hc2968006, 32'h4100cae0, 32'h42b11b45, 32'h42b9a30e, 32'hc24f82e1, 32'h42b15039, 32'hc233cbe8, 32'h402c882e};
test_output[18472:18479] = '{32'h0, 32'h4100cae0, 32'h42b11b45, 32'h42b9a30e, 32'h0, 32'h42b15039, 32'h0, 32'h402c882e};
test_input[18480:18487] = '{32'h415cc9c2, 32'h42abd1c3, 32'h425e43de, 32'hc2237681, 32'hc2c2fbf2, 32'hc1be23b3, 32'h4299e7c4, 32'h4130f3fa};
test_output[18480:18487] = '{32'h415cc9c2, 32'h42abd1c3, 32'h425e43de, 32'h0, 32'h0, 32'h0, 32'h4299e7c4, 32'h4130f3fa};
test_input[18488:18495] = '{32'hc2a122b9, 32'hc2bc53ce, 32'h40dde779, 32'hc2835ccc, 32'hc2b1ca34, 32'hc2a98d91, 32'h41dca231, 32'hc25a87e4};
test_output[18488:18495] = '{32'h0, 32'h0, 32'h40dde779, 32'h0, 32'h0, 32'h0, 32'h41dca231, 32'h0};
test_input[18496:18503] = '{32'hc06afb20, 32'hc2b8b55e, 32'h4299c633, 32'h41e108e0, 32'hc29c2002, 32'h42bd3638, 32'hc2167aa0, 32'hc1c0b053};
test_output[18496:18503] = '{32'h0, 32'h0, 32'h4299c633, 32'h41e108e0, 32'h0, 32'h42bd3638, 32'h0, 32'h0};
test_input[18504:18511] = '{32'hc2bc78aa, 32'h42ac2c7c, 32'h424e8794, 32'hc2ace450, 32'h42a9a3c9, 32'h426e6e7f, 32'hc24f2be8, 32'h424bcac7};
test_output[18504:18511] = '{32'h0, 32'h42ac2c7c, 32'h424e8794, 32'h0, 32'h42a9a3c9, 32'h426e6e7f, 32'h0, 32'h424bcac7};
test_input[18512:18519] = '{32'hc2b8bcb6, 32'hc198ac5f, 32'hc2b333a9, 32'h4085410f, 32'hc246b61a, 32'h4204a059, 32'h403e5844, 32'h3f684c53};
test_output[18512:18519] = '{32'h0, 32'h0, 32'h0, 32'h4085410f, 32'h0, 32'h4204a059, 32'h403e5844, 32'h3f684c53};
test_input[18520:18527] = '{32'hc2bdce14, 32'h4294905d, 32'hc20d98cf, 32'hc254867b, 32'hc1a8164e, 32'hc22b2bcf, 32'h42bab927, 32'h416a2979};
test_output[18520:18527] = '{32'h0, 32'h4294905d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bab927, 32'h416a2979};
test_input[18528:18535] = '{32'h4253778e, 32'hc0f76273, 32'h42c0d003, 32'hc2bddbc9, 32'hc2c04dc1, 32'hc1948012, 32'h428492fb, 32'h4085d1d0};
test_output[18528:18535] = '{32'h4253778e, 32'h0, 32'h42c0d003, 32'h0, 32'h0, 32'h0, 32'h428492fb, 32'h4085d1d0};
test_input[18536:18543] = '{32'h420d6c13, 32'h42014ff4, 32'hc2c44d4b, 32'h422283f6, 32'hc228b032, 32'hc19e30cb, 32'h42a76b61, 32'hc10ee7a9};
test_output[18536:18543] = '{32'h420d6c13, 32'h42014ff4, 32'h0, 32'h422283f6, 32'h0, 32'h0, 32'h42a76b61, 32'h0};
test_input[18544:18551] = '{32'h42a61247, 32'h429f710e, 32'hc272de9f, 32'h42382a67, 32'hc249730a, 32'h4295658f, 32'hc05cf2c9, 32'hc24001c5};
test_output[18544:18551] = '{32'h42a61247, 32'h429f710e, 32'h0, 32'h42382a67, 32'h0, 32'h4295658f, 32'h0, 32'h0};
test_input[18552:18559] = '{32'hc28d29f0, 32'hc0231e7d, 32'h420b49b5, 32'hc1c59aeb, 32'h42b62c02, 32'h410ce6b8, 32'hc181aa44, 32'hc268d708};
test_output[18552:18559] = '{32'h0, 32'h0, 32'h420b49b5, 32'h0, 32'h42b62c02, 32'h410ce6b8, 32'h0, 32'h0};
test_input[18560:18567] = '{32'hc28c793f, 32'h42929b6f, 32'h41fde254, 32'h41b20113, 32'hc1ce55b5, 32'hc26fcd70, 32'h4299b88b, 32'hc2453db5};
test_output[18560:18567] = '{32'h0, 32'h42929b6f, 32'h41fde254, 32'h41b20113, 32'h0, 32'h0, 32'h4299b88b, 32'h0};
test_input[18568:18575] = '{32'hc22974a2, 32'hc2c350b3, 32'h41c2afc4, 32'h427cf032, 32'h41075946, 32'h4226b708, 32'h427a0b99, 32'h42934986};
test_output[18568:18575] = '{32'h0, 32'h0, 32'h41c2afc4, 32'h427cf032, 32'h41075946, 32'h4226b708, 32'h427a0b99, 32'h42934986};
test_input[18576:18583] = '{32'hc267a199, 32'hc2808499, 32'h4236eefb, 32'hc296ce05, 32'h42523006, 32'hc2354fff, 32'hc2b5e0fc, 32'hc26a19ab};
test_output[18576:18583] = '{32'h0, 32'h0, 32'h4236eefb, 32'h0, 32'h42523006, 32'h0, 32'h0, 32'h0};
test_input[18584:18591] = '{32'h4260c3ee, 32'h4291ac5f, 32'hc2a36aff, 32'h42b5c09c, 32'h425a9f87, 32'h426e5d22, 32'hc24bc9b7, 32'h4201b5c3};
test_output[18584:18591] = '{32'h4260c3ee, 32'h4291ac5f, 32'h0, 32'h42b5c09c, 32'h425a9f87, 32'h426e5d22, 32'h0, 32'h4201b5c3};
test_input[18592:18599] = '{32'hc1bcf77d, 32'hc23acd4a, 32'h4221c3a4, 32'h42854e40, 32'h3fc10cc5, 32'hc1be3126, 32'h42a150fc, 32'h42a0406e};
test_output[18592:18599] = '{32'h0, 32'h0, 32'h4221c3a4, 32'h42854e40, 32'h3fc10cc5, 32'h0, 32'h42a150fc, 32'h42a0406e};
test_input[18600:18607] = '{32'hc1b2c40f, 32'hc22e7efb, 32'hc1dc76de, 32'h41d8ba67, 32'hc2c0d23a, 32'h4297d489, 32'hc219cfde, 32'h422ed256};
test_output[18600:18607] = '{32'h0, 32'h0, 32'h0, 32'h41d8ba67, 32'h0, 32'h4297d489, 32'h0, 32'h422ed256};
test_input[18608:18615] = '{32'h4196247b, 32'hc0547d94, 32'h42935a4a, 32'h425482ef, 32'hc0f79201, 32'hc12d0780, 32'h418ce1b8, 32'h421d3d6c};
test_output[18608:18615] = '{32'h4196247b, 32'h0, 32'h42935a4a, 32'h425482ef, 32'h0, 32'h0, 32'h418ce1b8, 32'h421d3d6c};
test_input[18616:18623] = '{32'hc112e013, 32'h418fe1fe, 32'hc1b19e79, 32'h429abf23, 32'hc247a820, 32'h3fddd1e5, 32'h428d90a2, 32'hc2929560};
test_output[18616:18623] = '{32'h0, 32'h418fe1fe, 32'h0, 32'h429abf23, 32'h0, 32'h3fddd1e5, 32'h428d90a2, 32'h0};
test_input[18624:18631] = '{32'hbc0e03d5, 32'hc2623fef, 32'hc292582c, 32'hc29d366c, 32'hc2c68bb1, 32'hc2356272, 32'h408d7311, 32'hc28e3bee};
test_output[18624:18631] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h408d7311, 32'h0};
test_input[18632:18639] = '{32'hc033a6fa, 32'hc20fd5dc, 32'h4291e75e, 32'hc1d5ea2d, 32'h41c1123e, 32'hc2bf8b68, 32'h4287ed35, 32'hc2bbf268};
test_output[18632:18639] = '{32'h0, 32'h0, 32'h4291e75e, 32'h0, 32'h41c1123e, 32'h0, 32'h4287ed35, 32'h0};
test_input[18640:18647] = '{32'hc2849003, 32'h41a3f8a9, 32'h424031d3, 32'h41f1a8c8, 32'h42a55758, 32'hc294abbe, 32'h42b864f6, 32'hc28d46f4};
test_output[18640:18647] = '{32'h0, 32'h41a3f8a9, 32'h424031d3, 32'h41f1a8c8, 32'h42a55758, 32'h0, 32'h42b864f6, 32'h0};
test_input[18648:18655] = '{32'hc279c9a1, 32'hc2990a27, 32'hc23e0ce0, 32'h41f99ab3, 32'h42a8a5b8, 32'hc28af740, 32'h42006386, 32'h425135ff};
test_output[18648:18655] = '{32'h0, 32'h0, 32'h0, 32'h41f99ab3, 32'h42a8a5b8, 32'h0, 32'h42006386, 32'h425135ff};
test_input[18656:18663] = '{32'hc232fe55, 32'hc22f98ca, 32'hc1683567, 32'hc2ad49ff, 32'h42c26403, 32'hc2002d56, 32'hc262e22a, 32'h41f01296};
test_output[18656:18663] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42c26403, 32'h0, 32'h0, 32'h41f01296};
test_input[18664:18671] = '{32'h42bbed44, 32'h41ab4565, 32'h4255e32a, 32'hc2817e9d, 32'hc1ecd24e, 32'h41b5f668, 32'hc29715cf, 32'hc2ac5406};
test_output[18664:18671] = '{32'h42bbed44, 32'h41ab4565, 32'h4255e32a, 32'h0, 32'h0, 32'h41b5f668, 32'h0, 32'h0};
test_input[18672:18679] = '{32'hc2c00e19, 32'hc2aa4cc9, 32'hc2acd3a0, 32'hc267a30b, 32'hc2a606cf, 32'hc2c43960, 32'hc1d4053a, 32'h42bcfd8d};
test_output[18672:18679] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bcfd8d};
test_input[18680:18687] = '{32'hc2c2107f, 32'h42810631, 32'h42868d1c, 32'hc1d617bb, 32'h42a2db33, 32'hc205b96f, 32'h423eebc3, 32'hc2c6a7c1};
test_output[18680:18687] = '{32'h0, 32'h42810631, 32'h42868d1c, 32'h0, 32'h42a2db33, 32'h0, 32'h423eebc3, 32'h0};
test_input[18688:18695] = '{32'hc2b1e3a8, 32'hc1f2b394, 32'h423d5418, 32'h42c40730, 32'h425b7c08, 32'h41839af4, 32'h420a81bf, 32'hc22126d2};
test_output[18688:18695] = '{32'h0, 32'h0, 32'h423d5418, 32'h42c40730, 32'h425b7c08, 32'h41839af4, 32'h420a81bf, 32'h0};
test_input[18696:18703] = '{32'hc2159e95, 32'h41dcfdae, 32'h41820456, 32'h4282950d, 32'hc297a69a, 32'h42404f0d, 32'hc1cb1b8e, 32'hc1bb798a};
test_output[18696:18703] = '{32'h0, 32'h41dcfdae, 32'h41820456, 32'h4282950d, 32'h0, 32'h42404f0d, 32'h0, 32'h0};
test_input[18704:18711] = '{32'h4124b772, 32'hc12bfc8c, 32'hc22482b7, 32'hc2311304, 32'h42aeb17b, 32'h41a88047, 32'hc21fc352, 32'h42853109};
test_output[18704:18711] = '{32'h4124b772, 32'h0, 32'h0, 32'h0, 32'h42aeb17b, 32'h41a88047, 32'h0, 32'h42853109};
test_input[18712:18719] = '{32'hc2269e6f, 32'h41b52ebf, 32'h42a872e9, 32'h42c0c022, 32'hc29f9334, 32'h41dc7c37, 32'hc1e97de0, 32'h42a3ac7c};
test_output[18712:18719] = '{32'h0, 32'h41b52ebf, 32'h42a872e9, 32'h42c0c022, 32'h0, 32'h41dc7c37, 32'h0, 32'h42a3ac7c};
test_input[18720:18727] = '{32'h41971b2a, 32'hc2abdd86, 32'h40cf1d71, 32'hc2878106, 32'hc0d475f6, 32'hc2c43499, 32'hc1e46dcb, 32'hc29ebf8b};
test_output[18720:18727] = '{32'h41971b2a, 32'h0, 32'h40cf1d71, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18728:18735] = '{32'hc2c0264d, 32'h425aefd8, 32'h40e70861, 32'h421da5ef, 32'h41a4a967, 32'hc10b4c43, 32'h42acbf30, 32'h4241e49e};
test_output[18728:18735] = '{32'h0, 32'h425aefd8, 32'h40e70861, 32'h421da5ef, 32'h41a4a967, 32'h0, 32'h42acbf30, 32'h4241e49e};
test_input[18736:18743] = '{32'hc28074cb, 32'h42595857, 32'h42af1f7f, 32'hc25cbd87, 32'h4024a0ff, 32'hc25632f5, 32'hc16de108, 32'h4287e9b5};
test_output[18736:18743] = '{32'h0, 32'h42595857, 32'h42af1f7f, 32'h0, 32'h4024a0ff, 32'h0, 32'h0, 32'h4287e9b5};
test_input[18744:18751] = '{32'hc2ac4441, 32'hc25e10d1, 32'h428e6fd2, 32'h423f83e2, 32'h41ea1c16, 32'hc2b0a964, 32'hc20bf381, 32'h4271ef98};
test_output[18744:18751] = '{32'h0, 32'h0, 32'h428e6fd2, 32'h423f83e2, 32'h41ea1c16, 32'h0, 32'h0, 32'h4271ef98};
test_input[18752:18759] = '{32'h428f1180, 32'hc2a59c4d, 32'h41fc33a3, 32'h42a23168, 32'h420bd3bf, 32'hc2b530a3, 32'h4255482a, 32'hc2addba6};
test_output[18752:18759] = '{32'h428f1180, 32'h0, 32'h41fc33a3, 32'h42a23168, 32'h420bd3bf, 32'h0, 32'h4255482a, 32'h0};
test_input[18760:18767] = '{32'h416f579d, 32'h42bcebd7, 32'hc294f1a7, 32'hc1f78e4c, 32'hc21ccf9c, 32'hc286123c, 32'hc29899fc, 32'hc17e30d8};
test_output[18760:18767] = '{32'h416f579d, 32'h42bcebd7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18768:18775] = '{32'h4291b42f, 32'h40de2134, 32'h41cfaec5, 32'h42a60093, 32'h42236f61, 32'hc27e5d4d, 32'h4288434f, 32'hc26b7fdb};
test_output[18768:18775] = '{32'h4291b42f, 32'h40de2134, 32'h41cfaec5, 32'h42a60093, 32'h42236f61, 32'h0, 32'h4288434f, 32'h0};
test_input[18776:18783] = '{32'h4245d95a, 32'hc294bff7, 32'h4213ba72, 32'hc2bb5032, 32'h428739f9, 32'h40cd33c8, 32'hc1fd56e4, 32'hc2c200ce};
test_output[18776:18783] = '{32'h4245d95a, 32'h0, 32'h4213ba72, 32'h0, 32'h428739f9, 32'h40cd33c8, 32'h0, 32'h0};
test_input[18784:18791] = '{32'h42425099, 32'hc2449279, 32'hc258a365, 32'hc292b7ab, 32'h40ce4029, 32'h429996b3, 32'h41ce7a79, 32'hc2505cab};
test_output[18784:18791] = '{32'h42425099, 32'h0, 32'h0, 32'h0, 32'h40ce4029, 32'h429996b3, 32'h41ce7a79, 32'h0};
test_input[18792:18799] = '{32'h42b1983a, 32'hc246d2f5, 32'hc2b4e6af, 32'h429ef711, 32'hc2bcd8c9, 32'h42a4c160, 32'h41e2571c, 32'hc2691b63};
test_output[18792:18799] = '{32'h42b1983a, 32'h0, 32'h0, 32'h429ef711, 32'h0, 32'h42a4c160, 32'h41e2571c, 32'h0};
test_input[18800:18807] = '{32'h428d3ecb, 32'hc28f9945, 32'h4202d5d2, 32'h42be3085, 32'h41d0f64f, 32'h4212eb7f, 32'h3f403cfe, 32'h418286c0};
test_output[18800:18807] = '{32'h428d3ecb, 32'h0, 32'h4202d5d2, 32'h42be3085, 32'h41d0f64f, 32'h4212eb7f, 32'h3f403cfe, 32'h418286c0};
test_input[18808:18815] = '{32'hc11f58ec, 32'hc2aa38c5, 32'h41e2388d, 32'hc2ba1612, 32'h429477a9, 32'hc2bafce3, 32'hc1ad78f1, 32'hc15e6cd4};
test_output[18808:18815] = '{32'h0, 32'h0, 32'h41e2388d, 32'h0, 32'h429477a9, 32'h0, 32'h0, 32'h0};
test_input[18816:18823] = '{32'h4289de9b, 32'h4298dc55, 32'h426c76cd, 32'hc01fc614, 32'h420a2720, 32'h42bc40e6, 32'hc28b8906, 32'h415aafed};
test_output[18816:18823] = '{32'h4289de9b, 32'h4298dc55, 32'h426c76cd, 32'h0, 32'h420a2720, 32'h42bc40e6, 32'h0, 32'h415aafed};
test_input[18824:18831] = '{32'hc28e9145, 32'hc24a82ff, 32'h41bfa6df, 32'hc1de387c, 32'h429eced4, 32'hbf83af76, 32'h4225f3bc, 32'hc287d672};
test_output[18824:18831] = '{32'h0, 32'h0, 32'h41bfa6df, 32'h0, 32'h429eced4, 32'h0, 32'h4225f3bc, 32'h0};
test_input[18832:18839] = '{32'hc0e23fb6, 32'hc19c1ed4, 32'hc2bfb929, 32'h42a8d1e1, 32'h41ec3de1, 32'h417bf243, 32'hc261d3e3, 32'hc213d02a};
test_output[18832:18839] = '{32'h0, 32'h0, 32'h0, 32'h42a8d1e1, 32'h41ec3de1, 32'h417bf243, 32'h0, 32'h0};
test_input[18840:18847] = '{32'hc285f59f, 32'h4293f3c6, 32'hc1a60668, 32'hc2087c3d, 32'hc14eae2b, 32'hc195c775, 32'hc299486e, 32'hc0259714};
test_output[18840:18847] = '{32'h0, 32'h4293f3c6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[18848:18855] = '{32'hc1ffbb99, 32'hc13acb83, 32'hc268dad6, 32'h41f8fde7, 32'hc23a6532, 32'hc1e1ad62, 32'hc2ae14aa, 32'h42bd3a99};
test_output[18848:18855] = '{32'h0, 32'h0, 32'h0, 32'h41f8fde7, 32'h0, 32'h0, 32'h0, 32'h42bd3a99};
test_input[18856:18863] = '{32'h429b24e1, 32'h42a87b89, 32'hc29eff51, 32'h4113d592, 32'h41a0fc5b, 32'hc231b281, 32'h42999c82, 32'h41399c02};
test_output[18856:18863] = '{32'h429b24e1, 32'h42a87b89, 32'h0, 32'h4113d592, 32'h41a0fc5b, 32'h0, 32'h42999c82, 32'h41399c02};
test_input[18864:18871] = '{32'hc013039e, 32'h4290a601, 32'hc2b8a2a2, 32'hc27ea6dc, 32'hc27881e7, 32'hc2c23606, 32'h42712c26, 32'h42a24ac6};
test_output[18864:18871] = '{32'h0, 32'h4290a601, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42712c26, 32'h42a24ac6};
test_input[18872:18879] = '{32'h41975dda, 32'hc2277878, 32'h4142308a, 32'h40a1698d, 32'hc223c6eb, 32'h42012224, 32'h41841cee, 32'h41937103};
test_output[18872:18879] = '{32'h41975dda, 32'h0, 32'h4142308a, 32'h40a1698d, 32'h0, 32'h42012224, 32'h41841cee, 32'h41937103};
test_input[18880:18887] = '{32'hc227d65e, 32'hc1023381, 32'h42991159, 32'h424b4e6a, 32'hc2a6ac68, 32'hc28507db, 32'h41d700ad, 32'h41958da5};
test_output[18880:18887] = '{32'h0, 32'h0, 32'h42991159, 32'h424b4e6a, 32'h0, 32'h0, 32'h41d700ad, 32'h41958da5};
test_input[18888:18895] = '{32'hc24aeece, 32'h42390a1c, 32'h42393224, 32'hc1ca0330, 32'hc2265cdf, 32'h41cd5ac0, 32'h428db966, 32'h4211bd0b};
test_output[18888:18895] = '{32'h0, 32'h42390a1c, 32'h42393224, 32'h0, 32'h0, 32'h41cd5ac0, 32'h428db966, 32'h4211bd0b};
test_input[18896:18903] = '{32'hc2baf366, 32'h41a0546d, 32'hc2894519, 32'h41b97e8b, 32'hc134b9e3, 32'h4264172a, 32'h41714a98, 32'h42ad8684};
test_output[18896:18903] = '{32'h0, 32'h41a0546d, 32'h0, 32'h41b97e8b, 32'h0, 32'h4264172a, 32'h41714a98, 32'h42ad8684};
test_input[18904:18911] = '{32'h411d6a8b, 32'h42b8ea6f, 32'h41076fbb, 32'hc2a19e71, 32'h3fc8f9e7, 32'hc169f9df, 32'h42ad09eb, 32'hc0d9b8ca};
test_output[18904:18911] = '{32'h411d6a8b, 32'h42b8ea6f, 32'h41076fbb, 32'h0, 32'h3fc8f9e7, 32'h0, 32'h42ad09eb, 32'h0};
test_input[18912:18919] = '{32'h42915f25, 32'hc1a980d3, 32'h42461d61, 32'hc085ef24, 32'h425443bc, 32'hc248f29d, 32'hc1520c2d, 32'h41297084};
test_output[18912:18919] = '{32'h42915f25, 32'h0, 32'h42461d61, 32'h0, 32'h425443bc, 32'h0, 32'h0, 32'h41297084};
test_input[18920:18927] = '{32'hc2738a7b, 32'hc283802d, 32'h421ffc1c, 32'h429fe59f, 32'h429cbf66, 32'h42a6ec2e, 32'h4285d15b, 32'h412ed556};
test_output[18920:18927] = '{32'h0, 32'h0, 32'h421ffc1c, 32'h429fe59f, 32'h429cbf66, 32'h42a6ec2e, 32'h4285d15b, 32'h412ed556};
test_input[18928:18935] = '{32'h4273c229, 32'h42848a10, 32'hc2665efe, 32'hc262a855, 32'h429ce148, 32'hc254fca5, 32'h4238c3a7, 32'hc242a5d1};
test_output[18928:18935] = '{32'h4273c229, 32'h42848a10, 32'h0, 32'h0, 32'h429ce148, 32'h0, 32'h4238c3a7, 32'h0};
test_input[18936:18943] = '{32'h4233d42f, 32'hc238d571, 32'h41ee416d, 32'hc088152c, 32'h426663a1, 32'hc28bee27, 32'hc2756a90, 32'hc003c9fd};
test_output[18936:18943] = '{32'h4233d42f, 32'h0, 32'h41ee416d, 32'h0, 32'h426663a1, 32'h0, 32'h0, 32'h0};
test_input[18944:18951] = '{32'hc2bcb031, 32'hc20a3f6e, 32'hbf4cdccb, 32'hc2abcd0b, 32'h41913cf4, 32'h421f8b2a, 32'hc297157d, 32'h429690ef};
test_output[18944:18951] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41913cf4, 32'h421f8b2a, 32'h0, 32'h429690ef};
test_input[18952:18959] = '{32'h42724673, 32'hc19d892f, 32'h420a6ff4, 32'h4268cd4f, 32'h42badd5f, 32'h42827fa7, 32'h41ada7e7, 32'hc21e7a63};
test_output[18952:18959] = '{32'h42724673, 32'h0, 32'h420a6ff4, 32'h4268cd4f, 32'h42badd5f, 32'h42827fa7, 32'h41ada7e7, 32'h0};
test_input[18960:18967] = '{32'hc2420674, 32'h42686850, 32'hc1c3cdb8, 32'h420895ef, 32'hc2275412, 32'h42946c59, 32'h4291f48a, 32'hc25b1bbe};
test_output[18960:18967] = '{32'h0, 32'h42686850, 32'h0, 32'h420895ef, 32'h0, 32'h42946c59, 32'h4291f48a, 32'h0};
test_input[18968:18975] = '{32'hc2ab43e2, 32'h4293713e, 32'h409ea44a, 32'h41a09081, 32'hc244399f, 32'hc2763c6c, 32'h428c694c, 32'h41cfb562};
test_output[18968:18975] = '{32'h0, 32'h4293713e, 32'h409ea44a, 32'h41a09081, 32'h0, 32'h0, 32'h428c694c, 32'h41cfb562};
test_input[18976:18983] = '{32'h41c80fcd, 32'h42bfbb25, 32'hc1a7ecb4, 32'h422cd80f, 32'h4249d9d7, 32'h419f064a, 32'h416bb85a, 32'hc2522064};
test_output[18976:18983] = '{32'h41c80fcd, 32'h42bfbb25, 32'h0, 32'h422cd80f, 32'h4249d9d7, 32'h419f064a, 32'h416bb85a, 32'h0};
test_input[18984:18991] = '{32'h4201bbb3, 32'h42c53d2b, 32'hc161ae19, 32'hc0bd5a2e, 32'h41616a1b, 32'h42ad3d62, 32'h41bfffab, 32'h42b4ab21};
test_output[18984:18991] = '{32'h4201bbb3, 32'h42c53d2b, 32'h0, 32'h0, 32'h41616a1b, 32'h42ad3d62, 32'h41bfffab, 32'h42b4ab21};
test_input[18992:18999] = '{32'hc2bd2fab, 32'h427bba25, 32'h428c30d3, 32'h42c3be8a, 32'hc03486cf, 32'hc224b1c1, 32'h422e158e, 32'hc280f427};
test_output[18992:18999] = '{32'h0, 32'h427bba25, 32'h428c30d3, 32'h42c3be8a, 32'h0, 32'h0, 32'h422e158e, 32'h0};
test_input[19000:19007] = '{32'h42adc5ad, 32'hc27eeae7, 32'hc24f8d44, 32'hc2bf5753, 32'h42bd5565, 32'h4286e8ed, 32'hc25cdba3, 32'h4231066d};
test_output[19000:19007] = '{32'h42adc5ad, 32'h0, 32'h0, 32'h0, 32'h42bd5565, 32'h4286e8ed, 32'h0, 32'h4231066d};
test_input[19008:19015] = '{32'hc2961d0f, 32'hc2411a07, 32'hc2b8326e, 32'hc22eb585, 32'hc23cdf3c, 32'h4194d658, 32'h4273a79d, 32'hc1fcd1a7};
test_output[19008:19015] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4194d658, 32'h4273a79d, 32'h0};
test_input[19016:19023] = '{32'h42347509, 32'hc16651f0, 32'hc2131b45, 32'h42bc512a, 32'hc23e4d9d, 32'h42a9e4b6, 32'h42b1d5fa, 32'hc10101f6};
test_output[19016:19023] = '{32'h42347509, 32'h0, 32'h0, 32'h42bc512a, 32'h0, 32'h42a9e4b6, 32'h42b1d5fa, 32'h0};
test_input[19024:19031] = '{32'hc2866d93, 32'hc281d4f2, 32'hc1598234, 32'h42144944, 32'hc2471a17, 32'h423224d6, 32'hc28902f6, 32'hc22d6280};
test_output[19024:19031] = '{32'h0, 32'h0, 32'h0, 32'h42144944, 32'h0, 32'h423224d6, 32'h0, 32'h0};
test_input[19032:19039] = '{32'hc201cc3e, 32'hc28f49cd, 32'hc296b5b6, 32'h41a56471, 32'hc23c73ba, 32'hc1a40f19, 32'hbfbb7a8e, 32'hc28c8f2d};
test_output[19032:19039] = '{32'h0, 32'h0, 32'h0, 32'h41a56471, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19040:19047] = '{32'hc28e3c9d, 32'h428f3174, 32'hc1d2986e, 32'h42bf21a5, 32'hc2b84fd5, 32'hc25bfc2a, 32'h42886c5a, 32'hc1915b96};
test_output[19040:19047] = '{32'h0, 32'h428f3174, 32'h0, 32'h42bf21a5, 32'h0, 32'h0, 32'h42886c5a, 32'h0};
test_input[19048:19055] = '{32'h40adf942, 32'h41b781f7, 32'h412933b9, 32'h41735410, 32'hc206a98f, 32'hc290f5f5, 32'h42270da2, 32'hc28f35f7};
test_output[19048:19055] = '{32'h40adf942, 32'h41b781f7, 32'h412933b9, 32'h41735410, 32'h0, 32'h0, 32'h42270da2, 32'h0};
test_input[19056:19063] = '{32'h41b68620, 32'hc2a513a4, 32'hc280fd71, 32'h42859100, 32'h42a40915, 32'hc221fd08, 32'h4229f9b7, 32'hc231735b};
test_output[19056:19063] = '{32'h41b68620, 32'h0, 32'h0, 32'h42859100, 32'h42a40915, 32'h0, 32'h4229f9b7, 32'h0};
test_input[19064:19071] = '{32'h42bd660f, 32'hc1794115, 32'h401fbd47, 32'hc28ffec9, 32'hc2979c0a, 32'h40a7e746, 32'hc28edf3d, 32'h42c0c34d};
test_output[19064:19071] = '{32'h42bd660f, 32'h0, 32'h401fbd47, 32'h0, 32'h0, 32'h40a7e746, 32'h0, 32'h42c0c34d};
test_input[19072:19079] = '{32'hc1e24a47, 32'hc183a423, 32'h429304ba, 32'hc2c2db5a, 32'hc288d7e5, 32'h42ae765c, 32'hc0793fd0, 32'h421ccf76};
test_output[19072:19079] = '{32'h0, 32'h0, 32'h429304ba, 32'h0, 32'h0, 32'h42ae765c, 32'h0, 32'h421ccf76};
test_input[19080:19087] = '{32'h4279fb5d, 32'hc1bd36a9, 32'h42686f4e, 32'h429965a2, 32'hc2917df4, 32'h4168393b, 32'hc08cdcad, 32'h428fde03};
test_output[19080:19087] = '{32'h4279fb5d, 32'h0, 32'h42686f4e, 32'h429965a2, 32'h0, 32'h4168393b, 32'h0, 32'h428fde03};
test_input[19088:19095] = '{32'hc2a52930, 32'h42bd5905, 32'hc26575e5, 32'h41485df1, 32'h427f90e5, 32'h41d870b6, 32'h4239cbdc, 32'hc11f8e07};
test_output[19088:19095] = '{32'h0, 32'h42bd5905, 32'h0, 32'h41485df1, 32'h427f90e5, 32'h41d870b6, 32'h4239cbdc, 32'h0};
test_input[19096:19103] = '{32'h4281a885, 32'hc1b3657c, 32'h424cd1e0, 32'h42bd49ea, 32'h4297cb3d, 32'h4106a245, 32'hc2a7758a, 32'hc266aa7a};
test_output[19096:19103] = '{32'h4281a885, 32'h0, 32'h424cd1e0, 32'h42bd49ea, 32'h4297cb3d, 32'h4106a245, 32'h0, 32'h0};
test_input[19104:19111] = '{32'hc243554e, 32'hc25a04f3, 32'h41fd73cb, 32'hc29c5e36, 32'hc2c724b8, 32'h40625b0f, 32'hc0ca25b6, 32'hc22a4a49};
test_output[19104:19111] = '{32'h0, 32'h0, 32'h41fd73cb, 32'h0, 32'h0, 32'h40625b0f, 32'h0, 32'h0};
test_input[19112:19119] = '{32'hc299c6bd, 32'hc21b91fd, 32'hc293ac7c, 32'h424c48c1, 32'h40a68b78, 32'hc1eb6298, 32'h420373c3, 32'h425eb34e};
test_output[19112:19119] = '{32'h0, 32'h0, 32'h0, 32'h424c48c1, 32'h40a68b78, 32'h0, 32'h420373c3, 32'h425eb34e};
test_input[19120:19127] = '{32'hc2751b18, 32'h42c0ca69, 32'hc1ddef77, 32'hc2869415, 32'hc2be236e, 32'hc245c93a, 32'h41b5e96e, 32'h429c2123};
test_output[19120:19127] = '{32'h0, 32'h42c0ca69, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b5e96e, 32'h429c2123};
test_input[19128:19135] = '{32'h42833fb2, 32'h4297d089, 32'hc2463884, 32'h42c0a160, 32'h42aa57db, 32'hc2430066, 32'hc2c0b79e, 32'hc281f934};
test_output[19128:19135] = '{32'h42833fb2, 32'h4297d089, 32'h0, 32'h42c0a160, 32'h42aa57db, 32'h0, 32'h0, 32'h0};
test_input[19136:19143] = '{32'hc1843cd5, 32'h428a62f6, 32'h42c73482, 32'hbfb575da, 32'hc29b08e8, 32'h420a5a8f, 32'hc285be36, 32'hc1239843};
test_output[19136:19143] = '{32'h0, 32'h428a62f6, 32'h42c73482, 32'h0, 32'h0, 32'h420a5a8f, 32'h0, 32'h0};
test_input[19144:19151] = '{32'hc2ae5a68, 32'h423fca8b, 32'h4226dc23, 32'hc27eb36e, 32'h4067864f, 32'h42c5fdfc, 32'hc014c285, 32'h4245b02c};
test_output[19144:19151] = '{32'h0, 32'h423fca8b, 32'h4226dc23, 32'h0, 32'h4067864f, 32'h42c5fdfc, 32'h0, 32'h4245b02c};
test_input[19152:19159] = '{32'hc23f8196, 32'h42a7de82, 32'h4281956c, 32'hc1f5fbe5, 32'h42253d31, 32'hc2745dfd, 32'h4270a74d, 32'hc26d423c};
test_output[19152:19159] = '{32'h0, 32'h42a7de82, 32'h4281956c, 32'h0, 32'h42253d31, 32'h0, 32'h4270a74d, 32'h0};
test_input[19160:19167] = '{32'hc236ece8, 32'hc2b41924, 32'hc2088a12, 32'hc211e0dd, 32'h42b98fe1, 32'hc2b1cf5e, 32'h42a91d45, 32'hc19a22ff};
test_output[19160:19167] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42b98fe1, 32'h0, 32'h42a91d45, 32'h0};
test_input[19168:19175] = '{32'h42aaaeae, 32'h426fbd0e, 32'h425030a6, 32'h42aa3733, 32'hc2af45ff, 32'hc2c48a99, 32'h42359527, 32'hc26d6d9a};
test_output[19168:19175] = '{32'h42aaaeae, 32'h426fbd0e, 32'h425030a6, 32'h42aa3733, 32'h0, 32'h0, 32'h42359527, 32'h0};
test_input[19176:19183] = '{32'hc2a8faec, 32'h425af0a3, 32'h4201ef6a, 32'h4241ba59, 32'h4185265b, 32'hc13e6378, 32'h42ad0dab, 32'h42a8dbea};
test_output[19176:19183] = '{32'h0, 32'h425af0a3, 32'h4201ef6a, 32'h4241ba59, 32'h4185265b, 32'h0, 32'h42ad0dab, 32'h42a8dbea};
test_input[19184:19191] = '{32'h42b1c8cd, 32'hc2bfc3aa, 32'hc1ac1d1b, 32'h426e80c5, 32'hc21f931b, 32'h42381b3b, 32'hc2ba92ec, 32'h41e2b419};
test_output[19184:19191] = '{32'h42b1c8cd, 32'h0, 32'h0, 32'h426e80c5, 32'h0, 32'h42381b3b, 32'h0, 32'h41e2b419};
test_input[19192:19199] = '{32'hc2378c7f, 32'h426a2728, 32'h429ebb8b, 32'hc2c2217d, 32'hc26446bf, 32'h424e8cd3, 32'h40b68c67, 32'h400c2d12};
test_output[19192:19199] = '{32'h0, 32'h426a2728, 32'h429ebb8b, 32'h0, 32'h0, 32'h424e8cd3, 32'h40b68c67, 32'h400c2d12};
test_input[19200:19207] = '{32'hc2838084, 32'h4234a1b5, 32'hc18fb777, 32'h413503ed, 32'h41791d50, 32'hc22223e5, 32'hc2964dbe, 32'hc2b2a415};
test_output[19200:19207] = '{32'h0, 32'h4234a1b5, 32'h0, 32'h413503ed, 32'h41791d50, 32'h0, 32'h0, 32'h0};
test_input[19208:19215] = '{32'hc23ef2a8, 32'hc12dcce2, 32'hc2ad6dc4, 32'hc07f1536, 32'h42696936, 32'h41bf84c0, 32'h42a56853, 32'hc246de3e};
test_output[19208:19215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42696936, 32'h41bf84c0, 32'h42a56853, 32'h0};
test_input[19216:19223] = '{32'h42b36056, 32'h41f11b01, 32'h429c532a, 32'h42a81e78, 32'h4291be8e, 32'hc298e3e1, 32'h4225aa5c, 32'hc2b801be};
test_output[19216:19223] = '{32'h42b36056, 32'h41f11b01, 32'h429c532a, 32'h42a81e78, 32'h4291be8e, 32'h0, 32'h4225aa5c, 32'h0};
test_input[19224:19231] = '{32'hc26fe628, 32'h41216776, 32'h422d654b, 32'h428c2a17, 32'hc2531792, 32'hc226205a, 32'h429d8ee2, 32'h420fcfa8};
test_output[19224:19231] = '{32'h0, 32'h41216776, 32'h422d654b, 32'h428c2a17, 32'h0, 32'h0, 32'h429d8ee2, 32'h420fcfa8};
test_input[19232:19239] = '{32'h42bd337f, 32'hc0183bab, 32'h42214aac, 32'h429a61be, 32'hc118c0ec, 32'h421b206b, 32'h42be1eea, 32'h425c2f62};
test_output[19232:19239] = '{32'h42bd337f, 32'h0, 32'h42214aac, 32'h429a61be, 32'h0, 32'h421b206b, 32'h42be1eea, 32'h425c2f62};
test_input[19240:19247] = '{32'hc2b5fe57, 32'hc2842a8c, 32'h4106bef4, 32'hc289a608, 32'h4217420a, 32'h41fdb9fe, 32'h42bfbd20, 32'hc2b8f77a};
test_output[19240:19247] = '{32'h0, 32'h0, 32'h4106bef4, 32'h0, 32'h4217420a, 32'h41fdb9fe, 32'h42bfbd20, 32'h0};
test_input[19248:19255] = '{32'h42b73307, 32'h42ab0d64, 32'h420c19b8, 32'hc24c000d, 32'h42c35bdf, 32'hbf697946, 32'h41053dde, 32'h42921980};
test_output[19248:19255] = '{32'h42b73307, 32'h42ab0d64, 32'h420c19b8, 32'h0, 32'h42c35bdf, 32'h0, 32'h41053dde, 32'h42921980};
test_input[19256:19263] = '{32'hc1a1c846, 32'h4212afa9, 32'h42c32eb3, 32'h42a11667, 32'hc20f4ae0, 32'hc237adf3, 32'hc260a74c, 32'h42b00125};
test_output[19256:19263] = '{32'h0, 32'h4212afa9, 32'h42c32eb3, 32'h42a11667, 32'h0, 32'h0, 32'h0, 32'h42b00125};
test_input[19264:19271] = '{32'hc28311a3, 32'hc2bdc49a, 32'hc18d12dd, 32'h415c748d, 32'hc1a93522, 32'hc201374e, 32'h42b592bb, 32'hc24d1d57};
test_output[19264:19271] = '{32'h0, 32'h0, 32'h0, 32'h415c748d, 32'h0, 32'h0, 32'h42b592bb, 32'h0};
test_input[19272:19279] = '{32'h419a5440, 32'hc2b770fc, 32'hc1b194b1, 32'h417ab1f9, 32'hc195f722, 32'hc288eea4, 32'hc268d206, 32'hc17587fb};
test_output[19272:19279] = '{32'h419a5440, 32'h0, 32'h0, 32'h417ab1f9, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19280:19287] = '{32'hc0c7edfe, 32'h4189b29e, 32'hc28b1d1f, 32'h416a2f82, 32'h42981efe, 32'h42794499, 32'hc2b0d8ae, 32'hc273d195};
test_output[19280:19287] = '{32'h0, 32'h4189b29e, 32'h0, 32'h416a2f82, 32'h42981efe, 32'h42794499, 32'h0, 32'h0};
test_input[19288:19295] = '{32'hc29d2768, 32'h428c8ed9, 32'h418d7f3b, 32'hc25373c1, 32'h418bc9b7, 32'hc2816c14, 32'h42a32629, 32'hc0bf51a5};
test_output[19288:19295] = '{32'h0, 32'h428c8ed9, 32'h418d7f3b, 32'h0, 32'h418bc9b7, 32'h0, 32'h42a32629, 32'h0};
test_input[19296:19303] = '{32'h41afe2af, 32'hc24c11eb, 32'h428e1641, 32'hc24dcfd0, 32'h423c14f5, 32'hc284a2f8, 32'h426da19c, 32'h4265c1b6};
test_output[19296:19303] = '{32'h41afe2af, 32'h0, 32'h428e1641, 32'h0, 32'h423c14f5, 32'h0, 32'h426da19c, 32'h4265c1b6};
test_input[19304:19311] = '{32'h42a9be37, 32'h4287dc94, 32'hc1f1c92b, 32'h42acbb49, 32'hc2ab19f0, 32'hc20d4c13, 32'hc126f83d, 32'h41e125fc};
test_output[19304:19311] = '{32'h42a9be37, 32'h4287dc94, 32'h0, 32'h42acbb49, 32'h0, 32'h0, 32'h0, 32'h41e125fc};
test_input[19312:19319] = '{32'hc1b0e7a2, 32'h428ba625, 32'h42c781af, 32'h41e36c30, 32'hc2610ef8, 32'hc1124f5b, 32'h418107c9, 32'h41568053};
test_output[19312:19319] = '{32'h0, 32'h428ba625, 32'h42c781af, 32'h41e36c30, 32'h0, 32'h0, 32'h418107c9, 32'h41568053};
test_input[19320:19327] = '{32'h41c8a114, 32'hc2886835, 32'hc284c7f9, 32'hc2b21861, 32'h42585509, 32'hc2b011bd, 32'h428e5656, 32'hc0b03ced};
test_output[19320:19327] = '{32'h41c8a114, 32'h0, 32'h0, 32'h0, 32'h42585509, 32'h0, 32'h428e5656, 32'h0};
test_input[19328:19335] = '{32'hc1f55787, 32'hc2a2edc5, 32'hc24a0f12, 32'hc2446c70, 32'hc1b07bef, 32'h42102b77, 32'hc25be2ca, 32'h4168ed0c};
test_output[19328:19335] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42102b77, 32'h0, 32'h4168ed0c};
test_input[19336:19343] = '{32'h4299becc, 32'hc283f418, 32'h428b35cb, 32'h42ab33b3, 32'hc171fe22, 32'hc2271d5a, 32'hc29ea6cf, 32'h41c33b8a};
test_output[19336:19343] = '{32'h4299becc, 32'h0, 32'h428b35cb, 32'h42ab33b3, 32'h0, 32'h0, 32'h0, 32'h41c33b8a};
test_input[19344:19351] = '{32'h4209dd35, 32'h426eef17, 32'h42a98f83, 32'hc192608d, 32'h4204175a, 32'hc2c796a2, 32'h41154087, 32'h422f3ea9};
test_output[19344:19351] = '{32'h4209dd35, 32'h426eef17, 32'h42a98f83, 32'h0, 32'h4204175a, 32'h0, 32'h41154087, 32'h422f3ea9};
test_input[19352:19359] = '{32'h4104d943, 32'hc22e5bad, 32'hc24b7175, 32'h4195a689, 32'h4207a9e6, 32'h42b58357, 32'h423857f6, 32'h4278c336};
test_output[19352:19359] = '{32'h4104d943, 32'h0, 32'h0, 32'h4195a689, 32'h4207a9e6, 32'h42b58357, 32'h423857f6, 32'h4278c336};
test_input[19360:19367] = '{32'hc2807887, 32'hc25585c3, 32'h428da027, 32'hbdea7944, 32'h42944885, 32'hc2913213, 32'h4135618c, 32'h40861e02};
test_output[19360:19367] = '{32'h0, 32'h0, 32'h428da027, 32'h0, 32'h42944885, 32'h0, 32'h4135618c, 32'h40861e02};
test_input[19368:19375] = '{32'h421e52de, 32'h42bf0ca5, 32'h42abe341, 32'h42be7ef0, 32'hc1fa6566, 32'h4299e8bb, 32'hc1ef11cd, 32'h4215f008};
test_output[19368:19375] = '{32'h421e52de, 32'h42bf0ca5, 32'h42abe341, 32'h42be7ef0, 32'h0, 32'h4299e8bb, 32'h0, 32'h4215f008};
test_input[19376:19383] = '{32'hc259b66e, 32'hc223001e, 32'h42451e2d, 32'hc2b645e8, 32'h42a117f0, 32'hc1349617, 32'h41a2993b, 32'hbf31a0f1};
test_output[19376:19383] = '{32'h0, 32'h0, 32'h42451e2d, 32'h0, 32'h42a117f0, 32'h0, 32'h41a2993b, 32'h0};
test_input[19384:19391] = '{32'hc26f2f0c, 32'h4287f417, 32'hc28be904, 32'h4201de12, 32'h426e5e74, 32'hc234b40e, 32'h4162e291, 32'hc25b8a51};
test_output[19384:19391] = '{32'h0, 32'h4287f417, 32'h0, 32'h4201de12, 32'h426e5e74, 32'h0, 32'h4162e291, 32'h0};
test_input[19392:19399] = '{32'hc2bd5b6d, 32'hc1bd4a7c, 32'h42a88705, 32'h4150eb5d, 32'hc0856bad, 32'h42bc18b0, 32'h42bd4337, 32'hc119a1d6};
test_output[19392:19399] = '{32'h0, 32'h0, 32'h42a88705, 32'h4150eb5d, 32'h0, 32'h42bc18b0, 32'h42bd4337, 32'h0};
test_input[19400:19407] = '{32'h40c5fce8, 32'h42437268, 32'h426e7dda, 32'hc2ab5621, 32'hc0ca06d0, 32'h40dfe9cd, 32'h428d8752, 32'hbf9330bd};
test_output[19400:19407] = '{32'h40c5fce8, 32'h42437268, 32'h426e7dda, 32'h0, 32'h0, 32'h40dfe9cd, 32'h428d8752, 32'h0};
test_input[19408:19415] = '{32'hc1a71f27, 32'hc2a33c7e, 32'h402111f0, 32'hc017d878, 32'h41f6dcef, 32'h41b3aa69, 32'h4263825b, 32'hc20e8b6e};
test_output[19408:19415] = '{32'h0, 32'h0, 32'h402111f0, 32'h0, 32'h41f6dcef, 32'h41b3aa69, 32'h4263825b, 32'h0};
test_input[19416:19423] = '{32'hc2b4438f, 32'h42952ad2, 32'h42667ade, 32'h42a128d2, 32'hc1d959e6, 32'h4272d9a6, 32'h425b64f6, 32'h409bf1aa};
test_output[19416:19423] = '{32'h0, 32'h42952ad2, 32'h42667ade, 32'h42a128d2, 32'h0, 32'h4272d9a6, 32'h425b64f6, 32'h409bf1aa};
test_input[19424:19431] = '{32'hc2ac2c12, 32'h4210994a, 32'hc2b55efb, 32'hc23ccf3c, 32'h42bc3730, 32'hc29f27a8, 32'h425cb974, 32'hc2877e8a};
test_output[19424:19431] = '{32'h0, 32'h4210994a, 32'h0, 32'h0, 32'h42bc3730, 32'h0, 32'h425cb974, 32'h0};
test_input[19432:19439] = '{32'hc14cb888, 32'h42c6f40d, 32'hc253a1c3, 32'h42161aa4, 32'hc1fba47d, 32'hc20b1182, 32'hc21e5ec1, 32'h4216cef7};
test_output[19432:19439] = '{32'h0, 32'h42c6f40d, 32'h0, 32'h42161aa4, 32'h0, 32'h0, 32'h0, 32'h4216cef7};
test_input[19440:19447] = '{32'hc2338e67, 32'h4217450c, 32'h422e3d74, 32'h4233d03e, 32'hc288951f, 32'h422529f1, 32'h42bd3648, 32'hc211a5b1};
test_output[19440:19447] = '{32'h0, 32'h4217450c, 32'h422e3d74, 32'h4233d03e, 32'h0, 32'h422529f1, 32'h42bd3648, 32'h0};
test_input[19448:19455] = '{32'hc2b3f334, 32'h42b16b8e, 32'h42ad595a, 32'hc2a0a447, 32'hc2a00af2, 32'h42b99873, 32'h4196e928, 32'h42312127};
test_output[19448:19455] = '{32'h0, 32'h42b16b8e, 32'h42ad595a, 32'h0, 32'h0, 32'h42b99873, 32'h4196e928, 32'h42312127};
test_input[19456:19463] = '{32'h41b87997, 32'hc2102e7a, 32'h420766da, 32'hc29cc3f0, 32'h42c2874b, 32'h42ae21dd, 32'hc23339b3, 32'h41fa0908};
test_output[19456:19463] = '{32'h41b87997, 32'h0, 32'h420766da, 32'h0, 32'h42c2874b, 32'h42ae21dd, 32'h0, 32'h41fa0908};
test_input[19464:19471] = '{32'h42c5677b, 32'h428c5ed3, 32'hc108525d, 32'hc1e789aa, 32'h426910f4, 32'hc2beb27c, 32'h419643f1, 32'h4185bf3c};
test_output[19464:19471] = '{32'h42c5677b, 32'h428c5ed3, 32'h0, 32'h0, 32'h426910f4, 32'h0, 32'h419643f1, 32'h4185bf3c};
test_input[19472:19479] = '{32'h413dbbdd, 32'hc24fa54c, 32'h42808085, 32'hc146fb75, 32'h420962cf, 32'h4293a1fb, 32'h42218b51, 32'hc1e1ccad};
test_output[19472:19479] = '{32'h413dbbdd, 32'h0, 32'h42808085, 32'h0, 32'h420962cf, 32'h4293a1fb, 32'h42218b51, 32'h0};
test_input[19480:19487] = '{32'h42bf49f1, 32'hc1a78bfe, 32'h42029cef, 32'hc209a6d9, 32'h41991f18, 32'h429e4c5d, 32'h3e8925a4, 32'h4248b0c8};
test_output[19480:19487] = '{32'h42bf49f1, 32'h0, 32'h42029cef, 32'h0, 32'h41991f18, 32'h429e4c5d, 32'h3e8925a4, 32'h4248b0c8};
test_input[19488:19495] = '{32'hc2b6357a, 32'h42895ffa, 32'hc224bea7, 32'hc1c1ccb0, 32'h411774ea, 32'hc2a734c9, 32'h427be2e3, 32'hc2b322a9};
test_output[19488:19495] = '{32'h0, 32'h42895ffa, 32'h0, 32'h0, 32'h411774ea, 32'h0, 32'h427be2e3, 32'h0};
test_input[19496:19503] = '{32'hc2c7f3e8, 32'hc22903aa, 32'h42678bf4, 32'h41f5ac85, 32'h418c7a03, 32'hc19ed7bb, 32'hc29170b8, 32'hc1d2951f};
test_output[19496:19503] = '{32'h0, 32'h0, 32'h42678bf4, 32'h41f5ac85, 32'h418c7a03, 32'h0, 32'h0, 32'h0};
test_input[19504:19511] = '{32'hc2557cc9, 32'h420f4030, 32'h40d0e9ec, 32'h41b4996f, 32'h4289c40d, 32'h42beca60, 32'hc24b7d84, 32'hc2a03af3};
test_output[19504:19511] = '{32'h0, 32'h420f4030, 32'h40d0e9ec, 32'h41b4996f, 32'h4289c40d, 32'h42beca60, 32'h0, 32'h0};
test_input[19512:19519] = '{32'h4239ee91, 32'hc2a3911b, 32'h4290353e, 32'hc27e8194, 32'hc272a335, 32'hc0845c61, 32'hc28b1b60, 32'hc2b62c73};
test_output[19512:19519] = '{32'h4239ee91, 32'h0, 32'h4290353e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19520:19527] = '{32'hc292825a, 32'h42b8caa2, 32'hc29f6361, 32'h422ecdb8, 32'hc2b9f88b, 32'hc2b9131a, 32'h42088e22, 32'h42887428};
test_output[19520:19527] = '{32'h0, 32'h42b8caa2, 32'h0, 32'h422ecdb8, 32'h0, 32'h0, 32'h42088e22, 32'h42887428};
test_input[19528:19535] = '{32'hc29380fc, 32'hc24eee34, 32'hc200fa81, 32'h42545d3c, 32'hc0e36158, 32'hc10247a3, 32'h42a064ce, 32'h426c1ee1};
test_output[19528:19535] = '{32'h0, 32'h0, 32'h0, 32'h42545d3c, 32'h0, 32'h0, 32'h42a064ce, 32'h426c1ee1};
test_input[19536:19543] = '{32'hc1d2156a, 32'h41d1fbab, 32'h427cf579, 32'hc1ae5a11, 32'h426fd2ea, 32'h42a0714a, 32'h420274ce, 32'h42052556};
test_output[19536:19543] = '{32'h0, 32'h41d1fbab, 32'h427cf579, 32'h0, 32'h426fd2ea, 32'h42a0714a, 32'h420274ce, 32'h42052556};
test_input[19544:19551] = '{32'hc0e11b7c, 32'h426c0e5c, 32'hc29aae0e, 32'hbf63d741, 32'h4160fd8b, 32'hc07fa59d, 32'hc2ab18ad, 32'h42669c47};
test_output[19544:19551] = '{32'h0, 32'h426c0e5c, 32'h0, 32'h0, 32'h4160fd8b, 32'h0, 32'h0, 32'h42669c47};
test_input[19552:19559] = '{32'hc2b44c2c, 32'h42251c50, 32'hc2afc34f, 32'hc24f470e, 32'hbfa5bb34, 32'hc20b90e8, 32'h4190db65, 32'h42a446e4};
test_output[19552:19559] = '{32'h0, 32'h42251c50, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4190db65, 32'h42a446e4};
test_input[19560:19567] = '{32'hc2c13406, 32'hc20e8ce1, 32'h42858388, 32'h4125410c, 32'h422b1a43, 32'hc2035314, 32'h4283f4d8, 32'hc2a11394};
test_output[19560:19567] = '{32'h0, 32'h0, 32'h42858388, 32'h4125410c, 32'h422b1a43, 32'h0, 32'h4283f4d8, 32'h0};
test_input[19568:19575] = '{32'hc28f392b, 32'h423a0637, 32'hc21c5994, 32'hc1a654a9, 32'h4039db08, 32'hc22bd154, 32'hc2a4e861, 32'h428468cb};
test_output[19568:19575] = '{32'h0, 32'h423a0637, 32'h0, 32'h0, 32'h4039db08, 32'h0, 32'h0, 32'h428468cb};
test_input[19576:19583] = '{32'hc274557e, 32'hc25739cb, 32'hc137bde3, 32'h429d40b2, 32'hc169412b, 32'hc1c2def9, 32'hc24a4075, 32'hc2bceaec};
test_output[19576:19583] = '{32'h0, 32'h0, 32'h0, 32'h429d40b2, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19584:19591] = '{32'h4187507f, 32'h417e91bb, 32'h410b229f, 32'h41946b0f, 32'hc299cf9c, 32'hc21ef7db, 32'h428ac4d3, 32'hc2bb0a77};
test_output[19584:19591] = '{32'h4187507f, 32'h417e91bb, 32'h410b229f, 32'h41946b0f, 32'h0, 32'h0, 32'h428ac4d3, 32'h0};
test_input[19592:19599] = '{32'h425a4fe4, 32'hc2474b55, 32'hc298b85f, 32'hc2bdf6bd, 32'hc14d1b11, 32'hc2a67650, 32'hc1cb2597, 32'hc1a4eb01};
test_output[19592:19599] = '{32'h425a4fe4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19600:19607] = '{32'hc27d5331, 32'hc2813e4e, 32'hc2951cda, 32'hc2c3a3ce, 32'hc231fa14, 32'h41b8d562, 32'h42bd26d7, 32'hc21fc8a5};
test_output[19600:19607] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b8d562, 32'h42bd26d7, 32'h0};
test_input[19608:19615] = '{32'hc27380dc, 32'hc2b7d125, 32'h41935d6f, 32'h42169d87, 32'h420d1210, 32'h4104fdf9, 32'hc17919b9, 32'h422135a8};
test_output[19608:19615] = '{32'h0, 32'h0, 32'h41935d6f, 32'h42169d87, 32'h420d1210, 32'h4104fdf9, 32'h0, 32'h422135a8};
test_input[19616:19623] = '{32'h425d21cc, 32'hc2b6d866, 32'h41d8e8d6, 32'hc21a9468, 32'h42334d09, 32'h42c42479, 32'hc2b19ab5, 32'hc1aa0e96};
test_output[19616:19623] = '{32'h425d21cc, 32'h0, 32'h41d8e8d6, 32'h0, 32'h42334d09, 32'h42c42479, 32'h0, 32'h0};
test_input[19624:19631] = '{32'h42a5bfeb, 32'hc29c8ac5, 32'h42906a5e, 32'h4272bb03, 32'hc22c7d82, 32'h428d7db6, 32'hc2ba5777, 32'h4241a028};
test_output[19624:19631] = '{32'h42a5bfeb, 32'h0, 32'h42906a5e, 32'h4272bb03, 32'h0, 32'h428d7db6, 32'h0, 32'h4241a028};
test_input[19632:19639] = '{32'hc2956043, 32'hc20edbf2, 32'hc2ad1f02, 32'hc26abc96, 32'hc2b3290d, 32'hc2c740d5, 32'hc090524d, 32'hc2006d78};
test_output[19632:19639] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19640:19647] = '{32'hc2a01c0c, 32'h42b9b96b, 32'h42b62e2d, 32'hc1a202d9, 32'h428aae25, 32'h428c0121, 32'h4276a928, 32'h42b8522f};
test_output[19640:19647] = '{32'h0, 32'h42b9b96b, 32'h42b62e2d, 32'h0, 32'h428aae25, 32'h428c0121, 32'h4276a928, 32'h42b8522f};
test_input[19648:19655] = '{32'hc1cd3260, 32'hc293f62b, 32'hc19a4eb5, 32'h41f40b70, 32'h42a74af1, 32'h423bd86e, 32'hc2c09dcd, 32'hc2b0a864};
test_output[19648:19655] = '{32'h0, 32'h0, 32'h0, 32'h41f40b70, 32'h42a74af1, 32'h423bd86e, 32'h0, 32'h0};
test_input[19656:19663] = '{32'h42ae2799, 32'h425368b3, 32'hc263028d, 32'hc1ac86ac, 32'h429ff4e7, 32'hc1b4fdfc, 32'hc2c2638c, 32'hc2088bef};
test_output[19656:19663] = '{32'h42ae2799, 32'h425368b3, 32'h0, 32'h0, 32'h429ff4e7, 32'h0, 32'h0, 32'h0};
test_input[19664:19671] = '{32'hc296c47d, 32'hc29af253, 32'hc14dd9ee, 32'hc24ba08c, 32'hc29d221f, 32'h429f0e70, 32'hc0874800, 32'hc12b71cb};
test_output[19664:19671] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429f0e70, 32'h0, 32'h0};
test_input[19672:19679] = '{32'hc2bd47ba, 32'hc23ca64c, 32'hc199e005, 32'hc131cbea, 32'hc0fa2f6a, 32'hc27f111c, 32'h42a3bf40, 32'hc2a46da1};
test_output[19672:19679] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a3bf40, 32'h0};
test_input[19680:19687] = '{32'h4291a92a, 32'hc28ac7e4, 32'hc20559c6, 32'h421f62e4, 32'h42629c51, 32'h401fbdac, 32'h424c4bcf, 32'h41b49fcc};
test_output[19680:19687] = '{32'h4291a92a, 32'h0, 32'h0, 32'h421f62e4, 32'h42629c51, 32'h401fbdac, 32'h424c4bcf, 32'h41b49fcc};
test_input[19688:19695] = '{32'h41b247d0, 32'h428d2357, 32'h40ea0edf, 32'hc21a15fe, 32'hc09440a2, 32'h41d4be35, 32'h4249ed4f, 32'h42157462};
test_output[19688:19695] = '{32'h41b247d0, 32'h428d2357, 32'h40ea0edf, 32'h0, 32'h0, 32'h41d4be35, 32'h4249ed4f, 32'h42157462};
test_input[19696:19703] = '{32'hc28eb32d, 32'h4275e440, 32'hc2767240, 32'hc233e574, 32'hc287cfd8, 32'hc2a4d726, 32'hc2986cd9, 32'hc2a62bdc};
test_output[19696:19703] = '{32'h0, 32'h4275e440, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19704:19711] = '{32'h42710e5f, 32'h42814b16, 32'hc16e559f, 32'h41f99ba8, 32'hc2a642ad, 32'hc2ab95b8, 32'h42bdde24, 32'h4272e8a3};
test_output[19704:19711] = '{32'h42710e5f, 32'h42814b16, 32'h0, 32'h41f99ba8, 32'h0, 32'h0, 32'h42bdde24, 32'h4272e8a3};
test_input[19712:19719] = '{32'h41ae4bbd, 32'hc28024a7, 32'h41162e3b, 32'h4291c969, 32'h42246c3e, 32'hc201abe5, 32'h428af7d7, 32'hc107ee30};
test_output[19712:19719] = '{32'h41ae4bbd, 32'h0, 32'h41162e3b, 32'h4291c969, 32'h42246c3e, 32'h0, 32'h428af7d7, 32'h0};
test_input[19720:19727] = '{32'hc1a227db, 32'h427c3937, 32'hc293e948, 32'h41084c93, 32'h42130e07, 32'h42827c11, 32'h410cc4c2, 32'hc28a18b0};
test_output[19720:19727] = '{32'h0, 32'h427c3937, 32'h0, 32'h41084c93, 32'h42130e07, 32'h42827c11, 32'h410cc4c2, 32'h0};
test_input[19728:19735] = '{32'hc28c96c4, 32'h42c2efd2, 32'h423c4b24, 32'h42411f02, 32'hc2a5ceb9, 32'hc19c4b34, 32'h42b75cfe, 32'h40d1865c};
test_output[19728:19735] = '{32'h0, 32'h42c2efd2, 32'h423c4b24, 32'h42411f02, 32'h0, 32'h0, 32'h42b75cfe, 32'h40d1865c};
test_input[19736:19743] = '{32'h420dc705, 32'h42b41c0a, 32'hc13e0e85, 32'h4231a982, 32'hc27e2e05, 32'hc2b2ff62, 32'hc29a977c, 32'hbf2f19b6};
test_output[19736:19743] = '{32'h420dc705, 32'h42b41c0a, 32'h0, 32'h4231a982, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19744:19751] = '{32'h42c2c047, 32'hc1ec9efd, 32'hc19a517d, 32'hc256cb6d, 32'h414cce5a, 32'h42a8ae4a, 32'hc25b0c32, 32'hc28b3095};
test_output[19744:19751] = '{32'h42c2c047, 32'h0, 32'h0, 32'h0, 32'h414cce5a, 32'h42a8ae4a, 32'h0, 32'h0};
test_input[19752:19759] = '{32'hc20cfef9, 32'h42b45e8a, 32'hc2c7bbf1, 32'h42bf515a, 32'h422ee5d4, 32'hc0f140b8, 32'hc2b136a6, 32'h42175e64};
test_output[19752:19759] = '{32'h0, 32'h42b45e8a, 32'h0, 32'h42bf515a, 32'h422ee5d4, 32'h0, 32'h0, 32'h42175e64};
test_input[19760:19767] = '{32'h42bf3aa3, 32'hc0aacd57, 32'h42b3c89f, 32'hc20e4170, 32'hc01111c4, 32'hc1a7b024, 32'hc1dba673, 32'hc29f1437};
test_output[19760:19767] = '{32'h42bf3aa3, 32'h0, 32'h42b3c89f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19768:19775] = '{32'h418494d1, 32'h41c06aa9, 32'h42ba7312, 32'h42768b2d, 32'h40102e17, 32'h40b03fe5, 32'hc2c7b4ac, 32'hc186320f};
test_output[19768:19775] = '{32'h418494d1, 32'h41c06aa9, 32'h42ba7312, 32'h42768b2d, 32'h40102e17, 32'h40b03fe5, 32'h0, 32'h0};
test_input[19776:19783] = '{32'hc24c533e, 32'hc29dc2bf, 32'h40853b05, 32'hc26c588e, 32'hc0c244ac, 32'h4228f8f9, 32'hc2139fa0, 32'h42582c3f};
test_output[19776:19783] = '{32'h0, 32'h0, 32'h40853b05, 32'h0, 32'h0, 32'h4228f8f9, 32'h0, 32'h42582c3f};
test_input[19784:19791] = '{32'hc16a367a, 32'h425ba315, 32'hc283d179, 32'hc292fff3, 32'hc2707dff, 32'hc2413cfd, 32'hc2bde3e8, 32'h42afb371};
test_output[19784:19791] = '{32'h0, 32'h425ba315, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42afb371};
test_input[19792:19799] = '{32'hc1c7542f, 32'hc22bde02, 32'hc2c0b85e, 32'h41acf930, 32'h423b35bf, 32'h41467265, 32'hc29094e8, 32'hc1fecfdf};
test_output[19792:19799] = '{32'h0, 32'h0, 32'h0, 32'h41acf930, 32'h423b35bf, 32'h41467265, 32'h0, 32'h0};
test_input[19800:19807] = '{32'h421427ea, 32'hc28b33e3, 32'hc2be3544, 32'hc2a296fa, 32'hc2b28560, 32'hc078ca06, 32'hc2a4858e, 32'hc2be7bb0};
test_output[19800:19807] = '{32'h421427ea, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19808:19815] = '{32'hc293eb87, 32'h42666fe4, 32'h424f0443, 32'h427f8ec6, 32'hc2620edc, 32'h41dab743, 32'h41d1762d, 32'h41e49139};
test_output[19808:19815] = '{32'h0, 32'h42666fe4, 32'h424f0443, 32'h427f8ec6, 32'h0, 32'h41dab743, 32'h41d1762d, 32'h41e49139};
test_input[19816:19823] = '{32'h4227934d, 32'hc2be64af, 32'h4230aa51, 32'hc29bbe77, 32'hc266264a, 32'hc2706a89, 32'hc23655a3, 32'hc2940d60};
test_output[19816:19823] = '{32'h4227934d, 32'h0, 32'h4230aa51, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[19824:19831] = '{32'hc2ae60d5, 32'h423cd14e, 32'h42a582cf, 32'h4241cbc5, 32'h3ff55cfb, 32'h42b81fda, 32'hc27c6b71, 32'hc29cd89f};
test_output[19824:19831] = '{32'h0, 32'h423cd14e, 32'h42a582cf, 32'h4241cbc5, 32'h3ff55cfb, 32'h42b81fda, 32'h0, 32'h0};
test_input[19832:19839] = '{32'h425e9b55, 32'h428f97c5, 32'h4187dacc, 32'h41ffaa75, 32'hc0f34da4, 32'hc21c65c4, 32'h417822b0, 32'hc1b84359};
test_output[19832:19839] = '{32'h425e9b55, 32'h428f97c5, 32'h4187dacc, 32'h41ffaa75, 32'h0, 32'h0, 32'h417822b0, 32'h0};
test_input[19840:19847] = '{32'hc2a25dc1, 32'hc25b758f, 32'h422829c9, 32'h416db065, 32'h4157ab3d, 32'hc282ea83, 32'hc11df160, 32'h42595d58};
test_output[19840:19847] = '{32'h0, 32'h0, 32'h422829c9, 32'h416db065, 32'h4157ab3d, 32'h0, 32'h0, 32'h42595d58};
test_input[19848:19855] = '{32'h4216ffa8, 32'h42abc6c5, 32'hc29cb5ea, 32'h4191fcc2, 32'h41c3b572, 32'hc2339b1b, 32'h422aca71, 32'hc1b9ace1};
test_output[19848:19855] = '{32'h4216ffa8, 32'h42abc6c5, 32'h0, 32'h4191fcc2, 32'h41c3b572, 32'h0, 32'h422aca71, 32'h0};
test_input[19856:19863] = '{32'h4210ba05, 32'hc2c418a1, 32'h41c796ae, 32'h4177d237, 32'hc21917f3, 32'h41c72519, 32'hc298392f, 32'hc2bf986d};
test_output[19856:19863] = '{32'h4210ba05, 32'h0, 32'h41c796ae, 32'h4177d237, 32'h0, 32'h41c72519, 32'h0, 32'h0};
test_input[19864:19871] = '{32'h41ee54ca, 32'h42b6e7bf, 32'h428b4c79, 32'h42c17c0c, 32'h4231ac3d, 32'h42603987, 32'h42278527, 32'hc241faf0};
test_output[19864:19871] = '{32'h41ee54ca, 32'h42b6e7bf, 32'h428b4c79, 32'h42c17c0c, 32'h4231ac3d, 32'h42603987, 32'h42278527, 32'h0};
test_input[19872:19879] = '{32'hc2c718c2, 32'h42aa7af2, 32'hc286fe84, 32'hc0ff265e, 32'hc2aa8f63, 32'h416e2d2c, 32'hc230d941, 32'hc09ae54c};
test_output[19872:19879] = '{32'h0, 32'h42aa7af2, 32'h0, 32'h0, 32'h0, 32'h416e2d2c, 32'h0, 32'h0};
test_input[19880:19887] = '{32'h424fc4dd, 32'h42389b30, 32'h42c16f7c, 32'h41dd1b59, 32'h42ba89e7, 32'hc255649a, 32'hc1efc752, 32'hc2248c1b};
test_output[19880:19887] = '{32'h424fc4dd, 32'h42389b30, 32'h42c16f7c, 32'h41dd1b59, 32'h42ba89e7, 32'h0, 32'h0, 32'h0};
test_input[19888:19895] = '{32'hc284aade, 32'hc275f4ef, 32'hc29171c5, 32'hc206c36d, 32'hc297646d, 32'hc252a4c0, 32'hc2169dc5, 32'h42ba81fd};
test_output[19888:19895] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ba81fd};
test_input[19896:19903] = '{32'hc2a29d21, 32'hbff53a36, 32'hc225617d, 32'h42b2ee73, 32'hc2bf471d, 32'hc210f48a, 32'h42067b06, 32'hc1c7ad62};
test_output[19896:19903] = '{32'h0, 32'h0, 32'h0, 32'h42b2ee73, 32'h0, 32'h0, 32'h42067b06, 32'h0};
test_input[19904:19911] = '{32'h41b0d01c, 32'h4162f2e7, 32'hc297d504, 32'h41df6dad, 32'h416c4e4d, 32'hc2806d14, 32'hc2a0e683, 32'hc18a2122};
test_output[19904:19911] = '{32'h41b0d01c, 32'h4162f2e7, 32'h0, 32'h41df6dad, 32'h416c4e4d, 32'h0, 32'h0, 32'h0};
test_input[19912:19919] = '{32'h418aade7, 32'hc05931fd, 32'h42185979, 32'h42a8f81e, 32'h42490857, 32'hc19baee0, 32'h42a20330, 32'hc1c4893d};
test_output[19912:19919] = '{32'h418aade7, 32'h0, 32'h42185979, 32'h42a8f81e, 32'h42490857, 32'h0, 32'h42a20330, 32'h0};
test_input[19920:19927] = '{32'hc201d1b8, 32'h4208ce8c, 32'hc1731607, 32'hc1e0eee0, 32'h41dd457b, 32'h42735086, 32'hc1bc285a, 32'h42153841};
test_output[19920:19927] = '{32'h0, 32'h4208ce8c, 32'h0, 32'h0, 32'h41dd457b, 32'h42735086, 32'h0, 32'h42153841};
test_input[19928:19935] = '{32'h4213890d, 32'hc29676df, 32'h42c0ca57, 32'h4287db21, 32'hc28e9726, 32'h4267e505, 32'h429fde1f, 32'h4183a39a};
test_output[19928:19935] = '{32'h4213890d, 32'h0, 32'h42c0ca57, 32'h4287db21, 32'h0, 32'h4267e505, 32'h429fde1f, 32'h4183a39a};
test_input[19936:19943] = '{32'h424e70da, 32'hc217f789, 32'h427ca8aa, 32'h41feaad1, 32'hc29f7e9b, 32'hc2ae7fb4, 32'h40ddfa54, 32'hc2802874};
test_output[19936:19943] = '{32'h424e70da, 32'h0, 32'h427ca8aa, 32'h41feaad1, 32'h0, 32'h0, 32'h40ddfa54, 32'h0};
test_input[19944:19951] = '{32'hc0ced32c, 32'hc27c4403, 32'hc1fe6153, 32'hc2166d89, 32'hc19e1820, 32'hc2a24412, 32'hc25d8b5a, 32'h423fd3df};
test_output[19944:19951] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423fd3df};
test_input[19952:19959] = '{32'h41d4b05b, 32'h4258f6ea, 32'h42735e96, 32'h42b3ffd2, 32'h418cf11c, 32'hc056fafb, 32'h412133a7, 32'hc2ab819c};
test_output[19952:19959] = '{32'h41d4b05b, 32'h4258f6ea, 32'h42735e96, 32'h42b3ffd2, 32'h418cf11c, 32'h0, 32'h412133a7, 32'h0};
test_input[19960:19967] = '{32'h4292d17b, 32'hc2c1a376, 32'h4094173e, 32'h40dbb518, 32'hc2a6f84e, 32'hc1968145, 32'hc2819677, 32'h426405a3};
test_output[19960:19967] = '{32'h4292d17b, 32'h0, 32'h4094173e, 32'h40dbb518, 32'h0, 32'h0, 32'h0, 32'h426405a3};
test_input[19968:19975] = '{32'h42c1e9a3, 32'h42562d7a, 32'hc26df69d, 32'h420dca53, 32'h422f75dd, 32'h427c5927, 32'h423dba38, 32'h423380a1};
test_output[19968:19975] = '{32'h42c1e9a3, 32'h42562d7a, 32'h0, 32'h420dca53, 32'h422f75dd, 32'h427c5927, 32'h423dba38, 32'h423380a1};
test_input[19976:19983] = '{32'h41fb2fa8, 32'hc0ca58eb, 32'hc239d306, 32'h41b0cf45, 32'h41748b14, 32'hc24483a6, 32'h41c33b9a, 32'h422ad156};
test_output[19976:19983] = '{32'h41fb2fa8, 32'h0, 32'h0, 32'h41b0cf45, 32'h41748b14, 32'h0, 32'h41c33b9a, 32'h422ad156};
test_input[19984:19991] = '{32'h41691d87, 32'h426a41c7, 32'hc2b7fc3d, 32'hc2c529f6, 32'hc1634681, 32'hc031e0bf, 32'h4288458f, 32'h420fc540};
test_output[19984:19991] = '{32'h41691d87, 32'h426a41c7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4288458f, 32'h420fc540};
test_input[19992:19999] = '{32'h4215cacc, 32'h4280b042, 32'hc29c6e2a, 32'hc1ba50d1, 32'hc25f1b76, 32'h41971550, 32'h42741cb7, 32'hc2b04893};
test_output[19992:19999] = '{32'h4215cacc, 32'h4280b042, 32'h0, 32'h0, 32'h0, 32'h41971550, 32'h42741cb7, 32'h0};
test_input[20000:20007] = '{32'h42b613c1, 32'hc211fdff, 32'hc2bf0a2a, 32'hc15708c0, 32'hc2c6f77f, 32'h428f9dcb, 32'h42aa4d60, 32'hc242b717};
test_output[20000:20007] = '{32'h42b613c1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428f9dcb, 32'h42aa4d60, 32'h0};
test_input[20008:20015] = '{32'h40fb38e8, 32'hc2b025c5, 32'h42b187d6, 32'hc2a3f42b, 32'hbf04e0c2, 32'h4296813f, 32'h423d7969, 32'h425d3189};
test_output[20008:20015] = '{32'h40fb38e8, 32'h0, 32'h42b187d6, 32'h0, 32'h0, 32'h4296813f, 32'h423d7969, 32'h425d3189};
test_input[20016:20023] = '{32'h42ac876a, 32'hc2732d1b, 32'hc0a1901c, 32'h42ae5ab0, 32'h413fe718, 32'h42c208ed, 32'h425622f3, 32'hc2b605e2};
test_output[20016:20023] = '{32'h42ac876a, 32'h0, 32'h0, 32'h42ae5ab0, 32'h413fe718, 32'h42c208ed, 32'h425622f3, 32'h0};
test_input[20024:20031] = '{32'h411bd45a, 32'h42897f5e, 32'hc297bc35, 32'hc22f501a, 32'h41a87bd6, 32'hc2aa37be, 32'hc1598ffe, 32'h428b5a64};
test_output[20024:20031] = '{32'h411bd45a, 32'h42897f5e, 32'h0, 32'h0, 32'h41a87bd6, 32'h0, 32'h0, 32'h428b5a64};
test_input[20032:20039] = '{32'hc204e3ec, 32'hc2ade922, 32'hc2a5ba11, 32'h427f3ff6, 32'hc24aec69, 32'h42c1a02f, 32'hc2b741e5, 32'h42910c26};
test_output[20032:20039] = '{32'h0, 32'h0, 32'h0, 32'h427f3ff6, 32'h0, 32'h42c1a02f, 32'h0, 32'h42910c26};
test_input[20040:20047] = '{32'h41cedf57, 32'h411eb92d, 32'hc2a02bfe, 32'h428871bc, 32'hc2ae6195, 32'hc070f81e, 32'hc1554039, 32'hc2b781be};
test_output[20040:20047] = '{32'h41cedf57, 32'h411eb92d, 32'h0, 32'h428871bc, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20048:20055] = '{32'hc2c377ed, 32'h4267233e, 32'hc292937e, 32'hc2b8203b, 32'h423307b2, 32'h42002e77, 32'hc25bf82c, 32'hc234ac53};
test_output[20048:20055] = '{32'h0, 32'h4267233e, 32'h0, 32'h0, 32'h423307b2, 32'h42002e77, 32'h0, 32'h0};
test_input[20056:20063] = '{32'h41c40ee9, 32'h4095240d, 32'h42c2c8ef, 32'h41bfa59b, 32'hc2848862, 32'h41d1c4bb, 32'h420f56b2, 32'hc2959a35};
test_output[20056:20063] = '{32'h41c40ee9, 32'h4095240d, 32'h42c2c8ef, 32'h41bfa59b, 32'h0, 32'h41d1c4bb, 32'h420f56b2, 32'h0};
test_input[20064:20071] = '{32'h42a73f06, 32'hc1a0b5c7, 32'h422d4b1b, 32'h42a9ca69, 32'h4287f08e, 32'hc141f165, 32'hc294f0ba, 32'h427ce00c};
test_output[20064:20071] = '{32'h42a73f06, 32'h0, 32'h422d4b1b, 32'h42a9ca69, 32'h4287f08e, 32'h0, 32'h0, 32'h427ce00c};
test_input[20072:20079] = '{32'h415c1736, 32'h420a3334, 32'hc28760cf, 32'hc2b2130b, 32'hc0bc211f, 32'h42c43270, 32'h41bf152f, 32'h409a32ea};
test_output[20072:20079] = '{32'h415c1736, 32'h420a3334, 32'h0, 32'h0, 32'h0, 32'h42c43270, 32'h41bf152f, 32'h409a32ea};
test_input[20080:20087] = '{32'hc24ac08e, 32'hc1624b22, 32'hc044ba6a, 32'hc2c5470f, 32'h420d6604, 32'h429f7e96, 32'hc2465bae, 32'hc2bc01bb};
test_output[20080:20087] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h420d6604, 32'h429f7e96, 32'h0, 32'h0};
test_input[20088:20095] = '{32'h429bb45b, 32'hc21f48e8, 32'h42a91a1a, 32'hc1839439, 32'h4212d4db, 32'hc1de82a2, 32'h426aba00, 32'hc10f983b};
test_output[20088:20095] = '{32'h429bb45b, 32'h0, 32'h42a91a1a, 32'h0, 32'h4212d4db, 32'h0, 32'h426aba00, 32'h0};
test_input[20096:20103] = '{32'hc1f75714, 32'hc2a08b3d, 32'h42612cf9, 32'hc254fef8, 32'hc104590a, 32'h421e1b49, 32'h421a7a14, 32'h42b221c9};
test_output[20096:20103] = '{32'h0, 32'h0, 32'h42612cf9, 32'h0, 32'h0, 32'h421e1b49, 32'h421a7a14, 32'h42b221c9};
test_input[20104:20111] = '{32'h42c6177e, 32'h42c225be, 32'hc1717ecc, 32'h42a8c6bb, 32'hc22b0b03, 32'h425733aa, 32'h42a033f5, 32'hc21442ea};
test_output[20104:20111] = '{32'h42c6177e, 32'h42c225be, 32'h0, 32'h42a8c6bb, 32'h0, 32'h425733aa, 32'h42a033f5, 32'h0};
test_input[20112:20119] = '{32'h4279e65d, 32'hc23350d0, 32'h419ae22a, 32'h423b06ff, 32'hc2b8654d, 32'h42b3e6f5, 32'hc1b1e9a2, 32'h418f075c};
test_output[20112:20119] = '{32'h4279e65d, 32'h0, 32'h419ae22a, 32'h423b06ff, 32'h0, 32'h42b3e6f5, 32'h0, 32'h418f075c};
test_input[20120:20127] = '{32'h4298f419, 32'hc20e4068, 32'hc196aae5, 32'hc21fd852, 32'hc1982541, 32'hc0c73ded, 32'hc237f473, 32'h42172ef6};
test_output[20120:20127] = '{32'h4298f419, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42172ef6};
test_input[20128:20135] = '{32'hc2c5d802, 32'hc20870c0, 32'h42c7c2ae, 32'hc28485a1, 32'h41f92665, 32'hc2553818, 32'hc1542585, 32'hc0988e16};
test_output[20128:20135] = '{32'h0, 32'h0, 32'h42c7c2ae, 32'h0, 32'h41f92665, 32'h0, 32'h0, 32'h0};
test_input[20136:20143] = '{32'hc2931277, 32'hc1c5c51e, 32'hc28856b2, 32'hc2a0f06a, 32'h42a34009, 32'hc187e126, 32'h41ceafb6, 32'h41982d54};
test_output[20136:20143] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a34009, 32'h0, 32'h41ceafb6, 32'h41982d54};
test_input[20144:20151] = '{32'hc15adc53, 32'hc183c166, 32'h4179623b, 32'h4248bd0d, 32'h42c775ec, 32'hc22e00da, 32'h420fcd22, 32'hc2b47140};
test_output[20144:20151] = '{32'h0, 32'h0, 32'h4179623b, 32'h4248bd0d, 32'h42c775ec, 32'h0, 32'h420fcd22, 32'h0};
test_input[20152:20159] = '{32'h4294de57, 32'hc093acc5, 32'h4291f8bb, 32'h41b30576, 32'hc252c65a, 32'h4291af40, 32'h42534277, 32'hc28b80dd};
test_output[20152:20159] = '{32'h4294de57, 32'h0, 32'h4291f8bb, 32'h41b30576, 32'h0, 32'h4291af40, 32'h42534277, 32'h0};
test_input[20160:20167] = '{32'hc2c7171b, 32'h42a2f1a2, 32'hc0ade6e7, 32'hc2c3d844, 32'h42bb3f54, 32'h41f16ac9, 32'h428594c7, 32'hc2c4f9bd};
test_output[20160:20167] = '{32'h0, 32'h42a2f1a2, 32'h0, 32'h0, 32'h42bb3f54, 32'h41f16ac9, 32'h428594c7, 32'h0};
test_input[20168:20175] = '{32'hc1bc6c7d, 32'h420dd68c, 32'hc1c1232e, 32'h4239a3be, 32'hc2bf5c01, 32'h427cd455, 32'h420babe3, 32'hc2871d27};
test_output[20168:20175] = '{32'h0, 32'h420dd68c, 32'h0, 32'h4239a3be, 32'h0, 32'h427cd455, 32'h420babe3, 32'h0};
test_input[20176:20183] = '{32'h4217b1ef, 32'hc25941ae, 32'h414e775c, 32'hc1a78cc2, 32'hc296d0fd, 32'h42a4ab43, 32'h41b10d78, 32'hc2434d07};
test_output[20176:20183] = '{32'h4217b1ef, 32'h0, 32'h414e775c, 32'h0, 32'h0, 32'h42a4ab43, 32'h41b10d78, 32'h0};
test_input[20184:20191] = '{32'hc2c061f1, 32'h42b8b489, 32'hc2b2dcc0, 32'h4278877c, 32'h429c8e91, 32'hc29c2027, 32'hc2974630, 32'h422c7e31};
test_output[20184:20191] = '{32'h0, 32'h42b8b489, 32'h0, 32'h4278877c, 32'h429c8e91, 32'h0, 32'h0, 32'h422c7e31};
test_input[20192:20199] = '{32'h421e2073, 32'h41917f08, 32'h411c702b, 32'hc2385dd5, 32'h41ecfb63, 32'hc289bd5e, 32'h40426599, 32'hc1947ee2};
test_output[20192:20199] = '{32'h421e2073, 32'h41917f08, 32'h411c702b, 32'h0, 32'h41ecfb63, 32'h0, 32'h40426599, 32'h0};
test_input[20200:20207] = '{32'hc26cbfc3, 32'hc1a1c30d, 32'hc20604c2, 32'h42a14bb6, 32'hc26e08ff, 32'hc2404136, 32'hc28e67cc, 32'hc241c472};
test_output[20200:20207] = '{32'h0, 32'h0, 32'h0, 32'h42a14bb6, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20208:20215] = '{32'h4284c906, 32'hc24256b5, 32'hc298372a, 32'h3fa8463b, 32'h42261ab2, 32'hc29836d2, 32'h40ae0077, 32'hc2a370c8};
test_output[20208:20215] = '{32'h4284c906, 32'h0, 32'h0, 32'h3fa8463b, 32'h42261ab2, 32'h0, 32'h40ae0077, 32'h0};
test_input[20216:20223] = '{32'h3f3a5457, 32'h411caa5d, 32'h419bc782, 32'h42236646, 32'hc18d0528, 32'hc1326c64, 32'hc2179579, 32'h4299a0f1};
test_output[20216:20223] = '{32'h3f3a5457, 32'h411caa5d, 32'h419bc782, 32'h42236646, 32'h0, 32'h0, 32'h0, 32'h4299a0f1};
test_input[20224:20231] = '{32'hc086af05, 32'h422ee2ff, 32'h4234f7a6, 32'h40ac5d43, 32'hc28a0691, 32'h4224ea0b, 32'hc2883e4c, 32'hc1148b0c};
test_output[20224:20231] = '{32'h0, 32'h422ee2ff, 32'h4234f7a6, 32'h40ac5d43, 32'h0, 32'h4224ea0b, 32'h0, 32'h0};
test_input[20232:20239] = '{32'h4207a301, 32'hc1ae12dd, 32'h42a06da8, 32'hc288307d, 32'hc1f778e4, 32'h42bcc52c, 32'h4294982e, 32'hc1dde9ab};
test_output[20232:20239] = '{32'h4207a301, 32'h0, 32'h42a06da8, 32'h0, 32'h0, 32'h42bcc52c, 32'h4294982e, 32'h0};
test_input[20240:20247] = '{32'h4292523b, 32'hc204ad34, 32'hc1c0f249, 32'hbf7f0b90, 32'hc2c6e6c1, 32'hc29781e8, 32'h4268d498, 32'hc27aa572};
test_output[20240:20247] = '{32'h4292523b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4268d498, 32'h0};
test_input[20248:20255] = '{32'h417b3d7c, 32'h41e2b10a, 32'hc2953ab7, 32'h41f31dfc, 32'h42a119bb, 32'hc28d770d, 32'hc2334d91, 32'hc2c4ba93};
test_output[20248:20255] = '{32'h417b3d7c, 32'h41e2b10a, 32'h0, 32'h41f31dfc, 32'h42a119bb, 32'h0, 32'h0, 32'h0};
test_input[20256:20263] = '{32'hc18d9a3d, 32'hc2961140, 32'h421fd3f3, 32'h42a4a7fa, 32'h42846b56, 32'h419c8f9c, 32'hbfd75e18, 32'hc2c3e490};
test_output[20256:20263] = '{32'h0, 32'h0, 32'h421fd3f3, 32'h42a4a7fa, 32'h42846b56, 32'h419c8f9c, 32'h0, 32'h0};
test_input[20264:20271] = '{32'hc27eb304, 32'h42117538, 32'hc24ca52d, 32'hc1d3b763, 32'hc2b26048, 32'hbdd31834, 32'hc24bfaf8, 32'hc2913ca7};
test_output[20264:20271] = '{32'h0, 32'h42117538, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20272:20279] = '{32'h423bc923, 32'hc2bded81, 32'h41f01812, 32'hc282d57b, 32'h42839792, 32'hc27eafd5, 32'hc2b39ecb, 32'hc2b861f8};
test_output[20272:20279] = '{32'h423bc923, 32'h0, 32'h41f01812, 32'h0, 32'h42839792, 32'h0, 32'h0, 32'h0};
test_input[20280:20287] = '{32'h42b37516, 32'hc1d780b5, 32'hc122927c, 32'h42aabe43, 32'hc28c8a44, 32'h4231df8c, 32'hc2104391, 32'h42751530};
test_output[20280:20287] = '{32'h42b37516, 32'h0, 32'h0, 32'h42aabe43, 32'h0, 32'h4231df8c, 32'h0, 32'h42751530};
test_input[20288:20295] = '{32'hc0d7e81e, 32'hc2c135b8, 32'h4254bd8f, 32'h416b8425, 32'hc26818a6, 32'h4292718c, 32'h4269161c, 32'h41610a59};
test_output[20288:20295] = '{32'h0, 32'h0, 32'h4254bd8f, 32'h416b8425, 32'h0, 32'h4292718c, 32'h4269161c, 32'h41610a59};
test_input[20296:20303] = '{32'h41f76ef2, 32'hbd9a7deb, 32'hc2956e20, 32'hc2c23ee4, 32'hc222df4a, 32'hc286e229, 32'h410a1b6a, 32'h42692e37};
test_output[20296:20303] = '{32'h41f76ef2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h410a1b6a, 32'h42692e37};
test_input[20304:20311] = '{32'h42bfd47c, 32'hc17ab653, 32'hc245c462, 32'hc28ee540, 32'hc28359e6, 32'hc280bb35, 32'hc2042565, 32'hc2a02c57};
test_output[20304:20311] = '{32'h42bfd47c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20312:20319] = '{32'hc28ca66e, 32'hc16196bb, 32'hc1c715c2, 32'hc2b50bbb, 32'hc2899f17, 32'hc2bd0408, 32'hc208cd94, 32'h42bd7bc2};
test_output[20312:20319] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bd7bc2};
test_input[20320:20327] = '{32'hc2774f3d, 32'h426c83c5, 32'h42187618, 32'h429e3d95, 32'hc158be65, 32'hc2bb113a, 32'hc1983838, 32'hc29a9236};
test_output[20320:20327] = '{32'h0, 32'h426c83c5, 32'h42187618, 32'h429e3d95, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20328:20335] = '{32'h40b1fd35, 32'hc045b9c0, 32'hc16b3b0d, 32'h42c351c6, 32'hc2592698, 32'hc17a31cf, 32'hc2382b1c, 32'h429c9283};
test_output[20328:20335] = '{32'h40b1fd35, 32'h0, 32'h0, 32'h42c351c6, 32'h0, 32'h0, 32'h0, 32'h429c9283};
test_input[20336:20343] = '{32'hc25d8739, 32'h4288c9be, 32'hc182d8d0, 32'h4283be04, 32'hc07791aa, 32'h40a77e77, 32'h429fbf5b, 32'hc20f7642};
test_output[20336:20343] = '{32'h0, 32'h4288c9be, 32'h0, 32'h4283be04, 32'h0, 32'h40a77e77, 32'h429fbf5b, 32'h0};
test_input[20344:20351] = '{32'hc2ab0894, 32'h41bbaabe, 32'h42bccf26, 32'hc2240aca, 32'h420fd55c, 32'hc2bd29a9, 32'hc20eb9b1, 32'hc14f7059};
test_output[20344:20351] = '{32'h0, 32'h41bbaabe, 32'h42bccf26, 32'h0, 32'h420fd55c, 32'h0, 32'h0, 32'h0};
test_input[20352:20359] = '{32'h41fa8c1f, 32'hc03f6dd2, 32'hc203a7c4, 32'h4256fc70, 32'h429ee10c, 32'h423055a0, 32'h41da8d34, 32'hc2b8695a};
test_output[20352:20359] = '{32'h41fa8c1f, 32'h0, 32'h0, 32'h4256fc70, 32'h429ee10c, 32'h423055a0, 32'h41da8d34, 32'h0};
test_input[20360:20367] = '{32'h42b09627, 32'h427cc6ac, 32'h4241b01b, 32'h420e650f, 32'hc2a79893, 32'h42319b33, 32'h42903467, 32'hc12af49e};
test_output[20360:20367] = '{32'h42b09627, 32'h427cc6ac, 32'h4241b01b, 32'h420e650f, 32'h0, 32'h42319b33, 32'h42903467, 32'h0};
test_input[20368:20375] = '{32'hc2a895d7, 32'h41f190e9, 32'hc1641341, 32'hc08db4e4, 32'h42b25539, 32'h421bea37, 32'h41f8a90a, 32'hc20231f3};
test_output[20368:20375] = '{32'h0, 32'h41f190e9, 32'h0, 32'h0, 32'h42b25539, 32'h421bea37, 32'h41f8a90a, 32'h0};
test_input[20376:20383] = '{32'h421e3185, 32'h426e5170, 32'h418d90fa, 32'h42575042, 32'hbeb805ac, 32'h42b78fc3, 32'hc2c63753, 32'hc17c42f8};
test_output[20376:20383] = '{32'h421e3185, 32'h426e5170, 32'h418d90fa, 32'h42575042, 32'h0, 32'h42b78fc3, 32'h0, 32'h0};
test_input[20384:20391] = '{32'h4249ccff, 32'h428bc9a2, 32'hc282fd96, 32'hc2c79232, 32'hc13df8f6, 32'h42a29786, 32'hc24c650c, 32'h42a3b164};
test_output[20384:20391] = '{32'h4249ccff, 32'h428bc9a2, 32'h0, 32'h0, 32'h0, 32'h42a29786, 32'h0, 32'h42a3b164};
test_input[20392:20399] = '{32'hc20a2bbd, 32'hbfc94fbf, 32'hc1fc4a3e, 32'h4270c7ed, 32'h42be3e9c, 32'hc1e23512, 32'hc248f7fb, 32'hc1ba3ac9};
test_output[20392:20399] = '{32'h0, 32'h0, 32'h0, 32'h4270c7ed, 32'h42be3e9c, 32'h0, 32'h0, 32'h0};
test_input[20400:20407] = '{32'hc2bc008f, 32'hc213eaf5, 32'hc1978799, 32'hc22dc110, 32'h42a11431, 32'h422e47b1, 32'hc23c5681, 32'hc2513c16};
test_output[20400:20407] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a11431, 32'h422e47b1, 32'h0, 32'h0};
test_input[20408:20415] = '{32'hc28c1cf6, 32'h426cdd7d, 32'h42b55e4f, 32'hc201bf19, 32'hc2a98d0c, 32'hc1545810, 32'h42bdc788, 32'hc29c227e};
test_output[20408:20415] = '{32'h0, 32'h426cdd7d, 32'h42b55e4f, 32'h0, 32'h0, 32'h0, 32'h42bdc788, 32'h0};
test_input[20416:20423] = '{32'hc2166d5f, 32'hc1c29a23, 32'h40cf9773, 32'hc235214a, 32'h42935df4, 32'hc223567d, 32'hc175bfee, 32'h41e026b6};
test_output[20416:20423] = '{32'h0, 32'h0, 32'h40cf9773, 32'h0, 32'h42935df4, 32'h0, 32'h0, 32'h41e026b6};
test_input[20424:20431] = '{32'h4148207e, 32'hc291a9f6, 32'h41eabd70, 32'h4039b833, 32'hc1e67d08, 32'hc229d136, 32'h408213b1, 32'h4296971e};
test_output[20424:20431] = '{32'h4148207e, 32'h0, 32'h41eabd70, 32'h4039b833, 32'h0, 32'h0, 32'h408213b1, 32'h4296971e};
test_input[20432:20439] = '{32'h41a73561, 32'hc0e45f01, 32'h42117cf0, 32'h41ca7f12, 32'h42aea4c1, 32'h4173470e, 32'h40df51c8, 32'h419a1094};
test_output[20432:20439] = '{32'h41a73561, 32'h0, 32'h42117cf0, 32'h41ca7f12, 32'h42aea4c1, 32'h4173470e, 32'h40df51c8, 32'h419a1094};
test_input[20440:20447] = '{32'hc209bfef, 32'h4237ed68, 32'h427ad1cb, 32'hc0331324, 32'hc2a59c48, 32'hc263cabe, 32'h421d5aa5, 32'hc11b6c6e};
test_output[20440:20447] = '{32'h0, 32'h4237ed68, 32'h427ad1cb, 32'h0, 32'h0, 32'h0, 32'h421d5aa5, 32'h0};
test_input[20448:20455] = '{32'h4120e242, 32'hc25ca589, 32'h429d4bce, 32'hc2a404a8, 32'h4167a542, 32'h426714cd, 32'hc2bef87a, 32'hc29934ea};
test_output[20448:20455] = '{32'h4120e242, 32'h0, 32'h429d4bce, 32'h0, 32'h4167a542, 32'h426714cd, 32'h0, 32'h0};
test_input[20456:20463] = '{32'h420ce5c1, 32'hc29b9fb5, 32'hc2084b5b, 32'h41b519e1, 32'hc20d581c, 32'h42aa499e, 32'hbef9fa79, 32'h4298dfbe};
test_output[20456:20463] = '{32'h420ce5c1, 32'h0, 32'h0, 32'h41b519e1, 32'h0, 32'h42aa499e, 32'h0, 32'h4298dfbe};
test_input[20464:20471] = '{32'h42a38e2b, 32'h42b6fc8c, 32'h427f9018, 32'hc1c2cb2d, 32'hc2b15521, 32'h424363b3, 32'hc1ff6294, 32'h429a5470};
test_output[20464:20471] = '{32'h42a38e2b, 32'h42b6fc8c, 32'h427f9018, 32'h0, 32'h0, 32'h424363b3, 32'h0, 32'h429a5470};
test_input[20472:20479] = '{32'hc1a928d4, 32'h4213627a, 32'hc2b91b48, 32'h421a43e9, 32'h427ec263, 32'hc28f2656, 32'h4298b78b, 32'h42692d9e};
test_output[20472:20479] = '{32'h0, 32'h4213627a, 32'h0, 32'h421a43e9, 32'h427ec263, 32'h0, 32'h4298b78b, 32'h42692d9e};
test_input[20480:20487] = '{32'hc1a839b0, 32'h41d1dc32, 32'hc1b331e1, 32'hc1393f81, 32'hc11d84dc, 32'hc1eb5aff, 32'hc26bb733, 32'h41afc6e1};
test_output[20480:20487] = '{32'h0, 32'h41d1dc32, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41afc6e1};
test_input[20488:20495] = '{32'hc18426b3, 32'hc1b14036, 32'hc2b46bc7, 32'hc1d50b8c, 32'hc2147602, 32'h42892528, 32'h42a618a9, 32'hc21259b8};
test_output[20488:20495] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42892528, 32'h42a618a9, 32'h0};
test_input[20496:20503] = '{32'hc20e490d, 32'hc28cb704, 32'h427704e0, 32'h42679e29, 32'hc2022d83, 32'h4250639e, 32'h42949aca, 32'h425854be};
test_output[20496:20503] = '{32'h0, 32'h0, 32'h427704e0, 32'h42679e29, 32'h0, 32'h4250639e, 32'h42949aca, 32'h425854be};
test_input[20504:20511] = '{32'hc2a9b4a3, 32'h4142de81, 32'hc257fe3f, 32'h42927268, 32'hc2ac6048, 32'hc22515e0, 32'hc2a44592, 32'h40f1f54a};
test_output[20504:20511] = '{32'h0, 32'h4142de81, 32'h0, 32'h42927268, 32'h0, 32'h0, 32'h0, 32'h40f1f54a};
test_input[20512:20519] = '{32'hc27ebbc5, 32'h42a226f7, 32'hc1b09118, 32'hc2abc061, 32'hc24ddeb6, 32'hc2c4f53a, 32'h4207ca99, 32'h40e7ea43};
test_output[20512:20519] = '{32'h0, 32'h42a226f7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4207ca99, 32'h40e7ea43};
test_input[20520:20527] = '{32'hc24423f4, 32'h424d9a5b, 32'h428e4224, 32'h42bf3b43, 32'hc1de6a7a, 32'hc2678a75, 32'h429e89e3, 32'hc18d3ee4};
test_output[20520:20527] = '{32'h0, 32'h424d9a5b, 32'h428e4224, 32'h42bf3b43, 32'h0, 32'h0, 32'h429e89e3, 32'h0};
test_input[20528:20535] = '{32'h42887e1d, 32'h41ae5660, 32'hc293574a, 32'h427afeb4, 32'hc2ba72db, 32'h426765c3, 32'hc0956066, 32'h4270591a};
test_output[20528:20535] = '{32'h42887e1d, 32'h41ae5660, 32'h0, 32'h427afeb4, 32'h0, 32'h426765c3, 32'h0, 32'h4270591a};
test_input[20536:20543] = '{32'h423e085f, 32'h42ab1082, 32'h41e88c57, 32'hc28ffd35, 32'h42a7fa5b, 32'h424380d3, 32'h42ba24b7, 32'h41ef4c4e};
test_output[20536:20543] = '{32'h423e085f, 32'h42ab1082, 32'h41e88c57, 32'h0, 32'h42a7fa5b, 32'h424380d3, 32'h42ba24b7, 32'h41ef4c4e};
test_input[20544:20551] = '{32'hc2290593, 32'h42b1cdc2, 32'h42ab1f85, 32'hc1347ebb, 32'hc21637b8, 32'hc27f7571, 32'hc1df486a, 32'h42b41dc0};
test_output[20544:20551] = '{32'h0, 32'h42b1cdc2, 32'h42ab1f85, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b41dc0};
test_input[20552:20559] = '{32'hc28148bd, 32'hc084dcec, 32'hc24276f1, 32'hc1a25238, 32'hc299d608, 32'hc283e9d3, 32'hc1bbd4aa, 32'hc21d5404};
test_output[20552:20559] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20560:20567] = '{32'hc293d379, 32'hc0a866e3, 32'hc1bd0eeb, 32'h42a2a59b, 32'hc243369a, 32'h42aab378, 32'h42b45b20, 32'hc1ce5488};
test_output[20560:20567] = '{32'h0, 32'h0, 32'h0, 32'h42a2a59b, 32'h0, 32'h42aab378, 32'h42b45b20, 32'h0};
test_input[20568:20575] = '{32'hc254969f, 32'hc2b9b935, 32'hc24dc5ba, 32'hc29094b5, 32'hc2a67a67, 32'h4033aba5, 32'h42930ebe, 32'h42b3efe6};
test_output[20568:20575] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4033aba5, 32'h42930ebe, 32'h42b3efe6};
test_input[20576:20583] = '{32'h4234b511, 32'hc2938b05, 32'h3f4e1a55, 32'hc2745f70, 32'hc113d441, 32'h4267c7a1, 32'hbf50e5f6, 32'h42a06318};
test_output[20576:20583] = '{32'h4234b511, 32'h0, 32'h3f4e1a55, 32'h0, 32'h0, 32'h4267c7a1, 32'h0, 32'h42a06318};
test_input[20584:20591] = '{32'h40eaebfb, 32'hc1c5123f, 32'h428de9c7, 32'hc2bec719, 32'h42a24369, 32'h42a0dd3a, 32'hc21a53db, 32'h426b6a99};
test_output[20584:20591] = '{32'h40eaebfb, 32'h0, 32'h428de9c7, 32'h0, 32'h42a24369, 32'h42a0dd3a, 32'h0, 32'h426b6a99};
test_input[20592:20599] = '{32'hc1c192d8, 32'h422de148, 32'hc2a630c8, 32'hc2963c5f, 32'h42230456, 32'hc24cb7b5, 32'h42bfa7fd, 32'h42ba17d3};
test_output[20592:20599] = '{32'h0, 32'h422de148, 32'h0, 32'h0, 32'h42230456, 32'h0, 32'h42bfa7fd, 32'h42ba17d3};
test_input[20600:20607] = '{32'h4215cd37, 32'h427e0fd7, 32'h4292824b, 32'h429f7ff4, 32'h41ac14d8, 32'h42c151b7, 32'h420676a3, 32'hbfaa50a2};
test_output[20600:20607] = '{32'h4215cd37, 32'h427e0fd7, 32'h4292824b, 32'h429f7ff4, 32'h41ac14d8, 32'h42c151b7, 32'h420676a3, 32'h0};
test_input[20608:20615] = '{32'h4203c64f, 32'hc18a5030, 32'h41c7eccc, 32'h4213a13b, 32'hc1a286b8, 32'h42b7fbce, 32'h41e0c39b, 32'h42a2c8ce};
test_output[20608:20615] = '{32'h4203c64f, 32'h0, 32'h41c7eccc, 32'h4213a13b, 32'h0, 32'h42b7fbce, 32'h41e0c39b, 32'h42a2c8ce};
test_input[20616:20623] = '{32'hc2afc7ac, 32'h429edce1, 32'h41000e42, 32'h41732ffd, 32'hc16f5894, 32'hbf82d932, 32'hc2a015fb, 32'h426e3572};
test_output[20616:20623] = '{32'h0, 32'h429edce1, 32'h41000e42, 32'h41732ffd, 32'h0, 32'h0, 32'h0, 32'h426e3572};
test_input[20624:20631] = '{32'h422f22fe, 32'h41a3f587, 32'h424b9130, 32'h41e8664d, 32'h4268a43d, 32'h42252933, 32'hc23ad746, 32'h42898848};
test_output[20624:20631] = '{32'h422f22fe, 32'h41a3f587, 32'h424b9130, 32'h41e8664d, 32'h4268a43d, 32'h42252933, 32'h0, 32'h42898848};
test_input[20632:20639] = '{32'h428a39e4, 32'h4256768c, 32'hc201dadb, 32'h40f8b563, 32'hc15958e8, 32'hc238a9ce, 32'h3f945f25, 32'hc2b2c080};
test_output[20632:20639] = '{32'h428a39e4, 32'h4256768c, 32'h0, 32'h40f8b563, 32'h0, 32'h0, 32'h3f945f25, 32'h0};
test_input[20640:20647] = '{32'h427352cd, 32'h42515561, 32'hc292c40f, 32'hc18a5aa0, 32'h4249a3da, 32'h40a0fbc8, 32'h42b18a51, 32'hc262118b};
test_output[20640:20647] = '{32'h427352cd, 32'h42515561, 32'h0, 32'h0, 32'h4249a3da, 32'h40a0fbc8, 32'h42b18a51, 32'h0};
test_input[20648:20655] = '{32'h42866b5b, 32'hc2850f5a, 32'h4191fe64, 32'h429c4bc9, 32'h4258fb50, 32'h4268e995, 32'h42409415, 32'h3f00dd84};
test_output[20648:20655] = '{32'h42866b5b, 32'h0, 32'h4191fe64, 32'h429c4bc9, 32'h4258fb50, 32'h4268e995, 32'h42409415, 32'h3f00dd84};
test_input[20656:20663] = '{32'h41d762c6, 32'h41d9a967, 32'hc275e821, 32'h41ae0888, 32'h4294624d, 32'hc1f9e1bd, 32'hc1dad8b2, 32'h4120801d};
test_output[20656:20663] = '{32'h41d762c6, 32'h41d9a967, 32'h0, 32'h41ae0888, 32'h4294624d, 32'h0, 32'h0, 32'h4120801d};
test_input[20664:20671] = '{32'hc18ed0dd, 32'h4059a4b6, 32'h428a5fc4, 32'hc2b3c8ee, 32'h428d45af, 32'hc282d1ff, 32'h42b1da9f, 32'h4285e263};
test_output[20664:20671] = '{32'h0, 32'h4059a4b6, 32'h428a5fc4, 32'h0, 32'h428d45af, 32'h0, 32'h42b1da9f, 32'h4285e263};
test_input[20672:20679] = '{32'h412fabfd, 32'h427738a0, 32'h4283c57b, 32'h41826b43, 32'hc18076ef, 32'hc226598d, 32'h41d7084b, 32'h426c52e6};
test_output[20672:20679] = '{32'h412fabfd, 32'h427738a0, 32'h4283c57b, 32'h41826b43, 32'h0, 32'h0, 32'h41d7084b, 32'h426c52e6};
test_input[20680:20687] = '{32'h41bcaf10, 32'h423110cd, 32'h42808985, 32'h41df2b3f, 32'hc1cfdf5e, 32'hc263797d, 32'h4298b350, 32'h3fae5830};
test_output[20680:20687] = '{32'h41bcaf10, 32'h423110cd, 32'h42808985, 32'h41df2b3f, 32'h0, 32'h0, 32'h4298b350, 32'h3fae5830};
test_input[20688:20695] = '{32'hc2b2d389, 32'h4291093c, 32'hc2917c62, 32'hc227836f, 32'hc1b84317, 32'hc193440f, 32'hc2b698f4, 32'h42a775dc};
test_output[20688:20695] = '{32'h0, 32'h4291093c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a775dc};
test_input[20696:20703] = '{32'hc2a231ef, 32'hc2865ea9, 32'h42b1300f, 32'hc1aa6a60, 32'h42a983f4, 32'h420e499c, 32'hc16e77a4, 32'h429a3bc2};
test_output[20696:20703] = '{32'h0, 32'h0, 32'h42b1300f, 32'h0, 32'h42a983f4, 32'h420e499c, 32'h0, 32'h429a3bc2};
test_input[20704:20711] = '{32'h424edd60, 32'h423ca43d, 32'h4225090c, 32'h42376f67, 32'h41d975d5, 32'h42bfcc53, 32'h40804ec4, 32'h410d4a1b};
test_output[20704:20711] = '{32'h424edd60, 32'h423ca43d, 32'h4225090c, 32'h42376f67, 32'h41d975d5, 32'h42bfcc53, 32'h40804ec4, 32'h410d4a1b};
test_input[20712:20719] = '{32'hc1eb6342, 32'h3f32e6ca, 32'hc24976c7, 32'h411f8e21, 32'hc28511c1, 32'h4124b398, 32'h42c5636e, 32'h42a5820b};
test_output[20712:20719] = '{32'h0, 32'h3f32e6ca, 32'h0, 32'h411f8e21, 32'h0, 32'h4124b398, 32'h42c5636e, 32'h42a5820b};
test_input[20720:20727] = '{32'h426b6b65, 32'hc289b896, 32'h424d4f7a, 32'hc2bbd2b7, 32'hc2a234e2, 32'hc172aef7, 32'hc1735ef5, 32'h42c7f6ed};
test_output[20720:20727] = '{32'h426b6b65, 32'h0, 32'h424d4f7a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c7f6ed};
test_input[20728:20735] = '{32'h411307f6, 32'h410d1fa1, 32'h42c7eedb, 32'hc18bfb00, 32'h3dcdb46e, 32'h42a8176c, 32'h42bff763, 32'h42866f11};
test_output[20728:20735] = '{32'h411307f6, 32'h410d1fa1, 32'h42c7eedb, 32'h0, 32'h3dcdb46e, 32'h42a8176c, 32'h42bff763, 32'h42866f11};
test_input[20736:20743] = '{32'hc2b9bdcd, 32'hbfbb3aa6, 32'hc1aca430, 32'h422c5775, 32'hc2b2da63, 32'h42c147bb, 32'h428998bc, 32'hc25714ad};
test_output[20736:20743] = '{32'h0, 32'h0, 32'h0, 32'h422c5775, 32'h0, 32'h42c147bb, 32'h428998bc, 32'h0};
test_input[20744:20751] = '{32'h429c00b7, 32'hc28ae6ce, 32'h4174a785, 32'h425cc7d6, 32'hc29eef85, 32'hc236e157, 32'h4278010e, 32'h4223f51e};
test_output[20744:20751] = '{32'h429c00b7, 32'h0, 32'h4174a785, 32'h425cc7d6, 32'h0, 32'h0, 32'h4278010e, 32'h4223f51e};
test_input[20752:20759] = '{32'hc1f97aad, 32'h42bdd1e1, 32'h4279d7c0, 32'hc210713f, 32'h4286d4d7, 32'h41947af5, 32'hc29bb6c4, 32'hc287964c};
test_output[20752:20759] = '{32'h0, 32'h42bdd1e1, 32'h4279d7c0, 32'h0, 32'h4286d4d7, 32'h41947af5, 32'h0, 32'h0};
test_input[20760:20767] = '{32'hc0d6893d, 32'hc2051a74, 32'h428f2f00, 32'h41925557, 32'h42a3191b, 32'hc2917e8f, 32'h4268106b, 32'hc216d548};
test_output[20760:20767] = '{32'h0, 32'h0, 32'h428f2f00, 32'h41925557, 32'h42a3191b, 32'h0, 32'h4268106b, 32'h0};
test_input[20768:20775] = '{32'hc26391d1, 32'hc1fce2dc, 32'hc1bf056a, 32'h41cc0ecb, 32'h428f5167, 32'hc291d0b2, 32'hc20f3f43, 32'h41f29cf5};
test_output[20768:20775] = '{32'h0, 32'h0, 32'h0, 32'h41cc0ecb, 32'h428f5167, 32'h0, 32'h0, 32'h41f29cf5};
test_input[20776:20783] = '{32'hc1ad49aa, 32'h42c3f478, 32'h422d7061, 32'h428dbf55, 32'h421eea75, 32'hc24ad053, 32'h42800fad, 32'hc23a7159};
test_output[20776:20783] = '{32'h0, 32'h42c3f478, 32'h422d7061, 32'h428dbf55, 32'h421eea75, 32'h0, 32'h42800fad, 32'h0};
test_input[20784:20791] = '{32'h42acb0ae, 32'hc2bf2e54, 32'hbf44da8f, 32'hc13bbb18, 32'h424f1222, 32'h428bcd48, 32'h42728388, 32'h42887b81};
test_output[20784:20791] = '{32'h42acb0ae, 32'h0, 32'h0, 32'h0, 32'h424f1222, 32'h428bcd48, 32'h42728388, 32'h42887b81};
test_input[20792:20799] = '{32'h42bc2dd0, 32'hc2be44b5, 32'hc27ef54b, 32'hc2391f76, 32'h42c191b3, 32'hc1d5a36b, 32'h42a782d8, 32'h42447498};
test_output[20792:20799] = '{32'h42bc2dd0, 32'h0, 32'h0, 32'h0, 32'h42c191b3, 32'h0, 32'h42a782d8, 32'h42447498};
test_input[20800:20807] = '{32'h4165e7ef, 32'hc2027490, 32'hc18574f4, 32'hc2bc631f, 32'hc1302848, 32'h42715d30, 32'h422315ec, 32'h422b383b};
test_output[20800:20807] = '{32'h4165e7ef, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42715d30, 32'h422315ec, 32'h422b383b};
test_input[20808:20815] = '{32'hc203e0b8, 32'hc2673999, 32'h42851510, 32'h425e08e1, 32'hc2795c49, 32'hc1b786fb, 32'hc2a99dc3, 32'h3f03bbf1};
test_output[20808:20815] = '{32'h0, 32'h0, 32'h42851510, 32'h425e08e1, 32'h0, 32'h0, 32'h0, 32'h3f03bbf1};
test_input[20816:20823] = '{32'h42922954, 32'hc215d0be, 32'hc2bbb0be, 32'hc13f4431, 32'h423d2eaa, 32'h41d61606, 32'h42a2e98f, 32'h41e6fc3a};
test_output[20816:20823] = '{32'h42922954, 32'h0, 32'h0, 32'h0, 32'h423d2eaa, 32'h41d61606, 32'h42a2e98f, 32'h41e6fc3a};
test_input[20824:20831] = '{32'h42a93065, 32'h423de387, 32'h42a00e5b, 32'h3f89b0fe, 32'hc2a06937, 32'hc1f02646, 32'hc23865d0, 32'hc046007d};
test_output[20824:20831] = '{32'h42a93065, 32'h423de387, 32'h42a00e5b, 32'h3f89b0fe, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20832:20839] = '{32'hbf8eae13, 32'h42c136cc, 32'h4236834e, 32'h40b38308, 32'hc1bcac9e, 32'h428a6af3, 32'hc18020ca, 32'hc0cf70e4};
test_output[20832:20839] = '{32'h0, 32'h42c136cc, 32'h4236834e, 32'h40b38308, 32'h0, 32'h428a6af3, 32'h0, 32'h0};
test_input[20840:20847] = '{32'hc2918941, 32'hc08e66a3, 32'hc1073754, 32'h41a329d7, 32'hc28a22bb, 32'hc20d3a13, 32'hc2952868, 32'hc207a64d};
test_output[20840:20847] = '{32'h0, 32'h0, 32'h0, 32'h41a329d7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[20848:20855] = '{32'h40c77866, 32'hc2a55e0c, 32'hc2c5d5c8, 32'hc25885b3, 32'hc13767f5, 32'h3f54e90a, 32'h41ec889b, 32'h41ed67d9};
test_output[20848:20855] = '{32'h40c77866, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3f54e90a, 32'h41ec889b, 32'h41ed67d9};
test_input[20856:20863] = '{32'h42c31da9, 32'h41187c28, 32'h4181d36f, 32'h4205d60d, 32'h401ffc2e, 32'h424d6094, 32'hc23e337a, 32'h423bc4db};
test_output[20856:20863] = '{32'h42c31da9, 32'h41187c28, 32'h4181d36f, 32'h4205d60d, 32'h401ffc2e, 32'h424d6094, 32'h0, 32'h423bc4db};
test_input[20864:20871] = '{32'h419fdd9a, 32'h4281b81d, 32'hc237ad44, 32'h42c1a7c2, 32'hc2a76c9b, 32'h42a9ca90, 32'h4158ac42, 32'hc1772bd2};
test_output[20864:20871] = '{32'h419fdd9a, 32'h4281b81d, 32'h0, 32'h42c1a7c2, 32'h0, 32'h42a9ca90, 32'h4158ac42, 32'h0};
test_input[20872:20879] = '{32'hc23263d7, 32'h4027935d, 32'h409ed89f, 32'h41946460, 32'h41f6cf62, 32'hc27873bd, 32'hc1f87428, 32'hc2c0a92d};
test_output[20872:20879] = '{32'h0, 32'h4027935d, 32'h409ed89f, 32'h41946460, 32'h41f6cf62, 32'h0, 32'h0, 32'h0};
test_input[20880:20887] = '{32'hbfeafdd7, 32'hc19c2c3b, 32'h42790467, 32'hc14ab0f2, 32'hc252e611, 32'h3fd080ed, 32'h41483efc, 32'hc2a8a0b6};
test_output[20880:20887] = '{32'h0, 32'h0, 32'h42790467, 32'h0, 32'h0, 32'h3fd080ed, 32'h41483efc, 32'h0};
test_input[20888:20895] = '{32'hc1e6d1b2, 32'hc2ba14a9, 32'hc20f9839, 32'h42839eb3, 32'hc28e201a, 32'h4207e180, 32'hc122ba03, 32'h42b2f439};
test_output[20888:20895] = '{32'h0, 32'h0, 32'h0, 32'h42839eb3, 32'h0, 32'h4207e180, 32'h0, 32'h42b2f439};
test_input[20896:20903] = '{32'h4262fd75, 32'hc2ab6887, 32'h4197c0f3, 32'hc25b6471, 32'h42800852, 32'h4174edc8, 32'h421e2aae, 32'h41b0e3ef};
test_output[20896:20903] = '{32'h4262fd75, 32'h0, 32'h4197c0f3, 32'h0, 32'h42800852, 32'h4174edc8, 32'h421e2aae, 32'h41b0e3ef};
test_input[20904:20911] = '{32'hc255a27c, 32'hc26eace2, 32'h4171cfd4, 32'h4170235c, 32'h422ecd10, 32'hc0e6e7b1, 32'hc255a7f9, 32'hc1fc6556};
test_output[20904:20911] = '{32'h0, 32'h0, 32'h4171cfd4, 32'h4170235c, 32'h422ecd10, 32'h0, 32'h0, 32'h0};
test_input[20912:20919] = '{32'hc2b686dd, 32'h428d7b30, 32'hc29bcc00, 32'h42831f5d, 32'h42917a0f, 32'h424d2fbf, 32'hc2a774d4, 32'h41c52451};
test_output[20912:20919] = '{32'h0, 32'h428d7b30, 32'h0, 32'h42831f5d, 32'h42917a0f, 32'h424d2fbf, 32'h0, 32'h41c52451};
test_input[20920:20927] = '{32'h40e62fcc, 32'hc2b8d1bb, 32'hc1b5914a, 32'h420e873b, 32'h42b39274, 32'hc22992a1, 32'h4156e45b, 32'hc2485104};
test_output[20920:20927] = '{32'h40e62fcc, 32'h0, 32'h0, 32'h420e873b, 32'h42b39274, 32'h0, 32'h4156e45b, 32'h0};
test_input[20928:20935] = '{32'h428a639b, 32'hc26431f3, 32'hc0231189, 32'h40e8d1f6, 32'h4201d46f, 32'hc21b7f44, 32'h4295f26c, 32'hc28434b7};
test_output[20928:20935] = '{32'h428a639b, 32'h0, 32'h0, 32'h40e8d1f6, 32'h4201d46f, 32'h0, 32'h4295f26c, 32'h0};
test_input[20936:20943] = '{32'hc276b872, 32'h41d5d311, 32'h4298e574, 32'h4171e783, 32'h41d3366c, 32'hc1afcc49, 32'hbfbe45ed, 32'hc280d2fb};
test_output[20936:20943] = '{32'h0, 32'h41d5d311, 32'h4298e574, 32'h4171e783, 32'h41d3366c, 32'h0, 32'h0, 32'h0};
test_input[20944:20951] = '{32'h4190727e, 32'h421115ec, 32'hc14fe942, 32'hc2748dad, 32'hc1262a1b, 32'hc2a45fc5, 32'hc255ba8b, 32'h4269e404};
test_output[20944:20951] = '{32'h4190727e, 32'h421115ec, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4269e404};
test_input[20952:20959] = '{32'hc2532919, 32'hc2943882, 32'hc25e1377, 32'h41400925, 32'h405b6ec6, 32'hbfa85719, 32'hc2b8e9c2, 32'h4258c5af};
test_output[20952:20959] = '{32'h0, 32'h0, 32'h0, 32'h41400925, 32'h405b6ec6, 32'h0, 32'h0, 32'h4258c5af};
test_input[20960:20967] = '{32'hc2318a1c, 32'hc19529a8, 32'hc21df1e9, 32'hc1a95c7c, 32'hc29f1f8d, 32'h42acdab4, 32'h40c9b0c7, 32'h42a485ee};
test_output[20960:20967] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42acdab4, 32'h40c9b0c7, 32'h42a485ee};
test_input[20968:20975] = '{32'hc1de0d0a, 32'h426be555, 32'hc2b8edd9, 32'hc1d4e2b1, 32'hc2af93cc, 32'hc12f9f20, 32'h42b11cd8, 32'hc1f5779e};
test_output[20968:20975] = '{32'h0, 32'h426be555, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b11cd8, 32'h0};
test_input[20976:20983] = '{32'hc1a62c2d, 32'hc20721dd, 32'hc27819a6, 32'h42a2f6c4, 32'h42a11988, 32'hc21352c0, 32'h4159e6d7, 32'hc2c44fd1};
test_output[20976:20983] = '{32'h0, 32'h0, 32'h0, 32'h42a2f6c4, 32'h42a11988, 32'h0, 32'h4159e6d7, 32'h0};
test_input[20984:20991] = '{32'hc24949b8, 32'h42b1e1ee, 32'hc2c42ea5, 32'hc26c8b9f, 32'h429b0b02, 32'hbf86224f, 32'hc278d492, 32'h41cbd926};
test_output[20984:20991] = '{32'h0, 32'h42b1e1ee, 32'h0, 32'h0, 32'h429b0b02, 32'h0, 32'h0, 32'h41cbd926};
test_input[20992:20999] = '{32'hc2062aa5, 32'h42894f8d, 32'h4213c79c, 32'hc2bbf668, 32'hc0f1d389, 32'h418d51af, 32'h42070a1e, 32'h423570e7};
test_output[20992:20999] = '{32'h0, 32'h42894f8d, 32'h4213c79c, 32'h0, 32'h0, 32'h418d51af, 32'h42070a1e, 32'h423570e7};
test_input[21000:21007] = '{32'hc2c36988, 32'hc27addc8, 32'hc2608210, 32'h4150ba6a, 32'hc22686f9, 32'hc2173fce, 32'hc2184b99, 32'hc20ca331};
test_output[21000:21007] = '{32'h0, 32'h0, 32'h0, 32'h4150ba6a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21008:21015] = '{32'h42aaacef, 32'hc2ab04ab, 32'hc2823c93, 32'h41f0fc7c, 32'hc1cd41ce, 32'h427e4cde, 32'hc1dd2f39, 32'h42651e92};
test_output[21008:21015] = '{32'h42aaacef, 32'h0, 32'h0, 32'h41f0fc7c, 32'h0, 32'h427e4cde, 32'h0, 32'h42651e92};
test_input[21016:21023] = '{32'h428b4d6c, 32'h4201abce, 32'h4270478f, 32'hc2b8c5b1, 32'hc146751a, 32'h41428f1d, 32'h4237fea5, 32'h42891488};
test_output[21016:21023] = '{32'h428b4d6c, 32'h4201abce, 32'h4270478f, 32'h0, 32'h0, 32'h41428f1d, 32'h4237fea5, 32'h42891488};
test_input[21024:21031] = '{32'hc236669e, 32'hc17207b2, 32'h427791e5, 32'h4261d68d, 32'h42689aa9, 32'h429b62bd, 32'hc2a11c8b, 32'hc0a5561b};
test_output[21024:21031] = '{32'h0, 32'h0, 32'h427791e5, 32'h4261d68d, 32'h42689aa9, 32'h429b62bd, 32'h0, 32'h0};
test_input[21032:21039] = '{32'hc284dfd9, 32'hc29a3e38, 32'hbfbbbd8b, 32'hc0d9a839, 32'hc1fa34e1, 32'hc2906071, 32'hc2692381, 32'hc088314b};
test_output[21032:21039] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21040:21047] = '{32'h41070d00, 32'h3fc24098, 32'hc29e79ba, 32'h422e73de, 32'h42acfca8, 32'hc24b7ef3, 32'hc264b9cc, 32'h40c09e26};
test_output[21040:21047] = '{32'h41070d00, 32'h3fc24098, 32'h0, 32'h422e73de, 32'h42acfca8, 32'h0, 32'h0, 32'h40c09e26};
test_input[21048:21055] = '{32'hc128d170, 32'h41a4be7d, 32'h427d8056, 32'hc287d7a6, 32'h42349d17, 32'h41629532, 32'hc2ada4c6, 32'h429cae3b};
test_output[21048:21055] = '{32'h0, 32'h41a4be7d, 32'h427d8056, 32'h0, 32'h42349d17, 32'h41629532, 32'h0, 32'h429cae3b};
test_input[21056:21063] = '{32'hc2b04a85, 32'hc2652763, 32'h42c41317, 32'hc2a731e0, 32'hc12292ab, 32'h4230a547, 32'h427cc1fd, 32'hc2aef287};
test_output[21056:21063] = '{32'h0, 32'h0, 32'h42c41317, 32'h0, 32'h0, 32'h4230a547, 32'h427cc1fd, 32'h0};
test_input[21064:21071] = '{32'hc20bebc0, 32'h420b4a8e, 32'hc1e4e8d1, 32'hc217f017, 32'h41916edb, 32'hc29eebe2, 32'hc2c6a601, 32'hc2b46ac8};
test_output[21064:21071] = '{32'h0, 32'h420b4a8e, 32'h0, 32'h0, 32'h41916edb, 32'h0, 32'h0, 32'h0};
test_input[21072:21079] = '{32'h42849b79, 32'h40c82c3e, 32'hc1fef7a3, 32'hc2bdd866, 32'h410c6c03, 32'h428281d2, 32'h429776d0, 32'h420aef2c};
test_output[21072:21079] = '{32'h42849b79, 32'h40c82c3e, 32'h0, 32'h0, 32'h410c6c03, 32'h428281d2, 32'h429776d0, 32'h420aef2c};
test_input[21080:21087] = '{32'hc27afdc6, 32'h4040b1d5, 32'hc1d82e6d, 32'hc2385f3f, 32'h42893e1b, 32'hc2bb9437, 32'hc2984b55, 32'hc2c4157c};
test_output[21080:21087] = '{32'h0, 32'h4040b1d5, 32'h0, 32'h0, 32'h42893e1b, 32'h0, 32'h0, 32'h0};
test_input[21088:21095] = '{32'hc2811eac, 32'hc1b765cb, 32'hc29c8b76, 32'h427cdfae, 32'h4201521c, 32'h40a50ad5, 32'h4245d42f, 32'h42c08cad};
test_output[21088:21095] = '{32'h0, 32'h0, 32'h0, 32'h427cdfae, 32'h4201521c, 32'h40a50ad5, 32'h4245d42f, 32'h42c08cad};
test_input[21096:21103] = '{32'h42916f12, 32'hc290c0fa, 32'h3faa252e, 32'h42828c52, 32'h422a7640, 32'h42ae331c, 32'h41bbde33, 32'hc231fe04};
test_output[21096:21103] = '{32'h42916f12, 32'h0, 32'h3faa252e, 32'h42828c52, 32'h422a7640, 32'h42ae331c, 32'h41bbde33, 32'h0};
test_input[21104:21111] = '{32'h40d45b85, 32'h4296ee1a, 32'hc22880f0, 32'hc229266c, 32'hc122590d, 32'hc2295121, 32'h42b1bb8e, 32'h42a0a065};
test_output[21104:21111] = '{32'h40d45b85, 32'h4296ee1a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b1bb8e, 32'h42a0a065};
test_input[21112:21119] = '{32'hc2a33faa, 32'h428c63ab, 32'hbeba759d, 32'hc28b3f5d, 32'h42825fd5, 32'hc247a5b0, 32'h42171816, 32'hc298039c};
test_output[21112:21119] = '{32'h0, 32'h428c63ab, 32'h0, 32'h0, 32'h42825fd5, 32'h0, 32'h42171816, 32'h0};
test_input[21120:21127] = '{32'hc2501829, 32'h429d38ff, 32'h41c2662f, 32'hc29512e0, 32'hc18e41d7, 32'hc1f5c298, 32'hc2b7b920, 32'h42a17f23};
test_output[21120:21127] = '{32'h0, 32'h429d38ff, 32'h41c2662f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a17f23};
test_input[21128:21135] = '{32'hc2a48a52, 32'hc2638ea0, 32'h423d8b00, 32'hc0918515, 32'h4291598e, 32'hc2b87d42, 32'hc29c0b9c, 32'h42a5193c};
test_output[21128:21135] = '{32'h0, 32'h0, 32'h423d8b00, 32'h0, 32'h4291598e, 32'h0, 32'h0, 32'h42a5193c};
test_input[21136:21143] = '{32'h4213624b, 32'h41a25c58, 32'hc2aeac40, 32'hc19c1065, 32'hc2474239, 32'hc284a00e, 32'hc2320b66, 32'h42328097};
test_output[21136:21143] = '{32'h4213624b, 32'h41a25c58, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42328097};
test_input[21144:21151] = '{32'h4232d64b, 32'h429cd44b, 32'h3e6ecc33, 32'h42798b92, 32'h429dc1f8, 32'hc256299a, 32'hc2a51e51, 32'hc2c40776};
test_output[21144:21151] = '{32'h4232d64b, 32'h429cd44b, 32'h3e6ecc33, 32'h42798b92, 32'h429dc1f8, 32'h0, 32'h0, 32'h0};
test_input[21152:21159] = '{32'h4110ae98, 32'hc2531803, 32'h42551abb, 32'hc2c20d98, 32'h4152bf9c, 32'hc187bf09, 32'hc2a6970c, 32'hc2524652};
test_output[21152:21159] = '{32'h4110ae98, 32'h0, 32'h42551abb, 32'h0, 32'h4152bf9c, 32'h0, 32'h0, 32'h0};
test_input[21160:21167] = '{32'hc223f26e, 32'hc2b40041, 32'hc2be39ef, 32'hc289b57e, 32'h42aa7bfd, 32'h4230e750, 32'h42bed01f, 32'hc298d347};
test_output[21160:21167] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42aa7bfd, 32'h4230e750, 32'h42bed01f, 32'h0};
test_input[21168:21175] = '{32'h41775c1c, 32'h4270aaba, 32'h4087c6f5, 32'hc299d484, 32'h4252bd72, 32'hc1016bbc, 32'h429bf2bf, 32'h42464aa3};
test_output[21168:21175] = '{32'h41775c1c, 32'h4270aaba, 32'h4087c6f5, 32'h0, 32'h4252bd72, 32'h0, 32'h429bf2bf, 32'h42464aa3};
test_input[21176:21183] = '{32'h4263855d, 32'h4268a824, 32'h4293dcc8, 32'hc222bd59, 32'hc2ae7d82, 32'hc0836362, 32'h42594e84, 32'h42a21bd1};
test_output[21176:21183] = '{32'h4263855d, 32'h4268a824, 32'h4293dcc8, 32'h0, 32'h0, 32'h0, 32'h42594e84, 32'h42a21bd1};
test_input[21184:21191] = '{32'hc225144d, 32'h42b44ce7, 32'hc17905e9, 32'h41481713, 32'hc25d89a5, 32'hc2a5a098, 32'hc0e3baa6, 32'h41c79ee7};
test_output[21184:21191] = '{32'h0, 32'h42b44ce7, 32'h0, 32'h41481713, 32'h0, 32'h0, 32'h0, 32'h41c79ee7};
test_input[21192:21199] = '{32'hbfd1592b, 32'hc2016dc4, 32'hc182ba15, 32'h413ae2ae, 32'h42517748, 32'h426e5451, 32'hc2035ce6, 32'h419747d1};
test_output[21192:21199] = '{32'h0, 32'h0, 32'h0, 32'h413ae2ae, 32'h42517748, 32'h426e5451, 32'h0, 32'h419747d1};
test_input[21200:21207] = '{32'hc28df9b8, 32'hc2a0b443, 32'hc2add68b, 32'h42764450, 32'hc1f31f7a, 32'hc25c5525, 32'h42b9089b, 32'h42669009};
test_output[21200:21207] = '{32'h0, 32'h0, 32'h0, 32'h42764450, 32'h0, 32'h0, 32'h42b9089b, 32'h42669009};
test_input[21208:21215] = '{32'hc27e6c61, 32'hc0050be6, 32'h42a17750, 32'hc211b9cd, 32'hc236b9e0, 32'hc26ec0d4, 32'hc1a24386, 32'h425c1ba1};
test_output[21208:21215] = '{32'h0, 32'h0, 32'h42a17750, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425c1ba1};
test_input[21216:21223] = '{32'hc099e6a3, 32'h428be5e9, 32'h42ba0a47, 32'hc2995428, 32'h40e125e5, 32'hc2446786, 32'hc21f67df, 32'h4285149a};
test_output[21216:21223] = '{32'h0, 32'h428be5e9, 32'h42ba0a47, 32'h0, 32'h40e125e5, 32'h0, 32'h0, 32'h4285149a};
test_input[21224:21231] = '{32'hbfdc0728, 32'h42458c8b, 32'h426f47ff, 32'hc2b13b9e, 32'hc2947802, 32'hc29565af, 32'hc26c4b50, 32'h42136b3a};
test_output[21224:21231] = '{32'h0, 32'h42458c8b, 32'h426f47ff, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42136b3a};
test_input[21232:21239] = '{32'hc1780459, 32'h41358a12, 32'h4230cbdd, 32'hc2c49371, 32'hc296bcc5, 32'hc2a9d5f6, 32'h416ec80e, 32'hc16d5876};
test_output[21232:21239] = '{32'h0, 32'h41358a12, 32'h4230cbdd, 32'h0, 32'h0, 32'h0, 32'h416ec80e, 32'h0};
test_input[21240:21247] = '{32'hc28c2263, 32'hc2b9705a, 32'h424f7485, 32'h422547cc, 32'hc20eb220, 32'hc2515568, 32'hc265900b, 32'hc2c087e2};
test_output[21240:21247] = '{32'h0, 32'h0, 32'h424f7485, 32'h422547cc, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21248:21255] = '{32'h417bc3a4, 32'h4275582e, 32'h4250a1e8, 32'h413fa2d0, 32'hc28c6152, 32'hc1dbb124, 32'hc21d548e, 32'h42b1af23};
test_output[21248:21255] = '{32'h417bc3a4, 32'h4275582e, 32'h4250a1e8, 32'h413fa2d0, 32'h0, 32'h0, 32'h0, 32'h42b1af23};
test_input[21256:21263] = '{32'h40c1822f, 32'h42184ee0, 32'h42c38fff, 32'h426822c5, 32'hc247c6a6, 32'h42b51eac, 32'h425cd9c3, 32'h42040ef9};
test_output[21256:21263] = '{32'h40c1822f, 32'h42184ee0, 32'h42c38fff, 32'h426822c5, 32'h0, 32'h42b51eac, 32'h425cd9c3, 32'h42040ef9};
test_input[21264:21271] = '{32'hc119c3e0, 32'h41e558e1, 32'hc1802a10, 32'hc15ef063, 32'h4298a4a0, 32'hc2ad42a1, 32'h423f447c, 32'h42281885};
test_output[21264:21271] = '{32'h0, 32'h41e558e1, 32'h0, 32'h0, 32'h4298a4a0, 32'h0, 32'h423f447c, 32'h42281885};
test_input[21272:21279] = '{32'hc27584d6, 32'hc28dc587, 32'h42bafb51, 32'h42c3c05d, 32'hc1923097, 32'hc20e88aa, 32'h41a2c01e, 32'hc2b42b79};
test_output[21272:21279] = '{32'h0, 32'h0, 32'h42bafb51, 32'h42c3c05d, 32'h0, 32'h0, 32'h41a2c01e, 32'h0};
test_input[21280:21287] = '{32'h41c95aa7, 32'h412a1e94, 32'hc2808be0, 32'hc2afe491, 32'hc28cfa39, 32'hc16c2051, 32'h42b0291b, 32'hc0a044fe};
test_output[21280:21287] = '{32'h41c95aa7, 32'h412a1e94, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b0291b, 32'h0};
test_input[21288:21295] = '{32'h4236319b, 32'h42a82460, 32'hc237d7f7, 32'hc28c49c2, 32'hc282d679, 32'hc2c20091, 32'hc28ce0d9, 32'h41d70a8c};
test_output[21288:21295] = '{32'h4236319b, 32'h42a82460, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41d70a8c};
test_input[21296:21303] = '{32'h421edf07, 32'h42825f13, 32'h42a57039, 32'hc1a23809, 32'hc29a4154, 32'h4283498a, 32'h429b0710, 32'hbfd678c4};
test_output[21296:21303] = '{32'h421edf07, 32'h42825f13, 32'h42a57039, 32'h0, 32'h0, 32'h4283498a, 32'h429b0710, 32'h0};
test_input[21304:21311] = '{32'h41f387e2, 32'h42a405f8, 32'hc1fae93f, 32'hc17cc242, 32'hc2924443, 32'h422cbcb0, 32'hc2ab010f, 32'hc0c08a00};
test_output[21304:21311] = '{32'h41f387e2, 32'h42a405f8, 32'h0, 32'h0, 32'h0, 32'h422cbcb0, 32'h0, 32'h0};
test_input[21312:21319] = '{32'h40f86653, 32'hc18f3d0b, 32'hc2989401, 32'h40c144cd, 32'hc2a1a03b, 32'h4294e499, 32'h40a570e5, 32'h40987fa1};
test_output[21312:21319] = '{32'h40f86653, 32'h0, 32'h0, 32'h40c144cd, 32'h0, 32'h4294e499, 32'h40a570e5, 32'h40987fa1};
test_input[21320:21327] = '{32'h420180fe, 32'hc26ab408, 32'h4265c103, 32'h4276e6b1, 32'hc1092eaa, 32'h411d18b9, 32'h420d7142, 32'hc2ab987f};
test_output[21320:21327] = '{32'h420180fe, 32'h0, 32'h4265c103, 32'h4276e6b1, 32'h0, 32'h411d18b9, 32'h420d7142, 32'h0};
test_input[21328:21335] = '{32'h42aeab21, 32'hc12b1a84, 32'h41fdf095, 32'h4211db57, 32'hc23b6dad, 32'h42be3673, 32'h423cf454, 32'h42550e82};
test_output[21328:21335] = '{32'h42aeab21, 32'h0, 32'h41fdf095, 32'h4211db57, 32'h0, 32'h42be3673, 32'h423cf454, 32'h42550e82};
test_input[21336:21343] = '{32'h424c7a6f, 32'h41fd164b, 32'hc2840d5f, 32'h422d58f4, 32'hc2b0a515, 32'h42419c6a, 32'hc1166925, 32'hc2468cc7};
test_output[21336:21343] = '{32'h424c7a6f, 32'h41fd164b, 32'h0, 32'h422d58f4, 32'h0, 32'h42419c6a, 32'h0, 32'h0};
test_input[21344:21351] = '{32'h4104b8e6, 32'hc2b36e49, 32'hc089ab47, 32'h42a80a18, 32'hc27674e6, 32'hc24abbe9, 32'hc2886b70, 32'h4298f0e0};
test_output[21344:21351] = '{32'h4104b8e6, 32'h0, 32'h0, 32'h42a80a18, 32'h0, 32'h0, 32'h0, 32'h4298f0e0};
test_input[21352:21359] = '{32'h42bcb5e2, 32'hc1e850f0, 32'hc27737cf, 32'h41e4a009, 32'hc282371f, 32'h4245a4bb, 32'h41db4f3b, 32'h41a5e811};
test_output[21352:21359] = '{32'h42bcb5e2, 32'h0, 32'h0, 32'h41e4a009, 32'h0, 32'h4245a4bb, 32'h41db4f3b, 32'h41a5e811};
test_input[21360:21367] = '{32'hc28fe6d8, 32'h42abd6a4, 32'hc23916b3, 32'h42507a88, 32'h42009a15, 32'h428d0a5f, 32'h4293c062, 32'h42359e02};
test_output[21360:21367] = '{32'h0, 32'h42abd6a4, 32'h0, 32'h42507a88, 32'h42009a15, 32'h428d0a5f, 32'h4293c062, 32'h42359e02};
test_input[21368:21375] = '{32'hc242993d, 32'h41867946, 32'hc16e1485, 32'h423fc366, 32'hc29ef5ac, 32'hc222b1ed, 32'h429542ca, 32'hc1f21bd8};
test_output[21368:21375] = '{32'h0, 32'h41867946, 32'h0, 32'h423fc366, 32'h0, 32'h0, 32'h429542ca, 32'h0};
test_input[21376:21383] = '{32'h42c0a5e5, 32'hc27d6d6e, 32'hc2b18ac6, 32'hc16c8ada, 32'h424baa0c, 32'hc2a2f1ec, 32'h42994756, 32'h4104755f};
test_output[21376:21383] = '{32'h42c0a5e5, 32'h0, 32'h0, 32'h0, 32'h424baa0c, 32'h0, 32'h42994756, 32'h4104755f};
test_input[21384:21391] = '{32'hc10513e5, 32'hc2ba968a, 32'h42be8ed2, 32'hc25999fc, 32'hc288fa2e, 32'h425f9f0b, 32'h4204244a, 32'h4295ab31};
test_output[21384:21391] = '{32'h0, 32'h0, 32'h42be8ed2, 32'h0, 32'h0, 32'h425f9f0b, 32'h4204244a, 32'h4295ab31};
test_input[21392:21399] = '{32'h4141479d, 32'h42c16539, 32'h42769e34, 32'hc1f67b91, 32'h41bc25d0, 32'hc29af727, 32'h428d85b1, 32'h4098a447};
test_output[21392:21399] = '{32'h4141479d, 32'h42c16539, 32'h42769e34, 32'h0, 32'h41bc25d0, 32'h0, 32'h428d85b1, 32'h4098a447};
test_input[21400:21407] = '{32'h42a2c67b, 32'h42ab9450, 32'hc2998b67, 32'h429f34b6, 32'hc21e918f, 32'h429bdbdc, 32'hc2b40d6f, 32'hc2b8d537};
test_output[21400:21407] = '{32'h42a2c67b, 32'h42ab9450, 32'h0, 32'h429f34b6, 32'h0, 32'h429bdbdc, 32'h0, 32'h0};
test_input[21408:21415] = '{32'h425bf0bc, 32'h42196379, 32'hc196b7bd, 32'hc29bfda8, 32'hc0f5b2c0, 32'h42587887, 32'hc26dd47c, 32'hc2c0cd74};
test_output[21408:21415] = '{32'h425bf0bc, 32'h42196379, 32'h0, 32'h0, 32'h0, 32'h42587887, 32'h0, 32'h0};
test_input[21416:21423] = '{32'h4272fca9, 32'h42b342c0, 32'h42799389, 32'h4168010c, 32'h4247b501, 32'hc2aca9a8, 32'h423bee65, 32'hc08d859a};
test_output[21416:21423] = '{32'h4272fca9, 32'h42b342c0, 32'h42799389, 32'h4168010c, 32'h4247b501, 32'h0, 32'h423bee65, 32'h0};
test_input[21424:21431] = '{32'hc100347d, 32'h4295f4d5, 32'hc277fa47, 32'hc072c869, 32'h418c4d15, 32'hc2562eb5, 32'h423edcdd, 32'h4281f904};
test_output[21424:21431] = '{32'h0, 32'h4295f4d5, 32'h0, 32'h0, 32'h418c4d15, 32'h0, 32'h423edcdd, 32'h4281f904};
test_input[21432:21439] = '{32'hc1e54d0c, 32'hc2359e6b, 32'h42b43180, 32'h42048780, 32'h428b860c, 32'h42297236, 32'hc2bcb03b, 32'h429790c1};
test_output[21432:21439] = '{32'h0, 32'h0, 32'h42b43180, 32'h42048780, 32'h428b860c, 32'h42297236, 32'h0, 32'h429790c1};
test_input[21440:21447] = '{32'h4248b744, 32'hc0cae12b, 32'hc281d1a7, 32'hc23eaee2, 32'hc22174e9, 32'h41981c88, 32'h4298dd7d, 32'h428d559e};
test_output[21440:21447] = '{32'h4248b744, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41981c88, 32'h4298dd7d, 32'h428d559e};
test_input[21448:21455] = '{32'h4280e0b9, 32'hc10cc72b, 32'hc20a9a73, 32'hc1cf870b, 32'h42a12cc2, 32'h42b5eefe, 32'hc20c5b57, 32'h414d1a49};
test_output[21448:21455] = '{32'h4280e0b9, 32'h0, 32'h0, 32'h0, 32'h42a12cc2, 32'h42b5eefe, 32'h0, 32'h414d1a49};
test_input[21456:21463] = '{32'hc2ac18de, 32'h4100cdbf, 32'h42ae3cb4, 32'hc207eb70, 32'hc2b5337a, 32'h42a38c1a, 32'h41974c65, 32'h42c27ae7};
test_output[21456:21463] = '{32'h0, 32'h4100cdbf, 32'h42ae3cb4, 32'h0, 32'h0, 32'h42a38c1a, 32'h41974c65, 32'h42c27ae7};
test_input[21464:21471] = '{32'hc2a732de, 32'h4223d41c, 32'h42610fee, 32'hc2b57f89, 32'hc199d32b, 32'h42c7da36, 32'hc290b420, 32'h4275bbd6};
test_output[21464:21471] = '{32'h0, 32'h4223d41c, 32'h42610fee, 32'h0, 32'h0, 32'h42c7da36, 32'h0, 32'h4275bbd6};
test_input[21472:21479] = '{32'h428a5314, 32'hc05dc138, 32'hc19af765, 32'h42b02015, 32'hc1b56385, 32'h42b8e6f9, 32'h42c7a87c, 32'h42899207};
test_output[21472:21479] = '{32'h428a5314, 32'h0, 32'h0, 32'h42b02015, 32'h0, 32'h42b8e6f9, 32'h42c7a87c, 32'h42899207};
test_input[21480:21487] = '{32'hc2325feb, 32'hc2991643, 32'h42bb0097, 32'h42134ce1, 32'hc1ffcbb7, 32'h414696a0, 32'h42966bfc, 32'hc22fe416};
test_output[21480:21487] = '{32'h0, 32'h0, 32'h42bb0097, 32'h42134ce1, 32'h0, 32'h414696a0, 32'h42966bfc, 32'h0};
test_input[21488:21495] = '{32'h41a6212b, 32'h3ec8ed1e, 32'h41f405f9, 32'hc28a287b, 32'hc1a85d7e, 32'hc0b01489, 32'h40a6b6f2, 32'h4205aeac};
test_output[21488:21495] = '{32'h41a6212b, 32'h3ec8ed1e, 32'h41f405f9, 32'h0, 32'h0, 32'h0, 32'h40a6b6f2, 32'h4205aeac};
test_input[21496:21503] = '{32'h4224c60d, 32'hc2a0beec, 32'hc29fcc76, 32'h41cd2821, 32'hc223e7de, 32'h3e6aa695, 32'h4298de9b, 32'h421299ab};
test_output[21496:21503] = '{32'h4224c60d, 32'h0, 32'h0, 32'h41cd2821, 32'h0, 32'h3e6aa695, 32'h4298de9b, 32'h421299ab};
test_input[21504:21511] = '{32'hc17b1c98, 32'h4286572f, 32'h41afd444, 32'hc2b995c3, 32'hc0491031, 32'hc210ea07, 32'h42118158, 32'hc201f446};
test_output[21504:21511] = '{32'h0, 32'h4286572f, 32'h41afd444, 32'h0, 32'h0, 32'h0, 32'h42118158, 32'h0};
test_input[21512:21519] = '{32'hc2886243, 32'hc13ef210, 32'h420edf13, 32'h4211ae9d, 32'h423f23f8, 32'h421ee057, 32'hc1c0e802, 32'hc28bb850};
test_output[21512:21519] = '{32'h0, 32'h0, 32'h420edf13, 32'h4211ae9d, 32'h423f23f8, 32'h421ee057, 32'h0, 32'h0};
test_input[21520:21527] = '{32'hc233b0d7, 32'h42a57735, 32'hc241c353, 32'hc20e5fe4, 32'h42c004b3, 32'h406e6b1b, 32'h428e4e01, 32'hc1770408};
test_output[21520:21527] = '{32'h0, 32'h42a57735, 32'h0, 32'h0, 32'h42c004b3, 32'h406e6b1b, 32'h428e4e01, 32'h0};
test_input[21528:21535] = '{32'hc216bb63, 32'h41d299b9, 32'h42bcf840, 32'h42179f58, 32'h42c63e5c, 32'h419efddd, 32'hc28b450d, 32'h4290d90f};
test_output[21528:21535] = '{32'h0, 32'h41d299b9, 32'h42bcf840, 32'h42179f58, 32'h42c63e5c, 32'h419efddd, 32'h0, 32'h4290d90f};
test_input[21536:21543] = '{32'hc2c5647a, 32'hc279800a, 32'hc217ed2d, 32'hc2a86608, 32'hc1363054, 32'h4112b4e1, 32'h41a1f2b4, 32'h42a70717};
test_output[21536:21543] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4112b4e1, 32'h41a1f2b4, 32'h42a70717};
test_input[21544:21551] = '{32'h427f6bdc, 32'h422fa948, 32'hc23bdc08, 32'h4177e014, 32'h413c6bdf, 32'h42adeb94, 32'hc2275087, 32'hc2aa746b};
test_output[21544:21551] = '{32'h427f6bdc, 32'h422fa948, 32'h0, 32'h4177e014, 32'h413c6bdf, 32'h42adeb94, 32'h0, 32'h0};
test_input[21552:21559] = '{32'hc297f14b, 32'hc01870bd, 32'h428eb639, 32'hc2482021, 32'hc290ac6e, 32'hc20acaa0, 32'h4292a258, 32'h423bf186};
test_output[21552:21559] = '{32'h0, 32'h0, 32'h428eb639, 32'h0, 32'h0, 32'h0, 32'h4292a258, 32'h423bf186};
test_input[21560:21567] = '{32'h42974d67, 32'h418bcf3f, 32'hc2646b10, 32'h428a1798, 32'hc28c201a, 32'hc2a3f31b, 32'hbf8b425d, 32'h421a0ea7};
test_output[21560:21567] = '{32'h42974d67, 32'h418bcf3f, 32'h0, 32'h428a1798, 32'h0, 32'h0, 32'h0, 32'h421a0ea7};
test_input[21568:21575] = '{32'h41d8128b, 32'h422f9c5a, 32'h42090a73, 32'h428f7403, 32'h41f82ec1, 32'hc19ab5bc, 32'h424dcb0c, 32'h418b96fa};
test_output[21568:21575] = '{32'h41d8128b, 32'h422f9c5a, 32'h42090a73, 32'h428f7403, 32'h41f82ec1, 32'h0, 32'h424dcb0c, 32'h418b96fa};
test_input[21576:21583] = '{32'hc2407cf1, 32'hc2b2b04f, 32'h41c992e5, 32'hc2a4e36d, 32'h41d440c6, 32'h42a7f093, 32'hc270434b, 32'h42c54d90};
test_output[21576:21583] = '{32'h0, 32'h0, 32'h41c992e5, 32'h0, 32'h41d440c6, 32'h42a7f093, 32'h0, 32'h42c54d90};
test_input[21584:21591] = '{32'h42750e3a, 32'h42acb538, 32'h424d179b, 32'hc234492b, 32'h41605756, 32'hc2bd3e64, 32'hc0f9d70c, 32'hc245d687};
test_output[21584:21591] = '{32'h42750e3a, 32'h42acb538, 32'h424d179b, 32'h0, 32'h41605756, 32'h0, 32'h0, 32'h0};
test_input[21592:21599] = '{32'h424756e2, 32'h42ad7bd9, 32'hc1e5ea7f, 32'hc2c38aaf, 32'h42bbbb7b, 32'h4291268c, 32'hc28bf902, 32'h4208b2de};
test_output[21592:21599] = '{32'h424756e2, 32'h42ad7bd9, 32'h0, 32'h0, 32'h42bbbb7b, 32'h4291268c, 32'h0, 32'h4208b2de};
test_input[21600:21607] = '{32'h41508265, 32'hc20cfdd4, 32'h4299f8f5, 32'hc2c07cfe, 32'h42bd4971, 32'h41c7e314, 32'h425826fc, 32'hc106d662};
test_output[21600:21607] = '{32'h41508265, 32'h0, 32'h4299f8f5, 32'h0, 32'h42bd4971, 32'h41c7e314, 32'h425826fc, 32'h0};
test_input[21608:21615] = '{32'hc2752f2a, 32'h42676733, 32'h42bce5a3, 32'hc2108646, 32'h416b62ec, 32'hc29d2407, 32'hc1fbcd3a, 32'hc2a06a08};
test_output[21608:21615] = '{32'h0, 32'h42676733, 32'h42bce5a3, 32'h0, 32'h416b62ec, 32'h0, 32'h0, 32'h0};
test_input[21616:21623] = '{32'hc297cc71, 32'hc1ecd7c0, 32'hc299a507, 32'h42a11f78, 32'hc263bd76, 32'h4132ed68, 32'hc2117b44, 32'hc2b48b1b};
test_output[21616:21623] = '{32'h0, 32'h0, 32'h0, 32'h42a11f78, 32'h0, 32'h4132ed68, 32'h0, 32'h0};
test_input[21624:21631] = '{32'h42c57b18, 32'h42a1d686, 32'hc2a9cb00, 32'h42804afb, 32'h42c25c9e, 32'h42806ab6, 32'h41fc36ee, 32'hc0b0369f};
test_output[21624:21631] = '{32'h42c57b18, 32'h42a1d686, 32'h0, 32'h42804afb, 32'h42c25c9e, 32'h42806ab6, 32'h41fc36ee, 32'h0};
test_input[21632:21639] = '{32'h41f5ed98, 32'hc284b256, 32'h41f54ce0, 32'hc1bcf64b, 32'hc1a2c6f2, 32'h42478b35, 32'hc29660f4, 32'h4267861f};
test_output[21632:21639] = '{32'h41f5ed98, 32'h0, 32'h41f54ce0, 32'h0, 32'h0, 32'h42478b35, 32'h0, 32'h4267861f};
test_input[21640:21647] = '{32'h427c9583, 32'h414484e4, 32'h4200fb5a, 32'hc1cd9762, 32'hc2a902ca, 32'hc22020cd, 32'h421e4b37, 32'hc286e6c4};
test_output[21640:21647] = '{32'h427c9583, 32'h414484e4, 32'h4200fb5a, 32'h0, 32'h0, 32'h0, 32'h421e4b37, 32'h0};
test_input[21648:21655] = '{32'h41be654e, 32'h413a2e69, 32'h427ff44c, 32'hc2aaf04d, 32'hc265b127, 32'h4285da2e, 32'h4268a800, 32'hc2b0c862};
test_output[21648:21655] = '{32'h41be654e, 32'h413a2e69, 32'h427ff44c, 32'h0, 32'h0, 32'h4285da2e, 32'h4268a800, 32'h0};
test_input[21656:21663] = '{32'hc20e1dd9, 32'hc1962afa, 32'hc18a3376, 32'h42bbf3a5, 32'h4299dbc7, 32'h418e840a, 32'hc24f26b1, 32'h42ad1ca4};
test_output[21656:21663] = '{32'h0, 32'h0, 32'h0, 32'h42bbf3a5, 32'h4299dbc7, 32'h418e840a, 32'h0, 32'h42ad1ca4};
test_input[21664:21671] = '{32'hc2526d0f, 32'h41f29876, 32'h4277be67, 32'hc2b61348, 32'h42b0546c, 32'hbf01dbe8, 32'hc1824045, 32'h427c9244};
test_output[21664:21671] = '{32'h0, 32'h41f29876, 32'h4277be67, 32'h0, 32'h42b0546c, 32'h0, 32'h0, 32'h427c9244};
test_input[21672:21679] = '{32'hc25bed1c, 32'hc1c42aef, 32'hc1b7a4ab, 32'h419c2b7e, 32'hc29b6720, 32'h42b0c6a9, 32'hc2a5f6ed, 32'h3f535188};
test_output[21672:21679] = '{32'h0, 32'h0, 32'h0, 32'h419c2b7e, 32'h0, 32'h42b0c6a9, 32'h0, 32'h3f535188};
test_input[21680:21687] = '{32'hc27b67a1, 32'h428729c5, 32'h42c379a1, 32'hc165d5e7, 32'hc22182ff, 32'hc1d20588, 32'h426b14e7, 32'h419f7480};
test_output[21680:21687] = '{32'h0, 32'h428729c5, 32'h42c379a1, 32'h0, 32'h0, 32'h0, 32'h426b14e7, 32'h419f7480};
test_input[21688:21695] = '{32'h419c2372, 32'h427602f7, 32'h41e8ee16, 32'h422e86dc, 32'h425a1e86, 32'hc21bd874, 32'hc21517e6, 32'hc29641f6};
test_output[21688:21695] = '{32'h419c2372, 32'h427602f7, 32'h41e8ee16, 32'h422e86dc, 32'h425a1e86, 32'h0, 32'h0, 32'h0};
test_input[21696:21703] = '{32'h42546abc, 32'h4246a611, 32'hc12e0228, 32'hc276fe5b, 32'hc243f1b3, 32'hc0af33e7, 32'h42a94a6d, 32'hc25aeefd};
test_output[21696:21703] = '{32'h42546abc, 32'h4246a611, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a94a6d, 32'h0};
test_input[21704:21711] = '{32'hc2bcec78, 32'h422717bf, 32'h42c13f85, 32'hc29b83df, 32'hc234f6dc, 32'hc2494327, 32'h419b8ef2, 32'h4286462b};
test_output[21704:21711] = '{32'h0, 32'h422717bf, 32'h42c13f85, 32'h0, 32'h0, 32'h0, 32'h419b8ef2, 32'h4286462b};
test_input[21712:21719] = '{32'h42c46689, 32'hc1dafe0e, 32'hc290bd63, 32'h4271da35, 32'h41b3990e, 32'hc18ec0b8, 32'h42aa9d0f, 32'h4216877c};
test_output[21712:21719] = '{32'h42c46689, 32'h0, 32'h0, 32'h4271da35, 32'h41b3990e, 32'h0, 32'h42aa9d0f, 32'h4216877c};
test_input[21720:21727] = '{32'h42813619, 32'hc2933efa, 32'h40f22bab, 32'hc297caa4, 32'hc2630747, 32'h428fea69, 32'h42bb913f, 32'h42a99b27};
test_output[21720:21727] = '{32'h42813619, 32'h0, 32'h40f22bab, 32'h0, 32'h0, 32'h428fea69, 32'h42bb913f, 32'h42a99b27};
test_input[21728:21735] = '{32'h4289b268, 32'h3f2cc740, 32'hbf47fce4, 32'h4232e14f, 32'hc0a87906, 32'hc11ba4b5, 32'h429d040a, 32'hc11dc354};
test_output[21728:21735] = '{32'h4289b268, 32'h3f2cc740, 32'h0, 32'h4232e14f, 32'h0, 32'h0, 32'h429d040a, 32'h0};
test_input[21736:21743] = '{32'h412b3567, 32'h42b932c8, 32'hc2bb6807, 32'h4274bee2, 32'hc1fbc163, 32'hc2941a63, 32'hc1b2dd86, 32'h4229ec4c};
test_output[21736:21743] = '{32'h412b3567, 32'h42b932c8, 32'h0, 32'h4274bee2, 32'h0, 32'h0, 32'h0, 32'h4229ec4c};
test_input[21744:21751] = '{32'hc234acf7, 32'h41ed065d, 32'h428cc22d, 32'hc2af6f7d, 32'h4236f8ae, 32'hc29f57b1, 32'hc24e6ae4, 32'h42ba4e05};
test_output[21744:21751] = '{32'h0, 32'h41ed065d, 32'h428cc22d, 32'h0, 32'h4236f8ae, 32'h0, 32'h0, 32'h42ba4e05};
test_input[21752:21759] = '{32'h417e0228, 32'h42079ffd, 32'hc27d6c10, 32'h413f444e, 32'hc1d21929, 32'hc2a032c8, 32'hc0e5041d, 32'hc288987d};
test_output[21752:21759] = '{32'h417e0228, 32'h42079ffd, 32'h0, 32'h413f444e, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[21760:21767] = '{32'h42ad03fa, 32'h42aa0273, 32'h42ae1925, 32'hc2850250, 32'hc1a129bf, 32'hc2af61a0, 32'h428db55d, 32'hc2c5eb28};
test_output[21760:21767] = '{32'h42ad03fa, 32'h42aa0273, 32'h42ae1925, 32'h0, 32'h0, 32'h0, 32'h428db55d, 32'h0};
test_input[21768:21775] = '{32'h423cb397, 32'hc2b2098e, 32'h4130fc43, 32'h421f7d1b, 32'h418b91d1, 32'hc1b2ad1d, 32'h40be9caa, 32'hc2ba2807};
test_output[21768:21775] = '{32'h423cb397, 32'h0, 32'h4130fc43, 32'h421f7d1b, 32'h418b91d1, 32'h0, 32'h40be9caa, 32'h0};
test_input[21776:21783] = '{32'hc23a38ac, 32'h428dc3e7, 32'h42a30940, 32'hc26de97c, 32'h42ac4fd1, 32'hc181c95b, 32'hc2a57bbc, 32'h41bbec65};
test_output[21776:21783] = '{32'h0, 32'h428dc3e7, 32'h42a30940, 32'h0, 32'h42ac4fd1, 32'h0, 32'h0, 32'h41bbec65};
test_input[21784:21791] = '{32'hc2302d59, 32'h429dad49, 32'h41a32229, 32'hc1a0ee04, 32'h42aae4ad, 32'hc284bff7, 32'hc1e96322, 32'hc2c58236};
test_output[21784:21791] = '{32'h0, 32'h429dad49, 32'h41a32229, 32'h0, 32'h42aae4ad, 32'h0, 32'h0, 32'h0};
test_input[21792:21799] = '{32'hc1e0133d, 32'hc06984dd, 32'hc2a9441c, 32'h4223855e, 32'h429f4f62, 32'h428cd72f, 32'hc2a91b2c, 32'hc2318699};
test_output[21792:21799] = '{32'h0, 32'h0, 32'h0, 32'h4223855e, 32'h429f4f62, 32'h428cd72f, 32'h0, 32'h0};
test_input[21800:21807] = '{32'hc2965967, 32'hc22e1231, 32'hc2918861, 32'hc1b77265, 32'h3f998316, 32'hc1998f2c, 32'h42893049, 32'hc2852bdf};
test_output[21800:21807] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h3f998316, 32'h0, 32'h42893049, 32'h0};
test_input[21808:21815] = '{32'h42c4e823, 32'hc0974cb8, 32'hc1b478da, 32'hc2a29e8a, 32'hc180849a, 32'h4258633c, 32'hc206c200, 32'hc12ef3b6};
test_output[21808:21815] = '{32'h42c4e823, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4258633c, 32'h0, 32'h0};
test_input[21816:21823] = '{32'h42433d3b, 32'hc122f1c0, 32'h41ce3173, 32'hc2880f7b, 32'hc24365ba, 32'h429b88b6, 32'hc2b9b3f1, 32'h42a2cf43};
test_output[21816:21823] = '{32'h42433d3b, 32'h0, 32'h41ce3173, 32'h0, 32'h0, 32'h429b88b6, 32'h0, 32'h42a2cf43};
test_input[21824:21831] = '{32'h403258c4, 32'hc1e29007, 32'h425fff2b, 32'hc2c1899b, 32'h424635a8, 32'h42021882, 32'hc2626aff, 32'h4230ea3e};
test_output[21824:21831] = '{32'h403258c4, 32'h0, 32'h425fff2b, 32'h0, 32'h424635a8, 32'h42021882, 32'h0, 32'h4230ea3e};
test_input[21832:21839] = '{32'h41a9e856, 32'hc1dfe42e, 32'hc0b7b42b, 32'h42879d83, 32'h42c62a43, 32'hc1f9420d, 32'h40d75836, 32'h42afcb82};
test_output[21832:21839] = '{32'h41a9e856, 32'h0, 32'h0, 32'h42879d83, 32'h42c62a43, 32'h0, 32'h40d75836, 32'h42afcb82};
test_input[21840:21847] = '{32'h42a0155d, 32'h41842d71, 32'hc2882b3d, 32'h428835b6, 32'hc15307b4, 32'h427e8f13, 32'h427e9985, 32'hc26a9856};
test_output[21840:21847] = '{32'h42a0155d, 32'h41842d71, 32'h0, 32'h428835b6, 32'h0, 32'h427e8f13, 32'h427e9985, 32'h0};
test_input[21848:21855] = '{32'h42219fc3, 32'hc052623e, 32'h4295edee, 32'h423b75ab, 32'hc251901a, 32'hc2ac9993, 32'h422031d4, 32'h414330c3};
test_output[21848:21855] = '{32'h42219fc3, 32'h0, 32'h4295edee, 32'h423b75ab, 32'h0, 32'h0, 32'h422031d4, 32'h414330c3};
test_input[21856:21863] = '{32'hc2c78f61, 32'hc2ad4d79, 32'hc20a949a, 32'hc1683fb3, 32'hc251d003, 32'hc2474c45, 32'hc0cfc76a, 32'h429c4bc7};
test_output[21856:21863] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429c4bc7};
test_input[21864:21871] = '{32'hc2a09ce4, 32'hc1ddaf31, 32'hc1a36ad3, 32'hc1b48a44, 32'h40eda3cf, 32'hc203eeb3, 32'hc2885690, 32'h41a28a40};
test_output[21864:21871] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40eda3cf, 32'h0, 32'h0, 32'h41a28a40};
test_input[21872:21879] = '{32'h3fdcebc3, 32'hc00bba81, 32'h42c71c12, 32'h3fa07b0c, 32'h425864dd, 32'hbfa5e7af, 32'h40d0711f, 32'h429d6a49};
test_output[21872:21879] = '{32'h3fdcebc3, 32'h0, 32'h42c71c12, 32'h3fa07b0c, 32'h425864dd, 32'h0, 32'h40d0711f, 32'h429d6a49};
test_input[21880:21887] = '{32'h4219bbc5, 32'hc2484cd6, 32'hc2c1b4a6, 32'h42c65e65, 32'h42afdba3, 32'hc2978c6a, 32'hc23533ac, 32'hc2b93c70};
test_output[21880:21887] = '{32'h4219bbc5, 32'h0, 32'h0, 32'h42c65e65, 32'h42afdba3, 32'h0, 32'h0, 32'h0};
test_input[21888:21895] = '{32'hc2625442, 32'h41b6193d, 32'h42236ca3, 32'hc285ac5d, 32'h4196d239, 32'hc0ad4661, 32'h4283f33b, 32'h42b8a1c1};
test_output[21888:21895] = '{32'h0, 32'h41b6193d, 32'h42236ca3, 32'h0, 32'h4196d239, 32'h0, 32'h4283f33b, 32'h42b8a1c1};
test_input[21896:21903] = '{32'hc001535b, 32'h42ac3aa1, 32'h42c6bc55, 32'h42a21757, 32'h40ea646b, 32'h4128e078, 32'hc2a465ae, 32'h42458189};
test_output[21896:21903] = '{32'h0, 32'h42ac3aa1, 32'h42c6bc55, 32'h42a21757, 32'h40ea646b, 32'h4128e078, 32'h0, 32'h42458189};
test_input[21904:21911] = '{32'hc1630f14, 32'h4144ecef, 32'h42392471, 32'hc2a2d2ee, 32'h4088073f, 32'hc2a6118b, 32'h4242b820, 32'hc19d5aef};
test_output[21904:21911] = '{32'h0, 32'h4144ecef, 32'h42392471, 32'h0, 32'h4088073f, 32'h0, 32'h4242b820, 32'h0};
test_input[21912:21919] = '{32'h421cc645, 32'hc1a7d8f1, 32'h4130521f, 32'h410d4f8c, 32'h423ce7ff, 32'hc243c157, 32'h41aacff4, 32'h42a1d268};
test_output[21912:21919] = '{32'h421cc645, 32'h0, 32'h4130521f, 32'h410d4f8c, 32'h423ce7ff, 32'h0, 32'h41aacff4, 32'h42a1d268};
test_input[21920:21927] = '{32'h42302f53, 32'h4282cb12, 32'hc2a4e690, 32'h4280dd8a, 32'hc21f6807, 32'h40fbf6c0, 32'hc2aa3bc9, 32'h40dad0de};
test_output[21920:21927] = '{32'h42302f53, 32'h4282cb12, 32'h0, 32'h4280dd8a, 32'h0, 32'h40fbf6c0, 32'h0, 32'h40dad0de};
test_input[21928:21935] = '{32'hc1c68f3f, 32'hc204b94e, 32'hc27d13c3, 32'h428d63e6, 32'h42261deb, 32'h42a28b51, 32'h42a6d71e, 32'h424630a5};
test_output[21928:21935] = '{32'h0, 32'h0, 32'h0, 32'h428d63e6, 32'h42261deb, 32'h42a28b51, 32'h42a6d71e, 32'h424630a5};
test_input[21936:21943] = '{32'hc195daee, 32'h4216c295, 32'h3fbf8d91, 32'h42b6ddaf, 32'hc245a125, 32'hc207a181, 32'hc2937b02, 32'h40c7c5ac};
test_output[21936:21943] = '{32'h0, 32'h4216c295, 32'h3fbf8d91, 32'h42b6ddaf, 32'h0, 32'h0, 32'h0, 32'h40c7c5ac};
test_input[21944:21951] = '{32'h420c7b27, 32'hc16d80d4, 32'hc1d1b5f3, 32'hc2882fc9, 32'h41a2f0bd, 32'hc2b071e2, 32'h426b07f4, 32'hc139cf06};
test_output[21944:21951] = '{32'h420c7b27, 32'h0, 32'h0, 32'h0, 32'h41a2f0bd, 32'h0, 32'h426b07f4, 32'h0};
test_input[21952:21959] = '{32'h42a6a49b, 32'hc2abcb59, 32'hc2a92189, 32'hc25e8fa7, 32'hc1743393, 32'hc29d106f, 32'h42b4b3b2, 32'h4264ef59};
test_output[21952:21959] = '{32'h42a6a49b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b4b3b2, 32'h4264ef59};
test_input[21960:21967] = '{32'hc2202150, 32'hc2557718, 32'h429d87db, 32'hc196c12c, 32'h42b81723, 32'hc28f47d0, 32'hc2a4075d, 32'hc2a2679a};
test_output[21960:21967] = '{32'h0, 32'h0, 32'h429d87db, 32'h0, 32'h42b81723, 32'h0, 32'h0, 32'h0};
test_input[21968:21975] = '{32'hc24e2f6c, 32'h42b4c525, 32'h42b43ce5, 32'hc282db1d, 32'h40bad75d, 32'h4292c656, 32'h4187983c, 32'h41552fc0};
test_output[21968:21975] = '{32'h0, 32'h42b4c525, 32'h42b43ce5, 32'h0, 32'h40bad75d, 32'h4292c656, 32'h4187983c, 32'h41552fc0};
test_input[21976:21983] = '{32'hc2b8ba2b, 32'hc2a6a5d4, 32'h4291b2c5, 32'h41959224, 32'h417a5e31, 32'hc275939b, 32'h42a10fcd, 32'h429afa2c};
test_output[21976:21983] = '{32'h0, 32'h0, 32'h4291b2c5, 32'h41959224, 32'h417a5e31, 32'h0, 32'h42a10fcd, 32'h429afa2c};
test_input[21984:21991] = '{32'h42a45245, 32'hc26d23ca, 32'hc18f1367, 32'h41261730, 32'h4251aa4f, 32'h42a381bd, 32'hc2416510, 32'hc260796f};
test_output[21984:21991] = '{32'h42a45245, 32'h0, 32'h0, 32'h41261730, 32'h4251aa4f, 32'h42a381bd, 32'h0, 32'h0};
test_input[21992:21999] = '{32'hc29c5a81, 32'hc14ad254, 32'h424730e0, 32'hc2b10f2f, 32'h413a27e2, 32'h41dd7e39, 32'h42ac7116, 32'hc2b3e990};
test_output[21992:21999] = '{32'h0, 32'h0, 32'h424730e0, 32'h0, 32'h413a27e2, 32'h41dd7e39, 32'h42ac7116, 32'h0};
test_input[22000:22007] = '{32'hc2c5ac16, 32'hc0fdf242, 32'h422f80c0, 32'hc1d65ca6, 32'h41ede194, 32'h4275d668, 32'h42a0ab8b, 32'hc248ef99};
test_output[22000:22007] = '{32'h0, 32'h0, 32'h422f80c0, 32'h0, 32'h41ede194, 32'h4275d668, 32'h42a0ab8b, 32'h0};
test_input[22008:22015] = '{32'h41e36e3d, 32'h42bcd57d, 32'hc13b864d, 32'hc1a2e62d, 32'h428e545c, 32'hc0e20532, 32'h42b8c746, 32'h40befcaf};
test_output[22008:22015] = '{32'h41e36e3d, 32'h42bcd57d, 32'h0, 32'h0, 32'h428e545c, 32'h0, 32'h42b8c746, 32'h40befcaf};
test_input[22016:22023] = '{32'h42c4480e, 32'hc24b11d4, 32'hc28aee1a, 32'hc22a9a0c, 32'hc0d2f03b, 32'hc11ecd28, 32'hc24db8ba, 32'hc2b735ae};
test_output[22016:22023] = '{32'h42c4480e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22024:22031] = '{32'h41ff5a30, 32'h419f3fd9, 32'hc21c0c56, 32'hc1708f67, 32'hc27ad0b5, 32'h428241cd, 32'hc2218091, 32'hc2640598};
test_output[22024:22031] = '{32'h41ff5a30, 32'h419f3fd9, 32'h0, 32'h0, 32'h0, 32'h428241cd, 32'h0, 32'h0};
test_input[22032:22039] = '{32'hc122bdfc, 32'h42356e19, 32'h428f2f44, 32'h420bce7a, 32'h42a4cd8d, 32'hc29933ad, 32'hc28c89e8, 32'hc2668a12};
test_output[22032:22039] = '{32'h0, 32'h42356e19, 32'h428f2f44, 32'h420bce7a, 32'h42a4cd8d, 32'h0, 32'h0, 32'h0};
test_input[22040:22047] = '{32'h41df0895, 32'h41d30f4b, 32'h4261fbb8, 32'hc27e321f, 32'h424be3f5, 32'h410f0f7d, 32'hc0f61a25, 32'h41c49924};
test_output[22040:22047] = '{32'h41df0895, 32'h41d30f4b, 32'h4261fbb8, 32'h0, 32'h424be3f5, 32'h410f0f7d, 32'h0, 32'h41c49924};
test_input[22048:22055] = '{32'h4217b732, 32'hc230750f, 32'h42bb0c8d, 32'hc29c334a, 32'hc2617169, 32'hbfe81290, 32'h4067a66a, 32'hc22078ed};
test_output[22048:22055] = '{32'h4217b732, 32'h0, 32'h42bb0c8d, 32'h0, 32'h0, 32'h0, 32'h4067a66a, 32'h0};
test_input[22056:22063] = '{32'h4180940f, 32'hc272b2af, 32'h42170200, 32'hc23881be, 32'hc042f139, 32'hc2190c29, 32'h42c0ca2d, 32'hc28838eb};
test_output[22056:22063] = '{32'h4180940f, 32'h0, 32'h42170200, 32'h0, 32'h0, 32'h0, 32'h42c0ca2d, 32'h0};
test_input[22064:22071] = '{32'h428e39aa, 32'hc26a03bf, 32'h41bdd790, 32'h426f86f1, 32'hc25da8ff, 32'h42109745, 32'h41b98ca2, 32'hc25a7ccf};
test_output[22064:22071] = '{32'h428e39aa, 32'h0, 32'h41bdd790, 32'h426f86f1, 32'h0, 32'h42109745, 32'h41b98ca2, 32'h0};
test_input[22072:22079] = '{32'h429ae668, 32'h421b74a8, 32'h42831a72, 32'hc212c048, 32'hc2a1c753, 32'h41b42b9f, 32'hc278b68b, 32'h40834f41};
test_output[22072:22079] = '{32'h429ae668, 32'h421b74a8, 32'h42831a72, 32'h0, 32'h0, 32'h41b42b9f, 32'h0, 32'h40834f41};
test_input[22080:22087] = '{32'h4250c36a, 32'hc2a3af63, 32'hc0c27db8, 32'h4225bfcd, 32'hc1922b71, 32'h42568bb1, 32'h40432d9a, 32'h429831de};
test_output[22080:22087] = '{32'h4250c36a, 32'h0, 32'h0, 32'h4225bfcd, 32'h0, 32'h42568bb1, 32'h40432d9a, 32'h429831de};
test_input[22088:22095] = '{32'h42bd6097, 32'h42baa71e, 32'hc224f755, 32'hc2977b5d, 32'hc1bd7c3d, 32'h42779b22, 32'hc227f044, 32'hc0a77336};
test_output[22088:22095] = '{32'h42bd6097, 32'h42baa71e, 32'h0, 32'h0, 32'h0, 32'h42779b22, 32'h0, 32'h0};
test_input[22096:22103] = '{32'hc22f6c16, 32'h425204e3, 32'h42973bd9, 32'hc2c3df80, 32'h417c7fcc, 32'h4295ff21, 32'hc20b15f8, 32'h428ff618};
test_output[22096:22103] = '{32'h0, 32'h425204e3, 32'h42973bd9, 32'h0, 32'h417c7fcc, 32'h4295ff21, 32'h0, 32'h428ff618};
test_input[22104:22111] = '{32'hc0fccbf9, 32'hc11fadb9, 32'h42b37ef8, 32'h4292e24c, 32'h42a4834d, 32'h42a87118, 32'h42841bd3, 32'h42084b25};
test_output[22104:22111] = '{32'h0, 32'h0, 32'h42b37ef8, 32'h4292e24c, 32'h42a4834d, 32'h42a87118, 32'h42841bd3, 32'h42084b25};
test_input[22112:22119] = '{32'h40337e0f, 32'hc2a3eb76, 32'hc27b8ab9, 32'hc2c24023, 32'h426146e2, 32'hc2604683, 32'h41d2d77d, 32'hc2aec73d};
test_output[22112:22119] = '{32'h40337e0f, 32'h0, 32'h0, 32'h0, 32'h426146e2, 32'h0, 32'h41d2d77d, 32'h0};
test_input[22120:22127] = '{32'h42b02cd6, 32'h42a38f4a, 32'hc1ae4e5b, 32'hc28f0e02, 32'h42af0738, 32'hc28243c9, 32'h42713921, 32'hc20e2f01};
test_output[22120:22127] = '{32'h42b02cd6, 32'h42a38f4a, 32'h0, 32'h0, 32'h42af0738, 32'h0, 32'h42713921, 32'h0};
test_input[22128:22135] = '{32'hc14205db, 32'hc2ad0b6c, 32'hc15fa8ba, 32'h42a5ab21, 32'hc23417a7, 32'hc263db0d, 32'hc1b0388a, 32'hc2a0cef5};
test_output[22128:22135] = '{32'h0, 32'h0, 32'h0, 32'h42a5ab21, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22136:22143] = '{32'h4159c7d5, 32'hc2018c99, 32'hc2a8262d, 32'hc24a31a7, 32'hc28d15fa, 32'hc177b439, 32'hc1394571, 32'h4255c774};
test_output[22136:22143] = '{32'h4159c7d5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4255c774};
test_input[22144:22151] = '{32'h4264df0d, 32'h41e07ce2, 32'hc18af5f5, 32'h4216e042, 32'h4122ac70, 32'hc282cf9b, 32'hc2438b61, 32'hc10175b2};
test_output[22144:22151] = '{32'h4264df0d, 32'h41e07ce2, 32'h0, 32'h4216e042, 32'h4122ac70, 32'h0, 32'h0, 32'h0};
test_input[22152:22159] = '{32'h42b789fb, 32'h42b39bfe, 32'h4150599b, 32'hc118a7dd, 32'hc0a0a969, 32'hc29a58aa, 32'hc12e6a1e, 32'h41648a4b};
test_output[22152:22159] = '{32'h42b789fb, 32'h42b39bfe, 32'h4150599b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41648a4b};
test_input[22160:22167] = '{32'h40b06bb1, 32'h428aae85, 32'h3ff99e8c, 32'h4287014c, 32'h4182df1c, 32'h42aa14d9, 32'hc1acdcb1, 32'h40dcb6e2};
test_output[22160:22167] = '{32'h40b06bb1, 32'h428aae85, 32'h3ff99e8c, 32'h4287014c, 32'h4182df1c, 32'h42aa14d9, 32'h0, 32'h40dcb6e2};
test_input[22168:22175] = '{32'hc2980c10, 32'hc25e356d, 32'h41df19e6, 32'hc209bdcc, 32'hc27440e9, 32'h42aef5c0, 32'hc28351e1, 32'h423449cf};
test_output[22168:22175] = '{32'h0, 32'h0, 32'h41df19e6, 32'h0, 32'h0, 32'h42aef5c0, 32'h0, 32'h423449cf};
test_input[22176:22183] = '{32'h41bd3a53, 32'hc25cd5f1, 32'hc279a486, 32'hc2a1c145, 32'h42bb29c7, 32'h42977521, 32'h429f461e, 32'hc2a1199b};
test_output[22176:22183] = '{32'h41bd3a53, 32'h0, 32'h0, 32'h0, 32'h42bb29c7, 32'h42977521, 32'h429f461e, 32'h0};
test_input[22184:22191] = '{32'hc1c8eade, 32'h419dfd74, 32'hc2bea398, 32'h418fd101, 32'hc0c2fb87, 32'h425a6a66, 32'h4111b97b, 32'h41e69013};
test_output[22184:22191] = '{32'h0, 32'h419dfd74, 32'h0, 32'h418fd101, 32'h0, 32'h425a6a66, 32'h4111b97b, 32'h41e69013};
test_input[22192:22199] = '{32'hc0ceaafb, 32'hc21aa8aa, 32'h3f3c6a8e, 32'h42095088, 32'h42c798fb, 32'h41f04acf, 32'hc2c3e8c9, 32'hc1d1ee8b};
test_output[22192:22199] = '{32'h0, 32'h0, 32'h3f3c6a8e, 32'h42095088, 32'h42c798fb, 32'h41f04acf, 32'h0, 32'h0};
test_input[22200:22207] = '{32'hc0ae377b, 32'h429fd6a8, 32'hc2ab0e12, 32'hc218e358, 32'h42339cd2, 32'h410cf80c, 32'h4217c4e3, 32'h428e7f36};
test_output[22200:22207] = '{32'h0, 32'h429fd6a8, 32'h0, 32'h0, 32'h42339cd2, 32'h410cf80c, 32'h4217c4e3, 32'h428e7f36};
test_input[22208:22215] = '{32'h429cd454, 32'h426630eb, 32'h4294cb26, 32'hc2941524, 32'hc235cf75, 32'hc18b7c33, 32'h42c2a09d, 32'hc25957c5};
test_output[22208:22215] = '{32'h429cd454, 32'h426630eb, 32'h4294cb26, 32'h0, 32'h0, 32'h0, 32'h42c2a09d, 32'h0};
test_input[22216:22223] = '{32'h42b83c2f, 32'h41347022, 32'hc24f536c, 32'hc15b35e0, 32'h426a04e4, 32'h42b52c26, 32'h418420c7, 32'hc1d6b8af};
test_output[22216:22223] = '{32'h42b83c2f, 32'h41347022, 32'h0, 32'h0, 32'h426a04e4, 32'h42b52c26, 32'h418420c7, 32'h0};
test_input[22224:22231] = '{32'hc2afbbd4, 32'hc28e6dee, 32'hc1c7bca3, 32'hc28d0079, 32'hc1bbdd2f, 32'hc232ad5f, 32'h425673d4, 32'hc21f9a7a};
test_output[22224:22231] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425673d4, 32'h0};
test_input[22232:22239] = '{32'h426a72b1, 32'h428e1e31, 32'hc22eb178, 32'hc15c9cdc, 32'hc2a161da, 32'h42ad212b, 32'hc2001fe7, 32'h417f14c4};
test_output[22232:22239] = '{32'h426a72b1, 32'h428e1e31, 32'h0, 32'h0, 32'h0, 32'h42ad212b, 32'h0, 32'h417f14c4};
test_input[22240:22247] = '{32'h42074fef, 32'h4209c897, 32'h42283277, 32'h41ac38ee, 32'hc29f8641, 32'h428ed496, 32'h425fb7fb, 32'h41f3a484};
test_output[22240:22247] = '{32'h42074fef, 32'h4209c897, 32'h42283277, 32'h41ac38ee, 32'h0, 32'h428ed496, 32'h425fb7fb, 32'h41f3a484};
test_input[22248:22255] = '{32'hc1d39e7f, 32'hc1864b55, 32'h425e5d73, 32'hc20611c1, 32'hc13fee32, 32'h42b14adb, 32'h42821d18, 32'hc2c5828a};
test_output[22248:22255] = '{32'h0, 32'h0, 32'h425e5d73, 32'h0, 32'h0, 32'h42b14adb, 32'h42821d18, 32'h0};
test_input[22256:22263] = '{32'hc2bc9eae, 32'hc0bd7549, 32'h41a991fd, 32'h42a71f55, 32'hc2c4dcc9, 32'hc292b873, 32'hc185aeb3, 32'hc1d8c6ef};
test_output[22256:22263] = '{32'h0, 32'h0, 32'h41a991fd, 32'h42a71f55, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22264:22271] = '{32'h4249906d, 32'hc2af2bcc, 32'hc25c2c83, 32'h422cb13a, 32'hc2a12a44, 32'h4248972b, 32'hbf17339e, 32'hc2311a6b};
test_output[22264:22271] = '{32'h4249906d, 32'h0, 32'h0, 32'h422cb13a, 32'h0, 32'h4248972b, 32'h0, 32'h0};
test_input[22272:22279] = '{32'h424eb30e, 32'h414d4c07, 32'h4238f8eb, 32'hc25c20f2, 32'h40813282, 32'h42878453, 32'hc21a7f3d, 32'hc2c0ce32};
test_output[22272:22279] = '{32'h424eb30e, 32'h414d4c07, 32'h4238f8eb, 32'h0, 32'h40813282, 32'h42878453, 32'h0, 32'h0};
test_input[22280:22287] = '{32'h428d9124, 32'h418eedc0, 32'hc2734215, 32'h428f1d4a, 32'h420c6719, 32'hc1c2533f, 32'h42b0059d, 32'h427b6c7c};
test_output[22280:22287] = '{32'h428d9124, 32'h418eedc0, 32'h0, 32'h428f1d4a, 32'h420c6719, 32'h0, 32'h42b0059d, 32'h427b6c7c};
test_input[22288:22295] = '{32'h41b111f7, 32'hc2809eee, 32'h424475e7, 32'hc2980108, 32'hc2b1c265, 32'h42b56cfb, 32'hc29f850e, 32'hc2386fd4};
test_output[22288:22295] = '{32'h41b111f7, 32'h0, 32'h424475e7, 32'h0, 32'h0, 32'h42b56cfb, 32'h0, 32'h0};
test_input[22296:22303] = '{32'h410f81b3, 32'h42431796, 32'h42a50132, 32'hc02af97d, 32'h42a9166f, 32'hc28e7ffa, 32'h425b5015, 32'h41e1c163};
test_output[22296:22303] = '{32'h410f81b3, 32'h42431796, 32'h42a50132, 32'h0, 32'h42a9166f, 32'h0, 32'h425b5015, 32'h41e1c163};
test_input[22304:22311] = '{32'hc0c5e71d, 32'h4262f7b3, 32'h421ae811, 32'h4255b8a2, 32'h4034e923, 32'hc0d4140c, 32'hc1bcd44f, 32'h42b1fc87};
test_output[22304:22311] = '{32'h0, 32'h4262f7b3, 32'h421ae811, 32'h4255b8a2, 32'h4034e923, 32'h0, 32'h0, 32'h42b1fc87};
test_input[22312:22319] = '{32'hc139281c, 32'h42a0aab8, 32'h42b082da, 32'hc2be8f00, 32'hc2177388, 32'h4278a3ba, 32'hc1c782b4, 32'hc1a233bb};
test_output[22312:22319] = '{32'h0, 32'h42a0aab8, 32'h42b082da, 32'h0, 32'h0, 32'h4278a3ba, 32'h0, 32'h0};
test_input[22320:22327] = '{32'h428e30a0, 32'h4205dbfc, 32'hc074c099, 32'hc046d478, 32'h41aafb82, 32'hc18bc0db, 32'hc182efee, 32'hc275ca31};
test_output[22320:22327] = '{32'h428e30a0, 32'h4205dbfc, 32'h0, 32'h0, 32'h41aafb82, 32'h0, 32'h0, 32'h0};
test_input[22328:22335] = '{32'h40bda41b, 32'hc1be9e87, 32'h42833c8b, 32'h429fa5e7, 32'hc20c249a, 32'h3f33aa43, 32'h42725952, 32'h423b08aa};
test_output[22328:22335] = '{32'h40bda41b, 32'h0, 32'h42833c8b, 32'h429fa5e7, 32'h0, 32'h3f33aa43, 32'h42725952, 32'h423b08aa};
test_input[22336:22343] = '{32'hc0d55a6f, 32'hc1a6cb28, 32'hc164d2ff, 32'hc28c16f5, 32'h41effb93, 32'h4264c0fd, 32'hc2559a40, 32'h42181131};
test_output[22336:22343] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41effb93, 32'h4264c0fd, 32'h0, 32'h42181131};
test_input[22344:22351] = '{32'h4254cd2d, 32'hc29cf8b9, 32'h4283857e, 32'h42b8b3d2, 32'h42b97e01, 32'hc2500088, 32'hc29831ea, 32'hc1db899e};
test_output[22344:22351] = '{32'h4254cd2d, 32'h0, 32'h4283857e, 32'h42b8b3d2, 32'h42b97e01, 32'h0, 32'h0, 32'h0};
test_input[22352:22359] = '{32'hc20c4d68, 32'h41fa5fc4, 32'hc1ff0306, 32'hc1eb5ced, 32'hc284b8f3, 32'hc292ba8b, 32'h42407515, 32'hc1baed16};
test_output[22352:22359] = '{32'h0, 32'h41fa5fc4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42407515, 32'h0};
test_input[22360:22367] = '{32'h40ce0213, 32'h42a105ad, 32'h40ea12e6, 32'h424d2c2f, 32'h42bf6890, 32'hc22c7a7a, 32'h42c4702d, 32'hc23f7afc};
test_output[22360:22367] = '{32'h40ce0213, 32'h42a105ad, 32'h40ea12e6, 32'h424d2c2f, 32'h42bf6890, 32'h0, 32'h42c4702d, 32'h0};
test_input[22368:22375] = '{32'h41a97b99, 32'hc280c32c, 32'hc29c7a93, 32'h4237b642, 32'h428bc557, 32'h412efe28, 32'hc213c066, 32'hc2a89200};
test_output[22368:22375] = '{32'h41a97b99, 32'h0, 32'h0, 32'h4237b642, 32'h428bc557, 32'h412efe28, 32'h0, 32'h0};
test_input[22376:22383] = '{32'hc2a4c8e6, 32'h427058d4, 32'hc2b79b97, 32'hc2104046, 32'h40b7f45c, 32'h41a905b0, 32'h423497c8, 32'hc2987f37};
test_output[22376:22383] = '{32'h0, 32'h427058d4, 32'h0, 32'h0, 32'h40b7f45c, 32'h41a905b0, 32'h423497c8, 32'h0};
test_input[22384:22391] = '{32'hc2b6969b, 32'h42ad4c90, 32'hc2b6ec60, 32'hc0a17040, 32'h41ca562a, 32'h42aeaac3, 32'h410be316, 32'hc24ae1eb};
test_output[22384:22391] = '{32'h0, 32'h42ad4c90, 32'h0, 32'h0, 32'h41ca562a, 32'h42aeaac3, 32'h410be316, 32'h0};
test_input[22392:22399] = '{32'hc25fea74, 32'hc2c5b24f, 32'h418ead3d, 32'h4262f046, 32'hc244d6e9, 32'h42c003e4, 32'hc268686f, 32'h41bd3850};
test_output[22392:22399] = '{32'h0, 32'h0, 32'h418ead3d, 32'h4262f046, 32'h0, 32'h42c003e4, 32'h0, 32'h41bd3850};
test_input[22400:22407] = '{32'h42a0be71, 32'hc28efc18, 32'h42178bfb, 32'h425d2f41, 32'hc2a8c2f0, 32'hc20e3797, 32'h423c227c, 32'h41c8d2de};
test_output[22400:22407] = '{32'h42a0be71, 32'h0, 32'h42178bfb, 32'h425d2f41, 32'h0, 32'h0, 32'h423c227c, 32'h41c8d2de};
test_input[22408:22415] = '{32'h424d6be5, 32'h42bc1182, 32'hc1c401b9, 32'h40d5ebc7, 32'h4173da0a, 32'h42968882, 32'hc2a7eb66, 32'hc2b93aac};
test_output[22408:22415] = '{32'h424d6be5, 32'h42bc1182, 32'h0, 32'h40d5ebc7, 32'h4173da0a, 32'h42968882, 32'h0, 32'h0};
test_input[22416:22423] = '{32'hc24674b6, 32'h4234a39b, 32'h42abb15c, 32'hc1843761, 32'hc2029bcc, 32'hc2577879, 32'hc22d7bd6, 32'hc18992a4};
test_output[22416:22423] = '{32'h0, 32'h4234a39b, 32'h42abb15c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22424:22431] = '{32'hc2a35035, 32'hc231450a, 32'h42bf9649, 32'h424e3457, 32'hc155532e, 32'hc2b00f27, 32'h426eda29, 32'h422839c4};
test_output[22424:22431] = '{32'h0, 32'h0, 32'h42bf9649, 32'h424e3457, 32'h0, 32'h0, 32'h426eda29, 32'h422839c4};
test_input[22432:22439] = '{32'hc1188ff2, 32'hc19d72ce, 32'h41c6dfd5, 32'h42c56e54, 32'hc22e09e9, 32'hc26c923e, 32'h40304bf7, 32'hc21eb432};
test_output[22432:22439] = '{32'h0, 32'h0, 32'h41c6dfd5, 32'h42c56e54, 32'h0, 32'h0, 32'h40304bf7, 32'h0};
test_input[22440:22447] = '{32'hc2024b6d, 32'hc1a55f80, 32'h423d888a, 32'hc2766fc6, 32'h42929f02, 32'h4256071f, 32'hc1d84170, 32'h423ba129};
test_output[22440:22447] = '{32'h0, 32'h0, 32'h423d888a, 32'h0, 32'h42929f02, 32'h4256071f, 32'h0, 32'h423ba129};
test_input[22448:22455] = '{32'hc22f2394, 32'h41b5d1b2, 32'h428e0da7, 32'h428c5662, 32'h42138a0c, 32'hc24499c7, 32'hc2c0959c, 32'h42b4618b};
test_output[22448:22455] = '{32'h0, 32'h41b5d1b2, 32'h428e0da7, 32'h428c5662, 32'h42138a0c, 32'h0, 32'h0, 32'h42b4618b};
test_input[22456:22463] = '{32'hc212aa16, 32'hc0c239ad, 32'hc183e9f2, 32'h421397fd, 32'hc216d66e, 32'hc14e53ec, 32'hc27ab9b2, 32'hc24e162a};
test_output[22456:22463] = '{32'h0, 32'h0, 32'h0, 32'h421397fd, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22464:22471] = '{32'hc0d86169, 32'hc2bd5392, 32'hc2b12844, 32'h429f6460, 32'hc1c4b22a, 32'hc28ea49a, 32'h4249581d, 32'hc215787d};
test_output[22464:22471] = '{32'h0, 32'h0, 32'h0, 32'h429f6460, 32'h0, 32'h0, 32'h4249581d, 32'h0};
test_input[22472:22479] = '{32'h40c57fca, 32'hc2c4b7d4, 32'hc271c957, 32'h41c99098, 32'h3fd154dc, 32'hc04b501a, 32'h412d7109, 32'h42bd6502};
test_output[22472:22479] = '{32'h40c57fca, 32'h0, 32'h0, 32'h41c99098, 32'h3fd154dc, 32'h0, 32'h412d7109, 32'h42bd6502};
test_input[22480:22487] = '{32'hc29f1e83, 32'hc2a5983a, 32'hc1f8b591, 32'h425ca844, 32'hc0a74039, 32'hc213a4f5, 32'hc2c1f4b7, 32'hc134f106};
test_output[22480:22487] = '{32'h0, 32'h0, 32'h0, 32'h425ca844, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22488:22495] = '{32'h4142126e, 32'hc2968fb0, 32'hc122ad71, 32'hc08dc2ce, 32'h4298ebc0, 32'hc25ec637, 32'hc14a397e, 32'h427783cb};
test_output[22488:22495] = '{32'h4142126e, 32'h0, 32'h0, 32'h0, 32'h4298ebc0, 32'h0, 32'h0, 32'h427783cb};
test_input[22496:22503] = '{32'h420a43c2, 32'hc264fd30, 32'h42718587, 32'hc2c659a9, 32'h40345a4b, 32'hc142d8e4, 32'h429a54bb, 32'h4127c669};
test_output[22496:22503] = '{32'h420a43c2, 32'h0, 32'h42718587, 32'h0, 32'h40345a4b, 32'h0, 32'h429a54bb, 32'h4127c669};
test_input[22504:22511] = '{32'hc28d61e0, 32'hc00f262d, 32'hc29bb42b, 32'h42207828, 32'h427b1f12, 32'h41932d34, 32'hc288f1ae, 32'h4205945a};
test_output[22504:22511] = '{32'h0, 32'h0, 32'h0, 32'h42207828, 32'h427b1f12, 32'h41932d34, 32'h0, 32'h4205945a};
test_input[22512:22519] = '{32'h42c30559, 32'hc04d3ed4, 32'h41813b58, 32'hc23e1555, 32'h41ce6d96, 32'hc17f1035, 32'h426ad962, 32'h41f756bd};
test_output[22512:22519] = '{32'h42c30559, 32'h0, 32'h41813b58, 32'h0, 32'h41ce6d96, 32'h0, 32'h426ad962, 32'h41f756bd};
test_input[22520:22527] = '{32'hc1f0314f, 32'hc193318b, 32'hc2b9657b, 32'h41884469, 32'hc1c297fd, 32'h422c6e7a, 32'hc10d4a29, 32'h41af0bdc};
test_output[22520:22527] = '{32'h0, 32'h0, 32'h0, 32'h41884469, 32'h0, 32'h422c6e7a, 32'h0, 32'h41af0bdc};
test_input[22528:22535] = '{32'h421abde8, 32'hc1765cac, 32'h42c204cc, 32'h42652ed8, 32'hc28bb150, 32'h42078957, 32'hc1b64482, 32'h41a22b01};
test_output[22528:22535] = '{32'h421abde8, 32'h0, 32'h42c204cc, 32'h42652ed8, 32'h0, 32'h42078957, 32'h0, 32'h41a22b01};
test_input[22536:22543] = '{32'h42b7f4c6, 32'h427d26c1, 32'hc1b2c42f, 32'h410fff70, 32'h4232f1a8, 32'hc1b31c1e, 32'h4244928b, 32'h42821fac};
test_output[22536:22543] = '{32'h42b7f4c6, 32'h427d26c1, 32'h0, 32'h410fff70, 32'h4232f1a8, 32'h0, 32'h4244928b, 32'h42821fac};
test_input[22544:22551] = '{32'h42567d9b, 32'hc1be2b27, 32'h4203dec0, 32'h41f2dd66, 32'h40c1ff25, 32'hc28d8510, 32'h4244807d, 32'hc2374033};
test_output[22544:22551] = '{32'h42567d9b, 32'h0, 32'h4203dec0, 32'h41f2dd66, 32'h40c1ff25, 32'h0, 32'h4244807d, 32'h0};
test_input[22552:22559] = '{32'hc2b44287, 32'hc2a4a4fe, 32'hc1e58801, 32'h421594ef, 32'hc2990964, 32'hc1a949b7, 32'h42b1415f, 32'h4232a475};
test_output[22552:22559] = '{32'h0, 32'h0, 32'h0, 32'h421594ef, 32'h0, 32'h0, 32'h42b1415f, 32'h4232a475};
test_input[22560:22567] = '{32'hc2acb720, 32'h428582cc, 32'h3fab447a, 32'hc28a495f, 32'h41620cf7, 32'h42394c91, 32'h41f1d49a, 32'h3f60efc1};
test_output[22560:22567] = '{32'h0, 32'h428582cc, 32'h3fab447a, 32'h0, 32'h41620cf7, 32'h42394c91, 32'h41f1d49a, 32'h3f60efc1};
test_input[22568:22575] = '{32'hc29a09e6, 32'h40a154d6, 32'h428a5167, 32'hc2b81dcb, 32'hc2a14a9d, 32'hc2a6f51c, 32'hc2a8b8bc, 32'hc1f5620d};
test_output[22568:22575] = '{32'h0, 32'h40a154d6, 32'h428a5167, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22576:22583] = '{32'hc22acc66, 32'hc25e0d01, 32'hc1ae470d, 32'hc282532c, 32'h41d5dac4, 32'hc245a787, 32'h41d87138, 32'hc2b39f04};
test_output[22576:22583] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41d5dac4, 32'h0, 32'h41d87138, 32'h0};
test_input[22584:22591] = '{32'hc2c1dc72, 32'h42526998, 32'h42bc0585, 32'hc071f309, 32'h42a416f2, 32'hc16db953, 32'h41548349, 32'hc0f8701d};
test_output[22584:22591] = '{32'h0, 32'h42526998, 32'h42bc0585, 32'h0, 32'h42a416f2, 32'h0, 32'h41548349, 32'h0};
test_input[22592:22599] = '{32'h42203b4c, 32'h41dc2430, 32'hc1f57e84, 32'h42916be1, 32'hc2847951, 32'hc1ba9644, 32'h42b7f4c9, 32'h414d2d0f};
test_output[22592:22599] = '{32'h42203b4c, 32'h41dc2430, 32'h0, 32'h42916be1, 32'h0, 32'h0, 32'h42b7f4c9, 32'h414d2d0f};
test_input[22600:22607] = '{32'h42a3a900, 32'h4277d5a2, 32'hc2b7eae6, 32'hc2401797, 32'h427a1410, 32'h42b316e7, 32'hc2a55fb7, 32'h41c64d64};
test_output[22600:22607] = '{32'h42a3a900, 32'h4277d5a2, 32'h0, 32'h0, 32'h427a1410, 32'h42b316e7, 32'h0, 32'h41c64d64};
test_input[22608:22615] = '{32'h40d347aa, 32'hc22c548a, 32'hc1af2d2a, 32'h42838b4f, 32'h42647439, 32'h42b9b7fd, 32'h42ac2d8d, 32'h42148804};
test_output[22608:22615] = '{32'h40d347aa, 32'h0, 32'h0, 32'h42838b4f, 32'h42647439, 32'h42b9b7fd, 32'h42ac2d8d, 32'h42148804};
test_input[22616:22623] = '{32'h423f4d52, 32'hc237bb35, 32'hc2c7637a, 32'hc2c758c5, 32'hc1f658c2, 32'hc09cd2f1, 32'h422e507d, 32'h41f4e5fc};
test_output[22616:22623] = '{32'h423f4d52, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422e507d, 32'h41f4e5fc};
test_input[22624:22631] = '{32'h42ae979a, 32'hc15a72bb, 32'h42a95dee, 32'h42b5938b, 32'h41eb9ec6, 32'hc16108e4, 32'hc28af372, 32'hc2440bba};
test_output[22624:22631] = '{32'h42ae979a, 32'h0, 32'h42a95dee, 32'h42b5938b, 32'h41eb9ec6, 32'h0, 32'h0, 32'h0};
test_input[22632:22639] = '{32'h42b4ecdf, 32'hc0c8106a, 32'h40ee1882, 32'hc1fbc023, 32'hc1a05dec, 32'h40e78e76, 32'h408c9163, 32'h427d6f8d};
test_output[22632:22639] = '{32'h42b4ecdf, 32'h0, 32'h40ee1882, 32'h0, 32'h0, 32'h40e78e76, 32'h408c9163, 32'h427d6f8d};
test_input[22640:22647] = '{32'hc13cdd4a, 32'h422db441, 32'hc2a5bf26, 32'h403c219c, 32'hc236ce03, 32'h41973975, 32'h42a6cb86, 32'hc267e2f9};
test_output[22640:22647] = '{32'h0, 32'h422db441, 32'h0, 32'h403c219c, 32'h0, 32'h41973975, 32'h42a6cb86, 32'h0};
test_input[22648:22655] = '{32'h41fee4c1, 32'hc22752c9, 32'h42c45d5e, 32'hc2c12430, 32'hc11f5255, 32'hc26e9ddc, 32'h4294feb2, 32'h42a4c474};
test_output[22648:22655] = '{32'h41fee4c1, 32'h0, 32'h42c45d5e, 32'h0, 32'h0, 32'h0, 32'h4294feb2, 32'h42a4c474};
test_input[22656:22663] = '{32'h40b8593d, 32'h4188b509, 32'h42157bd4, 32'hc2349256, 32'h4208b676, 32'hc20d8ca7, 32'h4101dc55, 32'hc25936a1};
test_output[22656:22663] = '{32'h40b8593d, 32'h4188b509, 32'h42157bd4, 32'h0, 32'h4208b676, 32'h0, 32'h4101dc55, 32'h0};
test_input[22664:22671] = '{32'h42bcf67f, 32'hc25f99a6, 32'h428911f7, 32'hc2899b70, 32'hc090b5f8, 32'hc18f3988, 32'hc1723c4a, 32'hc2461f01};
test_output[22664:22671] = '{32'h42bcf67f, 32'h0, 32'h428911f7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22672:22679] = '{32'h4290c6a3, 32'h41d2656c, 32'hc28a193f, 32'h42c766fe, 32'h42c4f2a7, 32'h3f23eff7, 32'h41dbda26, 32'h429d71fc};
test_output[22672:22679] = '{32'h4290c6a3, 32'h41d2656c, 32'h0, 32'h42c766fe, 32'h42c4f2a7, 32'h3f23eff7, 32'h41dbda26, 32'h429d71fc};
test_input[22680:22687] = '{32'hc2bcffc9, 32'h423535a7, 32'h4214ebef, 32'hc0a03c7d, 32'hc2c23d1c, 32'hc067e86b, 32'hc2ab5de7, 32'h41959356};
test_output[22680:22687] = '{32'h0, 32'h423535a7, 32'h4214ebef, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41959356};
test_input[22688:22695] = '{32'hc28a1983, 32'hc15baea9, 32'h4225378f, 32'hc22ecbab, 32'h41b4f243, 32'h41916da2, 32'h42810866, 32'h4198716b};
test_output[22688:22695] = '{32'h0, 32'h0, 32'h4225378f, 32'h0, 32'h41b4f243, 32'h41916da2, 32'h42810866, 32'h4198716b};
test_input[22696:22703] = '{32'hc128095f, 32'hc012771e, 32'h4248e4ab, 32'hc295ecb7, 32'h428ae8e0, 32'h428adf12, 32'hc2024e88, 32'hc1c5c2ac};
test_output[22696:22703] = '{32'h0, 32'h0, 32'h4248e4ab, 32'h0, 32'h428ae8e0, 32'h428adf12, 32'h0, 32'h0};
test_input[22704:22711] = '{32'hc29f5eeb, 32'hc295c18a, 32'hc283a179, 32'hc294bd36, 32'hc1e44ba9, 32'hc2a6296a, 32'h42a1cd20, 32'hc2673784};
test_output[22704:22711] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a1cd20, 32'h0};
test_input[22712:22719] = '{32'hc25edbac, 32'h42467432, 32'h41a3cf55, 32'hc0754cce, 32'hc2382635, 32'h42bde264, 32'h417fbeb6, 32'hc218fdb6};
test_output[22712:22719] = '{32'h0, 32'h42467432, 32'h41a3cf55, 32'h0, 32'h0, 32'h42bde264, 32'h417fbeb6, 32'h0};
test_input[22720:22727] = '{32'h427600ba, 32'h42be14fa, 32'h42366b31, 32'hc218bc67, 32'h421d9eea, 32'h42764059, 32'h41c3f01b, 32'h422a0043};
test_output[22720:22727] = '{32'h427600ba, 32'h42be14fa, 32'h42366b31, 32'h0, 32'h421d9eea, 32'h42764059, 32'h41c3f01b, 32'h422a0043};
test_input[22728:22735] = '{32'hc209e66f, 32'h428271a8, 32'h4027a110, 32'h42a66d13, 32'h42106244, 32'h42c7c5b2, 32'hc260b7e2, 32'hc27f4edc};
test_output[22728:22735] = '{32'h0, 32'h428271a8, 32'h4027a110, 32'h42a66d13, 32'h42106244, 32'h42c7c5b2, 32'h0, 32'h0};
test_input[22736:22743] = '{32'h426fc6fa, 32'hc2355e9d, 32'hc2503975, 32'hc15c6d01, 32'hc0a9847b, 32'hc269b684, 32'hc2c49924, 32'hc2469636};
test_output[22736:22743] = '{32'h426fc6fa, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22744:22751] = '{32'hc2a442da, 32'h42980214, 32'h42390056, 32'h419ec69f, 32'hc2b6324d, 32'h42870d28, 32'hc1a40bc6, 32'h429b4938};
test_output[22744:22751] = '{32'h0, 32'h42980214, 32'h42390056, 32'h419ec69f, 32'h0, 32'h42870d28, 32'h0, 32'h429b4938};
test_input[22752:22759] = '{32'h42abd514, 32'h41302955, 32'hc2bf9481, 32'h42193ddb, 32'hc2bf2332, 32'h429775c9, 32'hc2a87eab, 32'hc28813ce};
test_output[22752:22759] = '{32'h42abd514, 32'h41302955, 32'h0, 32'h42193ddb, 32'h0, 32'h429775c9, 32'h0, 32'h0};
test_input[22760:22767] = '{32'hc22d7391, 32'hc2b9e807, 32'hc286b889, 32'hc22ddb66, 32'hc0327413, 32'hc29694c2, 32'h419eebc4, 32'hc1a1c020};
test_output[22760:22767] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h419eebc4, 32'h0};
test_input[22768:22775] = '{32'h429170d2, 32'h42268732, 32'h4263dcf4, 32'hc2339567, 32'hc207c65e, 32'hc2365a00, 32'hc278bbdf, 32'h4158c3c4};
test_output[22768:22775] = '{32'h429170d2, 32'h42268732, 32'h4263dcf4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4158c3c4};
test_input[22776:22783] = '{32'hc2a475a5, 32'h4276faf6, 32'hc1b51cbc, 32'hbffac2cb, 32'h40a069f1, 32'h4241971c, 32'h42bace49, 32'h4220ed93};
test_output[22776:22783] = '{32'h0, 32'h4276faf6, 32'h0, 32'h0, 32'h40a069f1, 32'h4241971c, 32'h42bace49, 32'h4220ed93};
test_input[22784:22791] = '{32'hc27cc53a, 32'hc2479c1d, 32'h421a4b25, 32'hc2ac7f46, 32'h41c326e9, 32'hc277dd4b, 32'hc232b5c7, 32'h42718021};
test_output[22784:22791] = '{32'h0, 32'h0, 32'h421a4b25, 32'h0, 32'h41c326e9, 32'h0, 32'h0, 32'h42718021};
test_input[22792:22799] = '{32'hc06e2735, 32'hc28dbd5b, 32'hc1d8197e, 32'hc299c74c, 32'h426e86e3, 32'h42c4321c, 32'h42abfbee, 32'h400ca615};
test_output[22792:22799] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h426e86e3, 32'h42c4321c, 32'h42abfbee, 32'h400ca615};
test_input[22800:22807] = '{32'h429c6481, 32'h424173a4, 32'h428e1946, 32'hc226b9a7, 32'h410557c6, 32'h42ab0982, 32'h41db1c28, 32'hc14f5ba4};
test_output[22800:22807] = '{32'h429c6481, 32'h424173a4, 32'h428e1946, 32'h0, 32'h410557c6, 32'h42ab0982, 32'h41db1c28, 32'h0};
test_input[22808:22815] = '{32'h40dd6ba4, 32'h42653029, 32'hc1a6aceb, 32'h4288b4d5, 32'h41c8bb91, 32'hc19a86bb, 32'h4206b5c7, 32'h42325526};
test_output[22808:22815] = '{32'h40dd6ba4, 32'h42653029, 32'h0, 32'h4288b4d5, 32'h41c8bb91, 32'h0, 32'h4206b5c7, 32'h42325526};
test_input[22816:22823] = '{32'hc2c47208, 32'h42193890, 32'hc1072144, 32'hc1914141, 32'hc1eff820, 32'hc281f696, 32'h429c0fae, 32'h4244a039};
test_output[22816:22823] = '{32'h0, 32'h42193890, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429c0fae, 32'h4244a039};
test_input[22824:22831] = '{32'h421f3639, 32'hc2411265, 32'hc2b5765e, 32'hc21a9cfe, 32'hc23427dc, 32'hc1645d49, 32'h4159a18f, 32'hc1efa1de};
test_output[22824:22831] = '{32'h421f3639, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4159a18f, 32'h0};
test_input[22832:22839] = '{32'h42484fd6, 32'h424c5ae9, 32'h425f4694, 32'hc26ab4bf, 32'hc28945ae, 32'hc04a4e8b, 32'hc19a6456, 32'hc29d8c02};
test_output[22832:22839] = '{32'h42484fd6, 32'h424c5ae9, 32'h425f4694, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[22840:22847] = '{32'h4191df7f, 32'hc1a84cce, 32'h427ed659, 32'h42acf305, 32'h4221cd6e, 32'h42a4295e, 32'h407cdfa9, 32'h417edb31};
test_output[22840:22847] = '{32'h4191df7f, 32'h0, 32'h427ed659, 32'h42acf305, 32'h4221cd6e, 32'h42a4295e, 32'h407cdfa9, 32'h417edb31};
test_input[22848:22855] = '{32'h427aadfb, 32'hc218a5bf, 32'hc1adba0d, 32'h42a27ddf, 32'h42444155, 32'h416bcf80, 32'hc1784365, 32'h3f570251};
test_output[22848:22855] = '{32'h427aadfb, 32'h0, 32'h0, 32'h42a27ddf, 32'h42444155, 32'h416bcf80, 32'h0, 32'h3f570251};
test_input[22856:22863] = '{32'h42c270be, 32'hc29b11ee, 32'h42448c4a, 32'hbff16d23, 32'hc25a1cc2, 32'h4236d127, 32'h42b50749, 32'hc16dcf5d};
test_output[22856:22863] = '{32'h42c270be, 32'h0, 32'h42448c4a, 32'h0, 32'h0, 32'h4236d127, 32'h42b50749, 32'h0};
test_input[22864:22871] = '{32'hc27e0991, 32'hc2be9716, 32'h41d9b61a, 32'h42548f09, 32'h42bcded2, 32'hc2308cc3, 32'hc013465a, 32'h424e70c2};
test_output[22864:22871] = '{32'h0, 32'h0, 32'h41d9b61a, 32'h42548f09, 32'h42bcded2, 32'h0, 32'h0, 32'h424e70c2};
test_input[22872:22879] = '{32'hc1a46ea7, 32'h42254f4e, 32'hc214c297, 32'h423460f8, 32'hc2a9c887, 32'hc24b156f, 32'h42465ac0, 32'hc2b8670a};
test_output[22872:22879] = '{32'h0, 32'h42254f4e, 32'h0, 32'h423460f8, 32'h0, 32'h0, 32'h42465ac0, 32'h0};
test_input[22880:22887] = '{32'h42921d83, 32'hc1033bcd, 32'h4279502a, 32'h41bab93a, 32'h418e9122, 32'h422399ca, 32'hc2a0d892, 32'h41ef1ca0};
test_output[22880:22887] = '{32'h42921d83, 32'h0, 32'h4279502a, 32'h41bab93a, 32'h418e9122, 32'h422399ca, 32'h0, 32'h41ef1ca0};
test_input[22888:22895] = '{32'h429511da, 32'hc1ec274b, 32'hc2787700, 32'hc2610827, 32'h411a403b, 32'hc2a40e12, 32'h42a03a96, 32'hc2c4dcca};
test_output[22888:22895] = '{32'h429511da, 32'h0, 32'h0, 32'h0, 32'h411a403b, 32'h0, 32'h42a03a96, 32'h0};
test_input[22896:22903] = '{32'hc285fd73, 32'h42774824, 32'h417735d2, 32'h4206140e, 32'h425490ad, 32'h407fce82, 32'h42a06475, 32'hc2a4e141};
test_output[22896:22903] = '{32'h0, 32'h42774824, 32'h417735d2, 32'h4206140e, 32'h425490ad, 32'h407fce82, 32'h42a06475, 32'h0};
test_input[22904:22911] = '{32'hc2bc21dd, 32'h4282d79d, 32'h42974237, 32'h42c456ba, 32'hc276244c, 32'hc17a4a5b, 32'hc11da040, 32'h428eba3e};
test_output[22904:22911] = '{32'h0, 32'h4282d79d, 32'h42974237, 32'h42c456ba, 32'h0, 32'h0, 32'h0, 32'h428eba3e};
test_input[22912:22919] = '{32'hc1acd7e9, 32'hc18c0869, 32'h41a0afd7, 32'h4215553d, 32'h4228d7fb, 32'h42bd8171, 32'hc164ca7b, 32'h425ce0e1};
test_output[22912:22919] = '{32'h0, 32'h0, 32'h41a0afd7, 32'h4215553d, 32'h4228d7fb, 32'h42bd8171, 32'h0, 32'h425ce0e1};
test_input[22920:22927] = '{32'h42693c02, 32'hc1b4f95c, 32'h413364cd, 32'h41db85e8, 32'h42a4bcc2, 32'h41b695a2, 32'hc246940d, 32'h41d8025c};
test_output[22920:22927] = '{32'h42693c02, 32'h0, 32'h413364cd, 32'h41db85e8, 32'h42a4bcc2, 32'h41b695a2, 32'h0, 32'h41d8025c};
test_input[22928:22935] = '{32'h42a874d9, 32'hc216a532, 32'h41dcc72e, 32'h4275d8f0, 32'h429c5926, 32'h426db246, 32'h4238e792, 32'hc13a4ac6};
test_output[22928:22935] = '{32'h42a874d9, 32'h0, 32'h41dcc72e, 32'h4275d8f0, 32'h429c5926, 32'h426db246, 32'h4238e792, 32'h0};
test_input[22936:22943] = '{32'h42a95fed, 32'h4200abd0, 32'hc2b996ce, 32'hc19636ca, 32'h424e8714, 32'hc29f4a08, 32'hc1d372c6, 32'hc2871ae2};
test_output[22936:22943] = '{32'h42a95fed, 32'h4200abd0, 32'h0, 32'h0, 32'h424e8714, 32'h0, 32'h0, 32'h0};
test_input[22944:22951] = '{32'h41cc239d, 32'h427ccbbd, 32'h4288c204, 32'h41de1845, 32'h428b6ce0, 32'h429c90a8, 32'h429f271c, 32'hc297b80f};
test_output[22944:22951] = '{32'h41cc239d, 32'h427ccbbd, 32'h4288c204, 32'h41de1845, 32'h428b6ce0, 32'h429c90a8, 32'h429f271c, 32'h0};
test_input[22952:22959] = '{32'h419f1448, 32'h42ad699c, 32'h420661ea, 32'hc2922ac5, 32'h428267a2, 32'hc1c9f427, 32'h423a8e04, 32'hc2154422};
test_output[22952:22959] = '{32'h419f1448, 32'h42ad699c, 32'h420661ea, 32'h0, 32'h428267a2, 32'h0, 32'h423a8e04, 32'h0};
test_input[22960:22967] = '{32'hc111e184, 32'hc27c4b9d, 32'h42a43d40, 32'h427e9eae, 32'h41ca303f, 32'h4047207f, 32'h41b016b7, 32'hc14865c6};
test_output[22960:22967] = '{32'h0, 32'h0, 32'h42a43d40, 32'h427e9eae, 32'h41ca303f, 32'h4047207f, 32'h41b016b7, 32'h0};
test_input[22968:22975] = '{32'hc2880b2a, 32'hc2466727, 32'h41a26156, 32'h411bc46e, 32'hc14ad288, 32'hc2b26599, 32'h42207e41, 32'hc2a51ee1};
test_output[22968:22975] = '{32'h0, 32'h0, 32'h41a26156, 32'h411bc46e, 32'h0, 32'h0, 32'h42207e41, 32'h0};
test_input[22976:22983] = '{32'h410fefa4, 32'hc2a5c8e0, 32'hc29a4d66, 32'h4265752d, 32'h42b87af1, 32'h4231875a, 32'h42acaab9, 32'h4262608e};
test_output[22976:22983] = '{32'h410fefa4, 32'h0, 32'h0, 32'h4265752d, 32'h42b87af1, 32'h4231875a, 32'h42acaab9, 32'h4262608e};
test_input[22984:22991] = '{32'h42954445, 32'h416df7b6, 32'h42a31a18, 32'h422012e6, 32'hc2c33388, 32'h428c2b0b, 32'hc1be9b3e, 32'hc21a977c};
test_output[22984:22991] = '{32'h42954445, 32'h416df7b6, 32'h42a31a18, 32'h422012e6, 32'h0, 32'h428c2b0b, 32'h0, 32'h0};
test_input[22992:22999] = '{32'hc29e3fd6, 32'h4229065a, 32'h42c086b0, 32'hc2ab6c81, 32'h42872ebf, 32'hc1e27d4e, 32'hc234c842, 32'h42831c88};
test_output[22992:22999] = '{32'h0, 32'h4229065a, 32'h42c086b0, 32'h0, 32'h42872ebf, 32'h0, 32'h0, 32'h42831c88};
test_input[23000:23007] = '{32'h41a0d7d2, 32'hc1a7a61a, 32'h418ee975, 32'h4270cc26, 32'hc2961edb, 32'hc29c6b05, 32'hc2873f8b, 32'h4294c612};
test_output[23000:23007] = '{32'h41a0d7d2, 32'h0, 32'h418ee975, 32'h4270cc26, 32'h0, 32'h0, 32'h0, 32'h4294c612};
test_input[23008:23015] = '{32'h41988509, 32'h41e9a3ca, 32'h42c15a31, 32'h4183f781, 32'hc264defb, 32'h42341f14, 32'hc2896584, 32'h3fd3d364};
test_output[23008:23015] = '{32'h41988509, 32'h41e9a3ca, 32'h42c15a31, 32'h4183f781, 32'h0, 32'h42341f14, 32'h0, 32'h3fd3d364};
test_input[23016:23023] = '{32'h42b4ecf4, 32'h42c47e3e, 32'hc20923e2, 32'hc22eaffd, 32'h417e90e8, 32'h41059e16, 32'h42c79a33, 32'h428390a9};
test_output[23016:23023] = '{32'h42b4ecf4, 32'h42c47e3e, 32'h0, 32'h0, 32'h417e90e8, 32'h41059e16, 32'h42c79a33, 32'h428390a9};
test_input[23024:23031] = '{32'h4239a8e4, 32'hc2b72c51, 32'h42533777, 32'h428f6d46, 32'hc1a8eb82, 32'hc294a537, 32'hc1a0c984, 32'h426ff694};
test_output[23024:23031] = '{32'h4239a8e4, 32'h0, 32'h42533777, 32'h428f6d46, 32'h0, 32'h0, 32'h0, 32'h426ff694};
test_input[23032:23039] = '{32'h41ad725e, 32'h425845bb, 32'h42918aa5, 32'h4248f94b, 32'hc20673d4, 32'hc1a4dcb4, 32'h420d937a, 32'hc28e9ab6};
test_output[23032:23039] = '{32'h41ad725e, 32'h425845bb, 32'h42918aa5, 32'h4248f94b, 32'h0, 32'h0, 32'h420d937a, 32'h0};
test_input[23040:23047] = '{32'hc087fccb, 32'hc1d8e4c1, 32'h428f35c6, 32'h42825b7a, 32'hc1a3a566, 32'hc1fae8b1, 32'h420b498d, 32'h42a717d2};
test_output[23040:23047] = '{32'h0, 32'h0, 32'h428f35c6, 32'h42825b7a, 32'h0, 32'h0, 32'h420b498d, 32'h42a717d2};
test_input[23048:23055] = '{32'hc2a12acf, 32'hc227811f, 32'h42310311, 32'h42c271a3, 32'hc11f75ab, 32'h42593f89, 32'h425ed061, 32'h4296faa2};
test_output[23048:23055] = '{32'h0, 32'h0, 32'h42310311, 32'h42c271a3, 32'h0, 32'h42593f89, 32'h425ed061, 32'h4296faa2};
test_input[23056:23063] = '{32'hc26bacf7, 32'hc21ca494, 32'h42929527, 32'hc0d1b5e5, 32'h3f44bc3c, 32'hc2820161, 32'hc1c2f6a0, 32'hc25149cc};
test_output[23056:23063] = '{32'h0, 32'h0, 32'h42929527, 32'h0, 32'h3f44bc3c, 32'h0, 32'h0, 32'h0};
test_input[23064:23071] = '{32'h428d7044, 32'hc2b638a1, 32'h42a47355, 32'hc264255d, 32'h42c28ae7, 32'h42841191, 32'hc20d35b9, 32'hc1fff317};
test_output[23064:23071] = '{32'h428d7044, 32'h0, 32'h42a47355, 32'h0, 32'h42c28ae7, 32'h42841191, 32'h0, 32'h0};
test_input[23072:23079] = '{32'h41a65806, 32'hc2113d38, 32'hc2961598, 32'hc243838f, 32'h42a87340, 32'hc2ba1ccb, 32'hc16f402a, 32'hc12afe0d};
test_output[23072:23079] = '{32'h41a65806, 32'h0, 32'h0, 32'h0, 32'h42a87340, 32'h0, 32'h0, 32'h0};
test_input[23080:23087] = '{32'h41380483, 32'hc29cb23e, 32'hc28e23f2, 32'h42907939, 32'hc2011e7e, 32'hc1f572b1, 32'hc297b7f1, 32'h4293284c};
test_output[23080:23087] = '{32'h41380483, 32'h0, 32'h0, 32'h42907939, 32'h0, 32'h0, 32'h0, 32'h4293284c};
test_input[23088:23095] = '{32'h4285c727, 32'hc03f6941, 32'h42b7ecfe, 32'hc1686b40, 32'h421e6640, 32'hc2929084, 32'h4293a75c, 32'hc25e7ab9};
test_output[23088:23095] = '{32'h4285c727, 32'h0, 32'h42b7ecfe, 32'h0, 32'h421e6640, 32'h0, 32'h4293a75c, 32'h0};
test_input[23096:23103] = '{32'hc1a00752, 32'h42c157f7, 32'hc2a267da, 32'hc2764593, 32'h429aae46, 32'hc26922ad, 32'h3fcf0137, 32'hc2b07f6a};
test_output[23096:23103] = '{32'h0, 32'h42c157f7, 32'h0, 32'h0, 32'h429aae46, 32'h0, 32'h3fcf0137, 32'h0};
test_input[23104:23111] = '{32'h42074340, 32'h4266655f, 32'hc06eb18b, 32'h42b38833, 32'hc2914ef1, 32'hc12af7d7, 32'h41a3e8bc, 32'hc20b5b7b};
test_output[23104:23111] = '{32'h42074340, 32'h4266655f, 32'h0, 32'h42b38833, 32'h0, 32'h0, 32'h41a3e8bc, 32'h0};
test_input[23112:23119] = '{32'h42c6b0ae, 32'hc1deaed3, 32'hc293b35d, 32'h428b6262, 32'hc2a5b536, 32'h41e13c58, 32'hc2bd833c, 32'h42badb27};
test_output[23112:23119] = '{32'h42c6b0ae, 32'h0, 32'h0, 32'h428b6262, 32'h0, 32'h41e13c58, 32'h0, 32'h42badb27};
test_input[23120:23127] = '{32'hc2a607fb, 32'h42963888, 32'hc248db54, 32'hc22eb31c, 32'hc1e3838e, 32'h41897041, 32'hc2acbd65, 32'h4258671d};
test_output[23120:23127] = '{32'h0, 32'h42963888, 32'h0, 32'h0, 32'h0, 32'h41897041, 32'h0, 32'h4258671d};
test_input[23128:23135] = '{32'hc18e5e5f, 32'h41f30ba3, 32'hc16b0945, 32'hc28e9b45, 32'hc24a54ae, 32'hc25db8e0, 32'hc20a8d16, 32'hc2818a6b};
test_output[23128:23135] = '{32'h0, 32'h41f30ba3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23136:23143] = '{32'hc169f464, 32'h417f31b5, 32'hc247cf89, 32'h4292965e, 32'hc26965f4, 32'hc1146719, 32'h40629be0, 32'hc1d0d58f};
test_output[23136:23143] = '{32'h0, 32'h417f31b5, 32'h0, 32'h4292965e, 32'h0, 32'h0, 32'h40629be0, 32'h0};
test_input[23144:23151] = '{32'h42bd3de9, 32'h428d67bf, 32'hc141193c, 32'h4252409a, 32'h424dd507, 32'hc1c5b147, 32'hc0016847, 32'h3fa59236};
test_output[23144:23151] = '{32'h42bd3de9, 32'h428d67bf, 32'h0, 32'h4252409a, 32'h424dd507, 32'h0, 32'h0, 32'h3fa59236};
test_input[23152:23159] = '{32'h4287a829, 32'h40d68d6c, 32'hc0ce156a, 32'h42ae693c, 32'hc2c4daac, 32'hc1122b49, 32'h4282f75f, 32'h42a008eb};
test_output[23152:23159] = '{32'h4287a829, 32'h40d68d6c, 32'h0, 32'h42ae693c, 32'h0, 32'h0, 32'h4282f75f, 32'h42a008eb};
test_input[23160:23167] = '{32'hc2ab081e, 32'hc29956ce, 32'h429e53cb, 32'hc2301f0f, 32'hc0dc77e7, 32'h42ad185e, 32'hc168736e, 32'h4235ad1d};
test_output[23160:23167] = '{32'h0, 32'h0, 32'h429e53cb, 32'h0, 32'h0, 32'h42ad185e, 32'h0, 32'h4235ad1d};
test_input[23168:23175] = '{32'h428d615e, 32'h429ab6d5, 32'h42025266, 32'h428a31b6, 32'hc2360a72, 32'h3f2bd084, 32'hc2c4fd71, 32'hc2aa3d1b};
test_output[23168:23175] = '{32'h428d615e, 32'h429ab6d5, 32'h42025266, 32'h428a31b6, 32'h0, 32'h3f2bd084, 32'h0, 32'h0};
test_input[23176:23183] = '{32'hc22c40cb, 32'h4270a680, 32'h42b8fb79, 32'hc23cfa01, 32'h42c008ac, 32'h422c75a1, 32'hc25946af, 32'hc2c0fa5b};
test_output[23176:23183] = '{32'h0, 32'h4270a680, 32'h42b8fb79, 32'h0, 32'h42c008ac, 32'h422c75a1, 32'h0, 32'h0};
test_input[23184:23191] = '{32'hc10cfdf2, 32'h427da3a2, 32'hc1aaf823, 32'hc17f94e8, 32'h4287f1ec, 32'hc1896e09, 32'h4265c15a, 32'hc2c09578};
test_output[23184:23191] = '{32'h0, 32'h427da3a2, 32'h0, 32'h0, 32'h4287f1ec, 32'h0, 32'h4265c15a, 32'h0};
test_input[23192:23199] = '{32'hc2c3f79f, 32'hc2a8d8b9, 32'hc275ab5f, 32'h422a457f, 32'h429e052d, 32'h423eea28, 32'hc2c6c554, 32'h42bc8758};
test_output[23192:23199] = '{32'h0, 32'h0, 32'h0, 32'h422a457f, 32'h429e052d, 32'h423eea28, 32'h0, 32'h42bc8758};
test_input[23200:23207] = '{32'hc034cc6e, 32'h42690b1f, 32'hc262ebf1, 32'hc2b0c5a1, 32'h4157db1e, 32'h4218bae7, 32'h42a01999, 32'h419ee7b1};
test_output[23200:23207] = '{32'h0, 32'h42690b1f, 32'h0, 32'h0, 32'h4157db1e, 32'h4218bae7, 32'h42a01999, 32'h419ee7b1};
test_input[23208:23215] = '{32'hc17ad5e2, 32'h41dd26f7, 32'h429d95d8, 32'hc1a64a5a, 32'hc2c1cbdc, 32'hc2bd8ac1, 32'h42b54f66, 32'h4290b8fc};
test_output[23208:23215] = '{32'h0, 32'h41dd26f7, 32'h429d95d8, 32'h0, 32'h0, 32'h0, 32'h42b54f66, 32'h4290b8fc};
test_input[23216:23223] = '{32'hc1ead420, 32'hc24eac14, 32'hc1328755, 32'h42c7718a, 32'h429ea4b0, 32'h41f1edfb, 32'hc1048c35, 32'hc257dc86};
test_output[23216:23223] = '{32'h0, 32'h0, 32'h0, 32'h42c7718a, 32'h429ea4b0, 32'h41f1edfb, 32'h0, 32'h0};
test_input[23224:23231] = '{32'h411922ea, 32'hc217be30, 32'hc2b48224, 32'h42861346, 32'hc2afec30, 32'h42240e16, 32'hc2938e22, 32'hc23a15c6};
test_output[23224:23231] = '{32'h411922ea, 32'h0, 32'h0, 32'h42861346, 32'h0, 32'h42240e16, 32'h0, 32'h0};
test_input[23232:23239] = '{32'h4228517a, 32'h418f635a, 32'hc2b558b6, 32'h412616ec, 32'hc12ca40c, 32'h4209fb29, 32'hc2891d60, 32'hc1d997d6};
test_output[23232:23239] = '{32'h4228517a, 32'h418f635a, 32'h0, 32'h412616ec, 32'h0, 32'h4209fb29, 32'h0, 32'h0};
test_input[23240:23247] = '{32'hc2aa04f3, 32'h420bc9f5, 32'h428c7c1a, 32'hc28cef9d, 32'hc1ac97e4, 32'h4203181a, 32'hc1ac20fa, 32'h413ceb8f};
test_output[23240:23247] = '{32'h0, 32'h420bc9f5, 32'h428c7c1a, 32'h0, 32'h0, 32'h4203181a, 32'h0, 32'h413ceb8f};
test_input[23248:23255] = '{32'hc233bf60, 32'h42731225, 32'hc0367b44, 32'hc29c26d3, 32'hc23025e2, 32'hc1074bd5, 32'h422f1f3d, 32'h42c22280};
test_output[23248:23255] = '{32'h0, 32'h42731225, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422f1f3d, 32'h42c22280};
test_input[23256:23263] = '{32'hc2529d56, 32'hc282e194, 32'h42b91bf4, 32'hc235e7a0, 32'h4295a5e7, 32'h4297b202, 32'h41e6a145, 32'hc260ca2d};
test_output[23256:23263] = '{32'h0, 32'h0, 32'h42b91bf4, 32'h0, 32'h4295a5e7, 32'h4297b202, 32'h41e6a145, 32'h0};
test_input[23264:23271] = '{32'h40429b41, 32'hc128eaa4, 32'hbf92e5a8, 32'hc272c5fd, 32'hc2b3cd1e, 32'h42a3646e, 32'hc2b49e08, 32'hbedbbae3};
test_output[23264:23271] = '{32'h40429b41, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a3646e, 32'h0, 32'h0};
test_input[23272:23279] = '{32'hc296bcd6, 32'h41e014ff, 32'h42c309e7, 32'hc2bc2e21, 32'h42b704cb, 32'hc2b2d053, 32'h41f687c0, 32'h42a120e2};
test_output[23272:23279] = '{32'h0, 32'h41e014ff, 32'h42c309e7, 32'h0, 32'h42b704cb, 32'h0, 32'h41f687c0, 32'h42a120e2};
test_input[23280:23287] = '{32'h42a2a091, 32'hc08c83ab, 32'hc263a582, 32'hc16e154d, 32'hbe9dc0e3, 32'hc2bb6234, 32'h429993c1, 32'hc1e03a9f};
test_output[23280:23287] = '{32'h42a2a091, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429993c1, 32'h0};
test_input[23288:23295] = '{32'h42bc45f0, 32'h42677f8c, 32'h40bf848f, 32'hc1c859b5, 32'h429671fd, 32'h4137822c, 32'hc2800fc2, 32'h425e90a1};
test_output[23288:23295] = '{32'h42bc45f0, 32'h42677f8c, 32'h40bf848f, 32'h0, 32'h429671fd, 32'h4137822c, 32'h0, 32'h425e90a1};
test_input[23296:23303] = '{32'hc2c072b9, 32'hc1d71567, 32'h420d07ac, 32'h4271f97d, 32'hc2ab9c19, 32'h42b33e08, 32'h40ea7497, 32'h424ca586};
test_output[23296:23303] = '{32'h0, 32'h0, 32'h420d07ac, 32'h4271f97d, 32'h0, 32'h42b33e08, 32'h40ea7497, 32'h424ca586};
test_input[23304:23311] = '{32'hc18e9138, 32'h426f3848, 32'h41bf4fe9, 32'h403c316c, 32'h4208bd16, 32'hc2b8ce59, 32'hc24eb026, 32'h42baa290};
test_output[23304:23311] = '{32'h0, 32'h426f3848, 32'h41bf4fe9, 32'h403c316c, 32'h4208bd16, 32'h0, 32'h0, 32'h42baa290};
test_input[23312:23319] = '{32'hc2a1851d, 32'h42814cff, 32'hc10fcc0b, 32'hc2b01f44, 32'hc296557b, 32'h418a3d33, 32'hc2b2d7e3, 32'hc1b73fe6};
test_output[23312:23319] = '{32'h0, 32'h42814cff, 32'h0, 32'h0, 32'h0, 32'h418a3d33, 32'h0, 32'h0};
test_input[23320:23327] = '{32'h428c6043, 32'hc1f30b60, 32'h42bebe38, 32'hc2914c67, 32'hc2b6b0c6, 32'hc2003ecc, 32'hc2add075, 32'hc2bf7631};
test_output[23320:23327] = '{32'h428c6043, 32'h0, 32'h42bebe38, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23328:23335] = '{32'hc1d85746, 32'h4137c841, 32'hc2727fe7, 32'hc25e92b7, 32'h42b19c27, 32'h42ac89c8, 32'h41d804f5, 32'hc2b9ad3f};
test_output[23328:23335] = '{32'h0, 32'h4137c841, 32'h0, 32'h0, 32'h42b19c27, 32'h42ac89c8, 32'h41d804f5, 32'h0};
test_input[23336:23343] = '{32'h41fce3dd, 32'h4123bd04, 32'h42417d75, 32'hc1f442df, 32'h423b99b9, 32'hc1816dfa, 32'h42a75918, 32'h421f42c7};
test_output[23336:23343] = '{32'h41fce3dd, 32'h4123bd04, 32'h42417d75, 32'h0, 32'h423b99b9, 32'h0, 32'h42a75918, 32'h421f42c7};
test_input[23344:23351] = '{32'hc268d959, 32'hc28c2cb3, 32'h409af5b4, 32'hc28311a3, 32'h420eceac, 32'hc1ed902f, 32'hc2a2b2b4, 32'hc2aef0a5};
test_output[23344:23351] = '{32'h0, 32'h0, 32'h409af5b4, 32'h0, 32'h420eceac, 32'h0, 32'h0, 32'h0};
test_input[23352:23359] = '{32'hc1a44861, 32'hc29d5671, 32'h42bfe751, 32'hc24c4b8d, 32'hc24d59de, 32'hc0c7c9a2, 32'h41d16ade, 32'hc2c42117};
test_output[23352:23359] = '{32'h0, 32'h0, 32'h42bfe751, 32'h0, 32'h0, 32'h0, 32'h41d16ade, 32'h0};
test_input[23360:23367] = '{32'h425e223c, 32'hc2ae3d98, 32'hc21a1a20, 32'h426d5667, 32'hc146eff5, 32'h415fb48c, 32'hc2777b90, 32'h426da096};
test_output[23360:23367] = '{32'h425e223c, 32'h0, 32'h0, 32'h426d5667, 32'h0, 32'h415fb48c, 32'h0, 32'h426da096};
test_input[23368:23375] = '{32'hc1bf9b93, 32'h41fa3672, 32'hc0d33037, 32'h4236c9de, 32'h42a5943a, 32'hc1ea19b4, 32'h41b7c296, 32'hc29b8b8d};
test_output[23368:23375] = '{32'h0, 32'h41fa3672, 32'h0, 32'h4236c9de, 32'h42a5943a, 32'h0, 32'h41b7c296, 32'h0};
test_input[23376:23383] = '{32'h42995152, 32'h42b15142, 32'hc29321fc, 32'h428dcd36, 32'h41b162f1, 32'hc14487ed, 32'hc18d07c8, 32'hc287ce36};
test_output[23376:23383] = '{32'h42995152, 32'h42b15142, 32'h0, 32'h428dcd36, 32'h41b162f1, 32'h0, 32'h0, 32'h0};
test_input[23384:23391] = '{32'hc273be7e, 32'h4256f527, 32'hc22d962d, 32'hc195ba5e, 32'hc16c8eb6, 32'hc24634bb, 32'hc1acd619, 32'hc252469c};
test_output[23384:23391] = '{32'h0, 32'h4256f527, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23392:23399] = '{32'hc2564178, 32'hc2172688, 32'h3f77ea8f, 32'hc278ad42, 32'hc2a22cca, 32'hc21a2b6c, 32'hc29c2350, 32'h4256c53e};
test_output[23392:23399] = '{32'h0, 32'h0, 32'h3f77ea8f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4256c53e};
test_input[23400:23407] = '{32'hc287b576, 32'h4241d1f5, 32'hc1b93a5f, 32'h42be83f2, 32'hc1f7cbec, 32'h4263d499, 32'hc29156df, 32'hc278a86f};
test_output[23400:23407] = '{32'h0, 32'h4241d1f5, 32'h0, 32'h42be83f2, 32'h0, 32'h4263d499, 32'h0, 32'h0};
test_input[23408:23415] = '{32'hc1b078c0, 32'h428494fd, 32'h421cefef, 32'h41ba3099, 32'h42bbb5d1, 32'h4200c1b4, 32'h42323ff7, 32'hc27fb3a5};
test_output[23408:23415] = '{32'h0, 32'h428494fd, 32'h421cefef, 32'h41ba3099, 32'h42bbb5d1, 32'h4200c1b4, 32'h42323ff7, 32'h0};
test_input[23416:23423] = '{32'h42b1ff8a, 32'h4100741b, 32'h421b4bc5, 32'hc161d5ca, 32'hc1a9fc6a, 32'hc293b944, 32'h426ad98b, 32'h41b92d47};
test_output[23416:23423] = '{32'h42b1ff8a, 32'h4100741b, 32'h421b4bc5, 32'h0, 32'h0, 32'h0, 32'h426ad98b, 32'h41b92d47};
test_input[23424:23431] = '{32'hc1a101df, 32'h42c0e4e5, 32'hc2055792, 32'hc2988375, 32'hc251a663, 32'h421345d6, 32'hc213b7dc, 32'h42b2b844};
test_output[23424:23431] = '{32'h0, 32'h42c0e4e5, 32'h0, 32'h0, 32'h0, 32'h421345d6, 32'h0, 32'h42b2b844};
test_input[23432:23439] = '{32'h429a178e, 32'h41e205ca, 32'h4241d82b, 32'hc2b37eed, 32'hc2c63ffa, 32'hc2870de0, 32'hc14c4732, 32'hc190fed3};
test_output[23432:23439] = '{32'h429a178e, 32'h41e205ca, 32'h4241d82b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23440:23447] = '{32'h4297ffee, 32'h4266fcc4, 32'h42498ada, 32'hc21032b1, 32'h42c4e82a, 32'h42735ad2, 32'hc2b5dee5, 32'hc2aa648a};
test_output[23440:23447] = '{32'h4297ffee, 32'h4266fcc4, 32'h42498ada, 32'h0, 32'h42c4e82a, 32'h42735ad2, 32'h0, 32'h0};
test_input[23448:23455] = '{32'h421bb2e2, 32'h416c89d5, 32'hc2159da6, 32'hc2b146ec, 32'h41cef8e4, 32'hc29b5afc, 32'h411be645, 32'h421f2e4c};
test_output[23448:23455] = '{32'h421bb2e2, 32'h416c89d5, 32'h0, 32'h0, 32'h41cef8e4, 32'h0, 32'h411be645, 32'h421f2e4c};
test_input[23456:23463] = '{32'hc18af919, 32'hc29d5c67, 32'h420ee69e, 32'hc2af11f6, 32'h3fb3dd56, 32'h4288e0a5, 32'h42801ff4, 32'hc18f7cf1};
test_output[23456:23463] = '{32'h0, 32'h0, 32'h420ee69e, 32'h0, 32'h3fb3dd56, 32'h4288e0a5, 32'h42801ff4, 32'h0};
test_input[23464:23471] = '{32'h41b6800c, 32'hc0188585, 32'hc2998d23, 32'hc290b9a8, 32'hc2b3cc39, 32'hc2ae6d6a, 32'h412fc9f3, 32'hc279865a};
test_output[23464:23471] = '{32'h41b6800c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h412fc9f3, 32'h0};
test_input[23472:23479] = '{32'hc2b673b3, 32'h425dea21, 32'hc14bf312, 32'hc26ca10f, 32'hc1bc8e9f, 32'h42b34161, 32'hc23b5436, 32'hc1785109};
test_output[23472:23479] = '{32'h0, 32'h425dea21, 32'h0, 32'h0, 32'h0, 32'h42b34161, 32'h0, 32'h0};
test_input[23480:23487] = '{32'h413621d5, 32'h4222399e, 32'hc2a089ff, 32'h42ac5882, 32'h418a378e, 32'h42a3a7ff, 32'h42badc6d, 32'h42575481};
test_output[23480:23487] = '{32'h413621d5, 32'h4222399e, 32'h0, 32'h42ac5882, 32'h418a378e, 32'h42a3a7ff, 32'h42badc6d, 32'h42575481};
test_input[23488:23495] = '{32'h420c48f1, 32'hc2abb063, 32'h427a8d1b, 32'hc2bbe87e, 32'h3f91b14f, 32'hc09cb5a1, 32'h41ad02b8, 32'h4123b694};
test_output[23488:23495] = '{32'h420c48f1, 32'h0, 32'h427a8d1b, 32'h0, 32'h3f91b14f, 32'h0, 32'h41ad02b8, 32'h4123b694};
test_input[23496:23503] = '{32'hc101d4bf, 32'hc1acef67, 32'h42994f44, 32'h42b52d3f, 32'h42bf2250, 32'h42b0b5e3, 32'h4124997d, 32'h41e54422};
test_output[23496:23503] = '{32'h0, 32'h0, 32'h42994f44, 32'h42b52d3f, 32'h42bf2250, 32'h42b0b5e3, 32'h4124997d, 32'h41e54422};
test_input[23504:23511] = '{32'hc213e36f, 32'hc2b20fc1, 32'hc262b599, 32'hc15b42bc, 32'h420cd6fa, 32'h4288c7f8, 32'hc247029c, 32'h4207cc18};
test_output[23504:23511] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h420cd6fa, 32'h4288c7f8, 32'h0, 32'h4207cc18};
test_input[23512:23519] = '{32'hc2c155f2, 32'hc2a078d6, 32'h419413b7, 32'hc22e5655, 32'hc11f446c, 32'h42a51fad, 32'hc2026221, 32'h42b94869};
test_output[23512:23519] = '{32'h0, 32'h0, 32'h419413b7, 32'h0, 32'h0, 32'h42a51fad, 32'h0, 32'h42b94869};
test_input[23520:23527] = '{32'h42a5aca5, 32'h41fd6c25, 32'h42640834, 32'h41ae703f, 32'h411db90e, 32'h419e3726, 32'hc1b59397, 32'hc28b728c};
test_output[23520:23527] = '{32'h42a5aca5, 32'h41fd6c25, 32'h42640834, 32'h41ae703f, 32'h411db90e, 32'h419e3726, 32'h0, 32'h0};
test_input[23528:23535] = '{32'h42b75cc0, 32'h427c09ee, 32'h428380b8, 32'hc27430bd, 32'hc27719ca, 32'hc28463d6, 32'hc2afa94f, 32'hc215925d};
test_output[23528:23535] = '{32'h42b75cc0, 32'h427c09ee, 32'h428380b8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23536:23543] = '{32'h41425a6d, 32'h429de151, 32'h412bc75a, 32'h42786864, 32'hc2251f72, 32'hc23b75a8, 32'hc2a56e6d, 32'hc1e3ec70};
test_output[23536:23543] = '{32'h41425a6d, 32'h429de151, 32'h412bc75a, 32'h42786864, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23544:23551] = '{32'hc2b3c457, 32'h42ae9c7d, 32'hc26a8b19, 32'hc1ca10c2, 32'hc2a9e5be, 32'h42b4ed59, 32'h4210b56c, 32'h42a26955};
test_output[23544:23551] = '{32'h0, 32'h42ae9c7d, 32'h0, 32'h0, 32'h0, 32'h42b4ed59, 32'h4210b56c, 32'h42a26955};
test_input[23552:23559] = '{32'h42768bec, 32'h41edecc6, 32'h42a4193a, 32'h422169ed, 32'hc283e8c6, 32'hc2b52c99, 32'h4235edd4, 32'h42b43e39};
test_output[23552:23559] = '{32'h42768bec, 32'h41edecc6, 32'h42a4193a, 32'h422169ed, 32'h0, 32'h0, 32'h4235edd4, 32'h42b43e39};
test_input[23560:23567] = '{32'hc2abdb14, 32'hc249810f, 32'hc21a7323, 32'hc2b64e03, 32'hc28f4ba1, 32'hc2bcb23f, 32'h42821d41, 32'hc21d7af8};
test_output[23560:23567] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42821d41, 32'h0};
test_input[23568:23575] = '{32'h42b4f78d, 32'hc1a7176a, 32'h42b18a44, 32'hc12424d4, 32'hc2c2c42b, 32'hc288fa55, 32'h424946c6, 32'h423d429a};
test_output[23568:23575] = '{32'h42b4f78d, 32'h0, 32'h42b18a44, 32'h0, 32'h0, 32'h0, 32'h424946c6, 32'h423d429a};
test_input[23576:23583] = '{32'h3fd2a4b8, 32'h40d74f4f, 32'hc22f8b71, 32'h421367e8, 32'hc26e5d43, 32'h41911363, 32'h4202340d, 32'hc2c5fdf9};
test_output[23576:23583] = '{32'h3fd2a4b8, 32'h40d74f4f, 32'h0, 32'h421367e8, 32'h0, 32'h41911363, 32'h4202340d, 32'h0};
test_input[23584:23591] = '{32'h42c725e7, 32'h4283d3b7, 32'h42bb7844, 32'hc18a54a7, 32'h428624da, 32'h426695a2, 32'h3f865277, 32'h42331c60};
test_output[23584:23591] = '{32'h42c725e7, 32'h4283d3b7, 32'h42bb7844, 32'h0, 32'h428624da, 32'h426695a2, 32'h3f865277, 32'h42331c60};
test_input[23592:23599] = '{32'hc2622786, 32'h42728549, 32'h429f2a59, 32'h422b8cb9, 32'h42271f76, 32'h422a8387, 32'hc288b984, 32'h4254f613};
test_output[23592:23599] = '{32'h0, 32'h42728549, 32'h429f2a59, 32'h422b8cb9, 32'h42271f76, 32'h422a8387, 32'h0, 32'h4254f613};
test_input[23600:23607] = '{32'h421f4e8b, 32'h409eab54, 32'hc2b9fbd8, 32'hc2488430, 32'hc286693b, 32'hbffd5c85, 32'hc2c3650b, 32'hc0cc64d9};
test_output[23600:23607] = '{32'h421f4e8b, 32'h409eab54, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23608:23615] = '{32'hc212d933, 32'h42bd348f, 32'hc1d10094, 32'h3fd56982, 32'h4292daa8, 32'h400e8008, 32'hc2bbf7d7, 32'h42512205};
test_output[23608:23615] = '{32'h0, 32'h42bd348f, 32'h0, 32'h3fd56982, 32'h4292daa8, 32'h400e8008, 32'h0, 32'h42512205};
test_input[23616:23623] = '{32'hc2627188, 32'h428a6a54, 32'hc2c52cef, 32'h42bb62dd, 32'hc294734f, 32'hc29a39af, 32'hc1c644ab, 32'hc2242061};
test_output[23616:23623] = '{32'h0, 32'h428a6a54, 32'h0, 32'h42bb62dd, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23624:23631] = '{32'hc139d134, 32'h415b4412, 32'h42854ed3, 32'h419fb92d, 32'hc2b026c4, 32'hc2c5a35b, 32'h42ab92b1, 32'hc2977172};
test_output[23624:23631] = '{32'h0, 32'h415b4412, 32'h42854ed3, 32'h419fb92d, 32'h0, 32'h0, 32'h42ab92b1, 32'h0};
test_input[23632:23639] = '{32'hc298f868, 32'h41040f2c, 32'hc0a35074, 32'h4192039b, 32'h42c21d71, 32'hc2c69243, 32'h4200ffb2, 32'h42af97a1};
test_output[23632:23639] = '{32'h0, 32'h41040f2c, 32'h0, 32'h4192039b, 32'h42c21d71, 32'h0, 32'h4200ffb2, 32'h42af97a1};
test_input[23640:23647] = '{32'h427b7446, 32'hc1aa5efa, 32'h41dd8381, 32'hc27bbd59, 32'hc292f755, 32'h40619ede, 32'hc226a2ff, 32'h41d75478};
test_output[23640:23647] = '{32'h427b7446, 32'h0, 32'h41dd8381, 32'h0, 32'h0, 32'h40619ede, 32'h0, 32'h41d75478};
test_input[23648:23655] = '{32'hc2b5c5d3, 32'h4227c718, 32'hc2c61bc9, 32'hc2b9c595, 32'h40e83151, 32'hc1a1b306, 32'hc29eb77c, 32'h42c425c4};
test_output[23648:23655] = '{32'h0, 32'h4227c718, 32'h0, 32'h0, 32'h40e83151, 32'h0, 32'h0, 32'h42c425c4};
test_input[23656:23663] = '{32'hc259f6a1, 32'hc2a01a8b, 32'hc2c1b023, 32'h427d5c56, 32'hc2b62357, 32'h40747053, 32'hc2c6115b, 32'hc2b7346d};
test_output[23656:23663] = '{32'h0, 32'h0, 32'h0, 32'h427d5c56, 32'h0, 32'h40747053, 32'h0, 32'h0};
test_input[23664:23671] = '{32'h423fc2e1, 32'hc2a075ad, 32'h416e7f6a, 32'hc22ed75e, 32'h4007c360, 32'h425812fb, 32'hc2493afc, 32'h41378df7};
test_output[23664:23671] = '{32'h423fc2e1, 32'h0, 32'h416e7f6a, 32'h0, 32'h4007c360, 32'h425812fb, 32'h0, 32'h41378df7};
test_input[23672:23679] = '{32'h4220530d, 32'hc1a42669, 32'hc24e6826, 32'hc290b041, 32'hc2c0843e, 32'h4250d036, 32'h4249a705, 32'h420c316a};
test_output[23672:23679] = '{32'h4220530d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4250d036, 32'h4249a705, 32'h420c316a};
test_input[23680:23687] = '{32'h421266ee, 32'h429ffb99, 32'hc1884226, 32'h422fe7e7, 32'hc2bbdda2, 32'hc24e3d62, 32'hc29f4cba, 32'hc26d5a4e};
test_output[23680:23687] = '{32'h421266ee, 32'h429ffb99, 32'h0, 32'h422fe7e7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23688:23695] = '{32'h421d024c, 32'hc1afbd5f, 32'h427b2dad, 32'hc2a1e7b3, 32'hc2bc39cc, 32'h42819393, 32'h410971cc, 32'h42804396};
test_output[23688:23695] = '{32'h421d024c, 32'h0, 32'h427b2dad, 32'h0, 32'h0, 32'h42819393, 32'h410971cc, 32'h42804396};
test_input[23696:23703] = '{32'h423ecdc6, 32'h40d790b3, 32'h419e71be, 32'h42bf6d39, 32'hc100ff9c, 32'h428a9f6b, 32'hc23a0a33, 32'hc23f224d};
test_output[23696:23703] = '{32'h423ecdc6, 32'h40d790b3, 32'h419e71be, 32'h42bf6d39, 32'h0, 32'h428a9f6b, 32'h0, 32'h0};
test_input[23704:23711] = '{32'hc1cd1a63, 32'hc1eed681, 32'h42c38f24, 32'hc28c3662, 32'h42be346b, 32'hc2564b48, 32'hc10a0fd5, 32'hc2a13d88};
test_output[23704:23711] = '{32'h0, 32'h0, 32'h42c38f24, 32'h0, 32'h42be346b, 32'h0, 32'h0, 32'h0};
test_input[23712:23719] = '{32'hc27cf3c7, 32'h425b43a2, 32'h4270a122, 32'hc246a976, 32'hc2b8dce4, 32'hc2815063, 32'hc2bf2602, 32'h3f97556f};
test_output[23712:23719] = '{32'h0, 32'h425b43a2, 32'h4270a122, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3f97556f};
test_input[23720:23727] = '{32'h42b025bf, 32'hc2af4e3c, 32'h42ae4356, 32'hc1aae012, 32'hc275fb1d, 32'h427abd0a, 32'hc1ceef9d, 32'h41c510c7};
test_output[23720:23727] = '{32'h42b025bf, 32'h0, 32'h42ae4356, 32'h0, 32'h0, 32'h427abd0a, 32'h0, 32'h41c510c7};
test_input[23728:23735] = '{32'h41fbeead, 32'h426bc515, 32'hc127d073, 32'hc23c55c5, 32'h412202f9, 32'h4288a96b, 32'hc234769a, 32'hc2354b2a};
test_output[23728:23735] = '{32'h41fbeead, 32'h426bc515, 32'h0, 32'h0, 32'h412202f9, 32'h4288a96b, 32'h0, 32'h0};
test_input[23736:23743] = '{32'hc28bf748, 32'h42ab6459, 32'h42aa07f9, 32'hc1b83cde, 32'hc270fb69, 32'h4254b59b, 32'h412f3a41, 32'hc12d2976};
test_output[23736:23743] = '{32'h0, 32'h42ab6459, 32'h42aa07f9, 32'h0, 32'h0, 32'h4254b59b, 32'h412f3a41, 32'h0};
test_input[23744:23751] = '{32'hc2267fc6, 32'hc21660b4, 32'h42c17404, 32'hc252dfc4, 32'h4119b4c9, 32'hc27bba0e, 32'hc1e0b0bc, 32'h42a8f33a};
test_output[23744:23751] = '{32'h0, 32'h0, 32'h42c17404, 32'h0, 32'h4119b4c9, 32'h0, 32'h0, 32'h42a8f33a};
test_input[23752:23759] = '{32'h42a7fdf6, 32'hc25a8afb, 32'h42974907, 32'h42734fc4, 32'h4244e253, 32'hc2baf5c4, 32'hc26926d7, 32'h428d16c3};
test_output[23752:23759] = '{32'h42a7fdf6, 32'h0, 32'h42974907, 32'h42734fc4, 32'h4244e253, 32'h0, 32'h0, 32'h428d16c3};
test_input[23760:23767] = '{32'hc281ddb9, 32'h42692995, 32'hc2a1eb4f, 32'hc28df6b8, 32'hc1a10599, 32'h41bffcd9, 32'h41e4f9a3, 32'h42a84dbb};
test_output[23760:23767] = '{32'h0, 32'h42692995, 32'h0, 32'h0, 32'h0, 32'h41bffcd9, 32'h41e4f9a3, 32'h42a84dbb};
test_input[23768:23775] = '{32'hc281e6c2, 32'hc2a75458, 32'h4286503f, 32'hc246b96e, 32'hc2653203, 32'hc22facc8, 32'h422d003b, 32'hc1f651aa};
test_output[23768:23775] = '{32'h0, 32'h0, 32'h4286503f, 32'h0, 32'h0, 32'h0, 32'h422d003b, 32'h0};
test_input[23776:23783] = '{32'hc29a5972, 32'hc241aba5, 32'hc25c5f18, 32'hc2ad14a1, 32'hc12cfb6b, 32'hc2894001, 32'hc01bf948, 32'hc265ede1};
test_output[23776:23783] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23784:23791] = '{32'h424e1e0b, 32'h42816cee, 32'h426cd367, 32'hc1de71f3, 32'h4151f928, 32'h42b626fb, 32'h429a741d, 32'h42159279};
test_output[23784:23791] = '{32'h424e1e0b, 32'h42816cee, 32'h426cd367, 32'h0, 32'h4151f928, 32'h42b626fb, 32'h429a741d, 32'h42159279};
test_input[23792:23799] = '{32'h423f4fba, 32'h41b34685, 32'h423983e0, 32'h429f7ae8, 32'hc2779802, 32'hc2215d21, 32'hc2a80c24, 32'hc29d5323};
test_output[23792:23799] = '{32'h423f4fba, 32'h41b34685, 32'h423983e0, 32'h429f7ae8, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23800:23807] = '{32'h42bbd367, 32'hc2116d5b, 32'h42baccf7, 32'hc19e8c12, 32'hc2233136, 32'h41f8057b, 32'hc201178b, 32'h422b2ebe};
test_output[23800:23807] = '{32'h42bbd367, 32'h0, 32'h42baccf7, 32'h0, 32'h0, 32'h41f8057b, 32'h0, 32'h422b2ebe};
test_input[23808:23815] = '{32'hc1249fdb, 32'hc1d3feae, 32'hc2b7c658, 32'h428ceb98, 32'hc2b61e30, 32'hc2087d4d, 32'hc2b3bdc7, 32'hc2b3d282};
test_output[23808:23815] = '{32'h0, 32'h0, 32'h0, 32'h428ceb98, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[23816:23823] = '{32'hc23e66bb, 32'h41a224fd, 32'hc0a77421, 32'h429f2a7d, 32'h4174d85f, 32'h429c002a, 32'h4205006c, 32'h4115821a};
test_output[23816:23823] = '{32'h0, 32'h41a224fd, 32'h0, 32'h429f2a7d, 32'h4174d85f, 32'h429c002a, 32'h4205006c, 32'h4115821a};
test_input[23824:23831] = '{32'h42beae36, 32'hbf577129, 32'hc1c83fa2, 32'hc0ba4291, 32'h41a48fd6, 32'hc0dc28d2, 32'h42939b16, 32'h42a5e54e};
test_output[23824:23831] = '{32'h42beae36, 32'h0, 32'h0, 32'h0, 32'h41a48fd6, 32'h0, 32'h42939b16, 32'h42a5e54e};
test_input[23832:23839] = '{32'h42bcb63c, 32'hc02b3536, 32'h4251ed7c, 32'hc2a88773, 32'h41926881, 32'h42837987, 32'hc27eb36d, 32'h421f2d75};
test_output[23832:23839] = '{32'h42bcb63c, 32'h0, 32'h4251ed7c, 32'h0, 32'h41926881, 32'h42837987, 32'h0, 32'h421f2d75};
test_input[23840:23847] = '{32'h3fcd5045, 32'hc23afdbe, 32'h42a5b402, 32'hc19708d9, 32'h42bc5346, 32'h42bf4a33, 32'hc2980ff3, 32'hc1b9f4e5};
test_output[23840:23847] = '{32'h3fcd5045, 32'h0, 32'h42a5b402, 32'h0, 32'h42bc5346, 32'h42bf4a33, 32'h0, 32'h0};
test_input[23848:23855] = '{32'h41d54386, 32'hc2988fd1, 32'hc2a2d3c6, 32'h42c0f08d, 32'h421dba41, 32'h4233e46a, 32'hc2c51ff2, 32'hc259ff61};
test_output[23848:23855] = '{32'h41d54386, 32'h0, 32'h0, 32'h42c0f08d, 32'h421dba41, 32'h4233e46a, 32'h0, 32'h0};
test_input[23856:23863] = '{32'hc120be2d, 32'hc1c06ec9, 32'hc2641ae1, 32'hc243e11b, 32'h41ea08b6, 32'hc23f2b30, 32'h41b24975, 32'hbf341cf2};
test_output[23856:23863] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41ea08b6, 32'h0, 32'h41b24975, 32'h0};
test_input[23864:23871] = '{32'hc243b9a7, 32'hc0a4e14e, 32'h4211cc75, 32'h4290a383, 32'h4190d8c6, 32'h4251c45e, 32'h42b6417f, 32'h4141f9e5};
test_output[23864:23871] = '{32'h0, 32'h0, 32'h4211cc75, 32'h4290a383, 32'h4190d8c6, 32'h4251c45e, 32'h42b6417f, 32'h4141f9e5};
test_input[23872:23879] = '{32'hc0380743, 32'hc196b772, 32'hc28b4ebf, 32'hc2073c69, 32'h429c1b69, 32'h42204bea, 32'h424e12b1, 32'h425c05c7};
test_output[23872:23879] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429c1b69, 32'h42204bea, 32'h424e12b1, 32'h425c05c7};
test_input[23880:23887] = '{32'h40403a27, 32'hc228609a, 32'h4082ac71, 32'h41a5e9fb, 32'hc12ff763, 32'hc2af5a74, 32'h42b8fab8, 32'hc166e70c};
test_output[23880:23887] = '{32'h40403a27, 32'h0, 32'h4082ac71, 32'h41a5e9fb, 32'h0, 32'h0, 32'h42b8fab8, 32'h0};
test_input[23888:23895] = '{32'hc1babc95, 32'hc29432bb, 32'hc278f1ca, 32'hc29ae9d3, 32'hc2b897c6, 32'h4212e2b4, 32'h421a6bd6, 32'hc235b269};
test_output[23888:23895] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4212e2b4, 32'h421a6bd6, 32'h0};
test_input[23896:23903] = '{32'h42c709ff, 32'h42527e35, 32'hc19edbd8, 32'hbfb636a7, 32'h4191c0a2, 32'h3fe8510f, 32'hc0fe7edb, 32'h427bef55};
test_output[23896:23903] = '{32'h42c709ff, 32'h42527e35, 32'h0, 32'h0, 32'h4191c0a2, 32'h3fe8510f, 32'h0, 32'h427bef55};
test_input[23904:23911] = '{32'h424012e1, 32'hc25db47e, 32'hc25db8f7, 32'hc2927ccd, 32'hc235e749, 32'hc23d22bd, 32'hc2393e10, 32'h41e0278c};
test_output[23904:23911] = '{32'h424012e1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41e0278c};
test_input[23912:23919] = '{32'hc1e27069, 32'hc18c6c4b, 32'hc0f5915e, 32'h4210d1bf, 32'h42c0600f, 32'h42abc2c3, 32'hc21e2cb9, 32'h420bd63c};
test_output[23912:23919] = '{32'h0, 32'h0, 32'h0, 32'h4210d1bf, 32'h42c0600f, 32'h42abc2c3, 32'h0, 32'h420bd63c};
test_input[23920:23927] = '{32'hc283476f, 32'hc2a1b0c0, 32'h42b4a9e3, 32'hc2c1a488, 32'hc2560588, 32'h4115ea30, 32'h42868764, 32'h4284333e};
test_output[23920:23927] = '{32'h0, 32'h0, 32'h42b4a9e3, 32'h0, 32'h0, 32'h4115ea30, 32'h42868764, 32'h4284333e};
test_input[23928:23935] = '{32'hc1efe344, 32'hc2bb989c, 32'hc28a5e0c, 32'hc1f59417, 32'h42b2d5bd, 32'h42afa45a, 32'hc1887294, 32'h426be53b};
test_output[23928:23935] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42b2d5bd, 32'h42afa45a, 32'h0, 32'h426be53b};
test_input[23936:23943] = '{32'h428c83a0, 32'h42a0f738, 32'hc2b7bf8f, 32'h42935b14, 32'h42c5f8a9, 32'hc2b950c4, 32'h40cb7692, 32'hc22c4d0d};
test_output[23936:23943] = '{32'h428c83a0, 32'h42a0f738, 32'h0, 32'h42935b14, 32'h42c5f8a9, 32'h0, 32'h40cb7692, 32'h0};
test_input[23944:23951] = '{32'hc16c0285, 32'h4292be75, 32'hc0c7a57c, 32'hc16fdc5f, 32'hc1ff8adc, 32'hc24dc289, 32'hc1ee5408, 32'h41d28a4d};
test_output[23944:23951] = '{32'h0, 32'h4292be75, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41d28a4d};
test_input[23952:23959] = '{32'h40d8ec70, 32'hc1746d1c, 32'hc1a88493, 32'h422685c9, 32'hc240b6dd, 32'h42106b54, 32'hc29df856, 32'h41c945f9};
test_output[23952:23959] = '{32'h40d8ec70, 32'h0, 32'h0, 32'h422685c9, 32'h0, 32'h42106b54, 32'h0, 32'h41c945f9};
test_input[23960:23967] = '{32'h42b6b808, 32'h428a86c0, 32'h42a57d51, 32'h4202f7b4, 32'h41f8199f, 32'hc1513089, 32'hc202a5a5, 32'hc1c14fe3};
test_output[23960:23967] = '{32'h42b6b808, 32'h428a86c0, 32'h42a57d51, 32'h4202f7b4, 32'h41f8199f, 32'h0, 32'h0, 32'h0};
test_input[23968:23975] = '{32'h429d423b, 32'hc00e703a, 32'hc28bed78, 32'hc16375e6, 32'hc12302fd, 32'hc06bba37, 32'h422592b7, 32'hc2a600fe};
test_output[23968:23975] = '{32'h429d423b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422592b7, 32'h0};
test_input[23976:23983] = '{32'h41bb73d3, 32'hc2a9e652, 32'hc19802d0, 32'h42939344, 32'hc128d0f8, 32'h42504d84, 32'h423a9b20, 32'h41683682};
test_output[23976:23983] = '{32'h41bb73d3, 32'h0, 32'h0, 32'h42939344, 32'h0, 32'h42504d84, 32'h423a9b20, 32'h41683682};
test_input[23984:23991] = '{32'hc2445c44, 32'h42bc9b74, 32'h42079ebb, 32'h42032ec4, 32'hc1337780, 32'hc0f0ba4f, 32'hc2b2c225, 32'h42c37486};
test_output[23984:23991] = '{32'h0, 32'h42bc9b74, 32'h42079ebb, 32'h42032ec4, 32'h0, 32'h0, 32'h0, 32'h42c37486};
test_input[23992:23999] = '{32'h41e23850, 32'hc15a3781, 32'h406d28c4, 32'hc22f7701, 32'hc21743cb, 32'hc0830809, 32'h427ff1d1, 32'h42525afa};
test_output[23992:23999] = '{32'h41e23850, 32'h0, 32'h406d28c4, 32'h0, 32'h0, 32'h0, 32'h427ff1d1, 32'h42525afa};
test_input[24000:24007] = '{32'hc2744957, 32'hc2447a92, 32'hc23e38e4, 32'h4281ea7a, 32'h42b7c41e, 32'hc24dd12a, 32'hc2ad8f14, 32'hc232407d};
test_output[24000:24007] = '{32'h0, 32'h0, 32'h0, 32'h4281ea7a, 32'h42b7c41e, 32'h0, 32'h0, 32'h0};
test_input[24008:24015] = '{32'hc1854585, 32'hc28c5302, 32'hc26e0da8, 32'h415f88a2, 32'hc2ae4418, 32'h423a2a64, 32'h429a22b7, 32'h429c6bd5};
test_output[24008:24015] = '{32'h0, 32'h0, 32'h0, 32'h415f88a2, 32'h0, 32'h423a2a64, 32'h429a22b7, 32'h429c6bd5};
test_input[24016:24023] = '{32'h3e8bc844, 32'hc2b1ac93, 32'hc2bab720, 32'hc20136d2, 32'h413436b5, 32'hc1878b4a, 32'h42108e71, 32'h4122a3fc};
test_output[24016:24023] = '{32'h3e8bc844, 32'h0, 32'h0, 32'h0, 32'h413436b5, 32'h0, 32'h42108e71, 32'h4122a3fc};
test_input[24024:24031] = '{32'hc289ca59, 32'hc28120e0, 32'hc190e2ba, 32'h42a9d6d2, 32'h40653373, 32'hc1dd0862, 32'hc240c5ed, 32'hc0ea2896};
test_output[24024:24031] = '{32'h0, 32'h0, 32'h0, 32'h42a9d6d2, 32'h40653373, 32'h0, 32'h0, 32'h0};
test_input[24032:24039] = '{32'hc248012f, 32'h419cc187, 32'hc0872a75, 32'hc2998ab1, 32'hc2a8a2a3, 32'hc2819699, 32'hc0647cd2, 32'h41ffc732};
test_output[24032:24039] = '{32'h0, 32'h419cc187, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ffc732};
test_input[24040:24047] = '{32'h42a7799b, 32'hc111feed, 32'hc0d070ac, 32'h42b5e126, 32'h4065a9be, 32'hc1a5d6e0, 32'h411b44e5, 32'h42632a95};
test_output[24040:24047] = '{32'h42a7799b, 32'h0, 32'h0, 32'h42b5e126, 32'h4065a9be, 32'h0, 32'h411b44e5, 32'h42632a95};
test_input[24048:24055] = '{32'hc1fdc927, 32'hc2135ea5, 32'hc0ac3abe, 32'hc1cb6ee0, 32'hc285d1ab, 32'hc1cb63e4, 32'hc207e7a8, 32'h423adcb7};
test_output[24048:24055] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423adcb7};
test_input[24056:24063] = '{32'hc2633203, 32'h4254e201, 32'h4255ed30, 32'hc2871e78, 32'hc21504f6, 32'h411490a3, 32'h4229d92d, 32'hbf0f5dc2};
test_output[24056:24063] = '{32'h0, 32'h4254e201, 32'h4255ed30, 32'h0, 32'h0, 32'h411490a3, 32'h4229d92d, 32'h0};
test_input[24064:24071] = '{32'hc23ab442, 32'h420453ff, 32'h42106c29, 32'h42bddf99, 32'hc289a50f, 32'h428d4cc7, 32'h42624695, 32'h41f59574};
test_output[24064:24071] = '{32'h0, 32'h420453ff, 32'h42106c29, 32'h42bddf99, 32'h0, 32'h428d4cc7, 32'h42624695, 32'h41f59574};
test_input[24072:24079] = '{32'hc2246e84, 32'h41aa8977, 32'h4059f62b, 32'hc0ed4d3f, 32'h42b5e9ac, 32'hc2958c93, 32'hc0516bf6, 32'hc28eb97d};
test_output[24072:24079] = '{32'h0, 32'h41aa8977, 32'h4059f62b, 32'h0, 32'h42b5e9ac, 32'h0, 32'h0, 32'h0};
test_input[24080:24087] = '{32'h428d8198, 32'hc2613d9f, 32'hc252afc6, 32'hc20919dd, 32'hc1784b4e, 32'h42aa388b, 32'h4299c484, 32'h42bfd44b};
test_output[24080:24087] = '{32'h428d8198, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42aa388b, 32'h4299c484, 32'h42bfd44b};
test_input[24088:24095] = '{32'hc2c757bc, 32'h4221a83f, 32'h42710a8d, 32'hc2462a75, 32'hc218555d, 32'hc27ea7b1, 32'h42054d84, 32'hc2986b6f};
test_output[24088:24095] = '{32'h0, 32'h4221a83f, 32'h42710a8d, 32'h0, 32'h0, 32'h0, 32'h42054d84, 32'h0};
test_input[24096:24103] = '{32'h420c1c2e, 32'hc0cbd053, 32'hc115d71d, 32'hc24740d0, 32'h42bcf213, 32'h42a2e906, 32'h42426fc8, 32'h3f37a28e};
test_output[24096:24103] = '{32'h420c1c2e, 32'h0, 32'h0, 32'h0, 32'h42bcf213, 32'h42a2e906, 32'h42426fc8, 32'h3f37a28e};
test_input[24104:24111] = '{32'hc2776537, 32'h4216abe3, 32'hc180d664, 32'h42927dea, 32'hc257fd90, 32'hc2ba8f0e, 32'h41da8f6c, 32'hc2617604};
test_output[24104:24111] = '{32'h0, 32'h4216abe3, 32'h0, 32'h42927dea, 32'h0, 32'h0, 32'h41da8f6c, 32'h0};
test_input[24112:24119] = '{32'h427e39ce, 32'hc2732d50, 32'hc25dcd11, 32'hc2aa227b, 32'h42bcac23, 32'hc00db267, 32'hc2698507, 32'hc29198a8};
test_output[24112:24119] = '{32'h427e39ce, 32'h0, 32'h0, 32'h0, 32'h42bcac23, 32'h0, 32'h0, 32'h0};
test_input[24120:24127] = '{32'h420bb234, 32'hc28b4e67, 32'h421a0b98, 32'h42be9530, 32'h4221101c, 32'hc1f08fa5, 32'h41c8d697, 32'hc124af22};
test_output[24120:24127] = '{32'h420bb234, 32'h0, 32'h421a0b98, 32'h42be9530, 32'h4221101c, 32'h0, 32'h41c8d697, 32'h0};
test_input[24128:24135] = '{32'h42c16604, 32'hc1b6b03e, 32'h42471a26, 32'h411b24a5, 32'h428f9aa6, 32'hc297bf5d, 32'hc2364249, 32'h42aec0f2};
test_output[24128:24135] = '{32'h42c16604, 32'h0, 32'h42471a26, 32'h411b24a5, 32'h428f9aa6, 32'h0, 32'h0, 32'h42aec0f2};
test_input[24136:24143] = '{32'h42a70b38, 32'hc222e119, 32'h428a8b32, 32'h42248696, 32'h41144f16, 32'h42c6ce81, 32'hc208672d, 32'hc2ade6d6};
test_output[24136:24143] = '{32'h42a70b38, 32'h0, 32'h428a8b32, 32'h42248696, 32'h41144f16, 32'h42c6ce81, 32'h0, 32'h0};
test_input[24144:24151] = '{32'h41e42e61, 32'hc2a3c4d6, 32'h40e0f405, 32'h42077315, 32'h42aa0362, 32'hc22dd995, 32'hc1aac244, 32'hc23cf631};
test_output[24144:24151] = '{32'h41e42e61, 32'h0, 32'h40e0f405, 32'h42077315, 32'h42aa0362, 32'h0, 32'h0, 32'h0};
test_input[24152:24159] = '{32'h42a81a10, 32'hc2742c4f, 32'h4264d1b3, 32'h3e461a86, 32'h42bd8fff, 32'h4239fb70, 32'hc27d9f35, 32'h427fd1da};
test_output[24152:24159] = '{32'h42a81a10, 32'h0, 32'h4264d1b3, 32'h3e461a86, 32'h42bd8fff, 32'h4239fb70, 32'h0, 32'h427fd1da};
test_input[24160:24167] = '{32'hc28137f6, 32'hc1e94e74, 32'hc2b3b3e6, 32'hc2b4c96f, 32'hc286d998, 32'hc1cbbc39, 32'hc2a2c1c1, 32'hc2c0e211};
test_output[24160:24167] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24168:24175] = '{32'h42afcce2, 32'hc28e535d, 32'hc26f67fc, 32'hc0a620e5, 32'h426be60d, 32'hc24b50c2, 32'hc224891d, 32'h3e856050};
test_output[24168:24175] = '{32'h42afcce2, 32'h0, 32'h0, 32'h0, 32'h426be60d, 32'h0, 32'h0, 32'h3e856050};
test_input[24176:24183] = '{32'h428a9e79, 32'h42ae08d7, 32'hc2258171, 32'h40f2abb9, 32'h40e38bbe, 32'h4281983f, 32'h4128dd7f, 32'h422383f1};
test_output[24176:24183] = '{32'h428a9e79, 32'h42ae08d7, 32'h0, 32'h40f2abb9, 32'h40e38bbe, 32'h4281983f, 32'h4128dd7f, 32'h422383f1};
test_input[24184:24191] = '{32'hc28d09b3, 32'h41d29a68, 32'hc2ad3e36, 32'h41e6c926, 32'hc20fc498, 32'h42a90170, 32'hc242b1a4, 32'hbf038418};
test_output[24184:24191] = '{32'h0, 32'h41d29a68, 32'h0, 32'h41e6c926, 32'h0, 32'h42a90170, 32'h0, 32'h0};
test_input[24192:24199] = '{32'h42b676b7, 32'h41966c93, 32'h3f6431ea, 32'hc29abca3, 32'h42083619, 32'h428d7a17, 32'h4184dac4, 32'hc2894de1};
test_output[24192:24199] = '{32'h42b676b7, 32'h41966c93, 32'h3f6431ea, 32'h0, 32'h42083619, 32'h428d7a17, 32'h4184dac4, 32'h0};
test_input[24200:24207] = '{32'hc008929a, 32'h4276f1f0, 32'h42bb7a29, 32'hc2a64173, 32'h41b1e327, 32'hc2951b92, 32'h423dac5f, 32'h416f973c};
test_output[24200:24207] = '{32'h0, 32'h4276f1f0, 32'h42bb7a29, 32'h0, 32'h41b1e327, 32'h0, 32'h423dac5f, 32'h416f973c};
test_input[24208:24215] = '{32'h42bb31e9, 32'hc163bc5f, 32'h41ecec3e, 32'hc104c503, 32'hc1444c77, 32'h424be78e, 32'hc2061ada, 32'h41f9e1b3};
test_output[24208:24215] = '{32'h42bb31e9, 32'h0, 32'h41ecec3e, 32'h0, 32'h0, 32'h424be78e, 32'h0, 32'h41f9e1b3};
test_input[24216:24223] = '{32'hc21b6d25, 32'h42823707, 32'h426e012d, 32'h4202b397, 32'hc09c406d, 32'h41b366a9, 32'h4259d26e, 32'hc2ae7e51};
test_output[24216:24223] = '{32'h0, 32'h42823707, 32'h426e012d, 32'h4202b397, 32'h0, 32'h41b366a9, 32'h4259d26e, 32'h0};
test_input[24224:24231] = '{32'hc2968130, 32'hc2c20c06, 32'h42a68794, 32'h425b4c8a, 32'h42adb85c, 32'h3f804ab1, 32'h4277d363, 32'h42ac48a7};
test_output[24224:24231] = '{32'h0, 32'h0, 32'h42a68794, 32'h425b4c8a, 32'h42adb85c, 32'h3f804ab1, 32'h4277d363, 32'h42ac48a7};
test_input[24232:24239] = '{32'h3f3a9b8d, 32'h42bc0f31, 32'h4270c558, 32'h42164e8c, 32'h429c04b9, 32'h42aa58ae, 32'h419e7d5c, 32'h42bf96aa};
test_output[24232:24239] = '{32'h3f3a9b8d, 32'h42bc0f31, 32'h4270c558, 32'h42164e8c, 32'h429c04b9, 32'h42aa58ae, 32'h419e7d5c, 32'h42bf96aa};
test_input[24240:24247] = '{32'hc2af7235, 32'h424c7626, 32'h423bb3db, 32'h41dbdea2, 32'h41781ee0, 32'h424a1f46, 32'hc229f251, 32'hc1e692e2};
test_output[24240:24247] = '{32'h0, 32'h424c7626, 32'h423bb3db, 32'h41dbdea2, 32'h41781ee0, 32'h424a1f46, 32'h0, 32'h0};
test_input[24248:24255] = '{32'hc28a3356, 32'hc2806fd3, 32'h428178db, 32'h416b5e96, 32'h41b43375, 32'hc0e87d00, 32'h428df5e6, 32'h427b09a4};
test_output[24248:24255] = '{32'h0, 32'h0, 32'h428178db, 32'h416b5e96, 32'h41b43375, 32'h0, 32'h428df5e6, 32'h427b09a4};
test_input[24256:24263] = '{32'hc2c2914e, 32'h42aadb97, 32'h422f3afe, 32'hc23928f7, 32'hc2aba42d, 32'hc25af2c1, 32'h42330765, 32'h41ba3efc};
test_output[24256:24263] = '{32'h0, 32'h42aadb97, 32'h422f3afe, 32'h0, 32'h0, 32'h0, 32'h42330765, 32'h41ba3efc};
test_input[24264:24271] = '{32'h421bc31b, 32'hc29597d0, 32'h4297a0a0, 32'h429c7fb5, 32'hc257fbce, 32'hc228d823, 32'h420fe722, 32'h42c52229};
test_output[24264:24271] = '{32'h421bc31b, 32'h0, 32'h4297a0a0, 32'h429c7fb5, 32'h0, 32'h0, 32'h420fe722, 32'h42c52229};
test_input[24272:24279] = '{32'h424d9155, 32'h413f1d8a, 32'hc2199815, 32'h428a426f, 32'hc260a905, 32'h42ba2281, 32'hc2971d61, 32'h4241dd98};
test_output[24272:24279] = '{32'h424d9155, 32'h413f1d8a, 32'h0, 32'h428a426f, 32'h0, 32'h42ba2281, 32'h0, 32'h4241dd98};
test_input[24280:24287] = '{32'hc27fffbf, 32'h42adf8e0, 32'hc1d065a6, 32'h4280564b, 32'h413d7369, 32'hc2a50e8e, 32'hc1a29aa6, 32'h420e8bde};
test_output[24280:24287] = '{32'h0, 32'h42adf8e0, 32'h0, 32'h4280564b, 32'h413d7369, 32'h0, 32'h0, 32'h420e8bde};
test_input[24288:24295] = '{32'h41b2f99d, 32'h42184b58, 32'hc1c89e7e, 32'h41b53d9d, 32'h42af0176, 32'h4009434e, 32'hc2a8faa3, 32'hc22e79ef};
test_output[24288:24295] = '{32'h41b2f99d, 32'h42184b58, 32'h0, 32'h41b53d9d, 32'h42af0176, 32'h4009434e, 32'h0, 32'h0};
test_input[24296:24303] = '{32'hc295edc6, 32'h41bf05c9, 32'h428bba55, 32'hc2316dce, 32'hc295393b, 32'hc289e8f7, 32'hc226c81c, 32'h41acca6e};
test_output[24296:24303] = '{32'h0, 32'h41bf05c9, 32'h428bba55, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41acca6e};
test_input[24304:24311] = '{32'h420f063e, 32'h42145bc8, 32'h41e333b6, 32'hc2b6ab3b, 32'hc1ba33bd, 32'hc216d854, 32'hc20f1088, 32'h42604800};
test_output[24304:24311] = '{32'h420f063e, 32'h42145bc8, 32'h41e333b6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42604800};
test_input[24312:24319] = '{32'h42bf6e4a, 32'h429dd6f3, 32'h41c07250, 32'h42980738, 32'h427e9fb1, 32'hbfd1d891, 32'hc27e1f7b, 32'h41b90dc2};
test_output[24312:24319] = '{32'h42bf6e4a, 32'h429dd6f3, 32'h41c07250, 32'h42980738, 32'h427e9fb1, 32'h0, 32'h0, 32'h41b90dc2};
test_input[24320:24327] = '{32'hc183080f, 32'h41f09a62, 32'h420a536d, 32'hc27a3b6b, 32'h426ba0f4, 32'h4265a183, 32'hc2981a63, 32'hc1b702c9};
test_output[24320:24327] = '{32'h0, 32'h41f09a62, 32'h420a536d, 32'h0, 32'h426ba0f4, 32'h4265a183, 32'h0, 32'h0};
test_input[24328:24335] = '{32'hc11b45e3, 32'hc19d3a47, 32'h40deac00, 32'h41ccc08c, 32'hc1da41ab, 32'hc1dd7b4d, 32'h42b346d4, 32'h3ea71923};
test_output[24328:24335] = '{32'h0, 32'h0, 32'h40deac00, 32'h41ccc08c, 32'h0, 32'h0, 32'h42b346d4, 32'h3ea71923};
test_input[24336:24343] = '{32'hc2b1bf9b, 32'hc26f8c04, 32'h416a04ce, 32'h400e76bd, 32'h429c6d1b, 32'hc2a1adca, 32'hc29fbb2e, 32'hc2b89a12};
test_output[24336:24343] = '{32'h0, 32'h0, 32'h416a04ce, 32'h400e76bd, 32'h429c6d1b, 32'h0, 32'h0, 32'h0};
test_input[24344:24351] = '{32'h40fe3c1d, 32'h428912eb, 32'hc291df28, 32'h4272403a, 32'h42b69865, 32'h424cd8c6, 32'hc248f29e, 32'hc21d6488};
test_output[24344:24351] = '{32'h40fe3c1d, 32'h428912eb, 32'h0, 32'h4272403a, 32'h42b69865, 32'h424cd8c6, 32'h0, 32'h0};
test_input[24352:24359] = '{32'hc21c78ab, 32'h42bceaa9, 32'hc2b475b4, 32'hc18a2a97, 32'h424144e8, 32'h42ab68c4, 32'hc2be13e4, 32'hc28eb776};
test_output[24352:24359] = '{32'h0, 32'h42bceaa9, 32'h0, 32'h0, 32'h424144e8, 32'h42ab68c4, 32'h0, 32'h0};
test_input[24360:24367] = '{32'hc296e0dc, 32'hc2b0ed0f, 32'h42a76eed, 32'h41c3f343, 32'h422f1624, 32'hc24fb45e, 32'hc1b17a6c, 32'h42b7ab42};
test_output[24360:24367] = '{32'h0, 32'h0, 32'h42a76eed, 32'h41c3f343, 32'h422f1624, 32'h0, 32'h0, 32'h42b7ab42};
test_input[24368:24375] = '{32'hc18bd8e3, 32'hc2bb1cfc, 32'h42998aca, 32'hc2c1aa59, 32'h422b3203, 32'hc11a3ee8, 32'hc053cc0d, 32'h42b9be1f};
test_output[24368:24375] = '{32'h0, 32'h0, 32'h42998aca, 32'h0, 32'h422b3203, 32'h0, 32'h0, 32'h42b9be1f};
test_input[24376:24383] = '{32'h42a32c15, 32'h426c7bb4, 32'h4199192c, 32'h4265dd3f, 32'hc0c1a49b, 32'h42540d3b, 32'h427faa88, 32'h41dd85a0};
test_output[24376:24383] = '{32'h42a32c15, 32'h426c7bb4, 32'h4199192c, 32'h4265dd3f, 32'h0, 32'h42540d3b, 32'h427faa88, 32'h41dd85a0};
test_input[24384:24391] = '{32'h4253fcd9, 32'h423733ad, 32'h412d0283, 32'hc21a09b5, 32'h42244c6b, 32'h426764bc, 32'hc29f0031, 32'hc215b19f};
test_output[24384:24391] = '{32'h4253fcd9, 32'h423733ad, 32'h412d0283, 32'h0, 32'h42244c6b, 32'h426764bc, 32'h0, 32'h0};
test_input[24392:24399] = '{32'h41905b72, 32'hc2b34bd9, 32'h424893b5, 32'hc2951370, 32'h41dbb909, 32'h42137437, 32'h427221f3, 32'h4178748d};
test_output[24392:24399] = '{32'h41905b72, 32'h0, 32'h424893b5, 32'h0, 32'h41dbb909, 32'h42137437, 32'h427221f3, 32'h4178748d};
test_input[24400:24407] = '{32'h425e5cab, 32'hc264f31a, 32'h425152dc, 32'hc2b8171e, 32'h42976d93, 32'hc196abb8, 32'h42c2c035, 32'hc196931e};
test_output[24400:24407] = '{32'h425e5cab, 32'h0, 32'h425152dc, 32'h0, 32'h42976d93, 32'h0, 32'h42c2c035, 32'h0};
test_input[24408:24415] = '{32'hbfba1432, 32'hc2b87c62, 32'h422d5a77, 32'hc155b706, 32'h4287684f, 32'h427fe7c8, 32'h42649240, 32'hc2bb9e76};
test_output[24408:24415] = '{32'h0, 32'h0, 32'h422d5a77, 32'h0, 32'h4287684f, 32'h427fe7c8, 32'h42649240, 32'h0};
test_input[24416:24423] = '{32'h4263d1b3, 32'hc1fa8cd3, 32'hc29c0a3d, 32'hc295ae0d, 32'hc215295e, 32'h3f8f5eb2, 32'hc1e2a5de, 32'h4264aed3};
test_output[24416:24423] = '{32'h4263d1b3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3f8f5eb2, 32'h0, 32'h4264aed3};
test_input[24424:24431] = '{32'h42c65617, 32'h42271ae7, 32'h424b2a63, 32'h411ffc69, 32'h414d4670, 32'h4272b601, 32'h41878af8, 32'h42acb12c};
test_output[24424:24431] = '{32'h42c65617, 32'h42271ae7, 32'h424b2a63, 32'h411ffc69, 32'h414d4670, 32'h4272b601, 32'h41878af8, 32'h42acb12c};
test_input[24432:24439] = '{32'hc10e47d8, 32'h418aa19b, 32'h41c2f7b5, 32'h410c6382, 32'hc297e644, 32'h41e77bda, 32'hc186616f, 32'hc29d0b19};
test_output[24432:24439] = '{32'h0, 32'h418aa19b, 32'h41c2f7b5, 32'h410c6382, 32'h0, 32'h41e77bda, 32'h0, 32'h0};
test_input[24440:24447] = '{32'h42bc8fe5, 32'h422f5dc8, 32'h424349f9, 32'h42175fd2, 32'hc2aa71ea, 32'hc118c8ee, 32'hc27d38bf, 32'hc2835e7a};
test_output[24440:24447] = '{32'h42bc8fe5, 32'h422f5dc8, 32'h424349f9, 32'h42175fd2, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24448:24455] = '{32'h41bed3ec, 32'hc2994ee2, 32'h3fe20a13, 32'h42931576, 32'h429dc001, 32'h424659ad, 32'hc2c5eca3, 32'hc2a5f04b};
test_output[24448:24455] = '{32'h41bed3ec, 32'h0, 32'h3fe20a13, 32'h42931576, 32'h429dc001, 32'h424659ad, 32'h0, 32'h0};
test_input[24456:24463] = '{32'h429acc5d, 32'hc1623b75, 32'h42b18847, 32'h42ad32ac, 32'h429bf3ea, 32'hc14eb15d, 32'hc2bb2aed, 32'h4249f222};
test_output[24456:24463] = '{32'h429acc5d, 32'h0, 32'h42b18847, 32'h42ad32ac, 32'h429bf3ea, 32'h0, 32'h0, 32'h4249f222};
test_input[24464:24471] = '{32'h4160f574, 32'h428b82a2, 32'h4195efde, 32'h40d4f211, 32'h42483582, 32'hc1d40536, 32'h421ed611, 32'h42a05c72};
test_output[24464:24471] = '{32'h4160f574, 32'h428b82a2, 32'h4195efde, 32'h40d4f211, 32'h42483582, 32'h0, 32'h421ed611, 32'h42a05c72};
test_input[24472:24479] = '{32'hc28f16f2, 32'h42a59aa3, 32'hc1ec7880, 32'hc259e6e6, 32'h419e371c, 32'h423308a3, 32'h42939922, 32'hc2c44e23};
test_output[24472:24479] = '{32'h0, 32'h42a59aa3, 32'h0, 32'h0, 32'h419e371c, 32'h423308a3, 32'h42939922, 32'h0};
test_input[24480:24487] = '{32'h41bb241a, 32'h41b5a046, 32'h4222bd7a, 32'h40bf980d, 32'h411c2d40, 32'hc2840c51, 32'h420b7102, 32'hc24384d6};
test_output[24480:24487] = '{32'h41bb241a, 32'h41b5a046, 32'h4222bd7a, 32'h40bf980d, 32'h411c2d40, 32'h0, 32'h420b7102, 32'h0};
test_input[24488:24495] = '{32'h41758061, 32'hc28e7ce9, 32'h424c22f0, 32'hc2a89d2c, 32'hc2977087, 32'h42188b0a, 32'hc0321d50, 32'hc2b73b93};
test_output[24488:24495] = '{32'h41758061, 32'h0, 32'h424c22f0, 32'h0, 32'h0, 32'h42188b0a, 32'h0, 32'h0};
test_input[24496:24503] = '{32'hc1e7f88d, 32'hc05b8447, 32'h42ba1b85, 32'h421faae9, 32'hc2936b7e, 32'hc2843ba8, 32'h429667dc, 32'h42721dad};
test_output[24496:24503] = '{32'h0, 32'h0, 32'h42ba1b85, 32'h421faae9, 32'h0, 32'h0, 32'h429667dc, 32'h42721dad};
test_input[24504:24511] = '{32'hc160051c, 32'h41d1e59b, 32'h415ed46d, 32'h426df9b1, 32'h42b4e191, 32'hc2536372, 32'hc2b81854, 32'hc23e99b8};
test_output[24504:24511] = '{32'h0, 32'h41d1e59b, 32'h415ed46d, 32'h426df9b1, 32'h42b4e191, 32'h0, 32'h0, 32'h0};
test_input[24512:24519] = '{32'hc22c4a3b, 32'h42459ba8, 32'h42ac61df, 32'h42552ccf, 32'h41d7a06a, 32'hbfd75819, 32'h4259b662, 32'h4021347c};
test_output[24512:24519] = '{32'h0, 32'h42459ba8, 32'h42ac61df, 32'h42552ccf, 32'h41d7a06a, 32'h0, 32'h4259b662, 32'h4021347c};
test_input[24520:24527] = '{32'hc1e7b61d, 32'hc15ea30f, 32'h41fa8c60, 32'hc2a10094, 32'h42910fca, 32'hc27e1092, 32'h411b346e, 32'hc25698ab};
test_output[24520:24527] = '{32'h0, 32'h0, 32'h41fa8c60, 32'h0, 32'h42910fca, 32'h0, 32'h411b346e, 32'h0};
test_input[24528:24535] = '{32'hc099e840, 32'hc2bd3a35, 32'h42b683e0, 32'h42636b0b, 32'hc2af9a10, 32'h427518a3, 32'h427e381a, 32'h423b88e7};
test_output[24528:24535] = '{32'h0, 32'h0, 32'h42b683e0, 32'h42636b0b, 32'h0, 32'h427518a3, 32'h427e381a, 32'h423b88e7};
test_input[24536:24543] = '{32'h42bd135a, 32'h41bffe36, 32'h42c0d027, 32'hc239888d, 32'hc27836cb, 32'h42a66831, 32'h41b71656, 32'hc16ac555};
test_output[24536:24543] = '{32'h42bd135a, 32'h41bffe36, 32'h42c0d027, 32'h0, 32'h0, 32'h42a66831, 32'h41b71656, 32'h0};
test_input[24544:24551] = '{32'h429103dd, 32'hc244ae8e, 32'hc229fab6, 32'hc296aa5f, 32'h42915593, 32'hc1a9be0b, 32'h41e7be75, 32'hc2310340};
test_output[24544:24551] = '{32'h429103dd, 32'h0, 32'h0, 32'h0, 32'h42915593, 32'h0, 32'h41e7be75, 32'h0};
test_input[24552:24559] = '{32'h42ad3469, 32'hc2834fef, 32'hc2ba74be, 32'h422614fb, 32'hc23f3615, 32'hc2269439, 32'h42a000a5, 32'h41660db6};
test_output[24552:24559] = '{32'h42ad3469, 32'h0, 32'h0, 32'h422614fb, 32'h0, 32'h0, 32'h42a000a5, 32'h41660db6};
test_input[24560:24567] = '{32'hc1befac5, 32'hc0d1d19c, 32'h41e08190, 32'h428f3f5d, 32'h42c550a4, 32'hc1546fea, 32'hc29fc11e, 32'h427ebabd};
test_output[24560:24567] = '{32'h0, 32'h0, 32'h41e08190, 32'h428f3f5d, 32'h42c550a4, 32'h0, 32'h0, 32'h427ebabd};
test_input[24568:24575] = '{32'hc1c8bbea, 32'h428f8de3, 32'h4253fe8d, 32'hc26e0b00, 32'h424a7a00, 32'hc29e341c, 32'h407bdc4b, 32'hc1e0f7de};
test_output[24568:24575] = '{32'h0, 32'h428f8de3, 32'h4253fe8d, 32'h0, 32'h424a7a00, 32'h0, 32'h407bdc4b, 32'h0};
test_input[24576:24583] = '{32'h42a2f358, 32'h424f5fdd, 32'hc2b9648a, 32'h411e31ca, 32'hc21e530b, 32'hc2b7ef93, 32'h41ed114d, 32'h422250c0};
test_output[24576:24583] = '{32'h42a2f358, 32'h424f5fdd, 32'h0, 32'h411e31ca, 32'h0, 32'h0, 32'h41ed114d, 32'h422250c0};
test_input[24584:24591] = '{32'h429d8303, 32'hc288946b, 32'h41ffb50e, 32'hbef22eaa, 32'h4214c12c, 32'h420ccfe2, 32'h42b7ea06, 32'hc28eb8d3};
test_output[24584:24591] = '{32'h429d8303, 32'h0, 32'h41ffb50e, 32'h0, 32'h4214c12c, 32'h420ccfe2, 32'h42b7ea06, 32'h0};
test_input[24592:24599] = '{32'hc18db621, 32'hc0b6938d, 32'h42ade0d6, 32'h419d1058, 32'hc2522614, 32'hc1fa59e9, 32'h4223ccff, 32'hc2b70d0d};
test_output[24592:24599] = '{32'h0, 32'h0, 32'h42ade0d6, 32'h419d1058, 32'h0, 32'h0, 32'h4223ccff, 32'h0};
test_input[24600:24607] = '{32'hc21883e7, 32'hc27843a7, 32'h4100066e, 32'h41f8c7b2, 32'h42349413, 32'h42086d32, 32'h41855590, 32'h42a7a5f5};
test_output[24600:24607] = '{32'h0, 32'h0, 32'h4100066e, 32'h41f8c7b2, 32'h42349413, 32'h42086d32, 32'h41855590, 32'h42a7a5f5};
test_input[24608:24615] = '{32'hc29263ec, 32'h4157acb1, 32'h42671076, 32'hc2151b83, 32'h422bc977, 32'h421df216, 32'hc256b501, 32'hc259bd63};
test_output[24608:24615] = '{32'h0, 32'h4157acb1, 32'h42671076, 32'h0, 32'h422bc977, 32'h421df216, 32'h0, 32'h0};
test_input[24616:24623] = '{32'h419669f1, 32'hc2a59228, 32'h424edaf0, 32'hc260279f, 32'h420c2c2e, 32'h4287cb85, 32'h411fca43, 32'h41d834d1};
test_output[24616:24623] = '{32'h419669f1, 32'h0, 32'h424edaf0, 32'h0, 32'h420c2c2e, 32'h4287cb85, 32'h411fca43, 32'h41d834d1};
test_input[24624:24631] = '{32'hc27e23fc, 32'h4270242f, 32'h41983346, 32'hc250059d, 32'hc2a02e42, 32'h4257392c, 32'h408908f9, 32'h425f4359};
test_output[24624:24631] = '{32'h0, 32'h4270242f, 32'h41983346, 32'h0, 32'h0, 32'h4257392c, 32'h408908f9, 32'h425f4359};
test_input[24632:24639] = '{32'h41b95c8a, 32'h419814f5, 32'h41522122, 32'h42a18243, 32'h40997141, 32'hc1e2d124, 32'h4225683c, 32'hc29ca4a2};
test_output[24632:24639] = '{32'h41b95c8a, 32'h419814f5, 32'h41522122, 32'h42a18243, 32'h40997141, 32'h0, 32'h4225683c, 32'h0};
test_input[24640:24647] = '{32'hc251eb80, 32'h4248c017, 32'h428f1ac7, 32'h42997488, 32'h408ba857, 32'h429678cd, 32'h42b1b7ac, 32'h420f2673};
test_output[24640:24647] = '{32'h0, 32'h4248c017, 32'h428f1ac7, 32'h42997488, 32'h408ba857, 32'h429678cd, 32'h42b1b7ac, 32'h420f2673};
test_input[24648:24655] = '{32'h42a63b03, 32'hc1af620c, 32'hc2ab6b92, 32'h416365ab, 32'h4092a7a5, 32'h422bf920, 32'h418f4527, 32'h402cb3fb};
test_output[24648:24655] = '{32'h42a63b03, 32'h0, 32'h0, 32'h416365ab, 32'h4092a7a5, 32'h422bf920, 32'h418f4527, 32'h402cb3fb};
test_input[24656:24663] = '{32'hc2a418fd, 32'h421f503f, 32'h41afcbec, 32'h423628f9, 32'h42004fbd, 32'hc2b23c30, 32'hc268d36f, 32'h42a72ad9};
test_output[24656:24663] = '{32'h0, 32'h421f503f, 32'h41afcbec, 32'h423628f9, 32'h42004fbd, 32'h0, 32'h0, 32'h42a72ad9};
test_input[24664:24671] = '{32'hc12a805f, 32'h425282cc, 32'h4119da7a, 32'h420abd2c, 32'hc2399e54, 32'h42c6a10e, 32'hc1c93dc0, 32'h4266d398};
test_output[24664:24671] = '{32'h0, 32'h425282cc, 32'h4119da7a, 32'h420abd2c, 32'h0, 32'h42c6a10e, 32'h0, 32'h4266d398};
test_input[24672:24679] = '{32'h40d995a0, 32'hbf884d64, 32'h41a9af8e, 32'h41157479, 32'h420b3a91, 32'h40f9a3ee, 32'h41fb4eea, 32'hc1a22709};
test_output[24672:24679] = '{32'h40d995a0, 32'h0, 32'h41a9af8e, 32'h41157479, 32'h420b3a91, 32'h40f9a3ee, 32'h41fb4eea, 32'h0};
test_input[24680:24687] = '{32'h42b00b4d, 32'hc2c70a11, 32'h42b499cd, 32'h416e5026, 32'h42b0168c, 32'h41dad1f7, 32'h422f02f0, 32'h4234d443};
test_output[24680:24687] = '{32'h42b00b4d, 32'h0, 32'h42b499cd, 32'h416e5026, 32'h42b0168c, 32'h41dad1f7, 32'h422f02f0, 32'h4234d443};
test_input[24688:24695] = '{32'hc2aa3653, 32'h4220e701, 32'hc27201f8, 32'h423fcaeb, 32'hc19ea15b, 32'hc242ae88, 32'hc1d979c8, 32'h41707617};
test_output[24688:24695] = '{32'h0, 32'h4220e701, 32'h0, 32'h423fcaeb, 32'h0, 32'h0, 32'h0, 32'h41707617};
test_input[24696:24703] = '{32'h423aa4be, 32'hc22898ed, 32'h42af610c, 32'h42c682f8, 32'hc1232ae3, 32'h4281c503, 32'h42878d93, 32'hc2426866};
test_output[24696:24703] = '{32'h423aa4be, 32'h0, 32'h42af610c, 32'h42c682f8, 32'h0, 32'h4281c503, 32'h42878d93, 32'h0};
test_input[24704:24711] = '{32'hc2b299cd, 32'hc21ee4b0, 32'hc290c941, 32'h42382ba5, 32'h427d4278, 32'hc2828d57, 32'hc2c5ecb3, 32'h422439d6};
test_output[24704:24711] = '{32'h0, 32'h0, 32'h0, 32'h42382ba5, 32'h427d4278, 32'h0, 32'h0, 32'h422439d6};
test_input[24712:24719] = '{32'hc11201c0, 32'hc23447f3, 32'h4210c7ff, 32'hc1ec03d4, 32'hc1c8b125, 32'hc2720f3f, 32'h427b2b95, 32'h424c39fa};
test_output[24712:24719] = '{32'h0, 32'h0, 32'h4210c7ff, 32'h0, 32'h0, 32'h0, 32'h427b2b95, 32'h424c39fa};
test_input[24720:24727] = '{32'h41c4c55c, 32'hc2941926, 32'hc253d5b6, 32'h3f508f0d, 32'hc23f9519, 32'h42c443d4, 32'hc22d4ccc, 32'hc257e057};
test_output[24720:24727] = '{32'h41c4c55c, 32'h0, 32'h0, 32'h3f508f0d, 32'h0, 32'h42c443d4, 32'h0, 32'h0};
test_input[24728:24735] = '{32'hc223f0dd, 32'h4243be85, 32'h4216d2ca, 32'h42469de6, 32'hc0c705e0, 32'hc27c8667, 32'h42bdfbea, 32'hc19c0567};
test_output[24728:24735] = '{32'h0, 32'h4243be85, 32'h4216d2ca, 32'h42469de6, 32'h0, 32'h0, 32'h42bdfbea, 32'h0};
test_input[24736:24743] = '{32'h4299153d, 32'hc1873efb, 32'h4285dcb3, 32'h4002014c, 32'h426c6e31, 32'hc2388b4e, 32'h426864d6, 32'h41df53bc};
test_output[24736:24743] = '{32'h4299153d, 32'h0, 32'h4285dcb3, 32'h4002014c, 32'h426c6e31, 32'h0, 32'h426864d6, 32'h41df53bc};
test_input[24744:24751] = '{32'hc2b66ad4, 32'hc2a1a090, 32'h426aa13c, 32'hc1461e62, 32'hc2bfb485, 32'h41a1e31c, 32'h3f5945ec, 32'hc2c6aa89};
test_output[24744:24751] = '{32'h0, 32'h0, 32'h426aa13c, 32'h0, 32'h0, 32'h41a1e31c, 32'h3f5945ec, 32'h0};
test_input[24752:24759] = '{32'hc2acf164, 32'hc28f1bb4, 32'h42876218, 32'hc2593b47, 32'hc18ffb06, 32'hc274ce59, 32'h42a6c291, 32'h42ac5a0b};
test_output[24752:24759] = '{32'h0, 32'h0, 32'h42876218, 32'h0, 32'h0, 32'h0, 32'h42a6c291, 32'h42ac5a0b};
test_input[24760:24767] = '{32'hc28f909b, 32'h428e9d42, 32'h420c213e, 32'h415ab511, 32'hc1800268, 32'h427f60ec, 32'h424da715, 32'hc181f14c};
test_output[24760:24767] = '{32'h0, 32'h428e9d42, 32'h420c213e, 32'h415ab511, 32'h0, 32'h427f60ec, 32'h424da715, 32'h0};
test_input[24768:24775] = '{32'h4248a816, 32'h42382166, 32'h41929b5a, 32'hc2b61ddd, 32'h426be67c, 32'hc00f512f, 32'h411bdfe9, 32'hc1e81244};
test_output[24768:24775] = '{32'h4248a816, 32'h42382166, 32'h41929b5a, 32'h0, 32'h426be67c, 32'h0, 32'h411bdfe9, 32'h0};
test_input[24776:24783] = '{32'hc1de41da, 32'hc21838db, 32'h40d22e16, 32'hc1dc12d6, 32'h42c12d99, 32'h42ac38fe, 32'hc1d95494, 32'hc28435f0};
test_output[24776:24783] = '{32'h0, 32'h0, 32'h40d22e16, 32'h0, 32'h42c12d99, 32'h42ac38fe, 32'h0, 32'h0};
test_input[24784:24791] = '{32'h401e745e, 32'h411d4514, 32'hc2bfc71a, 32'hc2964acd, 32'hc1e86dca, 32'h428f7c50, 32'h42998201, 32'hc18842ef};
test_output[24784:24791] = '{32'h401e745e, 32'h411d4514, 32'h0, 32'h0, 32'h0, 32'h428f7c50, 32'h42998201, 32'h0};
test_input[24792:24799] = '{32'hc178efb2, 32'h4296cbf6, 32'hc2b11174, 32'h42b34879, 32'h42184461, 32'h4272b36d, 32'h42a15267, 32'hc2903d3f};
test_output[24792:24799] = '{32'h0, 32'h4296cbf6, 32'h0, 32'h42b34879, 32'h42184461, 32'h4272b36d, 32'h42a15267, 32'h0};
test_input[24800:24807] = '{32'h426cce88, 32'h423909fa, 32'h4115331a, 32'h427e2443, 32'hc2ad4cc3, 32'hc0fd0588, 32'hc28f28ee, 32'hc1b585c0};
test_output[24800:24807] = '{32'h426cce88, 32'h423909fa, 32'h4115331a, 32'h427e2443, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24808:24815] = '{32'hc2051718, 32'hc18662c0, 32'hc28d2341, 32'h42333b2f, 32'hc24ed6d6, 32'h418d0804, 32'h427f7e5c, 32'h41914242};
test_output[24808:24815] = '{32'h0, 32'h0, 32'h0, 32'h42333b2f, 32'h0, 32'h418d0804, 32'h427f7e5c, 32'h41914242};
test_input[24816:24823] = '{32'h41b648ad, 32'hc2303a9f, 32'hc28324f7, 32'h428c1365, 32'hc2a05c9c, 32'h42aea645, 32'h42b961e1, 32'hc29ed5b8};
test_output[24816:24823] = '{32'h41b648ad, 32'h0, 32'h0, 32'h428c1365, 32'h0, 32'h42aea645, 32'h42b961e1, 32'h0};
test_input[24824:24831] = '{32'hc2c334ab, 32'hc0aedc24, 32'h42be69ae, 32'hc26b21d9, 32'hc2bad3c2, 32'h428ecb5f, 32'hc28bd030, 32'hc2c31a67};
test_output[24824:24831] = '{32'h0, 32'h0, 32'h42be69ae, 32'h0, 32'h0, 32'h428ecb5f, 32'h0, 32'h0};
test_input[24832:24839] = '{32'h422e49e4, 32'h42830e07, 32'h42b5d932, 32'h4293bede, 32'h41012fc4, 32'hc241b176, 32'h422c41a5, 32'hc2931406};
test_output[24832:24839] = '{32'h422e49e4, 32'h42830e07, 32'h42b5d932, 32'h4293bede, 32'h41012fc4, 32'h0, 32'h422c41a5, 32'h0};
test_input[24840:24847] = '{32'h40cd1e38, 32'h4233d0e9, 32'h422967bc, 32'hc196d17d, 32'hc229b99d, 32'h424dc8f3, 32'hc22a2020, 32'h4235e7a1};
test_output[24840:24847] = '{32'h40cd1e38, 32'h4233d0e9, 32'h422967bc, 32'h0, 32'h0, 32'h424dc8f3, 32'h0, 32'h4235e7a1};
test_input[24848:24855] = '{32'hc240f7d5, 32'hc28c3240, 32'h42890aa1, 32'hc2a721ea, 32'hc283a499, 32'h4285a71e, 32'hc23325ec, 32'hc2abdd94};
test_output[24848:24855] = '{32'h0, 32'h0, 32'h42890aa1, 32'h0, 32'h0, 32'h4285a71e, 32'h0, 32'h0};
test_input[24856:24863] = '{32'hc286fe05, 32'hc1b7fab0, 32'hc1bc3cf1, 32'hc269d562, 32'h42961a87, 32'h41a8a713, 32'hc1d59f7b, 32'h429db689};
test_output[24856:24863] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42961a87, 32'h41a8a713, 32'h0, 32'h429db689};
test_input[24864:24871] = '{32'hc136818a, 32'h42909ec5, 32'hc2aff29e, 32'h42894f4e, 32'h42c5bf32, 32'h42afce7d, 32'h42a1defc, 32'hc1db91d9};
test_output[24864:24871] = '{32'h0, 32'h42909ec5, 32'h0, 32'h42894f4e, 32'h42c5bf32, 32'h42afce7d, 32'h42a1defc, 32'h0};
test_input[24872:24879] = '{32'hc1024c2e, 32'h4272ac3a, 32'hc1af59a5, 32'h423f7abe, 32'hc20e03e8, 32'h421a562f, 32'hc1a1f0c9, 32'h42bf7dd5};
test_output[24872:24879] = '{32'h0, 32'h4272ac3a, 32'h0, 32'h423f7abe, 32'h0, 32'h421a562f, 32'h0, 32'h42bf7dd5};
test_input[24880:24887] = '{32'h42abc1fb, 32'hc25d08f9, 32'hc2290fb8, 32'hc133e9ad, 32'h42b73c49, 32'h409cbb61, 32'hc2b1e5a8, 32'h42b26103};
test_output[24880:24887] = '{32'h42abc1fb, 32'h0, 32'h0, 32'h0, 32'h42b73c49, 32'h409cbb61, 32'h0, 32'h42b26103};
test_input[24888:24895] = '{32'h41984f7f, 32'hc2c2d681, 32'h412f19be, 32'hc20f4c5b, 32'h425002cf, 32'hc18e6ec2, 32'hc29cbbc6, 32'hc28bdfd5};
test_output[24888:24895] = '{32'h41984f7f, 32'h0, 32'h412f19be, 32'h0, 32'h425002cf, 32'h0, 32'h0, 32'h0};
test_input[24896:24903] = '{32'h425fee5c, 32'hc21e28bd, 32'h42a46861, 32'h428949b1, 32'hc1e92875, 32'hc260e422, 32'hc232ee92, 32'hc140003d};
test_output[24896:24903] = '{32'h425fee5c, 32'h0, 32'h42a46861, 32'h428949b1, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24904:24911] = '{32'hc0950a94, 32'hc22cbf76, 32'hc29d48ad, 32'hc2921529, 32'h42af5bde, 32'h41361f2a, 32'h41b8f3b2, 32'hc29c5ac9};
test_output[24904:24911] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42af5bde, 32'h41361f2a, 32'h41b8f3b2, 32'h0};
test_input[24912:24919] = '{32'hc1b0a71c, 32'hc24631a5, 32'h41c616bc, 32'hc2267131, 32'hc1fee037, 32'h422d9d70, 32'h42204089, 32'h42becb1d};
test_output[24912:24919] = '{32'h0, 32'h0, 32'h41c616bc, 32'h0, 32'h0, 32'h422d9d70, 32'h42204089, 32'h42becb1d};
test_input[24920:24927] = '{32'hc28c4b03, 32'h42119c9a, 32'h429f5ac5, 32'hc2b07ca8, 32'h428a3ac5, 32'h420ad8cb, 32'h421a3414, 32'hc12bdd77};
test_output[24920:24927] = '{32'h0, 32'h42119c9a, 32'h429f5ac5, 32'h0, 32'h428a3ac5, 32'h420ad8cb, 32'h421a3414, 32'h0};
test_input[24928:24935] = '{32'hc23f7de7, 32'h419ee99e, 32'h41b8caaf, 32'hc2b752d8, 32'h42368e16, 32'h425335e1, 32'hc2bc18f6, 32'hc2981dd8};
test_output[24928:24935] = '{32'h0, 32'h419ee99e, 32'h41b8caaf, 32'h0, 32'h42368e16, 32'h425335e1, 32'h0, 32'h0};
test_input[24936:24943] = '{32'hc12e1567, 32'hc280e2f2, 32'hc2ab60a4, 32'hc1dcfe1e, 32'hc2756ccd, 32'h4230459c, 32'hc296119f, 32'hc20daf7d};
test_output[24936:24943] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4230459c, 32'h0, 32'h0};
test_input[24944:24951] = '{32'h42b0bd7f, 32'hc216f695, 32'h428f83db, 32'h427d517d, 32'hc2aae9d4, 32'hc29831d5, 32'h42a70342, 32'hc1be60c5};
test_output[24944:24951] = '{32'h42b0bd7f, 32'h0, 32'h428f83db, 32'h427d517d, 32'h0, 32'h0, 32'h42a70342, 32'h0};
test_input[24952:24959] = '{32'hc23862f9, 32'hc293b2dd, 32'hc199bb84, 32'h41b0ef80, 32'hc2a0d76d, 32'h42bcbe74, 32'h40de27df, 32'h4244a4c0};
test_output[24952:24959] = '{32'h0, 32'h0, 32'h0, 32'h41b0ef80, 32'h0, 32'h42bcbe74, 32'h40de27df, 32'h4244a4c0};
test_input[24960:24967] = '{32'hc22cf664, 32'hc20bca31, 32'hc1811149, 32'hc1d8a97c, 32'hc28a142a, 32'h4209c9a2, 32'h418ab8b3, 32'hc21a88b9};
test_output[24960:24967] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4209c9a2, 32'h418ab8b3, 32'h0};
test_input[24968:24975] = '{32'hc2c1c854, 32'hc27e9f52, 32'hc2441fcc, 32'hc29e459a, 32'h42900677, 32'h40a83067, 32'hc1e3a8d9, 32'hc2818464};
test_output[24968:24975] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42900677, 32'h40a83067, 32'h0, 32'h0};
test_input[24976:24983] = '{32'h4293697d, 32'h41f1128c, 32'hc1cc430a, 32'h42c023ae, 32'hc127e4f1, 32'hc29740bb, 32'hc2a57959, 32'hc18db284};
test_output[24976:24983] = '{32'h4293697d, 32'h41f1128c, 32'h0, 32'h42c023ae, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[24984:24991] = '{32'h42bbdeb7, 32'h42557bfb, 32'h42a864b8, 32'hc1922557, 32'hc2305fba, 32'hc130da33, 32'hc2c4da76, 32'h427fffd3};
test_output[24984:24991] = '{32'h42bbdeb7, 32'h42557bfb, 32'h42a864b8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427fffd3};
test_input[24992:24999] = '{32'hc1dc0ee2, 32'hc0193984, 32'hc2933337, 32'h4231fabe, 32'h41d0c7bb, 32'hc096cd84, 32'hc21b0dbf, 32'h4092aaf8};
test_output[24992:24999] = '{32'h0, 32'h0, 32'h0, 32'h4231fabe, 32'h41d0c7bb, 32'h0, 32'h0, 32'h4092aaf8};
test_input[25000:25007] = '{32'hc2775812, 32'hc2684e21, 32'h41874261, 32'hc1f1fad7, 32'hc2b439af, 32'h416b7e53, 32'hc2bdc10d, 32'h42be1c22};
test_output[25000:25007] = '{32'h0, 32'h0, 32'h41874261, 32'h0, 32'h0, 32'h416b7e53, 32'h0, 32'h42be1c22};
test_input[25008:25015] = '{32'hc2ba1725, 32'h42802fb3, 32'hc2c61797, 32'hc227861d, 32'hc1ff2711, 32'hc28a31dc, 32'hc28eaf13, 32'hc29319ab};
test_output[25008:25015] = '{32'h0, 32'h42802fb3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25016:25023] = '{32'hc213fa93, 32'h4191c9be, 32'hc17cbffd, 32'hc14bf5f2, 32'hc135ae84, 32'h429281ba, 32'hc2a9fe33, 32'hc23743e7};
test_output[25016:25023] = '{32'h0, 32'h4191c9be, 32'h0, 32'h0, 32'h0, 32'h429281ba, 32'h0, 32'h0};
test_input[25024:25031] = '{32'h42be8907, 32'h4173b169, 32'hc2b6dcad, 32'h4289ff6b, 32'h421d5739, 32'hc2803682, 32'h4127143c, 32'hc2ab0227};
test_output[25024:25031] = '{32'h42be8907, 32'h4173b169, 32'h0, 32'h4289ff6b, 32'h421d5739, 32'h0, 32'h4127143c, 32'h0};
test_input[25032:25039] = '{32'hc19b243f, 32'h41da691c, 32'hc240e847, 32'hc2886213, 32'hc2c3b35d, 32'hc2a55ad1, 32'hc1edcf94, 32'h422b5898};
test_output[25032:25039] = '{32'h0, 32'h41da691c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422b5898};
test_input[25040:25047] = '{32'hc28f10ce, 32'h42b130a1, 32'h4268ceaa, 32'h424efe81, 32'hc260dcb6, 32'hc2ac36bd, 32'hbf93bda0, 32'hc2864bf3};
test_output[25040:25047] = '{32'h0, 32'h42b130a1, 32'h4268ceaa, 32'h424efe81, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25048:25055] = '{32'hc2c5fa7a, 32'h418e68bc, 32'h420841ed, 32'hc251aa52, 32'hc2349250, 32'h4223074f, 32'hc1ad0b58, 32'h42773a08};
test_output[25048:25055] = '{32'h0, 32'h418e68bc, 32'h420841ed, 32'h0, 32'h0, 32'h4223074f, 32'h0, 32'h42773a08};
test_input[25056:25063] = '{32'hc29a33b8, 32'hc21f2d7f, 32'h42c58f51, 32'hc2bf5951, 32'hc25f6439, 32'hc200a6d8, 32'hc26e6734, 32'h42b5c323};
test_output[25056:25063] = '{32'h0, 32'h0, 32'h42c58f51, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b5c323};
test_input[25064:25071] = '{32'h42b0ee3c, 32'h42afd141, 32'h41a1b328, 32'hc2548252, 32'h42afdcec, 32'hc21cc165, 32'hc1f5b165, 32'h42696cb1};
test_output[25064:25071] = '{32'h42b0ee3c, 32'h42afd141, 32'h41a1b328, 32'h0, 32'h42afdcec, 32'h0, 32'h0, 32'h42696cb1};
test_input[25072:25079] = '{32'hc280b54a, 32'hc2ba41af, 32'h425a8b9b, 32'h41f77084, 32'h42944b83, 32'h423176ec, 32'h42454140, 32'h42010fc7};
test_output[25072:25079] = '{32'h0, 32'h0, 32'h425a8b9b, 32'h41f77084, 32'h42944b83, 32'h423176ec, 32'h42454140, 32'h42010fc7};
test_input[25080:25087] = '{32'hc1b6d4e7, 32'h41cefb5b, 32'h41dc14a9, 32'h41acec10, 32'h404fb22c, 32'h41aef64a, 32'hc1f62c41, 32'h41f526db};
test_output[25080:25087] = '{32'h0, 32'h41cefb5b, 32'h41dc14a9, 32'h41acec10, 32'h404fb22c, 32'h41aef64a, 32'h0, 32'h41f526db};
test_input[25088:25095] = '{32'hc1d66cb9, 32'hc27e15cf, 32'hc29ae7f1, 32'hc22eb7f8, 32'h42a71095, 32'hc25a1eac, 32'h42c4e568, 32'h42062ecc};
test_output[25088:25095] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a71095, 32'h0, 32'h42c4e568, 32'h42062ecc};
test_input[25096:25103] = '{32'hc13f5c12, 32'hc2b40a0f, 32'hc0861be2, 32'h4221b3ef, 32'hc2a52c8e, 32'hc1b726a9, 32'h429c6695, 32'h41ef6a76};
test_output[25096:25103] = '{32'h0, 32'h0, 32'h0, 32'h4221b3ef, 32'h0, 32'h0, 32'h429c6695, 32'h41ef6a76};
test_input[25104:25111] = '{32'h417902e4, 32'h40d35e5b, 32'hc2347cfd, 32'hc255dec0, 32'h42a08eb4, 32'h42b31ed3, 32'h4111b7ea, 32'h4104aa39};
test_output[25104:25111] = '{32'h417902e4, 32'h40d35e5b, 32'h0, 32'h0, 32'h42a08eb4, 32'h42b31ed3, 32'h4111b7ea, 32'h4104aa39};
test_input[25112:25119] = '{32'hbf29efb7, 32'hc24cab8b, 32'h3f4c5bf6, 32'hbf8c1791, 32'h424b71d3, 32'hc2b8d0a7, 32'h429591c0, 32'hc2b3758d};
test_output[25112:25119] = '{32'h0, 32'h0, 32'h3f4c5bf6, 32'h0, 32'h424b71d3, 32'h0, 32'h429591c0, 32'h0};
test_input[25120:25127] = '{32'hc19944b3, 32'hc12c3ab0, 32'h42327425, 32'hc239b98d, 32'h419e4d39, 32'h415a8f7a, 32'hc2b9ebaf, 32'h41ad8a13};
test_output[25120:25127] = '{32'h0, 32'h0, 32'h42327425, 32'h0, 32'h419e4d39, 32'h415a8f7a, 32'h0, 32'h41ad8a13};
test_input[25128:25135] = '{32'hc1dba466, 32'hc2801d43, 32'hc2ac0aa2, 32'hc1aab5ff, 32'hc2264826, 32'hc2a4ca85, 32'h420cde1c, 32'hc0ee1688};
test_output[25128:25135] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h420cde1c, 32'h0};
test_input[25136:25143] = '{32'h42b5013d, 32'hc135fb19, 32'h428fc55c, 32'hbe98b371, 32'hc2c14e9f, 32'h4260aea1, 32'hc22cb5f5, 32'h42b01655};
test_output[25136:25143] = '{32'h42b5013d, 32'h0, 32'h428fc55c, 32'h0, 32'h0, 32'h4260aea1, 32'h0, 32'h42b01655};
test_input[25144:25151] = '{32'h40abb06d, 32'hc0226974, 32'hc29d1a6e, 32'h41fd7d15, 32'h419dd963, 32'hc1355741, 32'hc1ddee9e, 32'hc2545e4a};
test_output[25144:25151] = '{32'h40abb06d, 32'h0, 32'h0, 32'h41fd7d15, 32'h419dd963, 32'h0, 32'h0, 32'h0};
test_input[25152:25159] = '{32'hc275cfdc, 32'hc2a12ca9, 32'hc1c49055, 32'hc2689be5, 32'hc2730280, 32'hc26f73a0, 32'hc214a30b, 32'hc1fea5fd};
test_output[25152:25159] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25160:25167] = '{32'hc29b66e1, 32'hc2a4050b, 32'h42c31e79, 32'h42659df2, 32'hc25a258d, 32'h424c8f12, 32'hc2b9be41, 32'hc2b2e6b2};
test_output[25160:25167] = '{32'h0, 32'h0, 32'h42c31e79, 32'h42659df2, 32'h0, 32'h424c8f12, 32'h0, 32'h0};
test_input[25168:25175] = '{32'hc26c7464, 32'h4211ebc6, 32'h426a47dd, 32'h426f2fe4, 32'hc2a26800, 32'hc2909813, 32'hbfbf9a55, 32'h42b0d330};
test_output[25168:25175] = '{32'h0, 32'h4211ebc6, 32'h426a47dd, 32'h426f2fe4, 32'h0, 32'h0, 32'h0, 32'h42b0d330};
test_input[25176:25183] = '{32'hc1311c28, 32'h42947e7d, 32'h418af7ec, 32'h42bf3eb9, 32'hc2ba1e32, 32'h41f06836, 32'hc1fa4d0c, 32'hc2b5a99e};
test_output[25176:25183] = '{32'h0, 32'h42947e7d, 32'h418af7ec, 32'h42bf3eb9, 32'h0, 32'h41f06836, 32'h0, 32'h0};
test_input[25184:25191] = '{32'h42bb998e, 32'hc27af2ec, 32'hc1bbdeb8, 32'h4286383a, 32'hc0780cf4, 32'hc18fffd6, 32'h42c6f45d, 32'hc287d61a};
test_output[25184:25191] = '{32'h42bb998e, 32'h0, 32'h0, 32'h4286383a, 32'h0, 32'h0, 32'h42c6f45d, 32'h0};
test_input[25192:25199] = '{32'h4255698b, 32'h4253a290, 32'hc14b628e, 32'hc285b780, 32'h41f4839c, 32'hc2890fa1, 32'hc1917608, 32'hc23c898a};
test_output[25192:25199] = '{32'h4255698b, 32'h4253a290, 32'h0, 32'h0, 32'h41f4839c, 32'h0, 32'h0, 32'h0};
test_input[25200:25207] = '{32'hc194142b, 32'h428c993f, 32'h428217d1, 32'h3ed07235, 32'h422bbafb, 32'h4047f419, 32'h428d3aff, 32'h42a47284};
test_output[25200:25207] = '{32'h0, 32'h428c993f, 32'h428217d1, 32'h3ed07235, 32'h422bbafb, 32'h4047f419, 32'h428d3aff, 32'h42a47284};
test_input[25208:25215] = '{32'h410086a6, 32'h4253df85, 32'hc28628c0, 32'h427ca612, 32'hc20e24bc, 32'h4031599c, 32'hc18a0286, 32'h42b1403d};
test_output[25208:25215] = '{32'h410086a6, 32'h4253df85, 32'h0, 32'h427ca612, 32'h0, 32'h4031599c, 32'h0, 32'h42b1403d};
test_input[25216:25223] = '{32'hc2b8d263, 32'h425a587d, 32'hc212c493, 32'h42c691fc, 32'h427d6d44, 32'h418711f8, 32'hc21d256a, 32'h42665144};
test_output[25216:25223] = '{32'h0, 32'h425a587d, 32'h0, 32'h42c691fc, 32'h427d6d44, 32'h418711f8, 32'h0, 32'h42665144};
test_input[25224:25231] = '{32'hc194537d, 32'hc2830727, 32'hc15fc302, 32'hc188f22c, 32'h425c458b, 32'h419d98fa, 32'h4240e087, 32'h42a9b03d};
test_output[25224:25231] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h425c458b, 32'h419d98fa, 32'h4240e087, 32'h42a9b03d};
test_input[25232:25239] = '{32'h41db3c41, 32'h429b7cf2, 32'hc29afd5e, 32'hc18c304b, 32'hc2b9a59b, 32'h424fed68, 32'h42c4ad92, 32'hc288fb7b};
test_output[25232:25239] = '{32'h41db3c41, 32'h429b7cf2, 32'h0, 32'h0, 32'h0, 32'h424fed68, 32'h42c4ad92, 32'h0};
test_input[25240:25247] = '{32'h42b02fbd, 32'hc2b5e90e, 32'hc29dd8e6, 32'hc1efc0ba, 32'h42913082, 32'h427f0b24, 32'h42690fbe, 32'h425c521f};
test_output[25240:25247] = '{32'h42b02fbd, 32'h0, 32'h0, 32'h0, 32'h42913082, 32'h427f0b24, 32'h42690fbe, 32'h425c521f};
test_input[25248:25255] = '{32'hc2ae3d00, 32'h42bd88ac, 32'hc253da19, 32'hc287319d, 32'hc2298202, 32'hc245881c, 32'hc2287350, 32'h422457fb};
test_output[25248:25255] = '{32'h0, 32'h42bd88ac, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422457fb};
test_input[25256:25263] = '{32'h4196b69b, 32'hc2932b30, 32'h403ab224, 32'h4295ff56, 32'hc1b194ab, 32'h41d070ef, 32'hc2452c88, 32'h41b70bf3};
test_output[25256:25263] = '{32'h4196b69b, 32'h0, 32'h403ab224, 32'h4295ff56, 32'h0, 32'h41d070ef, 32'h0, 32'h41b70bf3};
test_input[25264:25271] = '{32'hc29d499d, 32'hc27279f3, 32'hc203f9ea, 32'hc244f1e6, 32'hc2957583, 32'hc2015aef, 32'hc28e1841, 32'h428677c1};
test_output[25264:25271] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428677c1};
test_input[25272:25279] = '{32'hc1d6cd49, 32'hc273cfc0, 32'h423ffc21, 32'h42819546, 32'hc0c3890e, 32'hc14b7432, 32'hc269ff75, 32'hc2b6c15f};
test_output[25272:25279] = '{32'h0, 32'h0, 32'h423ffc21, 32'h42819546, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25280:25287] = '{32'hc2793edb, 32'hc27a5318, 32'h409286a1, 32'h42392722, 32'h41060546, 32'h42ae3ae2, 32'h41e56650, 32'h420a7f1e};
test_output[25280:25287] = '{32'h0, 32'h0, 32'h409286a1, 32'h42392722, 32'h41060546, 32'h42ae3ae2, 32'h41e56650, 32'h420a7f1e};
test_input[25288:25295] = '{32'hc230b90d, 32'h420f2644, 32'h4205e1fc, 32'h4240fb7e, 32'h41f48653, 32'h429020cc, 32'h41e067b0, 32'hc2b2f7e6};
test_output[25288:25295] = '{32'h0, 32'h420f2644, 32'h4205e1fc, 32'h4240fb7e, 32'h41f48653, 32'h429020cc, 32'h41e067b0, 32'h0};
test_input[25296:25303] = '{32'hc21d4a40, 32'hc2a97093, 32'h426a9e0e, 32'h429c44ad, 32'h4243da5a, 32'hc234a948, 32'h4290a6e3, 32'h42c7c118};
test_output[25296:25303] = '{32'h0, 32'h0, 32'h426a9e0e, 32'h429c44ad, 32'h4243da5a, 32'h0, 32'h4290a6e3, 32'h42c7c118};
test_input[25304:25311] = '{32'h426f82b6, 32'h42171fe7, 32'hc29316cf, 32'h42bc99bd, 32'h41fb4529, 32'h422291b0, 32'h425755e2, 32'h42511bca};
test_output[25304:25311] = '{32'h426f82b6, 32'h42171fe7, 32'h0, 32'h42bc99bd, 32'h41fb4529, 32'h422291b0, 32'h425755e2, 32'h42511bca};
test_input[25312:25319] = '{32'h424e22d1, 32'hc2af82f9, 32'h422057da, 32'hc2297527, 32'hc29c899e, 32'hc2969cbd, 32'hc2a885e7, 32'hc206b269};
test_output[25312:25319] = '{32'h424e22d1, 32'h0, 32'h422057da, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25320:25327] = '{32'h42c1ee34, 32'h428d3313, 32'h42046cfa, 32'h41ecbd69, 32'hc23d7d2b, 32'h42b6b9e4, 32'h4117fc9e, 32'hc200d182};
test_output[25320:25327] = '{32'h42c1ee34, 32'h428d3313, 32'h42046cfa, 32'h41ecbd69, 32'h0, 32'h42b6b9e4, 32'h4117fc9e, 32'h0};
test_input[25328:25335] = '{32'h41a110ef, 32'hc2bbac57, 32'hc18ee80b, 32'h42c0ec09, 32'hc247a9cf, 32'hc2b2a096, 32'h423bbef5, 32'hc0e8bd42};
test_output[25328:25335] = '{32'h41a110ef, 32'h0, 32'h0, 32'h42c0ec09, 32'h0, 32'h0, 32'h423bbef5, 32'h0};
test_input[25336:25343] = '{32'hc280eadf, 32'h42a8eb07, 32'hc2594565, 32'h42997b67, 32'hc254ee4f, 32'hc20bd3c5, 32'hc27aec5c, 32'hc17043b0};
test_output[25336:25343] = '{32'h0, 32'h42a8eb07, 32'h0, 32'h42997b67, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25344:25351] = '{32'h42502be7, 32'h424af5ce, 32'hc2ad159b, 32'h42578162, 32'h425e4dc1, 32'h428a33a2, 32'h42146922, 32'h42ac5fa1};
test_output[25344:25351] = '{32'h42502be7, 32'h424af5ce, 32'h0, 32'h42578162, 32'h425e4dc1, 32'h428a33a2, 32'h42146922, 32'h42ac5fa1};
test_input[25352:25359] = '{32'h421ba628, 32'h42151f9b, 32'h42ab97d9, 32'hc2a41f07, 32'h4282b6c7, 32'h419058d1, 32'h4247be9e, 32'h3fd6b248};
test_output[25352:25359] = '{32'h421ba628, 32'h42151f9b, 32'h42ab97d9, 32'h0, 32'h4282b6c7, 32'h419058d1, 32'h4247be9e, 32'h3fd6b248};
test_input[25360:25367] = '{32'h40b19887, 32'h4207ce00, 32'h4231c771, 32'h41eac7a6, 32'hc15d232b, 32'h42651250, 32'h42612eda, 32'hc1866985};
test_output[25360:25367] = '{32'h40b19887, 32'h4207ce00, 32'h4231c771, 32'h41eac7a6, 32'h0, 32'h42651250, 32'h42612eda, 32'h0};
test_input[25368:25375] = '{32'hc2be8edf, 32'h41f1794d, 32'h4298c68e, 32'h4171a1ae, 32'h421a8503, 32'hc1f968d0, 32'hc04b49d5, 32'h42061546};
test_output[25368:25375] = '{32'h0, 32'h41f1794d, 32'h4298c68e, 32'h4171a1ae, 32'h421a8503, 32'h0, 32'h0, 32'h42061546};
test_input[25376:25383] = '{32'h3f1f9bfe, 32'hc1bc3bab, 32'h42aca19f, 32'hc1e2d1a4, 32'h42a89fbf, 32'h413d3b62, 32'hc1b075c2, 32'h4253c2fd};
test_output[25376:25383] = '{32'h3f1f9bfe, 32'h0, 32'h42aca19f, 32'h0, 32'h42a89fbf, 32'h413d3b62, 32'h0, 32'h4253c2fd};
test_input[25384:25391] = '{32'hc2933344, 32'h413291f2, 32'hc250b5ab, 32'hc284d23f, 32'hc27f304e, 32'hc0c4a416, 32'h423f2343, 32'h42457bef};
test_output[25384:25391] = '{32'h0, 32'h413291f2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423f2343, 32'h42457bef};
test_input[25392:25399] = '{32'hc2babb25, 32'hc1e9d4ac, 32'hc117b0d7, 32'h4098111a, 32'hc17adb25, 32'h420d5958, 32'h42bd582d, 32'hc20f17d2};
test_output[25392:25399] = '{32'h0, 32'h0, 32'h0, 32'h4098111a, 32'h0, 32'h420d5958, 32'h42bd582d, 32'h0};
test_input[25400:25407] = '{32'hc242ff45, 32'hc2187a6d, 32'h4212d321, 32'hc2916d21, 32'hc225a9eb, 32'h427b6729, 32'hc2344a90, 32'h41d79b9a};
test_output[25400:25407] = '{32'h0, 32'h0, 32'h4212d321, 32'h0, 32'h0, 32'h427b6729, 32'h0, 32'h41d79b9a};
test_input[25408:25415] = '{32'h42bf4917, 32'hc2b7c051, 32'hc29be1dd, 32'hc1d5a3db, 32'h40493d72, 32'hc2a68b3f, 32'h41cefd08, 32'h4219fd9f};
test_output[25408:25415] = '{32'h42bf4917, 32'h0, 32'h0, 32'h0, 32'h40493d72, 32'h0, 32'h41cefd08, 32'h4219fd9f};
test_input[25416:25423] = '{32'hbd67b65c, 32'hc26c4500, 32'h3fc65efb, 32'hc1b006cb, 32'h42764043, 32'h428a5851, 32'h428832d3, 32'hc23d1cdf};
test_output[25416:25423] = '{32'h0, 32'h0, 32'h3fc65efb, 32'h0, 32'h42764043, 32'h428a5851, 32'h428832d3, 32'h0};
test_input[25424:25431] = '{32'h41a897fa, 32'hc26dc316, 32'hc274be54, 32'h429a9f1c, 32'h423f7506, 32'h42331018, 32'hc2079585, 32'h4198a58d};
test_output[25424:25431] = '{32'h41a897fa, 32'h0, 32'h0, 32'h429a9f1c, 32'h423f7506, 32'h42331018, 32'h0, 32'h4198a58d};
test_input[25432:25439] = '{32'h3fc0a82f, 32'hc1a574b9, 32'h42034a27, 32'h429ea162, 32'hc0306085, 32'hc0f0c8dd, 32'h4224bcd7, 32'h42684b0b};
test_output[25432:25439] = '{32'h3fc0a82f, 32'h0, 32'h42034a27, 32'h429ea162, 32'h0, 32'h0, 32'h4224bcd7, 32'h42684b0b};
test_input[25440:25447] = '{32'h423025f1, 32'hc280fa50, 32'h42454fe2, 32'hc29e43f0, 32'h4234bb37, 32'h42b4dac4, 32'hc2307aa3, 32'h4290ede1};
test_output[25440:25447] = '{32'h423025f1, 32'h0, 32'h42454fe2, 32'h0, 32'h4234bb37, 32'h42b4dac4, 32'h0, 32'h4290ede1};
test_input[25448:25455] = '{32'h42c796c4, 32'h42ad7acf, 32'hc2bcbe32, 32'h42349b97, 32'hc1a2adc1, 32'h420347b0, 32'h412edb2e, 32'h423f4f1f};
test_output[25448:25455] = '{32'h42c796c4, 32'h42ad7acf, 32'h0, 32'h42349b97, 32'h0, 32'h420347b0, 32'h412edb2e, 32'h423f4f1f};
test_input[25456:25463] = '{32'hc2ae890f, 32'h42662e5d, 32'hc21ae1b9, 32'hc2b018fa, 32'hc239d121, 32'hc25a708b, 32'h42234384, 32'h42448b7d};
test_output[25456:25463] = '{32'h0, 32'h42662e5d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42234384, 32'h42448b7d};
test_input[25464:25471] = '{32'hc2bb6bd1, 32'hc179db97, 32'h424e9ffd, 32'hc287f376, 32'hc1c4d6ca, 32'hc1bcad81, 32'h418b2765, 32'hc27b2081};
test_output[25464:25471] = '{32'h0, 32'h0, 32'h424e9ffd, 32'h0, 32'h0, 32'h0, 32'h418b2765, 32'h0};
test_input[25472:25479] = '{32'hc23531a9, 32'h40bea878, 32'h42876d73, 32'hc2208ccd, 32'hc10672dc, 32'hc2b0061b, 32'h42432207, 32'hc28e18c8};
test_output[25472:25479] = '{32'h0, 32'h40bea878, 32'h42876d73, 32'h0, 32'h0, 32'h0, 32'h42432207, 32'h0};
test_input[25480:25487] = '{32'h42c6e54c, 32'h42823624, 32'h4187527e, 32'h422593cf, 32'h4297cbc7, 32'hc1167edc, 32'h42c13e87, 32'hc29557a1};
test_output[25480:25487] = '{32'h42c6e54c, 32'h42823624, 32'h4187527e, 32'h422593cf, 32'h4297cbc7, 32'h0, 32'h42c13e87, 32'h0};
test_input[25488:25495] = '{32'h429a4b04, 32'h3d26955c, 32'hc2c015b6, 32'h421a1a37, 32'hc184c775, 32'h428a2223, 32'h420663ae, 32'hc2c1894f};
test_output[25488:25495] = '{32'h429a4b04, 32'h3d26955c, 32'h0, 32'h421a1a37, 32'h0, 32'h428a2223, 32'h420663ae, 32'h0};
test_input[25496:25503] = '{32'hc1af2e29, 32'hc2585742, 32'h4091ce25, 32'h4225fd26, 32'h42b652a3, 32'hc185c5b5, 32'h42749178, 32'h42af0aef};
test_output[25496:25503] = '{32'h0, 32'h0, 32'h4091ce25, 32'h4225fd26, 32'h42b652a3, 32'h0, 32'h42749178, 32'h42af0aef};
test_input[25504:25511] = '{32'h4273ef23, 32'hc27e2eaa, 32'hc1923e76, 32'h424bb06f, 32'h3f573b83, 32'h42ae3922, 32'h4206d24f, 32'h4204ab6f};
test_output[25504:25511] = '{32'h4273ef23, 32'h0, 32'h0, 32'h424bb06f, 32'h3f573b83, 32'h42ae3922, 32'h4206d24f, 32'h4204ab6f};
test_input[25512:25519] = '{32'h4250320d, 32'h4284ec06, 32'h41fc4ade, 32'h42a56f7d, 32'hc2860024, 32'h411d5fb0, 32'hbed59036, 32'h42682c84};
test_output[25512:25519] = '{32'h4250320d, 32'h4284ec06, 32'h41fc4ade, 32'h42a56f7d, 32'h0, 32'h411d5fb0, 32'h0, 32'h42682c84};
test_input[25520:25527] = '{32'hc2bdd5ac, 32'hc2b73021, 32'h429dd05f, 32'hc19c8578, 32'hc248ac5c, 32'h428c5597, 32'hc29f8541, 32'h41285886};
test_output[25520:25527] = '{32'h0, 32'h0, 32'h429dd05f, 32'h0, 32'h0, 32'h428c5597, 32'h0, 32'h41285886};
test_input[25528:25535] = '{32'hc290c048, 32'hc0bc5383, 32'h4283d35b, 32'hbf7ac9dd, 32'hc16b6ac2, 32'h420a0c82, 32'hc1de32ab, 32'h41e4be88};
test_output[25528:25535] = '{32'h0, 32'h0, 32'h4283d35b, 32'h0, 32'h0, 32'h420a0c82, 32'h0, 32'h41e4be88};
test_input[25536:25543] = '{32'hc099d63a, 32'hc28d5658, 32'hc28d9586, 32'h4257d5b9, 32'hc2c08ce7, 32'hc0ebe991, 32'hc21885af, 32'h412e3348};
test_output[25536:25543] = '{32'h0, 32'h0, 32'h0, 32'h4257d5b9, 32'h0, 32'h0, 32'h0, 32'h412e3348};
test_input[25544:25551] = '{32'h428d4656, 32'hc1e7eccf, 32'hc161b067, 32'h41859f2d, 32'hc23e5b16, 32'hc22c002c, 32'h42373cf9, 32'hc1e65663};
test_output[25544:25551] = '{32'h428d4656, 32'h0, 32'h0, 32'h41859f2d, 32'h0, 32'h0, 32'h42373cf9, 32'h0};
test_input[25552:25559] = '{32'hc2695059, 32'hc1817146, 32'hbf08fd22, 32'h42c21306, 32'h42a3cebf, 32'h42a86097, 32'hc2228fad, 32'hc1441837};
test_output[25552:25559] = '{32'h0, 32'h0, 32'h0, 32'h42c21306, 32'h42a3cebf, 32'h42a86097, 32'h0, 32'h0};
test_input[25560:25567] = '{32'hc1bda7d0, 32'hc28a99af, 32'hc29dc2e3, 32'h42826af5, 32'hc0ee4408, 32'h41e5deb6, 32'hc20e404c, 32'h41e30d2a};
test_output[25560:25567] = '{32'h0, 32'h0, 32'h0, 32'h42826af5, 32'h0, 32'h41e5deb6, 32'h0, 32'h41e30d2a};
test_input[25568:25575] = '{32'h42b5b270, 32'hc24a182a, 32'hc0db291b, 32'h41ed5ddd, 32'hc02c1c91, 32'hc252a0b8, 32'h41553e7e, 32'h42a8b413};
test_output[25568:25575] = '{32'h42b5b270, 32'h0, 32'h0, 32'h41ed5ddd, 32'h0, 32'h0, 32'h41553e7e, 32'h42a8b413};
test_input[25576:25583] = '{32'hc1d2eddc, 32'hc1d8f189, 32'hc2872a4d, 32'hc0a34cf3, 32'h418dcf6b, 32'hc1e1ea5e, 32'hc25ed17b, 32'hc1a89121};
test_output[25576:25583] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h418dcf6b, 32'h0, 32'h0, 32'h0};
test_input[25584:25591] = '{32'hc1185444, 32'h41112a84, 32'hc2bbaf40, 32'h42a782d9, 32'hc246f6d9, 32'h41af382e, 32'hc2833163, 32'hc2a79666};
test_output[25584:25591] = '{32'h0, 32'h41112a84, 32'h0, 32'h42a782d9, 32'h0, 32'h41af382e, 32'h0, 32'h0};
test_input[25592:25599] = '{32'hc27daa51, 32'hc2950805, 32'hc2c15300, 32'h42b5df66, 32'hc205f2b4, 32'hc1fc05ec, 32'hc206fd83, 32'h429579a3};
test_output[25592:25599] = '{32'h0, 32'h0, 32'h0, 32'h42b5df66, 32'h0, 32'h0, 32'h0, 32'h429579a3};
test_input[25600:25607] = '{32'hc0bdd330, 32'h4218f77e, 32'hc0d66979, 32'h4286c0b8, 32'h4233467b, 32'h4264680a, 32'h41952729, 32'hc00b34cb};
test_output[25600:25607] = '{32'h0, 32'h4218f77e, 32'h0, 32'h4286c0b8, 32'h4233467b, 32'h4264680a, 32'h41952729, 32'h0};
test_input[25608:25615] = '{32'hc1058090, 32'hc13bb7e4, 32'h41b6d766, 32'hc27fa62b, 32'h42a40902, 32'h4144a2da, 32'h42118440, 32'hc29ced89};
test_output[25608:25615] = '{32'h0, 32'h0, 32'h41b6d766, 32'h0, 32'h42a40902, 32'h4144a2da, 32'h42118440, 32'h0};
test_input[25616:25623] = '{32'h41cd9e31, 32'h429fdb51, 32'h422dbd27, 32'hc2820128, 32'hc201b194, 32'hc10e5880, 32'hc26c1413, 32'h427d9990};
test_output[25616:25623] = '{32'h41cd9e31, 32'h429fdb51, 32'h422dbd27, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427d9990};
test_input[25624:25631] = '{32'h4233627a, 32'hc10baeba, 32'h42b4ca88, 32'hc2aff1f7, 32'hc224ea5e, 32'h410161f8, 32'hc2a4f0af, 32'hc28828b1};
test_output[25624:25631] = '{32'h4233627a, 32'h0, 32'h42b4ca88, 32'h0, 32'h0, 32'h410161f8, 32'h0, 32'h0};
test_input[25632:25639] = '{32'h40e1364f, 32'hbfe421ce, 32'h42729c0c, 32'hc21fb930, 32'h429d8075, 32'h42c1a4a0, 32'hc2aae8b8, 32'h4287ff74};
test_output[25632:25639] = '{32'h40e1364f, 32'h0, 32'h42729c0c, 32'h0, 32'h429d8075, 32'h42c1a4a0, 32'h0, 32'h4287ff74};
test_input[25640:25647] = '{32'h42af9de1, 32'hbf7bc230, 32'hc2890cec, 32'h425623d1, 32'h42c7936b, 32'hc2a88f50, 32'hc0f3d89e, 32'h426595f2};
test_output[25640:25647] = '{32'h42af9de1, 32'h0, 32'h0, 32'h425623d1, 32'h42c7936b, 32'h0, 32'h0, 32'h426595f2};
test_input[25648:25655] = '{32'hc2423aff, 32'h4292ccc9, 32'hc2b68df4, 32'h42a4535a, 32'hc2bd47a7, 32'h42298835, 32'h426f87a2, 32'h414ea70b};
test_output[25648:25655] = '{32'h0, 32'h4292ccc9, 32'h0, 32'h42a4535a, 32'h0, 32'h42298835, 32'h426f87a2, 32'h414ea70b};
test_input[25656:25663] = '{32'hc2a751c1, 32'h424b04ee, 32'h4284d2c4, 32'hc2241aa9, 32'h4159bcca, 32'h42034b77, 32'hc1b0d960, 32'h40d1cd2c};
test_output[25656:25663] = '{32'h0, 32'h424b04ee, 32'h4284d2c4, 32'h0, 32'h4159bcca, 32'h42034b77, 32'h0, 32'h40d1cd2c};
test_input[25664:25671] = '{32'h41392e98, 32'hc1f74bab, 32'hc2366370, 32'h41a29002, 32'h42be046b, 32'hc14be4ae, 32'hc29061e7, 32'hc29ea9b7};
test_output[25664:25671] = '{32'h41392e98, 32'h0, 32'h0, 32'h41a29002, 32'h42be046b, 32'h0, 32'h0, 32'h0};
test_input[25672:25679] = '{32'hc2185328, 32'h41e016a3, 32'hc25fd570, 32'hc246a3da, 32'hc2ab0ef0, 32'h4209bf18, 32'h42b75bed, 32'h4107112f};
test_output[25672:25679] = '{32'h0, 32'h41e016a3, 32'h0, 32'h0, 32'h0, 32'h4209bf18, 32'h42b75bed, 32'h4107112f};
test_input[25680:25687] = '{32'hc296ee94, 32'hc2bcf024, 32'hc1271db7, 32'h42a991d0, 32'hc20d2416, 32'h41e486e3, 32'h42019de0, 32'hc27ea8fa};
test_output[25680:25687] = '{32'h0, 32'h0, 32'h0, 32'h42a991d0, 32'h0, 32'h41e486e3, 32'h42019de0, 32'h0};
test_input[25688:25695] = '{32'hc1dea61e, 32'hc2b6f65a, 32'h3efee890, 32'hc2c2d50d, 32'h41c2e40b, 32'hc2128555, 32'h428e61da, 32'h42a5a2c8};
test_output[25688:25695] = '{32'h0, 32'h0, 32'h3efee890, 32'h0, 32'h41c2e40b, 32'h0, 32'h428e61da, 32'h42a5a2c8};
test_input[25696:25703] = '{32'hc238bc57, 32'hc21dea77, 32'h41b3aa16, 32'h42a162fc, 32'hc2149945, 32'h42130bac, 32'hc0ede914, 32'h419845e4};
test_output[25696:25703] = '{32'h0, 32'h0, 32'h41b3aa16, 32'h42a162fc, 32'h0, 32'h42130bac, 32'h0, 32'h419845e4};
test_input[25704:25711] = '{32'h42b75c5a, 32'hc1b33f6a, 32'hc27287aa, 32'hc254c67d, 32'h429f8b88, 32'hc2c085be, 32'h42b5b427, 32'h414ec759};
test_output[25704:25711] = '{32'h42b75c5a, 32'h0, 32'h0, 32'h0, 32'h429f8b88, 32'h0, 32'h42b5b427, 32'h414ec759};
test_input[25712:25719] = '{32'hc2bbde16, 32'hc29488ec, 32'h42bc9fc4, 32'hc299c079, 32'hc16a0dfd, 32'h42567e9f, 32'h423c93eb, 32'hc227c019};
test_output[25712:25719] = '{32'h0, 32'h0, 32'h42bc9fc4, 32'h0, 32'h0, 32'h42567e9f, 32'h423c93eb, 32'h0};
test_input[25720:25727] = '{32'h41aca80e, 32'h4296a99c, 32'h4279a017, 32'hc2078c51, 32'h4253d6ef, 32'h41820118, 32'hc2c3a041, 32'hc277223c};
test_output[25720:25727] = '{32'h41aca80e, 32'h4296a99c, 32'h4279a017, 32'h0, 32'h4253d6ef, 32'h41820118, 32'h0, 32'h0};
test_input[25728:25735] = '{32'hc1dedc39, 32'h42851d5f, 32'h4282a0ab, 32'hc26196a3, 32'h41518926, 32'hc20c7d6b, 32'hc2baf058, 32'h4123baf1};
test_output[25728:25735] = '{32'h0, 32'h42851d5f, 32'h4282a0ab, 32'h0, 32'h41518926, 32'h0, 32'h0, 32'h4123baf1};
test_input[25736:25743] = '{32'h429591cf, 32'hc2bfa1c5, 32'h42272e9d, 32'hc1ab5dba, 32'hc2912c11, 32'hc2a7f283, 32'h42373719, 32'hc0dad17b};
test_output[25736:25743] = '{32'h429591cf, 32'h0, 32'h42272e9d, 32'h0, 32'h0, 32'h0, 32'h42373719, 32'h0};
test_input[25744:25751] = '{32'hc25e1e5e, 32'h42ba821d, 32'h42c26d6f, 32'hc1a491e2, 32'hc29e8d3b, 32'h425f1955, 32'h42a968c5, 32'hc183ded8};
test_output[25744:25751] = '{32'h0, 32'h42ba821d, 32'h42c26d6f, 32'h0, 32'h0, 32'h425f1955, 32'h42a968c5, 32'h0};
test_input[25752:25759] = '{32'h4201d697, 32'hc2367b80, 32'h41bc96d1, 32'hc180a6d9, 32'h42825c71, 32'h419d7526, 32'hc2b9b02c, 32'h4234d0ea};
test_output[25752:25759] = '{32'h4201d697, 32'h0, 32'h41bc96d1, 32'h0, 32'h42825c71, 32'h419d7526, 32'h0, 32'h4234d0ea};
test_input[25760:25767] = '{32'hc1c4979c, 32'h419dc319, 32'hc248ccc8, 32'hc262cd95, 32'h41ac706f, 32'hc290709e, 32'hc1918f9d, 32'hc14805ec};
test_output[25760:25767] = '{32'h0, 32'h419dc319, 32'h0, 32'h0, 32'h41ac706f, 32'h0, 32'h0, 32'h0};
test_input[25768:25775] = '{32'h42792a56, 32'h42339c8a, 32'hc2ae25d9, 32'h41fbd1ab, 32'h4204ae19, 32'hc1cf3fc1, 32'hc28aac08, 32'h42bba6ea};
test_output[25768:25775] = '{32'h42792a56, 32'h42339c8a, 32'h0, 32'h41fbd1ab, 32'h4204ae19, 32'h0, 32'h0, 32'h42bba6ea};
test_input[25776:25783] = '{32'hc2661052, 32'h421ec12d, 32'h41e3ac2a, 32'h4254861d, 32'hc2b803b8, 32'h41e81a3b, 32'h41289be8, 32'hc267f939};
test_output[25776:25783] = '{32'h0, 32'h421ec12d, 32'h41e3ac2a, 32'h4254861d, 32'h0, 32'h41e81a3b, 32'h41289be8, 32'h0};
test_input[25784:25791] = '{32'h3fd47a9d, 32'hc246ee1d, 32'hc28d4f1a, 32'h40f4c26e, 32'hc28acd9c, 32'hc2788a66, 32'hc1ba18f0, 32'h42854453};
test_output[25784:25791] = '{32'h3fd47a9d, 32'h0, 32'h0, 32'h40f4c26e, 32'h0, 32'h0, 32'h0, 32'h42854453};
test_input[25792:25799] = '{32'hc28c6f4d, 32'h42bf7b21, 32'hc281c984, 32'h4282ebf8, 32'hc1c2b4f3, 32'h42346c14, 32'h429a1ed7, 32'h42b35e8d};
test_output[25792:25799] = '{32'h0, 32'h42bf7b21, 32'h0, 32'h4282ebf8, 32'h0, 32'h42346c14, 32'h429a1ed7, 32'h42b35e8d};
test_input[25800:25807] = '{32'h42b06ea3, 32'hc18c36cc, 32'h420df885, 32'h42b55f18, 32'h42b100f7, 32'h417d4031, 32'h42a7bf56, 32'h42a18e44};
test_output[25800:25807] = '{32'h42b06ea3, 32'h0, 32'h420df885, 32'h42b55f18, 32'h42b100f7, 32'h417d4031, 32'h42a7bf56, 32'h42a18e44};
test_input[25808:25815] = '{32'hc28bae76, 32'hc204e588, 32'hc2a7ea33, 32'hc2371908, 32'h4284f502, 32'h42443130, 32'h4250cda5, 32'h41bd16e5};
test_output[25808:25815] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4284f502, 32'h42443130, 32'h4250cda5, 32'h41bd16e5};
test_input[25816:25823] = '{32'h42154062, 32'h424cc158, 32'hc2419c99, 32'hc1a14616, 32'h428b3c5d, 32'hc0c3f97b, 32'hc22dfa92, 32'hc1dc1f68};
test_output[25816:25823] = '{32'h42154062, 32'h424cc158, 32'h0, 32'h0, 32'h428b3c5d, 32'h0, 32'h0, 32'h0};
test_input[25824:25831] = '{32'hc2a368b7, 32'h42863162, 32'hc21ef380, 32'hc232d3b5, 32'h428bf096, 32'hbea4dd5b, 32'h42419e68, 32'h425706c6};
test_output[25824:25831] = '{32'h0, 32'h42863162, 32'h0, 32'h0, 32'h428bf096, 32'h0, 32'h42419e68, 32'h425706c6};
test_input[25832:25839] = '{32'hc286d90a, 32'hc27f14da, 32'hc28692ea, 32'h42496a5b, 32'h412c6287, 32'h41b69c53, 32'h4245b443, 32'h424b8603};
test_output[25832:25839] = '{32'h0, 32'h0, 32'h0, 32'h42496a5b, 32'h412c6287, 32'h41b69c53, 32'h4245b443, 32'h424b8603};
test_input[25840:25847] = '{32'hc28e5514, 32'hc29272bb, 32'h42b442c4, 32'h423b789b, 32'hc19a54d2, 32'hc2a29032, 32'h42b11168, 32'hc26fbd2f};
test_output[25840:25847] = '{32'h0, 32'h0, 32'h42b442c4, 32'h423b789b, 32'h0, 32'h0, 32'h42b11168, 32'h0};
test_input[25848:25855] = '{32'hc0d9403c, 32'hc183937a, 32'h4244335b, 32'hc1c46e5a, 32'h42245529, 32'h4208f84a, 32'hc154a119, 32'hc12b0f81};
test_output[25848:25855] = '{32'h0, 32'h0, 32'h4244335b, 32'h0, 32'h42245529, 32'h4208f84a, 32'h0, 32'h0};
test_input[25856:25863] = '{32'hc284869d, 32'hc1cdfee6, 32'h4263d8e4, 32'hc2a8f65c, 32'h42949920, 32'hc136c522, 32'h424d3c94, 32'hc1a77d47};
test_output[25856:25863] = '{32'h0, 32'h0, 32'h4263d8e4, 32'h0, 32'h42949920, 32'h0, 32'h424d3c94, 32'h0};
test_input[25864:25871] = '{32'h421c21d1, 32'hc250ca9d, 32'h413d0157, 32'h427285af, 32'h3ffd0b49, 32'h42993bdc, 32'hc1533cfe, 32'h4261a7f0};
test_output[25864:25871] = '{32'h421c21d1, 32'h0, 32'h413d0157, 32'h427285af, 32'h3ffd0b49, 32'h42993bdc, 32'h0, 32'h4261a7f0};
test_input[25872:25879] = '{32'h413177f5, 32'h4009ac3b, 32'h42aaeb34, 32'h421ff852, 32'h42bcf997, 32'h41d51673, 32'h42ad2e19, 32'h42a2b8c1};
test_output[25872:25879] = '{32'h413177f5, 32'h4009ac3b, 32'h42aaeb34, 32'h421ff852, 32'h42bcf997, 32'h41d51673, 32'h42ad2e19, 32'h42a2b8c1};
test_input[25880:25887] = '{32'hc1ddd5ed, 32'h41dccff4, 32'hc1d7a55d, 32'hc1c689c0, 32'hc1111a4d, 32'hc1d353ae, 32'hc23fc135, 32'hc263a34c};
test_output[25880:25887] = '{32'h0, 32'h41dccff4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[25888:25895] = '{32'hc2969e21, 32'hc2a98e0c, 32'hc1cbe674, 32'h41d1190b, 32'h421831a9, 32'hc23f0ef3, 32'hc2053e56, 32'h42b3812b};
test_output[25888:25895] = '{32'h0, 32'h0, 32'h0, 32'h41d1190b, 32'h421831a9, 32'h0, 32'h0, 32'h42b3812b};
test_input[25896:25903] = '{32'hc2699b64, 32'hc2319924, 32'hc1a8bc8f, 32'hc1d7a1ac, 32'hc2aeeba4, 32'hc295e192, 32'hc28c9dcf, 32'h4220ef42};
test_output[25896:25903] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4220ef42};
test_input[25904:25911] = '{32'h427bc69a, 32'h42651247, 32'h4229347b, 32'h42af8f26, 32'hc23a36f6, 32'h4295e275, 32'h429b1ae7, 32'h42adeb5c};
test_output[25904:25911] = '{32'h427bc69a, 32'h42651247, 32'h4229347b, 32'h42af8f26, 32'h0, 32'h4295e275, 32'h429b1ae7, 32'h42adeb5c};
test_input[25912:25919] = '{32'hc17f4746, 32'hc2823d1a, 32'hc2aa158c, 32'h42791ce9, 32'hc100b1c0, 32'h41f475e1, 32'h423a30a8, 32'h41514ade};
test_output[25912:25919] = '{32'h0, 32'h0, 32'h0, 32'h42791ce9, 32'h0, 32'h41f475e1, 32'h423a30a8, 32'h41514ade};
test_input[25920:25927] = '{32'hc1e0254f, 32'hc2a127e4, 32'hc20c29ba, 32'hc2954035, 32'h413f99ef, 32'hc1d56418, 32'hc201d18f, 32'h42a14300};
test_output[25920:25927] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h413f99ef, 32'h0, 32'h0, 32'h42a14300};
test_input[25928:25935] = '{32'hc0637090, 32'hc20590f8, 32'h422208cf, 32'hc211aed1, 32'hc0acb5dc, 32'h42837c92, 32'h42bed935, 32'hc18f6c7e};
test_output[25928:25935] = '{32'h0, 32'h0, 32'h422208cf, 32'h0, 32'h0, 32'h42837c92, 32'h42bed935, 32'h0};
test_input[25936:25943] = '{32'h429e0af0, 32'hc1e49a60, 32'hc02f5d88, 32'hc2b1cbb8, 32'h41cf8b6b, 32'hc247f596, 32'hc28b8e97, 32'h410734ea};
test_output[25936:25943] = '{32'h429e0af0, 32'h0, 32'h0, 32'h0, 32'h41cf8b6b, 32'h0, 32'h0, 32'h410734ea};
test_input[25944:25951] = '{32'h4292aadb, 32'h4122cbb8, 32'h41d5dd60, 32'h42bd4de2, 32'h42a98ab0, 32'hc29de9aa, 32'hc29d8a98, 32'h4221c69b};
test_output[25944:25951] = '{32'h4292aadb, 32'h4122cbb8, 32'h41d5dd60, 32'h42bd4de2, 32'h42a98ab0, 32'h0, 32'h0, 32'h4221c69b};
test_input[25952:25959] = '{32'h42690328, 32'h426ce6d1, 32'h42a87361, 32'hc2654ad5, 32'hc27c562e, 32'hc1ca6207, 32'hc20cd0a5, 32'h429b9e59};
test_output[25952:25959] = '{32'h42690328, 32'h426ce6d1, 32'h42a87361, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429b9e59};
test_input[25960:25967] = '{32'h42b52b0b, 32'h42676a91, 32'h421c2491, 32'hc19a12e8, 32'h419a27ad, 32'hc2ab72c6, 32'h428cf756, 32'hbf896cab};
test_output[25960:25967] = '{32'h42b52b0b, 32'h42676a91, 32'h421c2491, 32'h0, 32'h419a27ad, 32'h0, 32'h428cf756, 32'h0};
test_input[25968:25975] = '{32'hc278a285, 32'h42a54209, 32'hc1372cfb, 32'hc2957420, 32'h4186294e, 32'h42c15184, 32'h4203cee8, 32'h427c0fc2};
test_output[25968:25975] = '{32'h0, 32'h42a54209, 32'h0, 32'h0, 32'h4186294e, 32'h42c15184, 32'h4203cee8, 32'h427c0fc2};
test_input[25976:25983] = '{32'hc052f32f, 32'hc1c81862, 32'h417e1949, 32'h42289443, 32'h4210f61d, 32'h42a59f4f, 32'h41a1bc31, 32'hc21a7ba0};
test_output[25976:25983] = '{32'h0, 32'h0, 32'h417e1949, 32'h42289443, 32'h4210f61d, 32'h42a59f4f, 32'h41a1bc31, 32'h0};
test_input[25984:25991] = '{32'h425e2893, 32'h41d31f0c, 32'h42225f89, 32'h41d05f2f, 32'h422b456d, 32'hc25e6179, 32'h42118102, 32'hc1a9f67c};
test_output[25984:25991] = '{32'h425e2893, 32'h41d31f0c, 32'h42225f89, 32'h41d05f2f, 32'h422b456d, 32'h0, 32'h42118102, 32'h0};
test_input[25992:25999] = '{32'hc29487d1, 32'hc280dff4, 32'hc22229a6, 32'h41fd2730, 32'h4248875a, 32'h42a27fe5, 32'hc1fd0c36, 32'hc1aeba9d};
test_output[25992:25999] = '{32'h0, 32'h0, 32'h0, 32'h41fd2730, 32'h4248875a, 32'h42a27fe5, 32'h0, 32'h0};
test_input[26000:26007] = '{32'h428f3bac, 32'h4277e0ee, 32'h4243355c, 32'h41953206, 32'hc20e7ad9, 32'hc06d163e, 32'hc16013c5, 32'hc067274e};
test_output[26000:26007] = '{32'h428f3bac, 32'h4277e0ee, 32'h4243355c, 32'h41953206, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26008:26015] = '{32'hc2045510, 32'h41bb0910, 32'hc29024b4, 32'hc298f2d4, 32'hc1ee8b83, 32'h4226c2ea, 32'hc26b7e96, 32'h4168f817};
test_output[26008:26015] = '{32'h0, 32'h41bb0910, 32'h0, 32'h0, 32'h0, 32'h4226c2ea, 32'h0, 32'h4168f817};
test_input[26016:26023] = '{32'hc184a3a6, 32'h409684cf, 32'h42a68b8b, 32'hc2ac06d2, 32'hc1fdbbec, 32'h42afa6eb, 32'h42889864, 32'hc2afc351};
test_output[26016:26023] = '{32'h0, 32'h409684cf, 32'h42a68b8b, 32'h0, 32'h0, 32'h42afa6eb, 32'h42889864, 32'h0};
test_input[26024:26031] = '{32'h42a03ccb, 32'hc2abf3e6, 32'h42982025, 32'h4154a691, 32'h4212d786, 32'hc290f319, 32'h41a17163, 32'hc2a8c586};
test_output[26024:26031] = '{32'h42a03ccb, 32'h0, 32'h42982025, 32'h4154a691, 32'h4212d786, 32'h0, 32'h41a17163, 32'h0};
test_input[26032:26039] = '{32'h42480f39, 32'hc2860d05, 32'hc1d597c4, 32'h42bce559, 32'h423113ac, 32'h40d8c55b, 32'hc29ec416, 32'hc19997ab};
test_output[26032:26039] = '{32'h42480f39, 32'h0, 32'h0, 32'h42bce559, 32'h423113ac, 32'h40d8c55b, 32'h0, 32'h0};
test_input[26040:26047] = '{32'hc2a9e548, 32'hc0f50c3a, 32'h423a5333, 32'h426f1d53, 32'hc2856f66, 32'h42b8a2d5, 32'hc2bbb43b, 32'h4224a303};
test_output[26040:26047] = '{32'h0, 32'h0, 32'h423a5333, 32'h426f1d53, 32'h0, 32'h42b8a2d5, 32'h0, 32'h4224a303};
test_input[26048:26055] = '{32'hc224f6e9, 32'hc2af5e13, 32'h42555911, 32'h411f90e4, 32'hc25dc758, 32'h414f3ce8, 32'hc24b23ed, 32'hc22febcd};
test_output[26048:26055] = '{32'h0, 32'h0, 32'h42555911, 32'h411f90e4, 32'h0, 32'h414f3ce8, 32'h0, 32'h0};
test_input[26056:26063] = '{32'h3fa163a1, 32'h41f05045, 32'h42bf71bb, 32'hc2718f72, 32'hc2c29ba5, 32'h421eca4a, 32'hc2b6ba84, 32'h4215e6ad};
test_output[26056:26063] = '{32'h3fa163a1, 32'h41f05045, 32'h42bf71bb, 32'h0, 32'h0, 32'h421eca4a, 32'h0, 32'h4215e6ad};
test_input[26064:26071] = '{32'hc27efd23, 32'hc1c8fab3, 32'hc295f6b2, 32'hc28d09fb, 32'hc19d4873, 32'hc1a8ed84, 32'hc291d389, 32'hc2800ab0};
test_output[26064:26071] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26072:26079] = '{32'h4190c975, 32'hc2be80ef, 32'h4130bbaf, 32'hc21cdfc2, 32'hc112ea4a, 32'hc28564e6, 32'h4235d980, 32'hc1fcaa6c};
test_output[26072:26079] = '{32'h4190c975, 32'h0, 32'h4130bbaf, 32'h0, 32'h0, 32'h0, 32'h4235d980, 32'h0};
test_input[26080:26087] = '{32'h4105a49a, 32'hc09d9c3d, 32'hc2718d1b, 32'hc2bcb409, 32'h4181b21f, 32'hc14ce582, 32'h428d521b, 32'hc29d20db};
test_output[26080:26087] = '{32'h4105a49a, 32'h0, 32'h0, 32'h0, 32'h4181b21f, 32'h0, 32'h428d521b, 32'h0};
test_input[26088:26095] = '{32'h42804602, 32'hc24ae81d, 32'h4175df80, 32'hc2b4baf9, 32'h42b4eba7, 32'h42837eca, 32'hc1eed81f, 32'hc2b994ce};
test_output[26088:26095] = '{32'h42804602, 32'h0, 32'h4175df80, 32'h0, 32'h42b4eba7, 32'h42837eca, 32'h0, 32'h0};
test_input[26096:26103] = '{32'h428a5a13, 32'h41728939, 32'h416f6828, 32'h41b3f1d8, 32'hc294ee17, 32'h412bdd92, 32'hc293f436, 32'h4229712e};
test_output[26096:26103] = '{32'h428a5a13, 32'h41728939, 32'h416f6828, 32'h41b3f1d8, 32'h0, 32'h412bdd92, 32'h0, 32'h4229712e};
test_input[26104:26111] = '{32'h4274b8eb, 32'hc2a949cd, 32'h42c1276d, 32'h4250af28, 32'h4239ea14, 32'hc18330c6, 32'hc223c0eb, 32'hc239a0da};
test_output[26104:26111] = '{32'h4274b8eb, 32'h0, 32'h42c1276d, 32'h4250af28, 32'h4239ea14, 32'h0, 32'h0, 32'h0};
test_input[26112:26119] = '{32'h40111949, 32'hc22419dd, 32'hc179fd10, 32'hc1211e42, 32'h42c235cc, 32'h4202025c, 32'hc148d153, 32'hc2bf2565};
test_output[26112:26119] = '{32'h40111949, 32'h0, 32'h0, 32'h0, 32'h42c235cc, 32'h4202025c, 32'h0, 32'h0};
test_input[26120:26127] = '{32'hc29c7d69, 32'h428a8510, 32'h42042243, 32'hc10accf8, 32'h4278151a, 32'h41aabb25, 32'hc28d7980, 32'hc2b71056};
test_output[26120:26127] = '{32'h0, 32'h428a8510, 32'h42042243, 32'h0, 32'h4278151a, 32'h41aabb25, 32'h0, 32'h0};
test_input[26128:26135] = '{32'h4289333c, 32'h421d6b0e, 32'hc2bf8002, 32'hc2bbbe59, 32'hc2b96ef0, 32'h42c06887, 32'h41e03a57, 32'hc2113081};
test_output[26128:26135] = '{32'h4289333c, 32'h421d6b0e, 32'h0, 32'h0, 32'h0, 32'h42c06887, 32'h41e03a57, 32'h0};
test_input[26136:26143] = '{32'hc2c35f10, 32'hc0d168fb, 32'hc1e16014, 32'h42bf7a7f, 32'hc276a1d0, 32'h422f2bd0, 32'h4299b9cd, 32'hc2b88d94};
test_output[26136:26143] = '{32'h0, 32'h0, 32'h0, 32'h42bf7a7f, 32'h0, 32'h422f2bd0, 32'h4299b9cd, 32'h0};
test_input[26144:26151] = '{32'hc21710ee, 32'hc2c5a91f, 32'h42a98538, 32'hc2bc6197, 32'h429fc8de, 32'h40da4930, 32'hc1bbdd8d, 32'hc2506b96};
test_output[26144:26151] = '{32'h0, 32'h0, 32'h42a98538, 32'h0, 32'h429fc8de, 32'h40da4930, 32'h0, 32'h0};
test_input[26152:26159] = '{32'hc1d997c7, 32'hc0faf8d2, 32'h429d446c, 32'h42a2ef64, 32'h41e55313, 32'h42654d8e, 32'h4184c267, 32'h410bc42b};
test_output[26152:26159] = '{32'h0, 32'h0, 32'h429d446c, 32'h42a2ef64, 32'h41e55313, 32'h42654d8e, 32'h4184c267, 32'h410bc42b};
test_input[26160:26167] = '{32'hc2743702, 32'hc1841711, 32'hc23b8552, 32'hc216e085, 32'h42b67a98, 32'h40f8b0f4, 32'hc29c58e8, 32'h3e8d1e03};
test_output[26160:26167] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42b67a98, 32'h40f8b0f4, 32'h0, 32'h3e8d1e03};
test_input[26168:26175] = '{32'h42c1afe9, 32'h42b9ec69, 32'h42b16766, 32'hc2a2d444, 32'hc28b4816, 32'h415060db, 32'h42afb3c2, 32'h42665a5f};
test_output[26168:26175] = '{32'h42c1afe9, 32'h42b9ec69, 32'h42b16766, 32'h0, 32'h0, 32'h415060db, 32'h42afb3c2, 32'h42665a5f};
test_input[26176:26183] = '{32'hc1096c79, 32'hbf4ebf84, 32'h42c0cecf, 32'h41af2a58, 32'hc13b0631, 32'hc2506702, 32'h42ad4716, 32'h42acf56c};
test_output[26176:26183] = '{32'h0, 32'h0, 32'h42c0cecf, 32'h41af2a58, 32'h0, 32'h0, 32'h42ad4716, 32'h42acf56c};
test_input[26184:26191] = '{32'hc2c06c17, 32'h42103332, 32'hc2775a58, 32'hc10156e9, 32'h425562f1, 32'hc1d7975d, 32'hc1da4318, 32'h420e7c88};
test_output[26184:26191] = '{32'h0, 32'h42103332, 32'h0, 32'h0, 32'h425562f1, 32'h0, 32'h0, 32'h420e7c88};
test_input[26192:26199] = '{32'h41a99311, 32'hc21b06c7, 32'h428342a4, 32'h428c82d7, 32'hc18e52de, 32'hc2beaadd, 32'h42af45d4, 32'h4276354e};
test_output[26192:26199] = '{32'h41a99311, 32'h0, 32'h428342a4, 32'h428c82d7, 32'h0, 32'h0, 32'h42af45d4, 32'h4276354e};
test_input[26200:26207] = '{32'h42b37f68, 32'h42af0f67, 32'hc247a1bd, 32'hc298ac52, 32'hc140016f, 32'h42955893, 32'h41c162fc, 32'h42583107};
test_output[26200:26207] = '{32'h42b37f68, 32'h42af0f67, 32'h0, 32'h0, 32'h0, 32'h42955893, 32'h41c162fc, 32'h42583107};
test_input[26208:26215] = '{32'h4104c44e, 32'hc1296377, 32'h41f8f937, 32'h42a11b0f, 32'h42670f39, 32'h42b8cde6, 32'hc2839632, 32'hc29ebc99};
test_output[26208:26215] = '{32'h4104c44e, 32'h0, 32'h41f8f937, 32'h42a11b0f, 32'h42670f39, 32'h42b8cde6, 32'h0, 32'h0};
test_input[26216:26223] = '{32'hc00d7a5e, 32'hc2925a6b, 32'hc2c294d7, 32'hc0f41842, 32'h421e31f6, 32'h4190cda0, 32'hc219e71d, 32'hc2be73fe};
test_output[26216:26223] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h421e31f6, 32'h4190cda0, 32'h0, 32'h0};
test_input[26224:26231] = '{32'hc21cc3df, 32'hc292274f, 32'hc1cf1b79, 32'h425eca86, 32'h409a82da, 32'h42907381, 32'hc1af96b5, 32'hc0736c32};
test_output[26224:26231] = '{32'h0, 32'h0, 32'h0, 32'h425eca86, 32'h409a82da, 32'h42907381, 32'h0, 32'h0};
test_input[26232:26239] = '{32'hc1b0fdf1, 32'h4290e2bc, 32'hc203f307, 32'hbf720090, 32'h41688aea, 32'h42882b20, 32'h42ae5f56, 32'h4265bedf};
test_output[26232:26239] = '{32'h0, 32'h4290e2bc, 32'h0, 32'h0, 32'h41688aea, 32'h42882b20, 32'h42ae5f56, 32'h4265bedf};
test_input[26240:26247] = '{32'hc2805e4f, 32'h4231e9a0, 32'hc16b6271, 32'hc24bcd70, 32'hc295b2fc, 32'h4106b70b, 32'h413c7682, 32'hc247ab5f};
test_output[26240:26247] = '{32'h0, 32'h4231e9a0, 32'h0, 32'h0, 32'h0, 32'h4106b70b, 32'h413c7682, 32'h0};
test_input[26248:26255] = '{32'hc195a43f, 32'h42c0cdc6, 32'h409c3603, 32'hc1880fac, 32'h40c42c87, 32'hc10274f5, 32'hc2b53c72, 32'h42ba9165};
test_output[26248:26255] = '{32'h0, 32'h42c0cdc6, 32'h409c3603, 32'h0, 32'h40c42c87, 32'h0, 32'h0, 32'h42ba9165};
test_input[26256:26263] = '{32'h41adf4a4, 32'hc285d762, 32'hc222dad5, 32'hc2aacac3, 32'h42bad7e8, 32'h41a00ab9, 32'hc1dabbb9, 32'hc2936daf};
test_output[26256:26263] = '{32'h41adf4a4, 32'h0, 32'h0, 32'h0, 32'h42bad7e8, 32'h41a00ab9, 32'h0, 32'h0};
test_input[26264:26271] = '{32'hc17bdf4f, 32'hc11780d0, 32'hc2a09c49, 32'h42ae7583, 32'hc1422213, 32'hc095ae5b, 32'h42a26b1c, 32'hc205d654};
test_output[26264:26271] = '{32'h0, 32'h0, 32'h0, 32'h42ae7583, 32'h0, 32'h0, 32'h42a26b1c, 32'h0};
test_input[26272:26279] = '{32'h41d86f73, 32'h41a42d5e, 32'h4298b430, 32'hc2adf458, 32'hc29e6706, 32'hc2870b71, 32'h429fe84a, 32'hc1c4f012};
test_output[26272:26279] = '{32'h41d86f73, 32'h41a42d5e, 32'h4298b430, 32'h0, 32'h0, 32'h0, 32'h429fe84a, 32'h0};
test_input[26280:26287] = '{32'hc23a21aa, 32'hbfd9b9b4, 32'h42b6882d, 32'hc0b83241, 32'hc29dacd8, 32'h42168bd1, 32'h42c7a719, 32'h42c39514};
test_output[26280:26287] = '{32'h0, 32'h0, 32'h42b6882d, 32'h0, 32'h0, 32'h42168bd1, 32'h42c7a719, 32'h42c39514};
test_input[26288:26295] = '{32'hc293831c, 32'hc287b9c4, 32'h411a207f, 32'hc1a7da4d, 32'h4169e03a, 32'hc21f2e0d, 32'hc1704122, 32'h42324774};
test_output[26288:26295] = '{32'h0, 32'h0, 32'h411a207f, 32'h0, 32'h4169e03a, 32'h0, 32'h0, 32'h42324774};
test_input[26296:26303] = '{32'h4083e5a2, 32'hc20a6502, 32'hc179f1e5, 32'hc18a900a, 32'h4288880e, 32'h4229a69a, 32'h42663f41, 32'h42c6b8b0};
test_output[26296:26303] = '{32'h4083e5a2, 32'h0, 32'h0, 32'h0, 32'h4288880e, 32'h4229a69a, 32'h42663f41, 32'h42c6b8b0};
test_input[26304:26311] = '{32'hc2abc461, 32'hc1ad709e, 32'hc184e6f2, 32'hc27011b6, 32'hc21e91ac, 32'h409934b4, 32'hc2118b11, 32'hc2a8b00a};
test_output[26304:26311] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h409934b4, 32'h0, 32'h0};
test_input[26312:26319] = '{32'hc24f090d, 32'hc21023e6, 32'h42a6c49c, 32'h42337b75, 32'hc2bd9d2a, 32'hc292d83b, 32'h4255ea25, 32'h4262c96b};
test_output[26312:26319] = '{32'h0, 32'h0, 32'h42a6c49c, 32'h42337b75, 32'h0, 32'h0, 32'h4255ea25, 32'h4262c96b};
test_input[26320:26327] = '{32'hc226fd48, 32'h41e97c08, 32'hbff555f8, 32'hc23b91f0, 32'h420ad632, 32'h41231ae7, 32'h42b1df34, 32'h409b0e4e};
test_output[26320:26327] = '{32'h0, 32'h41e97c08, 32'h0, 32'h0, 32'h420ad632, 32'h41231ae7, 32'h42b1df34, 32'h409b0e4e};
test_input[26328:26335] = '{32'h42845571, 32'h42a17018, 32'hc2b18c99, 32'h41ce99c5, 32'hc2306f19, 32'h424897e5, 32'h4247f6d7, 32'h41a65837};
test_output[26328:26335] = '{32'h42845571, 32'h42a17018, 32'h0, 32'h41ce99c5, 32'h0, 32'h424897e5, 32'h4247f6d7, 32'h41a65837};
test_input[26336:26343] = '{32'hc213dbe9, 32'hc2ab8234, 32'h428d3bc6, 32'h42214aaa, 32'h424134c4, 32'h42ba00f1, 32'hc2bbb6cc, 32'h423ccc86};
test_output[26336:26343] = '{32'h0, 32'h0, 32'h428d3bc6, 32'h42214aaa, 32'h424134c4, 32'h42ba00f1, 32'h0, 32'h423ccc86};
test_input[26344:26351] = '{32'hc2c5b34c, 32'h41420a45, 32'h41e816eb, 32'h421e65ca, 32'h41efa712, 32'hbe83d41c, 32'hc18d3501, 32'hc1f2d2e9};
test_output[26344:26351] = '{32'h0, 32'h41420a45, 32'h41e816eb, 32'h421e65ca, 32'h41efa712, 32'h0, 32'h0, 32'h0};
test_input[26352:26359] = '{32'hc2012ffc, 32'hc1966235, 32'h427d68a8, 32'hc1f25c44, 32'h429e5455, 32'h42ad4036, 32'h418d51f4, 32'hc217b940};
test_output[26352:26359] = '{32'h0, 32'h0, 32'h427d68a8, 32'h0, 32'h429e5455, 32'h42ad4036, 32'h418d51f4, 32'h0};
test_input[26360:26367] = '{32'hc203079f, 32'hc1c5d61d, 32'hc1b7bc44, 32'hc26523ac, 32'h420e52d5, 32'h3fc27d06, 32'h42b8307f, 32'h428534e7};
test_output[26360:26367] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h420e52d5, 32'h3fc27d06, 32'h42b8307f, 32'h428534e7};
test_input[26368:26375] = '{32'h411d8a16, 32'hc1274352, 32'h4107975f, 32'h421c9c17, 32'hc1be080f, 32'hc29718bd, 32'h4242a159, 32'hc2669a76};
test_output[26368:26375] = '{32'h411d8a16, 32'h0, 32'h4107975f, 32'h421c9c17, 32'h0, 32'h0, 32'h4242a159, 32'h0};
test_input[26376:26383] = '{32'h42952a42, 32'hc205a0ee, 32'h415b4763, 32'hc24a95e2, 32'hc233b90d, 32'h422478bd, 32'h42593d8a, 32'h42660e16};
test_output[26376:26383] = '{32'h42952a42, 32'h0, 32'h415b4763, 32'h0, 32'h0, 32'h422478bd, 32'h42593d8a, 32'h42660e16};
test_input[26384:26391] = '{32'h41e97604, 32'h426bc792, 32'h42c2212c, 32'h42a2f5ad, 32'hc2a27198, 32'h42495717, 32'h41607f8b, 32'hc13c6fc5};
test_output[26384:26391] = '{32'h41e97604, 32'h426bc792, 32'h42c2212c, 32'h42a2f5ad, 32'h0, 32'h42495717, 32'h41607f8b, 32'h0};
test_input[26392:26399] = '{32'hc24bbd03, 32'hc29ab3ab, 32'hc27a0b7e, 32'h41d2b5ab, 32'hc1b88e8a, 32'h42578a97, 32'hc1b7a6d1, 32'hc208fbab};
test_output[26392:26399] = '{32'h0, 32'h0, 32'h0, 32'h41d2b5ab, 32'h0, 32'h42578a97, 32'h0, 32'h0};
test_input[26400:26407] = '{32'hc1b3ba05, 32'h426a3c69, 32'h415e30e1, 32'hc26e800c, 32'h41ec5c2b, 32'h42b56426, 32'hc2470730, 32'h4183945e};
test_output[26400:26407] = '{32'h0, 32'h426a3c69, 32'h415e30e1, 32'h0, 32'h41ec5c2b, 32'h42b56426, 32'h0, 32'h4183945e};
test_input[26408:26415] = '{32'h41c2970b, 32'hc2c47743, 32'hc2af45ef, 32'hc0617bdc, 32'hc18d6c22, 32'h42a8e86e, 32'h40312b37, 32'hc1e5781e};
test_output[26408:26415] = '{32'h41c2970b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a8e86e, 32'h40312b37, 32'h0};
test_input[26416:26423] = '{32'h42c70106, 32'h40d1a2e0, 32'h42bebb2c, 32'h42bf5e79, 32'h42173594, 32'h42c3ec7f, 32'hc14cf9ec, 32'h424f3e84};
test_output[26416:26423] = '{32'h42c70106, 32'h40d1a2e0, 32'h42bebb2c, 32'h42bf5e79, 32'h42173594, 32'h42c3ec7f, 32'h0, 32'h424f3e84};
test_input[26424:26431] = '{32'h42a4633d, 32'hc18d1692, 32'h42837788, 32'h41a1f005, 32'hc200c64f, 32'hc0f8ec18, 32'hc17109e5, 32'h429e4e76};
test_output[26424:26431] = '{32'h42a4633d, 32'h0, 32'h42837788, 32'h41a1f005, 32'h0, 32'h0, 32'h0, 32'h429e4e76};
test_input[26432:26439] = '{32'h427b4759, 32'h41b67a0f, 32'hc2aa077f, 32'h41e39996, 32'hc281e9e6, 32'hc2099b4e, 32'hc2782845, 32'h42c58d1a};
test_output[26432:26439] = '{32'h427b4759, 32'h41b67a0f, 32'h0, 32'h41e39996, 32'h0, 32'h0, 32'h0, 32'h42c58d1a};
test_input[26440:26447] = '{32'hc13f9f15, 32'h4228fff7, 32'hc07bf06a, 32'hc20b2ebb, 32'hc2a62e9e, 32'h41556856, 32'h419e323b, 32'h405f9598};
test_output[26440:26447] = '{32'h0, 32'h4228fff7, 32'h0, 32'h0, 32'h0, 32'h41556856, 32'h419e323b, 32'h405f9598};
test_input[26448:26455] = '{32'h4041f8b0, 32'h3ff4a366, 32'h422a2907, 32'hc1bd85c0, 32'h406e8920, 32'h41b23453, 32'hc200b854, 32'hc29721f6};
test_output[26448:26455] = '{32'h4041f8b0, 32'h3ff4a366, 32'h422a2907, 32'h0, 32'h406e8920, 32'h41b23453, 32'h0, 32'h0};
test_input[26456:26463] = '{32'h428435d4, 32'h42b59f6a, 32'hc1492193, 32'h428c683f, 32'h420b0e4a, 32'h41a75086, 32'hc0eb574b, 32'hc099cc21};
test_output[26456:26463] = '{32'h428435d4, 32'h42b59f6a, 32'h0, 32'h428c683f, 32'h420b0e4a, 32'h41a75086, 32'h0, 32'h0};
test_input[26464:26471] = '{32'h4250115b, 32'hc2beadd8, 32'h42bf0241, 32'h425f50f3, 32'hc19abd52, 32'h4262e4a6, 32'h4141375d, 32'h4105e60a};
test_output[26464:26471] = '{32'h4250115b, 32'h0, 32'h42bf0241, 32'h425f50f3, 32'h0, 32'h4262e4a6, 32'h4141375d, 32'h4105e60a};
test_input[26472:26479] = '{32'h42c697a5, 32'h428ca85d, 32'hc2bfc720, 32'hc1cfe9b0, 32'hc29f05d4, 32'hc05b57d2, 32'h41d698db, 32'hc165b264};
test_output[26472:26479] = '{32'h42c697a5, 32'h428ca85d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41d698db, 32'h0};
test_input[26480:26487] = '{32'h4282a509, 32'h4186d676, 32'hc2c40d2f, 32'hc27f275d, 32'h429b9148, 32'hc257d721, 32'h41cbfa55, 32'h42b83de5};
test_output[26480:26487] = '{32'h4282a509, 32'h4186d676, 32'h0, 32'h0, 32'h429b9148, 32'h0, 32'h41cbfa55, 32'h42b83de5};
test_input[26488:26495] = '{32'h4226c4a7, 32'h422153fc, 32'h42c05a8f, 32'hc2193103, 32'hc285c272, 32'h4014e2c5, 32'h41a34a6f, 32'hc15d7458};
test_output[26488:26495] = '{32'h4226c4a7, 32'h422153fc, 32'h42c05a8f, 32'h0, 32'h0, 32'h4014e2c5, 32'h41a34a6f, 32'h0};
test_input[26496:26503] = '{32'hc2c4e772, 32'h42bf8ca2, 32'h41f5ec92, 32'hc266e737, 32'hc0af6da9, 32'h4295583e, 32'hc1b176d0, 32'h422313e1};
test_output[26496:26503] = '{32'h0, 32'h42bf8ca2, 32'h41f5ec92, 32'h0, 32'h0, 32'h4295583e, 32'h0, 32'h422313e1};
test_input[26504:26511] = '{32'hc2b14452, 32'h42b56366, 32'hc29d3cfd, 32'hc2332ba7, 32'h41be8fe7, 32'h4290bc5e, 32'hc2bef98c, 32'h42581d8a};
test_output[26504:26511] = '{32'h0, 32'h42b56366, 32'h0, 32'h0, 32'h41be8fe7, 32'h4290bc5e, 32'h0, 32'h42581d8a};
test_input[26512:26519] = '{32'hc2c3b182, 32'hc2a35d41, 32'h4209de01, 32'hc24c535a, 32'h4248a5aa, 32'hc1a0ceaf, 32'h40a1060f, 32'hc2c3781b};
test_output[26512:26519] = '{32'h0, 32'h0, 32'h4209de01, 32'h0, 32'h4248a5aa, 32'h0, 32'h40a1060f, 32'h0};
test_input[26520:26527] = '{32'hc1da8d01, 32'hc29bc2ac, 32'hc1f2f53d, 32'hc25c6983, 32'h41cf506b, 32'h4202b84e, 32'h419ba67d, 32'h425c66c5};
test_output[26520:26527] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41cf506b, 32'h4202b84e, 32'h419ba67d, 32'h425c66c5};
test_input[26528:26535] = '{32'h42b4181b, 32'h419e615f, 32'hc2b22112, 32'hc21dac26, 32'h42781700, 32'hc1a44182, 32'h42a27858, 32'hc23718b9};
test_output[26528:26535] = '{32'h42b4181b, 32'h419e615f, 32'h0, 32'h0, 32'h42781700, 32'h0, 32'h42a27858, 32'h0};
test_input[26536:26543] = '{32'h4242afce, 32'hc0f096f0, 32'hc1ce7419, 32'h420e98e5, 32'hc2c0ffa3, 32'h42609006, 32'hc28d450c, 32'h422053b4};
test_output[26536:26543] = '{32'h4242afce, 32'h0, 32'h0, 32'h420e98e5, 32'h0, 32'h42609006, 32'h0, 32'h422053b4};
test_input[26544:26551] = '{32'h4228674b, 32'hc24dafd0, 32'h419fbd35, 32'h40a98e05, 32'hc24e9c97, 32'hc2725a64, 32'h42ab69db, 32'hc1a79531};
test_output[26544:26551] = '{32'h4228674b, 32'h0, 32'h419fbd35, 32'h40a98e05, 32'h0, 32'h0, 32'h42ab69db, 32'h0};
test_input[26552:26559] = '{32'h402254ce, 32'hc2313251, 32'h42c386aa, 32'h42b3b72a, 32'hc2af7df0, 32'hc2a0a9bc, 32'hc24b0728, 32'hc292ed5f};
test_output[26552:26559] = '{32'h402254ce, 32'h0, 32'h42c386aa, 32'h42b3b72a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26560:26567] = '{32'h42109990, 32'h426b4218, 32'hc12d0a39, 32'h426303aa, 32'hc11c4f03, 32'h42a43b19, 32'hc2c1d008, 32'h42544bca};
test_output[26560:26567] = '{32'h42109990, 32'h426b4218, 32'h0, 32'h426303aa, 32'h0, 32'h42a43b19, 32'h0, 32'h42544bca};
test_input[26568:26575] = '{32'hc27090bc, 32'h42ac3ed7, 32'h4294618e, 32'hc226d4b7, 32'h42957ba8, 32'h416dae55, 32'h421ffd4a, 32'hc29157b4};
test_output[26568:26575] = '{32'h0, 32'h42ac3ed7, 32'h4294618e, 32'h0, 32'h42957ba8, 32'h416dae55, 32'h421ffd4a, 32'h0};
test_input[26576:26583] = '{32'hc2323f1f, 32'hc20db2d1, 32'hc1bd06d5, 32'h4179d3b2, 32'h42682cb4, 32'h40b43528, 32'h428bebd6, 32'hc193d3fe};
test_output[26576:26583] = '{32'h0, 32'h0, 32'h0, 32'h4179d3b2, 32'h42682cb4, 32'h40b43528, 32'h428bebd6, 32'h0};
test_input[26584:26591] = '{32'hc2b5f166, 32'hc28740f2, 32'hc2656720, 32'h41e7b30b, 32'h4292f3b5, 32'h41a69acc, 32'hc2239879, 32'hc0d3eb63};
test_output[26584:26591] = '{32'h0, 32'h0, 32'h0, 32'h41e7b30b, 32'h4292f3b5, 32'h41a69acc, 32'h0, 32'h0};
test_input[26592:26599] = '{32'h40691117, 32'h4227d08d, 32'hc201d0ac, 32'hc208a04b, 32'hc28953fc, 32'h41359472, 32'h428e7984, 32'hc23d501d};
test_output[26592:26599] = '{32'h40691117, 32'h4227d08d, 32'h0, 32'h0, 32'h0, 32'h41359472, 32'h428e7984, 32'h0};
test_input[26600:26607] = '{32'h4257d72d, 32'h41c1f4a6, 32'h42a1bf7e, 32'hc2a3be3c, 32'hc21d1b5b, 32'hc0a3a59e, 32'h41e57777, 32'hc1f86a9c};
test_output[26600:26607] = '{32'h4257d72d, 32'h41c1f4a6, 32'h42a1bf7e, 32'h0, 32'h0, 32'h0, 32'h41e57777, 32'h0};
test_input[26608:26615] = '{32'h428f0a91, 32'h4135c860, 32'hc0e8a129, 32'h421c6de5, 32'hc2c0a06c, 32'h425d0f77, 32'hc130100d, 32'h41b50a48};
test_output[26608:26615] = '{32'h428f0a91, 32'h4135c860, 32'h0, 32'h421c6de5, 32'h0, 32'h425d0f77, 32'h0, 32'h41b50a48};
test_input[26616:26623] = '{32'h428abc87, 32'hc2c57d8d, 32'hc21714f6, 32'h42148d5f, 32'hc2947d2a, 32'hc294be0d, 32'hc2708317, 32'h41987251};
test_output[26616:26623] = '{32'h428abc87, 32'h0, 32'h0, 32'h42148d5f, 32'h0, 32'h0, 32'h0, 32'h41987251};
test_input[26624:26631] = '{32'hc03ec358, 32'h41890220, 32'h41f1ac4b, 32'hc2a92b09, 32'h42957b55, 32'h429691b8, 32'hc125f6bd, 32'h42c2ba0d};
test_output[26624:26631] = '{32'h0, 32'h41890220, 32'h41f1ac4b, 32'h0, 32'h42957b55, 32'h429691b8, 32'h0, 32'h42c2ba0d};
test_input[26632:26639] = '{32'hc211ce12, 32'h42af62a1, 32'hc14ed3c7, 32'h40737d17, 32'h40d7a3d0, 32'h42b0b45f, 32'h4189a879, 32'h42adaae2};
test_output[26632:26639] = '{32'h0, 32'h42af62a1, 32'h0, 32'h40737d17, 32'h40d7a3d0, 32'h42b0b45f, 32'h4189a879, 32'h42adaae2};
test_input[26640:26647] = '{32'h42a2acbb, 32'hc290f550, 32'h4295de2a, 32'hc217926b, 32'hc2adc34d, 32'h3eccbe35, 32'h41bb5b17, 32'hc16d4e3e};
test_output[26640:26647] = '{32'h42a2acbb, 32'h0, 32'h4295de2a, 32'h0, 32'h0, 32'h3eccbe35, 32'h41bb5b17, 32'h0};
test_input[26648:26655] = '{32'h428d76c4, 32'hc1357a3c, 32'hc29d372b, 32'h42a10ef5, 32'h429a5a04, 32'hbf8e4553, 32'hc28c1160, 32'hc25f34f1};
test_output[26648:26655] = '{32'h428d76c4, 32'h0, 32'h0, 32'h42a10ef5, 32'h429a5a04, 32'h0, 32'h0, 32'h0};
test_input[26656:26663] = '{32'h42b660de, 32'hc1d4c747, 32'h40fcbe13, 32'h400eb174, 32'h425c09f0, 32'h411ef49f, 32'h40b19e9e, 32'hc249a6f0};
test_output[26656:26663] = '{32'h42b660de, 32'h0, 32'h40fcbe13, 32'h400eb174, 32'h425c09f0, 32'h411ef49f, 32'h40b19e9e, 32'h0};
test_input[26664:26671] = '{32'hc1e214a5, 32'h42180e47, 32'h42bcc32e, 32'hc2861f4d, 32'hc23252de, 32'h411da1ff, 32'h415b0c6b, 32'h42759a8b};
test_output[26664:26671] = '{32'h0, 32'h42180e47, 32'h42bcc32e, 32'h0, 32'h0, 32'h411da1ff, 32'h415b0c6b, 32'h42759a8b};
test_input[26672:26679] = '{32'hc26885bf, 32'h4226432b, 32'hc2ac7aea, 32'h4298e0de, 32'hc270668e, 32'hc2243605, 32'hc2c15044, 32'h42a97f2c};
test_output[26672:26679] = '{32'h0, 32'h4226432b, 32'h0, 32'h4298e0de, 32'h0, 32'h0, 32'h0, 32'h42a97f2c};
test_input[26680:26687] = '{32'hc1969203, 32'hc124c3d9, 32'hc28f1a28, 32'hc2b1aba2, 32'h426e2740, 32'hc2a66f36, 32'hc2a0592b, 32'h428ea756};
test_output[26680:26687] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h426e2740, 32'h0, 32'h0, 32'h428ea756};
test_input[26688:26695] = '{32'hc2ae0f65, 32'hc29f659c, 32'hc2aab9b8, 32'h421ca4e7, 32'hc1c71805, 32'h42ade9fc, 32'h42a1ed80, 32'hc2135ce3};
test_output[26688:26695] = '{32'h0, 32'h0, 32'h0, 32'h421ca4e7, 32'h0, 32'h42ade9fc, 32'h42a1ed80, 32'h0};
test_input[26696:26703] = '{32'hc2a15f34, 32'h424f90ba, 32'hc2803088, 32'h41c978ab, 32'hc1b9a920, 32'hc209f768, 32'h4181c29f, 32'h41b9d101};
test_output[26696:26703] = '{32'h0, 32'h424f90ba, 32'h0, 32'h41c978ab, 32'h0, 32'h0, 32'h4181c29f, 32'h41b9d101};
test_input[26704:26711] = '{32'h42a385c3, 32'hc2b61781, 32'hc263a7d3, 32'hc2b467b6, 32'h426b10eb, 32'hc275f3b4, 32'hc1eb64a3, 32'hc22e9ad6};
test_output[26704:26711] = '{32'h42a385c3, 32'h0, 32'h0, 32'h0, 32'h426b10eb, 32'h0, 32'h0, 32'h0};
test_input[26712:26719] = '{32'hc080d766, 32'h42ac33fa, 32'h403073d6, 32'h41e0959b, 32'hc2bcf165, 32'h4280bb9f, 32'h42ba2374, 32'h41fc6951};
test_output[26712:26719] = '{32'h0, 32'h42ac33fa, 32'h403073d6, 32'h41e0959b, 32'h0, 32'h4280bb9f, 32'h42ba2374, 32'h41fc6951};
test_input[26720:26727] = '{32'h419038d2, 32'h423d8e6b, 32'hc0c77801, 32'hc22104a5, 32'hc0fcc288, 32'hc2beef51, 32'h41dbc038, 32'hc1c32e2d};
test_output[26720:26727] = '{32'h419038d2, 32'h423d8e6b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41dbc038, 32'h0};
test_input[26728:26735] = '{32'h42bab9bb, 32'hc1b8cead, 32'h428a629b, 32'hc21087bc, 32'h42c5d779, 32'h426527ad, 32'hc16612b7, 32'hc0424df1};
test_output[26728:26735] = '{32'h42bab9bb, 32'h0, 32'h428a629b, 32'h0, 32'h42c5d779, 32'h426527ad, 32'h0, 32'h0};
test_input[26736:26743] = '{32'h4246756f, 32'h42b780ac, 32'hc23b2130, 32'hc1cd2f9c, 32'hc1f17f7b, 32'h401bc4a9, 32'hc2268976, 32'h42ba0c72};
test_output[26736:26743] = '{32'h4246756f, 32'h42b780ac, 32'h0, 32'h0, 32'h0, 32'h401bc4a9, 32'h0, 32'h42ba0c72};
test_input[26744:26751] = '{32'hc1e2a076, 32'hc28bf39a, 32'hc1ebe31b, 32'hc26df9c8, 32'hc1306b71, 32'h42a9e915, 32'h42879582, 32'h42979fdc};
test_output[26744:26751] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a9e915, 32'h42879582, 32'h42979fdc};
test_input[26752:26759] = '{32'h42375701, 32'h42393d4e, 32'hc20c91f6, 32'hc29c4edc, 32'hc2a31e9d, 32'h4280dd56, 32'h4288e2b0, 32'h42c14249};
test_output[26752:26759] = '{32'h42375701, 32'h42393d4e, 32'h0, 32'h0, 32'h0, 32'h4280dd56, 32'h4288e2b0, 32'h42c14249};
test_input[26760:26767] = '{32'hc23fc088, 32'hc237a510, 32'hc2a3e10c, 32'h429f3a9f, 32'hc2a9cef1, 32'hc213ac2e, 32'hc1f4f057, 32'hc1ff94b6};
test_output[26760:26767] = '{32'h0, 32'h0, 32'h0, 32'h429f3a9f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26768:26775] = '{32'h426dfa93, 32'hc1678402, 32'h42a6ecef, 32'hc236e2e6, 32'hc24917b6, 32'h429e3952, 32'hc27440cf, 32'h412f7f44};
test_output[26768:26775] = '{32'h426dfa93, 32'h0, 32'h42a6ecef, 32'h0, 32'h0, 32'h429e3952, 32'h0, 32'h412f7f44};
test_input[26776:26783] = '{32'hc1e68624, 32'hc277c39f, 32'hc2a48a87, 32'h42b1f0bb, 32'hc1790ec1, 32'h42a9f5db, 32'hc24a092f, 32'hc1e80970};
test_output[26776:26783] = '{32'h0, 32'h0, 32'h0, 32'h42b1f0bb, 32'h0, 32'h42a9f5db, 32'h0, 32'h0};
test_input[26784:26791] = '{32'h420f2a95, 32'hc25c3fa4, 32'h42a96880, 32'hc22797ea, 32'hc21d4a16, 32'hc2a90bf1, 32'hc27dcf02, 32'h418e4b11};
test_output[26784:26791] = '{32'h420f2a95, 32'h0, 32'h42a96880, 32'h0, 32'h0, 32'h0, 32'h0, 32'h418e4b11};
test_input[26792:26799] = '{32'hc24d646d, 32'h428346df, 32'h42976af6, 32'h42abe38b, 32'hc2992331, 32'hc2681955, 32'hc2a40425, 32'h42c6903f};
test_output[26792:26799] = '{32'h0, 32'h428346df, 32'h42976af6, 32'h42abe38b, 32'h0, 32'h0, 32'h0, 32'h42c6903f};
test_input[26800:26807] = '{32'hc09e9720, 32'h421e4d71, 32'h404b6ba1, 32'h409c9fb0, 32'hc19374c6, 32'h410047c4, 32'h424148d0, 32'h429b6288};
test_output[26800:26807] = '{32'h0, 32'h421e4d71, 32'h404b6ba1, 32'h409c9fb0, 32'h0, 32'h410047c4, 32'h424148d0, 32'h429b6288};
test_input[26808:26815] = '{32'hc2885ccf, 32'hc0a282bf, 32'h41b2819f, 32'hc247b366, 32'hc23dc9b1, 32'hc2c25ad8, 32'h42a1d00c, 32'h427bdc40};
test_output[26808:26815] = '{32'h0, 32'h0, 32'h41b2819f, 32'h0, 32'h0, 32'h0, 32'h42a1d00c, 32'h427bdc40};
test_input[26816:26823] = '{32'h420167d0, 32'h421cf352, 32'h42993224, 32'hc0949c24, 32'h41cf02f5, 32'hc1e1ce9d, 32'h4279d961, 32'h42a66aee};
test_output[26816:26823] = '{32'h420167d0, 32'h421cf352, 32'h42993224, 32'h0, 32'h41cf02f5, 32'h0, 32'h4279d961, 32'h42a66aee};
test_input[26824:26831] = '{32'h411785b6, 32'h427b768e, 32'h42911535, 32'h428ef115, 32'hc1dab72b, 32'h425c6b9c, 32'h42c0945d, 32'h4283a783};
test_output[26824:26831] = '{32'h411785b6, 32'h427b768e, 32'h42911535, 32'h428ef115, 32'h0, 32'h425c6b9c, 32'h42c0945d, 32'h4283a783};
test_input[26832:26839] = '{32'hc2871e02, 32'hc1e43369, 32'h429998e1, 32'h4125ed46, 32'h4296dd15, 32'hc1cb4f29, 32'hbf4c221e, 32'hc29ae8b8};
test_output[26832:26839] = '{32'h0, 32'h0, 32'h429998e1, 32'h4125ed46, 32'h4296dd15, 32'h0, 32'h0, 32'h0};
test_input[26840:26847] = '{32'hc16342df, 32'h41d948d8, 32'h42498010, 32'hc2953356, 32'hc24677df, 32'h4139213c, 32'h42acb593, 32'h425c855a};
test_output[26840:26847] = '{32'h0, 32'h41d948d8, 32'h42498010, 32'h0, 32'h0, 32'h4139213c, 32'h42acb593, 32'h425c855a};
test_input[26848:26855] = '{32'hc2029adb, 32'h4280991f, 32'h42a249f4, 32'hc260dcc9, 32'h42ae2893, 32'h4152ce2e, 32'hc05b22dc, 32'h40ca5f1f};
test_output[26848:26855] = '{32'h0, 32'h4280991f, 32'h42a249f4, 32'h0, 32'h42ae2893, 32'h4152ce2e, 32'h0, 32'h40ca5f1f};
test_input[26856:26863] = '{32'hc2ac58ce, 32'h42473f34, 32'hc2af0c84, 32'h41ab6066, 32'hc19bd52f, 32'hc0df2094, 32'h420decea, 32'hc2419107};
test_output[26856:26863] = '{32'h0, 32'h42473f34, 32'h0, 32'h41ab6066, 32'h0, 32'h0, 32'h420decea, 32'h0};
test_input[26864:26871] = '{32'hc10bf8f8, 32'h4191e55e, 32'h4101aafc, 32'h425f0627, 32'hc1fc59cd, 32'h42bade2c, 32'h4218648d, 32'h42c00a1a};
test_output[26864:26871] = '{32'h0, 32'h4191e55e, 32'h4101aafc, 32'h425f0627, 32'h0, 32'h42bade2c, 32'h4218648d, 32'h42c00a1a};
test_input[26872:26879] = '{32'h423a65d6, 32'hc20588ee, 32'h428f1cb8, 32'hc120fa13, 32'hc2b03a0d, 32'hc11b0d27, 32'h429435f5, 32'hc1b2daca};
test_output[26872:26879] = '{32'h423a65d6, 32'h0, 32'h428f1cb8, 32'h0, 32'h0, 32'h0, 32'h429435f5, 32'h0};
test_input[26880:26887] = '{32'h427dd6ac, 32'h428d186d, 32'hc283a624, 32'hc08cdc8b, 32'h423709a9, 32'h42b2ee8f, 32'h418c1d79, 32'hc2c2bb81};
test_output[26880:26887] = '{32'h427dd6ac, 32'h428d186d, 32'h0, 32'h0, 32'h423709a9, 32'h42b2ee8f, 32'h418c1d79, 32'h0};
test_input[26888:26895] = '{32'hc2060cea, 32'hc0faf960, 32'h420ac52a, 32'hc19b92e8, 32'h41e0b8e9, 32'hc29de5c4, 32'h42ba40a1, 32'h42bddde6};
test_output[26888:26895] = '{32'h0, 32'h0, 32'h420ac52a, 32'h0, 32'h41e0b8e9, 32'h0, 32'h42ba40a1, 32'h42bddde6};
test_input[26896:26903] = '{32'hc1642f87, 32'h41ea0c14, 32'hc21fd3ab, 32'hc1162836, 32'h42c1aec8, 32'hc03bae13, 32'hc21936c9, 32'hbeb0ba55};
test_output[26896:26903] = '{32'h0, 32'h41ea0c14, 32'h0, 32'h0, 32'h42c1aec8, 32'h0, 32'h0, 32'h0};
test_input[26904:26911] = '{32'h4292ebd1, 32'hc16b5f12, 32'hc26e780d, 32'h428153ee, 32'hc26211b0, 32'hc2c1a580, 32'hc1f40cd9, 32'hc0c7bb31};
test_output[26904:26911] = '{32'h4292ebd1, 32'h0, 32'h0, 32'h428153ee, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26912:26919] = '{32'hc20e9190, 32'hc2c63ecd, 32'hc21ac090, 32'hc15a4917, 32'hc229920d, 32'hc292a7ce, 32'hc1233162, 32'h4272f124};
test_output[26912:26919] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4272f124};
test_input[26920:26927] = '{32'hc2a96c28, 32'hc1c9623b, 32'hc296daac, 32'h42ae22be, 32'h42909725, 32'h413ad8df, 32'h428c00f9, 32'hc2708f9d};
test_output[26920:26927] = '{32'h0, 32'h0, 32'h0, 32'h42ae22be, 32'h42909725, 32'h413ad8df, 32'h428c00f9, 32'h0};
test_input[26928:26935] = '{32'h42555646, 32'h4223f8f8, 32'hc18f96d5, 32'hc1e0340d, 32'hc29db3f6, 32'hc29495aa, 32'h422c1d42, 32'hc2add5d0};
test_output[26928:26935] = '{32'h42555646, 32'h4223f8f8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422c1d42, 32'h0};
test_input[26936:26943] = '{32'hc2402cc4, 32'hc27559ca, 32'hc2a498a9, 32'h42aa49ff, 32'hc1389c5f, 32'hc20ff92c, 32'h429670e3, 32'hc2303c25};
test_output[26936:26943] = '{32'h0, 32'h0, 32'h0, 32'h42aa49ff, 32'h0, 32'h0, 32'h429670e3, 32'h0};
test_input[26944:26951] = '{32'hc13d4b59, 32'h42a76e4c, 32'h42a8a14e, 32'hc2306254, 32'h42770ec7, 32'h42c175c4, 32'h4235d90f, 32'h4263445a};
test_output[26944:26951] = '{32'h0, 32'h42a76e4c, 32'h42a8a14e, 32'h0, 32'h42770ec7, 32'h42c175c4, 32'h4235d90f, 32'h4263445a};
test_input[26952:26959] = '{32'hc11206ea, 32'hc2b258e5, 32'hc29e9032, 32'hc217abe6, 32'hc212b476, 32'hc2642a33, 32'hc291ab4f, 32'hc10f1651};
test_output[26952:26959] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[26960:26967] = '{32'hc2c02f6b, 32'h42886489, 32'hbe1de41b, 32'hc1966d32, 32'h42be94ed, 32'hc2a801df, 32'hc2640f7d, 32'h42a53bf1};
test_output[26960:26967] = '{32'h0, 32'h42886489, 32'h0, 32'h0, 32'h42be94ed, 32'h0, 32'h0, 32'h42a53bf1};
test_input[26968:26975] = '{32'h428973bc, 32'hc03f28d9, 32'h42988fef, 32'hc1ba48e3, 32'hc28439b5, 32'hc2943798, 32'hc1e4a859, 32'h42726cd8};
test_output[26968:26975] = '{32'h428973bc, 32'h0, 32'h42988fef, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42726cd8};
test_input[26976:26983] = '{32'hc2c389bb, 32'hc25a78f2, 32'h4287f191, 32'hc25fdf2f, 32'hc1e3a991, 32'hc2adf30d, 32'hc25d9c90, 32'h421b72bf};
test_output[26976:26983] = '{32'h0, 32'h0, 32'h4287f191, 32'h0, 32'h0, 32'h0, 32'h0, 32'h421b72bf};
test_input[26984:26991] = '{32'h42bf5b2d, 32'h41d635c1, 32'h422d91fc, 32'hc2608bb9, 32'hc281a07a, 32'h423265d4, 32'hbf80b296, 32'hc2b945ac};
test_output[26984:26991] = '{32'h42bf5b2d, 32'h41d635c1, 32'h422d91fc, 32'h0, 32'h0, 32'h423265d4, 32'h0, 32'h0};
test_input[26992:26999] = '{32'hc0cafd98, 32'h40fdb8bf, 32'h42b838b5, 32'h42b8fb4a, 32'h423c3d01, 32'hc2a279c1, 32'hc1123c58, 32'hc1763552};
test_output[26992:26999] = '{32'h0, 32'h40fdb8bf, 32'h42b838b5, 32'h42b8fb4a, 32'h423c3d01, 32'h0, 32'h0, 32'h0};
test_input[27000:27007] = '{32'h40c34e73, 32'hc2c22fe5, 32'h4208933c, 32'hc19785aa, 32'hc2646ad6, 32'h41938525, 32'hc26f05be, 32'hc165adf3};
test_output[27000:27007] = '{32'h40c34e73, 32'h0, 32'h4208933c, 32'h0, 32'h0, 32'h41938525, 32'h0, 32'h0};
test_input[27008:27015] = '{32'hc1a38f13, 32'h424d6bbe, 32'hc0f17ea7, 32'hc2063fbd, 32'hc18fa4df, 32'hc20a7159, 32'hc019b36d, 32'hc14f0649};
test_output[27008:27015] = '{32'h0, 32'h424d6bbe, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27016:27023] = '{32'h4258744c, 32'h42678a71, 32'h417cf3bd, 32'h426de340, 32'hc20780d0, 32'h4290258e, 32'h4181a8ec, 32'hc2abc463};
test_output[27016:27023] = '{32'h4258744c, 32'h42678a71, 32'h417cf3bd, 32'h426de340, 32'h0, 32'h4290258e, 32'h4181a8ec, 32'h0};
test_input[27024:27031] = '{32'h41a38b17, 32'hc2268d3d, 32'h42c1d55a, 32'hc2a33a47, 32'h42855f92, 32'h41ad7425, 32'h4215e72c, 32'hc2717c8d};
test_output[27024:27031] = '{32'h41a38b17, 32'h0, 32'h42c1d55a, 32'h0, 32'h42855f92, 32'h41ad7425, 32'h4215e72c, 32'h0};
test_input[27032:27039] = '{32'h418473bd, 32'h419cf229, 32'hc261a64d, 32'h42b84738, 32'h41c15729, 32'h42b3feef, 32'hc283f82b, 32'hc2830c3c};
test_output[27032:27039] = '{32'h418473bd, 32'h419cf229, 32'h0, 32'h42b84738, 32'h41c15729, 32'h42b3feef, 32'h0, 32'h0};
test_input[27040:27047] = '{32'h41857fd1, 32'hc20c54fa, 32'h42b37e84, 32'hc23a9955, 32'hc267933d, 32'h4119dc80, 32'h41847282, 32'hc1ca7d64};
test_output[27040:27047] = '{32'h41857fd1, 32'h0, 32'h42b37e84, 32'h0, 32'h0, 32'h4119dc80, 32'h41847282, 32'h0};
test_input[27048:27055] = '{32'hc2c450b1, 32'h40484f35, 32'h426ecdf1, 32'hc1790dc3, 32'hc2c6c485, 32'hbf56f13f, 32'hc269b7a8, 32'hc2245146};
test_output[27048:27055] = '{32'h0, 32'h40484f35, 32'h426ecdf1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27056:27063] = '{32'hc267fd1f, 32'h425345cc, 32'h41bc6222, 32'h41cdc13f, 32'h41fab27f, 32'hc20ba14b, 32'h423573a4, 32'hc258c8e6};
test_output[27056:27063] = '{32'h0, 32'h425345cc, 32'h41bc6222, 32'h41cdc13f, 32'h41fab27f, 32'h0, 32'h423573a4, 32'h0};
test_input[27064:27071] = '{32'h416817ee, 32'h42a3c37a, 32'hc25e0ef5, 32'hc21ea2b0, 32'h42b030b3, 32'hc2c2fbb8, 32'hc2844dbd, 32'h42749b01};
test_output[27064:27071] = '{32'h416817ee, 32'h42a3c37a, 32'h0, 32'h0, 32'h42b030b3, 32'h0, 32'h0, 32'h42749b01};
test_input[27072:27079] = '{32'h42a9ff77, 32'hc115d24e, 32'hc1d323b7, 32'h42b6b9b6, 32'hc230039a, 32'h423c6996, 32'hc1f39a3c, 32'hc23e2c07};
test_output[27072:27079] = '{32'h42a9ff77, 32'h0, 32'h0, 32'h42b6b9b6, 32'h0, 32'h423c6996, 32'h0, 32'h0};
test_input[27080:27087] = '{32'hc21cd01a, 32'h4192928a, 32'h42719e3f, 32'hc28a96b0, 32'hc2710e30, 32'h429dc928, 32'hc2acc749, 32'h42c5bd97};
test_output[27080:27087] = '{32'h0, 32'h4192928a, 32'h42719e3f, 32'h0, 32'h0, 32'h429dc928, 32'h0, 32'h42c5bd97};
test_input[27088:27095] = '{32'h3d99b6ce, 32'hc0f3a00c, 32'h42bfb3bb, 32'h428fd083, 32'hc1201799, 32'h428bf114, 32'hc1c46f77, 32'hc2179043};
test_output[27088:27095] = '{32'h3d99b6ce, 32'h0, 32'h42bfb3bb, 32'h428fd083, 32'h0, 32'h428bf114, 32'h0, 32'h0};
test_input[27096:27103] = '{32'h4280ad55, 32'hc2a46b6e, 32'h4133dd22, 32'h41bd2307, 32'h42a32a56, 32'h419ace74, 32'hc2a78197, 32'h4284d8ab};
test_output[27096:27103] = '{32'h4280ad55, 32'h0, 32'h4133dd22, 32'h41bd2307, 32'h42a32a56, 32'h419ace74, 32'h0, 32'h4284d8ab};
test_input[27104:27111] = '{32'h41e272d5, 32'h420fbe2d, 32'h427242f6, 32'hc262dd24, 32'h42a1694a, 32'h42b72315, 32'h414a9b74, 32'h42957ced};
test_output[27104:27111] = '{32'h41e272d5, 32'h420fbe2d, 32'h427242f6, 32'h0, 32'h42a1694a, 32'h42b72315, 32'h414a9b74, 32'h42957ced};
test_input[27112:27119] = '{32'hc2bdab93, 32'h426badcc, 32'hc2a7db19, 32'hc264d40b, 32'hc28d7197, 32'hc258610c, 32'hc2a5ba79, 32'h40b0f828};
test_output[27112:27119] = '{32'h0, 32'h426badcc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40b0f828};
test_input[27120:27127] = '{32'h42919843, 32'hc0afd04d, 32'hc23aa277, 32'h42b24ab1, 32'h429d33bd, 32'hc2ab8ee3, 32'h4279207f, 32'h429e186d};
test_output[27120:27127] = '{32'h42919843, 32'h0, 32'h0, 32'h42b24ab1, 32'h429d33bd, 32'h0, 32'h4279207f, 32'h429e186d};
test_input[27128:27135] = '{32'hc247c273, 32'h41e08339, 32'h4255330f, 32'hc2be538c, 32'hc2829757, 32'hc1b56619, 32'hc20c7c4d, 32'h426ef454};
test_output[27128:27135] = '{32'h0, 32'h41e08339, 32'h4255330f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426ef454};
test_input[27136:27143] = '{32'hc10ed6d0, 32'hc1199d26, 32'h417a7ac4, 32'hc2194b71, 32'h3fa6ecf3, 32'h42863223, 32'h42b7fb36, 32'hc19f3261};
test_output[27136:27143] = '{32'h0, 32'h0, 32'h417a7ac4, 32'h0, 32'h3fa6ecf3, 32'h42863223, 32'h42b7fb36, 32'h0};
test_input[27144:27151] = '{32'hc159561b, 32'hc1858488, 32'hc1a12aaf, 32'h427e6f7f, 32'h41b5cd3f, 32'h4249b87b, 32'hc28a6b79, 32'h42bc111d};
test_output[27144:27151] = '{32'h0, 32'h0, 32'h0, 32'h427e6f7f, 32'h41b5cd3f, 32'h4249b87b, 32'h0, 32'h42bc111d};
test_input[27152:27159] = '{32'hc1f65a8f, 32'h429f69a9, 32'h4210e79a, 32'h423c3f48, 32'hc26d5735, 32'hc1d7f085, 32'h42a32859, 32'h428995db};
test_output[27152:27159] = '{32'h0, 32'h429f69a9, 32'h4210e79a, 32'h423c3f48, 32'h0, 32'h0, 32'h42a32859, 32'h428995db};
test_input[27160:27167] = '{32'hc297be2a, 32'hc22eda6d, 32'hc292003a, 32'h42063bfe, 32'hc277d2d0, 32'h4138ba22, 32'hc10bb5d5, 32'hc15e8185};
test_output[27160:27167] = '{32'h0, 32'h0, 32'h0, 32'h42063bfe, 32'h0, 32'h4138ba22, 32'h0, 32'h0};
test_input[27168:27175] = '{32'h405edff3, 32'hc239e9f0, 32'h41c3a45c, 32'h41d7f447, 32'hc2039f81, 32'h4299252c, 32'h426c135a, 32'h4282cefd};
test_output[27168:27175] = '{32'h405edff3, 32'h0, 32'h41c3a45c, 32'h41d7f447, 32'h0, 32'h4299252c, 32'h426c135a, 32'h4282cefd};
test_input[27176:27183] = '{32'h4273a446, 32'hc1eede80, 32'hc17b4223, 32'h429ccb58, 32'hc294d0f2, 32'hc2673e60, 32'hc18ebd7e, 32'h418eee49};
test_output[27176:27183] = '{32'h4273a446, 32'h0, 32'h0, 32'h429ccb58, 32'h0, 32'h0, 32'h0, 32'h418eee49};
test_input[27184:27191] = '{32'hc24ea274, 32'hc21e717a, 32'h42be2fc2, 32'hc290c648, 32'hc21fa239, 32'h4270648a, 32'h42a84619, 32'hc22d5116};
test_output[27184:27191] = '{32'h0, 32'h0, 32'h42be2fc2, 32'h0, 32'h0, 32'h4270648a, 32'h42a84619, 32'h0};
test_input[27192:27199] = '{32'hc2c055c6, 32'hc28c55e0, 32'hc1eb2f1f, 32'hc29dcd7a, 32'h41fa4e99, 32'h42b8ab14, 32'hc24777da, 32'h425335e2};
test_output[27192:27199] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41fa4e99, 32'h42b8ab14, 32'h0, 32'h425335e2};
test_input[27200:27207] = '{32'hc2983c9e, 32'hc1b6bd66, 32'h4281609d, 32'h4264a5f8, 32'hc252f444, 32'hc294fcd3, 32'hc23319f4, 32'h42208fed};
test_output[27200:27207] = '{32'h0, 32'h0, 32'h4281609d, 32'h4264a5f8, 32'h0, 32'h0, 32'h0, 32'h42208fed};
test_input[27208:27215] = '{32'h425daf93, 32'h41e0eec5, 32'hc206a8ca, 32'hc2044ef3, 32'h42180880, 32'hc296a329, 32'hc1cb67ce, 32'h424fbf9e};
test_output[27208:27215] = '{32'h425daf93, 32'h41e0eec5, 32'h0, 32'h0, 32'h42180880, 32'h0, 32'h0, 32'h424fbf9e};
test_input[27216:27223] = '{32'hc228fc8c, 32'h42260665, 32'hc135b6d7, 32'hc2c33456, 32'h41e4a459, 32'h42a202aa, 32'hc1ecbc69, 32'hc2ac6309};
test_output[27216:27223] = '{32'h0, 32'h42260665, 32'h0, 32'h0, 32'h41e4a459, 32'h42a202aa, 32'h0, 32'h0};
test_input[27224:27231] = '{32'hc29b91d0, 32'h429421f6, 32'h421da83f, 32'hc1b1e864, 32'hc24e4a44, 32'hc2102d98, 32'hc2beefff, 32'hc1fbf437};
test_output[27224:27231] = '{32'h0, 32'h429421f6, 32'h421da83f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27232:27239] = '{32'h4293493b, 32'hc26de8e2, 32'h41cd7bec, 32'h421c36ef, 32'h42817bba, 32'hc189b06c, 32'h42988a53, 32'hc217d8e0};
test_output[27232:27239] = '{32'h4293493b, 32'h0, 32'h41cd7bec, 32'h421c36ef, 32'h42817bba, 32'h0, 32'h42988a53, 32'h0};
test_input[27240:27247] = '{32'h412a626f, 32'h41fd3d0b, 32'h418fa0d6, 32'hc20add5b, 32'h423f114b, 32'hc27778ef, 32'hc2958e08, 32'hc27eae15};
test_output[27240:27247] = '{32'h412a626f, 32'h41fd3d0b, 32'h418fa0d6, 32'h0, 32'h423f114b, 32'h0, 32'h0, 32'h0};
test_input[27248:27255] = '{32'h41ac20c9, 32'h42aeca51, 32'hc21aeab3, 32'hc210a675, 32'h42b08ae7, 32'h42995c67, 32'hc2830b26, 32'hc294da02};
test_output[27248:27255] = '{32'h41ac20c9, 32'h42aeca51, 32'h0, 32'h0, 32'h42b08ae7, 32'h42995c67, 32'h0, 32'h0};
test_input[27256:27263] = '{32'hc226887c, 32'hc2971c72, 32'hc2501f6d, 32'hc1959ecc, 32'h42616bdf, 32'hc162e2e2, 32'h40d749c4, 32'hc2a45c57};
test_output[27256:27263] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42616bdf, 32'h0, 32'h40d749c4, 32'h0};
test_input[27264:27271] = '{32'h4284d1b2, 32'h42c48bb8, 32'h411325d7, 32'hc09c2256, 32'h42a32dc0, 32'hc24c6780, 32'h42a77142, 32'h4283b052};
test_output[27264:27271] = '{32'h4284d1b2, 32'h42c48bb8, 32'h411325d7, 32'h0, 32'h42a32dc0, 32'h0, 32'h42a77142, 32'h4283b052};
test_input[27272:27279] = '{32'h4185bde0, 32'hc1f5ea98, 32'h42a98f8b, 32'hc26599e2, 32'h415bb8b5, 32'h413821b8, 32'h419f9abb, 32'h427556d1};
test_output[27272:27279] = '{32'h4185bde0, 32'h0, 32'h42a98f8b, 32'h0, 32'h415bb8b5, 32'h413821b8, 32'h419f9abb, 32'h427556d1};
test_input[27280:27287] = '{32'hc229cb81, 32'hc209fb10, 32'hc24e3f47, 32'hc2a9e2ef, 32'hc26ce77c, 32'h4258b743, 32'hc29355b7, 32'h413d0344};
test_output[27280:27287] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4258b743, 32'h0, 32'h413d0344};
test_input[27288:27295] = '{32'hc1d7ef80, 32'h4281afec, 32'h413df458, 32'hc2c0d788, 32'hc2842ac5, 32'h429a94ca, 32'h42aa4091, 32'hc026e39d};
test_output[27288:27295] = '{32'h0, 32'h4281afec, 32'h413df458, 32'h0, 32'h0, 32'h429a94ca, 32'h42aa4091, 32'h0};
test_input[27296:27303] = '{32'hc269735c, 32'hc19fd3e2, 32'h429af130, 32'h42779921, 32'hc1d19c8b, 32'h41e611e0, 32'hc2721db4, 32'h3e47fe45};
test_output[27296:27303] = '{32'h0, 32'h0, 32'h429af130, 32'h42779921, 32'h0, 32'h41e611e0, 32'h0, 32'h3e47fe45};
test_input[27304:27311] = '{32'h42b6b125, 32'hc2a6b349, 32'h419583d0, 32'hc2b9c244, 32'h4282a772, 32'hc29c43c7, 32'h417ef1a3, 32'h428becad};
test_output[27304:27311] = '{32'h42b6b125, 32'h0, 32'h419583d0, 32'h0, 32'h4282a772, 32'h0, 32'h417ef1a3, 32'h428becad};
test_input[27312:27319] = '{32'h42868c2c, 32'hc298681f, 32'hc1b2aea5, 32'hc29e6bfd, 32'h428c152c, 32'h426f9190, 32'h41f1205b, 32'hc179b607};
test_output[27312:27319] = '{32'h42868c2c, 32'h0, 32'h0, 32'h0, 32'h428c152c, 32'h426f9190, 32'h41f1205b, 32'h0};
test_input[27320:27327] = '{32'hc21076af, 32'h427a023b, 32'hc28d6b3f, 32'h428d6280, 32'h41e3b5b9, 32'hc259f54c, 32'hc1a9e304, 32'h42351cab};
test_output[27320:27327] = '{32'h0, 32'h427a023b, 32'h0, 32'h428d6280, 32'h41e3b5b9, 32'h0, 32'h0, 32'h42351cab};
test_input[27328:27335] = '{32'h4077ba2b, 32'h42bab154, 32'h42910b04, 32'h42903885, 32'hc25aaa72, 32'h424e9a11, 32'h42778957, 32'h428e399a};
test_output[27328:27335] = '{32'h4077ba2b, 32'h42bab154, 32'h42910b04, 32'h42903885, 32'h0, 32'h424e9a11, 32'h42778957, 32'h428e399a};
test_input[27336:27343] = '{32'hc20d41ee, 32'h42b1a5ab, 32'h41715e65, 32'hc2bb4d1a, 32'hc28e72b3, 32'h42bc7988, 32'hc10bb1b6, 32'h42aaf0c7};
test_output[27336:27343] = '{32'h0, 32'h42b1a5ab, 32'h41715e65, 32'h0, 32'h0, 32'h42bc7988, 32'h0, 32'h42aaf0c7};
test_input[27344:27351] = '{32'h42b1c782, 32'hc2348f1b, 32'h429192b0, 32'h41170188, 32'hc024809e, 32'h429a7bed, 32'hc2a15a6f, 32'hc24df580};
test_output[27344:27351] = '{32'h42b1c782, 32'h0, 32'h429192b0, 32'h41170188, 32'h0, 32'h429a7bed, 32'h0, 32'h0};
test_input[27352:27359] = '{32'h425deb2a, 32'hc1d97c62, 32'h41828c7b, 32'hc0df9e69, 32'hc295c9d6, 32'hc24131dd, 32'h428f505b, 32'hc151d369};
test_output[27352:27359] = '{32'h425deb2a, 32'h0, 32'h41828c7b, 32'h0, 32'h0, 32'h0, 32'h428f505b, 32'h0};
test_input[27360:27367] = '{32'hc1cf5b48, 32'h4010cc0b, 32'h41f0b506, 32'h42ab7cd8, 32'hc078ece0, 32'hc1fa8bc6, 32'hc2355064, 32'h4146450d};
test_output[27360:27367] = '{32'h0, 32'h4010cc0b, 32'h41f0b506, 32'h42ab7cd8, 32'h0, 32'h0, 32'h0, 32'h4146450d};
test_input[27368:27375] = '{32'hc11ae7a0, 32'h404060f0, 32'hbfc7fdb3, 32'hc272a147, 32'h42b15e1d, 32'hc262b4b2, 32'hc2b46fe2, 32'h42bb087f};
test_output[27368:27375] = '{32'h0, 32'h404060f0, 32'h0, 32'h0, 32'h42b15e1d, 32'h0, 32'h0, 32'h42bb087f};
test_input[27376:27383] = '{32'h428008b7, 32'h41cab07a, 32'hc29f6f06, 32'hc29cb450, 32'h425d34ad, 32'hc13ff1b6, 32'h42a1d1ea, 32'hc2be3a39};
test_output[27376:27383] = '{32'h428008b7, 32'h41cab07a, 32'h0, 32'h0, 32'h425d34ad, 32'h0, 32'h42a1d1ea, 32'h0};
test_input[27384:27391] = '{32'hc26332a1, 32'h42c4f765, 32'h4214c732, 32'h423421ac, 32'hc27745ed, 32'hc2aaa277, 32'hc2c3ff38, 32'h428fd8d1};
test_output[27384:27391] = '{32'h0, 32'h42c4f765, 32'h4214c732, 32'h423421ac, 32'h0, 32'h0, 32'h0, 32'h428fd8d1};
test_input[27392:27399] = '{32'h42b69f93, 32'hc2914267, 32'h42a33d98, 32'hc1de2252, 32'h42a0ea4c, 32'hbfafca27, 32'hc0446b68, 32'hc114630e};
test_output[27392:27399] = '{32'h42b69f93, 32'h0, 32'h42a33d98, 32'h0, 32'h42a0ea4c, 32'h0, 32'h0, 32'h0};
test_input[27400:27407] = '{32'hc281a977, 32'hbf91c83c, 32'hc280c315, 32'hc229ce0a, 32'h423ef63d, 32'hc238b3dd, 32'h4255276e, 32'hc23366e9};
test_output[27400:27407] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h423ef63d, 32'h0, 32'h4255276e, 32'h0};
test_input[27408:27415] = '{32'hc1738968, 32'h42b5231c, 32'h41b63a57, 32'h428caa0b, 32'hbf868b35, 32'hc2226e22, 32'hc2a8617a, 32'hc13e600e};
test_output[27408:27415] = '{32'h0, 32'h42b5231c, 32'h41b63a57, 32'h428caa0b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27416:27423] = '{32'hc1181549, 32'hc22a865c, 32'h42bcd720, 32'h416afc85, 32'h4195353c, 32'hc2b90034, 32'h42476ee6, 32'h4210bbbd};
test_output[27416:27423] = '{32'h0, 32'h0, 32'h42bcd720, 32'h416afc85, 32'h4195353c, 32'h0, 32'h42476ee6, 32'h4210bbbd};
test_input[27424:27431] = '{32'hc2c43634, 32'h42876ad6, 32'h41cf8ad3, 32'h4288495c, 32'hc1a5461c, 32'h41d6b5e5, 32'h42292a99, 32'h428f92b1};
test_output[27424:27431] = '{32'h0, 32'h42876ad6, 32'h41cf8ad3, 32'h4288495c, 32'h0, 32'h41d6b5e5, 32'h42292a99, 32'h428f92b1};
test_input[27432:27439] = '{32'h41dd8914, 32'h429aa0d5, 32'hc1c4b55b, 32'hc23b9830, 32'h420ebcfa, 32'h41f8ea5d, 32'hc22cd506, 32'hc19a46d7};
test_output[27432:27439] = '{32'h41dd8914, 32'h429aa0d5, 32'h0, 32'h0, 32'h420ebcfa, 32'h41f8ea5d, 32'h0, 32'h0};
test_input[27440:27447] = '{32'hc1d44177, 32'hc25db50b, 32'h42b2b613, 32'h42a9875e, 32'h410bfc49, 32'hc2787dd4, 32'h42b58ad7, 32'hc294aba4};
test_output[27440:27447] = '{32'h0, 32'h0, 32'h42b2b613, 32'h42a9875e, 32'h410bfc49, 32'h0, 32'h42b58ad7, 32'h0};
test_input[27448:27455] = '{32'h420890cb, 32'h42becc5a, 32'hc1b73819, 32'hc28c4512, 32'h40fb7029, 32'h428a7901, 32'h42940834, 32'hc26749bb};
test_output[27448:27455] = '{32'h420890cb, 32'h42becc5a, 32'h0, 32'h0, 32'h40fb7029, 32'h428a7901, 32'h42940834, 32'h0};
test_input[27456:27463] = '{32'h407f13a0, 32'hc2252a93, 32'h3e4fd2f5, 32'hc2b9fc99, 32'h412c22b4, 32'hc2055423, 32'hc252863f, 32'hc293613e};
test_output[27456:27463] = '{32'h407f13a0, 32'h0, 32'h3e4fd2f5, 32'h0, 32'h412c22b4, 32'h0, 32'h0, 32'h0};
test_input[27464:27471] = '{32'hc29b0b89, 32'hc2126f93, 32'h42927b94, 32'h42bcb73e, 32'h4245d148, 32'hc2b76aa2, 32'hc0543676, 32'hc114a73f};
test_output[27464:27471] = '{32'h0, 32'h0, 32'h42927b94, 32'h42bcb73e, 32'h4245d148, 32'h0, 32'h0, 32'h0};
test_input[27472:27479] = '{32'h427bbb03, 32'hc2b9b6ff, 32'h42832098, 32'hc0e30385, 32'hc24945b3, 32'h41fbf5ad, 32'hc29945d6, 32'hc230a147};
test_output[27472:27479] = '{32'h427bbb03, 32'h0, 32'h42832098, 32'h0, 32'h0, 32'h41fbf5ad, 32'h0, 32'h0};
test_input[27480:27487] = '{32'hc27a5753, 32'h42aa2088, 32'hc1d5190b, 32'hc250058c, 32'h42b8cb1f, 32'h4298c4c5, 32'hc22e6b44, 32'hc2131d3a};
test_output[27480:27487] = '{32'h0, 32'h42aa2088, 32'h0, 32'h0, 32'h42b8cb1f, 32'h4298c4c5, 32'h0, 32'h0};
test_input[27488:27495] = '{32'hc226db27, 32'h420eea8b, 32'hc1f98201, 32'h42bf8ef6, 32'h426abec7, 32'h428cc27e, 32'hc299c40a, 32'hc2970e71};
test_output[27488:27495] = '{32'h0, 32'h420eea8b, 32'h0, 32'h42bf8ef6, 32'h426abec7, 32'h428cc27e, 32'h0, 32'h0};
test_input[27496:27503] = '{32'h428c334e, 32'h42424466, 32'hc1e88afe, 32'h426f0624, 32'hc217b1ab, 32'hc286def2, 32'hbeb70aef, 32'h419fb53c};
test_output[27496:27503] = '{32'h428c334e, 32'h42424466, 32'h0, 32'h426f0624, 32'h0, 32'h0, 32'h0, 32'h419fb53c};
test_input[27504:27511] = '{32'h417bf4e4, 32'h412e6aea, 32'hc2524dd4, 32'hc29375bf, 32'h42b3b0aa, 32'h422ab1d0, 32'h4200677d, 32'h42c4b64d};
test_output[27504:27511] = '{32'h417bf4e4, 32'h412e6aea, 32'h0, 32'h0, 32'h42b3b0aa, 32'h422ab1d0, 32'h4200677d, 32'h42c4b64d};
test_input[27512:27519] = '{32'h4221b99e, 32'hc2a66446, 32'h42bed993, 32'hc2893cdf, 32'h42bd4e6c, 32'h428ddcad, 32'h40700c8d, 32'hc23003f2};
test_output[27512:27519] = '{32'h4221b99e, 32'h0, 32'h42bed993, 32'h0, 32'h42bd4e6c, 32'h428ddcad, 32'h40700c8d, 32'h0};
test_input[27520:27527] = '{32'hc1febbd8, 32'hc1aebdaf, 32'hc2a18667, 32'hbfb8a5da, 32'hc267c75a, 32'h40d9b3eb, 32'h42467a5c, 32'hc1a3e18b};
test_output[27520:27527] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40d9b3eb, 32'h42467a5c, 32'h0};
test_input[27528:27535] = '{32'h42c5766d, 32'hc26181fb, 32'h42b1eb20, 32'hc20cc715, 32'h421321a3, 32'h42835795, 32'hc226c82e, 32'h41897adb};
test_output[27528:27535] = '{32'h42c5766d, 32'h0, 32'h42b1eb20, 32'h0, 32'h421321a3, 32'h42835795, 32'h0, 32'h41897adb};
test_input[27536:27543] = '{32'hc2146afc, 32'hc27f7e08, 32'h427a6692, 32'hc10399f9, 32'h41f80e75, 32'h40deccc7, 32'hc236a40f, 32'hc217e3cb};
test_output[27536:27543] = '{32'h0, 32'h0, 32'h427a6692, 32'h0, 32'h41f80e75, 32'h40deccc7, 32'h0, 32'h0};
test_input[27544:27551] = '{32'h4266ee79, 32'h4258ba66, 32'hc175864c, 32'hc1f2755a, 32'h42b09f46, 32'hc180d5a4, 32'hc242b427, 32'h42209bb7};
test_output[27544:27551] = '{32'h4266ee79, 32'h4258ba66, 32'h0, 32'h0, 32'h42b09f46, 32'h0, 32'h0, 32'h42209bb7};
test_input[27552:27559] = '{32'hc263545f, 32'h4278b89b, 32'h4202b151, 32'h41bbdd42, 32'hc29bb766, 32'hc249dddd, 32'h42801c3e, 32'hc246e4b2};
test_output[27552:27559] = '{32'h0, 32'h4278b89b, 32'h4202b151, 32'h41bbdd42, 32'h0, 32'h0, 32'h42801c3e, 32'h0};
test_input[27560:27567] = '{32'hc2040670, 32'hc2050cfe, 32'hc28ad308, 32'hc26a03e3, 32'h41212b63, 32'h40f72285, 32'hc2442552, 32'hc2ae86e7};
test_output[27560:27567] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41212b63, 32'h40f72285, 32'h0, 32'h0};
test_input[27568:27575] = '{32'h418ac700, 32'h4228c771, 32'hc27d552e, 32'h4218dc8d, 32'hc22948a0, 32'h42470712, 32'hc283757b, 32'hc1b0c3eb};
test_output[27568:27575] = '{32'h418ac700, 32'h4228c771, 32'h0, 32'h4218dc8d, 32'h0, 32'h42470712, 32'h0, 32'h0};
test_input[27576:27583] = '{32'hc2354a4c, 32'h42563c81, 32'hc20cf5a6, 32'hc27921c1, 32'h42a04e74, 32'h40b7c1c0, 32'h4180dafc, 32'h4246b697};
test_output[27576:27583] = '{32'h0, 32'h42563c81, 32'h0, 32'h0, 32'h42a04e74, 32'h40b7c1c0, 32'h4180dafc, 32'h4246b697};
test_input[27584:27591] = '{32'hc1af8293, 32'hbff928d9, 32'hc221a15d, 32'h4280836e, 32'hc2c6c44a, 32'hc1ec8e63, 32'h42b1bfe4, 32'hc2c5e84c};
test_output[27584:27591] = '{32'h0, 32'h0, 32'h0, 32'h4280836e, 32'h0, 32'h0, 32'h42b1bfe4, 32'h0};
test_input[27592:27599] = '{32'hc2b4048d, 32'hc2c2d9d4, 32'hc1b95e6d, 32'h424822fe, 32'hc2a395b7, 32'hc1970802, 32'h428b7ba7, 32'hc2a5894b};
test_output[27592:27599] = '{32'h0, 32'h0, 32'h0, 32'h424822fe, 32'h0, 32'h0, 32'h428b7ba7, 32'h0};
test_input[27600:27607] = '{32'h427f8407, 32'hc2b27cfb, 32'h41112464, 32'hc1c98160, 32'h42784fe7, 32'h41a80591, 32'h419e2b9e, 32'h42be0b9d};
test_output[27600:27607] = '{32'h427f8407, 32'h0, 32'h41112464, 32'h0, 32'h42784fe7, 32'h41a80591, 32'h419e2b9e, 32'h42be0b9d};
test_input[27608:27615] = '{32'hc02edf06, 32'h422d36b0, 32'hc289c345, 32'hc1249bc5, 32'hc167ac99, 32'hc2607b70, 32'hc1ac01bf, 32'hc0d4575b};
test_output[27608:27615] = '{32'h0, 32'h422d36b0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27616:27623] = '{32'hc2c284a5, 32'h41d9be63, 32'hc28004dd, 32'h41ba0b22, 32'hc2a94fab, 32'hc2035890, 32'h41fe361f, 32'hc12ad2bc};
test_output[27616:27623] = '{32'h0, 32'h41d9be63, 32'h0, 32'h41ba0b22, 32'h0, 32'h0, 32'h41fe361f, 32'h0};
test_input[27624:27631] = '{32'h42b61958, 32'hc2868707, 32'h42ba0b05, 32'h4147cec9, 32'hc16088a8, 32'hc0ab2b06, 32'hc2837583, 32'hc2ba1b9c};
test_output[27624:27631] = '{32'h42b61958, 32'h0, 32'h42ba0b05, 32'h4147cec9, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27632:27639] = '{32'h4256f767, 32'hc228753f, 32'h4219714a, 32'h42c252b7, 32'hc29daf0a, 32'h42580994, 32'hc28c8926, 32'h42a4df91};
test_output[27632:27639] = '{32'h4256f767, 32'h0, 32'h4219714a, 32'h42c252b7, 32'h0, 32'h42580994, 32'h0, 32'h42a4df91};
test_input[27640:27647] = '{32'hc2c15fbb, 32'hc1a77d48, 32'hc1288b50, 32'h42c58c64, 32'h41e493ca, 32'h4226df72, 32'hc268c8e9, 32'h4180cb93};
test_output[27640:27647] = '{32'h0, 32'h0, 32'h0, 32'h42c58c64, 32'h41e493ca, 32'h4226df72, 32'h0, 32'h4180cb93};
test_input[27648:27655] = '{32'hc2ad6c7c, 32'hc24cada7, 32'hc255d903, 32'hc284d9bf, 32'hc0e00c00, 32'hc2203427, 32'h42653c44, 32'hc256fb6a};
test_output[27648:27655] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42653c44, 32'h0};
test_input[27656:27663] = '{32'h42163cb1, 32'hc2acda57, 32'hc18110b5, 32'h428c74b8, 32'hc2c1b7c4, 32'hc2891425, 32'hc2b2cc81, 32'hc2311b17};
test_output[27656:27663] = '{32'h42163cb1, 32'h0, 32'h0, 32'h428c74b8, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27664:27671] = '{32'h41ac1f05, 32'hc072f519, 32'h424bb868, 32'hc14b7a89, 32'hc19d0d5e, 32'hc0d687cf, 32'hc1484f4b, 32'hc2a305a2};
test_output[27664:27671] = '{32'h41ac1f05, 32'h0, 32'h424bb868, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27672:27679] = '{32'h421e1d76, 32'hc28bc563, 32'h401e25d6, 32'h41145ecf, 32'hc280460b, 32'h424b8392, 32'h42526228, 32'h41c57089};
test_output[27672:27679] = '{32'h421e1d76, 32'h0, 32'h401e25d6, 32'h41145ecf, 32'h0, 32'h424b8392, 32'h42526228, 32'h41c57089};
test_input[27680:27687] = '{32'h42832402, 32'h41d2fe62, 32'hc27ebf57, 32'h4272cb86, 32'h42905a65, 32'hc140b542, 32'h42afe269, 32'hc2297faa};
test_output[27680:27687] = '{32'h42832402, 32'h41d2fe62, 32'h0, 32'h4272cb86, 32'h42905a65, 32'h0, 32'h42afe269, 32'h0};
test_input[27688:27695] = '{32'h4263b6a3, 32'h412bc0fe, 32'h42bb9bee, 32'h41e69f5b, 32'h42a09fca, 32'hc27fc9ac, 32'h42ab9486, 32'h42c381e2};
test_output[27688:27695] = '{32'h4263b6a3, 32'h412bc0fe, 32'h42bb9bee, 32'h41e69f5b, 32'h42a09fca, 32'h0, 32'h42ab9486, 32'h42c381e2};
test_input[27696:27703] = '{32'h41858592, 32'h424425ff, 32'hc2005dba, 32'hc24ac3b0, 32'h429ce5ec, 32'h42b3937b, 32'hc1f715ce, 32'h423c1ede};
test_output[27696:27703] = '{32'h41858592, 32'h424425ff, 32'h0, 32'h0, 32'h429ce5ec, 32'h42b3937b, 32'h0, 32'h423c1ede};
test_input[27704:27711] = '{32'hc1bc34ee, 32'h426f3dca, 32'hc272cda3, 32'hc2698d18, 32'h42344b46, 32'hc2aaef06, 32'hc1869ed7, 32'h41ed08d3};
test_output[27704:27711] = '{32'h0, 32'h426f3dca, 32'h0, 32'h0, 32'h42344b46, 32'h0, 32'h0, 32'h41ed08d3};
test_input[27712:27719] = '{32'h42317688, 32'hc1091d95, 32'hc20b4a97, 32'h4237fd99, 32'h424a5ad0, 32'hc2128f98, 32'hc2859d16, 32'h4084352c};
test_output[27712:27719] = '{32'h42317688, 32'h0, 32'h0, 32'h4237fd99, 32'h424a5ad0, 32'h0, 32'h0, 32'h4084352c};
test_input[27720:27727] = '{32'hc2465432, 32'h41ac8aab, 32'hc1b3a0b9, 32'hc10e414b, 32'hc29324f6, 32'hc2310260, 32'hc1b69298, 32'hc1bc661d};
test_output[27720:27727] = '{32'h0, 32'h41ac8aab, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27728:27735] = '{32'h3e5dcd83, 32'h42bbf4ad, 32'hc189875b, 32'h42a83596, 32'h41c76715, 32'hc2a5c477, 32'hc2653414, 32'h42113b74};
test_output[27728:27735] = '{32'h3e5dcd83, 32'h42bbf4ad, 32'h0, 32'h42a83596, 32'h41c76715, 32'h0, 32'h0, 32'h42113b74};
test_input[27736:27743] = '{32'h425085b5, 32'hc29e4576, 32'hc23d0f7a, 32'h42915c5c, 32'h41a51bc3, 32'hc1c04321, 32'hc28ec823, 32'hc2341af1};
test_output[27736:27743] = '{32'h425085b5, 32'h0, 32'h0, 32'h42915c5c, 32'h41a51bc3, 32'h0, 32'h0, 32'h0};
test_input[27744:27751] = '{32'hc234b5bc, 32'hc2a0f5bb, 32'hc2171f73, 32'h41a09ece, 32'h42544b22, 32'hc2a499b0, 32'h4278b9d9, 32'hc2b53a7c};
test_output[27744:27751] = '{32'h0, 32'h0, 32'h0, 32'h41a09ece, 32'h42544b22, 32'h0, 32'h4278b9d9, 32'h0};
test_input[27752:27759] = '{32'hc2c64c1e, 32'hc04179bc, 32'hc2b0d5c8, 32'hc2a95588, 32'hc185fba8, 32'hc1bd3504, 32'hc269409b, 32'hc1961efb};
test_output[27752:27759] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27760:27767] = '{32'h4183eb4e, 32'h427a5fdd, 32'hc1526e5e, 32'hc29e9e17, 32'h42c05329, 32'h42149ce0, 32'h40ec988b, 32'h42c69f55};
test_output[27760:27767] = '{32'h4183eb4e, 32'h427a5fdd, 32'h0, 32'h0, 32'h42c05329, 32'h42149ce0, 32'h40ec988b, 32'h42c69f55};
test_input[27768:27775] = '{32'h42c6fe6c, 32'hc2a389d0, 32'hc28623f2, 32'hc1997de4, 32'h42768487, 32'hc166f5d5, 32'h4173bb52, 32'hc20a2055};
test_output[27768:27775] = '{32'h42c6fe6c, 32'h0, 32'h0, 32'h0, 32'h42768487, 32'h0, 32'h4173bb52, 32'h0};
test_input[27776:27783] = '{32'h429a8073, 32'hc205f064, 32'hc265be25, 32'h42a9f83a, 32'h424a6dc5, 32'hc2a8c5da, 32'h422003a5, 32'h41ac5a44};
test_output[27776:27783] = '{32'h429a8073, 32'h0, 32'h0, 32'h42a9f83a, 32'h424a6dc5, 32'h0, 32'h422003a5, 32'h41ac5a44};
test_input[27784:27791] = '{32'hc2b34553, 32'h4277dd2e, 32'hbfedd405, 32'hc23d7566, 32'hc208449f, 32'hc23cc87b, 32'hc22881b0, 32'h422a895c};
test_output[27784:27791] = '{32'h0, 32'h4277dd2e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422a895c};
test_input[27792:27799] = '{32'h41c6a211, 32'h41a14183, 32'hc28c6e43, 32'h41391c29, 32'h42c4f49b, 32'h4257da9f, 32'hc200d560, 32'hc233ee3b};
test_output[27792:27799] = '{32'h41c6a211, 32'h41a14183, 32'h0, 32'h41391c29, 32'h42c4f49b, 32'h4257da9f, 32'h0, 32'h0};
test_input[27800:27807] = '{32'h423ce7ff, 32'hc2a8cd24, 32'h424b98b1, 32'h40ce13dc, 32'h4213748c, 32'h41d467cf, 32'hc2b4b3a5, 32'hc18b2793};
test_output[27800:27807] = '{32'h423ce7ff, 32'h0, 32'h424b98b1, 32'h40ce13dc, 32'h4213748c, 32'h41d467cf, 32'h0, 32'h0};
test_input[27808:27815] = '{32'hc2b6ef84, 32'h429af306, 32'hc1274119, 32'h41b859fd, 32'hc2a010f0, 32'hc246c5ca, 32'hc282cd97, 32'h411dcaef};
test_output[27808:27815] = '{32'h0, 32'h429af306, 32'h0, 32'h41b859fd, 32'h0, 32'h0, 32'h0, 32'h411dcaef};
test_input[27816:27823] = '{32'h426bd4e5, 32'hc213da07, 32'h4267cb58, 32'hc2923608, 32'h41c4f793, 32'h428681a4, 32'hc241bd70, 32'hc22fb3ed};
test_output[27816:27823] = '{32'h426bd4e5, 32'h0, 32'h4267cb58, 32'h0, 32'h41c4f793, 32'h428681a4, 32'h0, 32'h0};
test_input[27824:27831] = '{32'hc29bc0bd, 32'h41164d1b, 32'h429fc8db, 32'hc28bddb2, 32'hc27c10c2, 32'hc2a2de3d, 32'h4110d5c0, 32'h425aed55};
test_output[27824:27831] = '{32'h0, 32'h41164d1b, 32'h429fc8db, 32'h0, 32'h0, 32'h0, 32'h4110d5c0, 32'h425aed55};
test_input[27832:27839] = '{32'h41cb6170, 32'hc28e0a2e, 32'h410eaae4, 32'h41c6de83, 32'h4208b386, 32'h4248ff1f, 32'h4180bcc8, 32'h42885862};
test_output[27832:27839] = '{32'h41cb6170, 32'h0, 32'h410eaae4, 32'h41c6de83, 32'h4208b386, 32'h4248ff1f, 32'h4180bcc8, 32'h42885862};
test_input[27840:27847] = '{32'hc2683dc7, 32'hc2aa3d98, 32'h42b95b87, 32'hc25d7527, 32'h42b73cdd, 32'h425434bb, 32'h42bbbbf2, 32'hc011e3df};
test_output[27840:27847] = '{32'h0, 32'h0, 32'h42b95b87, 32'h0, 32'h42b73cdd, 32'h425434bb, 32'h42bbbbf2, 32'h0};
test_input[27848:27855] = '{32'hc2bbedcd, 32'hc21d3786, 32'hc2964736, 32'h422e2fee, 32'hc2616b0b, 32'hc2954842, 32'h418fed0e, 32'hc1d07071};
test_output[27848:27855] = '{32'h0, 32'h0, 32'h0, 32'h422e2fee, 32'h0, 32'h0, 32'h418fed0e, 32'h0};
test_input[27856:27863] = '{32'hc24266b8, 32'h4026b639, 32'h4212b3fc, 32'hc2401dfc, 32'h41f5deeb, 32'h4193b632, 32'h42b7724a, 32'hc1be3d19};
test_output[27856:27863] = '{32'h0, 32'h4026b639, 32'h4212b3fc, 32'h0, 32'h41f5deeb, 32'h4193b632, 32'h42b7724a, 32'h0};
test_input[27864:27871] = '{32'hc1905ed2, 32'h419c2965, 32'hc2b85f3e, 32'h42298dfb, 32'h42a2cbf2, 32'h426d3a6d, 32'h424ed43f, 32'h4290cadd};
test_output[27864:27871] = '{32'h0, 32'h419c2965, 32'h0, 32'h42298dfb, 32'h42a2cbf2, 32'h426d3a6d, 32'h424ed43f, 32'h4290cadd};
test_input[27872:27879] = '{32'h42079cad, 32'h4233ea34, 32'h41d6a0c8, 32'h42b5c254, 32'hc2549e78, 32'h424dca2d, 32'hc1fb9314, 32'h423fb4a7};
test_output[27872:27879] = '{32'h42079cad, 32'h4233ea34, 32'h41d6a0c8, 32'h42b5c254, 32'h0, 32'h424dca2d, 32'h0, 32'h423fb4a7};
test_input[27880:27887] = '{32'h4102c3f8, 32'h4289088c, 32'h41e661c9, 32'h41c2d9cb, 32'hc1663b40, 32'h429a21c1, 32'h4223a3cb, 32'hc19f12c4};
test_output[27880:27887] = '{32'h4102c3f8, 32'h4289088c, 32'h41e661c9, 32'h41c2d9cb, 32'h0, 32'h429a21c1, 32'h4223a3cb, 32'h0};
test_input[27888:27895] = '{32'hc2a850fe, 32'h410efed7, 32'hc2899bc1, 32'h4250b149, 32'h42aef4e9, 32'h41cab257, 32'hc20f2dfa, 32'hc1428309};
test_output[27888:27895] = '{32'h0, 32'h410efed7, 32'h0, 32'h4250b149, 32'h42aef4e9, 32'h41cab257, 32'h0, 32'h0};
test_input[27896:27903] = '{32'h426dd9ff, 32'hc2a23e3c, 32'hc22316ee, 32'h407967bd, 32'h414ed628, 32'h419244e7, 32'hc27df871, 32'hc20d0c9d};
test_output[27896:27903] = '{32'h426dd9ff, 32'h0, 32'h0, 32'h407967bd, 32'h414ed628, 32'h419244e7, 32'h0, 32'h0};
test_input[27904:27911] = '{32'hc2c73f44, 32'hc24d3b1f, 32'h4265fc02, 32'hc008daca, 32'h41b061a8, 32'h4227262f, 32'h4136a9a0, 32'h4282c506};
test_output[27904:27911] = '{32'h0, 32'h0, 32'h4265fc02, 32'h0, 32'h41b061a8, 32'h4227262f, 32'h4136a9a0, 32'h4282c506};
test_input[27912:27919] = '{32'h420d75ac, 32'hc280a4c2, 32'hc14c3eae, 32'hc2c2f4e9, 32'h42b53806, 32'h409e4763, 32'hc293bc8b, 32'hc2934cc6};
test_output[27912:27919] = '{32'h420d75ac, 32'h0, 32'h0, 32'h0, 32'h42b53806, 32'h409e4763, 32'h0, 32'h0};
test_input[27920:27927] = '{32'hc2b2269f, 32'h42a599dc, 32'hc167a9c7, 32'h42858d29, 32'hc2943a92, 32'h41a908b8, 32'h42c30b56, 32'hc2a04d66};
test_output[27920:27927] = '{32'h0, 32'h42a599dc, 32'h0, 32'h42858d29, 32'h0, 32'h41a908b8, 32'h42c30b56, 32'h0};
test_input[27928:27935] = '{32'h4212d9d4, 32'h421fef35, 32'h42ba3142, 32'h41c64095, 32'h42309659, 32'h4226064a, 32'h42b7ce77, 32'h424f6d55};
test_output[27928:27935] = '{32'h4212d9d4, 32'h421fef35, 32'h42ba3142, 32'h41c64095, 32'h42309659, 32'h4226064a, 32'h42b7ce77, 32'h424f6d55};
test_input[27936:27943] = '{32'h42991b87, 32'h41d50237, 32'h42759476, 32'hc2657b3c, 32'h42bf5aa5, 32'h41b27b4d, 32'hc287ca18, 32'hc299f887};
test_output[27936:27943] = '{32'h42991b87, 32'h41d50237, 32'h42759476, 32'h0, 32'h42bf5aa5, 32'h41b27b4d, 32'h0, 32'h0};
test_input[27944:27951] = '{32'h42309906, 32'hc2a7d7e7, 32'h42bc68d1, 32'h42a449c8, 32'h415248ef, 32'hc2154b0d, 32'h4174476d, 32'h41c89a43};
test_output[27944:27951] = '{32'h42309906, 32'h0, 32'h42bc68d1, 32'h42a449c8, 32'h415248ef, 32'h0, 32'h4174476d, 32'h41c89a43};
test_input[27952:27959] = '{32'h41317a0d, 32'h41d16fec, 32'hc2877cd1, 32'h42b0ed6f, 32'h420b2870, 32'h4249fc37, 32'h41d12ef0, 32'hc2206432};
test_output[27952:27959] = '{32'h41317a0d, 32'h41d16fec, 32'h0, 32'h42b0ed6f, 32'h420b2870, 32'h4249fc37, 32'h41d12ef0, 32'h0};
test_input[27960:27967] = '{32'hc1d0fce2, 32'h41f0ed43, 32'hc2b485b6, 32'h42c49aad, 32'hc20a5ebb, 32'h42b05a45, 32'h4202cfc1, 32'h42b55130};
test_output[27960:27967] = '{32'h0, 32'h41f0ed43, 32'h0, 32'h42c49aad, 32'h0, 32'h42b05a45, 32'h4202cfc1, 32'h42b55130};
test_input[27968:27975] = '{32'hc2a6e476, 32'hc280a9c9, 32'h41d84455, 32'h4259f3be, 32'hc289f29e, 32'h4163b04e, 32'hc288d4e5, 32'hc12a2363};
test_output[27968:27975] = '{32'h0, 32'h0, 32'h41d84455, 32'h4259f3be, 32'h0, 32'h4163b04e, 32'h0, 32'h0};
test_input[27976:27983] = '{32'h42895a17, 32'hc26ab1ca, 32'h42949cd6, 32'hc1f33194, 32'hc1df5131, 32'hc2727e3d, 32'hc29a712a, 32'hc1b852ac};
test_output[27976:27983] = '{32'h42895a17, 32'h0, 32'h42949cd6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[27984:27991] = '{32'hc2062134, 32'hc29de3a7, 32'hc232c41e, 32'hc1cf64d2, 32'hc2bb9228, 32'hc2acdcca, 32'h41320b0f, 32'h42424fb2};
test_output[27984:27991] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41320b0f, 32'h42424fb2};
test_input[27992:27999] = '{32'h429d37de, 32'h42b88322, 32'hc1a2c0dd, 32'hc1fb0291, 32'h4224ee33, 32'h427ac609, 32'hc2aad785, 32'h4200286e};
test_output[27992:27999] = '{32'h429d37de, 32'h42b88322, 32'h0, 32'h0, 32'h4224ee33, 32'h427ac609, 32'h0, 32'h4200286e};
test_input[28000:28007] = '{32'h42179af5, 32'h421657fc, 32'h429b2121, 32'h425c7338, 32'h4206dd74, 32'hc20d03f1, 32'hc16b6394, 32'hc29fbd1e};
test_output[28000:28007] = '{32'h42179af5, 32'h421657fc, 32'h429b2121, 32'h425c7338, 32'h4206dd74, 32'h0, 32'h0, 32'h0};
test_input[28008:28015] = '{32'h42acca65, 32'h42aeca11, 32'hc06b74bd, 32'hc24a1305, 32'h42752dbb, 32'hc286d96c, 32'hc2b6555e, 32'h42c26e4c};
test_output[28008:28015] = '{32'h42acca65, 32'h42aeca11, 32'h0, 32'h0, 32'h42752dbb, 32'h0, 32'h0, 32'h42c26e4c};
test_input[28016:28023] = '{32'h4142d4ef, 32'h421e7db0, 32'hc21292d2, 32'h41f4a752, 32'hc21f7581, 32'hc0c02063, 32'hc19153ba, 32'hc0ec33be};
test_output[28016:28023] = '{32'h4142d4ef, 32'h421e7db0, 32'h0, 32'h41f4a752, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28024:28031] = '{32'h42301936, 32'h40a50888, 32'h4134e00a, 32'h40a8372b, 32'hc22c1b0d, 32'hc14cda3a, 32'hc27b3517, 32'hc14efea1};
test_output[28024:28031] = '{32'h42301936, 32'h40a50888, 32'h4134e00a, 32'h40a8372b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28032:28039] = '{32'h41de27f0, 32'h429fffb8, 32'hc137c6ee, 32'h4230db05, 32'hc2b25dca, 32'h422c85f5, 32'h4297bcac, 32'hc129fde6};
test_output[28032:28039] = '{32'h41de27f0, 32'h429fffb8, 32'h0, 32'h4230db05, 32'h0, 32'h422c85f5, 32'h4297bcac, 32'h0};
test_input[28040:28047] = '{32'h41dfaa1c, 32'hc0490f6f, 32'h427c0080, 32'hc27fa848, 32'hc2580f14, 32'h40ac6d90, 32'hc0416a1f, 32'hc2aab641};
test_output[28040:28047] = '{32'h41dfaa1c, 32'h0, 32'h427c0080, 32'h0, 32'h0, 32'h40ac6d90, 32'h0, 32'h0};
test_input[28048:28055] = '{32'h420abb5f, 32'hc217039a, 32'h4189d007, 32'h425479ec, 32'h424f194b, 32'hc072d55d, 32'hc254e3ed, 32'hc25c1f2d};
test_output[28048:28055] = '{32'h420abb5f, 32'h0, 32'h4189d007, 32'h425479ec, 32'h424f194b, 32'h0, 32'h0, 32'h0};
test_input[28056:28063] = '{32'hc1263753, 32'hc24899ee, 32'h4249bcb1, 32'hc0a847bd, 32'hc23cf24c, 32'h42a021af, 32'h42aeb1a0, 32'hc27c8288};
test_output[28056:28063] = '{32'h0, 32'h0, 32'h4249bcb1, 32'h0, 32'h0, 32'h42a021af, 32'h42aeb1a0, 32'h0};
test_input[28064:28071] = '{32'hc26d6cc7, 32'h42b19d27, 32'h42bdaae4, 32'h419cf0fa, 32'hc2253b47, 32'hc2ab4b3b, 32'hbfb00b2d, 32'hc04bcac1};
test_output[28064:28071] = '{32'h0, 32'h42b19d27, 32'h42bdaae4, 32'h419cf0fa, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28072:28079] = '{32'h41d41d40, 32'hc2a02a03, 32'hc0d8d7fb, 32'h41e4ba79, 32'h42478bfe, 32'hc17aaede, 32'h42b93fe8, 32'h421bb190};
test_output[28072:28079] = '{32'h41d41d40, 32'h0, 32'h0, 32'h41e4ba79, 32'h42478bfe, 32'h0, 32'h42b93fe8, 32'h421bb190};
test_input[28080:28087] = '{32'h426e0066, 32'hc2c315fc, 32'hc2723fc9, 32'hc2a5cbcc, 32'hc22919ba, 32'hc2461e03, 32'h42a89ec5, 32'h42bf366d};
test_output[28080:28087] = '{32'h426e0066, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a89ec5, 32'h42bf366d};
test_input[28088:28095] = '{32'h4208918a, 32'h42441272, 32'hc04dfd24, 32'h41882ccc, 32'hc0e2cd16, 32'h428958b9, 32'h41d10c33, 32'h41ffdd2b};
test_output[28088:28095] = '{32'h4208918a, 32'h42441272, 32'h0, 32'h41882ccc, 32'h0, 32'h428958b9, 32'h41d10c33, 32'h41ffdd2b};
test_input[28096:28103] = '{32'h42b08ba7, 32'h41aed4a8, 32'h414a551e, 32'hc20da994, 32'hc275b9f3, 32'h417cccb4, 32'h3f25ec5e, 32'hc2ad4201};
test_output[28096:28103] = '{32'h42b08ba7, 32'h41aed4a8, 32'h414a551e, 32'h0, 32'h0, 32'h417cccb4, 32'h3f25ec5e, 32'h0};
test_input[28104:28111] = '{32'hc208876c, 32'h418b7ad7, 32'h42a637f4, 32'hc296807e, 32'h42ab3bef, 32'h423ff6fd, 32'h40dac2ba, 32'hc20f9a65};
test_output[28104:28111] = '{32'h0, 32'h418b7ad7, 32'h42a637f4, 32'h0, 32'h42ab3bef, 32'h423ff6fd, 32'h40dac2ba, 32'h0};
test_input[28112:28119] = '{32'hc25bd3f3, 32'hc21d50cc, 32'hc2be8646, 32'hc0f6b9ea, 32'h423af525, 32'hc1cd06b4, 32'hc2a33e16, 32'h41c26877};
test_output[28112:28119] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h423af525, 32'h0, 32'h0, 32'h41c26877};
test_input[28120:28127] = '{32'hc18ba3da, 32'hc29bafec, 32'hc26f2129, 32'hc274e50d, 32'h4251d30e, 32'hc2b25e67, 32'hc2a9f0d2, 32'hc297113c};
test_output[28120:28127] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4251d30e, 32'h0, 32'h0, 32'h0};
test_input[28128:28135] = '{32'h42b520b6, 32'h41a0fa58, 32'hc20ed5b9, 32'hc1ba5d5d, 32'hc209355a, 32'h4210b2c2, 32'h422351e3, 32'hc289bfa1};
test_output[28128:28135] = '{32'h42b520b6, 32'h41a0fa58, 32'h0, 32'h0, 32'h0, 32'h4210b2c2, 32'h422351e3, 32'h0};
test_input[28136:28143] = '{32'h42ae1090, 32'hc1f9a89b, 32'h42882b2e, 32'hc20bb0b4, 32'hc296610c, 32'h4287101a, 32'h406bc130, 32'h413f5ab7};
test_output[28136:28143] = '{32'h42ae1090, 32'h0, 32'h42882b2e, 32'h0, 32'h0, 32'h4287101a, 32'h406bc130, 32'h413f5ab7};
test_input[28144:28151] = '{32'h41e91bd8, 32'hc242b00d, 32'hc1fe8b0b, 32'hc23225da, 32'h4224858e, 32'h40c3b896, 32'h418ff5a3, 32'h412c6a14};
test_output[28144:28151] = '{32'h41e91bd8, 32'h0, 32'h0, 32'h0, 32'h4224858e, 32'h40c3b896, 32'h418ff5a3, 32'h412c6a14};
test_input[28152:28159] = '{32'h42adfb5d, 32'h4261850d, 32'h428efe13, 32'hc22066da, 32'hc26c9cdf, 32'h410e1211, 32'h429dab37, 32'h4258a347};
test_output[28152:28159] = '{32'h42adfb5d, 32'h4261850d, 32'h428efe13, 32'h0, 32'h0, 32'h410e1211, 32'h429dab37, 32'h4258a347};
test_input[28160:28167] = '{32'h41f80eb7, 32'hc277f779, 32'hc248c45a, 32'h426a9330, 32'h427d0e1f, 32'h42c4d886, 32'hc2b50a48, 32'h4283d8d6};
test_output[28160:28167] = '{32'h41f80eb7, 32'h0, 32'h0, 32'h426a9330, 32'h427d0e1f, 32'h42c4d886, 32'h0, 32'h4283d8d6};
test_input[28168:28175] = '{32'h42871624, 32'h42c60c21, 32'hc2b96ef7, 32'h42993074, 32'h41f16ee4, 32'h425630a3, 32'hc2b80ef5, 32'h42c2e8cc};
test_output[28168:28175] = '{32'h42871624, 32'h42c60c21, 32'h0, 32'h42993074, 32'h41f16ee4, 32'h425630a3, 32'h0, 32'h42c2e8cc};
test_input[28176:28183] = '{32'hc204366e, 32'hc2944328, 32'hc2022332, 32'h41ed85c2, 32'hc253b093, 32'hc1e7f94b, 32'h3ef5a61a, 32'hc1a995e2};
test_output[28176:28183] = '{32'h0, 32'h0, 32'h0, 32'h41ed85c2, 32'h0, 32'h0, 32'h3ef5a61a, 32'h0};
test_input[28184:28191] = '{32'hc1b3a76e, 32'h42493767, 32'h416016f7, 32'hc29eecee, 32'hc2c4a475, 32'hc2992426, 32'hc200081c, 32'h427dc744};
test_output[28184:28191] = '{32'h0, 32'h42493767, 32'h416016f7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427dc744};
test_input[28192:28199] = '{32'hc156af67, 32'hc135dbd1, 32'h422e089e, 32'hbf24a306, 32'hc2b5a4ba, 32'h420bcffe, 32'hc29933ff, 32'hc248fb37};
test_output[28192:28199] = '{32'h0, 32'h0, 32'h422e089e, 32'h0, 32'h0, 32'h420bcffe, 32'h0, 32'h0};
test_input[28200:28207] = '{32'hbfb71fdc, 32'h405f65ac, 32'h42b27b4a, 32'h4109fa89, 32'h421b7d89, 32'h40482818, 32'hc2965a0a, 32'hc20e6915};
test_output[28200:28207] = '{32'h0, 32'h405f65ac, 32'h42b27b4a, 32'h4109fa89, 32'h421b7d89, 32'h40482818, 32'h0, 32'h0};
test_input[28208:28215] = '{32'hc28e357a, 32'hc2a2c22f, 32'h424bee25, 32'h417dfcc3, 32'h429b7e90, 32'hc0773c41, 32'h429f6dfc, 32'hc2875534};
test_output[28208:28215] = '{32'h0, 32'h0, 32'h424bee25, 32'h417dfcc3, 32'h429b7e90, 32'h0, 32'h429f6dfc, 32'h0};
test_input[28216:28223] = '{32'h41027155, 32'hc252c099, 32'hc2310900, 32'hc28cb488, 32'h425047c0, 32'h42897a54, 32'hc246df98, 32'hc1975bcb};
test_output[28216:28223] = '{32'h41027155, 32'h0, 32'h0, 32'h0, 32'h425047c0, 32'h42897a54, 32'h0, 32'h0};
test_input[28224:28231] = '{32'hc1d8fe34, 32'hc22c44fc, 32'h42ae4204, 32'h4280efb1, 32'h429f29f2, 32'hc2b800c8, 32'h41e4b346, 32'hc27039bf};
test_output[28224:28231] = '{32'h0, 32'h0, 32'h42ae4204, 32'h4280efb1, 32'h429f29f2, 32'h0, 32'h41e4b346, 32'h0};
test_input[28232:28239] = '{32'hc26ae1f1, 32'hc2c73011, 32'h428fbecf, 32'h421edabb, 32'hc284f5db, 32'h42ae52ca, 32'h41cae36f, 32'hc2b61cc7};
test_output[28232:28239] = '{32'h0, 32'h0, 32'h428fbecf, 32'h421edabb, 32'h0, 32'h42ae52ca, 32'h41cae36f, 32'h0};
test_input[28240:28247] = '{32'h42c491fd, 32'h428e8d04, 32'hc23ba824, 32'h40b29690, 32'h421bd549, 32'h4262e250, 32'h41d1d174, 32'h42810fd7};
test_output[28240:28247] = '{32'h42c491fd, 32'h428e8d04, 32'h0, 32'h40b29690, 32'h421bd549, 32'h4262e250, 32'h41d1d174, 32'h42810fd7};
test_input[28248:28255] = '{32'hc2a86870, 32'hc1afecb4, 32'hc20184dd, 32'hc2ae4d1c, 32'h4173e15c, 32'h426085da, 32'hc2a99fea, 32'h41d6be3f};
test_output[28248:28255] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4173e15c, 32'h426085da, 32'h0, 32'h41d6be3f};
test_input[28256:28263] = '{32'h429606c5, 32'hc2b8168c, 32'h428c8292, 32'h42779fc6, 32'h41b08280, 32'hc20a03f6, 32'h42b46aa3, 32'hc029e699};
test_output[28256:28263] = '{32'h429606c5, 32'h0, 32'h428c8292, 32'h42779fc6, 32'h41b08280, 32'h0, 32'h42b46aa3, 32'h0};
test_input[28264:28271] = '{32'hc29c850b, 32'h4153587d, 32'hc24ef364, 32'h41328092, 32'h40a190ff, 32'h42b5c65e, 32'hc13e4462, 32'hc2c49768};
test_output[28264:28271] = '{32'h0, 32'h4153587d, 32'h0, 32'h41328092, 32'h40a190ff, 32'h42b5c65e, 32'h0, 32'h0};
test_input[28272:28279] = '{32'h427bd8ea, 32'hc130314e, 32'hc227af98, 32'hc21390a8, 32'h42b2ab38, 32'h42b57c74, 32'hc29c517b, 32'h4274aa8c};
test_output[28272:28279] = '{32'h427bd8ea, 32'h0, 32'h0, 32'h0, 32'h42b2ab38, 32'h42b57c74, 32'h0, 32'h4274aa8c};
test_input[28280:28287] = '{32'h42a42361, 32'h41445bb1, 32'h423ad020, 32'hc20d8ab1, 32'h4270faa3, 32'hc07b9a5c, 32'hc2a1afca, 32'hc11d77e9};
test_output[28280:28287] = '{32'h42a42361, 32'h41445bb1, 32'h423ad020, 32'h0, 32'h4270faa3, 32'h0, 32'h0, 32'h0};
test_input[28288:28295] = '{32'h42bc9ac1, 32'h423d9976, 32'hc17367a2, 32'h4285b514, 32'hc2897706, 32'h42288000, 32'h419088a9, 32'hc182a075};
test_output[28288:28295] = '{32'h42bc9ac1, 32'h423d9976, 32'h0, 32'h4285b514, 32'h0, 32'h42288000, 32'h419088a9, 32'h0};
test_input[28296:28303] = '{32'hc29cb446, 32'h4273be94, 32'hc1eead97, 32'hc2917d5b, 32'h418db2b7, 32'hc2b154a4, 32'h42aae8f5, 32'h42319f13};
test_output[28296:28303] = '{32'h0, 32'h4273be94, 32'h0, 32'h0, 32'h418db2b7, 32'h0, 32'h42aae8f5, 32'h42319f13};
test_input[28304:28311] = '{32'hc269371e, 32'hc243e577, 32'hc2288e55, 32'hc265d6ee, 32'hc0596381, 32'hc1b8d514, 32'hc24e62f0, 32'hc2597ed7};
test_output[28304:28311] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28312:28319] = '{32'hc23104e2, 32'h41c4a0b6, 32'hc1b20272, 32'hc1b5774f, 32'hc280e49f, 32'hc1c7d7e4, 32'hc0a423a4, 32'h40b907a3};
test_output[28312:28319] = '{32'h0, 32'h41c4a0b6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40b907a3};
test_input[28320:28327] = '{32'h41824923, 32'h41d4514b, 32'h4286eb40, 32'hc1af841b, 32'h4259e9af, 32'h422d1b36, 32'h42b27608, 32'hc29645c2};
test_output[28320:28327] = '{32'h41824923, 32'h41d4514b, 32'h4286eb40, 32'h0, 32'h4259e9af, 32'h422d1b36, 32'h42b27608, 32'h0};
test_input[28328:28335] = '{32'hc28ea3f7, 32'h4291a3b7, 32'h413084c0, 32'h423b4a2f, 32'hc29b1028, 32'hc2a02fdd, 32'hc251c994, 32'hc1befe0d};
test_output[28328:28335] = '{32'h0, 32'h4291a3b7, 32'h413084c0, 32'h423b4a2f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28336:28343] = '{32'hc1980686, 32'hc1f3936f, 32'hc2b55d78, 32'hc29cc787, 32'hc25e1b34, 32'h4120b6d0, 32'h4283139a, 32'hc2019917};
test_output[28336:28343] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4120b6d0, 32'h4283139a, 32'h0};
test_input[28344:28351] = '{32'hc28505ee, 32'h42807769, 32'hc165a79a, 32'hc24cd1d1, 32'hc2961465, 32'hc1ebfb52, 32'hc0e8bfac, 32'h4258db75};
test_output[28344:28351] = '{32'h0, 32'h42807769, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4258db75};
test_input[28352:28359] = '{32'hc169e479, 32'h41367e94, 32'h429e9109, 32'h41bccb5b, 32'hc21bbe8e, 32'hc1ca194f, 32'h42a51722, 32'hc0bd8ff8};
test_output[28352:28359] = '{32'h0, 32'h41367e94, 32'h429e9109, 32'h41bccb5b, 32'h0, 32'h0, 32'h42a51722, 32'h0};
test_input[28360:28367] = '{32'hc2b88520, 32'h4215e237, 32'h4297477f, 32'h41adbded, 32'hc2990237, 32'hc26cb841, 32'h420507ba, 32'hc2462e87};
test_output[28360:28367] = '{32'h0, 32'h4215e237, 32'h4297477f, 32'h41adbded, 32'h0, 32'h0, 32'h420507ba, 32'h0};
test_input[28368:28375] = '{32'hc2468be9, 32'hc1e199d3, 32'hc1d200b5, 32'hc2853d95, 32'h426e569e, 32'hc1eea845, 32'h41d9f155, 32'h42bb6230};
test_output[28368:28375] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h426e569e, 32'h0, 32'h41d9f155, 32'h42bb6230};
test_input[28376:28383] = '{32'h42a72c7c, 32'h425d9b67, 32'h42601216, 32'h410849ce, 32'hbf8a3998, 32'hc189c69f, 32'hc1de08e1, 32'hc26c2eaa};
test_output[28376:28383] = '{32'h42a72c7c, 32'h425d9b67, 32'h42601216, 32'h410849ce, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28384:28391] = '{32'hc2907a8f, 32'h42154aa5, 32'hc23d9c65, 32'hc2b166fc, 32'h41265dc6, 32'hc256c9af, 32'h4007888f, 32'hc26b05fb};
test_output[28384:28391] = '{32'h0, 32'h42154aa5, 32'h0, 32'h0, 32'h41265dc6, 32'h0, 32'h4007888f, 32'h0};
test_input[28392:28399] = '{32'hc2c285bd, 32'h428ec423, 32'hc285e8bb, 32'h42928e38, 32'h42c27c8a, 32'hc259c595, 32'h41b47439, 32'hc23d266d};
test_output[28392:28399] = '{32'h0, 32'h428ec423, 32'h0, 32'h42928e38, 32'h42c27c8a, 32'h0, 32'h41b47439, 32'h0};
test_input[28400:28407] = '{32'hc24c5d7b, 32'h42c5b96f, 32'hc285b9fc, 32'hc260d019, 32'hbfe80ac1, 32'h426db5ec, 32'h427918d9, 32'h428d7492};
test_output[28400:28407] = '{32'h0, 32'h42c5b96f, 32'h0, 32'h0, 32'h0, 32'h426db5ec, 32'h427918d9, 32'h428d7492};
test_input[28408:28415] = '{32'hc22b1160, 32'hc104c00c, 32'hc2b4d8fc, 32'h3fcca0b5, 32'hc221c6f4, 32'hc2a7845d, 32'h4153b4f9, 32'hc18c1f72};
test_output[28408:28415] = '{32'h0, 32'h0, 32'h0, 32'h3fcca0b5, 32'h0, 32'h0, 32'h4153b4f9, 32'h0};
test_input[28416:28423] = '{32'h42b5ae02, 32'hc1c1dce8, 32'h41057d33, 32'hc267b939, 32'hc29fec6d, 32'h42115930, 32'h423fe95c, 32'h42a9fa09};
test_output[28416:28423] = '{32'h42b5ae02, 32'h0, 32'h41057d33, 32'h0, 32'h0, 32'h42115930, 32'h423fe95c, 32'h42a9fa09};
test_input[28424:28431] = '{32'hc28ff02c, 32'hc273aada, 32'hc24f3c10, 32'h42a635e8, 32'hc28c8db0, 32'h429a1582, 32'hc0bca752, 32'h4193ce52};
test_output[28424:28431] = '{32'h0, 32'h0, 32'h0, 32'h42a635e8, 32'h0, 32'h429a1582, 32'h0, 32'h4193ce52};
test_input[28432:28439] = '{32'hc2136a01, 32'h4212cc3f, 32'h420ce1f7, 32'hc1426ac2, 32'hc257929c, 32'hc1ba1b49, 32'hc1ac05a7, 32'hc13316b7};
test_output[28432:28439] = '{32'h0, 32'h4212cc3f, 32'h420ce1f7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28440:28447] = '{32'hc192978c, 32'hc25e01d6, 32'h418a9315, 32'hc2829f3a, 32'hc2c01631, 32'hc2ab2a27, 32'hc2c2ee91, 32'h4270174a};
test_output[28440:28447] = '{32'h0, 32'h0, 32'h418a9315, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4270174a};
test_input[28448:28455] = '{32'h42b856c3, 32'h42c4a875, 32'h4223226f, 32'hc2ae2784, 32'h4295ff7e, 32'hc20c3f9b, 32'h4286657d, 32'h429fc848};
test_output[28448:28455] = '{32'h42b856c3, 32'h42c4a875, 32'h4223226f, 32'h0, 32'h4295ff7e, 32'h0, 32'h4286657d, 32'h429fc848};
test_input[28456:28463] = '{32'hc27d7608, 32'hc28d3e2f, 32'h42835441, 32'h41bdc202, 32'hc2aa4974, 32'h41a9fb6d, 32'hc1e8c457, 32'hc1cf1e32};
test_output[28456:28463] = '{32'h0, 32'h0, 32'h42835441, 32'h41bdc202, 32'h0, 32'h41a9fb6d, 32'h0, 32'h0};
test_input[28464:28471] = '{32'hc25eb3ee, 32'hc1caa121, 32'hc28083b9, 32'hc27293e3, 32'hc2b8cdb7, 32'h42ba3a04, 32'h42902946, 32'hc2b6f0a9};
test_output[28464:28471] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42ba3a04, 32'h42902946, 32'h0};
test_input[28472:28479] = '{32'h4291b1e1, 32'h42718ad4, 32'h42c246c2, 32'h42990395, 32'h41884e8e, 32'h41c6f73c, 32'hc1525139, 32'hc208eb2b};
test_output[28472:28479] = '{32'h4291b1e1, 32'h42718ad4, 32'h42c246c2, 32'h42990395, 32'h41884e8e, 32'h41c6f73c, 32'h0, 32'h0};
test_input[28480:28487] = '{32'h4251fa1c, 32'hc0fc1d6e, 32'h42c3fd91, 32'hc2ab20e4, 32'h42b92543, 32'hc1829e0d, 32'hc1f9c6fc, 32'hc289fbd4};
test_output[28480:28487] = '{32'h4251fa1c, 32'h0, 32'h42c3fd91, 32'h0, 32'h42b92543, 32'h0, 32'h0, 32'h0};
test_input[28488:28495] = '{32'hc2ae42d2, 32'hc2c1ce6c, 32'hc2021feb, 32'h41abe6d8, 32'hc159927a, 32'h428d1bd1, 32'h405a82b8, 32'h4265a8a9};
test_output[28488:28495] = '{32'h0, 32'h0, 32'h0, 32'h41abe6d8, 32'h0, 32'h428d1bd1, 32'h405a82b8, 32'h4265a8a9};
test_input[28496:28503] = '{32'hc250ae1a, 32'hc2951078, 32'hc0fd8a9a, 32'hc2b5b498, 32'hc2bd6dae, 32'h425b2f60, 32'hc1c77a7a, 32'h420935ce};
test_output[28496:28503] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425b2f60, 32'h0, 32'h420935ce};
test_input[28504:28511] = '{32'hc16f7b1d, 32'hc1f9ece3, 32'hc218f523, 32'h4238a1e4, 32'hc23a1da6, 32'hc2ad02e4, 32'hc0ca222c, 32'hc2a339f7};
test_output[28504:28511] = '{32'h0, 32'h0, 32'h0, 32'h4238a1e4, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28512:28519] = '{32'h4212ddeb, 32'h419fd00d, 32'hc1d888be, 32'hc290355e, 32'hc232bcba, 32'hc1ce3443, 32'h41d198b6, 32'hc18004b5};
test_output[28512:28519] = '{32'h4212ddeb, 32'h419fd00d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41d198b6, 32'h0};
test_input[28520:28527] = '{32'hc1998c46, 32'hc2bc10c2, 32'hc26cffe8, 32'h429e03e5, 32'hc272d2dd, 32'h41da0774, 32'hc2b8a872, 32'hc12097e9};
test_output[28520:28527] = '{32'h0, 32'h0, 32'h0, 32'h429e03e5, 32'h0, 32'h41da0774, 32'h0, 32'h0};
test_input[28528:28535] = '{32'hc2bcd767, 32'hc259d2e7, 32'hc28ffada, 32'h42b3a1a7, 32'hc2955f0a, 32'hc2650894, 32'hc2822ee4, 32'hc26b7575};
test_output[28528:28535] = '{32'h0, 32'h0, 32'h0, 32'h42b3a1a7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28536:28543] = '{32'hc25528a8, 32'h41ee3b40, 32'hc2addadb, 32'hc11b9ac4, 32'hc27cdc75, 32'h418baf53, 32'hc2aca18a, 32'hc2988141};
test_output[28536:28543] = '{32'h0, 32'h41ee3b40, 32'h0, 32'h0, 32'h0, 32'h418baf53, 32'h0, 32'h0};
test_input[28544:28551] = '{32'h425d5612, 32'h4276b1c0, 32'h42affeaf, 32'h429ee2b6, 32'hc1e33405, 32'h42352bc2, 32'hc2942f1a, 32'h42664ca4};
test_output[28544:28551] = '{32'h425d5612, 32'h4276b1c0, 32'h42affeaf, 32'h429ee2b6, 32'h0, 32'h42352bc2, 32'h0, 32'h42664ca4};
test_input[28552:28559] = '{32'hc21e2e68, 32'hc293a7e6, 32'hc27a1ff4, 32'hc19a908b, 32'hc1ebdaf6, 32'hc273700f, 32'h429454c6, 32'hc223d701};
test_output[28552:28559] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429454c6, 32'h0};
test_input[28560:28567] = '{32'hc21dbaca, 32'h427719a0, 32'hc1a4a85d, 32'hc1e33eb2, 32'hc2667a15, 32'h4215d6e5, 32'hc1d8579f, 32'hc2a22014};
test_output[28560:28567] = '{32'h0, 32'h427719a0, 32'h0, 32'h0, 32'h0, 32'h4215d6e5, 32'h0, 32'h0};
test_input[28568:28575] = '{32'h42a2d1ca, 32'h426f8554, 32'h411e8624, 32'h429302a5, 32'hc1ace9c8, 32'h422fefc2, 32'hc1230f3f, 32'hc1b2d056};
test_output[28568:28575] = '{32'h42a2d1ca, 32'h426f8554, 32'h411e8624, 32'h429302a5, 32'h0, 32'h422fefc2, 32'h0, 32'h0};
test_input[28576:28583] = '{32'hc2ab2783, 32'h42a6f9eb, 32'h42ab4c0e, 32'hc2ab99af, 32'hc21c4edb, 32'h40372b04, 32'h4284083e, 32'hc2900001};
test_output[28576:28583] = '{32'h0, 32'h42a6f9eb, 32'h42ab4c0e, 32'h0, 32'h0, 32'h40372b04, 32'h4284083e, 32'h0};
test_input[28584:28591] = '{32'h422d7dff, 32'hc2a9fc40, 32'h425449c3, 32'hc17cffa5, 32'hc21a2904, 32'hc2bd5b91, 32'h41ff1e29, 32'hc0ca2b71};
test_output[28584:28591] = '{32'h422d7dff, 32'h0, 32'h425449c3, 32'h0, 32'h0, 32'h0, 32'h41ff1e29, 32'h0};
test_input[28592:28599] = '{32'h42b95aac, 32'hc111eda3, 32'h42b2ad9c, 32'hc292d608, 32'h427b13f6, 32'hc105e022, 32'hc24c3f96, 32'h42bed736};
test_output[28592:28599] = '{32'h42b95aac, 32'h0, 32'h42b2ad9c, 32'h0, 32'h427b13f6, 32'h0, 32'h0, 32'h42bed736};
test_input[28600:28607] = '{32'hc285e70f, 32'hc23c70d2, 32'h415e1c35, 32'h422107c3, 32'hc174e209, 32'hc25517eb, 32'hc2870405, 32'hc1f7ab65};
test_output[28600:28607] = '{32'h0, 32'h0, 32'h415e1c35, 32'h422107c3, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28608:28615] = '{32'h428b0e16, 32'hc2132a70, 32'hc2473609, 32'h42b04034, 32'hc2682aca, 32'hc210fda0, 32'hc29261d1, 32'h42126305};
test_output[28608:28615] = '{32'h428b0e16, 32'h0, 32'h0, 32'h42b04034, 32'h0, 32'h0, 32'h0, 32'h42126305};
test_input[28616:28623] = '{32'hc25bfa74, 32'hc2a7277c, 32'hc250b947, 32'hc1a1d426, 32'h41ba9bff, 32'hc1e4ae21, 32'h42759d72, 32'h41736989};
test_output[28616:28623] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41ba9bff, 32'h0, 32'h42759d72, 32'h41736989};
test_input[28624:28631] = '{32'hc2706733, 32'h4265b9d2, 32'hc276ec69, 32'hc1722394, 32'h42a2c7dd, 32'hc1d57a83, 32'h41c28e36, 32'hc2524425};
test_output[28624:28631] = '{32'h0, 32'h4265b9d2, 32'h0, 32'h0, 32'h42a2c7dd, 32'h0, 32'h41c28e36, 32'h0};
test_input[28632:28639] = '{32'hc18ea2d5, 32'h41c5e6a1, 32'h421b96ca, 32'h425794ce, 32'hc1735b09, 32'h41492c2c, 32'h419d333e, 32'hc1a01bcb};
test_output[28632:28639] = '{32'h0, 32'h41c5e6a1, 32'h421b96ca, 32'h425794ce, 32'h0, 32'h41492c2c, 32'h419d333e, 32'h0};
test_input[28640:28647] = '{32'h42c775d0, 32'h41aa2ea3, 32'hc1493781, 32'hc18c3836, 32'hc2bd090f, 32'hc263b9d4, 32'hc298304f, 32'hc0755777};
test_output[28640:28647] = '{32'h42c775d0, 32'h41aa2ea3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28648:28655] = '{32'hc1ba451e, 32'hc2449fdf, 32'h42954642, 32'h420d3df3, 32'h42a27c97, 32'hc2ba97ef, 32'hc27c4afe, 32'h421a3044};
test_output[28648:28655] = '{32'h0, 32'h0, 32'h42954642, 32'h420d3df3, 32'h42a27c97, 32'h0, 32'h0, 32'h421a3044};
test_input[28656:28663] = '{32'hc18850e3, 32'hc29d5a85, 32'hc2a2fafc, 32'hc27dbdc7, 32'h41939842, 32'hc1833694, 32'h418fdfe9, 32'h422fa72b};
test_output[28656:28663] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41939842, 32'h0, 32'h418fdfe9, 32'h422fa72b};
test_input[28664:28671] = '{32'hc28d5ac5, 32'h42a541bc, 32'hc1f928bc, 32'hc17dcd80, 32'h42a75127, 32'hc14ab8c2, 32'hc26f237e, 32'hc2a33a67};
test_output[28664:28671] = '{32'h0, 32'h42a541bc, 32'h0, 32'h0, 32'h42a75127, 32'h0, 32'h0, 32'h0};
test_input[28672:28679] = '{32'h429f2c44, 32'hc2803b5d, 32'h426ab7c2, 32'hc2a272b6, 32'hc2b02add, 32'hc2b042f9, 32'h41d8f96a, 32'hc24db432};
test_output[28672:28679] = '{32'h429f2c44, 32'h0, 32'h426ab7c2, 32'h0, 32'h0, 32'h0, 32'h41d8f96a, 32'h0};
test_input[28680:28687] = '{32'h41266e45, 32'h42907496, 32'h42695a92, 32'hc2c28a44, 32'h4211f516, 32'hc208be98, 32'h42b45ffe, 32'hc2a0dc22};
test_output[28680:28687] = '{32'h41266e45, 32'h42907496, 32'h42695a92, 32'h0, 32'h4211f516, 32'h0, 32'h42b45ffe, 32'h0};
test_input[28688:28695] = '{32'hc2b8bdfc, 32'h429b5bd8, 32'hc2ba5dd2, 32'h411c20f3, 32'h41d87a2b, 32'hc2299b93, 32'h42103581, 32'h42b023a4};
test_output[28688:28695] = '{32'h0, 32'h429b5bd8, 32'h0, 32'h411c20f3, 32'h41d87a2b, 32'h0, 32'h42103581, 32'h42b023a4};
test_input[28696:28703] = '{32'h42af323a, 32'hc2a58848, 32'hbfa29d37, 32'h42ab1cb1, 32'h4220ff72, 32'h41d1484a, 32'hc23487c3, 32'hc1fa8fae};
test_output[28696:28703] = '{32'h42af323a, 32'h0, 32'h0, 32'h42ab1cb1, 32'h4220ff72, 32'h41d1484a, 32'h0, 32'h0};
test_input[28704:28711] = '{32'hc2063415, 32'h42c1dd9a, 32'h42b256a6, 32'h4283954e, 32'h40d62e44, 32'hc1c649cb, 32'hc2684e45, 32'hc1b67a25};
test_output[28704:28711] = '{32'h0, 32'h42c1dd9a, 32'h42b256a6, 32'h4283954e, 32'h40d62e44, 32'h0, 32'h0, 32'h0};
test_input[28712:28719] = '{32'hc2bf9a6f, 32'h41774a22, 32'hc238f258, 32'h42bda164, 32'hc22c37e0, 32'h42518475, 32'hc21d0f68, 32'hc26b3a9c};
test_output[28712:28719] = '{32'h0, 32'h41774a22, 32'h0, 32'h42bda164, 32'h0, 32'h42518475, 32'h0, 32'h0};
test_input[28720:28727] = '{32'hc0091974, 32'hc231587b, 32'h41f74387, 32'h42aa2e16, 32'hc0de3d53, 32'h41730e88, 32'hc2b2006f, 32'h42b6a1f3};
test_output[28720:28727] = '{32'h0, 32'h0, 32'h41f74387, 32'h42aa2e16, 32'h0, 32'h41730e88, 32'h0, 32'h42b6a1f3};
test_input[28728:28735] = '{32'h4210eb1f, 32'hc24f7f2c, 32'hc22d4983, 32'hc2135b4c, 32'hc29fd354, 32'hc21cf0a7, 32'h410f628d, 32'h42740eb9};
test_output[28728:28735] = '{32'h4210eb1f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h410f628d, 32'h42740eb9};
test_input[28736:28743] = '{32'hc2433576, 32'h423406f6, 32'hc1b89613, 32'h4106a6dc, 32'h42308fb5, 32'h42afdbea, 32'h4206f11c, 32'h42b65d8a};
test_output[28736:28743] = '{32'h0, 32'h423406f6, 32'h0, 32'h4106a6dc, 32'h42308fb5, 32'h42afdbea, 32'h4206f11c, 32'h42b65d8a};
test_input[28744:28751] = '{32'h41baf536, 32'h41c92f17, 32'h41b1325b, 32'hc1a3e115, 32'h42835680, 32'h42b6e8f5, 32'hc21ff29d, 32'h41ebde0b};
test_output[28744:28751] = '{32'h41baf536, 32'h41c92f17, 32'h41b1325b, 32'h0, 32'h42835680, 32'h42b6e8f5, 32'h0, 32'h41ebde0b};
test_input[28752:28759] = '{32'hc181fd3c, 32'h426c5091, 32'hc0920d81, 32'h42c0876e, 32'hc2a12726, 32'h4268a27d, 32'hc26f4637, 32'h422ab1fa};
test_output[28752:28759] = '{32'h0, 32'h426c5091, 32'h0, 32'h42c0876e, 32'h0, 32'h4268a27d, 32'h0, 32'h422ab1fa};
test_input[28760:28767] = '{32'h4287e963, 32'h413d3bee, 32'h41bf324d, 32'hc21904c8, 32'hc2409845, 32'hc0c95c5e, 32'h40d6ea48, 32'h4191be67};
test_output[28760:28767] = '{32'h4287e963, 32'h413d3bee, 32'h41bf324d, 32'h0, 32'h0, 32'h0, 32'h40d6ea48, 32'h4191be67};
test_input[28768:28775] = '{32'h400846b5, 32'h4292d8dc, 32'h41aa65b2, 32'hc22f488b, 32'h428d252b, 32'h417dd8c9, 32'h42aaad74, 32'hc24fee36};
test_output[28768:28775] = '{32'h400846b5, 32'h4292d8dc, 32'h41aa65b2, 32'h0, 32'h428d252b, 32'h417dd8c9, 32'h42aaad74, 32'h0};
test_input[28776:28783] = '{32'hc26c9eaf, 32'h42161abe, 32'hc1bf2eef, 32'h4228f08a, 32'hc292a3fc, 32'h410fdc0c, 32'hc299334a, 32'hc18e5576};
test_output[28776:28783] = '{32'h0, 32'h42161abe, 32'h0, 32'h4228f08a, 32'h0, 32'h410fdc0c, 32'h0, 32'h0};
test_input[28784:28791] = '{32'h40a5df1d, 32'hc23c22cb, 32'h42917263, 32'hc2a9646f, 32'h42b20b9c, 32'h42c27fbb, 32'hc2123869, 32'hc1b722d1};
test_output[28784:28791] = '{32'h40a5df1d, 32'h0, 32'h42917263, 32'h0, 32'h42b20b9c, 32'h42c27fbb, 32'h0, 32'h0};
test_input[28792:28799] = '{32'h42a2138c, 32'hc214eb81, 32'h4248998d, 32'hc1ffd17b, 32'h41a8cd2a, 32'hc112070c, 32'hc29f903a, 32'hc20b8e26};
test_output[28792:28799] = '{32'h42a2138c, 32'h0, 32'h4248998d, 32'h0, 32'h41a8cd2a, 32'h0, 32'h0, 32'h0};
test_input[28800:28807] = '{32'hc2ba2bd2, 32'h42c772d7, 32'hc1d4405f, 32'hc1e370a7, 32'hc266b646, 32'hc279b5ea, 32'h42954875, 32'hc1bfb49d};
test_output[28800:28807] = '{32'h0, 32'h42c772d7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42954875, 32'h0};
test_input[28808:28815] = '{32'hc273b829, 32'hc1978c35, 32'hc1c964c0, 32'h4289e1f5, 32'hc1d42c75, 32'h42b7786d, 32'hc21c92f7, 32'hc28fe0fe};
test_output[28808:28815] = '{32'h0, 32'h0, 32'h0, 32'h4289e1f5, 32'h0, 32'h42b7786d, 32'h0, 32'h0};
test_input[28816:28823] = '{32'h41708cac, 32'hc297b98b, 32'h412944f5, 32'h41fd0c11, 32'h42c058a8, 32'h4234a2b7, 32'h4268296a, 32'hc1141ef4};
test_output[28816:28823] = '{32'h41708cac, 32'h0, 32'h412944f5, 32'h41fd0c11, 32'h42c058a8, 32'h4234a2b7, 32'h4268296a, 32'h0};
test_input[28824:28831] = '{32'h4134e232, 32'hc2989384, 32'hc1897996, 32'hc2989beb, 32'h417501a3, 32'hc28958a1, 32'h4268cd85, 32'h420508f7};
test_output[28824:28831] = '{32'h4134e232, 32'h0, 32'h0, 32'h0, 32'h417501a3, 32'h0, 32'h4268cd85, 32'h420508f7};
test_input[28832:28839] = '{32'hc2a9fa51, 32'h4107d449, 32'hc19fcfdb, 32'hc220242c, 32'hc2c5ef46, 32'hc1b878aa, 32'hc284684e, 32'hc0c6e4c1};
test_output[28832:28839] = '{32'h0, 32'h4107d449, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28840:28847] = '{32'hc216849c, 32'h4299e7ec, 32'h424a3f8c, 32'h42ba66f3, 32'h421405d2, 32'h424e7030, 32'hc24c4c12, 32'hc297ff8c};
test_output[28840:28847] = '{32'h0, 32'h4299e7ec, 32'h424a3f8c, 32'h42ba66f3, 32'h421405d2, 32'h424e7030, 32'h0, 32'h0};
test_input[28848:28855] = '{32'hc286b35f, 32'h42ad41ad, 32'h42801c79, 32'h4260a70c, 32'hc291bd7f, 32'hc274cb85, 32'h4222a0c5, 32'hc2466012};
test_output[28848:28855] = '{32'h0, 32'h42ad41ad, 32'h42801c79, 32'h4260a70c, 32'h0, 32'h0, 32'h4222a0c5, 32'h0};
test_input[28856:28863] = '{32'h422743ae, 32'h42b4d982, 32'h421a967f, 32'hc1be4e9f, 32'hc29457f6, 32'h403a56f7, 32'h4270094a, 32'hc28dfc66};
test_output[28856:28863] = '{32'h422743ae, 32'h42b4d982, 32'h421a967f, 32'h0, 32'h0, 32'h403a56f7, 32'h4270094a, 32'h0};
test_input[28864:28871] = '{32'hc254b68f, 32'hc1e0ea1b, 32'hc227556e, 32'h41c5a1b8, 32'hc2ab466e, 32'hc230748a, 32'hc0ed6b37, 32'hc2b092e5};
test_output[28864:28871] = '{32'h0, 32'h0, 32'h0, 32'h41c5a1b8, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28872:28879] = '{32'hc2b7b99b, 32'h427f7eea, 32'h42700db8, 32'hc296c539, 32'hc25925fc, 32'h42b6859a, 32'hc29f8c88, 32'hc20ba9ee};
test_output[28872:28879] = '{32'h0, 32'h427f7eea, 32'h42700db8, 32'h0, 32'h0, 32'h42b6859a, 32'h0, 32'h0};
test_input[28880:28887] = '{32'h4275ee76, 32'h424e3f63, 32'hc25e9682, 32'hc244d3ed, 32'h414da597, 32'h41e4ec4c, 32'h42a75f86, 32'hc271164d};
test_output[28880:28887] = '{32'h4275ee76, 32'h424e3f63, 32'h0, 32'h0, 32'h414da597, 32'h41e4ec4c, 32'h42a75f86, 32'h0};
test_input[28888:28895] = '{32'hc285b9da, 32'h41d1240f, 32'h425b3e25, 32'hc24c69b7, 32'h40811520, 32'hc23d7296, 32'h42973f79, 32'hc29268be};
test_output[28888:28895] = '{32'h0, 32'h41d1240f, 32'h425b3e25, 32'h0, 32'h40811520, 32'h0, 32'h42973f79, 32'h0};
test_input[28896:28903] = '{32'hc206bd0d, 32'h42b39d3f, 32'h429466a2, 32'h41f71b41, 32'h413e0373, 32'hc26bc72b, 32'h41cb1953, 32'hc2a0f781};
test_output[28896:28903] = '{32'h0, 32'h42b39d3f, 32'h429466a2, 32'h41f71b41, 32'h413e0373, 32'h0, 32'h41cb1953, 32'h0};
test_input[28904:28911] = '{32'h42a07298, 32'hc164b847, 32'h428e65db, 32'h424bf284, 32'h42b36e93, 32'hc2c0ffed, 32'h41c30b0a, 32'hc1ca4838};
test_output[28904:28911] = '{32'h42a07298, 32'h0, 32'h428e65db, 32'h424bf284, 32'h42b36e93, 32'h0, 32'h41c30b0a, 32'h0};
test_input[28912:28919] = '{32'hc1d7f875, 32'hc269186a, 32'hc29c618d, 32'hc287cdb9, 32'hc23ff2ac, 32'hc2c1acaa, 32'hbe32ca00, 32'hc18ca37a};
test_output[28912:28919] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[28920:28927] = '{32'h42754b01, 32'h42bd839d, 32'hc2b15a19, 32'h41fa76db, 32'h42bd0648, 32'h424b110e, 32'h4281c5ba, 32'h42b88891};
test_output[28920:28927] = '{32'h42754b01, 32'h42bd839d, 32'h0, 32'h41fa76db, 32'h42bd0648, 32'h424b110e, 32'h4281c5ba, 32'h42b88891};
test_input[28928:28935] = '{32'hc289ea3b, 32'h42c653bf, 32'h418578f5, 32'hc1b6e91a, 32'hc2c134ea, 32'hc242ffa3, 32'h41ae2e82, 32'h42013591};
test_output[28928:28935] = '{32'h0, 32'h42c653bf, 32'h418578f5, 32'h0, 32'h0, 32'h0, 32'h41ae2e82, 32'h42013591};
test_input[28936:28943] = '{32'hc29f61f9, 32'hc2c6a229, 32'hc2c4e84b, 32'hbf1fa0d3, 32'hc1987ff0, 32'h42bfedbc, 32'h42857b4d, 32'h4163a603};
test_output[28936:28943] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bfedbc, 32'h42857b4d, 32'h4163a603};
test_input[28944:28951] = '{32'h42a3917e, 32'hc25eb668, 32'hc241f45f, 32'h4244a479, 32'h4218ceff, 32'hc1ac43b9, 32'h424510c9, 32'hc22a5014};
test_output[28944:28951] = '{32'h42a3917e, 32'h0, 32'h0, 32'h4244a479, 32'h4218ceff, 32'h0, 32'h424510c9, 32'h0};
test_input[28952:28959] = '{32'hc1dcd32d, 32'hc20ff6c6, 32'hc23d41c3, 32'hc24eaddb, 32'hc29ffa62, 32'h41983d0d, 32'hc26a9e8c, 32'h40a4db09};
test_output[28952:28959] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41983d0d, 32'h0, 32'h40a4db09};
test_input[28960:28967] = '{32'h41889f90, 32'h40678f5f, 32'hc28b7190, 32'hc20798a5, 32'h3fc9f4e7, 32'h42749025, 32'h42553154, 32'hc28d6e88};
test_output[28960:28967] = '{32'h41889f90, 32'h40678f5f, 32'h0, 32'h0, 32'h3fc9f4e7, 32'h42749025, 32'h42553154, 32'h0};
test_input[28968:28975] = '{32'h42844ff0, 32'h42bda366, 32'h42179841, 32'h42c61d02, 32'hc2906c1e, 32'hc214973f, 32'h403165eb, 32'h41c75f56};
test_output[28968:28975] = '{32'h42844ff0, 32'h42bda366, 32'h42179841, 32'h42c61d02, 32'h0, 32'h0, 32'h403165eb, 32'h41c75f56};
test_input[28976:28983] = '{32'h429f6871, 32'hc2a54b4c, 32'h42336e26, 32'h424ac33f, 32'hc28323dc, 32'hc2203898, 32'h429e5673, 32'h42c7bcd1};
test_output[28976:28983] = '{32'h429f6871, 32'h0, 32'h42336e26, 32'h424ac33f, 32'h0, 32'h0, 32'h429e5673, 32'h42c7bcd1};
test_input[28984:28991] = '{32'h4294d8ab, 32'hc262c1aa, 32'h42c25608, 32'h417febfb, 32'h414ccde5, 32'h4149689c, 32'h420998e7, 32'h41bdf7db};
test_output[28984:28991] = '{32'h4294d8ab, 32'h0, 32'h42c25608, 32'h417febfb, 32'h414ccde5, 32'h4149689c, 32'h420998e7, 32'h41bdf7db};
test_input[28992:28999] = '{32'h42bf47c8, 32'h42452078, 32'h42aaa21c, 32'hc1721846, 32'hc0cd413f, 32'hc2510ed8, 32'h42bf6f25, 32'h429c7096};
test_output[28992:28999] = '{32'h42bf47c8, 32'h42452078, 32'h42aaa21c, 32'h0, 32'h0, 32'h0, 32'h42bf6f25, 32'h429c7096};
test_input[29000:29007] = '{32'h424206a4, 32'h419ced67, 32'hc246af30, 32'h420a777d, 32'h4284f008, 32'h41049f18, 32'h41cd455a, 32'h4198ad82};
test_output[29000:29007] = '{32'h424206a4, 32'h419ced67, 32'h0, 32'h420a777d, 32'h4284f008, 32'h41049f18, 32'h41cd455a, 32'h4198ad82};
test_input[29008:29015] = '{32'hc280bff0, 32'h41b3a54e, 32'hc218c2f7, 32'h42266dae, 32'hc2a5dad3, 32'h40e3eca8, 32'hc219ef22, 32'hc29449b3};
test_output[29008:29015] = '{32'h0, 32'h41b3a54e, 32'h0, 32'h42266dae, 32'h0, 32'h40e3eca8, 32'h0, 32'h0};
test_input[29016:29023] = '{32'h42058563, 32'hc2658529, 32'hc1ed6ec7, 32'hc11c38b3, 32'hc09615cb, 32'hc1f43f8e, 32'h40bd41d1, 32'h42460514};
test_output[29016:29023] = '{32'h42058563, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40bd41d1, 32'h42460514};
test_input[29024:29031] = '{32'h42c36fef, 32'hc2045ee8, 32'h429141b1, 32'hc106e625, 32'h410cbe34, 32'hc0672b19, 32'hbde047b1, 32'h424a58a5};
test_output[29024:29031] = '{32'h42c36fef, 32'h0, 32'h429141b1, 32'h0, 32'h410cbe34, 32'h0, 32'h0, 32'h424a58a5};
test_input[29032:29039] = '{32'hc28b685f, 32'h4158ffc1, 32'hc2774e01, 32'h42459834, 32'h40cda8e7, 32'hc2ad7acb, 32'h42bd8aa8, 32'h42905534};
test_output[29032:29039] = '{32'h0, 32'h4158ffc1, 32'h0, 32'h42459834, 32'h40cda8e7, 32'h0, 32'h42bd8aa8, 32'h42905534};
test_input[29040:29047] = '{32'hc1514a3a, 32'hc22c35ea, 32'hc2a6b2a2, 32'h41232b97, 32'hc04fda69, 32'h42b73753, 32'h4288a982, 32'h42483613};
test_output[29040:29047] = '{32'h0, 32'h0, 32'h0, 32'h41232b97, 32'h0, 32'h42b73753, 32'h4288a982, 32'h42483613};
test_input[29048:29055] = '{32'h42c786ef, 32'h427c8815, 32'hc1025e75, 32'h4284cdc5, 32'hc28e0b58, 32'hc2c1df85, 32'hc2a685e4, 32'hc2430503};
test_output[29048:29055] = '{32'h42c786ef, 32'h427c8815, 32'h0, 32'h4284cdc5, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29056:29063] = '{32'h426da601, 32'hc2b6c94e, 32'hc2123c92, 32'hc24d1922, 32'h420289fc, 32'hc22dcd24, 32'h4224141b, 32'h42920aee};
test_output[29056:29063] = '{32'h426da601, 32'h0, 32'h0, 32'h0, 32'h420289fc, 32'h0, 32'h4224141b, 32'h42920aee};
test_input[29064:29071] = '{32'hc2030f59, 32'h425f3f6f, 32'h42145004, 32'hc2885489, 32'hc1f84bed, 32'h3ef8d281, 32'hc23bc49c, 32'h423049ed};
test_output[29064:29071] = '{32'h0, 32'h425f3f6f, 32'h42145004, 32'h0, 32'h0, 32'h3ef8d281, 32'h0, 32'h423049ed};
test_input[29072:29079] = '{32'hc21c95a9, 32'h42800bf8, 32'hc2b9cd5a, 32'hc28f70b2, 32'h412967bb, 32'hc29addc0, 32'hc250cac5, 32'h4164434f};
test_output[29072:29079] = '{32'h0, 32'h42800bf8, 32'h0, 32'h0, 32'h412967bb, 32'h0, 32'h0, 32'h4164434f};
test_input[29080:29087] = '{32'h4244f4fb, 32'hc247138b, 32'h429c7a93, 32'h4203829c, 32'hc1d8ec83, 32'h429e2d58, 32'hc0ac739d, 32'h418656d0};
test_output[29080:29087] = '{32'h4244f4fb, 32'h0, 32'h429c7a93, 32'h4203829c, 32'h0, 32'h429e2d58, 32'h0, 32'h418656d0};
test_input[29088:29095] = '{32'hc2b9103c, 32'hc295943a, 32'h41f92685, 32'h4280a367, 32'hc148c3a2, 32'h428f4b68, 32'h42c734c3, 32'h4210152b};
test_output[29088:29095] = '{32'h0, 32'h0, 32'h41f92685, 32'h4280a367, 32'h0, 32'h428f4b68, 32'h42c734c3, 32'h4210152b};
test_input[29096:29103] = '{32'hc23e117e, 32'hc292e0a7, 32'hc1f1f0d9, 32'h42ac55ff, 32'hc283b876, 32'hc1efae1f, 32'h42ad1bc5, 32'h42b3a45a};
test_output[29096:29103] = '{32'h0, 32'h0, 32'h0, 32'h42ac55ff, 32'h0, 32'h0, 32'h42ad1bc5, 32'h42b3a45a};
test_input[29104:29111] = '{32'h423bc571, 32'hc15362a3, 32'h40f6a818, 32'hc204f15b, 32'hc29201b1, 32'hc296595a, 32'h42bad741, 32'h428425ad};
test_output[29104:29111] = '{32'h423bc571, 32'h0, 32'h40f6a818, 32'h0, 32'h0, 32'h0, 32'h42bad741, 32'h428425ad};
test_input[29112:29119] = '{32'hc280f8ed, 32'hc2160bb0, 32'hc1feb19f, 32'h4216d9a5, 32'h418b95b4, 32'hc2a8e872, 32'hc29f0a5a, 32'h42852367};
test_output[29112:29119] = '{32'h0, 32'h0, 32'h0, 32'h4216d9a5, 32'h418b95b4, 32'h0, 32'h0, 32'h42852367};
test_input[29120:29127] = '{32'hc2bb8fc8, 32'h4253416f, 32'h42a6019d, 32'h42720a8d, 32'h41686f2c, 32'hc17fb403, 32'hc294b64b, 32'hc1a44328};
test_output[29120:29127] = '{32'h0, 32'h4253416f, 32'h42a6019d, 32'h42720a8d, 32'h41686f2c, 32'h0, 32'h0, 32'h0};
test_input[29128:29135] = '{32'hc2b5def8, 32'h41133b48, 32'hc296ebac, 32'h41d3d873, 32'hc1b2aeb8, 32'h40cd173f, 32'hc2a311b1, 32'hc2a665ee};
test_output[29128:29135] = '{32'h0, 32'h41133b48, 32'h0, 32'h41d3d873, 32'h0, 32'h40cd173f, 32'h0, 32'h0};
test_input[29136:29143] = '{32'h425ca836, 32'hc2abfa46, 32'h428a4293, 32'hc2b12686, 32'hc0b603f6, 32'h4184241d, 32'h42b4c317, 32'h42aef95a};
test_output[29136:29143] = '{32'h425ca836, 32'h0, 32'h428a4293, 32'h0, 32'h0, 32'h4184241d, 32'h42b4c317, 32'h42aef95a};
test_input[29144:29151] = '{32'hc2c62fff, 32'h4279f517, 32'h41ff8173, 32'hc1faccdb, 32'h422ca8ab, 32'hc1d9556e, 32'h42c2c7cd, 32'h42194a39};
test_output[29144:29151] = '{32'h0, 32'h4279f517, 32'h41ff8173, 32'h0, 32'h422ca8ab, 32'h0, 32'h42c2c7cd, 32'h42194a39};
test_input[29152:29159] = '{32'hc28358a5, 32'hc268efd1, 32'h424f1c93, 32'h424a02a0, 32'h424f885f, 32'h42b130d5, 32'h4231a7f4, 32'hc2a16263};
test_output[29152:29159] = '{32'h0, 32'h0, 32'h424f1c93, 32'h424a02a0, 32'h424f885f, 32'h42b130d5, 32'h4231a7f4, 32'h0};
test_input[29160:29167] = '{32'hc1ac44d9, 32'hc1095ed1, 32'hc2ae9f30, 32'h41278973, 32'h4104f983, 32'h42924f9b, 32'h42701ae0, 32'hc2a99cd3};
test_output[29160:29167] = '{32'h0, 32'h0, 32'h0, 32'h41278973, 32'h4104f983, 32'h42924f9b, 32'h42701ae0, 32'h0};
test_input[29168:29175] = '{32'h423a4794, 32'hc25f0477, 32'hc1e14e94, 32'h4284060c, 32'hc24ab8cc, 32'h4278191f, 32'h4298a3ae, 32'h410ac78d};
test_output[29168:29175] = '{32'h423a4794, 32'h0, 32'h0, 32'h4284060c, 32'h0, 32'h4278191f, 32'h4298a3ae, 32'h410ac78d};
test_input[29176:29183] = '{32'hc25b93b6, 32'hc1b5ca78, 32'hc235c90c, 32'h427065ce, 32'h42b6c181, 32'h42838c37, 32'h3ed92e9e, 32'h41ed9d4f};
test_output[29176:29183] = '{32'h0, 32'h0, 32'h0, 32'h427065ce, 32'h42b6c181, 32'h42838c37, 32'h3ed92e9e, 32'h41ed9d4f};
test_input[29184:29191] = '{32'h42a1fbd8, 32'h411c6458, 32'hc21c7a1a, 32'h42488fc0, 32'hc21af6eb, 32'h427931cc, 32'h421e6650, 32'h421edb7b};
test_output[29184:29191] = '{32'h42a1fbd8, 32'h411c6458, 32'h0, 32'h42488fc0, 32'h0, 32'h427931cc, 32'h421e6650, 32'h421edb7b};
test_input[29192:29199] = '{32'h4214262e, 32'hc192ab15, 32'h42a35c89, 32'h42a676a5, 32'hc2bfdd05, 32'hc27c9d17, 32'h41a0acd8, 32'h422c8a2f};
test_output[29192:29199] = '{32'h4214262e, 32'h0, 32'h42a35c89, 32'h42a676a5, 32'h0, 32'h0, 32'h41a0acd8, 32'h422c8a2f};
test_input[29200:29207] = '{32'hc27bac57, 32'hc2b82719, 32'hc1fe37e2, 32'h42620315, 32'h41f5117b, 32'hc2b81a06, 32'hc2916147, 32'hc20bde33};
test_output[29200:29207] = '{32'h0, 32'h0, 32'h0, 32'h42620315, 32'h41f5117b, 32'h0, 32'h0, 32'h0};
test_input[29208:29215] = '{32'hc1dd58dc, 32'hc1b55cef, 32'hc2b28138, 32'hc2bd47b9, 32'hc0f1302e, 32'h40b3699c, 32'h40a90e35, 32'h424e1af2};
test_output[29208:29215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40b3699c, 32'h40a90e35, 32'h424e1af2};
test_input[29216:29223] = '{32'h4269f5e2, 32'h42376e12, 32'hc2844c16, 32'h42b952df, 32'h40f0ca69, 32'h427ea977, 32'hc29a318e, 32'h4216b0dc};
test_output[29216:29223] = '{32'h4269f5e2, 32'h42376e12, 32'h0, 32'h42b952df, 32'h40f0ca69, 32'h427ea977, 32'h0, 32'h4216b0dc};
test_input[29224:29231] = '{32'h41d3234a, 32'h428b8130, 32'h4172f6c6, 32'h42b34ab4, 32'hc21849bb, 32'h4287e7b0, 32'hc2608780, 32'hc1a4e195};
test_output[29224:29231] = '{32'h41d3234a, 32'h428b8130, 32'h4172f6c6, 32'h42b34ab4, 32'h0, 32'h4287e7b0, 32'h0, 32'h0};
test_input[29232:29239] = '{32'hc28a94b3, 32'hc08c30ba, 32'h42b9f471, 32'h427f7414, 32'hc2580cc3, 32'hc194674a, 32'hc28d3f27, 32'h4212d4f4};
test_output[29232:29239] = '{32'h0, 32'h0, 32'h42b9f471, 32'h427f7414, 32'h0, 32'h0, 32'h0, 32'h4212d4f4};
test_input[29240:29247] = '{32'hc213ef14, 32'h42838dcc, 32'h42095573, 32'h4068d7cc, 32'h42c596da, 32'h42823a11, 32'h423587d7, 32'hc0fda99d};
test_output[29240:29247] = '{32'h0, 32'h42838dcc, 32'h42095573, 32'h4068d7cc, 32'h42c596da, 32'h42823a11, 32'h423587d7, 32'h0};
test_input[29248:29255] = '{32'hc1193ada, 32'hbf1c34c4, 32'h41526645, 32'hc2233323, 32'h42889594, 32'h421d8f91, 32'h426f5f15, 32'h4178e4c3};
test_output[29248:29255] = '{32'h0, 32'h0, 32'h41526645, 32'h0, 32'h42889594, 32'h421d8f91, 32'h426f5f15, 32'h4178e4c3};
test_input[29256:29263] = '{32'hc29dfb6b, 32'h4298e7de, 32'hc282add2, 32'h42c776ff, 32'h421bbc8a, 32'hc2a4ba6a, 32'h41acd780, 32'hc20f76b4};
test_output[29256:29263] = '{32'h0, 32'h4298e7de, 32'h0, 32'h42c776ff, 32'h421bbc8a, 32'h0, 32'h41acd780, 32'h0};
test_input[29264:29271] = '{32'h427dd02c, 32'h4291385c, 32'hc222b795, 32'hc25e1534, 32'hc2b0ffd7, 32'hc2a5b867, 32'h42a5c205, 32'hc204e0ce};
test_output[29264:29271] = '{32'h427dd02c, 32'h4291385c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a5c205, 32'h0};
test_input[29272:29279] = '{32'h401eceb6, 32'h42b08bac, 32'h42339512, 32'h42909027, 32'h428219fc, 32'hc1fcde2e, 32'h42a45fca, 32'hc209dfa2};
test_output[29272:29279] = '{32'h401eceb6, 32'h42b08bac, 32'h42339512, 32'h42909027, 32'h428219fc, 32'h0, 32'h42a45fca, 32'h0};
test_input[29280:29287] = '{32'hc2570683, 32'hc23b6d1a, 32'hc282295e, 32'hc18dff7e, 32'h413e2330, 32'h40ad889c, 32'hc28245d0, 32'h4097157e};
test_output[29280:29287] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h413e2330, 32'h40ad889c, 32'h0, 32'h4097157e};
test_input[29288:29295] = '{32'h422485a6, 32'h42aa3c27, 32'h42ae726a, 32'hc264fcdc, 32'h419cfca2, 32'hc248a0a0, 32'h4281b306, 32'hc0ac5162};
test_output[29288:29295] = '{32'h422485a6, 32'h42aa3c27, 32'h42ae726a, 32'h0, 32'h419cfca2, 32'h0, 32'h4281b306, 32'h0};
test_input[29296:29303] = '{32'hc2b0d19b, 32'hc1599058, 32'hc297165c, 32'h41b30102, 32'hc1fad8c5, 32'hc2c00dcf, 32'h42aef51a, 32'hc2bf10ac};
test_output[29296:29303] = '{32'h0, 32'h0, 32'h0, 32'h41b30102, 32'h0, 32'h0, 32'h42aef51a, 32'h0};
test_input[29304:29311] = '{32'h41801f76, 32'hc2b824e0, 32'h41958939, 32'h42621288, 32'h42b043c4, 32'h41b73129, 32'hc22d256f, 32'hc208d2c6};
test_output[29304:29311] = '{32'h41801f76, 32'h0, 32'h41958939, 32'h42621288, 32'h42b043c4, 32'h41b73129, 32'h0, 32'h0};
test_input[29312:29319] = '{32'hc1e3b78a, 32'hc2b267f8, 32'h429bd6c1, 32'hc22df3db, 32'h4226223c, 32'hc25e71b2, 32'hc2a9a13e, 32'hc1b22c61};
test_output[29312:29319] = '{32'h0, 32'h0, 32'h429bd6c1, 32'h0, 32'h4226223c, 32'h0, 32'h0, 32'h0};
test_input[29320:29327] = '{32'hc2a05b0c, 32'h42b9eca9, 32'hc0aa6966, 32'h41fc9815, 32'h427610b9, 32'hc2b7ea85, 32'h4288af1b, 32'h426594d6};
test_output[29320:29327] = '{32'h0, 32'h42b9eca9, 32'h0, 32'h41fc9815, 32'h427610b9, 32'h0, 32'h4288af1b, 32'h426594d6};
test_input[29328:29335] = '{32'hc29363ff, 32'h423a3ab9, 32'h42441874, 32'hc2b620f5, 32'h418ea30d, 32'h41d39ffb, 32'h423a422f, 32'h424f2d1c};
test_output[29328:29335] = '{32'h0, 32'h423a3ab9, 32'h42441874, 32'h0, 32'h418ea30d, 32'h41d39ffb, 32'h423a422f, 32'h424f2d1c};
test_input[29336:29343] = '{32'hc21d6497, 32'hc253ef06, 32'hc270f407, 32'h40994f98, 32'hc267a28d, 32'h4250d643, 32'hc22665a6, 32'h4084c705};
test_output[29336:29343] = '{32'h0, 32'h0, 32'h0, 32'h40994f98, 32'h0, 32'h4250d643, 32'h0, 32'h4084c705};
test_input[29344:29351] = '{32'hc08b0cb0, 32'h42be2259, 32'hc296763c, 32'h42372162, 32'h42c16cb0, 32'h426e1832, 32'h41e583e6, 32'h4093b2ad};
test_output[29344:29351] = '{32'h0, 32'h42be2259, 32'h0, 32'h42372162, 32'h42c16cb0, 32'h426e1832, 32'h41e583e6, 32'h4093b2ad};
test_input[29352:29359] = '{32'hc24f8e4e, 32'hc27877c7, 32'h41a1fa4f, 32'h41d32dec, 32'h42902b32, 32'h42b6ed3b, 32'hc298ca00, 32'h423e7dbb};
test_output[29352:29359] = '{32'h0, 32'h0, 32'h41a1fa4f, 32'h41d32dec, 32'h42902b32, 32'h42b6ed3b, 32'h0, 32'h423e7dbb};
test_input[29360:29367] = '{32'h429add6d, 32'h42c32ddf, 32'hc19dbf07, 32'hc167b73b, 32'h4238f362, 32'hc269b60d, 32'hc26eb780, 32'hc2b98e91};
test_output[29360:29367] = '{32'h429add6d, 32'h42c32ddf, 32'h0, 32'h0, 32'h4238f362, 32'h0, 32'h0, 32'h0};
test_input[29368:29375] = '{32'hc2b3a8f6, 32'hbf959ab6, 32'h420ab42b, 32'hbf04dfe6, 32'hc236dadb, 32'hc2c527f7, 32'h4210d31e, 32'hc21eda92};
test_output[29368:29375] = '{32'h0, 32'h0, 32'h420ab42b, 32'h0, 32'h0, 32'h0, 32'h4210d31e, 32'h0};
test_input[29376:29383] = '{32'h42b8f74b, 32'h41ad60a6, 32'h415dd642, 32'h42b5ae7d, 32'h42bda8ab, 32'h41782a29, 32'h425207b6, 32'h41c82b74};
test_output[29376:29383] = '{32'h42b8f74b, 32'h41ad60a6, 32'h415dd642, 32'h42b5ae7d, 32'h42bda8ab, 32'h41782a29, 32'h425207b6, 32'h41c82b74};
test_input[29384:29391] = '{32'h41d86b69, 32'h41b462a9, 32'hc25a097b, 32'hc022b790, 32'hc28be698, 32'hc2941405, 32'h4140aa40, 32'h423f76c9};
test_output[29384:29391] = '{32'h41d86b69, 32'h41b462a9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4140aa40, 32'h423f76c9};
test_input[29392:29399] = '{32'h41b6d9a0, 32'hc1b79114, 32'h429f8044, 32'h41873e8c, 32'hc2b850b5, 32'hc2b3dd43, 32'h42a828b2, 32'h4265a71f};
test_output[29392:29399] = '{32'h41b6d9a0, 32'h0, 32'h429f8044, 32'h41873e8c, 32'h0, 32'h0, 32'h42a828b2, 32'h4265a71f};
test_input[29400:29407] = '{32'hc1e8eaa9, 32'hc28eb067, 32'hc2b78350, 32'h428581f4, 32'h42bc7031, 32'hc28e3244, 32'hc11f1cde, 32'hc271eb78};
test_output[29400:29407] = '{32'h0, 32'h0, 32'h0, 32'h428581f4, 32'h42bc7031, 32'h0, 32'h0, 32'h0};
test_input[29408:29415] = '{32'hc1e49caa, 32'h429fd0de, 32'h41a595bd, 32'hc20118cc, 32'hc10f78f0, 32'h41f2a6b2, 32'hc283c645, 32'hc253bab1};
test_output[29408:29415] = '{32'h0, 32'h429fd0de, 32'h41a595bd, 32'h0, 32'h0, 32'h41f2a6b2, 32'h0, 32'h0};
test_input[29416:29423] = '{32'hc1380952, 32'h40e56c36, 32'h4235c3e4, 32'h4114febf, 32'h42c53975, 32'h426515ed, 32'hc26a8843, 32'hc22ff724};
test_output[29416:29423] = '{32'h0, 32'h40e56c36, 32'h4235c3e4, 32'h4114febf, 32'h42c53975, 32'h426515ed, 32'h0, 32'h0};
test_input[29424:29431] = '{32'hc22e5356, 32'h41fe9444, 32'h4243d61e, 32'hc271081d, 32'hc2979d8c, 32'h3fddc00d, 32'h412c8c3b, 32'hc2619b10};
test_output[29424:29431] = '{32'h0, 32'h41fe9444, 32'h4243d61e, 32'h0, 32'h0, 32'h3fddc00d, 32'h412c8c3b, 32'h0};
test_input[29432:29439] = '{32'hc1926b6d, 32'hc101e6f4, 32'h401c1183, 32'h42188089, 32'h4237cede, 32'h427e1f77, 32'h42c3a6bf, 32'hc1f08ac0};
test_output[29432:29439] = '{32'h0, 32'h0, 32'h401c1183, 32'h42188089, 32'h4237cede, 32'h427e1f77, 32'h42c3a6bf, 32'h0};
test_input[29440:29447] = '{32'h423c1cfa, 32'hc23e2628, 32'h42557423, 32'hc2123763, 32'h42868707, 32'h42c3db44, 32'h3ffede50, 32'hc183fca4};
test_output[29440:29447] = '{32'h423c1cfa, 32'h0, 32'h42557423, 32'h0, 32'h42868707, 32'h42c3db44, 32'h3ffede50, 32'h0};
test_input[29448:29455] = '{32'h425e2ffb, 32'hc22fe8d8, 32'hc2af8f33, 32'hc1c6ed45, 32'hc0b94c3b, 32'hc2071475, 32'h4159583e, 32'h429bc7b5};
test_output[29448:29455] = '{32'h425e2ffb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4159583e, 32'h429bc7b5};
test_input[29456:29463] = '{32'h42a4a67b, 32'hc2174103, 32'h4240544d, 32'hc2b23094, 32'hc19b4471, 32'h428941ef, 32'hc2aeb79f, 32'hc2879a71};
test_output[29456:29463] = '{32'h42a4a67b, 32'h0, 32'h4240544d, 32'h0, 32'h0, 32'h428941ef, 32'h0, 32'h0};
test_input[29464:29471] = '{32'hc1187c94, 32'hc0faab90, 32'h41f367f3, 32'h421c1be9, 32'hc2bc7bb7, 32'hc1a2b8fb, 32'hc0b01989, 32'hc213d5b7};
test_output[29464:29471] = '{32'h0, 32'h0, 32'h41f367f3, 32'h421c1be9, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[29472:29479] = '{32'h42bb64ab, 32'hbeabea1e, 32'h41bb8ae6, 32'hc11442a5, 32'h4224bf7e, 32'hc28d02a9, 32'hc2483b8b, 32'h4293f26f};
test_output[29472:29479] = '{32'h42bb64ab, 32'h0, 32'h41bb8ae6, 32'h0, 32'h4224bf7e, 32'h0, 32'h0, 32'h4293f26f};
test_input[29480:29487] = '{32'h4271da98, 32'hc2b94f50, 32'hc274ae6a, 32'h4296fe7e, 32'hc2a7f8ea, 32'h3e99a8ab, 32'h4292adbe, 32'hc270f30d};
test_output[29480:29487] = '{32'h4271da98, 32'h0, 32'h0, 32'h4296fe7e, 32'h0, 32'h3e99a8ab, 32'h4292adbe, 32'h0};
test_input[29488:29495] = '{32'hc2aaebad, 32'hc2aaec44, 32'hc28ff9a0, 32'hc23b3aba, 32'hc0d351c1, 32'hc1a09ca5, 32'hc2c03e9d, 32'h41917e06};
test_output[29488:29495] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41917e06};
test_input[29496:29503] = '{32'hc23183d5, 32'h41ea87b8, 32'h41f7491e, 32'hc27d6370, 32'h42a74c0c, 32'h42b47873, 32'h403f934d, 32'h426867d8};
test_output[29496:29503] = '{32'h0, 32'h41ea87b8, 32'h41f7491e, 32'h0, 32'h42a74c0c, 32'h42b47873, 32'h403f934d, 32'h426867d8};
test_input[29504:29511] = '{32'h42a663cc, 32'h41ed6fdd, 32'hc28a02ca, 32'h423f58b9, 32'hc1bbb433, 32'h42c1f82c, 32'h41c863b5, 32'hc1b1711d};
test_output[29504:29511] = '{32'h42a663cc, 32'h41ed6fdd, 32'h0, 32'h423f58b9, 32'h0, 32'h42c1f82c, 32'h41c863b5, 32'h0};
test_input[29512:29519] = '{32'h420b6769, 32'h429b38b1, 32'h42c7b2ac, 32'hc2a6f256, 32'hc2c52fd0, 32'h42a6f48b, 32'h418ce15e, 32'hc218d566};
test_output[29512:29519] = '{32'h420b6769, 32'h429b38b1, 32'h42c7b2ac, 32'h0, 32'h0, 32'h42a6f48b, 32'h418ce15e, 32'h0};
test_input[29520:29527] = '{32'hc2a8a964, 32'h4123b20a, 32'hc22c8a88, 32'h41803f32, 32'hc0fa92f8, 32'hc2471be9, 32'hc2b46170, 32'h421a54ab};
test_output[29520:29527] = '{32'h0, 32'h4123b20a, 32'h0, 32'h41803f32, 32'h0, 32'h0, 32'h0, 32'h421a54ab};
test_input[29528:29535] = '{32'h41bb731a, 32'h4273bc2c, 32'hc2552d81, 32'hc074132a, 32'h4284056c, 32'h42a7e3d5, 32'hc02a743a, 32'h4239077b};
test_output[29528:29535] = '{32'h41bb731a, 32'h4273bc2c, 32'h0, 32'h0, 32'h4284056c, 32'h42a7e3d5, 32'h0, 32'h4239077b};
test_input[29536:29543] = '{32'hc245335b, 32'h424baf2d, 32'hc2615b54, 32'hc29f466f, 32'hc1d876b0, 32'h427d370b, 32'hc23ab89b, 32'h4260b715};
test_output[29536:29543] = '{32'h0, 32'h424baf2d, 32'h0, 32'h0, 32'h0, 32'h427d370b, 32'h0, 32'h4260b715};
test_input[29544:29551] = '{32'hc2a11d2f, 32'hc193e51a, 32'hc22562ff, 32'h41dabee8, 32'h4237aefa, 32'hc22bd8a1, 32'h41a63558, 32'h41a14db1};
test_output[29544:29551] = '{32'h0, 32'h0, 32'h0, 32'h41dabee8, 32'h4237aefa, 32'h0, 32'h41a63558, 32'h41a14db1};
test_input[29552:29559] = '{32'h42b51874, 32'h42b9486e, 32'h41ee4154, 32'h41de1c59, 32'h423474e1, 32'h41e62922, 32'h42578758, 32'h4287eaac};
test_output[29552:29559] = '{32'h42b51874, 32'h42b9486e, 32'h41ee4154, 32'h41de1c59, 32'h423474e1, 32'h41e62922, 32'h42578758, 32'h4287eaac};
test_input[29560:29567] = '{32'h4266a245, 32'h42390d34, 32'h419aedf8, 32'hc141b1a9, 32'hc227ff6f, 32'h41ff544b, 32'h4184df04, 32'h418aca1e};
test_output[29560:29567] = '{32'h4266a245, 32'h42390d34, 32'h419aedf8, 32'h0, 32'h0, 32'h41ff544b, 32'h4184df04, 32'h418aca1e};
test_input[29568:29575] = '{32'h42401ae6, 32'hc2c7a3bd, 32'h42a01c59, 32'h413a15fd, 32'hc2acf83e, 32'hc25edd50, 32'h42a6f21c, 32'hc1f360ac};
test_output[29568:29575] = '{32'h42401ae6, 32'h0, 32'h42a01c59, 32'h413a15fd, 32'h0, 32'h0, 32'h42a6f21c, 32'h0};
test_input[29576:29583] = '{32'hc2b07613, 32'hc2532e2c, 32'hc2912f95, 32'hc2765d68, 32'hc21d51cb, 32'h41ff1834, 32'h424952d1, 32'hc240453f};
test_output[29576:29583] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ff1834, 32'h424952d1, 32'h0};
test_input[29584:29591] = '{32'h41bca1a4, 32'hc29c6281, 32'h428df994, 32'hc2748b31, 32'hc298ba3c, 32'hc1d55788, 32'h42bae77f, 32'hc2676b86};
test_output[29584:29591] = '{32'h41bca1a4, 32'h0, 32'h428df994, 32'h0, 32'h0, 32'h0, 32'h42bae77f, 32'h0};
test_input[29592:29599] = '{32'h425cdcc2, 32'h423b59f0, 32'hc290d1da, 32'hc2a6b774, 32'h412e1dab, 32'hc244fb58, 32'hc2209f13, 32'h4227ba2b};
test_output[29592:29599] = '{32'h425cdcc2, 32'h423b59f0, 32'h0, 32'h0, 32'h412e1dab, 32'h0, 32'h0, 32'h4227ba2b};
test_input[29600:29607] = '{32'h429ba8df, 32'h420d893b, 32'h42a83833, 32'hc28a2503, 32'h42632a57, 32'h412e8f61, 32'hc1d42185, 32'hc2be1753};
test_output[29600:29607] = '{32'h429ba8df, 32'h420d893b, 32'h42a83833, 32'h0, 32'h42632a57, 32'h412e8f61, 32'h0, 32'h0};
test_input[29608:29615] = '{32'hc2b05fc6, 32'h42b67481, 32'h42192774, 32'hc141252f, 32'hc239e733, 32'hc209ff25, 32'hc23f4426, 32'h4273a650};
test_output[29608:29615] = '{32'h0, 32'h42b67481, 32'h42192774, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4273a650};
test_input[29616:29623] = '{32'hc225b79f, 32'hc1f70e97, 32'hc27af948, 32'h42aa084d, 32'hc211c4b7, 32'hc19809fd, 32'h42c18e74, 32'hc2a26207};
test_output[29616:29623] = '{32'h0, 32'h0, 32'h0, 32'h42aa084d, 32'h0, 32'h0, 32'h42c18e74, 32'h0};
test_input[29624:29631] = '{32'hc2b0f3a4, 32'h428d8950, 32'h41ecb013, 32'h41cda8e2, 32'h42901261, 32'h40acf89c, 32'h42af8244, 32'hc1b0b0f8};
test_output[29624:29631] = '{32'h0, 32'h428d8950, 32'h41ecb013, 32'h41cda8e2, 32'h42901261, 32'h40acf89c, 32'h42af8244, 32'h0};
test_input[29632:29639] = '{32'hc2c4c499, 32'hc2006905, 32'h42bca6dc, 32'h410b8ca1, 32'hc2646270, 32'hc2b73444, 32'h429cd647, 32'hc26ce4bd};
test_output[29632:29639] = '{32'h0, 32'h0, 32'h42bca6dc, 32'h410b8ca1, 32'h0, 32'h0, 32'h429cd647, 32'h0};
test_input[29640:29647] = '{32'h429beade, 32'h415f096f, 32'h419e240b, 32'hc1993fd2, 32'hc2999ef4, 32'hc2497336, 32'hc216e932, 32'h418ead43};
test_output[29640:29647] = '{32'h429beade, 32'h415f096f, 32'h419e240b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h418ead43};
test_input[29648:29655] = '{32'h417b8beb, 32'hc1cd63fb, 32'h4248f309, 32'hc19f055c, 32'hc00937ca, 32'hc20c1344, 32'h422c1560, 32'h429b9bd2};
test_output[29648:29655] = '{32'h417b8beb, 32'h0, 32'h4248f309, 32'h0, 32'h0, 32'h0, 32'h422c1560, 32'h429b9bd2};
test_input[29656:29663] = '{32'hc2865eb8, 32'hc285cde1, 32'h4217e33b, 32'hc0fd1796, 32'hc0d86768, 32'h423b504e, 32'hc1ea8a04, 32'hc23cddbc};
test_output[29656:29663] = '{32'h0, 32'h0, 32'h4217e33b, 32'h0, 32'h0, 32'h423b504e, 32'h0, 32'h0};
test_input[29664:29671] = '{32'h4285c9bf, 32'h428ccc50, 32'h41cbc9c7, 32'h418ddf28, 32'hc27ca568, 32'h41f7e801, 32'h42bf16e9, 32'hc282e45e};
test_output[29664:29671] = '{32'h4285c9bf, 32'h428ccc50, 32'h41cbc9c7, 32'h418ddf28, 32'h0, 32'h41f7e801, 32'h42bf16e9, 32'h0};
test_input[29672:29679] = '{32'h40044157, 32'h4272b536, 32'hc07f6f9f, 32'h42a4d10f, 32'h41d45f1b, 32'hc14729ab, 32'hc0b9189d, 32'hc2acf99c};
test_output[29672:29679] = '{32'h40044157, 32'h4272b536, 32'h0, 32'h42a4d10f, 32'h41d45f1b, 32'h0, 32'h0, 32'h0};
test_input[29680:29687] = '{32'hc2b32023, 32'h428aaa50, 32'h42058f79, 32'hc1a49a63, 32'h42b5bb43, 32'h42af3e36, 32'h427c8696, 32'hc19dc450};
test_output[29680:29687] = '{32'h0, 32'h428aaa50, 32'h42058f79, 32'h0, 32'h42b5bb43, 32'h42af3e36, 32'h427c8696, 32'h0};
test_input[29688:29695] = '{32'hc1c289b0, 32'hc237c4dc, 32'hc24e3c7a, 32'h429f3b0d, 32'h42717673, 32'h42619025, 32'hc0cde99e, 32'h40527f48};
test_output[29688:29695] = '{32'h0, 32'h0, 32'h0, 32'h429f3b0d, 32'h42717673, 32'h42619025, 32'h0, 32'h40527f48};
test_input[29696:29703] = '{32'hc2219bf4, 32'h4225495a, 32'hc28347e6, 32'h424c55c0, 32'h41a9831f, 32'hc0abf3e4, 32'hc279d8c7, 32'hc1c7d7d5};
test_output[29696:29703] = '{32'h0, 32'h4225495a, 32'h0, 32'h424c55c0, 32'h41a9831f, 32'h0, 32'h0, 32'h0};
test_input[29704:29711] = '{32'hc1c4cbb3, 32'hc1c00913, 32'hc2b934d8, 32'hc22e6c85, 32'h42a72599, 32'h4200d645, 32'hc0ddac16, 32'h4293e249};
test_output[29704:29711] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a72599, 32'h4200d645, 32'h0, 32'h4293e249};
test_input[29712:29719] = '{32'h40c95581, 32'hc267c026, 32'hc1fe975a, 32'hc248db71, 32'h4148ce88, 32'h4260a1aa, 32'hc23fa046, 32'h41bff041};
test_output[29712:29719] = '{32'h40c95581, 32'h0, 32'h0, 32'h0, 32'h4148ce88, 32'h4260a1aa, 32'h0, 32'h41bff041};
test_input[29720:29727] = '{32'h42a795bf, 32'hc2616bfc, 32'hc26d8470, 32'h41288676, 32'hc1dfd25b, 32'h428ef117, 32'hc1d3e7db, 32'hc2455e5c};
test_output[29720:29727] = '{32'h42a795bf, 32'h0, 32'h0, 32'h41288676, 32'h0, 32'h428ef117, 32'h0, 32'h0};
test_input[29728:29735] = '{32'hc2a26d2b, 32'hc18c73cb, 32'h427c77b8, 32'hc27ab176, 32'h42474a02, 32'h42309633, 32'hc1f0f6e4, 32'h41f2590f};
test_output[29728:29735] = '{32'h0, 32'h0, 32'h427c77b8, 32'h0, 32'h42474a02, 32'h42309633, 32'h0, 32'h41f2590f};
test_input[29736:29743] = '{32'h412b01e5, 32'h429ae859, 32'hc1f3cd77, 32'h406f657f, 32'hc1438150, 32'hc27aa0e9, 32'h42becc88, 32'h4246b6cc};
test_output[29736:29743] = '{32'h412b01e5, 32'h429ae859, 32'h0, 32'h406f657f, 32'h0, 32'h0, 32'h42becc88, 32'h4246b6cc};
test_input[29744:29751] = '{32'hc276dd8a, 32'h42814358, 32'hbfefea78, 32'hc29272b3, 32'h429978f8, 32'h42ae51f8, 32'hc2a964e5, 32'h428de425};
test_output[29744:29751] = '{32'h0, 32'h42814358, 32'h0, 32'h0, 32'h429978f8, 32'h42ae51f8, 32'h0, 32'h428de425};
test_input[29752:29759] = '{32'hc19b160d, 32'h41f8d5cd, 32'h42788d09, 32'hc25916a4, 32'hc2924370, 32'h429d9a00, 32'hc285e277, 32'hc1864f38};
test_output[29752:29759] = '{32'h0, 32'h41f8d5cd, 32'h42788d09, 32'h0, 32'h0, 32'h429d9a00, 32'h0, 32'h0};
test_input[29760:29767] = '{32'hc25e67f4, 32'h41de21e6, 32'h429930a2, 32'hc1a1cec4, 32'hbde00ec1, 32'h42c4942e, 32'h42950b2a, 32'h4294f006};
test_output[29760:29767] = '{32'h0, 32'h41de21e6, 32'h429930a2, 32'h0, 32'h0, 32'h42c4942e, 32'h42950b2a, 32'h4294f006};
test_input[29768:29775] = '{32'hc2a65797, 32'h42ab066f, 32'h41c7b2ae, 32'hc2a3ff91, 32'h4293c3ed, 32'h42a831d1, 32'h420e2bf9, 32'hc19a6522};
test_output[29768:29775] = '{32'h0, 32'h42ab066f, 32'h41c7b2ae, 32'h0, 32'h4293c3ed, 32'h42a831d1, 32'h420e2bf9, 32'h0};
test_input[29776:29783] = '{32'h428895af, 32'h421bf3a8, 32'h4178260a, 32'h4299f352, 32'h41bd79d4, 32'h429f3578, 32'h4221e714, 32'h424fce16};
test_output[29776:29783] = '{32'h428895af, 32'h421bf3a8, 32'h4178260a, 32'h4299f352, 32'h41bd79d4, 32'h429f3578, 32'h4221e714, 32'h424fce16};
test_input[29784:29791] = '{32'h41e81b53, 32'h42afe2c3, 32'h4227048b, 32'hc266999b, 32'hc1b789fc, 32'hc1bd1ae7, 32'h428a306b, 32'h428e0d7c};
test_output[29784:29791] = '{32'h41e81b53, 32'h42afe2c3, 32'h4227048b, 32'h0, 32'h0, 32'h0, 32'h428a306b, 32'h428e0d7c};
test_input[29792:29799] = '{32'hc24fc248, 32'hc29495c0, 32'h4226febb, 32'hc2af5324, 32'hc21ae448, 32'h42c1d9c8, 32'hc299d75d, 32'h404b9eed};
test_output[29792:29799] = '{32'h0, 32'h0, 32'h4226febb, 32'h0, 32'h0, 32'h42c1d9c8, 32'h0, 32'h404b9eed};
test_input[29800:29807] = '{32'h4298bdd5, 32'h41ad6db0, 32'hc2839e08, 32'h41a68fd4, 32'hc2942448, 32'hc286e976, 32'hc2102677, 32'h4262e622};
test_output[29800:29807] = '{32'h4298bdd5, 32'h41ad6db0, 32'h0, 32'h41a68fd4, 32'h0, 32'h0, 32'h0, 32'h4262e622};
test_input[29808:29815] = '{32'hc1e6cd14, 32'hc2964262, 32'h40ead328, 32'hc2bce656, 32'hc2c4f2db, 32'h428c6ec2, 32'hc25da7ba, 32'h42b4ba95};
test_output[29808:29815] = '{32'h0, 32'h0, 32'h40ead328, 32'h0, 32'h0, 32'h428c6ec2, 32'h0, 32'h42b4ba95};
test_input[29816:29823] = '{32'hc231808b, 32'h428a05db, 32'h42aefeab, 32'h42c66c2e, 32'h42bb80ff, 32'h42bcb6bb, 32'h420a5bab, 32'hc2bf8d47};
test_output[29816:29823] = '{32'h0, 32'h428a05db, 32'h42aefeab, 32'h42c66c2e, 32'h42bb80ff, 32'h42bcb6bb, 32'h420a5bab, 32'h0};
test_input[29824:29831] = '{32'hc0b72de5, 32'hc2192d6c, 32'h4251ebf3, 32'hc2b0d83c, 32'h423568e5, 32'hc115a462, 32'h429b9a68, 32'h429f76af};
test_output[29824:29831] = '{32'h0, 32'h0, 32'h4251ebf3, 32'h0, 32'h423568e5, 32'h0, 32'h429b9a68, 32'h429f76af};
test_input[29832:29839] = '{32'hc26c20f9, 32'h42bc4bf2, 32'h41c08067, 32'hc2c1fd51, 32'h42917d84, 32'h425c5936, 32'h422ecbe8, 32'hc2713cdc};
test_output[29832:29839] = '{32'h0, 32'h42bc4bf2, 32'h41c08067, 32'h0, 32'h42917d84, 32'h425c5936, 32'h422ecbe8, 32'h0};
test_input[29840:29847] = '{32'hc2bd36c3, 32'hc290fb05, 32'h409200c2, 32'h42b2324d, 32'h429c4fac, 32'hc204a03c, 32'h4287e741, 32'h40d46f5a};
test_output[29840:29847] = '{32'h0, 32'h0, 32'h409200c2, 32'h42b2324d, 32'h429c4fac, 32'h0, 32'h4287e741, 32'h40d46f5a};
test_input[29848:29855] = '{32'hc251ee7c, 32'hc19ba306, 32'hc0fe45cb, 32'hc2b94480, 32'h3f65c9c9, 32'hc23fbbf9, 32'h427dbd58, 32'hc2589a34};
test_output[29848:29855] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h3f65c9c9, 32'h0, 32'h427dbd58, 32'h0};
test_input[29856:29863] = '{32'hc271866d, 32'h4136107b, 32'h41b93600, 32'h3d18803e, 32'hc1feb68f, 32'h42205c35, 32'hc21516ee, 32'h41f0eb4c};
test_output[29856:29863] = '{32'h0, 32'h4136107b, 32'h41b93600, 32'h3d18803e, 32'h0, 32'h42205c35, 32'h0, 32'h41f0eb4c};
test_input[29864:29871] = '{32'hc2a1686c, 32'hc25c3f76, 32'h420ec187, 32'h4212467c, 32'hc2865b54, 32'h429f940a, 32'h429b2ad8, 32'hc1330d83};
test_output[29864:29871] = '{32'h0, 32'h0, 32'h420ec187, 32'h4212467c, 32'h0, 32'h429f940a, 32'h429b2ad8, 32'h0};
test_input[29872:29879] = '{32'h42943521, 32'h41518ea6, 32'hc2059d4b, 32'hc1ed289a, 32'hc212d47b, 32'hc2684860, 32'hc2c21172, 32'h415a6fb8};
test_output[29872:29879] = '{32'h42943521, 32'h41518ea6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h415a6fb8};
test_input[29880:29887] = '{32'hc2497cfd, 32'hc20c22b6, 32'h3e0df8bb, 32'hc295ee98, 32'hc29de543, 32'h42c2f450, 32'h423f0226, 32'hc02eff0f};
test_output[29880:29887] = '{32'h0, 32'h0, 32'h3e0df8bb, 32'h0, 32'h0, 32'h42c2f450, 32'h423f0226, 32'h0};
test_input[29888:29895] = '{32'hc28edf1e, 32'h4285cdd9, 32'hc018c938, 32'hc292f401, 32'hc2aa0dc3, 32'h42a68ec8, 32'hc299b19a, 32'hc1b4996e};
test_output[29888:29895] = '{32'h0, 32'h4285cdd9, 32'h0, 32'h0, 32'h0, 32'h42a68ec8, 32'h0, 32'h0};
test_input[29896:29903] = '{32'hc2b40514, 32'hc23b5ea8, 32'hc2353adb, 32'h42b76871, 32'h429c5b13, 32'h4269d516, 32'h4205fb78, 32'h429fdb48};
test_output[29896:29903] = '{32'h0, 32'h0, 32'h0, 32'h42b76871, 32'h429c5b13, 32'h4269d516, 32'h4205fb78, 32'h429fdb48};
test_input[29904:29911] = '{32'hc219e150, 32'hc2bf36b3, 32'h4092591f, 32'hc2a97916, 32'h41660885, 32'h421fb3ba, 32'hc1e9e8e1, 32'hc227dd86};
test_output[29904:29911] = '{32'h0, 32'h0, 32'h4092591f, 32'h0, 32'h41660885, 32'h421fb3ba, 32'h0, 32'h0};
test_input[29912:29919] = '{32'hc1f787dc, 32'hc0c7354b, 32'hc2103776, 32'hc2c12ced, 32'h4003b87a, 32'hc250f18b, 32'hc21c3daf, 32'hc0aae129};
test_output[29912:29919] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4003b87a, 32'h0, 32'h0, 32'h0};
test_input[29920:29927] = '{32'hc283845a, 32'hc2c0b2ac, 32'hc2546c31, 32'h414c20a5, 32'hc2b09a1a, 32'h41d43a1c, 32'hc28646f8, 32'h42a43787};
test_output[29920:29927] = '{32'h0, 32'h0, 32'h0, 32'h414c20a5, 32'h0, 32'h41d43a1c, 32'h0, 32'h42a43787};
test_input[29928:29935] = '{32'h42a2e0c1, 32'h418b4860, 32'hc151bc66, 32'h428fc6b4, 32'hc2832620, 32'h427bfb0d, 32'hc19d0e4b, 32'hc259a1eb};
test_output[29928:29935] = '{32'h42a2e0c1, 32'h418b4860, 32'h0, 32'h428fc6b4, 32'h0, 32'h427bfb0d, 32'h0, 32'h0};
test_input[29936:29943] = '{32'h41f88754, 32'hc288e172, 32'hc1719ee6, 32'h422e63fe, 32'h428d529f, 32'hc02f393a, 32'hc2bb6b8d, 32'hc2277d7e};
test_output[29936:29943] = '{32'h41f88754, 32'h0, 32'h0, 32'h422e63fe, 32'h428d529f, 32'h0, 32'h0, 32'h0};
test_input[29944:29951] = '{32'hc244a093, 32'h41832cbd, 32'hc2277b1f, 32'hc246f1a2, 32'hc2bb0566, 32'hc19af45c, 32'hc1d94eaf, 32'h4288a4f1};
test_output[29944:29951] = '{32'h0, 32'h41832cbd, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4288a4f1};
test_input[29952:29959] = '{32'hc14d86e3, 32'h429cf6c5, 32'hc21c9da6, 32'h41d3b433, 32'hc29397e7, 32'h429455af, 32'h426fe35b, 32'h428e3ea3};
test_output[29952:29959] = '{32'h0, 32'h429cf6c5, 32'h0, 32'h41d3b433, 32'h0, 32'h429455af, 32'h426fe35b, 32'h428e3ea3};
test_input[29960:29967] = '{32'hc0a366dc, 32'h40f473cd, 32'h42bfe803, 32'hc1e86056, 32'h423060e5, 32'h419fc76a, 32'hc270e1bd, 32'hc14d6b07};
test_output[29960:29967] = '{32'h0, 32'h40f473cd, 32'h42bfe803, 32'h0, 32'h423060e5, 32'h419fc76a, 32'h0, 32'h0};
test_input[29968:29975] = '{32'hc252ae97, 32'hc1c7fa68, 32'h425bc7d0, 32'hc15458cd, 32'h41c5f4bb, 32'hc237a098, 32'hc04f8959, 32'h42889a4f};
test_output[29968:29975] = '{32'h0, 32'h0, 32'h425bc7d0, 32'h0, 32'h41c5f4bb, 32'h0, 32'h0, 32'h42889a4f};
test_input[29976:29983] = '{32'hc210f605, 32'hc2bce746, 32'hc1c19465, 32'h415c5af2, 32'h42a88d2a, 32'hc2a9ca09, 32'h426f59e8, 32'h42337641};
test_output[29976:29983] = '{32'h0, 32'h0, 32'h0, 32'h415c5af2, 32'h42a88d2a, 32'h0, 32'h426f59e8, 32'h42337641};
test_input[29984:29991] = '{32'hc2721887, 32'hc0f82667, 32'hc2758472, 32'hc1b40af6, 32'h4234ddcf, 32'hc0e28d5f, 32'hc18ed1e7, 32'hc2666ab4};
test_output[29984:29991] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4234ddcf, 32'h0, 32'h0, 32'h0};
test_input[29992:29999] = '{32'hc1e43725, 32'hc220aecf, 32'h41e67039, 32'hc2353237, 32'h4178ca60, 32'hc28e0b39, 32'h40e8de1a, 32'h4238cd09};
test_output[29992:29999] = '{32'h0, 32'h0, 32'h41e67039, 32'h0, 32'h4178ca60, 32'h0, 32'h40e8de1a, 32'h4238cd09};
test_input[30000:30007] = '{32'hc26eb056, 32'h424ae0b5, 32'h4127a311, 32'hc252ca48, 32'hc24d9479, 32'h42068167, 32'h41d74dcd, 32'hc23cb717};
test_output[30000:30007] = '{32'h0, 32'h424ae0b5, 32'h4127a311, 32'h0, 32'h0, 32'h42068167, 32'h41d74dcd, 32'h0};
test_input[30008:30015] = '{32'h42970861, 32'h4117b914, 32'h42026629, 32'h4289efa8, 32'hc2739767, 32'hc12fae32, 32'hc259467a, 32'hc165fd60};
test_output[30008:30015] = '{32'h42970861, 32'h4117b914, 32'h42026629, 32'h4289efa8, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30016:30023] = '{32'h421518bc, 32'h41822ed2, 32'hc20a6b7c, 32'hc1c6c8d3, 32'hc21acfc7, 32'h41867570, 32'h4255fcf9, 32'h42aac608};
test_output[30016:30023] = '{32'h421518bc, 32'h41822ed2, 32'h0, 32'h0, 32'h0, 32'h41867570, 32'h4255fcf9, 32'h42aac608};
test_input[30024:30031] = '{32'h41ecb31f, 32'hc18b039b, 32'hc19a2118, 32'hc13eeec9, 32'h428edb87, 32'h42452713, 32'h428b017d, 32'h42699e63};
test_output[30024:30031] = '{32'h41ecb31f, 32'h0, 32'h0, 32'h0, 32'h428edb87, 32'h42452713, 32'h428b017d, 32'h42699e63};
test_input[30032:30039] = '{32'h41e8e21e, 32'h42a3e7ca, 32'h41a87741, 32'h40a82d21, 32'h41d8ea00, 32'hc21bf83d, 32'hc25e0655, 32'h414e4bea};
test_output[30032:30039] = '{32'h41e8e21e, 32'h42a3e7ca, 32'h41a87741, 32'h40a82d21, 32'h41d8ea00, 32'h0, 32'h0, 32'h414e4bea};
test_input[30040:30047] = '{32'hc28a80a2, 32'h40decb16, 32'hc269088f, 32'hc1edb1c9, 32'hc266c0f1, 32'h4103cf3c, 32'h414ce413, 32'h42bed3c7};
test_output[30040:30047] = '{32'h0, 32'h40decb16, 32'h0, 32'h0, 32'h0, 32'h4103cf3c, 32'h414ce413, 32'h42bed3c7};
test_input[30048:30055] = '{32'hc0e6a128, 32'hc2a9ddd0, 32'h42526d7c, 32'h422576a4, 32'hc285a5a6, 32'h426f08cd, 32'h42b27a0e, 32'h427bbb8b};
test_output[30048:30055] = '{32'h0, 32'h0, 32'h42526d7c, 32'h422576a4, 32'h0, 32'h426f08cd, 32'h42b27a0e, 32'h427bbb8b};
test_input[30056:30063] = '{32'h42656aa5, 32'hc2688e6c, 32'hc1f2ca79, 32'h421acaa5, 32'hc27caf5c, 32'hc233fdbe, 32'hbf40e564, 32'h4218f0d4};
test_output[30056:30063] = '{32'h42656aa5, 32'h0, 32'h0, 32'h421acaa5, 32'h0, 32'h0, 32'h0, 32'h4218f0d4};
test_input[30064:30071] = '{32'hc1c32327, 32'h428b2f51, 32'h42901d0c, 32'h429af515, 32'hc2870b2f, 32'hc2ae0606, 32'hc299d6fb, 32'hc29da35a};
test_output[30064:30071] = '{32'h0, 32'h428b2f51, 32'h42901d0c, 32'h429af515, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30072:30079] = '{32'hbf30ac84, 32'h4298e49c, 32'h42283419, 32'h4286e7df, 32'hc20d7745, 32'hbfd22a24, 32'hbf03c956, 32'hc1a533f4};
test_output[30072:30079] = '{32'h0, 32'h4298e49c, 32'h42283419, 32'h4286e7df, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30080:30087] = '{32'hc2891d5d, 32'hc11d9c77, 32'hc2b6c1b8, 32'h4269d4bb, 32'h42b35467, 32'hc27820cb, 32'hc1de74d6, 32'h4126f528};
test_output[30080:30087] = '{32'h0, 32'h0, 32'h0, 32'h4269d4bb, 32'h42b35467, 32'h0, 32'h0, 32'h4126f528};
test_input[30088:30095] = '{32'hc2b6b507, 32'h424e27ef, 32'hc2a32e67, 32'h412d3fc3, 32'hc2c59307, 32'hc2b4ea57, 32'hc28dd7c9, 32'h425d2120};
test_output[30088:30095] = '{32'h0, 32'h424e27ef, 32'h0, 32'h412d3fc3, 32'h0, 32'h0, 32'h0, 32'h425d2120};
test_input[30096:30103] = '{32'hc23a57b1, 32'h426eff58, 32'hc24e38c7, 32'hc1879a9c, 32'hc251fdd2, 32'hc2a651d7, 32'hc1c1e3a8, 32'h4288bee7};
test_output[30096:30103] = '{32'h0, 32'h426eff58, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4288bee7};
test_input[30104:30111] = '{32'h41b456f5, 32'hc260830b, 32'hc2797297, 32'h4295d49a, 32'hc26c926e, 32'hc2236386, 32'h4233bdac, 32'hc232067c};
test_output[30104:30111] = '{32'h41b456f5, 32'h0, 32'h0, 32'h4295d49a, 32'h0, 32'h0, 32'h4233bdac, 32'h0};
test_input[30112:30119] = '{32'hc2c3542f, 32'h4273e235, 32'hc21e30a4, 32'hc1ed670a, 32'h42a21879, 32'h429831b6, 32'hc242403b, 32'h41f667a0};
test_output[30112:30119] = '{32'h0, 32'h4273e235, 32'h0, 32'h0, 32'h42a21879, 32'h429831b6, 32'h0, 32'h41f667a0};
test_input[30120:30127] = '{32'h414e2ba1, 32'h42ab0442, 32'h4228689d, 32'hc01619d9, 32'h42521b08, 32'hc289d88b, 32'hc2b2cd4b, 32'hc201ea16};
test_output[30120:30127] = '{32'h414e2ba1, 32'h42ab0442, 32'h4228689d, 32'h0, 32'h42521b08, 32'h0, 32'h0, 32'h0};
test_input[30128:30135] = '{32'hc1cf7efd, 32'h4195ef13, 32'hc2bf9f6e, 32'h41e8350e, 32'h41045c93, 32'hc251cddb, 32'hc283f42a, 32'h41ee2d06};
test_output[30128:30135] = '{32'h0, 32'h4195ef13, 32'h0, 32'h41e8350e, 32'h41045c93, 32'h0, 32'h0, 32'h41ee2d06};
test_input[30136:30143] = '{32'hc2b70f77, 32'h423dfe9c, 32'h426750cb, 32'hc29f56ff, 32'h420e6648, 32'h42648ed0, 32'h42a50a3f, 32'h42ab38c4};
test_output[30136:30143] = '{32'h0, 32'h423dfe9c, 32'h426750cb, 32'h0, 32'h420e6648, 32'h42648ed0, 32'h42a50a3f, 32'h42ab38c4};
test_input[30144:30151] = '{32'h4278fdde, 32'h42c54d25, 32'h4150f46f, 32'hc288e168, 32'h42509be9, 32'hc21f5b49, 32'h4293ffc7, 32'hc2b83fc4};
test_output[30144:30151] = '{32'h4278fdde, 32'h42c54d25, 32'h4150f46f, 32'h0, 32'h42509be9, 32'h0, 32'h4293ffc7, 32'h0};
test_input[30152:30159] = '{32'hc2386e95, 32'h419b85c9, 32'h429039f9, 32'hc28fb4fd, 32'h42819e12, 32'h4249ccc9, 32'h4262daf1, 32'h428a971f};
test_output[30152:30159] = '{32'h0, 32'h419b85c9, 32'h429039f9, 32'h0, 32'h42819e12, 32'h4249ccc9, 32'h4262daf1, 32'h428a971f};
test_input[30160:30167] = '{32'hc0905557, 32'h429d6d88, 32'h4294d016, 32'hbe0f4f88, 32'hc249ea07, 32'h41ace55d, 32'h429701b1, 32'h427d85b9};
test_output[30160:30167] = '{32'h0, 32'h429d6d88, 32'h4294d016, 32'h0, 32'h0, 32'h41ace55d, 32'h429701b1, 32'h427d85b9};
test_input[30168:30175] = '{32'h41d4f01d, 32'h42aeb464, 32'hc1829b7d, 32'h41d3fd9d, 32'hc1a9c934, 32'hc169a030, 32'hc2a51c1f, 32'h42605886};
test_output[30168:30175] = '{32'h41d4f01d, 32'h42aeb464, 32'h0, 32'h41d3fd9d, 32'h0, 32'h0, 32'h0, 32'h42605886};
test_input[30176:30183] = '{32'h40fbd4dc, 32'h421c8838, 32'h4224f9fc, 32'hc20da00e, 32'h42480b7a, 32'h426f90cc, 32'h421bc8db, 32'h4200d637};
test_output[30176:30183] = '{32'h40fbd4dc, 32'h421c8838, 32'h4224f9fc, 32'h0, 32'h42480b7a, 32'h426f90cc, 32'h421bc8db, 32'h4200d637};
test_input[30184:30191] = '{32'h42a2e265, 32'h423de4cf, 32'hc2b609bb, 32'hc29f40d7, 32'hc2b230b1, 32'hc224160e, 32'hc11f11ed, 32'h409b4a04};
test_output[30184:30191] = '{32'h42a2e265, 32'h423de4cf, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h409b4a04};
test_input[30192:30199] = '{32'hc295cd4e, 32'hc24b54d6, 32'hc2210cc5, 32'h42ab6856, 32'hc29a6e41, 32'h4216d6a0, 32'hc21bdab7, 32'h42699bb1};
test_output[30192:30199] = '{32'h0, 32'h0, 32'h0, 32'h42ab6856, 32'h0, 32'h4216d6a0, 32'h0, 32'h42699bb1};
test_input[30200:30207] = '{32'h42c04f64, 32'h42acb403, 32'hc11034b6, 32'hc2053d5c, 32'hc2511e8b, 32'h42395ca2, 32'hc24bf548, 32'hc2a3aad1};
test_output[30200:30207] = '{32'h42c04f64, 32'h42acb403, 32'h0, 32'h0, 32'h0, 32'h42395ca2, 32'h0, 32'h0};
test_input[30208:30215] = '{32'h41bae092, 32'hbfd525c0, 32'h42447a60, 32'h42abfe01, 32'h42bc2aa8, 32'h41cd5abf, 32'h4281c2e2, 32'h42824047};
test_output[30208:30215] = '{32'h41bae092, 32'h0, 32'h42447a60, 32'h42abfe01, 32'h42bc2aa8, 32'h41cd5abf, 32'h4281c2e2, 32'h42824047};
test_input[30216:30223] = '{32'hc2a24e85, 32'h41909fb6, 32'h42aeb62a, 32'h421d8840, 32'hc06d9407, 32'h41f20265, 32'hc1f78ae7, 32'hc2a20c98};
test_output[30216:30223] = '{32'h0, 32'h41909fb6, 32'h42aeb62a, 32'h421d8840, 32'h0, 32'h41f20265, 32'h0, 32'h0};
test_input[30224:30231] = '{32'hc19c3125, 32'hc2b1422b, 32'hc2242b19, 32'h429c2d9f, 32'h4295f001, 32'h4238250a, 32'hc22fe338, 32'hc1b98e83};
test_output[30224:30231] = '{32'h0, 32'h0, 32'h0, 32'h429c2d9f, 32'h4295f001, 32'h4238250a, 32'h0, 32'h0};
test_input[30232:30239] = '{32'hc2b58963, 32'hc1d49ffb, 32'hc1b4ebb8, 32'hc1502e46, 32'h4222b574, 32'hc1d5694c, 32'hc2872298, 32'h42952a82};
test_output[30232:30239] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4222b574, 32'h0, 32'h0, 32'h42952a82};
test_input[30240:30247] = '{32'h424d5739, 32'h42a28bad, 32'hc200332f, 32'h420c866c, 32'hc2a820b9, 32'h428c6a43, 32'hc125f3cd, 32'hc28f179f};
test_output[30240:30247] = '{32'h424d5739, 32'h42a28bad, 32'h0, 32'h420c866c, 32'h0, 32'h428c6a43, 32'h0, 32'h0};
test_input[30248:30255] = '{32'h42c113ef, 32'h426004b4, 32'h416fa194, 32'hc1b182d3, 32'h40bb232e, 32'hc1b141b1, 32'hc1cc35e1, 32'hc2903c20};
test_output[30248:30255] = '{32'h42c113ef, 32'h426004b4, 32'h416fa194, 32'h0, 32'h40bb232e, 32'h0, 32'h0, 32'h0};
test_input[30256:30263] = '{32'h424bb3b0, 32'hc1bad2cb, 32'hc2068912, 32'hc0dedb8b, 32'hc20d2173, 32'h40a4234b, 32'h41a875a0, 32'h4290e095};
test_output[30256:30263] = '{32'h424bb3b0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40a4234b, 32'h41a875a0, 32'h4290e095};
test_input[30264:30271] = '{32'h414ba819, 32'h426e9ece, 32'h41f07151, 32'hc26c599c, 32'hc2b19ea4, 32'hc242814c, 32'h420c9277, 32'h4104489e};
test_output[30264:30271] = '{32'h414ba819, 32'h426e9ece, 32'h41f07151, 32'h0, 32'h0, 32'h0, 32'h420c9277, 32'h4104489e};
test_input[30272:30279] = '{32'h41f4512e, 32'hc17114b5, 32'hc21e5f4e, 32'h426573a6, 32'hc1b80e42, 32'h4204c3f3, 32'hc282e045, 32'h429f2ae7};
test_output[30272:30279] = '{32'h41f4512e, 32'h0, 32'h0, 32'h426573a6, 32'h0, 32'h4204c3f3, 32'h0, 32'h429f2ae7};
test_input[30280:30287] = '{32'h42767f79, 32'hc2c2730a, 32'h41e7c5a2, 32'hc2bd66bf, 32'h42aeff31, 32'hc1d75995, 32'hc2c20ea6, 32'hc11cbdfd};
test_output[30280:30287] = '{32'h42767f79, 32'h0, 32'h41e7c5a2, 32'h0, 32'h42aeff31, 32'h0, 32'h0, 32'h0};
test_input[30288:30295] = '{32'hc230e658, 32'hc1aeb936, 32'h4200e8b1, 32'h4293b623, 32'hc1e7f6ee, 32'hc187062f, 32'hc098e286, 32'h42025f36};
test_output[30288:30295] = '{32'h0, 32'h0, 32'h4200e8b1, 32'h4293b623, 32'h0, 32'h0, 32'h0, 32'h42025f36};
test_input[30296:30303] = '{32'hc0893441, 32'hc29d3dfe, 32'hc2a451c6, 32'h4222b569, 32'h41b21a99, 32'h42ad2aa2, 32'hc28d1155, 32'h42ae3981};
test_output[30296:30303] = '{32'h0, 32'h0, 32'h0, 32'h4222b569, 32'h41b21a99, 32'h42ad2aa2, 32'h0, 32'h42ae3981};
test_input[30304:30311] = '{32'hc28be409, 32'hc1ce2e27, 32'h42797b42, 32'hc2023bc1, 32'h426f9738, 32'h4287212d, 32'hc205c58c, 32'h42b8f5c8};
test_output[30304:30311] = '{32'h0, 32'h0, 32'h42797b42, 32'h0, 32'h426f9738, 32'h4287212d, 32'h0, 32'h42b8f5c8};
test_input[30312:30319] = '{32'h42a4ad8f, 32'h41f1b209, 32'h4290ca34, 32'hc201325f, 32'hc0d1925c, 32'h423e951d, 32'h3fce2768, 32'h42247c79};
test_output[30312:30319] = '{32'h42a4ad8f, 32'h41f1b209, 32'h4290ca34, 32'h0, 32'h0, 32'h423e951d, 32'h3fce2768, 32'h42247c79};
test_input[30320:30327] = '{32'h42278733, 32'h4280f963, 32'hc121df7c, 32'hc262386f, 32'h42b70053, 32'hc21eb85c, 32'h41edb44c, 32'hc263ff41};
test_output[30320:30327] = '{32'h42278733, 32'h4280f963, 32'h0, 32'h0, 32'h42b70053, 32'h0, 32'h41edb44c, 32'h0};
test_input[30328:30335] = '{32'h41c5e209, 32'hc28d3d84, 32'hc22f40b8, 32'hc26d860a, 32'hc2ab99da, 32'hc287a8e1, 32'hc2be4eb8, 32'hc1ff28fd};
test_output[30328:30335] = '{32'h41c5e209, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30336:30343] = '{32'hbff5131b, 32'h427bd46a, 32'hc25bbd07, 32'h42a426ad, 32'h42adb399, 32'h42b1e9e3, 32'h412f3a5f, 32'h41aa1c5b};
test_output[30336:30343] = '{32'h0, 32'h427bd46a, 32'h0, 32'h42a426ad, 32'h42adb399, 32'h42b1e9e3, 32'h412f3a5f, 32'h41aa1c5b};
test_input[30344:30351] = '{32'h42b9e995, 32'hc22632c2, 32'hc22f5fec, 32'h4238d7ca, 32'hc2a81669, 32'hc293100d, 32'hc2778658, 32'h40faea51};
test_output[30344:30351] = '{32'h42b9e995, 32'h0, 32'h0, 32'h4238d7ca, 32'h0, 32'h0, 32'h0, 32'h40faea51};
test_input[30352:30359] = '{32'h4258a8a4, 32'h41e5ec38, 32'hc23e6bc7, 32'h42070fc1, 32'hc2c753bb, 32'h426bb7b3, 32'hc295dcdf, 32'h41b0596c};
test_output[30352:30359] = '{32'h4258a8a4, 32'h41e5ec38, 32'h0, 32'h42070fc1, 32'h0, 32'h426bb7b3, 32'h0, 32'h41b0596c};
test_input[30360:30367] = '{32'hc274a56b, 32'hc0e28e8d, 32'hc29c08a9, 32'hc2a0aecf, 32'h426068eb, 32'h414d322e, 32'h4120b20d, 32'hc20a508b};
test_output[30360:30367] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h426068eb, 32'h414d322e, 32'h4120b20d, 32'h0};
test_input[30368:30375] = '{32'hc1c1eb20, 32'hc20f4e06, 32'hc2770d77, 32'h42940b3f, 32'h42708609, 32'hc0e1a89f, 32'h42890cb4, 32'h4125f036};
test_output[30368:30375] = '{32'h0, 32'h0, 32'h0, 32'h42940b3f, 32'h42708609, 32'h0, 32'h42890cb4, 32'h4125f036};
test_input[30376:30383] = '{32'h42479bf7, 32'h40cda9c5, 32'hbee1737e, 32'h4252b098, 32'hc25cc7f9, 32'hc28156fc, 32'h4252ccde, 32'h4269e1c9};
test_output[30376:30383] = '{32'h42479bf7, 32'h40cda9c5, 32'h0, 32'h4252b098, 32'h0, 32'h0, 32'h4252ccde, 32'h4269e1c9};
test_input[30384:30391] = '{32'h42274462, 32'h42502499, 32'h42af62bb, 32'hc2116980, 32'h40a8bdd4, 32'hc23a3cf9, 32'h4293a798, 32'h42c44b1d};
test_output[30384:30391] = '{32'h42274462, 32'h42502499, 32'h42af62bb, 32'h0, 32'h40a8bdd4, 32'h0, 32'h4293a798, 32'h42c44b1d};
test_input[30392:30399] = '{32'hc2aa39fb, 32'h42914982, 32'hc25e5a60, 32'h428e9615, 32'hc29e9e72, 32'hc271874e, 32'hc2b6f1c4, 32'hc268e1bb};
test_output[30392:30399] = '{32'h0, 32'h42914982, 32'h0, 32'h428e9615, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30400:30407] = '{32'h42161c76, 32'hc2a61930, 32'h413c2ec8, 32'h4291da8a, 32'h410a796e, 32'hc29eb66a, 32'hc2126544, 32'h41a50adc};
test_output[30400:30407] = '{32'h42161c76, 32'h0, 32'h413c2ec8, 32'h4291da8a, 32'h410a796e, 32'h0, 32'h0, 32'h41a50adc};
test_input[30408:30415] = '{32'h426927fe, 32'hc25897ec, 32'h4266ff4e, 32'hc2b27a90, 32'h4023f7bb, 32'h428b9833, 32'h41bc047e, 32'hc2968aef};
test_output[30408:30415] = '{32'h426927fe, 32'h0, 32'h4266ff4e, 32'h0, 32'h4023f7bb, 32'h428b9833, 32'h41bc047e, 32'h0};
test_input[30416:30423] = '{32'hc053d51c, 32'hc291e98d, 32'hc26c7f33, 32'hc2b3ec97, 32'h42c36e43, 32'hc0b0355b, 32'h42a2da61, 32'h429f667e};
test_output[30416:30423] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42c36e43, 32'h0, 32'h42a2da61, 32'h429f667e};
test_input[30424:30431] = '{32'hc282ddb2, 32'hc2562d6d, 32'h428d0ccb, 32'h429624da, 32'h42860a06, 32'hc245678a, 32'hc2c48e78, 32'hc2785012};
test_output[30424:30431] = '{32'h0, 32'h0, 32'h428d0ccb, 32'h429624da, 32'h42860a06, 32'h0, 32'h0, 32'h0};
test_input[30432:30439] = '{32'h42b48a35, 32'h4276becb, 32'hc260673d, 32'hc29f1b07, 32'hc1227b65, 32'hc2a9f03f, 32'hc0c87085, 32'hbf0d96ad};
test_output[30432:30439] = '{32'h42b48a35, 32'h4276becb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30440:30447] = '{32'hc08eb846, 32'hc0ce8dcb, 32'hc1d70e52, 32'hc2c1d3df, 32'hc28baa31, 32'hc1ff10b9, 32'hc27c78d7, 32'h422fd5b7};
test_output[30440:30447] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422fd5b7};
test_input[30448:30455] = '{32'hc1358312, 32'hc1f79f94, 32'hc256d075, 32'h41a99f89, 32'hc25c077f, 32'h41e3e60b, 32'h4265ec54, 32'hc1940c28};
test_output[30448:30455] = '{32'h0, 32'h0, 32'h0, 32'h41a99f89, 32'h0, 32'h41e3e60b, 32'h4265ec54, 32'h0};
test_input[30456:30463] = '{32'h42c56be5, 32'hc2934665, 32'hc28acaeb, 32'h41eabba4, 32'hc2c2d8cb, 32'h41513e26, 32'hc2bc926c, 32'hc1cd2f55};
test_output[30456:30463] = '{32'h42c56be5, 32'h0, 32'h0, 32'h41eabba4, 32'h0, 32'h41513e26, 32'h0, 32'h0};
test_input[30464:30471] = '{32'hc1324065, 32'h3ee48fc0, 32'hc1a77275, 32'hc209672f, 32'h42b5c520, 32'hc21c33fb, 32'hc01e0810, 32'h422eea4d};
test_output[30464:30471] = '{32'h0, 32'h3ee48fc0, 32'h0, 32'h0, 32'h42b5c520, 32'h0, 32'h0, 32'h422eea4d};
test_input[30472:30479] = '{32'hc22f883b, 32'h41b4f76c, 32'hc1cb762e, 32'h42b131ab, 32'h42914329, 32'hc2a6f112, 32'hc20890cc, 32'h42b2608e};
test_output[30472:30479] = '{32'h0, 32'h41b4f76c, 32'h0, 32'h42b131ab, 32'h42914329, 32'h0, 32'h0, 32'h42b2608e};
test_input[30480:30487] = '{32'h423f3d28, 32'h420b47f7, 32'h4229d38e, 32'hc2a7896e, 32'hc2b1058b, 32'hc11e2289, 32'hc19172b1, 32'hc158d565};
test_output[30480:30487] = '{32'h423f3d28, 32'h420b47f7, 32'h4229d38e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30488:30495] = '{32'h415984f2, 32'h423ecfa8, 32'h4237bdc7, 32'hc29e9761, 32'hc0e872d5, 32'hc24fe0cc, 32'h42ac9d66, 32'hc2b3ee14};
test_output[30488:30495] = '{32'h415984f2, 32'h423ecfa8, 32'h4237bdc7, 32'h0, 32'h0, 32'h0, 32'h42ac9d66, 32'h0};
test_input[30496:30503] = '{32'hc23c9b52, 32'hc214b241, 32'hc19b6c29, 32'h42490227, 32'hc0587562, 32'hc1097fbd, 32'hc10a3269, 32'hc2c41b57};
test_output[30496:30503] = '{32'h0, 32'h0, 32'h0, 32'h42490227, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30504:30511] = '{32'hc2070187, 32'hc22e3ad5, 32'hc2064b42, 32'h42225b4d, 32'hc26a8bca, 32'hc1b41e97, 32'h421bc654, 32'h41c75124};
test_output[30504:30511] = '{32'h0, 32'h0, 32'h0, 32'h42225b4d, 32'h0, 32'h0, 32'h421bc654, 32'h41c75124};
test_input[30512:30519] = '{32'h42a4af97, 32'hc23f8f9d, 32'h429c858c, 32'hc234bfce, 32'hc26a17a6, 32'hc0c89f5f, 32'h42684337, 32'h42b20cc6};
test_output[30512:30519] = '{32'h42a4af97, 32'h0, 32'h429c858c, 32'h0, 32'h0, 32'h0, 32'h42684337, 32'h42b20cc6};
test_input[30520:30527] = '{32'hc2a11f95, 32'hc2c45e98, 32'h41a82e9c, 32'hc2275841, 32'hc26ab59e, 32'h42c56c0e, 32'hc18bdc57, 32'hc11b7d34};
test_output[30520:30527] = '{32'h0, 32'h0, 32'h41a82e9c, 32'h0, 32'h0, 32'h42c56c0e, 32'h0, 32'h0};
test_input[30528:30535] = '{32'h42a4a07d, 32'h42887e94, 32'h4088a1a9, 32'hc2b785f6, 32'hc1c82f49, 32'hc22abfeb, 32'h42823fa0, 32'h4079a052};
test_output[30528:30535] = '{32'h42a4a07d, 32'h42887e94, 32'h4088a1a9, 32'h0, 32'h0, 32'h0, 32'h42823fa0, 32'h4079a052};
test_input[30536:30543] = '{32'hc2b09617, 32'hc22c167a, 32'hc066c89e, 32'hc097f4a2, 32'hc23c5beb, 32'hc2c5eab3, 32'h42764318, 32'h4255af4c};
test_output[30536:30543] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42764318, 32'h4255af4c};
test_input[30544:30551] = '{32'hc283bb9e, 32'h42b6cd53, 32'h4277dd6e, 32'h4281c983, 32'hc24c9344, 32'hc2999e01, 32'h42797e4d, 32'hbf31009e};
test_output[30544:30551] = '{32'h0, 32'h42b6cd53, 32'h4277dd6e, 32'h4281c983, 32'h0, 32'h0, 32'h42797e4d, 32'h0};
test_input[30552:30559] = '{32'hc2aadd76, 32'hc213742c, 32'h426c46f8, 32'hc284e6a0, 32'hc20818e0, 32'h418bd070, 32'h42876f8c, 32'hc0d9043d};
test_output[30552:30559] = '{32'h0, 32'h0, 32'h426c46f8, 32'h0, 32'h0, 32'h418bd070, 32'h42876f8c, 32'h0};
test_input[30560:30567] = '{32'h40d3003e, 32'h41812053, 32'h42336880, 32'hc2c5445b, 32'hc17beb68, 32'h424dab43, 32'h42a04689, 32'hc2c165d5};
test_output[30560:30567] = '{32'h40d3003e, 32'h41812053, 32'h42336880, 32'h0, 32'h0, 32'h424dab43, 32'h42a04689, 32'h0};
test_input[30568:30575] = '{32'h429d9732, 32'h420d6e41, 32'hc27c173d, 32'h42003d77, 32'hc0edc9db, 32'h41fcbd66, 32'hc0b9f9cb, 32'h429a3bc1};
test_output[30568:30575] = '{32'h429d9732, 32'h420d6e41, 32'h0, 32'h42003d77, 32'h0, 32'h41fcbd66, 32'h0, 32'h429a3bc1};
test_input[30576:30583] = '{32'hc2386459, 32'hc17ab7c1, 32'h42bbb153, 32'hc2703b0c, 32'hc0d61487, 32'h42227f23, 32'h4216eeb3, 32'hbfa979d4};
test_output[30576:30583] = '{32'h0, 32'h0, 32'h42bbb153, 32'h0, 32'h0, 32'h42227f23, 32'h4216eeb3, 32'h0};
test_input[30584:30591] = '{32'h4241ed2b, 32'hc248d8d1, 32'h4134d28a, 32'hc27c7f48, 32'h42081985, 32'h428a99a0, 32'hc2b7191d, 32'hc1a9c411};
test_output[30584:30591] = '{32'h4241ed2b, 32'h0, 32'h4134d28a, 32'h0, 32'h42081985, 32'h428a99a0, 32'h0, 32'h0};
test_input[30592:30599] = '{32'hc2aa2214, 32'h429c4530, 32'h42bc6d74, 32'hc1ef9a68, 32'h422a5442, 32'hc2bfb9d3, 32'h42466fc9, 32'hc2790a0b};
test_output[30592:30599] = '{32'h0, 32'h429c4530, 32'h42bc6d74, 32'h0, 32'h422a5442, 32'h0, 32'h42466fc9, 32'h0};
test_input[30600:30607] = '{32'hc2951581, 32'h42967abf, 32'hc228f308, 32'hc28c7809, 32'h4193015b, 32'h428e6b94, 32'h42b8dfeb, 32'hc187a38b};
test_output[30600:30607] = '{32'h0, 32'h42967abf, 32'h0, 32'h0, 32'h4193015b, 32'h428e6b94, 32'h42b8dfeb, 32'h0};
test_input[30608:30615] = '{32'h41dd7e6f, 32'h42588fdb, 32'hc1af01ae, 32'h42a9c660, 32'h42050a30, 32'hc2351eda, 32'h429b80d5, 32'h42a51ab9};
test_output[30608:30615] = '{32'h41dd7e6f, 32'h42588fdb, 32'h0, 32'h42a9c660, 32'h42050a30, 32'h0, 32'h429b80d5, 32'h42a51ab9};
test_input[30616:30623] = '{32'hc243284d, 32'h41f2c65e, 32'h41e19ba9, 32'h41481193, 32'hc251b5be, 32'hc249502e, 32'h418f1271, 32'h42a6a6d4};
test_output[30616:30623] = '{32'h0, 32'h41f2c65e, 32'h41e19ba9, 32'h41481193, 32'h0, 32'h0, 32'h418f1271, 32'h42a6a6d4};
test_input[30624:30631] = '{32'hc2bc5ee9, 32'hc0456e76, 32'hc1c4b3ef, 32'h42c0d2e2, 32'h4289fffe, 32'hc1e7423a, 32'hc2bcd3ab, 32'hc2379e09};
test_output[30624:30631] = '{32'h0, 32'h0, 32'h0, 32'h42c0d2e2, 32'h4289fffe, 32'h0, 32'h0, 32'h0};
test_input[30632:30639] = '{32'h428fc4e2, 32'hc200b38d, 32'hc2c258f6, 32'h419ec44e, 32'h425e77de, 32'hc290b46b, 32'h42ae335f, 32'h4245bf16};
test_output[30632:30639] = '{32'h428fc4e2, 32'h0, 32'h0, 32'h419ec44e, 32'h425e77de, 32'h0, 32'h42ae335f, 32'h4245bf16};
test_input[30640:30647] = '{32'h423a8f37, 32'hc17be802, 32'hc2a499f5, 32'hc1d68611, 32'hc1b64f03, 32'h4293274f, 32'hc1afe1fc, 32'hc1a5b4db};
test_output[30640:30647] = '{32'h423a8f37, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4293274f, 32'h0, 32'h0};
test_input[30648:30655] = '{32'h42b8af1f, 32'hc19efb41, 32'hc2927f9c, 32'h405cc882, 32'h42937fde, 32'h40133c15, 32'hc22aa848, 32'hc2858614};
test_output[30648:30655] = '{32'h42b8af1f, 32'h0, 32'h0, 32'h405cc882, 32'h42937fde, 32'h40133c15, 32'h0, 32'h0};
test_input[30656:30663] = '{32'h419b6b9e, 32'hc2887e42, 32'hc239d7cf, 32'h429fb7f8, 32'h42494716, 32'hc2beb6e2, 32'hc1ed66fb, 32'h4254d3e7};
test_output[30656:30663] = '{32'h419b6b9e, 32'h0, 32'h0, 32'h429fb7f8, 32'h42494716, 32'h0, 32'h0, 32'h4254d3e7};
test_input[30664:30671] = '{32'hc2c47fcb, 32'hbfc1b3a4, 32'hc2bf196f, 32'h42876d38, 32'h425fac5a, 32'hc2c4465a, 32'hc1c33b5d, 32'h4200c56a};
test_output[30664:30671] = '{32'h0, 32'h0, 32'h0, 32'h42876d38, 32'h425fac5a, 32'h0, 32'h0, 32'h4200c56a};
test_input[30672:30679] = '{32'h41a2acfa, 32'hc1f0d129, 32'hc1fea854, 32'h4295588e, 32'h423a5da2, 32'hc225a183, 32'hc28f95be, 32'h4235db45};
test_output[30672:30679] = '{32'h41a2acfa, 32'h0, 32'h0, 32'h4295588e, 32'h423a5da2, 32'h0, 32'h0, 32'h4235db45};
test_input[30680:30687] = '{32'hc237030c, 32'hc1954de4, 32'h4222340e, 32'hc2a80c11, 32'h427ca255, 32'hc1961982, 32'hc1ca0229, 32'hc153eed8};
test_output[30680:30687] = '{32'h0, 32'h0, 32'h4222340e, 32'h0, 32'h427ca255, 32'h0, 32'h0, 32'h0};
test_input[30688:30695] = '{32'hc0cb5333, 32'hc25ab382, 32'hc27733cf, 32'h42c317d7, 32'hbf8594e7, 32'hc29c942e, 32'h42a1bc3e, 32'h427ba2f4};
test_output[30688:30695] = '{32'h0, 32'h0, 32'h0, 32'h42c317d7, 32'h0, 32'h0, 32'h42a1bc3e, 32'h427ba2f4};
test_input[30696:30703] = '{32'h42208feb, 32'hc18975bf, 32'hc2b66144, 32'hc1b31ac1, 32'hc2b2b357, 32'hc1959cac, 32'hc201b0a7, 32'h428a2d36};
test_output[30696:30703] = '{32'h42208feb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428a2d36};
test_input[30704:30711] = '{32'hc29b36f7, 32'h4291dc92, 32'h41e86905, 32'hc2330441, 32'h42816729, 32'hc28f057f, 32'h41aa2d67, 32'h422cb748};
test_output[30704:30711] = '{32'h0, 32'h4291dc92, 32'h41e86905, 32'h0, 32'h42816729, 32'h0, 32'h41aa2d67, 32'h422cb748};
test_input[30712:30719] = '{32'h42a7ccb2, 32'hc2970c05, 32'h40b40803, 32'h41e1d867, 32'hc0345351, 32'h42b73557, 32'h4103423c, 32'h4203ba64};
test_output[30712:30719] = '{32'h42a7ccb2, 32'h0, 32'h40b40803, 32'h41e1d867, 32'h0, 32'h42b73557, 32'h4103423c, 32'h4203ba64};
test_input[30720:30727] = '{32'hc1f169ae, 32'hc24bbcae, 32'hc24c48e7, 32'hc2270f1e, 32'h40b06a66, 32'hc25c3aea, 32'h422b6b2f, 32'hc10ece87};
test_output[30720:30727] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h40b06a66, 32'h0, 32'h422b6b2f, 32'h0};
test_input[30728:30735] = '{32'h42b7e3dc, 32'hbfe6b002, 32'h4289767a, 32'h423c5f4d, 32'h42853971, 32'hc26f1642, 32'h4243c189, 32'hc2b82462};
test_output[30728:30735] = '{32'h42b7e3dc, 32'h0, 32'h4289767a, 32'h423c5f4d, 32'h42853971, 32'h0, 32'h4243c189, 32'h0};
test_input[30736:30743] = '{32'hc1d8a6d4, 32'h410b2d8c, 32'hc14c2f1f, 32'h4137c0c1, 32'hc2970b0c, 32'h42a88c42, 32'h41d42104, 32'hc22ceab2};
test_output[30736:30743] = '{32'h0, 32'h410b2d8c, 32'h0, 32'h4137c0c1, 32'h0, 32'h42a88c42, 32'h41d42104, 32'h0};
test_input[30744:30751] = '{32'h409a8d55, 32'hc2975b2d, 32'hc19e3cb9, 32'h42ae12f3, 32'h42be6bfd, 32'hc25322b1, 32'hc2989f57, 32'h42298dc7};
test_output[30744:30751] = '{32'h409a8d55, 32'h0, 32'h0, 32'h42ae12f3, 32'h42be6bfd, 32'h0, 32'h0, 32'h42298dc7};
test_input[30752:30759] = '{32'h4268b2c0, 32'h42bdc509, 32'hc2369215, 32'hc28f806b, 32'hc2bba9f7, 32'hc1a7cec7, 32'hc2c312b1, 32'h4206b0b6};
test_output[30752:30759] = '{32'h4268b2c0, 32'h42bdc509, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4206b0b6};
test_input[30760:30767] = '{32'h42c297b1, 32'hc1039a8c, 32'h4209365d, 32'hc268d30f, 32'hc2909c29, 32'h4260547d, 32'hc213eb26, 32'h3faa0773};
test_output[30760:30767] = '{32'h42c297b1, 32'h0, 32'h4209365d, 32'h0, 32'h0, 32'h4260547d, 32'h0, 32'h3faa0773};
test_input[30768:30775] = '{32'hc2822931, 32'hc1797152, 32'hc2624274, 32'h415f9c06, 32'hc04163a0, 32'hc2785cb1, 32'h428ea17d, 32'hc2b5699a};
test_output[30768:30775] = '{32'h0, 32'h0, 32'h0, 32'h415f9c06, 32'h0, 32'h0, 32'h428ea17d, 32'h0};
test_input[30776:30783] = '{32'h42af9395, 32'h429e3d9c, 32'hc19b9ae6, 32'h42a9deb3, 32'h41dc002f, 32'h42aebd8a, 32'hc2172dec, 32'hc26133ea};
test_output[30776:30783] = '{32'h42af9395, 32'h429e3d9c, 32'h0, 32'h42a9deb3, 32'h41dc002f, 32'h42aebd8a, 32'h0, 32'h0};
test_input[30784:30791] = '{32'h4253c465, 32'h40f30718, 32'h42a2fff5, 32'h4293b0d6, 32'h4230cee8, 32'hc28d1da8, 32'h41354adc, 32'hc2533b9c};
test_output[30784:30791] = '{32'h4253c465, 32'h40f30718, 32'h42a2fff5, 32'h4293b0d6, 32'h4230cee8, 32'h0, 32'h41354adc, 32'h0};
test_input[30792:30799] = '{32'h42256195, 32'h42a42d61, 32'hc04a75d2, 32'h422a78d7, 32'h4107c56f, 32'h421dd5b2, 32'h41d6a584, 32'hc2987fee};
test_output[30792:30799] = '{32'h42256195, 32'h42a42d61, 32'h0, 32'h422a78d7, 32'h4107c56f, 32'h421dd5b2, 32'h41d6a584, 32'h0};
test_input[30800:30807] = '{32'h427c4fe2, 32'h411c055d, 32'hc28591e5, 32'h408c8eab, 32'h4282182f, 32'hc1b94e97, 32'hc28147ea, 32'hc2a329b7};
test_output[30800:30807] = '{32'h427c4fe2, 32'h411c055d, 32'h0, 32'h408c8eab, 32'h4282182f, 32'h0, 32'h0, 32'h0};
test_input[30808:30815] = '{32'h4297da30, 32'hc2c0bde6, 32'h421db47d, 32'hc2c25841, 32'hc2120e84, 32'h428d7b7f, 32'h4258e79b, 32'h3e5e1bcc};
test_output[30808:30815] = '{32'h4297da30, 32'h0, 32'h421db47d, 32'h0, 32'h0, 32'h428d7b7f, 32'h4258e79b, 32'h3e5e1bcc};
test_input[30816:30823] = '{32'hc184a0ce, 32'h41f7d9a8, 32'h424936ff, 32'h42908c6b, 32'hc2657229, 32'hc1b5f499, 32'h4082e860, 32'hc2b49183};
test_output[30816:30823] = '{32'h0, 32'h41f7d9a8, 32'h424936ff, 32'h42908c6b, 32'h0, 32'h0, 32'h4082e860, 32'h0};
test_input[30824:30831] = '{32'hc28d792c, 32'h41341875, 32'h42754d06, 32'h420130ee, 32'hc24295bc, 32'hc2402a56, 32'hc09f30f4, 32'hc2492eab};
test_output[30824:30831] = '{32'h0, 32'h41341875, 32'h42754d06, 32'h420130ee, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30832:30839] = '{32'h4265e64d, 32'hc0dfb00a, 32'hc2203729, 32'h41b84207, 32'hc2a5a2bc, 32'h4294175e, 32'hc1e3db22, 32'h41fddce3};
test_output[30832:30839] = '{32'h4265e64d, 32'h0, 32'h0, 32'h41b84207, 32'h0, 32'h4294175e, 32'h0, 32'h41fddce3};
test_input[30840:30847] = '{32'h428e5c55, 32'h40c4bd44, 32'h423981c7, 32'hc14aa276, 32'hc2b485ab, 32'hc2a8fdbd, 32'hc26a3dba, 32'hc2bbdfa4};
test_output[30840:30847] = '{32'h428e5c55, 32'h40c4bd44, 32'h423981c7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[30848:30855] = '{32'h4263ffc0, 32'h424eba58, 32'h42ab79f3, 32'h4289424f, 32'hc2c2e7be, 32'h423ab3da, 32'h42be5db7, 32'h42a2d0d6};
test_output[30848:30855] = '{32'h4263ffc0, 32'h424eba58, 32'h42ab79f3, 32'h4289424f, 32'h0, 32'h423ab3da, 32'h42be5db7, 32'h42a2d0d6};
test_input[30856:30863] = '{32'h4264d5bd, 32'h422aab29, 32'hc23ef8ae, 32'h42084e59, 32'hc29f4edf, 32'h4298f692, 32'hc20ec4b0, 32'h42918764};
test_output[30856:30863] = '{32'h4264d5bd, 32'h422aab29, 32'h0, 32'h42084e59, 32'h0, 32'h4298f692, 32'h0, 32'h42918764};
test_input[30864:30871] = '{32'h4285646f, 32'hc1ff4b93, 32'h42bd2e1a, 32'hc2b47d22, 32'hc2b105ef, 32'h427231d2, 32'h4202023f, 32'hc1c576ef};
test_output[30864:30871] = '{32'h4285646f, 32'h0, 32'h42bd2e1a, 32'h0, 32'h0, 32'h427231d2, 32'h4202023f, 32'h0};
test_input[30872:30879] = '{32'h427d082a, 32'h42b630a9, 32'h3f8c1181, 32'hc23b9e78, 32'h42241717, 32'h4261f74f, 32'hc2023a9e, 32'h41b33685};
test_output[30872:30879] = '{32'h427d082a, 32'h42b630a9, 32'h3f8c1181, 32'h0, 32'h42241717, 32'h4261f74f, 32'h0, 32'h41b33685};
test_input[30880:30887] = '{32'hc2885899, 32'hc18b754c, 32'h42a0053c, 32'hc123da87, 32'h4180ca0c, 32'hc189e192, 32'h42abb98b, 32'h422a616e};
test_output[30880:30887] = '{32'h0, 32'h0, 32'h42a0053c, 32'h0, 32'h4180ca0c, 32'h0, 32'h42abb98b, 32'h422a616e};
test_input[30888:30895] = '{32'h427d60f2, 32'hc2b8d814, 32'h41cf3c33, 32'h42b66001, 32'h42c1dfe0, 32'hc073c153, 32'h4247f21c, 32'hc1b45c54};
test_output[30888:30895] = '{32'h427d60f2, 32'h0, 32'h41cf3c33, 32'h42b66001, 32'h42c1dfe0, 32'h0, 32'h4247f21c, 32'h0};
test_input[30896:30903] = '{32'hc202efbf, 32'h4288f931, 32'h42588d95, 32'hc1ca8223, 32'hc1d9a2cd, 32'hc291978c, 32'h42388439, 32'hc1e94f19};
test_output[30896:30903] = '{32'h0, 32'h4288f931, 32'h42588d95, 32'h0, 32'h0, 32'h0, 32'h42388439, 32'h0};
test_input[30904:30911] = '{32'hc1662bbe, 32'hc24ff0ad, 32'hc29fa69f, 32'h422d0b52, 32'h42c7f848, 32'hc195886f, 32'h41f40730, 32'hc0349365};
test_output[30904:30911] = '{32'h0, 32'h0, 32'h0, 32'h422d0b52, 32'h42c7f848, 32'h0, 32'h41f40730, 32'h0};
test_input[30912:30919] = '{32'h40ecd23e, 32'h42a5fef0, 32'hc154591a, 32'hc2ada5e5, 32'hc2b54b86, 32'hc1815a3f, 32'h42aed5e2, 32'hc2966f94};
test_output[30912:30919] = '{32'h40ecd23e, 32'h42a5fef0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42aed5e2, 32'h0};
test_input[30920:30927] = '{32'hc28994d6, 32'h4168ea8c, 32'h428d9ee0, 32'h422f516f, 32'h4229960f, 32'h4207d9d2, 32'h41c551f2, 32'h40e0b03e};
test_output[30920:30927] = '{32'h0, 32'h4168ea8c, 32'h428d9ee0, 32'h422f516f, 32'h4229960f, 32'h4207d9d2, 32'h41c551f2, 32'h40e0b03e};
test_input[30928:30935] = '{32'h40be1493, 32'h410d2d0b, 32'h41847756, 32'hc2c13be8, 32'hc20bd5eb, 32'hc205d9cc, 32'h429b4c28, 32'h410c7778};
test_output[30928:30935] = '{32'h40be1493, 32'h410d2d0b, 32'h41847756, 32'h0, 32'h0, 32'h0, 32'h429b4c28, 32'h410c7778};
test_input[30936:30943] = '{32'h42a19d39, 32'hc1d41239, 32'h42621d13, 32'hc12cb976, 32'h418878ef, 32'h426cc52d, 32'h42bdb4bd, 32'hc1953c97};
test_output[30936:30943] = '{32'h42a19d39, 32'h0, 32'h42621d13, 32'h0, 32'h418878ef, 32'h426cc52d, 32'h42bdb4bd, 32'h0};
test_input[30944:30951] = '{32'hc279f616, 32'h42c6bbc8, 32'h41976f25, 32'h42670ce5, 32'hc296e238, 32'hc2b772ff, 32'hc2886763, 32'h429f9ecd};
test_output[30944:30951] = '{32'h0, 32'h42c6bbc8, 32'h41976f25, 32'h42670ce5, 32'h0, 32'h0, 32'h0, 32'h429f9ecd};
test_input[30952:30959] = '{32'h41222c04, 32'hc29f8d5f, 32'hc1a7bd75, 32'h42601965, 32'h4218a85a, 32'h402caf65, 32'hc1abee81, 32'h4040279e};
test_output[30952:30959] = '{32'h41222c04, 32'h0, 32'h0, 32'h42601965, 32'h4218a85a, 32'h402caf65, 32'h0, 32'h4040279e};
test_input[30960:30967] = '{32'h42968185, 32'hc24bf739, 32'h427cd89c, 32'hc285bba4, 32'h420e83d9, 32'h42ac1610, 32'h42486edd, 32'h41147a41};
test_output[30960:30967] = '{32'h42968185, 32'h0, 32'h427cd89c, 32'h0, 32'h420e83d9, 32'h42ac1610, 32'h42486edd, 32'h41147a41};
test_input[30968:30975] = '{32'hc256edac, 32'hc130bfc5, 32'hc1cd9abc, 32'hc1c57271, 32'h4296c970, 32'hc12733b4, 32'hc2170f5a, 32'hc2b4e659};
test_output[30968:30975] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4296c970, 32'h0, 32'h0, 32'h0};
test_input[30976:30983] = '{32'h41c8e32d, 32'hc21c0181, 32'h426bfc04, 32'h4213f20a, 32'h41dca84c, 32'hc2c5fd0d, 32'hc29be8a9, 32'h422712e3};
test_output[30976:30983] = '{32'h41c8e32d, 32'h0, 32'h426bfc04, 32'h4213f20a, 32'h41dca84c, 32'h0, 32'h0, 32'h422712e3};
test_input[30984:30991] = '{32'h42227409, 32'hc28f544c, 32'h41429d94, 32'hc229e314, 32'hc2304fb7, 32'hc2b24f7f, 32'h41e2fbb5, 32'hc29c1e48};
test_output[30984:30991] = '{32'h42227409, 32'h0, 32'h41429d94, 32'h0, 32'h0, 32'h0, 32'h41e2fbb5, 32'h0};
test_input[30992:30999] = '{32'h4211eefc, 32'h412a5e43, 32'hbfb75c3d, 32'h40ec31bc, 32'hc0b5f60f, 32'h41f81000, 32'hc1d73484, 32'hc2096323};
test_output[30992:30999] = '{32'h4211eefc, 32'h412a5e43, 32'h0, 32'h40ec31bc, 32'h0, 32'h41f81000, 32'h0, 32'h0};
test_input[31000:31007] = '{32'hc0bf545d, 32'hc1be9beb, 32'h4270bf37, 32'h428c92c2, 32'hc195c0b2, 32'h4235be5e, 32'hc22351a6, 32'hc232baf9};
test_output[31000:31007] = '{32'h0, 32'h0, 32'h4270bf37, 32'h428c92c2, 32'h0, 32'h4235be5e, 32'h0, 32'h0};
test_input[31008:31015] = '{32'h424a58ab, 32'hc2b2a292, 32'h420c2523, 32'h405b7199, 32'hc2bfb3e0, 32'hc2c50c29, 32'h42ad9b25, 32'hc17144c4};
test_output[31008:31015] = '{32'h424a58ab, 32'h0, 32'h420c2523, 32'h405b7199, 32'h0, 32'h0, 32'h42ad9b25, 32'h0};
test_input[31016:31023] = '{32'h421efda8, 32'h42c17a07, 32'hc2c6b248, 32'h42933adf, 32'hc0850612, 32'hc22ec8ba, 32'hc2c386b4, 32'h41bebaf7};
test_output[31016:31023] = '{32'h421efda8, 32'h42c17a07, 32'h0, 32'h42933adf, 32'h0, 32'h0, 32'h0, 32'h41bebaf7};
test_input[31024:31031] = '{32'hc14795ee, 32'h421293a0, 32'hc28bde9f, 32'hc2893bb6, 32'hc2b0661c, 32'hc2c7a5f1, 32'hc288a6f2, 32'hc1a7e019};
test_output[31024:31031] = '{32'h0, 32'h421293a0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31032:31039] = '{32'h425ff056, 32'hc1d76136, 32'h42a1df1f, 32'h42b2f50c, 32'h4227614b, 32'h41d83bb0, 32'hc28b18e4, 32'h42b33851};
test_output[31032:31039] = '{32'h425ff056, 32'h0, 32'h42a1df1f, 32'h42b2f50c, 32'h4227614b, 32'h41d83bb0, 32'h0, 32'h42b33851};
test_input[31040:31047] = '{32'h419feb31, 32'h423d1be8, 32'h419cdb5f, 32'h41bcf041, 32'hc11b6c28, 32'h421359b5, 32'h3f0965cf, 32'hc2364505};
test_output[31040:31047] = '{32'h419feb31, 32'h423d1be8, 32'h419cdb5f, 32'h41bcf041, 32'h0, 32'h421359b5, 32'h3f0965cf, 32'h0};
test_input[31048:31055] = '{32'h42788f7f, 32'hc1ee1b6e, 32'h428287e2, 32'hc1005846, 32'hc24fc1a3, 32'h41dbc885, 32'hc221278a, 32'hc299c03b};
test_output[31048:31055] = '{32'h42788f7f, 32'h0, 32'h428287e2, 32'h0, 32'h0, 32'h41dbc885, 32'h0, 32'h0};
test_input[31056:31063] = '{32'h42ac0e79, 32'hc1a97ab9, 32'h42352cb8, 32'hc1b731ef, 32'hc28a757e, 32'hc21110d9, 32'hc23eb0a4, 32'h421f253b};
test_output[31056:31063] = '{32'h42ac0e79, 32'h0, 32'h42352cb8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h421f253b};
test_input[31064:31071] = '{32'hc1fd1c4e, 32'h41d091a1, 32'h41c002b0, 32'hc2a5745a, 32'hc29a0d54, 32'hc22d601a, 32'hc207db86, 32'h42af303b};
test_output[31064:31071] = '{32'h0, 32'h41d091a1, 32'h41c002b0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42af303b};
test_input[31072:31079] = '{32'hc2c7d2c7, 32'h4299d822, 32'hc25c6db9, 32'hc28d36a2, 32'h41ae4ce8, 32'hc20e8cde, 32'h4121cd2c, 32'h429f4a56};
test_output[31072:31079] = '{32'h0, 32'h4299d822, 32'h0, 32'h0, 32'h41ae4ce8, 32'h0, 32'h4121cd2c, 32'h429f4a56};
test_input[31080:31087] = '{32'h41de5690, 32'hc08ba840, 32'hc2290c04, 32'hc28cc839, 32'hc2b8b176, 32'hc0174bad, 32'h428bf99d, 32'hc199c74b};
test_output[31080:31087] = '{32'h41de5690, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428bf99d, 32'h0};
test_input[31088:31095] = '{32'hc0fc3078, 32'hc084875e, 32'h41d2d2e4, 32'hc1da2672, 32'hc1c9a461, 32'hc2b62bd8, 32'h41d9eda4, 32'h42960804};
test_output[31088:31095] = '{32'h0, 32'h0, 32'h41d2d2e4, 32'h0, 32'h0, 32'h0, 32'h41d9eda4, 32'h42960804};
test_input[31096:31103] = '{32'hc276ee1f, 32'h4282c189, 32'hc24cfc74, 32'h425fb55a, 32'h42c5e0a6, 32'h42933f42, 32'hc28278b0, 32'h42a9cadb};
test_output[31096:31103] = '{32'h0, 32'h4282c189, 32'h0, 32'h425fb55a, 32'h42c5e0a6, 32'h42933f42, 32'h0, 32'h42a9cadb};
test_input[31104:31111] = '{32'h4196ac93, 32'h42b5565c, 32'h4038fe8c, 32'hc2229543, 32'h421935ac, 32'hc2c03e03, 32'hc2924d62, 32'hc180e260};
test_output[31104:31111] = '{32'h4196ac93, 32'h42b5565c, 32'h4038fe8c, 32'h0, 32'h421935ac, 32'h0, 32'h0, 32'h0};
test_input[31112:31119] = '{32'hc283be4a, 32'h423853ea, 32'hc185ee7e, 32'hc20c74b1, 32'h410b79c0, 32'h42925ee3, 32'h420d86b8, 32'h4131a4ee};
test_output[31112:31119] = '{32'h0, 32'h423853ea, 32'h0, 32'h0, 32'h410b79c0, 32'h42925ee3, 32'h420d86b8, 32'h4131a4ee};
test_input[31120:31127] = '{32'hc2000ba3, 32'hc23d41da, 32'hc1845d7d, 32'h4144dba9, 32'hc28552dc, 32'hc1ba1d27, 32'h424c7732, 32'hc299b4d8};
test_output[31120:31127] = '{32'h0, 32'h0, 32'h0, 32'h4144dba9, 32'h0, 32'h0, 32'h424c7732, 32'h0};
test_input[31128:31135] = '{32'hc2258419, 32'hc29ebc43, 32'hc1dd3c85, 32'hc2a4d86d, 32'h421ef276, 32'h41a086e6, 32'h422c9fb2, 32'h409f3441};
test_output[31128:31135] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h421ef276, 32'h41a086e6, 32'h422c9fb2, 32'h409f3441};
test_input[31136:31143] = '{32'hc1551719, 32'hc2a2b71a, 32'h41247b24, 32'hc23d1674, 32'hc08e58c3, 32'hc25dd7a6, 32'hc29231d8, 32'hc24d26bc};
test_output[31136:31143] = '{32'h0, 32'h0, 32'h41247b24, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31144:31151] = '{32'hc25ee994, 32'h424dcda3, 32'hc2a654d6, 32'h42812e9f, 32'h42b790e7, 32'h42a30bea, 32'hc2912885, 32'h427a4464};
test_output[31144:31151] = '{32'h0, 32'h424dcda3, 32'h0, 32'h42812e9f, 32'h42b790e7, 32'h42a30bea, 32'h0, 32'h427a4464};
test_input[31152:31159] = '{32'hc2ae922a, 32'hc2b64cf5, 32'hc2b87256, 32'hc2bde590, 32'h4211cdf3, 32'hc2a615d9, 32'h422347a9, 32'h40f276e0};
test_output[31152:31159] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4211cdf3, 32'h0, 32'h422347a9, 32'h40f276e0};
test_input[31160:31167] = '{32'hc29da1bd, 32'h422e1fac, 32'h42454d49, 32'h41dcb38b, 32'hc26203df, 32'h42a84ed0, 32'hc23bb772, 32'h42b7097d};
test_output[31160:31167] = '{32'h0, 32'h422e1fac, 32'h42454d49, 32'h41dcb38b, 32'h0, 32'h42a84ed0, 32'h0, 32'h42b7097d};
test_input[31168:31175] = '{32'h3f67d21d, 32'h4229c494, 32'h42adc2c5, 32'h426d23df, 32'hc11d8034, 32'hc2923e97, 32'hc2837ec1, 32'hc20e380a};
test_output[31168:31175] = '{32'h3f67d21d, 32'h4229c494, 32'h42adc2c5, 32'h426d23df, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31176:31183] = '{32'hc200ca26, 32'hc15fbec9, 32'hc24b784f, 32'h42a884f7, 32'hc2c4ea84, 32'h4270e5ab, 32'h40b5d280, 32'h41ff8327};
test_output[31176:31183] = '{32'h0, 32'h0, 32'h0, 32'h42a884f7, 32'h0, 32'h4270e5ab, 32'h40b5d280, 32'h41ff8327};
test_input[31184:31191] = '{32'hc109cfd0, 32'hc1538783, 32'hc2a0112e, 32'h42c79946, 32'hbeaa0c98, 32'h428e67f5, 32'h424aa3c0, 32'h41ad9d39};
test_output[31184:31191] = '{32'h0, 32'h0, 32'h0, 32'h42c79946, 32'h0, 32'h428e67f5, 32'h424aa3c0, 32'h41ad9d39};
test_input[31192:31199] = '{32'hc03cd53b, 32'hc23e0672, 32'h425fe6ce, 32'h42aa2241, 32'h3efaebf6, 32'h41f78809, 32'hc20c4e2c, 32'h42b3f470};
test_output[31192:31199] = '{32'h0, 32'h0, 32'h425fe6ce, 32'h42aa2241, 32'h3efaebf6, 32'h41f78809, 32'h0, 32'h42b3f470};
test_input[31200:31207] = '{32'h42a9d43c, 32'h428410e6, 32'hc2219749, 32'hc1c5313a, 32'h426d22cf, 32'hc27d41df, 32'hc29d9a0f, 32'hc2b6be4f};
test_output[31200:31207] = '{32'h42a9d43c, 32'h428410e6, 32'h0, 32'h0, 32'h426d22cf, 32'h0, 32'h0, 32'h0};
test_input[31208:31215] = '{32'h4224aab6, 32'h42878e8a, 32'hc2576a8b, 32'h42b77855, 32'hc217f913, 32'h42234e1f, 32'h41bb6ba9, 32'hc1328280};
test_output[31208:31215] = '{32'h4224aab6, 32'h42878e8a, 32'h0, 32'h42b77855, 32'h0, 32'h42234e1f, 32'h41bb6ba9, 32'h0};
test_input[31216:31223] = '{32'hc2bdd714, 32'h41e08e11, 32'hc2923c6a, 32'hc29c2fa2, 32'hc24f9e5d, 32'h42a49fc3, 32'h42a5ad6e, 32'h41e4dbca};
test_output[31216:31223] = '{32'h0, 32'h41e08e11, 32'h0, 32'h0, 32'h0, 32'h42a49fc3, 32'h42a5ad6e, 32'h41e4dbca};
test_input[31224:31231] = '{32'h410bde76, 32'h3bef82ed, 32'hc2ac4f23, 32'hc22363f6, 32'hc23e3154, 32'hc26ab87c, 32'h41e7febf, 32'h429d0cdd};
test_output[31224:31231] = '{32'h410bde76, 32'h3bef82ed, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41e7febf, 32'h429d0cdd};
test_input[31232:31239] = '{32'h427762c0, 32'hc095a5d2, 32'hc2515e65, 32'h42618b60, 32'hc05f4481, 32'h4200e83d, 32'h429975e1, 32'hc2b5ec21};
test_output[31232:31239] = '{32'h427762c0, 32'h0, 32'h0, 32'h42618b60, 32'h0, 32'h4200e83d, 32'h429975e1, 32'h0};
test_input[31240:31247] = '{32'h41994965, 32'hc28c1b86, 32'hc2b7984f, 32'h42c39826, 32'h424d0cda, 32'h415d4cab, 32'hc25ab0c9, 32'h41cf738d};
test_output[31240:31247] = '{32'h41994965, 32'h0, 32'h0, 32'h42c39826, 32'h424d0cda, 32'h415d4cab, 32'h0, 32'h41cf738d};
test_input[31248:31255] = '{32'hc1453140, 32'h41d3be69, 32'h426472e7, 32'hc1da1502, 32'h42a2faa8, 32'hc1b6dcec, 32'hc28fa2c0, 32'hc26ea27c};
test_output[31248:31255] = '{32'h0, 32'h41d3be69, 32'h426472e7, 32'h0, 32'h42a2faa8, 32'h0, 32'h0, 32'h0};
test_input[31256:31263] = '{32'h42864b3b, 32'hc2a11fc7, 32'hc24f8baf, 32'h426b88a8, 32'hc1288c0a, 32'hc1eb7cac, 32'h42348161, 32'hc2492626};
test_output[31256:31263] = '{32'h42864b3b, 32'h0, 32'h0, 32'h426b88a8, 32'h0, 32'h0, 32'h42348161, 32'h0};
test_input[31264:31271] = '{32'hc198df1f, 32'h4223fbe7, 32'h42435a90, 32'h4202883f, 32'h428d10bf, 32'h42961da5, 32'h42af1b00, 32'h42a62f99};
test_output[31264:31271] = '{32'h0, 32'h4223fbe7, 32'h42435a90, 32'h4202883f, 32'h428d10bf, 32'h42961da5, 32'h42af1b00, 32'h42a62f99};
test_input[31272:31279] = '{32'hc2198e15, 32'hc1c38e62, 32'hc22c44f5, 32'hc2454805, 32'h410cae80, 32'hc29c5326, 32'hc23fac31, 32'hc2b8b2c8};
test_output[31272:31279] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h410cae80, 32'h0, 32'h0, 32'h0};
test_input[31280:31287] = '{32'hc2b882f7, 32'h42165ff8, 32'hc28140c9, 32'h4269ec9d, 32'h41bb2540, 32'hc204bd8f, 32'h4296bcc1, 32'hc2862fd7};
test_output[31280:31287] = '{32'h0, 32'h42165ff8, 32'h0, 32'h4269ec9d, 32'h41bb2540, 32'h0, 32'h4296bcc1, 32'h0};
test_input[31288:31295] = '{32'hc1778a21, 32'h4243bda9, 32'h41b5b954, 32'hc2a8433e, 32'hc290beac, 32'hc219bb18, 32'hc1b9a03a, 32'h4166e0b2};
test_output[31288:31295] = '{32'h0, 32'h4243bda9, 32'h41b5b954, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4166e0b2};
test_input[31296:31303] = '{32'h41860b67, 32'h42120e83, 32'hc28b4ce6, 32'hc253e7fa, 32'hc221f1c4, 32'hc2aa8fbb, 32'hc0d44860, 32'hc2541988};
test_output[31296:31303] = '{32'h41860b67, 32'h42120e83, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31304:31311] = '{32'h41e5a44a, 32'hc282d38e, 32'h42935468, 32'h42a2ec4c, 32'h42c5cf6c, 32'hc2c292d8, 32'hc29d28ec, 32'hc2c5a170};
test_output[31304:31311] = '{32'h41e5a44a, 32'h0, 32'h42935468, 32'h42a2ec4c, 32'h42c5cf6c, 32'h0, 32'h0, 32'h0};
test_input[31312:31319] = '{32'hc0861e46, 32'hc2441822, 32'h3f41a365, 32'hc1aa847c, 32'h4176130d, 32'hc2ba26a5, 32'h42125ed6, 32'hc256ac43};
test_output[31312:31319] = '{32'h0, 32'h0, 32'h3f41a365, 32'h0, 32'h4176130d, 32'h0, 32'h42125ed6, 32'h0};
test_input[31320:31327] = '{32'hc22290bc, 32'h41dc0949, 32'h428ce597, 32'hc29de932, 32'hc1590061, 32'h41ad9dff, 32'h428c6ede, 32'h41dfdd51};
test_output[31320:31327] = '{32'h0, 32'h41dc0949, 32'h428ce597, 32'h0, 32'h0, 32'h41ad9dff, 32'h428c6ede, 32'h41dfdd51};
test_input[31328:31335] = '{32'h42039785, 32'h403ab89a, 32'h4295e0f9, 32'h42c6683f, 32'hc2a6a117, 32'h422f9423, 32'hc29e5c1c, 32'hc23c0ae0};
test_output[31328:31335] = '{32'h42039785, 32'h403ab89a, 32'h4295e0f9, 32'h42c6683f, 32'h0, 32'h422f9423, 32'h0, 32'h0};
test_input[31336:31343] = '{32'h4203017a, 32'hc299e245, 32'hc24a6426, 32'h42582d60, 32'hc25a96f8, 32'h420bd1cb, 32'h4106fdec, 32'h42b9dc18};
test_output[31336:31343] = '{32'h4203017a, 32'h0, 32'h0, 32'h42582d60, 32'h0, 32'h420bd1cb, 32'h4106fdec, 32'h42b9dc18};
test_input[31344:31351] = '{32'h42a75941, 32'hc0a6981c, 32'h41726f65, 32'hc290a7f3, 32'h42a21c09, 32'h427e2dbb, 32'h3eeef422, 32'hc282e2bf};
test_output[31344:31351] = '{32'h42a75941, 32'h0, 32'h41726f65, 32'h0, 32'h42a21c09, 32'h427e2dbb, 32'h3eeef422, 32'h0};
test_input[31352:31359] = '{32'hc21eb87b, 32'h4296a0e8, 32'h42326f10, 32'hc1fd472f, 32'h427915e2, 32'h422bb3bf, 32'hc2475296, 32'h419f8dd5};
test_output[31352:31359] = '{32'h0, 32'h4296a0e8, 32'h42326f10, 32'h0, 32'h427915e2, 32'h422bb3bf, 32'h0, 32'h419f8dd5};
test_input[31360:31367] = '{32'hc2c322f1, 32'h41486de0, 32'hc2600c55, 32'hc26a5225, 32'hc2b03422, 32'h41e76b48, 32'h42af2c0a, 32'h42c3f505};
test_output[31360:31367] = '{32'h0, 32'h41486de0, 32'h0, 32'h0, 32'h0, 32'h41e76b48, 32'h42af2c0a, 32'h42c3f505};
test_input[31368:31375] = '{32'h429d2a5b, 32'hc15bc321, 32'h42b94b83, 32'hc21eae30, 32'h4178e3d0, 32'h42b578f8, 32'hc27d0f00, 32'h422914a7};
test_output[31368:31375] = '{32'h429d2a5b, 32'h0, 32'h42b94b83, 32'h0, 32'h4178e3d0, 32'h42b578f8, 32'h0, 32'h422914a7};
test_input[31376:31383] = '{32'hc29752e9, 32'hc2c5de72, 32'h42a9eb60, 32'h425d7f88, 32'hc29dc220, 32'h40e944e3, 32'h42b1cf53, 32'h42c4d7ec};
test_output[31376:31383] = '{32'h0, 32'h0, 32'h42a9eb60, 32'h425d7f88, 32'h0, 32'h40e944e3, 32'h42b1cf53, 32'h42c4d7ec};
test_input[31384:31391] = '{32'hc295661d, 32'h41fd8eed, 32'h4228a1d1, 32'h42572836, 32'h429dc7c8, 32'h42bfddb8, 32'h42063d88, 32'hc28f064e};
test_output[31384:31391] = '{32'h0, 32'h41fd8eed, 32'h4228a1d1, 32'h42572836, 32'h429dc7c8, 32'h42bfddb8, 32'h42063d88, 32'h0};
test_input[31392:31399] = '{32'hbf844569, 32'h42418970, 32'hc247f354, 32'hc161fe5c, 32'hc21d1cc6, 32'h42b1f571, 32'hc22fe5f4, 32'hc1d84e21};
test_output[31392:31399] = '{32'h0, 32'h42418970, 32'h0, 32'h0, 32'h0, 32'h42b1f571, 32'h0, 32'h0};
test_input[31400:31407] = '{32'h427d0df1, 32'h41c2074b, 32'h42be6da1, 32'h41f6df51, 32'hc1cf86c9, 32'hc2b0b07a, 32'hc0c89a84, 32'hbf83c736};
test_output[31400:31407] = '{32'h427d0df1, 32'h41c2074b, 32'h42be6da1, 32'h41f6df51, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31408:31415] = '{32'hc246b0ca, 32'h42601c97, 32'h41c10237, 32'hc28a9f14, 32'hc16a36eb, 32'hc2c45a96, 32'hc299d6b3, 32'hc202e733};
test_output[31408:31415] = '{32'h0, 32'h42601c97, 32'h41c10237, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31416:31423] = '{32'hc2bdd7d8, 32'h429ffb12, 32'hc1b510c1, 32'h42301b6e, 32'h422424e3, 32'h4020df07, 32'hc196cf11, 32'h427537fe};
test_output[31416:31423] = '{32'h0, 32'h429ffb12, 32'h0, 32'h42301b6e, 32'h422424e3, 32'h4020df07, 32'h0, 32'h427537fe};
test_input[31424:31431] = '{32'hc26c7df8, 32'hc2a5f38e, 32'hc23276d5, 32'hc1dc686a, 32'hc227d786, 32'h42357332, 32'h4288acff, 32'hc054b04b};
test_output[31424:31431] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42357332, 32'h4288acff, 32'h0};
test_input[31432:31439] = '{32'hc1ce76c3, 32'h42b5b58b, 32'hc281a542, 32'h4249c31f, 32'hc2c49bc0, 32'hc2c7f197, 32'h42831614, 32'hc29550d2};
test_output[31432:31439] = '{32'h0, 32'h42b5b58b, 32'h0, 32'h4249c31f, 32'h0, 32'h0, 32'h42831614, 32'h0};
test_input[31440:31447] = '{32'h429a419c, 32'h42c28497, 32'hc2a32823, 32'hc281fbe3, 32'hc1de929b, 32'hc2bbdaa9, 32'hc200f684, 32'hc2a81380};
test_output[31440:31447] = '{32'h429a419c, 32'h42c28497, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31448:31455] = '{32'h42adf68e, 32'hc27f6e2b, 32'h41c023d8, 32'h42279abe, 32'hc07a1a85, 32'h4193eeea, 32'h4293b927, 32'hc2996039};
test_output[31448:31455] = '{32'h42adf68e, 32'h0, 32'h41c023d8, 32'h42279abe, 32'h0, 32'h4193eeea, 32'h4293b927, 32'h0};
test_input[31456:31463] = '{32'hc15b888c, 32'h421100b0, 32'h42400487, 32'hc2bc20f5, 32'hc28168c9, 32'h41d3a049, 32'hc23139d1, 32'hc265df64};
test_output[31456:31463] = '{32'h0, 32'h421100b0, 32'h42400487, 32'h0, 32'h0, 32'h41d3a049, 32'h0, 32'h0};
test_input[31464:31471] = '{32'hc28d3e89, 32'h41713d48, 32'hc1c788d3, 32'h40e1dbbc, 32'h42bd5304, 32'h42c73a7b, 32'h40ce7af9, 32'hc28c837c};
test_output[31464:31471] = '{32'h0, 32'h41713d48, 32'h0, 32'h40e1dbbc, 32'h42bd5304, 32'h42c73a7b, 32'h40ce7af9, 32'h0};
test_input[31472:31479] = '{32'hc271f608, 32'hc21b3988, 32'h4098c94d, 32'h41603d91, 32'hc1a29bbd, 32'hc243c4e6, 32'h42838fd9, 32'h429b13ed};
test_output[31472:31479] = '{32'h0, 32'h0, 32'h4098c94d, 32'h41603d91, 32'h0, 32'h0, 32'h42838fd9, 32'h429b13ed};
test_input[31480:31487] = '{32'hc2913fad, 32'h425a5a58, 32'hc21e8cad, 32'h413728ea, 32'hc29963ba, 32'h40dce2e8, 32'h3e0bb3f0, 32'h42b1a0e0};
test_output[31480:31487] = '{32'h0, 32'h425a5a58, 32'h0, 32'h413728ea, 32'h0, 32'h40dce2e8, 32'h3e0bb3f0, 32'h42b1a0e0};
test_input[31488:31495] = '{32'hc2b83b4a, 32'hc291407e, 32'h425545a9, 32'h42c21dab, 32'hc23d24be, 32'hc05d607a, 32'hc2ac30fa, 32'hc243722e};
test_output[31488:31495] = '{32'h0, 32'h0, 32'h425545a9, 32'h42c21dab, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31496:31503] = '{32'h4209557c, 32'hc290befa, 32'h42a29f20, 32'h414e28d2, 32'hc24fcb04, 32'hc2b32145, 32'h420ab39a, 32'hc29401b4};
test_output[31496:31503] = '{32'h4209557c, 32'h0, 32'h42a29f20, 32'h414e28d2, 32'h0, 32'h0, 32'h420ab39a, 32'h0};
test_input[31504:31511] = '{32'h4280a651, 32'hc0adf106, 32'h42161e73, 32'hbfc4d423, 32'hc20d6724, 32'h42b67266, 32'hc0a4e199, 32'h425a7900};
test_output[31504:31511] = '{32'h4280a651, 32'h0, 32'h42161e73, 32'h0, 32'h0, 32'h42b67266, 32'h0, 32'h425a7900};
test_input[31512:31519] = '{32'hc29ce2a5, 32'h42808866, 32'h429c3823, 32'hc2c0953d, 32'h4225035d, 32'hc2c0372e, 32'h41ef8ac9, 32'hc0ba6d8d};
test_output[31512:31519] = '{32'h0, 32'h42808866, 32'h429c3823, 32'h0, 32'h4225035d, 32'h0, 32'h41ef8ac9, 32'h0};
test_input[31520:31527] = '{32'h40d2799a, 32'hc25b938f, 32'hc2a8691f, 32'hc1cf8d63, 32'h420c43b8, 32'h428cc6b1, 32'h42307f94, 32'hc20f4084};
test_output[31520:31527] = '{32'h40d2799a, 32'h0, 32'h0, 32'h0, 32'h420c43b8, 32'h428cc6b1, 32'h42307f94, 32'h0};
test_input[31528:31535] = '{32'hc2325cef, 32'h41f33f36, 32'hc0d143b7, 32'hc289273f, 32'hc24ae0c6, 32'h42b41e8a, 32'hc2b2554f, 32'hc28dc35a};
test_output[31528:31535] = '{32'h0, 32'h41f33f36, 32'h0, 32'h0, 32'h0, 32'h42b41e8a, 32'h0, 32'h0};
test_input[31536:31543] = '{32'h42844e6d, 32'h42850de5, 32'h42adf7cb, 32'hc1ed5a76, 32'hc28446da, 32'h413d0108, 32'hc2b4d00c, 32'h4288e854};
test_output[31536:31543] = '{32'h42844e6d, 32'h42850de5, 32'h42adf7cb, 32'h0, 32'h0, 32'h413d0108, 32'h0, 32'h4288e854};
test_input[31544:31551] = '{32'h42888a34, 32'h420b036c, 32'h42384fc3, 32'h4131328c, 32'hc2216c7f, 32'h425dd869, 32'hc1a14611, 32'h4294e0e1};
test_output[31544:31551] = '{32'h42888a34, 32'h420b036c, 32'h42384fc3, 32'h4131328c, 32'h0, 32'h425dd869, 32'h0, 32'h4294e0e1};
test_input[31552:31559] = '{32'hc2128734, 32'h4248ac4f, 32'h42a44343, 32'h41a2410c, 32'hc2b7c4c4, 32'hc1cabaa5, 32'h41c011f5, 32'h4244c15b};
test_output[31552:31559] = '{32'h0, 32'h4248ac4f, 32'h42a44343, 32'h41a2410c, 32'h0, 32'h0, 32'h41c011f5, 32'h4244c15b};
test_input[31560:31567] = '{32'hc28f5e86, 32'h4280d9c6, 32'h40b00354, 32'hbd826436, 32'h429a771c, 32'hc2009e7e, 32'hc245743c, 32'h42825b97};
test_output[31560:31567] = '{32'h0, 32'h4280d9c6, 32'h40b00354, 32'h0, 32'h429a771c, 32'h0, 32'h0, 32'h42825b97};
test_input[31568:31575] = '{32'hc2c2fd20, 32'hc1bbce7c, 32'hc27c54cc, 32'h42543d5c, 32'hc285ab53, 32'h424ef787, 32'h42589dd2, 32'h41331e95};
test_output[31568:31575] = '{32'h0, 32'h0, 32'h0, 32'h42543d5c, 32'h0, 32'h424ef787, 32'h42589dd2, 32'h41331e95};
test_input[31576:31583] = '{32'h41ebef52, 32'h42078993, 32'hc1a85dec, 32'hc2b63317, 32'hbf51f2cc, 32'h420e60f4, 32'hc1d2b427, 32'h411937ea};
test_output[31576:31583] = '{32'h41ebef52, 32'h42078993, 32'h0, 32'h0, 32'h0, 32'h420e60f4, 32'h0, 32'h411937ea};
test_input[31584:31591] = '{32'hc1f17371, 32'hc1590a9b, 32'hc1fe5f19, 32'h421dd64f, 32'hc2b36f7e, 32'h422e1792, 32'h42619aa1, 32'hc2309adb};
test_output[31584:31591] = '{32'h0, 32'h0, 32'h0, 32'h421dd64f, 32'h0, 32'h422e1792, 32'h42619aa1, 32'h0};
test_input[31592:31599] = '{32'hc1c52ef2, 32'hc12ab70f, 32'h428f19ce, 32'hc2c7f26a, 32'hc1d49cdc, 32'h42c0cae3, 32'h429abd0e, 32'hc213673e};
test_output[31592:31599] = '{32'h0, 32'h0, 32'h428f19ce, 32'h0, 32'h0, 32'h42c0cae3, 32'h429abd0e, 32'h0};
test_input[31600:31607] = '{32'hc22807de, 32'hc14594e7, 32'hc27a14d2, 32'hc1c597ef, 32'hc28717ef, 32'h4188170e, 32'h42693699, 32'hc2c4deeb};
test_output[31600:31607] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4188170e, 32'h42693699, 32'h0};
test_input[31608:31615] = '{32'h4280d3d5, 32'h42b09ed0, 32'hc29a1f66, 32'hc10198b5, 32'hc11a49b4, 32'hc29e6800, 32'h418ec7e1, 32'h41632d29};
test_output[31608:31615] = '{32'h4280d3d5, 32'h42b09ed0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h418ec7e1, 32'h41632d29};
test_input[31616:31623] = '{32'hc2311f1b, 32'h42285559, 32'hc2a55441, 32'h3fa386f2, 32'h426f02a4, 32'h423e2688, 32'h429d0495, 32'hc1d5eaff};
test_output[31616:31623] = '{32'h0, 32'h42285559, 32'h0, 32'h3fa386f2, 32'h426f02a4, 32'h423e2688, 32'h429d0495, 32'h0};
test_input[31624:31631] = '{32'h419d4afc, 32'hc2585cd5, 32'hc1bca84a, 32'h42bba950, 32'h4244c520, 32'hc25d89e5, 32'hc29e1e73, 32'hc2947a91};
test_output[31624:31631] = '{32'h419d4afc, 32'h0, 32'h0, 32'h42bba950, 32'h4244c520, 32'h0, 32'h0, 32'h0};
test_input[31632:31639] = '{32'h428b7eb3, 32'hc2a7ef2d, 32'h42be1846, 32'h426853a6, 32'hc24e7522, 32'hc28bf252, 32'h418c5d73, 32'h429fc9ff};
test_output[31632:31639] = '{32'h428b7eb3, 32'h0, 32'h42be1846, 32'h426853a6, 32'h0, 32'h0, 32'h418c5d73, 32'h429fc9ff};
test_input[31640:31647] = '{32'h41ca6d06, 32'h42a42229, 32'hc08960fe, 32'hc184bac3, 32'hc2bb9e89, 32'h42193aa2, 32'h41eab76b, 32'h418a445d};
test_output[31640:31647] = '{32'h41ca6d06, 32'h42a42229, 32'h0, 32'h0, 32'h0, 32'h42193aa2, 32'h41eab76b, 32'h418a445d};
test_input[31648:31655] = '{32'h40f55278, 32'h428b3d76, 32'hc0b4da3a, 32'hc2712362, 32'h416a7fe7, 32'h41fdfa49, 32'h4137735d, 32'h41b1ab63};
test_output[31648:31655] = '{32'h40f55278, 32'h428b3d76, 32'h0, 32'h0, 32'h416a7fe7, 32'h41fdfa49, 32'h4137735d, 32'h41b1ab63};
test_input[31656:31663] = '{32'hc102ee11, 32'hc2bcf88a, 32'hc2a7d1b1, 32'h42c42a53, 32'h42c6e421, 32'hc2972f23, 32'h42840f9a, 32'hc0a9d979};
test_output[31656:31663] = '{32'h0, 32'h0, 32'h0, 32'h42c42a53, 32'h42c6e421, 32'h0, 32'h42840f9a, 32'h0};
test_input[31664:31671] = '{32'hc154272c, 32'hc1a3f5e1, 32'h42b66520, 32'hc2318f6b, 32'h41ed7fed, 32'hc22aa9d6, 32'h42a54529, 32'h40be880a};
test_output[31664:31671] = '{32'h0, 32'h0, 32'h42b66520, 32'h0, 32'h41ed7fed, 32'h0, 32'h42a54529, 32'h40be880a};
test_input[31672:31679] = '{32'h4219fde8, 32'h4085aabd, 32'h41168460, 32'hc23f7e46, 32'hc1b285e4, 32'hc21c0295, 32'h4121f003, 32'h40e455fb};
test_output[31672:31679] = '{32'h4219fde8, 32'h4085aabd, 32'h41168460, 32'h0, 32'h0, 32'h0, 32'h4121f003, 32'h40e455fb};
test_input[31680:31687] = '{32'hc24b0be1, 32'hc265ac1c, 32'hc2b9e0c6, 32'hc2be8a60, 32'h41b3114a, 32'h4235209f, 32'hc2bdfcc2, 32'hc148cf34};
test_output[31680:31687] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41b3114a, 32'h4235209f, 32'h0, 32'h0};
test_input[31688:31695] = '{32'h42c37fd3, 32'hc1a22e03, 32'hc20b2e88, 32'hc257fe6d, 32'hc225551e, 32'hc26c1cea, 32'h41ad5b7d, 32'hc1e582e8};
test_output[31688:31695] = '{32'h42c37fd3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ad5b7d, 32'h0};
test_input[31696:31703] = '{32'hc23e98d2, 32'hc25bf1a5, 32'h42c36baa, 32'h425a2ce8, 32'hc2586daf, 32'hc0ab46ff, 32'h42686290, 32'h4250fce4};
test_output[31696:31703] = '{32'h0, 32'h0, 32'h42c36baa, 32'h425a2ce8, 32'h0, 32'h0, 32'h42686290, 32'h4250fce4};
test_input[31704:31711] = '{32'hc0bee6d6, 32'h419f6d7d, 32'hc24204bf, 32'hc112cfd6, 32'hc2b3e303, 32'hc173abab, 32'hc1c1990a, 32'h427fda36};
test_output[31704:31711] = '{32'h0, 32'h419f6d7d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427fda36};
test_input[31712:31719] = '{32'h4297ead1, 32'hc1d996a7, 32'h41da4f90, 32'h4282b972, 32'h413e3946, 32'h4044016b, 32'h4291629a, 32'h42bf676b};
test_output[31712:31719] = '{32'h4297ead1, 32'h0, 32'h41da4f90, 32'h4282b972, 32'h413e3946, 32'h4044016b, 32'h4291629a, 32'h42bf676b};
test_input[31720:31727] = '{32'hc2812166, 32'h42636061, 32'hc2b6fa8d, 32'h4273735d, 32'hc2b5bdde, 32'hc0ab00c1, 32'h409cd8f5, 32'hc259dfdc};
test_output[31720:31727] = '{32'h0, 32'h42636061, 32'h0, 32'h4273735d, 32'h0, 32'h0, 32'h409cd8f5, 32'h0};
test_input[31728:31735] = '{32'hc10e4dee, 32'hc2ad7755, 32'hc2c6a188, 32'h4242c115, 32'hc2b2e601, 32'h40ee30ad, 32'h4224fa9e, 32'h422d4f1a};
test_output[31728:31735] = '{32'h0, 32'h0, 32'h0, 32'h4242c115, 32'h0, 32'h40ee30ad, 32'h4224fa9e, 32'h422d4f1a};
test_input[31736:31743] = '{32'hc2220c82, 32'h4178cdbb, 32'hc2236be8, 32'h41fc56b3, 32'h41df8784, 32'h3fa58e44, 32'h41ad7702, 32'h422d2d04};
test_output[31736:31743] = '{32'h0, 32'h4178cdbb, 32'h0, 32'h41fc56b3, 32'h41df8784, 32'h3fa58e44, 32'h41ad7702, 32'h422d2d04};
test_input[31744:31751] = '{32'hc125bf71, 32'h4278aff4, 32'h421af53e, 32'h41cd12d0, 32'h4272a953, 32'h42177fd1, 32'h427763ec, 32'h429c8d7e};
test_output[31744:31751] = '{32'h0, 32'h4278aff4, 32'h421af53e, 32'h41cd12d0, 32'h4272a953, 32'h42177fd1, 32'h427763ec, 32'h429c8d7e};
test_input[31752:31759] = '{32'h42340690, 32'hc1fe7791, 32'h4211f9b3, 32'hbf84ed2c, 32'hc2950120, 32'h41f1113c, 32'hc29d179e, 32'hc27637e8};
test_output[31752:31759] = '{32'h42340690, 32'h0, 32'h4211f9b3, 32'h0, 32'h0, 32'h41f1113c, 32'h0, 32'h0};
test_input[31760:31767] = '{32'h42be2448, 32'hc2b740d1, 32'h421df426, 32'hc0a1ba6c, 32'hc2b56194, 32'h41e352fd, 32'h420257d1, 32'h421c8d1b};
test_output[31760:31767] = '{32'h42be2448, 32'h0, 32'h421df426, 32'h0, 32'h0, 32'h41e352fd, 32'h420257d1, 32'h421c8d1b};
test_input[31768:31775] = '{32'h42a8bef5, 32'h42ae6bb9, 32'h42bb44da, 32'h41d094d3, 32'hc2a64ecc, 32'hc106f675, 32'h42957922, 32'h42bd0e94};
test_output[31768:31775] = '{32'h42a8bef5, 32'h42ae6bb9, 32'h42bb44da, 32'h41d094d3, 32'h0, 32'h0, 32'h42957922, 32'h42bd0e94};
test_input[31776:31783] = '{32'hc1293c23, 32'hc0baae70, 32'h4179827e, 32'hc14d72ed, 32'h42ac573c, 32'hc292d5b3, 32'h4246ac69, 32'h428b170f};
test_output[31776:31783] = '{32'h0, 32'h0, 32'h4179827e, 32'h0, 32'h42ac573c, 32'h0, 32'h4246ac69, 32'h428b170f};
test_input[31784:31791] = '{32'hc2a443a9, 32'hc26b388b, 32'hc2aa54d1, 32'h4296d2c9, 32'h429e0596, 32'h429d1618, 32'hc2a68bdf, 32'h425dda71};
test_output[31784:31791] = '{32'h0, 32'h0, 32'h0, 32'h4296d2c9, 32'h429e0596, 32'h429d1618, 32'h0, 32'h425dda71};
test_input[31792:31799] = '{32'hc2aa38d6, 32'hc23cab58, 32'hc2011c1f, 32'h4255ce37, 32'hc1da3cf9, 32'hbffc2ee1, 32'h3efbc419, 32'h41e3aa71};
test_output[31792:31799] = '{32'h0, 32'h0, 32'h0, 32'h4255ce37, 32'h0, 32'h0, 32'h3efbc419, 32'h41e3aa71};
test_input[31800:31807] = '{32'hc2018540, 32'hc2be5cd6, 32'h41ce09ea, 32'h4156fcf6, 32'hc070084f, 32'hc2458331, 32'hc28cec84, 32'hc0eaa0ae};
test_output[31800:31807] = '{32'h0, 32'h0, 32'h41ce09ea, 32'h4156fcf6, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31808:31815] = '{32'h40e9d716, 32'h42b4c6a0, 32'hc192591f, 32'hc19c630d, 32'hc1e31ae0, 32'hc2020f59, 32'h429eccd1, 32'hc2a9ae8d};
test_output[31808:31815] = '{32'h40e9d716, 32'h42b4c6a0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429eccd1, 32'h0};
test_input[31816:31823] = '{32'h42337663, 32'hc2511012, 32'h42af3e9c, 32'h42aed897, 32'h42888b9b, 32'h41331ca7, 32'h42b4d3a5, 32'h423425a9};
test_output[31816:31823] = '{32'h42337663, 32'h0, 32'h42af3e9c, 32'h42aed897, 32'h42888b9b, 32'h41331ca7, 32'h42b4d3a5, 32'h423425a9};
test_input[31824:31831] = '{32'h41b6486b, 32'h4272e624, 32'hc204b0ec, 32'hc2241bc2, 32'hc2665f94, 32'h42a3c8ef, 32'h41dc5921, 32'h4185b29d};
test_output[31824:31831] = '{32'h41b6486b, 32'h4272e624, 32'h0, 32'h0, 32'h0, 32'h42a3c8ef, 32'h41dc5921, 32'h4185b29d};
test_input[31832:31839] = '{32'hc2828bb6, 32'h4298643e, 32'h429b66ab, 32'h428683ff, 32'hc1c53e50, 32'hc2b9a063, 32'h42b50756, 32'hc1f3316c};
test_output[31832:31839] = '{32'h0, 32'h4298643e, 32'h429b66ab, 32'h428683ff, 32'h0, 32'h0, 32'h42b50756, 32'h0};
test_input[31840:31847] = '{32'hc28b230f, 32'hc2866b8f, 32'hc1532b61, 32'hc1981aa7, 32'hc2bb9fc8, 32'hc2095c89, 32'h42028398, 32'hc224ea48};
test_output[31840:31847] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42028398, 32'h0};
test_input[31848:31855] = '{32'h42ba2c18, 32'h422e2442, 32'hc1a73249, 32'h428ed017, 32'hc1e9b676, 32'h42c1ba3b, 32'h4119db78, 32'hc283b8c3};
test_output[31848:31855] = '{32'h42ba2c18, 32'h422e2442, 32'h0, 32'h428ed017, 32'h0, 32'h42c1ba3b, 32'h4119db78, 32'h0};
test_input[31856:31863] = '{32'hc2aca9b2, 32'hc1e36fec, 32'h42967e18, 32'h3fd92ee3, 32'hc2b11295, 32'h4281bb58, 32'hc1881a8f, 32'h40ae4a8c};
test_output[31856:31863] = '{32'h0, 32'h0, 32'h42967e18, 32'h3fd92ee3, 32'h0, 32'h4281bb58, 32'h0, 32'h40ae4a8c};
test_input[31864:31871] = '{32'h429b6e8d, 32'h41c78a44, 32'h428d7052, 32'h42b4506a, 32'hc192bc52, 32'h41fdca37, 32'h4208f68e, 32'hc2962137};
test_output[31864:31871] = '{32'h429b6e8d, 32'h41c78a44, 32'h428d7052, 32'h42b4506a, 32'h0, 32'h41fdca37, 32'h4208f68e, 32'h0};
test_input[31872:31879] = '{32'hc1ff86c0, 32'hc208a23b, 32'hc26b9502, 32'h3ff634d0, 32'h419624cb, 32'hc18b714d, 32'h422e0197, 32'h420d0326};
test_output[31872:31879] = '{32'h0, 32'h0, 32'h0, 32'h3ff634d0, 32'h419624cb, 32'h0, 32'h422e0197, 32'h420d0326};
test_input[31880:31887] = '{32'h411b6a6d, 32'h4273af80, 32'hc0c4479a, 32'hc2ac4c6e, 32'h4100f319, 32'h42bd9ff7, 32'hc1a8a707, 32'hc2c50d16};
test_output[31880:31887] = '{32'h411b6a6d, 32'h4273af80, 32'h0, 32'h0, 32'h4100f319, 32'h42bd9ff7, 32'h0, 32'h0};
test_input[31888:31895] = '{32'h42aa2303, 32'h42bd565d, 32'h41d4f29e, 32'hc0322bfb, 32'h4292bc0d, 32'hc28888c0, 32'h4087f876, 32'hbf2b2999};
test_output[31888:31895] = '{32'h42aa2303, 32'h42bd565d, 32'h41d4f29e, 32'h0, 32'h4292bc0d, 32'h0, 32'h4087f876, 32'h0};
test_input[31896:31903] = '{32'hc222ea2c, 32'h42ab8092, 32'h4285b1ac, 32'h42c50aa2, 32'h4202f82a, 32'hc291ed92, 32'hc21c2152, 32'hc2a1fcb2};
test_output[31896:31903] = '{32'h0, 32'h42ab8092, 32'h4285b1ac, 32'h42c50aa2, 32'h4202f82a, 32'h0, 32'h0, 32'h0};
test_input[31904:31911] = '{32'hc26256c1, 32'hc20fc87e, 32'hc2329cf0, 32'hc1e31fd1, 32'h41e931e9, 32'hc086b0be, 32'h429420d8, 32'h42b93ccd};
test_output[31904:31911] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41e931e9, 32'h0, 32'h429420d8, 32'h42b93ccd};
test_input[31912:31919] = '{32'h425db3ee, 32'hc2a754ea, 32'hc2a01d02, 32'h42bab122, 32'hc0b2f3a4, 32'hc27a6f7c, 32'hc00ccffc, 32'h419e3db7};
test_output[31912:31919] = '{32'h425db3ee, 32'h0, 32'h0, 32'h42bab122, 32'h0, 32'h0, 32'h0, 32'h419e3db7};
test_input[31920:31927] = '{32'h42b363b1, 32'h426a11a5, 32'hc22748ff, 32'h40d44a5e, 32'h415ca5b8, 32'h42aedf7a, 32'hc18742f7, 32'h427748bd};
test_output[31920:31927] = '{32'h42b363b1, 32'h426a11a5, 32'h0, 32'h40d44a5e, 32'h415ca5b8, 32'h42aedf7a, 32'h0, 32'h427748bd};
test_input[31928:31935] = '{32'h42882574, 32'hc20703e6, 32'hc1c8712b, 32'hc05e6e78, 32'h42a83dd3, 32'hc17f7596, 32'h41814845, 32'h42b7c900};
test_output[31928:31935] = '{32'h42882574, 32'h0, 32'h0, 32'h0, 32'h42a83dd3, 32'h0, 32'h41814845, 32'h42b7c900};
test_input[31936:31943] = '{32'h42bf1658, 32'h429d42e8, 32'hc1a7e3e3, 32'h428d1ce8, 32'hc1794a76, 32'hc26d91e0, 32'h4039151f, 32'hc27930ea};
test_output[31936:31943] = '{32'h42bf1658, 32'h429d42e8, 32'h0, 32'h428d1ce8, 32'h0, 32'h0, 32'h4039151f, 32'h0};
test_input[31944:31951] = '{32'hc1c2bfb4, 32'h42ad7ab8, 32'h42c14c24, 32'hc249f36c, 32'hc0b6e1f1, 32'h40d5a7a4, 32'hc1586360, 32'h426340a0};
test_output[31944:31951] = '{32'h0, 32'h42ad7ab8, 32'h42c14c24, 32'h0, 32'h0, 32'h40d5a7a4, 32'h0, 32'h426340a0};
test_input[31952:31959] = '{32'h426ff42d, 32'hc29fceb7, 32'hc20f4193, 32'hc2a8a5c7, 32'hc2b67151, 32'hc2613811, 32'hc1ef2eaa, 32'hc13c946d};
test_output[31952:31959] = '{32'h426ff42d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[31960:31967] = '{32'h42b33465, 32'hc2872310, 32'h42bdef6e, 32'hc1aacc34, 32'hc2be1344, 32'hc2b35261, 32'h4248c6bb, 32'hc1a76d85};
test_output[31960:31967] = '{32'h42b33465, 32'h0, 32'h42bdef6e, 32'h0, 32'h0, 32'h0, 32'h4248c6bb, 32'h0};
test_input[31968:31975] = '{32'hc246d844, 32'h42585e0e, 32'hc2ba4c78, 32'hc282f19d, 32'h4205d61f, 32'hc27182a5, 32'h424abbf4, 32'h4118033f};
test_output[31968:31975] = '{32'h0, 32'h42585e0e, 32'h0, 32'h0, 32'h4205d61f, 32'h0, 32'h424abbf4, 32'h4118033f};
test_input[31976:31983] = '{32'h4237e3a6, 32'hc2256b7a, 32'hc1a0373c, 32'h42ba0109, 32'h42bfa36a, 32'h41bb2ba9, 32'hc2be840d, 32'h42c04a36};
test_output[31976:31983] = '{32'h4237e3a6, 32'h0, 32'h0, 32'h42ba0109, 32'h42bfa36a, 32'h41bb2ba9, 32'h0, 32'h42c04a36};
test_input[31984:31991] = '{32'h41fb9f50, 32'hc299d75d, 32'h429a00df, 32'hc286c9bb, 32'h42130feb, 32'h428bdc09, 32'hc2910ad6, 32'hc1820dd4};
test_output[31984:31991] = '{32'h41fb9f50, 32'h0, 32'h429a00df, 32'h0, 32'h42130feb, 32'h428bdc09, 32'h0, 32'h0};
test_input[31992:31999] = '{32'h41c8dd92, 32'h421db7f2, 32'h429aaf43, 32'hc2a0f8fd, 32'h42408c4f, 32'hc20c2d95, 32'hc295961a, 32'h42347d04};
test_output[31992:31999] = '{32'h41c8dd92, 32'h421db7f2, 32'h429aaf43, 32'h0, 32'h42408c4f, 32'h0, 32'h0, 32'h42347d04};
test_input[32000:32007] = '{32'h428c7f32, 32'hc1b2029c, 32'h422f3e06, 32'hc2a8983f, 32'h41921795, 32'h41fea496, 32'hc2a7ab59, 32'h4196bc2c};
test_output[32000:32007] = '{32'h428c7f32, 32'h0, 32'h422f3e06, 32'h0, 32'h41921795, 32'h41fea496, 32'h0, 32'h4196bc2c};
test_input[32008:32015] = '{32'h42878bb3, 32'hc17977c5, 32'h42571f99, 32'hc2645d84, 32'hc270f627, 32'h428d8b0b, 32'h428b4591, 32'h3dc7065f};
test_output[32008:32015] = '{32'h42878bb3, 32'h0, 32'h42571f99, 32'h0, 32'h0, 32'h428d8b0b, 32'h428b4591, 32'h3dc7065f};
test_input[32016:32023] = '{32'hc1920b7c, 32'hc233a354, 32'h42b8cd74, 32'h42bd737f, 32'h3fd3abbf, 32'hc26345b9, 32'hc2bb6508, 32'h42c7e790};
test_output[32016:32023] = '{32'h0, 32'h0, 32'h42b8cd74, 32'h42bd737f, 32'h3fd3abbf, 32'h0, 32'h0, 32'h42c7e790};
test_input[32024:32031] = '{32'hc1b50b76, 32'h4248a458, 32'hc20f60ba, 32'h422f4aaf, 32'h42179e26, 32'hc22b2217, 32'h410b0e6d, 32'h419f2a4d};
test_output[32024:32031] = '{32'h0, 32'h4248a458, 32'h0, 32'h422f4aaf, 32'h42179e26, 32'h0, 32'h410b0e6d, 32'h419f2a4d};
test_input[32032:32039] = '{32'hc2a33407, 32'h42827c4f, 32'hc1b767a3, 32'hc1c607f6, 32'h41996cf8, 32'h427b960f, 32'h3fc49f7a, 32'hc2164cf9};
test_output[32032:32039] = '{32'h0, 32'h42827c4f, 32'h0, 32'h0, 32'h41996cf8, 32'h427b960f, 32'h3fc49f7a, 32'h0};
test_input[32040:32047] = '{32'hc28272a4, 32'hc1325ac3, 32'hc24e7eb8, 32'h4280c666, 32'h42816445, 32'hc270534b, 32'h42c73fd2, 32'h421c9fc5};
test_output[32040:32047] = '{32'h0, 32'h0, 32'h0, 32'h4280c666, 32'h42816445, 32'h0, 32'h42c73fd2, 32'h421c9fc5};
test_input[32048:32055] = '{32'h4191ac9a, 32'hc2b75518, 32'h42a350d8, 32'h4250e5bc, 32'h41650dae, 32'hc20196ff, 32'h4231056e, 32'h4284d7b4};
test_output[32048:32055] = '{32'h4191ac9a, 32'h0, 32'h42a350d8, 32'h4250e5bc, 32'h41650dae, 32'h0, 32'h4231056e, 32'h4284d7b4};
test_input[32056:32063] = '{32'h41ad95d3, 32'h42bb7719, 32'h42a681f7, 32'hc0c9b497, 32'h4162a06c, 32'h42b4fea4, 32'hc29432bf, 32'h42b9a2c9};
test_output[32056:32063] = '{32'h41ad95d3, 32'h42bb7719, 32'h42a681f7, 32'h0, 32'h4162a06c, 32'h42b4fea4, 32'h0, 32'h42b9a2c9};
test_input[32064:32071] = '{32'hc2aa33b9, 32'hc2a1423b, 32'h424615ed, 32'h416f0f55, 32'h42352432, 32'h4291e5c5, 32'hc2c66505, 32'h429d2f31};
test_output[32064:32071] = '{32'h0, 32'h0, 32'h424615ed, 32'h416f0f55, 32'h42352432, 32'h4291e5c5, 32'h0, 32'h429d2f31};
test_input[32072:32079] = '{32'h421f5659, 32'hc1e40e51, 32'h42a24014, 32'h424e3d88, 32'h42b94327, 32'hc275daef, 32'hc24c2c36, 32'h42b2d731};
test_output[32072:32079] = '{32'h421f5659, 32'h0, 32'h42a24014, 32'h424e3d88, 32'h42b94327, 32'h0, 32'h0, 32'h42b2d731};
test_input[32080:32087] = '{32'h419b08ef, 32'hc2851371, 32'hc1afa0a1, 32'h42c2db2e, 32'h41ea0f47, 32'hc2a16d70, 32'hc15555c1, 32'h42728a9a};
test_output[32080:32087] = '{32'h419b08ef, 32'h0, 32'h0, 32'h42c2db2e, 32'h41ea0f47, 32'h0, 32'h0, 32'h42728a9a};
test_input[32088:32095] = '{32'h411a1994, 32'h42631cf5, 32'hc183fda3, 32'h428343f9, 32'hc2234818, 32'hc202dd23, 32'hc234170d, 32'h41a08d85};
test_output[32088:32095] = '{32'h411a1994, 32'h42631cf5, 32'h0, 32'h428343f9, 32'h0, 32'h0, 32'h0, 32'h41a08d85};
test_input[32096:32103] = '{32'h42c7bd00, 32'h4296775f, 32'hc2966270, 32'h4202c610, 32'hc096ff35, 32'hc11f8418, 32'h41ad2aef, 32'h4215f50a};
test_output[32096:32103] = '{32'h42c7bd00, 32'h4296775f, 32'h0, 32'h4202c610, 32'h0, 32'h0, 32'h41ad2aef, 32'h4215f50a};
test_input[32104:32111] = '{32'h426fb2ce, 32'h415ca971, 32'h42b1018d, 32'h4281d713, 32'hc2c01d0a, 32'h42a4ee49, 32'h42b57d5e, 32'h427ad2a0};
test_output[32104:32111] = '{32'h426fb2ce, 32'h415ca971, 32'h42b1018d, 32'h4281d713, 32'h0, 32'h42a4ee49, 32'h42b57d5e, 32'h427ad2a0};
test_input[32112:32119] = '{32'hc1ead445, 32'h41e0720d, 32'hc22fed48, 32'hc26106e8, 32'h42425daa, 32'h4271da46, 32'hc1bbd24b, 32'h42038330};
test_output[32112:32119] = '{32'h0, 32'h41e0720d, 32'h0, 32'h0, 32'h42425daa, 32'h4271da46, 32'h0, 32'h42038330};
test_input[32120:32127] = '{32'hc22b6e5e, 32'hc2bbd18d, 32'hbf0e641c, 32'h42a7a8bc, 32'hc23d97db, 32'hc2a79077, 32'hbf9c8533, 32'hc100a5fa};
test_output[32120:32127] = '{32'h0, 32'h0, 32'h0, 32'h42a7a8bc, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[32128:32135] = '{32'h40912a59, 32'hc20c0a30, 32'hc29e5202, 32'hc0e7bad4, 32'h429d446d, 32'h41dc905a, 32'hc1d2cc3a, 32'hc287405a};
test_output[32128:32135] = '{32'h40912a59, 32'h0, 32'h0, 32'h0, 32'h429d446d, 32'h41dc905a, 32'h0, 32'h0};
test_input[32136:32143] = '{32'h420cfeeb, 32'h424f0fb6, 32'hc1be778d, 32'h426f46b6, 32'h425d9b70, 32'h409d4877, 32'hc195891a, 32'h42248048};
test_output[32136:32143] = '{32'h420cfeeb, 32'h424f0fb6, 32'h0, 32'h426f46b6, 32'h425d9b70, 32'h409d4877, 32'h0, 32'h42248048};
test_input[32144:32151] = '{32'h42c1cabe, 32'h42c0f824, 32'h42a36e8a, 32'h42b59884, 32'hc1654f91, 32'h4273866a, 32'hc10de46c, 32'h427ffbcd};
test_output[32144:32151] = '{32'h42c1cabe, 32'h42c0f824, 32'h42a36e8a, 32'h42b59884, 32'h0, 32'h4273866a, 32'h0, 32'h427ffbcd};
test_input[32152:32159] = '{32'h42243967, 32'hc1dc30de, 32'h41f32cdd, 32'h41e1a50f, 32'h426a73e0, 32'hc2bf0a13, 32'h42166e8f, 32'hc2830ab5};
test_output[32152:32159] = '{32'h42243967, 32'h0, 32'h41f32cdd, 32'h41e1a50f, 32'h426a73e0, 32'h0, 32'h42166e8f, 32'h0};
test_input[32160:32167] = '{32'h4280cafb, 32'h4261c8de, 32'h42b3d583, 32'hc19aa240, 32'hc2c276d3, 32'h415207ef, 32'hc2a457e8, 32'hbfe8c31f};
test_output[32160:32167] = '{32'h4280cafb, 32'h4261c8de, 32'h42b3d583, 32'h0, 32'h0, 32'h415207ef, 32'h0, 32'h0};
test_input[32168:32175] = '{32'hc2af661a, 32'hc27074cf, 32'hc251de41, 32'hc24f6962, 32'hc20f29d1, 32'h410a0adb, 32'hc248be34, 32'h42252831};
test_output[32168:32175] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h410a0adb, 32'h0, 32'h42252831};
test_input[32176:32183] = '{32'hc19b92f7, 32'h42a32479, 32'hc149f076, 32'hc2c6b536, 32'h41da147d, 32'h42a6f56f, 32'hc24b29ea, 32'h4292b936};
test_output[32176:32183] = '{32'h0, 32'h42a32479, 32'h0, 32'h0, 32'h41da147d, 32'h42a6f56f, 32'h0, 32'h4292b936};
test_input[32184:32191] = '{32'hc257a33d, 32'hc25dfbbf, 32'h42c55a66, 32'h429a7f38, 32'hc22e9a20, 32'hc2abf468, 32'h426973c2, 32'hc2a577fc};
test_output[32184:32191] = '{32'h0, 32'h0, 32'h42c55a66, 32'h429a7f38, 32'h0, 32'h0, 32'h426973c2, 32'h0};
test_input[32192:32199] = '{32'h41e168fe, 32'hc2554dcb, 32'h423da5a4, 32'h4099f8d7, 32'h425cfed1, 32'h4223e735, 32'h423ab360, 32'hc2ac4724};
test_output[32192:32199] = '{32'h41e168fe, 32'h0, 32'h423da5a4, 32'h4099f8d7, 32'h425cfed1, 32'h4223e735, 32'h423ab360, 32'h0};
test_input[32200:32207] = '{32'h4283a4d7, 32'hc288609c, 32'hc2acaa39, 32'h42be7864, 32'hc227d46a, 32'h423a5ff1, 32'hc25a6413, 32'hc2a93b95};
test_output[32200:32207] = '{32'h4283a4d7, 32'h0, 32'h0, 32'h42be7864, 32'h0, 32'h423a5ff1, 32'h0, 32'h0};
test_input[32208:32215] = '{32'h42606f3e, 32'hc14cabaf, 32'h4098cfb8, 32'h4155788b, 32'h42955800, 32'h425bb200, 32'hc2a3023f, 32'hc1f874cf};
test_output[32208:32215] = '{32'h42606f3e, 32'h0, 32'h4098cfb8, 32'h4155788b, 32'h42955800, 32'h425bb200, 32'h0, 32'h0};
test_input[32216:32223] = '{32'h42be57ba, 32'hc298611d, 32'h429f9307, 32'hc257c2c7, 32'h42c113d3, 32'h4244c71a, 32'hc1fb6840, 32'hc15fe8bf};
test_output[32216:32223] = '{32'h42be57ba, 32'h0, 32'h429f9307, 32'h0, 32'h42c113d3, 32'h4244c71a, 32'h0, 32'h0};
test_input[32224:32231] = '{32'hc26fe62a, 32'hc0eac2e1, 32'h4290785a, 32'h4215106d, 32'hc263b7a9, 32'hc2a7f346, 32'h4019506f, 32'hc1b2836c};
test_output[32224:32231] = '{32'h0, 32'h0, 32'h4290785a, 32'h4215106d, 32'h0, 32'h0, 32'h4019506f, 32'h0};
test_input[32232:32239] = '{32'h42a206b9, 32'hc265163f, 32'h4294b836, 32'hc251025b, 32'hc2c62228, 32'hc273de6f, 32'hc1f4118c, 32'h41d62986};
test_output[32232:32239] = '{32'h42a206b9, 32'h0, 32'h4294b836, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41d62986};
test_input[32240:32247] = '{32'hc1a20cec, 32'hc2984cad, 32'hc206d509, 32'hc23a1286, 32'hc1751a67, 32'h419f965b, 32'h422504b2, 32'hc2b9a913};
test_output[32240:32247] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h419f965b, 32'h422504b2, 32'h0};
test_input[32248:32255] = '{32'h4268fe61, 32'h41a43c87, 32'hc27a98b6, 32'hc1069653, 32'h429cd78f, 32'hc1ae3c08, 32'hc2c1d8cf, 32'hc2728838};
test_output[32248:32255] = '{32'h4268fe61, 32'h41a43c87, 32'h0, 32'h0, 32'h429cd78f, 32'h0, 32'h0, 32'h0};
test_input[32256:32263] = '{32'hc2445782, 32'hc287dc90, 32'h41dc946d, 32'hc27c381d, 32'h42b2a04c, 32'hc10af209, 32'h42bba5dd, 32'hc2a4981c};
test_output[32256:32263] = '{32'h0, 32'h0, 32'h41dc946d, 32'h0, 32'h42b2a04c, 32'h0, 32'h42bba5dd, 32'h0};
test_input[32264:32271] = '{32'h421bad68, 32'hc1ad6522, 32'hc19f590e, 32'h42589aea, 32'h4208991d, 32'h4193a981, 32'h41d64de1, 32'h40932154};
test_output[32264:32271] = '{32'h421bad68, 32'h0, 32'h0, 32'h42589aea, 32'h4208991d, 32'h4193a981, 32'h41d64de1, 32'h40932154};
test_input[32272:32279] = '{32'hc2c356f0, 32'hc2998e94, 32'h40ce3bbd, 32'h42509d3f, 32'h416f9d0b, 32'h41a8c481, 32'h42c7441e, 32'hbe09ed5f};
test_output[32272:32279] = '{32'h0, 32'h0, 32'h40ce3bbd, 32'h42509d3f, 32'h416f9d0b, 32'h41a8c481, 32'h42c7441e, 32'h0};
test_input[32280:32287] = '{32'hc2815fdc, 32'h42c2fea2, 32'hc20e5297, 32'h419683a0, 32'hc1e18a67, 32'h42970734, 32'h428ba9f2, 32'h4297ae8d};
test_output[32280:32287] = '{32'h0, 32'h42c2fea2, 32'h0, 32'h419683a0, 32'h0, 32'h42970734, 32'h428ba9f2, 32'h4297ae8d};
test_input[32288:32295] = '{32'hbf3b3546, 32'hc1c2ea49, 32'h42476aea, 32'hc12d2fd9, 32'h4210a993, 32'hc2458ff5, 32'h426ba67d, 32'h4268285a};
test_output[32288:32295] = '{32'h0, 32'h0, 32'h42476aea, 32'h0, 32'h4210a993, 32'h0, 32'h426ba67d, 32'h4268285a};
test_input[32296:32303] = '{32'h4223b51c, 32'hc16f3d06, 32'hc27be4fc, 32'hc0d705fb, 32'h420a6f2d, 32'h42c0fa84, 32'h42b184de, 32'hbf4dd400};
test_output[32296:32303] = '{32'h4223b51c, 32'h0, 32'h0, 32'h0, 32'h420a6f2d, 32'h42c0fa84, 32'h42b184de, 32'h0};
test_input[32304:32311] = '{32'hc1b4363e, 32'hc20f2380, 32'hc2b8283e, 32'hc2c4e85a, 32'h41c214f2, 32'h418436b6, 32'hc1ee1778, 32'hc093c695};
test_output[32304:32311] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41c214f2, 32'h418436b6, 32'h0, 32'h0};
test_input[32312:32319] = '{32'hc2408b7c, 32'hc2233c8d, 32'h4135bb6b, 32'h42c6c5f9, 32'hc19a4d7a, 32'hc2beb6a8, 32'h42292a4a, 32'h422d0dc3};
test_output[32312:32319] = '{32'h0, 32'h0, 32'h4135bb6b, 32'h42c6c5f9, 32'h0, 32'h0, 32'h42292a4a, 32'h422d0dc3};
test_input[32320:32327] = '{32'hc2aaa978, 32'hc18c16a4, 32'h421b9cfa, 32'h427d77b5, 32'hc16cd34e, 32'hc220c4dc, 32'h42c6a197, 32'h42387e1c};
test_output[32320:32327] = '{32'h0, 32'h0, 32'h421b9cfa, 32'h427d77b5, 32'h0, 32'h0, 32'h42c6a197, 32'h42387e1c};
test_input[32328:32335] = '{32'hc071bc33, 32'h422dd476, 32'hc1d214e1, 32'h42008127, 32'hc1ea0709, 32'hc2af5c6f, 32'hc28751ef, 32'h42c3ed6f};
test_output[32328:32335] = '{32'h0, 32'h422dd476, 32'h0, 32'h42008127, 32'h0, 32'h0, 32'h0, 32'h42c3ed6f};
test_input[32336:32343] = '{32'h410085aa, 32'h424bcf56, 32'hc2222d4f, 32'hc12aacfc, 32'h41e080c0, 32'hc28881da, 32'hc16fd2b7, 32'h42196938};
test_output[32336:32343] = '{32'h410085aa, 32'h424bcf56, 32'h0, 32'h0, 32'h41e080c0, 32'h0, 32'h0, 32'h42196938};
test_input[32344:32351] = '{32'hc2aa586e, 32'h413a12aa, 32'hc2218298, 32'hc0fe8191, 32'h42644199, 32'h42b7c9ce, 32'hc261a643, 32'hc0c26a48};
test_output[32344:32351] = '{32'h0, 32'h413a12aa, 32'h0, 32'h0, 32'h42644199, 32'h42b7c9ce, 32'h0, 32'h0};
test_input[32352:32359] = '{32'h42332323, 32'hc27cacef, 32'hc1ff1b47, 32'hc28662a9, 32'h4227b07b, 32'hc2a2347d, 32'h3fcb48ab, 32'h41dd6320};
test_output[32352:32359] = '{32'h42332323, 32'h0, 32'h0, 32'h0, 32'h4227b07b, 32'h0, 32'h3fcb48ab, 32'h41dd6320};
test_input[32360:32367] = '{32'h410324de, 32'hc2afe85c, 32'h4109aaeb, 32'h42b6bf1d, 32'h4215e8b1, 32'h41b423ce, 32'hc26572b5, 32'h429d882b};
test_output[32360:32367] = '{32'h410324de, 32'h0, 32'h4109aaeb, 32'h42b6bf1d, 32'h4215e8b1, 32'h41b423ce, 32'h0, 32'h429d882b};
test_input[32368:32375] = '{32'hc2bab9b5, 32'h42617201, 32'hc244fea1, 32'h42b944ac, 32'hc120d05d, 32'hc2ba8c9d, 32'h42ad6e82, 32'hc131cda7};
test_output[32368:32375] = '{32'h0, 32'h42617201, 32'h0, 32'h42b944ac, 32'h0, 32'h0, 32'h42ad6e82, 32'h0};
test_input[32376:32383] = '{32'hc23f8ccd, 32'h4271dda7, 32'h40017384, 32'hc245aabf, 32'hc28cf8b0, 32'h42808ff9, 32'h41e82930, 32'h410c9c04};
test_output[32376:32383] = '{32'h0, 32'h4271dda7, 32'h40017384, 32'h0, 32'h0, 32'h42808ff9, 32'h41e82930, 32'h410c9c04};
test_input[32384:32391] = '{32'h4179492c, 32'h42956e75, 32'h419fcb02, 32'hc1b75b8c, 32'h4121e54a, 32'hc275270a, 32'hc253958a, 32'h429262ca};
test_output[32384:32391] = '{32'h4179492c, 32'h42956e75, 32'h419fcb02, 32'h0, 32'h4121e54a, 32'h0, 32'h0, 32'h429262ca};
test_input[32392:32399] = '{32'hc0005065, 32'hc2c49772, 32'h4292067a, 32'hc2c30b6d, 32'h41bf8c50, 32'hc1521f4d, 32'h4142a720, 32'h42b5838f};
test_output[32392:32399] = '{32'h0, 32'h0, 32'h4292067a, 32'h0, 32'h41bf8c50, 32'h0, 32'h4142a720, 32'h42b5838f};
test_input[32400:32407] = '{32'hc25b9709, 32'h42c4f10d, 32'h422fbdbd, 32'h426aa8d4, 32'h42c7692a, 32'h4254511c, 32'hc2994ade, 32'hc2a56350};
test_output[32400:32407] = '{32'h0, 32'h42c4f10d, 32'h422fbdbd, 32'h426aa8d4, 32'h42c7692a, 32'h4254511c, 32'h0, 32'h0};
test_input[32408:32415] = '{32'h429b725d, 32'h4187f96b, 32'hc285e1f9, 32'hc28c51fc, 32'hc10ed467, 32'hc210f030, 32'h4196bb86, 32'h428ca736};
test_output[32408:32415] = '{32'h429b725d, 32'h4187f96b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4196bb86, 32'h428ca736};
test_input[32416:32423] = '{32'hc088944a, 32'h42622304, 32'hc259ce2d, 32'h423cc4d0, 32'hc2787673, 32'h41b550a5, 32'hc05f225d, 32'h42b6fd5b};
test_output[32416:32423] = '{32'h0, 32'h42622304, 32'h0, 32'h423cc4d0, 32'h0, 32'h41b550a5, 32'h0, 32'h42b6fd5b};
test_input[32424:32431] = '{32'h425c4a22, 32'hc2c740aa, 32'hc2b786b0, 32'hc21e8d40, 32'hc29e6a47, 32'h4270e70d, 32'h41281fdb, 32'h421c75c3};
test_output[32424:32431] = '{32'h425c4a22, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4270e70d, 32'h41281fdb, 32'h421c75c3};
test_input[32432:32439] = '{32'h424283af, 32'hc2ad5166, 32'h42a4608a, 32'h42c066b4, 32'hc25737f1, 32'h42574c26, 32'h4285efbd, 32'hc2bb13d5};
test_output[32432:32439] = '{32'h424283af, 32'h0, 32'h42a4608a, 32'h42c066b4, 32'h0, 32'h42574c26, 32'h4285efbd, 32'h0};
test_input[32440:32447] = '{32'h42b91694, 32'hc2123cf9, 32'hc1d50ad8, 32'h42b31daa, 32'hc115cc53, 32'hc28e6ea6, 32'h3fecab65, 32'hc118eb37};
test_output[32440:32447] = '{32'h42b91694, 32'h0, 32'h0, 32'h42b31daa, 32'h0, 32'h0, 32'h3fecab65, 32'h0};
test_input[32448:32455] = '{32'hc2a18fdc, 32'hc2b6a8a3, 32'h422e4500, 32'h42a5384a, 32'hc2c36c29, 32'h4288ddb5, 32'h40d6d9b6, 32'hc10e314d};
test_output[32448:32455] = '{32'h0, 32'h0, 32'h422e4500, 32'h42a5384a, 32'h0, 32'h4288ddb5, 32'h40d6d9b6, 32'h0};
test_input[32456:32463] = '{32'h4184c8ed, 32'h41ea7301, 32'hc233129f, 32'h427332c6, 32'h41c1d091, 32'h42bfef44, 32'h42c5a3f2, 32'h427911ef};
test_output[32456:32463] = '{32'h4184c8ed, 32'h41ea7301, 32'h0, 32'h427332c6, 32'h41c1d091, 32'h42bfef44, 32'h42c5a3f2, 32'h427911ef};
test_input[32464:32471] = '{32'hc225cb13, 32'h429e1efb, 32'h42272b36, 32'hc251fdc5, 32'hc284991e, 32'hc2afcabf, 32'hc28adf51, 32'h42846d11};
test_output[32464:32471] = '{32'h0, 32'h429e1efb, 32'h42272b36, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42846d11};
test_input[32472:32479] = '{32'hc09a6178, 32'hc10eee58, 32'h414f0b5e, 32'hc0017f72, 32'h42a49230, 32'h413ec152, 32'h42bd995e, 32'hc2c157cb};
test_output[32472:32479] = '{32'h0, 32'h0, 32'h414f0b5e, 32'h0, 32'h42a49230, 32'h413ec152, 32'h42bd995e, 32'h0};
test_input[32480:32487] = '{32'hc2bb1217, 32'h420907bc, 32'h4238560f, 32'hbfc15ec1, 32'hc1404dac, 32'h428d4d46, 32'hc2bfac57, 32'h4239670a};
test_output[32480:32487] = '{32'h0, 32'h420907bc, 32'h4238560f, 32'h0, 32'h0, 32'h428d4d46, 32'h0, 32'h4239670a};
test_input[32488:32495] = '{32'h4222fe91, 32'hc250ff8d, 32'h428d720b, 32'hc243a4e5, 32'hc29b6e62, 32'hc2b9ac42, 32'hc2ab916d, 32'hc18b703d};
test_output[32488:32495] = '{32'h4222fe91, 32'h0, 32'h428d720b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[32496:32503] = '{32'h428e5c38, 32'h4263ceb3, 32'h4237f519, 32'hc1b549df, 32'hc18876a7, 32'hc214338f, 32'h4101ee91, 32'h428c5990};
test_output[32496:32503] = '{32'h428e5c38, 32'h4263ceb3, 32'h4237f519, 32'h0, 32'h0, 32'h0, 32'h4101ee91, 32'h428c5990};
test_input[32504:32511] = '{32'h4189f8ed, 32'h42b25729, 32'hc1948b34, 32'hc2298a69, 32'h42308a77, 32'hc2bc7039, 32'hc2b83202, 32'hc24070b3};
test_output[32504:32511] = '{32'h4189f8ed, 32'h42b25729, 32'h0, 32'h0, 32'h42308a77, 32'h0, 32'h0, 32'h0};
test_input[32512:32519] = '{32'hc08f854e, 32'hc12200e2, 32'hbfbdfea3, 32'hc14cdbd2, 32'hc18e3758, 32'hc220bc9b, 32'hc2a77171, 32'h413118d7};
test_output[32512:32519] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h413118d7};
test_input[32520:32527] = '{32'h41311894, 32'hc1f15054, 32'h3f490e36, 32'hc19082a1, 32'hc0c100b8, 32'hc08f6ee4, 32'h421593c5, 32'h420fac98};
test_output[32520:32527] = '{32'h41311894, 32'h0, 32'h3f490e36, 32'h0, 32'h0, 32'h0, 32'h421593c5, 32'h420fac98};
test_input[32528:32535] = '{32'h426af175, 32'hc270a251, 32'h4139ab44, 32'hc2a0e3f6, 32'hc2739d33, 32'hc2ba7e40, 32'hc2acf7b8, 32'h42456abc};
test_output[32528:32535] = '{32'h426af175, 32'h0, 32'h4139ab44, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42456abc};
test_input[32536:32543] = '{32'hc2c2d480, 32'hc1ae5b5a, 32'h42826a00, 32'h41c9fcd1, 32'hc0d64ff3, 32'h3f183b4c, 32'h41a8bb0d, 32'h42ab2bc8};
test_output[32536:32543] = '{32'h0, 32'h0, 32'h42826a00, 32'h41c9fcd1, 32'h0, 32'h3f183b4c, 32'h41a8bb0d, 32'h42ab2bc8};
test_input[32544:32551] = '{32'h41a66843, 32'hc1d4c863, 32'h41f0ccc1, 32'h427cbf1f, 32'hc29970ed, 32'hc1bbbadf, 32'hc2abf1f4, 32'h4230945e};
test_output[32544:32551] = '{32'h41a66843, 32'h0, 32'h41f0ccc1, 32'h427cbf1f, 32'h0, 32'h0, 32'h0, 32'h4230945e};
test_input[32552:32559] = '{32'hc2a7a5bd, 32'hc2ae896d, 32'hc215e6bd, 32'h4217f8c1, 32'hc1d5fe34, 32'hc14df796, 32'h422aeb92, 32'h40d98068};
test_output[32552:32559] = '{32'h0, 32'h0, 32'h0, 32'h4217f8c1, 32'h0, 32'h0, 32'h422aeb92, 32'h40d98068};
test_input[32560:32567] = '{32'h40f39d2c, 32'h42bd5e34, 32'hc1d10009, 32'hc21e5f1c, 32'hc28ba2f5, 32'hc281f24f, 32'h3f3725a5, 32'h41ab3272};
test_output[32560:32567] = '{32'h40f39d2c, 32'h42bd5e34, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3f3725a5, 32'h41ab3272};
test_input[32568:32575] = '{32'h42444c41, 32'h4191d424, 32'hc248e7a9, 32'hc1ee63f1, 32'hc23c5f5f, 32'hc2aceca4, 32'h4213d4ca, 32'h41fd736f};
test_output[32568:32575] = '{32'h42444c41, 32'h4191d424, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4213d4ca, 32'h41fd736f};
test_input[32576:32583] = '{32'h418d4e10, 32'hc23f431d, 32'h4229b6b6, 32'h42685286, 32'hc2bb02e9, 32'hc2a4f4e1, 32'hc2b65ae9, 32'h42b12328};
test_output[32576:32583] = '{32'h418d4e10, 32'h0, 32'h4229b6b6, 32'h42685286, 32'h0, 32'h0, 32'h0, 32'h42b12328};
test_input[32584:32591] = '{32'hc2092166, 32'hc2ad1ec2, 32'hc124626c, 32'hc1c3d0b1, 32'hc28c0edc, 32'hc2638489, 32'hc2c017a8, 32'h41ff5269};
test_output[32584:32591] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41ff5269};
test_input[32592:32599] = '{32'h42932f9f, 32'hc29c6ab1, 32'hc12a385e, 32'h4265df7a, 32'h42b772be, 32'hc1bf83f4, 32'h4238875f, 32'hc295aebc};
test_output[32592:32599] = '{32'h42932f9f, 32'h0, 32'h0, 32'h4265df7a, 32'h42b772be, 32'h0, 32'h4238875f, 32'h0};
test_input[32600:32607] = '{32'h428055f5, 32'hc215b56b, 32'h42aa52e9, 32'hc229edad, 32'h41cc6a13, 32'hc25855e3, 32'h41aa0503, 32'h4174f6eb};
test_output[32600:32607] = '{32'h428055f5, 32'h0, 32'h42aa52e9, 32'h0, 32'h41cc6a13, 32'h0, 32'h41aa0503, 32'h4174f6eb};
test_input[32608:32615] = '{32'hc1f035de, 32'h400de48f, 32'h42c71b77, 32'hc112ae4c, 32'h424a4059, 32'h406adee6, 32'h427f48e8, 32'h41833891};
test_output[32608:32615] = '{32'h0, 32'h400de48f, 32'h42c71b77, 32'h0, 32'h424a4059, 32'h406adee6, 32'h427f48e8, 32'h41833891};
test_input[32616:32623] = '{32'h426819a9, 32'h415ea2be, 32'h4223e848, 32'h42371fc2, 32'hc29d75a9, 32'h42aabcef, 32'h4221f713, 32'hc2c7ae5f};
test_output[32616:32623] = '{32'h426819a9, 32'h415ea2be, 32'h4223e848, 32'h42371fc2, 32'h0, 32'h42aabcef, 32'h4221f713, 32'h0};
test_input[32624:32631] = '{32'h42c1cc07, 32'h41af3d67, 32'hc274be9f, 32'hc2b8c9b4, 32'h42bdc860, 32'h428f24ce, 32'h4296151f, 32'hc2bba22d};
test_output[32624:32631] = '{32'h42c1cc07, 32'h41af3d67, 32'h0, 32'h0, 32'h42bdc860, 32'h428f24ce, 32'h4296151f, 32'h0};
test_input[32632:32639] = '{32'h423085f0, 32'hc291226e, 32'hc282c6e5, 32'hbf7d83e3, 32'h42bb5765, 32'h42347436, 32'h4273d6a3, 32'h42216cc3};
test_output[32632:32639] = '{32'h423085f0, 32'h0, 32'h0, 32'h0, 32'h42bb5765, 32'h42347436, 32'h4273d6a3, 32'h42216cc3};
test_input[32640:32647] = '{32'hc12c70cf, 32'hc25dc004, 32'h42b66f5d, 32'hc1faf198, 32'hc21a43c3, 32'h420d32e6, 32'h42c567e1, 32'h41f6ee28};
test_output[32640:32647] = '{32'h0, 32'h0, 32'h42b66f5d, 32'h0, 32'h0, 32'h420d32e6, 32'h42c567e1, 32'h41f6ee28};
test_input[32648:32655] = '{32'hc2a9611e, 32'h42a9f28d, 32'h4170b142, 32'hc297fe23, 32'h41db87fd, 32'h4206657d, 32'hc20d90c6, 32'h42b60891};
test_output[32648:32655] = '{32'h0, 32'h42a9f28d, 32'h4170b142, 32'h0, 32'h41db87fd, 32'h4206657d, 32'h0, 32'h42b60891};
test_input[32656:32663] = '{32'h42700c63, 32'h4225e9a2, 32'hc2432c18, 32'h4294f612, 32'hc29e3287, 32'hc1c18331, 32'h42710be4, 32'h42615bfe};
test_output[32656:32663] = '{32'h42700c63, 32'h4225e9a2, 32'h0, 32'h4294f612, 32'h0, 32'h0, 32'h42710be4, 32'h42615bfe};
test_input[32664:32671] = '{32'hc29b3057, 32'h41c6287e, 32'hc23bfa1e, 32'hc28b8cfc, 32'hc2c6d32a, 32'h41e9b097, 32'h41b09582, 32'h40bcc986};
test_output[32664:32671] = '{32'h0, 32'h41c6287e, 32'h0, 32'h0, 32'h0, 32'h41e9b097, 32'h41b09582, 32'h40bcc986};
test_input[32672:32679] = '{32'hc2a4d8be, 32'hc2a7c0e2, 32'hc1db0a84, 32'h41f62023, 32'h40f959ea, 32'h41cf7574, 32'hc22f5939, 32'hc29ce7fe};
test_output[32672:32679] = '{32'h0, 32'h0, 32'h0, 32'h41f62023, 32'h40f959ea, 32'h41cf7574, 32'h0, 32'h0};
test_input[32680:32687] = '{32'h429bac32, 32'h41ce0d7a, 32'h422d137b, 32'h419e22d7, 32'h42392819, 32'hc2b2575f, 32'h42104b8f, 32'hc2be5109};
test_output[32680:32687] = '{32'h429bac32, 32'h41ce0d7a, 32'h422d137b, 32'h419e22d7, 32'h42392819, 32'h0, 32'h42104b8f, 32'h0};
test_input[32688:32695] = '{32'h42302209, 32'h42856132, 32'hc2aecdf2, 32'h4255a6cb, 32'hc19f6ad9, 32'h42348dbb, 32'h4211f952, 32'hc2b7d147};
test_output[32688:32695] = '{32'h42302209, 32'h42856132, 32'h0, 32'h4255a6cb, 32'h0, 32'h42348dbb, 32'h4211f952, 32'h0};
test_input[32696:32703] = '{32'h42b201c8, 32'hc2b7acb8, 32'hc28a9932, 32'h41b648c0, 32'hc17c00de, 32'hc0dddbb1, 32'h41ef6007, 32'hc1a3b3fc};
test_output[32696:32703] = '{32'h42b201c8, 32'h0, 32'h0, 32'h41b648c0, 32'h0, 32'h0, 32'h41ef6007, 32'h0};
test_input[32704:32711] = '{32'h41de1262, 32'hc0c675ad, 32'hc2990d71, 32'hc0a8cae0, 32'h424d1ebc, 32'hc2b1a60d, 32'h425bee0b, 32'hc2b3aeb7};
test_output[32704:32711] = '{32'h41de1262, 32'h0, 32'h0, 32'h0, 32'h424d1ebc, 32'h0, 32'h425bee0b, 32'h0};
test_input[32712:32719] = '{32'h428135f0, 32'hc1927997, 32'hc24abc62, 32'hc2007d7b, 32'h4276ca64, 32'h41f42fcd, 32'hc181023c, 32'hc288879c};
test_output[32712:32719] = '{32'h428135f0, 32'h0, 32'h0, 32'h0, 32'h4276ca64, 32'h41f42fcd, 32'h0, 32'h0};
test_input[32720:32727] = '{32'h41e29a45, 32'hbfdbc1b4, 32'hc2c64b59, 32'hc1db2cd2, 32'hc26f0b3d, 32'h423d7169, 32'h415e76b7, 32'hc2b4cbbd};
test_output[32720:32727] = '{32'h41e29a45, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423d7169, 32'h415e76b7, 32'h0};
test_input[32728:32735] = '{32'h41f50cbe, 32'hc17d6987, 32'h4295fbb3, 32'hc2c360d9, 32'h42897e21, 32'hc191ec72, 32'hc1302c4c, 32'h42647f2b};
test_output[32728:32735] = '{32'h41f50cbe, 32'h0, 32'h4295fbb3, 32'h0, 32'h42897e21, 32'h0, 32'h0, 32'h42647f2b};
test_input[32736:32743] = '{32'h41dc3361, 32'hc2b447a1, 32'hc25db623, 32'hc2a55a5f, 32'h425bb928, 32'h402d1e76, 32'h42b2d49d, 32'h42825070};
test_output[32736:32743] = '{32'h41dc3361, 32'h0, 32'h0, 32'h0, 32'h425bb928, 32'h402d1e76, 32'h42b2d49d, 32'h42825070};
test_input[32744:32751] = '{32'hc0fd1e92, 32'hc2c018f5, 32'h41a55cc3, 32'hc243dcff, 32'hc2bc1856, 32'hc0c6dcb7, 32'h426f5944, 32'hc2842a85};
test_output[32744:32751] = '{32'h0, 32'h0, 32'h41a55cc3, 32'h0, 32'h0, 32'h0, 32'h426f5944, 32'h0};
test_input[32752:32759] = '{32'hc259d3e0, 32'hc241968d, 32'hc0927864, 32'h41dd3898, 32'hc2c21ff6, 32'h41fa6568, 32'h419fd264, 32'hc173ad48};
test_output[32752:32759] = '{32'h0, 32'h0, 32'h0, 32'h41dd3898, 32'h0, 32'h41fa6568, 32'h419fd264, 32'h0};
test_input[32760:32767] = '{32'hc2965dcf, 32'hc2842ad0, 32'h41ac24d0, 32'h41b51402, 32'h408e6346, 32'h42181135, 32'hc0a70b71, 32'hc209a964};
test_output[32760:32767] = '{32'h0, 32'h0, 32'h41ac24d0, 32'h41b51402, 32'h408e6346, 32'h42181135, 32'h0, 32'h0};
test_input[32768:32775] = '{32'h4228384b, 32'h402797f4, 32'hc266b9b9, 32'hc260c229, 32'hc1c7e1b2, 32'hc2a0bb21, 32'h421b206e, 32'h42802344};
test_output[32768:32775] = '{32'h4228384b, 32'h402797f4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h421b206e, 32'h42802344};
test_input[32776:32783] = '{32'hc25aaee8, 32'hc12d5a14, 32'hc27eb9eb, 32'hc2afb05a, 32'hc1e1484f, 32'hc179c103, 32'hc2c624a8, 32'hc214801d};
test_output[32776:32783] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[32784:32791] = '{32'h41af5d35, 32'h42c39e9a, 32'hc2a5b745, 32'h42999c21, 32'h422540f6, 32'hc2c0fa0a, 32'hc28f3c08, 32'hc2bcddf0};
test_output[32784:32791] = '{32'h41af5d35, 32'h42c39e9a, 32'h0, 32'h42999c21, 32'h422540f6, 32'h0, 32'h0, 32'h0};
test_input[32792:32799] = '{32'h4299af66, 32'hc1e17d85, 32'hc05aff4b, 32'h42ab04c5, 32'hc2468a7d, 32'hc2042315, 32'h3f86630c, 32'h425a866e};
test_output[32792:32799] = '{32'h4299af66, 32'h0, 32'h0, 32'h42ab04c5, 32'h0, 32'h0, 32'h3f86630c, 32'h425a866e};
test_input[32800:32807] = '{32'h412cfc45, 32'h4264da37, 32'hc26bb93a, 32'hc26466ca, 32'hc20c6c77, 32'h420e31be, 32'h424f3976, 32'hc2009a24};
test_output[32800:32807] = '{32'h412cfc45, 32'h4264da37, 32'h0, 32'h0, 32'h0, 32'h420e31be, 32'h424f3976, 32'h0};
test_input[32808:32815] = '{32'h42b6b93c, 32'hc1d4dffb, 32'hc278ba47, 32'hc29ad22e, 32'hc2a8cb29, 32'hc2b79561, 32'h41740419, 32'hc1e38ce6};
test_output[32808:32815] = '{32'h42b6b93c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41740419, 32'h0};
test_input[32816:32823] = '{32'h4293d250, 32'h42ab217f, 32'h423b708e, 32'hc2c73247, 32'hc251c553, 32'hc1d817dd, 32'h4084e461, 32'hc22673e2};
test_output[32816:32823] = '{32'h4293d250, 32'h42ab217f, 32'h423b708e, 32'h0, 32'h0, 32'h0, 32'h4084e461, 32'h0};
test_input[32824:32831] = '{32'h422035aa, 32'h40aea5d4, 32'h411b9a7b, 32'hc2aeed46, 32'h421f88ef, 32'hc25a1f5e, 32'hc28b304b, 32'hc2b2aed4};
test_output[32824:32831] = '{32'h422035aa, 32'h40aea5d4, 32'h411b9a7b, 32'h0, 32'h421f88ef, 32'h0, 32'h0, 32'h0};
test_input[32832:32839] = '{32'hc2012652, 32'hc28760f5, 32'hbf94e284, 32'hc2a3fbcd, 32'hc21af0c8, 32'hc2331177, 32'hc2b64494, 32'h419b2e99};
test_output[32832:32839] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h419b2e99};
test_input[32840:32847] = '{32'h4240c190, 32'hc2c0eb83, 32'h42b3c55f, 32'hc2652754, 32'hc28fc579, 32'hc2c6e7fa, 32'hc101f8a3, 32'h4237b7be};
test_output[32840:32847] = '{32'h4240c190, 32'h0, 32'h42b3c55f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4237b7be};
test_input[32848:32855] = '{32'h42b79925, 32'hc2a28586, 32'hc1dd3ded, 32'h429a27a1, 32'h42a2132a, 32'hc28739fe, 32'h426acf91, 32'hc12d75c2};
test_output[32848:32855] = '{32'h42b79925, 32'h0, 32'h0, 32'h429a27a1, 32'h42a2132a, 32'h0, 32'h426acf91, 32'h0};
test_input[32856:32863] = '{32'h42362646, 32'h42bf96e1, 32'h424560a4, 32'hc28036a5, 32'h41ef4bf0, 32'hc2016208, 32'h423f3376, 32'hc28721d6};
test_output[32856:32863] = '{32'h42362646, 32'h42bf96e1, 32'h424560a4, 32'h0, 32'h41ef4bf0, 32'h0, 32'h423f3376, 32'h0};
test_input[32864:32871] = '{32'h4290b2b1, 32'h41e4bddb, 32'hc15034e7, 32'h419404a5, 32'h41c14a84, 32'hc29dff8b, 32'h4142173a, 32'h42bfa9d8};
test_output[32864:32871] = '{32'h4290b2b1, 32'h41e4bddb, 32'h0, 32'h419404a5, 32'h41c14a84, 32'h0, 32'h4142173a, 32'h42bfa9d8};
test_input[32872:32879] = '{32'hc2817958, 32'hc2ae4f68, 32'hc2829729, 32'hc2b2348a, 32'h42ae28ba, 32'hc17a91d8, 32'h42b15613, 32'h429318c4};
test_output[32872:32879] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42ae28ba, 32'h0, 32'h42b15613, 32'h429318c4};
test_input[32880:32887] = '{32'hbf7addb7, 32'h42400e1f, 32'h42155ddc, 32'hc2757b51, 32'hc1f67166, 32'hc29cc086, 32'hc2bff9f6, 32'hc1dc5cee};
test_output[32880:32887] = '{32'h0, 32'h42400e1f, 32'h42155ddc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[32888:32895] = '{32'h41ad00ed, 32'h42253cca, 32'h414300b3, 32'h42aef24c, 32'hc148bc48, 32'h40e31cad, 32'h42804cfc, 32'h426136f1};
test_output[32888:32895] = '{32'h41ad00ed, 32'h42253cca, 32'h414300b3, 32'h42aef24c, 32'h0, 32'h40e31cad, 32'h42804cfc, 32'h426136f1};
test_input[32896:32903] = '{32'h40f57333, 32'hc169fc38, 32'hc1564319, 32'hc2a98986, 32'h423bc59c, 32'h42ae7237, 32'h423a57d1, 32'h4216325d};
test_output[32896:32903] = '{32'h40f57333, 32'h0, 32'h0, 32'h0, 32'h423bc59c, 32'h42ae7237, 32'h423a57d1, 32'h4216325d};
test_input[32904:32911] = '{32'hc2ba07c6, 32'hc21e48d0, 32'hc2a6948a, 32'hc05bb243, 32'hc2a126fc, 32'h42b74aab, 32'hc27fe48c, 32'hc2a03b8b};
test_output[32904:32911] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b74aab, 32'h0, 32'h0};
test_input[32912:32919] = '{32'hc2b6cc7a, 32'h42b7996e, 32'h414d778d, 32'hc200ad46, 32'hc27a3dec, 32'hc1c8fe66, 32'hc2aaef69, 32'h42bda08b};
test_output[32912:32919] = '{32'h0, 32'h42b7996e, 32'h414d778d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bda08b};
test_input[32920:32927] = '{32'h4278c44c, 32'hc1e23ef2, 32'hc271f13a, 32'hc03b0622, 32'h41ba2f92, 32'h4140b131, 32'h4213e419, 32'hc282f605};
test_output[32920:32927] = '{32'h4278c44c, 32'h0, 32'h0, 32'h0, 32'h41ba2f92, 32'h4140b131, 32'h4213e419, 32'h0};
test_input[32928:32935] = '{32'hc24329d0, 32'hc0cdf48b, 32'h42879c65, 32'hc1ef31a4, 32'h423ea49e, 32'hc2c1c187, 32'h42af86f3, 32'hc00af95d};
test_output[32928:32935] = '{32'h0, 32'h0, 32'h42879c65, 32'h0, 32'h423ea49e, 32'h0, 32'h42af86f3, 32'h0};
test_input[32936:32943] = '{32'h41f6bc39, 32'h40914531, 32'hc2ae37fc, 32'h41c7f8e3, 32'h411c0d11, 32'h41a7878f, 32'hc28f411f, 32'hc28d5e87};
test_output[32936:32943] = '{32'h41f6bc39, 32'h40914531, 32'h0, 32'h41c7f8e3, 32'h411c0d11, 32'h41a7878f, 32'h0, 32'h0};
test_input[32944:32951] = '{32'hc254a5d6, 32'hc1a280a4, 32'h42b32bc4, 32'h4273775a, 32'h42935127, 32'hc024573b, 32'hc181bec1, 32'h420f877e};
test_output[32944:32951] = '{32'h0, 32'h0, 32'h42b32bc4, 32'h4273775a, 32'h42935127, 32'h0, 32'h0, 32'h420f877e};
test_input[32952:32959] = '{32'h41eb263a, 32'hc240ce22, 32'hc22be0e3, 32'hc2755475, 32'hc1bcb776, 32'h42bb3bef, 32'h42a30e0b, 32'hc1510f99};
test_output[32952:32959] = '{32'h41eb263a, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bb3bef, 32'h42a30e0b, 32'h0};
test_input[32960:32967] = '{32'hc25cf11c, 32'h42a37906, 32'h4296bd25, 32'h416a9258, 32'h41e9447b, 32'h420bd29a, 32'h42c483a8, 32'hc2107f78};
test_output[32960:32967] = '{32'h0, 32'h42a37906, 32'h4296bd25, 32'h416a9258, 32'h41e9447b, 32'h420bd29a, 32'h42c483a8, 32'h0};
test_input[32968:32975] = '{32'h42b8b326, 32'h41701733, 32'hc08fa7c6, 32'hc2a55faf, 32'h40c92a88, 32'hc2551c97, 32'h423c919e, 32'h42b3c1aa};
test_output[32968:32975] = '{32'h42b8b326, 32'h41701733, 32'h0, 32'h0, 32'h40c92a88, 32'h0, 32'h423c919e, 32'h42b3c1aa};
test_input[32976:32983] = '{32'h4256160f, 32'h4175abee, 32'hc29a0004, 32'h41ba7fc0, 32'h3f023bfc, 32'hc1fdfcea, 32'hc2461f4d, 32'hc1259459};
test_output[32976:32983] = '{32'h4256160f, 32'h4175abee, 32'h0, 32'h41ba7fc0, 32'h3f023bfc, 32'h0, 32'h0, 32'h0};
test_input[32984:32991] = '{32'hc2959784, 32'h41e439c5, 32'hc105c7af, 32'hc2043f6f, 32'h42606cd6, 32'h42a251da, 32'hc1a6808b, 32'h41997a1d};
test_output[32984:32991] = '{32'h0, 32'h41e439c5, 32'h0, 32'h0, 32'h42606cd6, 32'h42a251da, 32'h0, 32'h41997a1d};
test_input[32992:32999] = '{32'h41266c0d, 32'h41d9feb4, 32'h42bc0777, 32'h42a4cdab, 32'hc2bd83d5, 32'h418eda82, 32'h429d5970, 32'h42549034};
test_output[32992:32999] = '{32'h41266c0d, 32'h41d9feb4, 32'h42bc0777, 32'h42a4cdab, 32'h0, 32'h418eda82, 32'h429d5970, 32'h42549034};
test_input[33000:33007] = '{32'hc28e0911, 32'hc2967be7, 32'hc25de65d, 32'hc1f1baf6, 32'hc213314f, 32'h4290c0fd, 32'hc271d6ae, 32'h427d4fe1};
test_output[33000:33007] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4290c0fd, 32'h0, 32'h427d4fe1};
test_input[33008:33015] = '{32'h4251a9bc, 32'h41cd22c8, 32'hc2583571, 32'h419924cf, 32'h41b7234d, 32'hc27f7ec3, 32'hc2a87c25, 32'h418c42d8};
test_output[33008:33015] = '{32'h4251a9bc, 32'h41cd22c8, 32'h0, 32'h419924cf, 32'h41b7234d, 32'h0, 32'h0, 32'h418c42d8};
test_input[33016:33023] = '{32'h421763dc, 32'hc1471ba7, 32'hc2747249, 32'hc0e83e08, 32'hc22486aa, 32'hc1a25f81, 32'h4272306f, 32'h41b67eba};
test_output[33016:33023] = '{32'h421763dc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4272306f, 32'h41b67eba};
test_input[33024:33031] = '{32'h3fbeba11, 32'hc271c24f, 32'hc2c37d63, 32'hc2611996, 32'h42aaa6eb, 32'h423da180, 32'h42bb5c18, 32'hc2a2a400};
test_output[33024:33031] = '{32'h3fbeba11, 32'h0, 32'h0, 32'h0, 32'h42aaa6eb, 32'h423da180, 32'h42bb5c18, 32'h0};
test_input[33032:33039] = '{32'hc209b0ed, 32'h4246f0e7, 32'h42a8b5bf, 32'hc15f95d4, 32'h428b9660, 32'h42302385, 32'h419fb44c, 32'h42739fad};
test_output[33032:33039] = '{32'h0, 32'h4246f0e7, 32'h42a8b5bf, 32'h0, 32'h428b9660, 32'h42302385, 32'h419fb44c, 32'h42739fad};
test_input[33040:33047] = '{32'hc20d22c7, 32'hc098757b, 32'h42b07909, 32'hc187c3c1, 32'hc2028f5d, 32'h42b8547c, 32'h41d14937, 32'h42119c8e};
test_output[33040:33047] = '{32'h0, 32'h0, 32'h42b07909, 32'h0, 32'h0, 32'h42b8547c, 32'h41d14937, 32'h42119c8e};
test_input[33048:33055] = '{32'hc298796a, 32'h41a5f979, 32'h422ac154, 32'hc2bef1c0, 32'hc2c76dfe, 32'hc2056bbf, 32'h42a2c08f, 32'h42219a34};
test_output[33048:33055] = '{32'h0, 32'h41a5f979, 32'h422ac154, 32'h0, 32'h0, 32'h0, 32'h42a2c08f, 32'h42219a34};
test_input[33056:33063] = '{32'h42a8ab1b, 32'hc165813f, 32'h4248f866, 32'h42342c35, 32'h4234acfb, 32'hc1f1e630, 32'hc25d1c33, 32'hc2a9b427};
test_output[33056:33063] = '{32'h42a8ab1b, 32'h0, 32'h4248f866, 32'h42342c35, 32'h4234acfb, 32'h0, 32'h0, 32'h0};
test_input[33064:33071] = '{32'h424d46f6, 32'h412398ca, 32'h41b24eeb, 32'hc219a048, 32'hc2695dd7, 32'hc2c4cfa2, 32'h414700ec, 32'hc22894ce};
test_output[33064:33071] = '{32'h424d46f6, 32'h412398ca, 32'h41b24eeb, 32'h0, 32'h0, 32'h0, 32'h414700ec, 32'h0};
test_input[33072:33079] = '{32'h4252c3d4, 32'hc2765d95, 32'h41deb689, 32'hc2a5613c, 32'hc21bb3ab, 32'h42696940, 32'hc0b78822, 32'hc1a2d6c6};
test_output[33072:33079] = '{32'h4252c3d4, 32'h0, 32'h41deb689, 32'h0, 32'h0, 32'h42696940, 32'h0, 32'h0};
test_input[33080:33087] = '{32'hc2984560, 32'hc133dab3, 32'hc17046a8, 32'h423bad91, 32'h41e4daf4, 32'h41486bf2, 32'hc275223d, 32'h42c6fabe};
test_output[33080:33087] = '{32'h0, 32'h0, 32'h0, 32'h423bad91, 32'h41e4daf4, 32'h41486bf2, 32'h0, 32'h42c6fabe};
test_input[33088:33095] = '{32'hc16a8185, 32'h42a44132, 32'hc20825df, 32'hc1cd3364, 32'hc14afe5f, 32'hc146ee5f, 32'h4293c41f, 32'h404f5c18};
test_output[33088:33095] = '{32'h0, 32'h42a44132, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4293c41f, 32'h404f5c18};
test_input[33096:33103] = '{32'hc270235c, 32'h4218b0f2, 32'h42c78644, 32'hc1bdd536, 32'h4270a4bf, 32'hc12a0cbb, 32'hc1124ab3, 32'h423213f0};
test_output[33096:33103] = '{32'h0, 32'h4218b0f2, 32'h42c78644, 32'h0, 32'h4270a4bf, 32'h0, 32'h0, 32'h423213f0};
test_input[33104:33111] = '{32'h4088d82d, 32'h41cf1d71, 32'hc1df8c09, 32'h42496ede, 32'h426ab07b, 32'hc29eeba8, 32'hc291b230, 32'hc2836adc};
test_output[33104:33111] = '{32'h4088d82d, 32'h41cf1d71, 32'h0, 32'h42496ede, 32'h426ab07b, 32'h0, 32'h0, 32'h0};
test_input[33112:33119] = '{32'hc1e0777f, 32'h42b967a8, 32'hc19480ec, 32'hc1e287b2, 32'hc29c5608, 32'h4031a20a, 32'hc22276f3, 32'hc2970f8e};
test_output[33112:33119] = '{32'h0, 32'h42b967a8, 32'h0, 32'h0, 32'h0, 32'h4031a20a, 32'h0, 32'h0};
test_input[33120:33127] = '{32'hc2a81a8c, 32'h429db3cc, 32'h41c475ee, 32'hc2abc614, 32'h4243104d, 32'hc1a25478, 32'hc2c4e0fa, 32'h42224683};
test_output[33120:33127] = '{32'h0, 32'h429db3cc, 32'h41c475ee, 32'h0, 32'h4243104d, 32'h0, 32'h0, 32'h42224683};
test_input[33128:33135] = '{32'hc2678fb6, 32'hc2b61e4d, 32'h41d861e8, 32'h42a2eed3, 32'h428a0c97, 32'h4287ca21, 32'h42b906db, 32'h4266f8df};
test_output[33128:33135] = '{32'h0, 32'h0, 32'h41d861e8, 32'h42a2eed3, 32'h428a0c97, 32'h4287ca21, 32'h42b906db, 32'h4266f8df};
test_input[33136:33143] = '{32'hc269432d, 32'h41558366, 32'h41c209a5, 32'hc28186a6, 32'h4239dc43, 32'hc2942b97, 32'hc25d14ea, 32'hc208de42};
test_output[33136:33143] = '{32'h0, 32'h41558366, 32'h41c209a5, 32'h0, 32'h4239dc43, 32'h0, 32'h0, 32'h0};
test_input[33144:33151] = '{32'hc22e9e68, 32'h42085438, 32'h426d8215, 32'hc2bea2e6, 32'hc1778ca5, 32'hc1edc728, 32'hc167fda9, 32'hc12f393d};
test_output[33144:33151] = '{32'h0, 32'h42085438, 32'h426d8215, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[33152:33159] = '{32'hc217b5db, 32'hc2465324, 32'h424318a5, 32'h41938774, 32'hc0cffcd3, 32'hc2a21c66, 32'h42607c77, 32'hc2c2384b};
test_output[33152:33159] = '{32'h0, 32'h0, 32'h424318a5, 32'h41938774, 32'h0, 32'h0, 32'h42607c77, 32'h0};
test_input[33160:33167] = '{32'h4209b455, 32'h429e9699, 32'h427cb37c, 32'hc0744de1, 32'hc2c2b22c, 32'hc10425d1, 32'h42bf76c7, 32'hc2bebecc};
test_output[33160:33167] = '{32'h4209b455, 32'h429e9699, 32'h427cb37c, 32'h0, 32'h0, 32'h0, 32'h42bf76c7, 32'h0};
test_input[33168:33175] = '{32'h422eefdd, 32'hc26abc6e, 32'hbf16db5e, 32'hc29cd867, 32'h4256a347, 32'hc2a8bd38, 32'h4205895b, 32'hc2b14b26};
test_output[33168:33175] = '{32'h422eefdd, 32'h0, 32'h0, 32'h0, 32'h4256a347, 32'h0, 32'h4205895b, 32'h0};
test_input[33176:33183] = '{32'hc27bfb37, 32'h42bdd48d, 32'h42037d35, 32'h41ebc194, 32'h417b216a, 32'hc2c6dc7b, 32'hc285b3f0, 32'h41418408};
test_output[33176:33183] = '{32'h0, 32'h42bdd48d, 32'h42037d35, 32'h41ebc194, 32'h417b216a, 32'h0, 32'h0, 32'h41418408};
test_input[33184:33191] = '{32'h429c77c2, 32'hc05d0a46, 32'h42c47da5, 32'h41e8d13e, 32'h41eb9b57, 32'hc25900ad, 32'h428f2005, 32'hc2285c4a};
test_output[33184:33191] = '{32'h429c77c2, 32'h0, 32'h42c47da5, 32'h41e8d13e, 32'h41eb9b57, 32'h0, 32'h428f2005, 32'h0};
test_input[33192:33199] = '{32'h41fcd3e6, 32'hc2baf17b, 32'h42840c85, 32'hc1b48e0f, 32'hc2382ae4, 32'h422351a8, 32'h423f7d75, 32'hc10e471c};
test_output[33192:33199] = '{32'h41fcd3e6, 32'h0, 32'h42840c85, 32'h0, 32'h0, 32'h422351a8, 32'h423f7d75, 32'h0};
test_input[33200:33207] = '{32'hc20abaa1, 32'h425bc701, 32'h42940491, 32'hc281bf22, 32'h42b25b96, 32'hc13ca4f7, 32'hc212e178, 32'h4236ca45};
test_output[33200:33207] = '{32'h0, 32'h425bc701, 32'h42940491, 32'h0, 32'h42b25b96, 32'h0, 32'h0, 32'h4236ca45};
test_input[33208:33215] = '{32'hc2649501, 32'h4282bc9e, 32'hc2b3a9c9, 32'hc271d74c, 32'h3f77041b, 32'h4284e482, 32'hc1849028, 32'h421100a5};
test_output[33208:33215] = '{32'h0, 32'h4282bc9e, 32'h0, 32'h0, 32'h3f77041b, 32'h4284e482, 32'h0, 32'h421100a5};
test_input[33216:33223] = '{32'h4112c4d4, 32'hc0d6c581, 32'h42094b54, 32'hc2094a75, 32'h416272ec, 32'hc29d36a7, 32'h410b73ad, 32'hc17e693a};
test_output[33216:33223] = '{32'h4112c4d4, 32'h0, 32'h42094b54, 32'h0, 32'h416272ec, 32'h0, 32'h410b73ad, 32'h0};
test_input[33224:33231] = '{32'h42810ca0, 32'h42ba3172, 32'hc22c5fe1, 32'h416f27cd, 32'hc18e1c7d, 32'h421b190e, 32'h421876ff, 32'hc2779ab2};
test_output[33224:33231] = '{32'h42810ca0, 32'h42ba3172, 32'h0, 32'h416f27cd, 32'h0, 32'h421b190e, 32'h421876ff, 32'h0};
test_input[33232:33239] = '{32'h416249f8, 32'h401c8d6e, 32'hc2a11492, 32'hc195a3d7, 32'hc222cdf6, 32'hc0f35b87, 32'hc0cf26b2, 32'h4169a412};
test_output[33232:33239] = '{32'h416249f8, 32'h401c8d6e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4169a412};
test_input[33240:33247] = '{32'hc28a6bf9, 32'h42c3c8b9, 32'hc2ad3bde, 32'h423ec7b2, 32'h42b28df1, 32'h4232edd5, 32'hc2b2e53c, 32'hc2c4235d};
test_output[33240:33247] = '{32'h0, 32'h42c3c8b9, 32'h0, 32'h423ec7b2, 32'h42b28df1, 32'h4232edd5, 32'h0, 32'h0};
test_input[33248:33255] = '{32'h426b63e1, 32'hc22fffad, 32'h42111f69, 32'hc28c7036, 32'hc27a2518, 32'hc2b75335, 32'hc23b1ed8, 32'h42c4e201};
test_output[33248:33255] = '{32'h426b63e1, 32'h0, 32'h42111f69, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c4e201};
test_input[33256:33263] = '{32'h42451c38, 32'h4287dcad, 32'h42803b27, 32'h41a8b32f, 32'hc27a3194, 32'h424c7c62, 32'h42282da3, 32'hc15f6274};
test_output[33256:33263] = '{32'h42451c38, 32'h4287dcad, 32'h42803b27, 32'h41a8b32f, 32'h0, 32'h424c7c62, 32'h42282da3, 32'h0};
test_input[33264:33271] = '{32'hc2b3fd5c, 32'h41b0673b, 32'hc257c779, 32'h4187e2ce, 32'h423a9bba, 32'hc2832433, 32'h420e20e5, 32'hc20350be};
test_output[33264:33271] = '{32'h0, 32'h41b0673b, 32'h0, 32'h4187e2ce, 32'h423a9bba, 32'h0, 32'h420e20e5, 32'h0};
test_input[33272:33279] = '{32'hc2a9b487, 32'hc2b71d73, 32'h42c53dcd, 32'hc2b07346, 32'hc2406291, 32'h417c2b99, 32'hc2763d16, 32'h426cd3fa};
test_output[33272:33279] = '{32'h0, 32'h0, 32'h42c53dcd, 32'h0, 32'h0, 32'h417c2b99, 32'h0, 32'h426cd3fa};
test_input[33280:33287] = '{32'h428ffe0f, 32'hc25b7d19, 32'hc1c67b4f, 32'h3fcdad51, 32'hc201a4e5, 32'h42005d04, 32'h42b53e58, 32'hc1980ba6};
test_output[33280:33287] = '{32'h428ffe0f, 32'h0, 32'h0, 32'h3fcdad51, 32'h0, 32'h42005d04, 32'h42b53e58, 32'h0};
test_input[33288:33295] = '{32'hc2ae7c11, 32'hc20ffb5e, 32'h425f5a80, 32'hc1c96e6e, 32'h40b7417e, 32'h42238fa6, 32'h4290b2be, 32'hc2881977};
test_output[33288:33295] = '{32'h0, 32'h0, 32'h425f5a80, 32'h0, 32'h40b7417e, 32'h42238fa6, 32'h4290b2be, 32'h0};
test_input[33296:33303] = '{32'h41a22f67, 32'hc2b56d7c, 32'h41d99378, 32'hc2b1a88d, 32'h42bf49bd, 32'hc246b8ac, 32'hc0e94edc, 32'hc282e773};
test_output[33296:33303] = '{32'h41a22f67, 32'h0, 32'h41d99378, 32'h0, 32'h42bf49bd, 32'h0, 32'h0, 32'h0};
test_input[33304:33311] = '{32'hc2474689, 32'hc2b29c48, 32'h41cc644c, 32'h42144da6, 32'h418564f7, 32'hc2059594, 32'h4234e7a6, 32'hc2bac5b2};
test_output[33304:33311] = '{32'h0, 32'h0, 32'h41cc644c, 32'h42144da6, 32'h418564f7, 32'h0, 32'h4234e7a6, 32'h0};
test_input[33312:33319] = '{32'h42c36d4f, 32'h423c2537, 32'hc2702fb6, 32'h42448792, 32'h410e7282, 32'h4292b6cd, 32'hc232fe21, 32'hc2a9d603};
test_output[33312:33319] = '{32'h42c36d4f, 32'h423c2537, 32'h0, 32'h42448792, 32'h410e7282, 32'h4292b6cd, 32'h0, 32'h0};
test_input[33320:33327] = '{32'h427fb80f, 32'h40ce45e3, 32'hc26458f5, 32'h42ace0f9, 32'hc13e574d, 32'h42b78a4c, 32'hc206816a, 32'hc246cb8a};
test_output[33320:33327] = '{32'h427fb80f, 32'h40ce45e3, 32'h0, 32'h42ace0f9, 32'h0, 32'h42b78a4c, 32'h0, 32'h0};
test_input[33328:33335] = '{32'hc1c67114, 32'hc2a9e7fe, 32'h41ef0eb7, 32'h427dd001, 32'h42821836, 32'hc251eb62, 32'hc206ee89, 32'h420c140e};
test_output[33328:33335] = '{32'h0, 32'h0, 32'h41ef0eb7, 32'h427dd001, 32'h42821836, 32'h0, 32'h0, 32'h420c140e};
test_input[33336:33343] = '{32'h41ac621d, 32'hc14dbfd3, 32'h429ebd61, 32'hc269fa18, 32'hc293b7cd, 32'h4138d74b, 32'hc2641a01, 32'hc26551f7};
test_output[33336:33343] = '{32'h41ac621d, 32'h0, 32'h429ebd61, 32'h0, 32'h0, 32'h4138d74b, 32'h0, 32'h0};
test_input[33344:33351] = '{32'h426a6a19, 32'hc244eb0a, 32'h4198481b, 32'hc13d70cc, 32'hc184c133, 32'hc111edc0, 32'hc18ba26f, 32'hc28c8e8f};
test_output[33344:33351] = '{32'h426a6a19, 32'h0, 32'h4198481b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[33352:33359] = '{32'h425d71f1, 32'h42557ed1, 32'h41b1c0dd, 32'h41f71938, 32'hc2aeae8f, 32'h414bcbd6, 32'hc23249d9, 32'hc2bce028};
test_output[33352:33359] = '{32'h425d71f1, 32'h42557ed1, 32'h41b1c0dd, 32'h41f71938, 32'h0, 32'h414bcbd6, 32'h0, 32'h0};
test_input[33360:33367] = '{32'hc281fadd, 32'hc1d13161, 32'h402cf848, 32'hc26e4b06, 32'h42c19855, 32'hc294c3e4, 32'hc18e7bf9, 32'h424efb60};
test_output[33360:33367] = '{32'h0, 32'h0, 32'h402cf848, 32'h0, 32'h42c19855, 32'h0, 32'h0, 32'h424efb60};
test_input[33368:33375] = '{32'h42a7bb9e, 32'hc2c622c6, 32'h42a20f8d, 32'h4232ba8a, 32'h40e5ece5, 32'hc248a62b, 32'hc08a9cff, 32'h4231e85a};
test_output[33368:33375] = '{32'h42a7bb9e, 32'h0, 32'h42a20f8d, 32'h4232ba8a, 32'h40e5ece5, 32'h0, 32'h0, 32'h4231e85a};
test_input[33376:33383] = '{32'hc1edc7aa, 32'h4221ecf8, 32'hc27aea7b, 32'h420e1918, 32'h420fe1ca, 32'hc1bdf7c4, 32'h42c46da9, 32'hc26e169a};
test_output[33376:33383] = '{32'h0, 32'h4221ecf8, 32'h0, 32'h420e1918, 32'h420fe1ca, 32'h0, 32'h42c46da9, 32'h0};
test_input[33384:33391] = '{32'h429aaccf, 32'hc20fd7e0, 32'h41e870ed, 32'h41e845c6, 32'h4159bdec, 32'hc1c6e58c, 32'hc23130db, 32'hc19ef5ef};
test_output[33384:33391] = '{32'h429aaccf, 32'h0, 32'h41e870ed, 32'h41e845c6, 32'h4159bdec, 32'h0, 32'h0, 32'h0};
test_input[33392:33399] = '{32'h411f2441, 32'hc2969ebb, 32'h4251a90c, 32'h427e72e9, 32'h42c4454a, 32'hc1781ebe, 32'hc20e78dd, 32'h42915172};
test_output[33392:33399] = '{32'h411f2441, 32'h0, 32'h4251a90c, 32'h427e72e9, 32'h42c4454a, 32'h0, 32'h0, 32'h42915172};
test_input[33400:33407] = '{32'h423fd676, 32'h42a32e07, 32'h41d467aa, 32'h422438b8, 32'hc21045c1, 32'hc1726965, 32'h4266fe3d, 32'hc2147814};
test_output[33400:33407] = '{32'h423fd676, 32'h42a32e07, 32'h41d467aa, 32'h422438b8, 32'h0, 32'h0, 32'h4266fe3d, 32'h0};
test_input[33408:33415] = '{32'hc28766db, 32'hc22f6f8a, 32'hc1e037f3, 32'hc2ac8607, 32'h416fadc1, 32'hc228c0f7, 32'h429ac436, 32'hc211901e};
test_output[33408:33415] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h416fadc1, 32'h0, 32'h429ac436, 32'h0};
test_input[33416:33423] = '{32'hc237406d, 32'h42880c76, 32'h4275d7a7, 32'hc2c5d6ce, 32'hc217ad1f, 32'hc2c25253, 32'h4228fd65, 32'h429dba07};
test_output[33416:33423] = '{32'h0, 32'h42880c76, 32'h4275d7a7, 32'h0, 32'h0, 32'h0, 32'h4228fd65, 32'h429dba07};
test_input[33424:33431] = '{32'hc1981416, 32'hc16df981, 32'h4221db70, 32'h4276ffa8, 32'h4207d80f, 32'h41f6ff4f, 32'h4285ae72, 32'hc1dcd0f3};
test_output[33424:33431] = '{32'h0, 32'h0, 32'h4221db70, 32'h4276ffa8, 32'h4207d80f, 32'h41f6ff4f, 32'h4285ae72, 32'h0};
test_input[33432:33439] = '{32'hc206aa51, 32'hc2488007, 32'hc2a626b5, 32'h40cb46f0, 32'h3c720231, 32'hc1f60921, 32'hc2c70d63, 32'hc15876d1};
test_output[33432:33439] = '{32'h0, 32'h0, 32'h0, 32'h40cb46f0, 32'h3c720231, 32'h0, 32'h0, 32'h0};
test_input[33440:33447] = '{32'hc20d1044, 32'hc1cbfb22, 32'hc1c68a31, 32'hc275667e, 32'hc20f2d04, 32'h42aac1bf, 32'h42bbc970, 32'hc2b57443};
test_output[33440:33447] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42aac1bf, 32'h42bbc970, 32'h0};
test_input[33448:33455] = '{32'hc217d7fa, 32'hc0ba17c9, 32'h41ae5ebc, 32'hc0bbd4e5, 32'h40c67398, 32'h42789f8e, 32'hc2ab7511, 32'hc2a21b95};
test_output[33448:33455] = '{32'h0, 32'h0, 32'h41ae5ebc, 32'h0, 32'h40c67398, 32'h42789f8e, 32'h0, 32'h0};
test_input[33456:33463] = '{32'h41aa82ca, 32'hc28e4592, 32'h41cbfadf, 32'h42375c62, 32'h41afb928, 32'hc1214436, 32'h40823a3e, 32'h42043b11};
test_output[33456:33463] = '{32'h41aa82ca, 32'h0, 32'h41cbfadf, 32'h42375c62, 32'h41afb928, 32'h0, 32'h40823a3e, 32'h42043b11};
test_input[33464:33471] = '{32'hc0995324, 32'h41f96da3, 32'h41f9592d, 32'h42c7755d, 32'h4071eb01, 32'h42aeb105, 32'h42a0fc7a, 32'h42ac1578};
test_output[33464:33471] = '{32'h0, 32'h41f96da3, 32'h41f9592d, 32'h42c7755d, 32'h4071eb01, 32'h42aeb105, 32'h42a0fc7a, 32'h42ac1578};
test_input[33472:33479] = '{32'hc287b5ec, 32'h42962b83, 32'hc2c6923b, 32'h41f8dd47, 32'h424e3890, 32'hc2afa422, 32'hc24d1e39, 32'h412ac8be};
test_output[33472:33479] = '{32'h0, 32'h42962b83, 32'h0, 32'h41f8dd47, 32'h424e3890, 32'h0, 32'h0, 32'h412ac8be};
test_input[33480:33487] = '{32'hc1f0f573, 32'h421de1ad, 32'hc19567d3, 32'hc23f20c2, 32'h41228d27, 32'hc2808fb7, 32'hc14fb839, 32'h428ec158};
test_output[33480:33487] = '{32'h0, 32'h421de1ad, 32'h0, 32'h0, 32'h41228d27, 32'h0, 32'h0, 32'h428ec158};
test_input[33488:33495] = '{32'hc2622d7b, 32'hc1b5a766, 32'h429d8f31, 32'h416cbb68, 32'hc1909806, 32'h40875483, 32'h42850bf7, 32'hc29127c6};
test_output[33488:33495] = '{32'h0, 32'h0, 32'h429d8f31, 32'h416cbb68, 32'h0, 32'h40875483, 32'h42850bf7, 32'h0};
test_input[33496:33503] = '{32'hc204a3ee, 32'hc1945e78, 32'hc23f1dbe, 32'hc22ff827, 32'hc12a14df, 32'h427f13b3, 32'h4296ca1a, 32'hc19de1dd};
test_output[33496:33503] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h427f13b3, 32'h4296ca1a, 32'h0};
test_input[33504:33511] = '{32'h42a96e1e, 32'h41851e91, 32'hc1f65973, 32'h42212f6d, 32'hc2571278, 32'h424185d7, 32'h41d899ef, 32'hc164e7a3};
test_output[33504:33511] = '{32'h42a96e1e, 32'h41851e91, 32'h0, 32'h42212f6d, 32'h0, 32'h424185d7, 32'h41d899ef, 32'h0};
test_input[33512:33519] = '{32'hc1cde598, 32'h42b8dd0e, 32'h42871a58, 32'h41e15228, 32'hc288ea04, 32'h411e4930, 32'h42891b58, 32'hc24c365e};
test_output[33512:33519] = '{32'h0, 32'h42b8dd0e, 32'h42871a58, 32'h41e15228, 32'h0, 32'h411e4930, 32'h42891b58, 32'h0};
test_input[33520:33527] = '{32'h428eea07, 32'h426e541e, 32'hc002c6be, 32'h428f099e, 32'h4241f965, 32'h41b564c5, 32'h42414c7a, 32'hc1d04a97};
test_output[33520:33527] = '{32'h428eea07, 32'h426e541e, 32'h0, 32'h428f099e, 32'h4241f965, 32'h41b564c5, 32'h42414c7a, 32'h0};
test_input[33528:33535] = '{32'h41f0fdc7, 32'h41f6f386, 32'h42a7d2aa, 32'hc2276397, 32'h3fa12f75, 32'hc0ea2d06, 32'h3fe3abd3, 32'h42748f25};
test_output[33528:33535] = '{32'h41f0fdc7, 32'h41f6f386, 32'h42a7d2aa, 32'h0, 32'h3fa12f75, 32'h0, 32'h3fe3abd3, 32'h42748f25};
test_input[33536:33543] = '{32'h423da570, 32'h41641a49, 32'hc234d62f, 32'h41f9c0b6, 32'hc2adcc9e, 32'hc2c4019f, 32'hc22f52e4, 32'h4298e549};
test_output[33536:33543] = '{32'h423da570, 32'h41641a49, 32'h0, 32'h41f9c0b6, 32'h0, 32'h0, 32'h0, 32'h4298e549};
test_input[33544:33551] = '{32'h411b6698, 32'h42c40886, 32'h42871cfb, 32'hc23506f3, 32'h428b5451, 32'h3f43cdf1, 32'hc25166c9, 32'h42b10757};
test_output[33544:33551] = '{32'h411b6698, 32'h42c40886, 32'h42871cfb, 32'h0, 32'h428b5451, 32'h3f43cdf1, 32'h0, 32'h42b10757};
test_input[33552:33559] = '{32'hc1e5d808, 32'hc294528d, 32'h4285d789, 32'hc247e185, 32'h3fc9a70e, 32'hc2ad0b61, 32'h42c1baa8, 32'h424dc08b};
test_output[33552:33559] = '{32'h0, 32'h0, 32'h4285d789, 32'h0, 32'h3fc9a70e, 32'h0, 32'h42c1baa8, 32'h424dc08b};
test_input[33560:33567] = '{32'h41060783, 32'hc2a516e7, 32'h42affd8b, 32'hc249b54a, 32'h4289ecf9, 32'hc2b0f5ce, 32'hc2962238, 32'hc2398427};
test_output[33560:33567] = '{32'h41060783, 32'h0, 32'h42affd8b, 32'h0, 32'h4289ecf9, 32'h0, 32'h0, 32'h0};
test_input[33568:33575] = '{32'hc2b73567, 32'h420b26b3, 32'hc138f76f, 32'hc19ec4d6, 32'h42a261d4, 32'hc28fa38d, 32'h42ae009f, 32'h428dc071};
test_output[33568:33575] = '{32'h0, 32'h420b26b3, 32'h0, 32'h0, 32'h42a261d4, 32'h0, 32'h42ae009f, 32'h428dc071};
test_input[33576:33583] = '{32'h42a10aa8, 32'hc244f55a, 32'hc1b7b0c0, 32'hc224e1a1, 32'hc1c47fbe, 32'hc24efd0c, 32'hc1c87326, 32'hc2b0f753};
test_output[33576:33583] = '{32'h42a10aa8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[33584:33591] = '{32'hc1bca10b, 32'h42a9a7df, 32'h402bf5bc, 32'h424a3731, 32'hc2a7b3c5, 32'hc2b2ca94, 32'hc2a1e76a, 32'h4206518a};
test_output[33584:33591] = '{32'h0, 32'h42a9a7df, 32'h402bf5bc, 32'h424a3731, 32'h0, 32'h0, 32'h0, 32'h4206518a};
test_input[33592:33599] = '{32'hc28547e2, 32'hc23cd1a9, 32'hc290d100, 32'hc2860a03, 32'hc277136a, 32'h4147ff9f, 32'h41070e12, 32'hc11ee04f};
test_output[33592:33599] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4147ff9f, 32'h41070e12, 32'h0};
test_input[33600:33607] = '{32'hc2ace8b9, 32'hc210d58b, 32'h42521afb, 32'hc281f801, 32'hc27508f4, 32'h41236021, 32'h423ffc95, 32'hc16fc095};
test_output[33600:33607] = '{32'h0, 32'h0, 32'h42521afb, 32'h0, 32'h0, 32'h41236021, 32'h423ffc95, 32'h0};
test_input[33608:33615] = '{32'h42ad9270, 32'hc1263a37, 32'h4283b393, 32'hc294ac4c, 32'hc25fee4c, 32'h42268e97, 32'hc2605997, 32'hc2c17635};
test_output[33608:33615] = '{32'h42ad9270, 32'h0, 32'h4283b393, 32'h0, 32'h0, 32'h42268e97, 32'h0, 32'h0};
test_input[33616:33623] = '{32'h41346c56, 32'h426b436d, 32'h429b7a09, 32'hc2aa7468, 32'h42986306, 32'hc1834fff, 32'h429835d7, 32'hc1e89808};
test_output[33616:33623] = '{32'h41346c56, 32'h426b436d, 32'h429b7a09, 32'h0, 32'h42986306, 32'h0, 32'h429835d7, 32'h0};
test_input[33624:33631] = '{32'hc286c2da, 32'hc238195c, 32'hc2a3af4f, 32'h42163d5f, 32'hc20ab09f, 32'h42057164, 32'hc28cc1a4, 32'hc2c71e32};
test_output[33624:33631] = '{32'h0, 32'h0, 32'h0, 32'h42163d5f, 32'h0, 32'h42057164, 32'h0, 32'h0};
test_input[33632:33639] = '{32'h4113a592, 32'hc202b4c5, 32'h4259ecfb, 32'hc2a5cfa7, 32'hc1db9508, 32'h421416aa, 32'hc2330809, 32'hc2bd51f5};
test_output[33632:33639] = '{32'h4113a592, 32'h0, 32'h4259ecfb, 32'h0, 32'h0, 32'h421416aa, 32'h0, 32'h0};
test_input[33640:33647] = '{32'h41a758dd, 32'h4273cd48, 32'hc258449b, 32'hc1f20100, 32'h42482543, 32'hc28d3ce6, 32'h42097449, 32'h4297996e};
test_output[33640:33647] = '{32'h41a758dd, 32'h4273cd48, 32'h0, 32'h0, 32'h42482543, 32'h0, 32'h42097449, 32'h4297996e};
test_input[33648:33655] = '{32'hc195a51b, 32'hc2795cdc, 32'h42c415c5, 32'hc2aa585c, 32'hc2309af7, 32'h42c51f03, 32'h4237b1cb, 32'h42afd815};
test_output[33648:33655] = '{32'h0, 32'h0, 32'h42c415c5, 32'h0, 32'h0, 32'h42c51f03, 32'h4237b1cb, 32'h42afd815};
test_input[33656:33663] = '{32'hc0c6a9a5, 32'h42bd548b, 32'hc1f000a5, 32'h4239d528, 32'h427e32d1, 32'hc2b572c6, 32'h428ca29b, 32'h426bd0e0};
test_output[33656:33663] = '{32'h0, 32'h42bd548b, 32'h0, 32'h4239d528, 32'h427e32d1, 32'h0, 32'h428ca29b, 32'h426bd0e0};
test_input[33664:33671] = '{32'h42b16e28, 32'hc1c2363b, 32'h413fbc3d, 32'hc195c878, 32'hc169ec5f, 32'hc2adcc2b, 32'hbf97d82d, 32'hc289520a};
test_output[33664:33671] = '{32'h42b16e28, 32'h0, 32'h413fbc3d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[33672:33679] = '{32'hc0735213, 32'hc2967099, 32'h42bb2a77, 32'h42343451, 32'hc1e8a469, 32'h4149e667, 32'h41a8fe12, 32'h4295f77c};
test_output[33672:33679] = '{32'h0, 32'h0, 32'h42bb2a77, 32'h42343451, 32'h0, 32'h4149e667, 32'h41a8fe12, 32'h4295f77c};
test_input[33680:33687] = '{32'hc2bca49b, 32'h41d62939, 32'hc01e2992, 32'hc28f883e, 32'hc296e924, 32'h41d76157, 32'h42795f6a, 32'hc2b86adb};
test_output[33680:33687] = '{32'h0, 32'h41d62939, 32'h0, 32'h0, 32'h0, 32'h41d76157, 32'h42795f6a, 32'h0};
test_input[33688:33695] = '{32'hc277d6a2, 32'h42a77963, 32'hc048f48f, 32'hc2014cc1, 32'h42a39d4d, 32'h428508e1, 32'h41d5c93a, 32'h421cfa8b};
test_output[33688:33695] = '{32'h0, 32'h42a77963, 32'h0, 32'h0, 32'h42a39d4d, 32'h428508e1, 32'h41d5c93a, 32'h421cfa8b};
test_input[33696:33703] = '{32'h427462a8, 32'h42be3c4d, 32'h4140e756, 32'hc2ba3c1e, 32'h428785e4, 32'h4297eb1b, 32'h42bb2150, 32'hc2500d90};
test_output[33696:33703] = '{32'h427462a8, 32'h42be3c4d, 32'h4140e756, 32'h0, 32'h428785e4, 32'h4297eb1b, 32'h42bb2150, 32'h0};
test_input[33704:33711] = '{32'h3f91f7e8, 32'h421aab80, 32'hc18502a1, 32'hc08f69c8, 32'hc18804ea, 32'hc282d1df, 32'h426c8ad4, 32'h41f8994f};
test_output[33704:33711] = '{32'h3f91f7e8, 32'h421aab80, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426c8ad4, 32'h41f8994f};
test_input[33712:33719] = '{32'hc2177dad, 32'hbf94cb36, 32'hc294a137, 32'h42678027, 32'hc2aecfdc, 32'hc1008055, 32'hc298e23f, 32'hc1b47a81};
test_output[33712:33719] = '{32'h0, 32'h0, 32'h0, 32'h42678027, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[33720:33727] = '{32'hc2a58195, 32'hc22ef1ad, 32'hc211a0b5, 32'hc2b82e30, 32'hc12bd040, 32'h4224eba7, 32'h427c01c5, 32'hc0b0523a};
test_output[33720:33727] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4224eba7, 32'h427c01c5, 32'h0};
test_input[33728:33735] = '{32'hc2a266d1, 32'hc2033709, 32'h4091fa87, 32'hc2b46f87, 32'h42b1087b, 32'h42b98983, 32'h42c72c99, 32'hc2584f0f};
test_output[33728:33735] = '{32'h0, 32'h0, 32'h4091fa87, 32'h0, 32'h42b1087b, 32'h42b98983, 32'h42c72c99, 32'h0};
test_input[33736:33743] = '{32'h429428fe, 32'hc1735825, 32'h427f9c93, 32'h41ff7c9c, 32'h4259e7a9, 32'hc160a702, 32'hc1dd1ad4, 32'h423d62c1};
test_output[33736:33743] = '{32'h429428fe, 32'h0, 32'h427f9c93, 32'h41ff7c9c, 32'h4259e7a9, 32'h0, 32'h0, 32'h423d62c1};
test_input[33744:33751] = '{32'hc252b7e3, 32'h4268e79e, 32'h42acb075, 32'hc2616560, 32'h42818fb3, 32'hc250d778, 32'h429677d8, 32'h424dcaf5};
test_output[33744:33751] = '{32'h0, 32'h4268e79e, 32'h42acb075, 32'h0, 32'h42818fb3, 32'h0, 32'h429677d8, 32'h424dcaf5};
test_input[33752:33759] = '{32'h42098ff3, 32'hc27b28e0, 32'h42ab7aa2, 32'h41064ce9, 32'hc20f5beb, 32'h4223c3e5, 32'hc14f8239, 32'hc1a9f090};
test_output[33752:33759] = '{32'h42098ff3, 32'h0, 32'h42ab7aa2, 32'h41064ce9, 32'h0, 32'h4223c3e5, 32'h0, 32'h0};
test_input[33760:33767] = '{32'h41bceb32, 32'h421f86ec, 32'h419c1c63, 32'h421be46c, 32'hc2b7da3b, 32'h425ddacb, 32'h427f6390, 32'h42659bc5};
test_output[33760:33767] = '{32'h41bceb32, 32'h421f86ec, 32'h419c1c63, 32'h421be46c, 32'h0, 32'h425ddacb, 32'h427f6390, 32'h42659bc5};
test_input[33768:33775] = '{32'h418ee4c6, 32'hc23e8f7a, 32'h42983f4e, 32'h41bc0677, 32'hc181f797, 32'hc2c14ccb, 32'h41dc862a, 32'h42404706};
test_output[33768:33775] = '{32'h418ee4c6, 32'h0, 32'h42983f4e, 32'h41bc0677, 32'h0, 32'h0, 32'h41dc862a, 32'h42404706};
test_input[33776:33783] = '{32'hc24d6a9b, 32'hc2a39208, 32'hc2919e9e, 32'hc28c1276, 32'h401f61fa, 32'hc2a9b2a5, 32'h4210d5c4, 32'hc1cac144};
test_output[33776:33783] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h401f61fa, 32'h0, 32'h4210d5c4, 32'h0};
test_input[33784:33791] = '{32'h3e917d71, 32'hc2b74432, 32'h4273b256, 32'hc1d59f42, 32'h411a54f1, 32'h42c361fd, 32'h420ed7c7, 32'hc2c2a247};
test_output[33784:33791] = '{32'h3e917d71, 32'h0, 32'h4273b256, 32'h0, 32'h411a54f1, 32'h42c361fd, 32'h420ed7c7, 32'h0};
test_input[33792:33799] = '{32'hc2af9538, 32'h4255d898, 32'hc2be873b, 32'hc137a0bf, 32'h42417a5e, 32'h42c18c2a, 32'hc2a64dac, 32'h42c3f35f};
test_output[33792:33799] = '{32'h0, 32'h4255d898, 32'h0, 32'h0, 32'h42417a5e, 32'h42c18c2a, 32'h0, 32'h42c3f35f};
test_input[33800:33807] = '{32'h42b394e8, 32'h4292e057, 32'h42bb43c2, 32'h41c51135, 32'hc2176b17, 32'hc2389bc9, 32'h40041569, 32'h4287b088};
test_output[33800:33807] = '{32'h42b394e8, 32'h4292e057, 32'h42bb43c2, 32'h41c51135, 32'h0, 32'h0, 32'h40041569, 32'h4287b088};
test_input[33808:33815] = '{32'h41ef41f4, 32'h41dbe26a, 32'h4287514c, 32'h41079157, 32'hc18e2f67, 32'hc2811620, 32'hc0ceccd7, 32'hc20ea1de};
test_output[33808:33815] = '{32'h41ef41f4, 32'h41dbe26a, 32'h4287514c, 32'h41079157, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[33816:33823] = '{32'h428df27f, 32'hc1f76b04, 32'hc0aefc10, 32'hc2854c4e, 32'hc2bdc3c1, 32'h425254ca, 32'h41ba4be4, 32'h4023f498};
test_output[33816:33823] = '{32'h428df27f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h425254ca, 32'h41ba4be4, 32'h4023f498};
test_input[33824:33831] = '{32'h41dedf87, 32'hc1229b2c, 32'hc255a08f, 32'hc27075b2, 32'h41a39111, 32'h4254c6ee, 32'h421edab6, 32'h428e8ec1};
test_output[33824:33831] = '{32'h41dedf87, 32'h0, 32'h0, 32'h0, 32'h41a39111, 32'h4254c6ee, 32'h421edab6, 32'h428e8ec1};
test_input[33832:33839] = '{32'hc2199533, 32'hc1c20d8d, 32'h412488cf, 32'h42abde8b, 32'h42227632, 32'h41120162, 32'hbea2c529, 32'h42a2cde9};
test_output[33832:33839] = '{32'h0, 32'h0, 32'h412488cf, 32'h42abde8b, 32'h42227632, 32'h41120162, 32'h0, 32'h42a2cde9};
test_input[33840:33847] = '{32'hc1f046bd, 32'h42b9df75, 32'h40b01aae, 32'h420fe6d9, 32'h406d3637, 32'h42aaa6ec, 32'h42b02a6e, 32'hc2c40693};
test_output[33840:33847] = '{32'h0, 32'h42b9df75, 32'h40b01aae, 32'h420fe6d9, 32'h406d3637, 32'h42aaa6ec, 32'h42b02a6e, 32'h0};
test_input[33848:33855] = '{32'h42712587, 32'hc281bf1f, 32'hc2a44fed, 32'hc1876a0b, 32'hc2641dab, 32'hc1b684a7, 32'hc23e2615, 32'hc1a4e79e};
test_output[33848:33855] = '{32'h42712587, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[33856:33863] = '{32'hc18d9903, 32'h413d02ee, 32'h423512d3, 32'h413a10cf, 32'hc2b98359, 32'hc29459ee, 32'h42ae2b2d, 32'hc2b151ac};
test_output[33856:33863] = '{32'h0, 32'h413d02ee, 32'h423512d3, 32'h413a10cf, 32'h0, 32'h0, 32'h42ae2b2d, 32'h0};
test_input[33864:33871] = '{32'hc2adc30e, 32'hc29dc153, 32'hc180fb83, 32'h42a849c9, 32'h41ab9a9f, 32'hc22fc832, 32'h4210410f, 32'hc2499f4b};
test_output[33864:33871] = '{32'h0, 32'h0, 32'h0, 32'h42a849c9, 32'h41ab9a9f, 32'h0, 32'h4210410f, 32'h0};
test_input[33872:33879] = '{32'hc2acf084, 32'h42a0b1af, 32'hc29c6762, 32'hc2a62c6f, 32'h42429c7d, 32'h42013d46, 32'h4102c6b2, 32'h42a1cf85};
test_output[33872:33879] = '{32'h0, 32'h42a0b1af, 32'h0, 32'h0, 32'h42429c7d, 32'h42013d46, 32'h4102c6b2, 32'h42a1cf85};
test_input[33880:33887] = '{32'h41af5ede, 32'h418f8039, 32'h4250a4fd, 32'hc215cfb9, 32'hc24e7c2b, 32'h41a14688, 32'h422e1f77, 32'hc2a14d41};
test_output[33880:33887] = '{32'h41af5ede, 32'h418f8039, 32'h4250a4fd, 32'h0, 32'h0, 32'h41a14688, 32'h422e1f77, 32'h0};
test_input[33888:33895] = '{32'hc1bc2d5d, 32'hc231f25c, 32'h4084968c, 32'hc18eb3df, 32'h4254b4a0, 32'hc1eca661, 32'h42ae81c7, 32'h42862780};
test_output[33888:33895] = '{32'h0, 32'h0, 32'h4084968c, 32'h0, 32'h4254b4a0, 32'h0, 32'h42ae81c7, 32'h42862780};
test_input[33896:33903] = '{32'h428510d7, 32'h4296568c, 32'hc29b8102, 32'h42898102, 32'hc29a1da0, 32'hc1ebc969, 32'hc2218fe3, 32'hc1344edf};
test_output[33896:33903] = '{32'h428510d7, 32'h4296568c, 32'h0, 32'h42898102, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[33904:33911] = '{32'h42a9563e, 32'hc2b894b9, 32'hc2503f7b, 32'hc22ea05a, 32'h429f5d19, 32'h413d47e3, 32'h429e893b, 32'h421d04bc};
test_output[33904:33911] = '{32'h42a9563e, 32'h0, 32'h0, 32'h0, 32'h429f5d19, 32'h413d47e3, 32'h429e893b, 32'h421d04bc};
test_input[33912:33919] = '{32'h419eda86, 32'hc07760d4, 32'hc283837e, 32'hc209920d, 32'h42be90c4, 32'h422f3bd4, 32'hc0f08ac0, 32'hc0a2d149};
test_output[33912:33919] = '{32'h419eda86, 32'h0, 32'h0, 32'h0, 32'h42be90c4, 32'h422f3bd4, 32'h0, 32'h0};
test_input[33920:33927] = '{32'h42a72cfd, 32'h4223b4c2, 32'h423b4443, 32'h428b21dc, 32'h4251abcc, 32'h424f9d47, 32'hc1a225d2, 32'hc2a76f00};
test_output[33920:33927] = '{32'h42a72cfd, 32'h4223b4c2, 32'h423b4443, 32'h428b21dc, 32'h4251abcc, 32'h424f9d47, 32'h0, 32'h0};
test_input[33928:33935] = '{32'hc0217b96, 32'hc21e746d, 32'hc2992812, 32'h426f774c, 32'h4241c6cb, 32'hc2830161, 32'h41066333, 32'h4119933a};
test_output[33928:33935] = '{32'h0, 32'h0, 32'h0, 32'h426f774c, 32'h4241c6cb, 32'h0, 32'h41066333, 32'h4119933a};
test_input[33936:33943] = '{32'hc1cd0bd2, 32'h41929fe3, 32'h428e6501, 32'h4288e080, 32'hc2aac93f, 32'h42495586, 32'h42276093, 32'hc29a13a5};
test_output[33936:33943] = '{32'h0, 32'h41929fe3, 32'h428e6501, 32'h4288e080, 32'h0, 32'h42495586, 32'h42276093, 32'h0};
test_input[33944:33951] = '{32'hc1d44bbe, 32'hc1f40b83, 32'hc10c1299, 32'hc2af0b92, 32'h41a7be0e, 32'h41a1b733, 32'h4277e4e2, 32'hbf3f4ac7};
test_output[33944:33951] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41a7be0e, 32'h41a1b733, 32'h4277e4e2, 32'h0};
test_input[33952:33959] = '{32'hc22943cb, 32'hc2348031, 32'h42090afc, 32'hc28b3138, 32'hc12fbe8a, 32'h42a10b0a, 32'hc2b7a8f8, 32'h418dac61};
test_output[33952:33959] = '{32'h0, 32'h0, 32'h42090afc, 32'h0, 32'h0, 32'h42a10b0a, 32'h0, 32'h418dac61};
test_input[33960:33967] = '{32'h417c57e4, 32'h42742d77, 32'h4281b769, 32'h419eeacf, 32'hc109acb5, 32'hc1c7382f, 32'h41c6eb37, 32'h42130336};
test_output[33960:33967] = '{32'h417c57e4, 32'h42742d77, 32'h4281b769, 32'h419eeacf, 32'h0, 32'h0, 32'h41c6eb37, 32'h42130336};
test_input[33968:33975] = '{32'h4291bb49, 32'hc23aa0f4, 32'hc2905d5d, 32'h427376be, 32'hc28c656b, 32'h41805701, 32'h4243f3b9, 32'hc2aa9b56};
test_output[33968:33975] = '{32'h4291bb49, 32'h0, 32'h0, 32'h427376be, 32'h0, 32'h41805701, 32'h4243f3b9, 32'h0};
test_input[33976:33983] = '{32'hc1423581, 32'hc0bcc5ed, 32'h41d70927, 32'h428810f8, 32'h424fae09, 32'hc190d7ea, 32'hc2445380, 32'hc2a5723a};
test_output[33976:33983] = '{32'h0, 32'h0, 32'h41d70927, 32'h428810f8, 32'h424fae09, 32'h0, 32'h0, 32'h0};
test_input[33984:33991] = '{32'hc26ef626, 32'hc2623085, 32'h42716fb7, 32'hc2bb3a69, 32'hc164e9a0, 32'hc211708d, 32'h428b621f, 32'h40535dc8};
test_output[33984:33991] = '{32'h0, 32'h0, 32'h42716fb7, 32'h0, 32'h0, 32'h0, 32'h428b621f, 32'h40535dc8};
test_input[33992:33999] = '{32'h4123308a, 32'hc2bd9bc3, 32'h42a1df97, 32'hc26a14b1, 32'hc2bf4de6, 32'h4142caff, 32'h40abbcbf, 32'h4067f3f4};
test_output[33992:33999] = '{32'h4123308a, 32'h0, 32'h42a1df97, 32'h0, 32'h0, 32'h4142caff, 32'h40abbcbf, 32'h4067f3f4};
test_input[34000:34007] = '{32'hc23684df, 32'h42928ff5, 32'hbe641cda, 32'hc2c796f1, 32'h4298c3db, 32'h419965d8, 32'hc23d59bf, 32'hc2806a1a};
test_output[34000:34007] = '{32'h0, 32'h42928ff5, 32'h0, 32'h0, 32'h4298c3db, 32'h419965d8, 32'h0, 32'h0};
test_input[34008:34015] = '{32'hc09d879e, 32'h4289e408, 32'hc0da4112, 32'h3f594390, 32'hbfd16b04, 32'h4285aa5d, 32'h420230ef, 32'hc21d96a9};
test_output[34008:34015] = '{32'h0, 32'h4289e408, 32'h0, 32'h3f594390, 32'h0, 32'h4285aa5d, 32'h420230ef, 32'h0};
test_input[34016:34023] = '{32'hc0e54692, 32'hc2b1007f, 32'hc2a7b352, 32'hc1d4dc86, 32'h4255a7f7, 32'hc2126bcb, 32'hc2adf02e, 32'h429f0e9e};
test_output[34016:34023] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4255a7f7, 32'h0, 32'h0, 32'h429f0e9e};
test_input[34024:34031] = '{32'hc2c61c71, 32'h4262c753, 32'h4273b853, 32'h427334b3, 32'h4274d5fc, 32'h42491599, 32'hc1e3cbb6, 32'hc031afe0};
test_output[34024:34031] = '{32'h0, 32'h4262c753, 32'h4273b853, 32'h427334b3, 32'h4274d5fc, 32'h42491599, 32'h0, 32'h0};
test_input[34032:34039] = '{32'hc23b736d, 32'h42384d41, 32'h41fa4043, 32'hc26526ba, 32'hc28704ee, 32'h40102663, 32'h423470d8, 32'hc24fbad5};
test_output[34032:34039] = '{32'h0, 32'h42384d41, 32'h41fa4043, 32'h0, 32'h0, 32'h40102663, 32'h423470d8, 32'h0};
test_input[34040:34047] = '{32'h42a7d236, 32'h4239ff6c, 32'hc299ada9, 32'h4207118b, 32'hc24c44ed, 32'hc231b5aa, 32'h42aa59ac, 32'hbfc7fff1};
test_output[34040:34047] = '{32'h42a7d236, 32'h4239ff6c, 32'h0, 32'h4207118b, 32'h0, 32'h0, 32'h42aa59ac, 32'h0};
test_input[34048:34055] = '{32'hc21357cc, 32'hc1460e22, 32'h41b46991, 32'hc2a17e8c, 32'hc2ba8f46, 32'h420b7f45, 32'hc24454df, 32'h41c89d0c};
test_output[34048:34055] = '{32'h0, 32'h0, 32'h41b46991, 32'h0, 32'h0, 32'h420b7f45, 32'h0, 32'h41c89d0c};
test_input[34056:34063] = '{32'hc2afdf5a, 32'hc245bf21, 32'h41a6da80, 32'h42a7f51f, 32'hc203011e, 32'h4160a7c2, 32'hc25e351d, 32'hc24b7c77};
test_output[34056:34063] = '{32'h0, 32'h0, 32'h41a6da80, 32'h42a7f51f, 32'h0, 32'h4160a7c2, 32'h0, 32'h0};
test_input[34064:34071] = '{32'h42572b01, 32'hc28f32ab, 32'h42130fa5, 32'h428816e0, 32'hc1b82184, 32'h425201c5, 32'h3fa1d744, 32'hc22534cf};
test_output[34064:34071] = '{32'h42572b01, 32'h0, 32'h42130fa5, 32'h428816e0, 32'h0, 32'h425201c5, 32'h3fa1d744, 32'h0};
test_input[34072:34079] = '{32'hc15a92b7, 32'h42762078, 32'hc275cfc3, 32'hc2c4221a, 32'h42a8597b, 32'hc211d3cd, 32'h426340bc, 32'h4224295d};
test_output[34072:34079] = '{32'h0, 32'h42762078, 32'h0, 32'h0, 32'h42a8597b, 32'h0, 32'h426340bc, 32'h4224295d};
test_input[34080:34087] = '{32'hc2a13fa7, 32'h42af89cf, 32'hc2a0f96b, 32'hc2a49f33, 32'h426fea92, 32'h429b7c3d, 32'h4295cbcd, 32'hc291d929};
test_output[34080:34087] = '{32'h0, 32'h42af89cf, 32'h0, 32'h0, 32'h426fea92, 32'h429b7c3d, 32'h4295cbcd, 32'h0};
test_input[34088:34095] = '{32'hc2ae9e2c, 32'hc2b62500, 32'hc29d7536, 32'hc240885d, 32'h419f555b, 32'hc2948371, 32'h41944917, 32'hc20bda3e};
test_output[34088:34095] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h419f555b, 32'h0, 32'h41944917, 32'h0};
test_input[34096:34103] = '{32'hbed08781, 32'hc28bb86f, 32'h4214e02e, 32'hc25e8d0a, 32'hc2a2fc95, 32'hc29c54b9, 32'h415b4a06, 32'h41d2aba2};
test_output[34096:34103] = '{32'h0, 32'h0, 32'h4214e02e, 32'h0, 32'h0, 32'h0, 32'h415b4a06, 32'h41d2aba2};
test_input[34104:34111] = '{32'hc2224e8d, 32'hc19628c0, 32'hc2108578, 32'h4248a2fb, 32'h417ba2b0, 32'hc11476af, 32'h42a6e5d0, 32'h41f250ab};
test_output[34104:34111] = '{32'h0, 32'h0, 32'h0, 32'h4248a2fb, 32'h417ba2b0, 32'h0, 32'h42a6e5d0, 32'h41f250ab};
test_input[34112:34119] = '{32'h41f99112, 32'h42830e31, 32'h42610dca, 32'hc2c4302b, 32'hc2b9977c, 32'hc0f99370, 32'hc20c2b3c, 32'hc2b69074};
test_output[34112:34119] = '{32'h41f99112, 32'h42830e31, 32'h42610dca, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[34120:34127] = '{32'hc196bd24, 32'h4201ba66, 32'hc208cd0d, 32'hc2a8404a, 32'hc24108b8, 32'h421bd2e4, 32'hc2a5ca80, 32'h42846b6a};
test_output[34120:34127] = '{32'h0, 32'h4201ba66, 32'h0, 32'h0, 32'h0, 32'h421bd2e4, 32'h0, 32'h42846b6a};
test_input[34128:34135] = '{32'hc2b539f9, 32'h41210f47, 32'hc2963382, 32'h42b163f6, 32'hc20c3f09, 32'hc2610739, 32'h4295746d, 32'h42c35bfe};
test_output[34128:34135] = '{32'h0, 32'h41210f47, 32'h0, 32'h42b163f6, 32'h0, 32'h0, 32'h4295746d, 32'h42c35bfe};
test_input[34136:34143] = '{32'h42ae2dd0, 32'h42ae1d25, 32'h428ebd4b, 32'hc29fdca8, 32'hc283970a, 32'h42bacb50, 32'h41cf20fa, 32'hc1e90f14};
test_output[34136:34143] = '{32'h42ae2dd0, 32'h42ae1d25, 32'h428ebd4b, 32'h0, 32'h0, 32'h42bacb50, 32'h41cf20fa, 32'h0};
test_input[34144:34151] = '{32'h41b4e90b, 32'h4033ead9, 32'hc2b45233, 32'h42309a67, 32'hc18ca25e, 32'hc246c1b8, 32'h427f0fc3, 32'h42a56849};
test_output[34144:34151] = '{32'h41b4e90b, 32'h4033ead9, 32'h0, 32'h42309a67, 32'h0, 32'h0, 32'h427f0fc3, 32'h42a56849};
test_input[34152:34159] = '{32'h409213d6, 32'h42b7f3f6, 32'hbf12ed7a, 32'hc1e17924, 32'h425cb73b, 32'hc2c7511d, 32'h41ca342a, 32'h423c3b9b};
test_output[34152:34159] = '{32'h409213d6, 32'h42b7f3f6, 32'h0, 32'h0, 32'h425cb73b, 32'h0, 32'h41ca342a, 32'h423c3b9b};
test_input[34160:34167] = '{32'h428f0810, 32'hc1d2dd1c, 32'hc1595f9e, 32'h413317a5, 32'h42c4580d, 32'h42a4edcf, 32'h427a0cf6, 32'hc2492962};
test_output[34160:34167] = '{32'h428f0810, 32'h0, 32'h0, 32'h413317a5, 32'h42c4580d, 32'h42a4edcf, 32'h427a0cf6, 32'h0};
test_input[34168:34175] = '{32'hc2b4fb00, 32'hc2854568, 32'hc2149705, 32'hc2b9b83b, 32'hc01127dd, 32'hc1e18bae, 32'hc296282b, 32'h4262edc3};
test_output[34168:34175] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4262edc3};
test_input[34176:34183] = '{32'h4285f7a4, 32'hc0747fae, 32'hc205b7c2, 32'h42ae8a48, 32'hc16238a5, 32'hc28d7976, 32'h424a0c4a, 32'h41e70653};
test_output[34176:34183] = '{32'h4285f7a4, 32'h0, 32'h0, 32'h42ae8a48, 32'h0, 32'h0, 32'h424a0c4a, 32'h41e70653};
test_input[34184:34191] = '{32'h429eb5e4, 32'hc182fd68, 32'hc2597f51, 32'h42595063, 32'h40e26ee2, 32'hc229a2f7, 32'hc26b9031, 32'hc1d1d896};
test_output[34184:34191] = '{32'h429eb5e4, 32'h0, 32'h0, 32'h42595063, 32'h40e26ee2, 32'h0, 32'h0, 32'h0};
test_input[34192:34199] = '{32'h423767bc, 32'h42bbbe3a, 32'h4292d80b, 32'h4291b097, 32'hc26ae9f2, 32'h41958b14, 32'h42782edf, 32'h429103e8};
test_output[34192:34199] = '{32'h423767bc, 32'h42bbbe3a, 32'h4292d80b, 32'h4291b097, 32'h0, 32'h41958b14, 32'h42782edf, 32'h429103e8};
test_input[34200:34207] = '{32'hc26651f7, 32'hc1f9ae23, 32'hc110ba44, 32'hc210cfb5, 32'hc28d68a5, 32'hc0c5dea7, 32'h423a6a72, 32'hc2c215af};
test_output[34200:34207] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423a6a72, 32'h0};
test_input[34208:34215] = '{32'hc18d65a7, 32'h40ca64cc, 32'hc1a80f96, 32'h42b6d403, 32'hc2bb81a9, 32'h4268dbf2, 32'hc254af5e, 32'hc28bf2e6};
test_output[34208:34215] = '{32'h0, 32'h40ca64cc, 32'h0, 32'h42b6d403, 32'h0, 32'h4268dbf2, 32'h0, 32'h0};
test_input[34216:34223] = '{32'h41df6edc, 32'h4207f36c, 32'h42946eb1, 32'hc2b9cbe0, 32'hc287c91c, 32'hc271d09a, 32'hc1b8cb65, 32'h4198b1de};
test_output[34216:34223] = '{32'h41df6edc, 32'h4207f36c, 32'h42946eb1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4198b1de};
test_input[34224:34231] = '{32'h42b385e9, 32'h423e01d2, 32'hc23bf779, 32'h418340c1, 32'hc045ecd7, 32'hc0948324, 32'hc28fcb44, 32'hbfc487ed};
test_output[34224:34231] = '{32'h42b385e9, 32'h423e01d2, 32'h0, 32'h418340c1, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[34232:34239] = '{32'h42baf9c8, 32'hc29f69ae, 32'hc216486f, 32'h428523d9, 32'hc29231ec, 32'h3e262844, 32'hc2086b04, 32'hc1d390fb};
test_output[34232:34239] = '{32'h42baf9c8, 32'h0, 32'h0, 32'h428523d9, 32'h0, 32'h3e262844, 32'h0, 32'h0};
test_input[34240:34247] = '{32'hc29d7668, 32'hc2b5d8ea, 32'hc2440320, 32'hc28b8e47, 32'hc2ac4774, 32'h4223e8f8, 32'h42319882, 32'h4233934e};
test_output[34240:34247] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4223e8f8, 32'h42319882, 32'h4233934e};
test_input[34248:34255] = '{32'hc14d0a8d, 32'hc29bed90, 32'hc1f226ec, 32'h42b66613, 32'hc29aaede, 32'hc282303a, 32'hc2b35190, 32'hc266b1d7};
test_output[34248:34255] = '{32'h0, 32'h0, 32'h0, 32'h42b66613, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[34256:34263] = '{32'h41a43d01, 32'h4233c224, 32'h42733bcd, 32'hc209df95, 32'hc2072a85, 32'hc29695db, 32'h429054d1, 32'hc2aa1deb};
test_output[34256:34263] = '{32'h41a43d01, 32'h4233c224, 32'h42733bcd, 32'h0, 32'h0, 32'h0, 32'h429054d1, 32'h0};
test_input[34264:34271] = '{32'hc2b48c11, 32'hc286b1e9, 32'hc1f5d9cb, 32'h424f3ced, 32'h41eab1c2, 32'h4244068e, 32'hc2bd4726, 32'h423014ee};
test_output[34264:34271] = '{32'h0, 32'h0, 32'h0, 32'h424f3ced, 32'h41eab1c2, 32'h4244068e, 32'h0, 32'h423014ee};
test_input[34272:34279] = '{32'h40c86d74, 32'h42a6c4ac, 32'hbfe9876f, 32'h427871da, 32'hc2129d73, 32'hc2b85618, 32'hc23b4f49, 32'h424e151c};
test_output[34272:34279] = '{32'h40c86d74, 32'h42a6c4ac, 32'h0, 32'h427871da, 32'h0, 32'h0, 32'h0, 32'h424e151c};
test_input[34280:34287] = '{32'hc28cd04b, 32'h4135065b, 32'hc289d6ad, 32'hc28121dd, 32'hc227e7cd, 32'hc1f009e0, 32'h42bf32d4, 32'h3e071679};
test_output[34280:34287] = '{32'h0, 32'h4135065b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bf32d4, 32'h3e071679};
test_input[34288:34295] = '{32'h41abdb42, 32'hc16d13c8, 32'hc2bc10d4, 32'hc299620b, 32'h428040d4, 32'h41fe90ab, 32'hc2c69ded, 32'h42be47d4};
test_output[34288:34295] = '{32'h41abdb42, 32'h0, 32'h0, 32'h0, 32'h428040d4, 32'h41fe90ab, 32'h0, 32'h42be47d4};
test_input[34296:34303] = '{32'hc1b233ca, 32'h42c30e6d, 32'hc1aedd90, 32'h4282f5f5, 32'hc2a18496, 32'h4214e162, 32'hc2a5b7e3, 32'hc2c0ef70};
test_output[34296:34303] = '{32'h0, 32'h42c30e6d, 32'h0, 32'h4282f5f5, 32'h0, 32'h4214e162, 32'h0, 32'h0};
test_input[34304:34311] = '{32'hc2b89a77, 32'hc22e6a05, 32'hc288b4d2, 32'h4237b686, 32'hc2556135, 32'h42a5399f, 32'h411b9ce8, 32'hc14d4298};
test_output[34304:34311] = '{32'h0, 32'h0, 32'h0, 32'h4237b686, 32'h0, 32'h42a5399f, 32'h411b9ce8, 32'h0};
test_input[34312:34319] = '{32'hc2a01955, 32'hc276ed5a, 32'h4262d643, 32'hc285d888, 32'h3f921e91, 32'hc24e85c7, 32'h42b27a15, 32'hc19b3071};
test_output[34312:34319] = '{32'h0, 32'h0, 32'h4262d643, 32'h0, 32'h3f921e91, 32'h0, 32'h42b27a15, 32'h0};
test_input[34320:34327] = '{32'hc1675bae, 32'h41f6ce38, 32'h41eef4db, 32'hc1271914, 32'h41073239, 32'hc1c81a08, 32'hc231504a, 32'h42081019};
test_output[34320:34327] = '{32'h0, 32'h41f6ce38, 32'h41eef4db, 32'h0, 32'h41073239, 32'h0, 32'h0, 32'h42081019};
test_input[34328:34335] = '{32'hc0bd71d6, 32'hc060715d, 32'hc262d2b0, 32'h42a18d6c, 32'hc2b9c1aa, 32'hc27bb68a, 32'h42452b03, 32'hc2a5c2cf};
test_output[34328:34335] = '{32'h0, 32'h0, 32'h0, 32'h42a18d6c, 32'h0, 32'h0, 32'h42452b03, 32'h0};
test_input[34336:34343] = '{32'hc2c2a187, 32'h429f82c0, 32'h428d8372, 32'hc24abe52, 32'hc23f1543, 32'hc1e0327a, 32'h42b7b0b3, 32'h41566b89};
test_output[34336:34343] = '{32'h0, 32'h429f82c0, 32'h428d8372, 32'h0, 32'h0, 32'h0, 32'h42b7b0b3, 32'h41566b89};
test_input[34344:34351] = '{32'h428debc0, 32'hc240daf0, 32'h41f53098, 32'hc1910822, 32'hc1251de2, 32'h422a871f, 32'hc251641e, 32'h424f49f0};
test_output[34344:34351] = '{32'h428debc0, 32'h0, 32'h41f53098, 32'h0, 32'h0, 32'h422a871f, 32'h0, 32'h424f49f0};
test_input[34352:34359] = '{32'hc221f3dc, 32'hc2b6b5f1, 32'h4205c16d, 32'hc2a98221, 32'hc1ad1c65, 32'hc2578cd8, 32'hc10a0112, 32'h42617c43};
test_output[34352:34359] = '{32'h0, 32'h0, 32'h4205c16d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42617c43};
test_input[34360:34367] = '{32'h42446002, 32'hc1b8b9d6, 32'hc2b98d5d, 32'hc2bcdb59, 32'h41d2f9fd, 32'h42364da8, 32'h41ce1356, 32'h41d0a7a4};
test_output[34360:34367] = '{32'h42446002, 32'h0, 32'h0, 32'h0, 32'h41d2f9fd, 32'h42364da8, 32'h41ce1356, 32'h41d0a7a4};
test_input[34368:34375] = '{32'hc245e353, 32'h41118d18, 32'hc280122b, 32'h42c5c618, 32'h4295b8ee, 32'hc0c780d0, 32'hc1bf9c73, 32'h4249ecd8};
test_output[34368:34375] = '{32'h0, 32'h41118d18, 32'h0, 32'h42c5c618, 32'h4295b8ee, 32'h0, 32'h0, 32'h4249ecd8};
test_input[34376:34383] = '{32'h4275d84a, 32'h4270f5ef, 32'hc29ce04c, 32'hc10a09ed, 32'hc2c540d4, 32'hc1d4e2ea, 32'hc07aaebe, 32'hc239d72d};
test_output[34376:34383] = '{32'h4275d84a, 32'h4270f5ef, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[34384:34391] = '{32'h41e1b262, 32'h42b24de3, 32'hc292ef2a, 32'h42c4c313, 32'h425e9ffe, 32'h42b7d74f, 32'h42ac0553, 32'h41359e25};
test_output[34384:34391] = '{32'h41e1b262, 32'h42b24de3, 32'h0, 32'h42c4c313, 32'h425e9ffe, 32'h42b7d74f, 32'h42ac0553, 32'h41359e25};
test_input[34392:34399] = '{32'hc16d3e45, 32'hc1dcd94b, 32'hc2270242, 32'hc18761ce, 32'h4296fc0c, 32'hc298d1a6, 32'hc23d051b, 32'hc2023eb0};
test_output[34392:34399] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4296fc0c, 32'h0, 32'h0, 32'h0};
test_input[34400:34407] = '{32'h41559ec3, 32'h4252f1d1, 32'hc1a28c75, 32'h4296bc81, 32'h42548784, 32'h4156b984, 32'hc2b70fff, 32'hc2893bb6};
test_output[34400:34407] = '{32'h41559ec3, 32'h4252f1d1, 32'h0, 32'h4296bc81, 32'h42548784, 32'h4156b984, 32'h0, 32'h0};
test_input[34408:34415] = '{32'hc281a98b, 32'hc1c31459, 32'h4079ddf9, 32'h4299cf73, 32'hc04aaa0d, 32'h42901dd7, 32'h411a9ba1, 32'hc18b7beb};
test_output[34408:34415] = '{32'h0, 32'h0, 32'h4079ddf9, 32'h4299cf73, 32'h0, 32'h42901dd7, 32'h411a9ba1, 32'h0};
test_input[34416:34423] = '{32'hc1867e82, 32'h4234e69e, 32'hc199c774, 32'h418018fc, 32'h42771b20, 32'hc191aaa3, 32'h42be1164, 32'hc1c499ff};
test_output[34416:34423] = '{32'h0, 32'h4234e69e, 32'h0, 32'h418018fc, 32'h42771b20, 32'h0, 32'h42be1164, 32'h0};
test_input[34424:34431] = '{32'h40d1490c, 32'h4152018f, 32'h4292eec0, 32'hc2c60abb, 32'h4268eade, 32'hc249b710, 32'hc0e94b68, 32'h4272820e};
test_output[34424:34431] = '{32'h40d1490c, 32'h4152018f, 32'h4292eec0, 32'h0, 32'h4268eade, 32'h0, 32'h0, 32'h4272820e};
test_input[34432:34439] = '{32'h420f0370, 32'h42be1860, 32'hc28b9cc3, 32'hbf4cc415, 32'hc1815f57, 32'hc2b6b0e5, 32'hc0e31de9, 32'hbfdb0153};
test_output[34432:34439] = '{32'h420f0370, 32'h42be1860, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[34440:34447] = '{32'hc251a70e, 32'h41acf57f, 32'hc0c8a018, 32'h42704824, 32'h41831801, 32'hc1d7eb46, 32'hc28001cb, 32'hc169d817};
test_output[34440:34447] = '{32'h0, 32'h41acf57f, 32'h0, 32'h42704824, 32'h41831801, 32'h0, 32'h0, 32'h0};
test_input[34448:34455] = '{32'h421017df, 32'hc27e4b88, 32'h417ab379, 32'hc296ae92, 32'h42b15423, 32'hc2a95062, 32'h41f7fab3, 32'h42bbc948};
test_output[34448:34455] = '{32'h421017df, 32'h0, 32'h417ab379, 32'h0, 32'h42b15423, 32'h0, 32'h41f7fab3, 32'h42bbc948};
test_input[34456:34463] = '{32'hc27418e4, 32'hc2941a99, 32'h4220f438, 32'h42b6b7c7, 32'h427f9707, 32'h420313aa, 32'hc285139f, 32'hc2548596};
test_output[34456:34463] = '{32'h0, 32'h0, 32'h4220f438, 32'h42b6b7c7, 32'h427f9707, 32'h420313aa, 32'h0, 32'h0};
test_input[34464:34471] = '{32'hc2c1e7a9, 32'hc1ec9c29, 32'h420da2d3, 32'hc22cb651, 32'hc1de7903, 32'h41d3ac87, 32'hc10d748b, 32'hc2836a34};
test_output[34464:34471] = '{32'h0, 32'h0, 32'h420da2d3, 32'h0, 32'h0, 32'h41d3ac87, 32'h0, 32'h0};
test_input[34472:34479] = '{32'hc29200f6, 32'hc2587ab4, 32'h42a5513e, 32'hc23233d9, 32'h4218a772, 32'h4197cd0b, 32'h4259fff3, 32'h429859a3};
test_output[34472:34479] = '{32'h0, 32'h0, 32'h42a5513e, 32'h0, 32'h4218a772, 32'h4197cd0b, 32'h4259fff3, 32'h429859a3};
test_input[34480:34487] = '{32'hc1cd6816, 32'h429a999e, 32'hc0b080e8, 32'h427e95bd, 32'hc2a78e3f, 32'hc28fd5e7, 32'h42ae57b6, 32'h4211d63f};
test_output[34480:34487] = '{32'h0, 32'h429a999e, 32'h0, 32'h427e95bd, 32'h0, 32'h0, 32'h42ae57b6, 32'h4211d63f};
test_input[34488:34495] = '{32'h414ac4f0, 32'h41d7557b, 32'hc2316b81, 32'h419765bb, 32'h402ea917, 32'h423138c8, 32'h42742310, 32'h4209df45};
test_output[34488:34495] = '{32'h414ac4f0, 32'h41d7557b, 32'h0, 32'h419765bb, 32'h402ea917, 32'h423138c8, 32'h42742310, 32'h4209df45};
test_input[34496:34503] = '{32'h4196410b, 32'hc211e5cb, 32'h4264d0a0, 32'hc25b9af0, 32'h4271ce74, 32'h424a2f72, 32'h4184d875, 32'h429c6819};
test_output[34496:34503] = '{32'h4196410b, 32'h0, 32'h4264d0a0, 32'h0, 32'h4271ce74, 32'h424a2f72, 32'h4184d875, 32'h429c6819};
test_input[34504:34511] = '{32'h41a296a7, 32'h422f4485, 32'hc19e1e4a, 32'hc23c65c3, 32'hbe08f02d, 32'h4298445d, 32'hc26b5d63, 32'h41e1486a};
test_output[34504:34511] = '{32'h41a296a7, 32'h422f4485, 32'h0, 32'h0, 32'h0, 32'h4298445d, 32'h0, 32'h41e1486a};
test_input[34512:34519] = '{32'h42ba064a, 32'h42a6c267, 32'hc2506fb3, 32'hc080a576, 32'h429cf7de, 32'hc2b49855, 32'hc259abfe, 32'hc09e7a5f};
test_output[34512:34519] = '{32'h42ba064a, 32'h42a6c267, 32'h0, 32'h0, 32'h429cf7de, 32'h0, 32'h0, 32'h0};
test_input[34520:34527] = '{32'h4223e35f, 32'h41da0bfa, 32'hc11f7521, 32'h42a41331, 32'h41da3e8c, 32'h4292487d, 32'h428c6192, 32'hc29296ac};
test_output[34520:34527] = '{32'h4223e35f, 32'h41da0bfa, 32'h0, 32'h42a41331, 32'h41da3e8c, 32'h4292487d, 32'h428c6192, 32'h0};
test_input[34528:34535] = '{32'hc2b753b7, 32'h42c3b35e, 32'hc0b8d3c6, 32'h41fb1c26, 32'hc28d7d7d, 32'hc28e8de4, 32'hc28287ee, 32'h42ab3fac};
test_output[34528:34535] = '{32'h0, 32'h42c3b35e, 32'h0, 32'h41fb1c26, 32'h0, 32'h0, 32'h0, 32'h42ab3fac};
test_input[34536:34543] = '{32'hc2951e96, 32'h42a24460, 32'h402aa5fd, 32'hc250a24c, 32'hc2b25d73, 32'h42bb05cb, 32'hc0cf5dfc, 32'h428eee3d};
test_output[34536:34543] = '{32'h0, 32'h42a24460, 32'h402aa5fd, 32'h0, 32'h0, 32'h42bb05cb, 32'h0, 32'h428eee3d};
test_input[34544:34551] = '{32'h4169010b, 32'hc252499d, 32'h42b2b750, 32'h40a62e9e, 32'hc2842e78, 32'h4245eaf1, 32'h427a6cd9, 32'h41736c77};
test_output[34544:34551] = '{32'h4169010b, 32'h0, 32'h42b2b750, 32'h40a62e9e, 32'h0, 32'h4245eaf1, 32'h427a6cd9, 32'h41736c77};
test_input[34552:34559] = '{32'h42aca658, 32'hc2c39b53, 32'h42bbc812, 32'h4151d03b, 32'hc25b26f1, 32'hc2345aab, 32'hc2c78819, 32'hc184698a};
test_output[34552:34559] = '{32'h42aca658, 32'h0, 32'h42bbc812, 32'h4151d03b, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[34560:34567] = '{32'h42ac382f, 32'h4277e88b, 32'h41dbca6f, 32'h42bb533a, 32'hc28c4b90, 32'hc21d6a3a, 32'hc17f0734, 32'h41ce01f9};
test_output[34560:34567] = '{32'h42ac382f, 32'h4277e88b, 32'h41dbca6f, 32'h42bb533a, 32'h0, 32'h0, 32'h0, 32'h41ce01f9};
test_input[34568:34575] = '{32'h4163fd5c, 32'hc1f5b494, 32'h4297d180, 32'hc280b723, 32'h41ab1733, 32'h4174af4a, 32'hc259a46e, 32'hc237083a};
test_output[34568:34575] = '{32'h4163fd5c, 32'h0, 32'h4297d180, 32'h0, 32'h41ab1733, 32'h4174af4a, 32'h0, 32'h0};
test_input[34576:34583] = '{32'h42a2f455, 32'hc2b1ae23, 32'hc250bc5a, 32'h429f71c0, 32'hc224c706, 32'h41688235, 32'hc2be583f, 32'h4030fae0};
test_output[34576:34583] = '{32'h42a2f455, 32'h0, 32'h0, 32'h429f71c0, 32'h0, 32'h41688235, 32'h0, 32'h4030fae0};
test_input[34584:34591] = '{32'h42c707a0, 32'hc24c9c5b, 32'hc29d62c2, 32'hc12a50a7, 32'hc28698f9, 32'h4285a789, 32'hc2b1e182, 32'h4240f011};
test_output[34584:34591] = '{32'h42c707a0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4285a789, 32'h0, 32'h4240f011};
test_input[34592:34599] = '{32'h4212179c, 32'h4275f10e, 32'hc1968738, 32'hc22c8a04, 32'hc27320bf, 32'h421b39ed, 32'h42847296, 32'hc2b9dcc3};
test_output[34592:34599] = '{32'h4212179c, 32'h4275f10e, 32'h0, 32'h0, 32'h0, 32'h421b39ed, 32'h42847296, 32'h0};
test_input[34600:34607] = '{32'hc2b030b3, 32'h42891c95, 32'hc2bed4b7, 32'hc1784b46, 32'h42bf70e1, 32'hc24e4aca, 32'h4298ec91, 32'hc20f81ff};
test_output[34600:34607] = '{32'h0, 32'h42891c95, 32'h0, 32'h0, 32'h42bf70e1, 32'h0, 32'h4298ec91, 32'h0};
test_input[34608:34615] = '{32'hc229bdd2, 32'h42a6b4e8, 32'hc2172ca8, 32'hc1e05250, 32'hc18c6263, 32'h418fb5cc, 32'h42a5dfe6, 32'h422d5cfd};
test_output[34608:34615] = '{32'h0, 32'h42a6b4e8, 32'h0, 32'h0, 32'h0, 32'h418fb5cc, 32'h42a5dfe6, 32'h422d5cfd};
test_input[34616:34623] = '{32'hc1d72436, 32'hc10d029d, 32'hc24d9a93, 32'hc171e344, 32'hc1070884, 32'h41623b31, 32'hc2199a37, 32'h42a33e68};
test_output[34616:34623] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41623b31, 32'h0, 32'h42a33e68};
test_input[34624:34631] = '{32'h40e38364, 32'h41b9361e, 32'hc0db60b5, 32'h41d1a763, 32'h429a4ec9, 32'h423490d9, 32'h423f4132, 32'hc288e1d3};
test_output[34624:34631] = '{32'h40e38364, 32'h41b9361e, 32'h0, 32'h41d1a763, 32'h429a4ec9, 32'h423490d9, 32'h423f4132, 32'h0};
test_input[34632:34639] = '{32'h40941992, 32'hc1e93fc3, 32'hc28d7876, 32'h40f31cd3, 32'h3f8d8708, 32'hc23982d3, 32'hc29fb090, 32'h42c3675b};
test_output[34632:34639] = '{32'h40941992, 32'h0, 32'h0, 32'h40f31cd3, 32'h3f8d8708, 32'h0, 32'h0, 32'h42c3675b};
test_input[34640:34647] = '{32'hc2a78936, 32'hc2339380, 32'hc21c2d77, 32'h416100b9, 32'h4269a851, 32'hc2658ae8, 32'hc10a83d6, 32'hc2664b69};
test_output[34640:34647] = '{32'h0, 32'h0, 32'h0, 32'h416100b9, 32'h4269a851, 32'h0, 32'h0, 32'h0};
test_input[34648:34655] = '{32'hbfd628c7, 32'h4294df73, 32'h42ae9642, 32'h42bd4040, 32'hc193c5b7, 32'hc28a2d07, 32'h42bea48f, 32'h42b85967};
test_output[34648:34655] = '{32'h0, 32'h4294df73, 32'h42ae9642, 32'h42bd4040, 32'h0, 32'h0, 32'h42bea48f, 32'h42b85967};
test_input[34656:34663] = '{32'h423e3ead, 32'h4291bb61, 32'h42b52c0c, 32'hc0e9af90, 32'hc286e18f, 32'h42abbcc3, 32'h42590c03, 32'hc2614912};
test_output[34656:34663] = '{32'h423e3ead, 32'h4291bb61, 32'h42b52c0c, 32'h0, 32'h0, 32'h42abbcc3, 32'h42590c03, 32'h0};
test_input[34664:34671] = '{32'hc240bc43, 32'hc2b6434c, 32'h41fc059b, 32'h41834da1, 32'h424d62da, 32'hc26c3486, 32'h427935a0, 32'h4210ad1d};
test_output[34664:34671] = '{32'h0, 32'h0, 32'h41fc059b, 32'h41834da1, 32'h424d62da, 32'h0, 32'h427935a0, 32'h4210ad1d};
test_input[34672:34679] = '{32'h417fbf0c, 32'hc1bcb11f, 32'h423cb654, 32'hc2a4c947, 32'h41c7f4ba, 32'h42c1b177, 32'h41ee1a07, 32'hc2954c03};
test_output[34672:34679] = '{32'h417fbf0c, 32'h0, 32'h423cb654, 32'h0, 32'h41c7f4ba, 32'h42c1b177, 32'h41ee1a07, 32'h0};
test_input[34680:34687] = '{32'hc211eec2, 32'hc2be6c5c, 32'hc26e7ab3, 32'hc27a294f, 32'h42c1f9a7, 32'h42937ca3, 32'h42aca21d, 32'h424ea738};
test_output[34680:34687] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42c1f9a7, 32'h42937ca3, 32'h42aca21d, 32'h424ea738};
test_input[34688:34695] = '{32'h429b779d, 32'h40e15eff, 32'hc10416b5, 32'hc0a8b551, 32'hc2842139, 32'h41be9b50, 32'hc296cd98, 32'hc208983f};
test_output[34688:34695] = '{32'h429b779d, 32'h40e15eff, 32'h0, 32'h0, 32'h0, 32'h41be9b50, 32'h0, 32'h0};
test_input[34696:34703] = '{32'h3f8506bd, 32'h41896146, 32'h42897758, 32'h41946c11, 32'hc292005e, 32'hbfd1eef7, 32'h4266064c, 32'hc1d41d2f};
test_output[34696:34703] = '{32'h3f8506bd, 32'h41896146, 32'h42897758, 32'h41946c11, 32'h0, 32'h0, 32'h4266064c, 32'h0};
test_input[34704:34711] = '{32'hc213146c, 32'hc2c01ff3, 32'h4272ebab, 32'h428d0a01, 32'h42014135, 32'h41aaf1ac, 32'h423f524a, 32'hc2465790};
test_output[34704:34711] = '{32'h0, 32'h0, 32'h4272ebab, 32'h428d0a01, 32'h42014135, 32'h41aaf1ac, 32'h423f524a, 32'h0};
test_input[34712:34719] = '{32'hc0e264a4, 32'h427cc3fb, 32'h42bfd2c0, 32'hc29b606d, 32'h42b8db4e, 32'h40260996, 32'h423e98c3, 32'hc21fdcfa};
test_output[34712:34719] = '{32'h0, 32'h427cc3fb, 32'h42bfd2c0, 32'h0, 32'h42b8db4e, 32'h40260996, 32'h423e98c3, 32'h0};
test_input[34720:34727] = '{32'hc19c983f, 32'h42571f19, 32'h42244a2d, 32'hbe8b4e18, 32'h41f22ef9, 32'h42b03fb4, 32'h42c5dda2, 32'h42b4cfd4};
test_output[34720:34727] = '{32'h0, 32'h42571f19, 32'h42244a2d, 32'h0, 32'h41f22ef9, 32'h42b03fb4, 32'h42c5dda2, 32'h42b4cfd4};
test_input[34728:34735] = '{32'h40e076ac, 32'h42bcc80e, 32'hc260ec31, 32'h40c157f8, 32'h42c44ab5, 32'hc2b42787, 32'hc2b7d6fe, 32'hc266a938};
test_output[34728:34735] = '{32'h40e076ac, 32'h42bcc80e, 32'h0, 32'h40c157f8, 32'h42c44ab5, 32'h0, 32'h0, 32'h0};
test_input[34736:34743] = '{32'hc1f68685, 32'hc1ce5775, 32'h42a52ca0, 32'h4274721e, 32'h42ab50d2, 32'h4133dfef, 32'hc22620dc, 32'h4237d5c5};
test_output[34736:34743] = '{32'h0, 32'h0, 32'h42a52ca0, 32'h4274721e, 32'h42ab50d2, 32'h4133dfef, 32'h0, 32'h4237d5c5};
test_input[34744:34751] = '{32'hc2b77072, 32'hc0dd11bb, 32'hc2bb1734, 32'h40831bed, 32'h426e1086, 32'hc2514059, 32'hc2200abb, 32'hc1061dd3};
test_output[34744:34751] = '{32'h0, 32'h0, 32'h0, 32'h40831bed, 32'h426e1086, 32'h0, 32'h0, 32'h0};
test_input[34752:34759] = '{32'h4205d037, 32'h42b89ca2, 32'hc24ef102, 32'h42598587, 32'hc1d8d84b, 32'hc1678bc2, 32'h3f9b352a, 32'hc259a96e};
test_output[34752:34759] = '{32'h4205d037, 32'h42b89ca2, 32'h0, 32'h42598587, 32'h0, 32'h0, 32'h3f9b352a, 32'h0};
test_input[34760:34767] = '{32'hc1a434f1, 32'hc2892f86, 32'hc2bcc68a, 32'h41d9390a, 32'hc2b261ce, 32'h42053667, 32'hc244b4e0, 32'h429d3a6a};
test_output[34760:34767] = '{32'h0, 32'h0, 32'h0, 32'h41d9390a, 32'h0, 32'h42053667, 32'h0, 32'h429d3a6a};
test_input[34768:34775] = '{32'hc2bda9b3, 32'h429970da, 32'hc2c04346, 32'h42be0b2e, 32'hc168df80, 32'h412679e9, 32'h429db92c, 32'h42c10458};
test_output[34768:34775] = '{32'h0, 32'h429970da, 32'h0, 32'h42be0b2e, 32'h0, 32'h412679e9, 32'h429db92c, 32'h42c10458};
test_input[34776:34783] = '{32'h4291c926, 32'h41f2d6c5, 32'h42399f68, 32'hc050ab9d, 32'hc2063dc7, 32'hc1e84087, 32'h42c7d9b3, 32'hc15e681b};
test_output[34776:34783] = '{32'h4291c926, 32'h41f2d6c5, 32'h42399f68, 32'h0, 32'h0, 32'h0, 32'h42c7d9b3, 32'h0};
test_input[34784:34791] = '{32'h41ef5209, 32'hc2bb9521, 32'hc162d0b9, 32'hc28f2ce0, 32'hc28e791d, 32'hc224f1b3, 32'h41eacb09, 32'hc25db360};
test_output[34784:34791] = '{32'h41ef5209, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41eacb09, 32'h0};
test_input[34792:34799] = '{32'hc124fdaf, 32'h414ee726, 32'hc29c0b9f, 32'h41c85e12, 32'hc1e0dbd9, 32'h420bcb31, 32'h428a47e5, 32'hc269e654};
test_output[34792:34799] = '{32'h0, 32'h414ee726, 32'h0, 32'h41c85e12, 32'h0, 32'h420bcb31, 32'h428a47e5, 32'h0};
test_input[34800:34807] = '{32'h42afd96c, 32'hc22cb84d, 32'h42269be0, 32'hc08d0512, 32'h41b2b339, 32'h4285d362, 32'h42aa030b, 32'hc2aaa228};
test_output[34800:34807] = '{32'h42afd96c, 32'h0, 32'h42269be0, 32'h0, 32'h41b2b339, 32'h4285d362, 32'h42aa030b, 32'h0};
test_input[34808:34815] = '{32'hc221c99a, 32'h423df1b1, 32'hc2385ed8, 32'hc24670bb, 32'hc2ab88d5, 32'h4220554d, 32'h42b2e71a, 32'h428111e8};
test_output[34808:34815] = '{32'h0, 32'h423df1b1, 32'h0, 32'h0, 32'h0, 32'h4220554d, 32'h42b2e71a, 32'h428111e8};
test_input[34816:34823] = '{32'hc2c25920, 32'h42bd1121, 32'hc00bdd39, 32'h424aace4, 32'hc22f41e8, 32'hc264c1ad, 32'hc2456574, 32'h40da17f9};
test_output[34816:34823] = '{32'h0, 32'h42bd1121, 32'h0, 32'h424aace4, 32'h0, 32'h0, 32'h0, 32'h40da17f9};
test_input[34824:34831] = '{32'h426eee20, 32'h42bb35e5, 32'h4269fee8, 32'h412c109d, 32'hc07fce5f, 32'hc1c635e2, 32'h41ea4c26, 32'h42018ff4};
test_output[34824:34831] = '{32'h426eee20, 32'h42bb35e5, 32'h4269fee8, 32'h412c109d, 32'h0, 32'h0, 32'h41ea4c26, 32'h42018ff4};
test_input[34832:34839] = '{32'hc25f82c1, 32'hc2702afa, 32'hbf7c3453, 32'h424efc60, 32'h419aa439, 32'hc237c7d0, 32'h4238d3cf, 32'hc29e9b27};
test_output[34832:34839] = '{32'h0, 32'h0, 32'h0, 32'h424efc60, 32'h419aa439, 32'h0, 32'h4238d3cf, 32'h0};
test_input[34840:34847] = '{32'h429c4345, 32'hc2bc916e, 32'hc1a5ed9e, 32'h42598886, 32'hc2c3728f, 32'h41f7a008, 32'h4166e347, 32'h42c52b39};
test_output[34840:34847] = '{32'h429c4345, 32'h0, 32'h0, 32'h42598886, 32'h0, 32'h41f7a008, 32'h4166e347, 32'h42c52b39};
test_input[34848:34855] = '{32'h426455bd, 32'hc2a84f10, 32'h421751e2, 32'hc2068374, 32'hc284d1f8, 32'h41a889ae, 32'h4291641a, 32'h429a49ac};
test_output[34848:34855] = '{32'h426455bd, 32'h0, 32'h421751e2, 32'h0, 32'h0, 32'h41a889ae, 32'h4291641a, 32'h429a49ac};
test_input[34856:34863] = '{32'hc285e9ba, 32'h3d21425a, 32'hc1db6222, 32'h41f12232, 32'hc29eb588, 32'hc22aff82, 32'h41f679bb, 32'hc004dd1c};
test_output[34856:34863] = '{32'h0, 32'h3d21425a, 32'h0, 32'h41f12232, 32'h0, 32'h0, 32'h41f679bb, 32'h0};
test_input[34864:34871] = '{32'hc2a81a82, 32'h4226656c, 32'hc279318c, 32'hc11ebcc6, 32'h428ece00, 32'h41df8a1c, 32'hc21e7d53, 32'hc270f22e};
test_output[34864:34871] = '{32'h0, 32'h4226656c, 32'h0, 32'h0, 32'h428ece00, 32'h41df8a1c, 32'h0, 32'h0};
test_input[34872:34879] = '{32'h41aa0393, 32'h422a0d2f, 32'hc19980b5, 32'hc21519b7, 32'h414ebc9e, 32'h4286a290, 32'h42233da6, 32'hc242c4f5};
test_output[34872:34879] = '{32'h41aa0393, 32'h422a0d2f, 32'h0, 32'h0, 32'h414ebc9e, 32'h4286a290, 32'h42233da6, 32'h0};
test_input[34880:34887] = '{32'hc2a82498, 32'hc2bb38b3, 32'hc2820b85, 32'h428758f2, 32'h4284c48b, 32'hc2443738, 32'h42ac3258, 32'h42be1a46};
test_output[34880:34887] = '{32'h0, 32'h0, 32'h0, 32'h428758f2, 32'h4284c48b, 32'h0, 32'h42ac3258, 32'h42be1a46};
test_input[34888:34895] = '{32'hc18cbdd8, 32'h40e8b3aa, 32'hc2a437f3, 32'hc23bc932, 32'hc2bb8f98, 32'h42c53514, 32'hc1ea2e9e, 32'hc203aa35};
test_output[34888:34895] = '{32'h0, 32'h40e8b3aa, 32'h0, 32'h0, 32'h0, 32'h42c53514, 32'h0, 32'h0};
test_input[34896:34903] = '{32'h41e59b5d, 32'hc2836617, 32'h429093ce, 32'hc1ada648, 32'hc1c9dcd1, 32'h42c5ee94, 32'hc27e6783, 32'hc0a22820};
test_output[34896:34903] = '{32'h41e59b5d, 32'h0, 32'h429093ce, 32'h0, 32'h0, 32'h42c5ee94, 32'h0, 32'h0};
test_input[34904:34911] = '{32'h4244620c, 32'h4202704d, 32'hc1b14e58, 32'h422df2d5, 32'hc2a8eb45, 32'hbfa97904, 32'h4278bf93, 32'hc28f3d0e};
test_output[34904:34911] = '{32'h4244620c, 32'h4202704d, 32'h0, 32'h422df2d5, 32'h0, 32'h0, 32'h4278bf93, 32'h0};
test_input[34912:34919] = '{32'h3fbdca45, 32'h418b2248, 32'h4278d0b7, 32'h41b7ae1f, 32'hc16c7201, 32'h4067423d, 32'h4286dafd, 32'hc13843e9};
test_output[34912:34919] = '{32'h3fbdca45, 32'h418b2248, 32'h4278d0b7, 32'h41b7ae1f, 32'h0, 32'h4067423d, 32'h4286dafd, 32'h0};
test_input[34920:34927] = '{32'hc2ac4e2f, 32'hc2a5ad22, 32'h421627bb, 32'h42b28130, 32'hc220ab5b, 32'hc2a44de3, 32'h41c69260, 32'hbf6b1939};
test_output[34920:34927] = '{32'h0, 32'h0, 32'h421627bb, 32'h42b28130, 32'h0, 32'h0, 32'h41c69260, 32'h0};
test_input[34928:34935] = '{32'h428ddf8d, 32'h41cdf24b, 32'h427f8b01, 32'h41ca06ae, 32'hc262909e, 32'h429a52a4, 32'h422c07e3, 32'h426866bf};
test_output[34928:34935] = '{32'h428ddf8d, 32'h41cdf24b, 32'h427f8b01, 32'h41ca06ae, 32'h0, 32'h429a52a4, 32'h422c07e3, 32'h426866bf};
test_input[34936:34943] = '{32'hc253f35b, 32'hc2930dbf, 32'h409183f8, 32'h413101d5, 32'h424bc648, 32'h41fcdca8, 32'h42ac93b0, 32'h422a2dc6};
test_output[34936:34943] = '{32'h0, 32'h0, 32'h409183f8, 32'h413101d5, 32'h424bc648, 32'h41fcdca8, 32'h42ac93b0, 32'h422a2dc6};
test_input[34944:34951] = '{32'h41be9a11, 32'hc1ae44ba, 32'h42b94a7c, 32'h412da778, 32'hc1d90861, 32'hc2884e56, 32'hc291d20e, 32'hc17bc626};
test_output[34944:34951] = '{32'h41be9a11, 32'h0, 32'h42b94a7c, 32'h412da778, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[34952:34959] = '{32'h429a9bfa, 32'hc2c0f651, 32'hc27e77c6, 32'hc28ded32, 32'hc1b54817, 32'hc28bd01c, 32'h414a6cc1, 32'hc284ccab};
test_output[34952:34959] = '{32'h429a9bfa, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h414a6cc1, 32'h0};
test_input[34960:34967] = '{32'hc1ec67c4, 32'hc1ed00f4, 32'h41c585c7, 32'h41d2ce78, 32'hc2b45db3, 32'hc295dc9a, 32'h4231918c, 32'h413f147a};
test_output[34960:34967] = '{32'h0, 32'h0, 32'h41c585c7, 32'h41d2ce78, 32'h0, 32'h0, 32'h4231918c, 32'h413f147a};
test_input[34968:34975] = '{32'hc20ca99e, 32'h4274b553, 32'hbf234ba0, 32'h4283a0c5, 32'hc1b7d700, 32'h427a2d7b, 32'h42a7abe0, 32'h42553798};
test_output[34968:34975] = '{32'h0, 32'h4274b553, 32'h0, 32'h4283a0c5, 32'h0, 32'h427a2d7b, 32'h42a7abe0, 32'h42553798};
test_input[34976:34983] = '{32'h42b02555, 32'hc2846fbb, 32'h403e0dc0, 32'hc13c2135, 32'h425a32bb, 32'hc2bb5517, 32'h41fcb71e, 32'h4289d5c0};
test_output[34976:34983] = '{32'h42b02555, 32'h0, 32'h403e0dc0, 32'h0, 32'h425a32bb, 32'h0, 32'h41fcb71e, 32'h4289d5c0};
test_input[34984:34991] = '{32'hc0a4bcaa, 32'hc1ca7b00, 32'hc175817e, 32'h427f9212, 32'hc064ef1f, 32'h420d85f4, 32'hc256689d, 32'h4288f4b9};
test_output[34984:34991] = '{32'h0, 32'h0, 32'h0, 32'h427f9212, 32'h0, 32'h420d85f4, 32'h0, 32'h4288f4b9};
test_input[34992:34999] = '{32'hc2b207af, 32'h40c0f2d7, 32'h41346bfb, 32'h41c0664d, 32'h4232e70b, 32'h41bbeea5, 32'h422257e8, 32'hc2a75675};
test_output[34992:34999] = '{32'h0, 32'h40c0f2d7, 32'h41346bfb, 32'h41c0664d, 32'h4232e70b, 32'h41bbeea5, 32'h422257e8, 32'h0};
test_input[35000:35007] = '{32'h413e5d5c, 32'h41855fbf, 32'h420cdad4, 32'hc23ea9c3, 32'hc26514ec, 32'hc2a4f811, 32'h4291e502, 32'hc20a4c61};
test_output[35000:35007] = '{32'h413e5d5c, 32'h41855fbf, 32'h420cdad4, 32'h0, 32'h0, 32'h0, 32'h4291e502, 32'h0};
test_input[35008:35015] = '{32'h428244d7, 32'hc2b67301, 32'hc2170efd, 32'hc2268c35, 32'h427d9f3b, 32'hc20bdb28, 32'h3f3c1363, 32'h413016ab};
test_output[35008:35015] = '{32'h428244d7, 32'h0, 32'h0, 32'h0, 32'h427d9f3b, 32'h0, 32'h3f3c1363, 32'h413016ab};
test_input[35016:35023] = '{32'h41885064, 32'hc2176c29, 32'h42b0394a, 32'h425f566a, 32'h423cfc8f, 32'hc2a21619, 32'hc286966c, 32'hc2316419};
test_output[35016:35023] = '{32'h41885064, 32'h0, 32'h42b0394a, 32'h425f566a, 32'h423cfc8f, 32'h0, 32'h0, 32'h0};
test_input[35024:35031] = '{32'hc2c2b187, 32'h4129101e, 32'hc2a90435, 32'hc27151dd, 32'hc2986f3a, 32'hc2a93211, 32'hc1a37b61, 32'hc2c6ac9c};
test_output[35024:35031] = '{32'h0, 32'h4129101e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35032:35039] = '{32'hc2103a9a, 32'h428d40de, 32'h42111017, 32'hc28b27d2, 32'hc2062910, 32'hc285cc97, 32'hc2c3cd67, 32'h4219336d};
test_output[35032:35039] = '{32'h0, 32'h428d40de, 32'h42111017, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4219336d};
test_input[35040:35047] = '{32'h42a24b96, 32'hc2ad3d1b, 32'hc21a2260, 32'h41daa6d7, 32'hc1932ada, 32'hc13c1ee7, 32'hc23e70f2, 32'hc1ee7d5a};
test_output[35040:35047] = '{32'h42a24b96, 32'h0, 32'h0, 32'h41daa6d7, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35048:35055] = '{32'hc1fb75c1, 32'h4222cf84, 32'hc278ad5f, 32'h4250fcc9, 32'h42007186, 32'hc1a63a6a, 32'h4290971c, 32'h41ee5310};
test_output[35048:35055] = '{32'h0, 32'h4222cf84, 32'h0, 32'h4250fcc9, 32'h42007186, 32'h0, 32'h4290971c, 32'h41ee5310};
test_input[35056:35063] = '{32'hc1b62232, 32'hc1281339, 32'h408e9bdc, 32'hc2742487, 32'h429243fe, 32'h42ae1a15, 32'hc2bda55a, 32'h427693be};
test_output[35056:35063] = '{32'h0, 32'h0, 32'h408e9bdc, 32'h0, 32'h429243fe, 32'h42ae1a15, 32'h0, 32'h427693be};
test_input[35064:35071] = '{32'h41acf993, 32'h429a93d0, 32'h4291dc9e, 32'h428b06fa, 32'h420e37dd, 32'hc1975c22, 32'h40b34376, 32'hc2208073};
test_output[35064:35071] = '{32'h41acf993, 32'h429a93d0, 32'h4291dc9e, 32'h428b06fa, 32'h420e37dd, 32'h0, 32'h40b34376, 32'h0};
test_input[35072:35079] = '{32'h428d2f52, 32'h4241c693, 32'h42a33e79, 32'hc29cbf0c, 32'h42039322, 32'h424daf0e, 32'hc282b167, 32'hc27b81d8};
test_output[35072:35079] = '{32'h428d2f52, 32'h4241c693, 32'h42a33e79, 32'h0, 32'h42039322, 32'h424daf0e, 32'h0, 32'h0};
test_input[35080:35087] = '{32'hc293e72a, 32'h415fa931, 32'hc24529cf, 32'hc0faffc4, 32'hc2c3c106, 32'h42a02baa, 32'h3fa637b2, 32'hc29442d6};
test_output[35080:35087] = '{32'h0, 32'h415fa931, 32'h0, 32'h0, 32'h0, 32'h42a02baa, 32'h3fa637b2, 32'h0};
test_input[35088:35095] = '{32'h4201be7c, 32'hc27d7f9b, 32'h421e3f03, 32'h400a4539, 32'hc25180cd, 32'hc2724904, 32'h422a4d08, 32'h41875b49};
test_output[35088:35095] = '{32'h4201be7c, 32'h0, 32'h421e3f03, 32'h400a4539, 32'h0, 32'h0, 32'h422a4d08, 32'h41875b49};
test_input[35096:35103] = '{32'h415d7e3f, 32'hc298fe12, 32'hc2241935, 32'h41fbc851, 32'h421e593f, 32'hc29ef056, 32'hc2398f83, 32'h41fb56f0};
test_output[35096:35103] = '{32'h415d7e3f, 32'h0, 32'h0, 32'h41fbc851, 32'h421e593f, 32'h0, 32'h0, 32'h41fb56f0};
test_input[35104:35111] = '{32'hc2369625, 32'hc176ee02, 32'h429234c0, 32'h3f0935c1, 32'hc2b9a095, 32'hc1bcde21, 32'hc25b903a, 32'hc2a51360};
test_output[35104:35111] = '{32'h0, 32'h0, 32'h429234c0, 32'h3f0935c1, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35112:35119] = '{32'h422ebe15, 32'h426ab6bf, 32'h40fd38b8, 32'h428ebc50, 32'hc29b1b20, 32'hc1aeb98b, 32'h40c8a5c6, 32'h429d0207};
test_output[35112:35119] = '{32'h422ebe15, 32'h426ab6bf, 32'h40fd38b8, 32'h428ebc50, 32'h0, 32'h0, 32'h40c8a5c6, 32'h429d0207};
test_input[35120:35127] = '{32'h419494e3, 32'hc18ea816, 32'h42859ffc, 32'h4114d13f, 32'hc135cb3e, 32'h424be50d, 32'hc028f71f, 32'hc28c24e4};
test_output[35120:35127] = '{32'h419494e3, 32'h0, 32'h42859ffc, 32'h4114d13f, 32'h0, 32'h424be50d, 32'h0, 32'h0};
test_input[35128:35135] = '{32'hc2a9d68c, 32'h4282f820, 32'h42a5a1f3, 32'hc25e2b91, 32'h425a401e, 32'hc18c8574, 32'hc08b86bb, 32'h42a6cf12};
test_output[35128:35135] = '{32'h0, 32'h4282f820, 32'h42a5a1f3, 32'h0, 32'h425a401e, 32'h0, 32'h0, 32'h42a6cf12};
test_input[35136:35143] = '{32'h418c1f38, 32'hc284ec8f, 32'h42a9a2ac, 32'hc28e9fb1, 32'h4293f71f, 32'hc215be1c, 32'hc1973716, 32'h413562a0};
test_output[35136:35143] = '{32'h418c1f38, 32'h0, 32'h42a9a2ac, 32'h0, 32'h4293f71f, 32'h0, 32'h0, 32'h413562a0};
test_input[35144:35151] = '{32'hc25b7eb8, 32'h42170d2e, 32'hc249df4a, 32'h421b9f30, 32'hc29ef172, 32'h407aad2f, 32'hc2986f93, 32'h429520f1};
test_output[35144:35151] = '{32'h0, 32'h42170d2e, 32'h0, 32'h421b9f30, 32'h0, 32'h407aad2f, 32'h0, 32'h429520f1};
test_input[35152:35159] = '{32'h427d2919, 32'hc2aaab1b, 32'h429bdb27, 32'h425f96a1, 32'hc25758de, 32'hc10ee4a0, 32'h41ce4a6f, 32'h41891a32};
test_output[35152:35159] = '{32'h427d2919, 32'h0, 32'h429bdb27, 32'h425f96a1, 32'h0, 32'h0, 32'h41ce4a6f, 32'h41891a32};
test_input[35160:35167] = '{32'h42be7b71, 32'hc234d4a4, 32'hc275c5d2, 32'hc29d32a1, 32'hc29f1a03, 32'h4242c634, 32'h425fae62, 32'h4201b0d5};
test_output[35160:35167] = '{32'h42be7b71, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4242c634, 32'h425fae62, 32'h4201b0d5};
test_input[35168:35175] = '{32'h429dbf2e, 32'h42abb2c0, 32'hc28564b2, 32'h4298dafb, 32'h42c796a9, 32'h428f95c5, 32'h4298b8b3, 32'hc1204798};
test_output[35168:35175] = '{32'h429dbf2e, 32'h42abb2c0, 32'h0, 32'h4298dafb, 32'h42c796a9, 32'h428f95c5, 32'h4298b8b3, 32'h0};
test_input[35176:35183] = '{32'h425725d7, 32'hbfb921a0, 32'h42247717, 32'hc1add4e3, 32'hc2b4b3ac, 32'hc249f9fd, 32'hc07ebb1d, 32'h42327087};
test_output[35176:35183] = '{32'h425725d7, 32'h0, 32'h42247717, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42327087};
test_input[35184:35191] = '{32'hc292c8b1, 32'hc2256802, 32'hc18c2079, 32'hc2465790, 32'hc289270c, 32'hc08c4503, 32'hc2bd06d6, 32'hc1029a33};
test_output[35184:35191] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35192:35199] = '{32'hc0f5417e, 32'h42947ef1, 32'hc1e3ae35, 32'hc1214dab, 32'hc28ae524, 32'h423fa000, 32'h41b55a5f, 32'h42a29bc1};
test_output[35192:35199] = '{32'h0, 32'h42947ef1, 32'h0, 32'h0, 32'h0, 32'h423fa000, 32'h41b55a5f, 32'h42a29bc1};
test_input[35200:35207] = '{32'hc1f34d9a, 32'hc164566f, 32'h429e3f63, 32'h42b81eaf, 32'h41fac0ec, 32'hc2802b33, 32'hc09ec746, 32'hc18069ad};
test_output[35200:35207] = '{32'h0, 32'h0, 32'h429e3f63, 32'h42b81eaf, 32'h41fac0ec, 32'h0, 32'h0, 32'h0};
test_input[35208:35215] = '{32'hc1e738b0, 32'h41c76918, 32'h4297ba9a, 32'h428cf0f6, 32'h42167b0c, 32'h4285ca88, 32'h41bae299, 32'h41667655};
test_output[35208:35215] = '{32'h0, 32'h41c76918, 32'h4297ba9a, 32'h428cf0f6, 32'h42167b0c, 32'h4285ca88, 32'h41bae299, 32'h41667655};
test_input[35216:35223] = '{32'hc23f7906, 32'hc271adbf, 32'hc2b23122, 32'h425bb24f, 32'hc2b28d86, 32'hc0a1f972, 32'hc294b49f, 32'h41568e79};
test_output[35216:35223] = '{32'h0, 32'h0, 32'h0, 32'h425bb24f, 32'h0, 32'h0, 32'h0, 32'h41568e79};
test_input[35224:35231] = '{32'h429697cc, 32'h42877a53, 32'h414bfd16, 32'h423de273, 32'hc258f04f, 32'h41afcbcc, 32'h42c3c825, 32'hc1848244};
test_output[35224:35231] = '{32'h429697cc, 32'h42877a53, 32'h414bfd16, 32'h423de273, 32'h0, 32'h41afcbcc, 32'h42c3c825, 32'h0};
test_input[35232:35239] = '{32'h420f16cf, 32'h41412f1e, 32'hc2a23a9b, 32'h4227a100, 32'hc2a976b2, 32'h4230e465, 32'h422e1704, 32'hc210deca};
test_output[35232:35239] = '{32'h420f16cf, 32'h41412f1e, 32'h0, 32'h4227a100, 32'h0, 32'h4230e465, 32'h422e1704, 32'h0};
test_input[35240:35247] = '{32'h42ab3cc5, 32'h41f716bc, 32'h4280d227, 32'hc29bd6b3, 32'h42060ecf, 32'h42274cad, 32'hc24fd247, 32'hc1fb84bd};
test_output[35240:35247] = '{32'h42ab3cc5, 32'h41f716bc, 32'h4280d227, 32'h0, 32'h42060ecf, 32'h42274cad, 32'h0, 32'h0};
test_input[35248:35255] = '{32'h41a90968, 32'hc259c9c1, 32'h42bbe0f9, 32'hc1c53238, 32'hc288bbb3, 32'hc2691a7f, 32'h422012cf, 32'hc283acf6};
test_output[35248:35255] = '{32'h41a90968, 32'h0, 32'h42bbe0f9, 32'h0, 32'h0, 32'h0, 32'h422012cf, 32'h0};
test_input[35256:35263] = '{32'hc0c43154, 32'h3fb15482, 32'h41cbab84, 32'hc2b4088e, 32'h42bb8f5d, 32'hc252c463, 32'h418830cd, 32'hc211c617};
test_output[35256:35263] = '{32'h0, 32'h3fb15482, 32'h41cbab84, 32'h0, 32'h42bb8f5d, 32'h0, 32'h418830cd, 32'h0};
test_input[35264:35271] = '{32'h424207a0, 32'hc1f03891, 32'hc27bb539, 32'hc23a5f60, 32'hc2668668, 32'hc282ae8f, 32'h422ccc81, 32'hc246e79b};
test_output[35264:35271] = '{32'h424207a0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h422ccc81, 32'h0};
test_input[35272:35279] = '{32'h41817d64, 32'h422fd68a, 32'hc0f44694, 32'hc21a8238, 32'h42c0e142, 32'h42a05839, 32'hc2b639d8, 32'h4186163a};
test_output[35272:35279] = '{32'h41817d64, 32'h422fd68a, 32'h0, 32'h0, 32'h42c0e142, 32'h42a05839, 32'h0, 32'h4186163a};
test_input[35280:35287] = '{32'h42b25415, 32'hc2911c4b, 32'hc0820893, 32'hc2a40c52, 32'h4245b866, 32'hc179a2d5, 32'hc2b35eea, 32'hc1fffb19};
test_output[35280:35287] = '{32'h42b25415, 32'h0, 32'h0, 32'h0, 32'h4245b866, 32'h0, 32'h0, 32'h0};
test_input[35288:35295] = '{32'hc28a4dfd, 32'hc253aa90, 32'hc2977a9f, 32'h42435034, 32'h418dced9, 32'hc159521b, 32'hc2887f28, 32'h416a4f42};
test_output[35288:35295] = '{32'h0, 32'h0, 32'h0, 32'h42435034, 32'h418dced9, 32'h0, 32'h0, 32'h416a4f42};
test_input[35296:35303] = '{32'hc2918ba7, 32'hc264ed43, 32'hc2c57c49, 32'hc296123d, 32'h402512c7, 32'hc291e8cd, 32'h42ab0287, 32'h429e4229};
test_output[35296:35303] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h402512c7, 32'h0, 32'h42ab0287, 32'h429e4229};
test_input[35304:35311] = '{32'h414f78e7, 32'h42c1a5e7, 32'hc2664a17, 32'hc1f4935d, 32'h42a1f88d, 32'hc181659d, 32'h427fd1c2, 32'hc28cbe09};
test_output[35304:35311] = '{32'h414f78e7, 32'h42c1a5e7, 32'h0, 32'h0, 32'h42a1f88d, 32'h0, 32'h427fd1c2, 32'h0};
test_input[35312:35319] = '{32'hc2c4ccb9, 32'h425e9817, 32'hc036c90b, 32'hc278c39b, 32'hc29cc995, 32'h4171657d, 32'h4256e5fa, 32'h42c1d924};
test_output[35312:35319] = '{32'h0, 32'h425e9817, 32'h0, 32'h0, 32'h0, 32'h4171657d, 32'h4256e5fa, 32'h42c1d924};
test_input[35320:35327] = '{32'hc271f63c, 32'hc211e3ff, 32'h41fb397e, 32'hc090746b, 32'hc28fd237, 32'h428c9e86, 32'hc211c51c, 32'h427c89c4};
test_output[35320:35327] = '{32'h0, 32'h0, 32'h41fb397e, 32'h0, 32'h0, 32'h428c9e86, 32'h0, 32'h427c89c4};
test_input[35328:35335] = '{32'h411f9306, 32'hc287e7eb, 32'h4200df3c, 32'h42210ecc, 32'h42c28644, 32'h41025b00, 32'hc2a433fb, 32'h423f85b5};
test_output[35328:35335] = '{32'h411f9306, 32'h0, 32'h4200df3c, 32'h42210ecc, 32'h42c28644, 32'h41025b00, 32'h0, 32'h423f85b5};
test_input[35336:35343] = '{32'hbe51c87a, 32'h421e7fbf, 32'hc275cae7, 32'h4291fde2, 32'h42487a22, 32'hc27cbc3a, 32'hc29e6f2d, 32'hc1daafe6};
test_output[35336:35343] = '{32'h0, 32'h421e7fbf, 32'h0, 32'h4291fde2, 32'h42487a22, 32'h0, 32'h0, 32'h0};
test_input[35344:35351] = '{32'hc148b382, 32'hc27d2f25, 32'hc29993af, 32'h429a0888, 32'h41cdc4ff, 32'h41700e23, 32'hc27cda10, 32'hc2954c7d};
test_output[35344:35351] = '{32'h0, 32'h0, 32'h0, 32'h429a0888, 32'h41cdc4ff, 32'h41700e23, 32'h0, 32'h0};
test_input[35352:35359] = '{32'h4233f31e, 32'h428ce780, 32'hc2b19694, 32'hc2169c71, 32'h4285f67a, 32'hc27967e0, 32'hc20e0a23, 32'h40c9779d};
test_output[35352:35359] = '{32'h4233f31e, 32'h428ce780, 32'h0, 32'h0, 32'h4285f67a, 32'h0, 32'h0, 32'h40c9779d};
test_input[35360:35367] = '{32'hc21d02d7, 32'h41bc2591, 32'h41b71b57, 32'hc2751460, 32'hc2859078, 32'hc2457769, 32'hc11b8c0b, 32'h42401f82};
test_output[35360:35367] = '{32'h0, 32'h41bc2591, 32'h41b71b57, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42401f82};
test_input[35368:35375] = '{32'hc21622f2, 32'hc27fa676, 32'hc25803bc, 32'h42170a8f, 32'h4083f3d8, 32'hc1f11f23, 32'hc2c6afce, 32'hc25128af};
test_output[35368:35375] = '{32'h0, 32'h0, 32'h0, 32'h42170a8f, 32'h4083f3d8, 32'h0, 32'h0, 32'h0};
test_input[35376:35383] = '{32'h428565a3, 32'h41d1c76b, 32'hc20c8533, 32'h41ccc5d4, 32'hc28c4278, 32'h42360c5d, 32'hc207baeb, 32'hc2aa9acf};
test_output[35376:35383] = '{32'h428565a3, 32'h41d1c76b, 32'h0, 32'h41ccc5d4, 32'h0, 32'h42360c5d, 32'h0, 32'h0};
test_input[35384:35391] = '{32'hc2a0d3ef, 32'h42459b71, 32'h421fadcb, 32'hc1913d1a, 32'hc21c9ea0, 32'hc1d6c471, 32'hc2588c03, 32'hbfcf3be3};
test_output[35384:35391] = '{32'h0, 32'h42459b71, 32'h421fadcb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35392:35399] = '{32'h40fe8d75, 32'h427f039e, 32'hc13b65cc, 32'h428c6a20, 32'h40b7e44f, 32'h4294ce03, 32'hc2964ad5, 32'hc26db715};
test_output[35392:35399] = '{32'h40fe8d75, 32'h427f039e, 32'h0, 32'h428c6a20, 32'h40b7e44f, 32'h4294ce03, 32'h0, 32'h0};
test_input[35400:35407] = '{32'hc22ad134, 32'hc2873583, 32'h42226477, 32'h429ef369, 32'hc23bf0d3, 32'h428c11c7, 32'hc1658c73, 32'hc2b3759a};
test_output[35400:35407] = '{32'h0, 32'h0, 32'h42226477, 32'h429ef369, 32'h0, 32'h428c11c7, 32'h0, 32'h0};
test_input[35408:35415] = '{32'h41d7de50, 32'h42827c57, 32'hc1a9d4fb, 32'h420284e3, 32'hc2120d94, 32'h425fd2b4, 32'h42737fcf, 32'h4285bd5b};
test_output[35408:35415] = '{32'h41d7de50, 32'h42827c57, 32'h0, 32'h420284e3, 32'h0, 32'h425fd2b4, 32'h42737fcf, 32'h4285bd5b};
test_input[35416:35423] = '{32'h41a37473, 32'h42c3a0de, 32'h42b27117, 32'h4165a172, 32'hc26c2685, 32'hc2979818, 32'hc2077c6c, 32'h41502e24};
test_output[35416:35423] = '{32'h41a37473, 32'h42c3a0de, 32'h42b27117, 32'h4165a172, 32'h0, 32'h0, 32'h0, 32'h41502e24};
test_input[35424:35431] = '{32'hc1c9c263, 32'hc233975b, 32'hc2b1577c, 32'h42b26290, 32'h3ea80a20, 32'h42a44580, 32'h42318427, 32'hc2203883};
test_output[35424:35431] = '{32'h0, 32'h0, 32'h0, 32'h42b26290, 32'h3ea80a20, 32'h42a44580, 32'h42318427, 32'h0};
test_input[35432:35439] = '{32'hc19fa18b, 32'hc2104bd8, 32'hc1e21a2d, 32'h41b3fa7d, 32'h42a0fdc5, 32'hc274dc98, 32'hc2bda0dc, 32'h425cb9ce};
test_output[35432:35439] = '{32'h0, 32'h0, 32'h0, 32'h41b3fa7d, 32'h42a0fdc5, 32'h0, 32'h0, 32'h425cb9ce};
test_input[35440:35447] = '{32'h414f6e5b, 32'hc2ae9549, 32'h42a22a1e, 32'hc27d0efd, 32'h426a7843, 32'h40e5bb4c, 32'h42bcd843, 32'hc2a889b4};
test_output[35440:35447] = '{32'h414f6e5b, 32'h0, 32'h42a22a1e, 32'h0, 32'h426a7843, 32'h40e5bb4c, 32'h42bcd843, 32'h0};
test_input[35448:35455] = '{32'h428740cf, 32'hc0cca559, 32'h426139b0, 32'h4265d6ef, 32'h428a0001, 32'h41ccf21b, 32'hc2990161, 32'hc1946910};
test_output[35448:35455] = '{32'h428740cf, 32'h0, 32'h426139b0, 32'h4265d6ef, 32'h428a0001, 32'h41ccf21b, 32'h0, 32'h0};
test_input[35456:35463] = '{32'hc2152c67, 32'h4218e69c, 32'hc288d230, 32'h429d5b61, 32'h42821deb, 32'hc203efd0, 32'hc26bd354, 32'hc0aabf44};
test_output[35456:35463] = '{32'h0, 32'h4218e69c, 32'h0, 32'h429d5b61, 32'h42821deb, 32'h0, 32'h0, 32'h0};
test_input[35464:35471] = '{32'h408aac3b, 32'h420fb48d, 32'hc296a938, 32'hc2a4965f, 32'hc28104e0, 32'hc2862be2, 32'h41f71398, 32'h42954b4f};
test_output[35464:35471] = '{32'h408aac3b, 32'h420fb48d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41f71398, 32'h42954b4f};
test_input[35472:35479] = '{32'h40fefaed, 32'hc27002e0, 32'h429d832d, 32'h42b74306, 32'hc2c0a25f, 32'h428d5c17, 32'hc22e3f39, 32'h41fa6250};
test_output[35472:35479] = '{32'h40fefaed, 32'h0, 32'h429d832d, 32'h42b74306, 32'h0, 32'h428d5c17, 32'h0, 32'h41fa6250};
test_input[35480:35487] = '{32'hc203366f, 32'h428994f7, 32'hc285bcd2, 32'h425270d8, 32'h4278c2f7, 32'h42be3279, 32'h415fda83, 32'h426a79aa};
test_output[35480:35487] = '{32'h0, 32'h428994f7, 32'h0, 32'h425270d8, 32'h4278c2f7, 32'h42be3279, 32'h415fda83, 32'h426a79aa};
test_input[35488:35495] = '{32'hc1485aed, 32'h4289971b, 32'h405692b1, 32'hc28cc4b0, 32'h4156e65c, 32'h424b4f12, 32'hc2a8852b, 32'hc2649f4f};
test_output[35488:35495] = '{32'h0, 32'h4289971b, 32'h405692b1, 32'h0, 32'h4156e65c, 32'h424b4f12, 32'h0, 32'h0};
test_input[35496:35503] = '{32'hc1d36bbc, 32'hc1c75fbb, 32'hc1b01f22, 32'h4278db3c, 32'h4226438e, 32'hc298381b, 32'h42b14d18, 32'hc29372be};
test_output[35496:35503] = '{32'h0, 32'h0, 32'h0, 32'h4278db3c, 32'h4226438e, 32'h0, 32'h42b14d18, 32'h0};
test_input[35504:35511] = '{32'h4171f16d, 32'h425b409b, 32'h41bd36b7, 32'h4273fa72, 32'hc2c378f1, 32'h429674a4, 32'h408bcfa7, 32'hc280ec80};
test_output[35504:35511] = '{32'h4171f16d, 32'h425b409b, 32'h41bd36b7, 32'h4273fa72, 32'h0, 32'h429674a4, 32'h408bcfa7, 32'h0};
test_input[35512:35519] = '{32'hc13d389b, 32'h4234b397, 32'h41eaa6a9, 32'hc2a8a340, 32'hc22182dd, 32'hc21cdb64, 32'h42bb80f7, 32'h42939a14};
test_output[35512:35519] = '{32'h0, 32'h4234b397, 32'h41eaa6a9, 32'h0, 32'h0, 32'h0, 32'h42bb80f7, 32'h42939a14};
test_input[35520:35527] = '{32'hc26cd506, 32'hc26c188a, 32'h42b6e5d7, 32'h42ab5048, 32'h424029a4, 32'hc1a30860, 32'hc1dcd1df, 32'h429ee497};
test_output[35520:35527] = '{32'h0, 32'h0, 32'h42b6e5d7, 32'h42ab5048, 32'h424029a4, 32'h0, 32'h0, 32'h429ee497};
test_input[35528:35535] = '{32'h429edb8b, 32'hc25a9c02, 32'hc2b8e4b2, 32'h41c78679, 32'h42163181, 32'hc2a0f4b4, 32'hc29285c1, 32'h41d55a09};
test_output[35528:35535] = '{32'h429edb8b, 32'h0, 32'h0, 32'h41c78679, 32'h42163181, 32'h0, 32'h0, 32'h41d55a09};
test_input[35536:35543] = '{32'h419afbed, 32'h4264a8e0, 32'h42b84392, 32'h41b334b6, 32'h42bb7a13, 32'hc1aae762, 32'h41826477, 32'h400d6dca};
test_output[35536:35543] = '{32'h419afbed, 32'h4264a8e0, 32'h42b84392, 32'h41b334b6, 32'h42bb7a13, 32'h0, 32'h41826477, 32'h400d6dca};
test_input[35544:35551] = '{32'h420b50ce, 32'h42843837, 32'h4297ab86, 32'hc2bdb720, 32'hc287ae7e, 32'h404f156f, 32'h426d2d2b, 32'hc1db47f2};
test_output[35544:35551] = '{32'h420b50ce, 32'h42843837, 32'h4297ab86, 32'h0, 32'h0, 32'h404f156f, 32'h426d2d2b, 32'h0};
test_input[35552:35559] = '{32'h421485d9, 32'hc219c71a, 32'hc2a457f6, 32'h41fdad7d, 32'hc25da999, 32'h42855359, 32'hc2bffa85, 32'hc23628c8};
test_output[35552:35559] = '{32'h421485d9, 32'h0, 32'h0, 32'h41fdad7d, 32'h0, 32'h42855359, 32'h0, 32'h0};
test_input[35560:35567] = '{32'h40629f18, 32'h4299bba9, 32'hc18ba037, 32'hc2281bde, 32'h4285a403, 32'hc14012ec, 32'hc1db9045, 32'h407ad79c};
test_output[35560:35567] = '{32'h40629f18, 32'h4299bba9, 32'h0, 32'h0, 32'h4285a403, 32'h0, 32'h0, 32'h407ad79c};
test_input[35568:35575] = '{32'h41db441c, 32'h4204e855, 32'hc0f108f4, 32'hc2b38785, 32'hc2724a2c, 32'hc1d2bee6, 32'hc285a01c, 32'hbf0fa596};
test_output[35568:35575] = '{32'h41db441c, 32'h4204e855, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35576:35583] = '{32'hc14c3a39, 32'hc22fda65, 32'h424c0ba7, 32'hc2ad72db, 32'h42619f7f, 32'hc18f2825, 32'h4218eaf3, 32'hc29781ab};
test_output[35576:35583] = '{32'h0, 32'h0, 32'h424c0ba7, 32'h0, 32'h42619f7f, 32'h0, 32'h4218eaf3, 32'h0};
test_input[35584:35591] = '{32'h4283f890, 32'h421ac0b4, 32'h410ef9de, 32'h413c3af3, 32'h42838b6b, 32'hc0ccb212, 32'hc2810a9c, 32'hc29a4501};
test_output[35584:35591] = '{32'h4283f890, 32'h421ac0b4, 32'h410ef9de, 32'h413c3af3, 32'h42838b6b, 32'h0, 32'h0, 32'h0};
test_input[35592:35599] = '{32'hc2c02e76, 32'hc21042f5, 32'hc23135e2, 32'hc177f953, 32'hc20c133d, 32'hc2999210, 32'hc29a4664, 32'h423ebc5e};
test_output[35592:35599] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423ebc5e};
test_input[35600:35607] = '{32'h4256f246, 32'hbe17a9df, 32'h4293b29b, 32'h42afe358, 32'hc2c73f0c, 32'h42732846, 32'hc187283f, 32'h412bc059};
test_output[35600:35607] = '{32'h4256f246, 32'h0, 32'h4293b29b, 32'h42afe358, 32'h0, 32'h42732846, 32'h0, 32'h412bc059};
test_input[35608:35615] = '{32'hc29ad99b, 32'hc18761f7, 32'h429bf621, 32'hc1870bd9, 32'h4294e6ea, 32'hc24c71db, 32'hc280e117, 32'hc2bcbb8d};
test_output[35608:35615] = '{32'h0, 32'h0, 32'h429bf621, 32'h0, 32'h4294e6ea, 32'h0, 32'h0, 32'h0};
test_input[35616:35623] = '{32'h42b53434, 32'hc284d711, 32'hc2a731d8, 32'hc2b830bb, 32'h41f065f6, 32'hc2a5747b, 32'hc1caa9c1, 32'h424843b9};
test_output[35616:35623] = '{32'h42b53434, 32'h0, 32'h0, 32'h0, 32'h41f065f6, 32'h0, 32'h0, 32'h424843b9};
test_input[35624:35631] = '{32'hc281c0fe, 32'h4299d350, 32'hc28e5b61, 32'h42c31e38, 32'hc23255c8, 32'hc1086629, 32'hc2ac7ceb, 32'h428102a3};
test_output[35624:35631] = '{32'h0, 32'h4299d350, 32'h0, 32'h42c31e38, 32'h0, 32'h0, 32'h0, 32'h428102a3};
test_input[35632:35639] = '{32'hc2c7a82c, 32'h4295b340, 32'hc29f2c81, 32'hc216e9b0, 32'hc0d2f3c9, 32'hc1f8d6a6, 32'h424aba08, 32'h419dccac};
test_output[35632:35639] = '{32'h0, 32'h4295b340, 32'h0, 32'h0, 32'h0, 32'h0, 32'h424aba08, 32'h419dccac};
test_input[35640:35647] = '{32'hc241cfb9, 32'h421d89ea, 32'h42984427, 32'hc216f6bd, 32'h42bb5ad0, 32'h429d7ad4, 32'hc217d7ed, 32'h411c2062};
test_output[35640:35647] = '{32'h0, 32'h421d89ea, 32'h42984427, 32'h0, 32'h42bb5ad0, 32'h429d7ad4, 32'h0, 32'h411c2062};
test_input[35648:35655] = '{32'hc212db36, 32'hc1649dae, 32'hc0ba424c, 32'h42c469ae, 32'hc224df9b, 32'h40fbab1a, 32'hc2754a0c, 32'hc1e9ec2e};
test_output[35648:35655] = '{32'h0, 32'h0, 32'h0, 32'h42c469ae, 32'h0, 32'h40fbab1a, 32'h0, 32'h0};
test_input[35656:35663] = '{32'h4210a2a3, 32'h4298f71b, 32'hc27633d6, 32'hc22512a4, 32'hc29d6d74, 32'hc2113196, 32'hc294ed5f, 32'hc1f2e3ee};
test_output[35656:35663] = '{32'h4210a2a3, 32'h4298f71b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35664:35671] = '{32'hbfc04008, 32'hc1c0e9dd, 32'hc0b53fdc, 32'hc1c591a4, 32'hc21764c9, 32'hc28925e5, 32'h42742cb8, 32'h420f6298};
test_output[35664:35671] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42742cb8, 32'h420f6298};
test_input[35672:35679] = '{32'hc27ca511, 32'hc28c79e2, 32'hc277e9c7, 32'h40956f24, 32'h42919c33, 32'h42a49807, 32'hc1b9daaf, 32'h42b7ec2a};
test_output[35672:35679] = '{32'h0, 32'h0, 32'h0, 32'h40956f24, 32'h42919c33, 32'h42a49807, 32'h0, 32'h42b7ec2a};
test_input[35680:35687] = '{32'hc1b2f2c6, 32'hc29b281f, 32'hc00a5a91, 32'h41b7349a, 32'hc2a85ec1, 32'hc2534f67, 32'hc20f7117, 32'hc2a126b8};
test_output[35680:35687] = '{32'h0, 32'h0, 32'h0, 32'h41b7349a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35688:35695] = '{32'h4224d267, 32'hc296a21c, 32'hc1ca1136, 32'h429d9ab7, 32'hc188756d, 32'hc24cc6a6, 32'h427ae08b, 32'hc2b631d5};
test_output[35688:35695] = '{32'h4224d267, 32'h0, 32'h0, 32'h429d9ab7, 32'h0, 32'h0, 32'h427ae08b, 32'h0};
test_input[35696:35703] = '{32'hc2bc7023, 32'hc2b15600, 32'h41b92c18, 32'hc298e832, 32'h420ac2c7, 32'h41a52fd8, 32'h42984fae, 32'hc299e8d0};
test_output[35696:35703] = '{32'h0, 32'h0, 32'h41b92c18, 32'h0, 32'h420ac2c7, 32'h41a52fd8, 32'h42984fae, 32'h0};
test_input[35704:35711] = '{32'hc1f8892a, 32'h42bd9b3b, 32'h41a09db7, 32'h42302173, 32'hc2b229f6, 32'h42b01917, 32'hbfbd3a0f, 32'hc1fd55f9};
test_output[35704:35711] = '{32'h0, 32'h42bd9b3b, 32'h41a09db7, 32'h42302173, 32'h0, 32'h42b01917, 32'h0, 32'h0};
test_input[35712:35719] = '{32'hc208c9ed, 32'h427aaca0, 32'h426ffe6f, 32'hc0eabaf9, 32'h41873101, 32'hc2297d3a, 32'h42024e35, 32'h40b7a17c};
test_output[35712:35719] = '{32'h0, 32'h427aaca0, 32'h426ffe6f, 32'h0, 32'h41873101, 32'h0, 32'h42024e35, 32'h40b7a17c};
test_input[35720:35727] = '{32'hc1f25993, 32'hc03cf820, 32'hc1ef55e4, 32'hc2adc3f3, 32'h4288a6e9, 32'h41c200ba, 32'h424879ca, 32'hc1dd8c75};
test_output[35720:35727] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4288a6e9, 32'h41c200ba, 32'h424879ca, 32'h0};
test_input[35728:35735] = '{32'hc21f3589, 32'hc2c03211, 32'hc2ab0f13, 32'h429eb5da, 32'h42c4ea99, 32'hc1f416e6, 32'hc2242cfd, 32'h4294e86f};
test_output[35728:35735] = '{32'h0, 32'h0, 32'h0, 32'h429eb5da, 32'h42c4ea99, 32'h0, 32'h0, 32'h4294e86f};
test_input[35736:35743] = '{32'h418c0756, 32'h412f9c76, 32'h41bff4b4, 32'h419c544a, 32'hc2a98b27, 32'hc27788b3, 32'hc28af7e2, 32'h42adf874};
test_output[35736:35743] = '{32'h418c0756, 32'h412f9c76, 32'h41bff4b4, 32'h419c544a, 32'h0, 32'h0, 32'h0, 32'h42adf874};
test_input[35744:35751] = '{32'hc273990a, 32'hc2ba810d, 32'h4295f419, 32'hc20af6f0, 32'h428bab0e, 32'h429d6a0e, 32'hc2bf9148, 32'h42c11f3e};
test_output[35744:35751] = '{32'h0, 32'h0, 32'h4295f419, 32'h0, 32'h428bab0e, 32'h429d6a0e, 32'h0, 32'h42c11f3e};
test_input[35752:35759] = '{32'h3fd54869, 32'h4244ced2, 32'h420e8cd8, 32'hc23d56cc, 32'hc089b061, 32'h422bedd0, 32'h415c9ffe, 32'h422427cc};
test_output[35752:35759] = '{32'h3fd54869, 32'h4244ced2, 32'h420e8cd8, 32'h0, 32'h0, 32'h422bedd0, 32'h415c9ffe, 32'h422427cc};
test_input[35760:35767] = '{32'hc248b3aa, 32'h42c6654b, 32'h42770370, 32'h42497809, 32'hc23c1234, 32'h42b816fc, 32'h421c8c71, 32'h42160377};
test_output[35760:35767] = '{32'h0, 32'h42c6654b, 32'h42770370, 32'h42497809, 32'h0, 32'h42b816fc, 32'h421c8c71, 32'h42160377};
test_input[35768:35775] = '{32'hc26dffe4, 32'h4264599b, 32'hc2a0948f, 32'h42114dd3, 32'h42b24b12, 32'h425328ef, 32'h4052fc27, 32'h42c426be};
test_output[35768:35775] = '{32'h0, 32'h4264599b, 32'h0, 32'h42114dd3, 32'h42b24b12, 32'h425328ef, 32'h4052fc27, 32'h42c426be};
test_input[35776:35783] = '{32'hc149e740, 32'hc1a64575, 32'hc29d39cc, 32'hc2b02e80, 32'hc193b673, 32'hc244cd03, 32'hc2b5aa47, 32'hc0fa56c3};
test_output[35776:35783] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35784:35791] = '{32'h42a5e7ec, 32'h429aca3c, 32'hc223a838, 32'h422d3459, 32'hc2004f53, 32'hc2b18587, 32'hc27e946f, 32'h423dda42};
test_output[35784:35791] = '{32'h42a5e7ec, 32'h429aca3c, 32'h0, 32'h422d3459, 32'h0, 32'h0, 32'h0, 32'h423dda42};
test_input[35792:35799] = '{32'h41a1efaf, 32'h4290f8cb, 32'hc216add6, 32'h40e02dc5, 32'h4201bdfb, 32'hc0b2488a, 32'hc2769167, 32'hc1392214};
test_output[35792:35799] = '{32'h41a1efaf, 32'h4290f8cb, 32'h0, 32'h40e02dc5, 32'h4201bdfb, 32'h0, 32'h0, 32'h0};
test_input[35800:35807] = '{32'hc1b06e8d, 32'h429b3ddb, 32'h4296cb7b, 32'hc22e0915, 32'hc00aab57, 32'hc2197f52, 32'hc2939389, 32'hc27bcafc};
test_output[35800:35807] = '{32'h0, 32'h429b3ddb, 32'h4296cb7b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35808:35815] = '{32'h42614667, 32'hc2bf4041, 32'h427f64e8, 32'h42afac37, 32'h428fd3e3, 32'h418e65ac, 32'h42afffc4, 32'h42ac612c};
test_output[35808:35815] = '{32'h42614667, 32'h0, 32'h427f64e8, 32'h42afac37, 32'h428fd3e3, 32'h418e65ac, 32'h42afffc4, 32'h42ac612c};
test_input[35816:35823] = '{32'h4266bd54, 32'h40d1ffa5, 32'h429233f0, 32'h4267adaa, 32'hc1bc0561, 32'hc0fc6756, 32'h4100edb6, 32'hc2c1b990};
test_output[35816:35823] = '{32'h4266bd54, 32'h40d1ffa5, 32'h429233f0, 32'h4267adaa, 32'h0, 32'h0, 32'h4100edb6, 32'h0};
test_input[35824:35831] = '{32'hc24738db, 32'h41be4d26, 32'hc28c938e, 32'h41f6ca33, 32'h42c0f191, 32'h41927000, 32'hc2817ec5, 32'hc28c1a30};
test_output[35824:35831] = '{32'h0, 32'h41be4d26, 32'h0, 32'h41f6ca33, 32'h42c0f191, 32'h41927000, 32'h0, 32'h0};
test_input[35832:35839] = '{32'h42a2ebde, 32'h422bb3ac, 32'h42beed84, 32'hc10642d6, 32'hc270e689, 32'h4214fcec, 32'hc2be19a5, 32'hc217c5a6};
test_output[35832:35839] = '{32'h42a2ebde, 32'h422bb3ac, 32'h42beed84, 32'h0, 32'h0, 32'h4214fcec, 32'h0, 32'h0};
test_input[35840:35847] = '{32'hc238ed63, 32'hc2a3869b, 32'h420803ab, 32'hc28cac3f, 32'h40391c3e, 32'h42a403e1, 32'hc1410d9f, 32'hc20b5b7e};
test_output[35840:35847] = '{32'h0, 32'h0, 32'h420803ab, 32'h0, 32'h40391c3e, 32'h42a403e1, 32'h0, 32'h0};
test_input[35848:35855] = '{32'h4095599c, 32'h42c24ff6, 32'h40bcbeaa, 32'hc0538c14, 32'h424fae42, 32'h4292f1eb, 32'h4283192f, 32'hc288440b};
test_output[35848:35855] = '{32'h4095599c, 32'h42c24ff6, 32'h40bcbeaa, 32'h0, 32'h424fae42, 32'h4292f1eb, 32'h4283192f, 32'h0};
test_input[35856:35863] = '{32'h4116c160, 32'h4217f239, 32'h42ac6ba4, 32'hc220d509, 32'hc24c5b84, 32'hc25a0551, 32'hc2a665bf, 32'hc25a3e9c};
test_output[35856:35863] = '{32'h4116c160, 32'h4217f239, 32'h42ac6ba4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35864:35871] = '{32'h414cdef1, 32'hc2a348cd, 32'h415628c2, 32'hc2a90b22, 32'h418a3a91, 32'h41ac7b41, 32'hc049ab83, 32'h428f4a26};
test_output[35864:35871] = '{32'h414cdef1, 32'h0, 32'h415628c2, 32'h0, 32'h418a3a91, 32'h41ac7b41, 32'h0, 32'h428f4a26};
test_input[35872:35879] = '{32'h421c9f9c, 32'hc20275e2, 32'h42ada7f9, 32'hc24eed87, 32'h420cc680, 32'hc28a0f5e, 32'h4220ef5a, 32'h42a35125};
test_output[35872:35879] = '{32'h421c9f9c, 32'h0, 32'h42ada7f9, 32'h0, 32'h420cc680, 32'h0, 32'h4220ef5a, 32'h42a35125};
test_input[35880:35887] = '{32'hc22b246a, 32'hc1bac006, 32'hc29566ba, 32'hc14bac86, 32'h419537ac, 32'hc29b65de, 32'hc12f481d, 32'h409bc9ef};
test_output[35880:35887] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h419537ac, 32'h0, 32'h0, 32'h409bc9ef};
test_input[35888:35895] = '{32'h4164c75e, 32'hc214376d, 32'hc20c6a6a, 32'hc21aafd1, 32'hc291576a, 32'hc2b68388, 32'h4119117d, 32'h4287ac2c};
test_output[35888:35895] = '{32'h4164c75e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4119117d, 32'h4287ac2c};
test_input[35896:35903] = '{32'h4287ed98, 32'h407b89c7, 32'hc29a7bfa, 32'h4205f687, 32'hc20cffea, 32'hc26a54a4, 32'h423a6414, 32'hc2c55098};
test_output[35896:35903] = '{32'h4287ed98, 32'h407b89c7, 32'h0, 32'h4205f687, 32'h0, 32'h0, 32'h423a6414, 32'h0};
test_input[35904:35911] = '{32'hc2836e2b, 32'h41e34138, 32'h428e15ea, 32'hc1252bd1, 32'h41fa5d26, 32'h41415209, 32'hc2279bda, 32'h41b28bd6};
test_output[35904:35911] = '{32'h0, 32'h41e34138, 32'h428e15ea, 32'h0, 32'h41fa5d26, 32'h41415209, 32'h0, 32'h41b28bd6};
test_input[35912:35919] = '{32'hc19fe707, 32'hc187c48f, 32'h418d1f10, 32'h4261e263, 32'h421d4f0e, 32'hc1fdcd41, 32'hc1cd31fb, 32'hc201e690};
test_output[35912:35919] = '{32'h0, 32'h0, 32'h418d1f10, 32'h4261e263, 32'h421d4f0e, 32'h0, 32'h0, 32'h0};
test_input[35920:35927] = '{32'h42a83dde, 32'h426e3c11, 32'hc224094c, 32'hc22871d5, 32'h42869e08, 32'hc2be8c04, 32'h429bb06e, 32'hc24d1388};
test_output[35920:35927] = '{32'h42a83dde, 32'h426e3c11, 32'h0, 32'h0, 32'h42869e08, 32'h0, 32'h429bb06e, 32'h0};
test_input[35928:35935] = '{32'h42715ca1, 32'hc2914a27, 32'hc1ee9e99, 32'h4213723f, 32'hc2c7d808, 32'h4212b636, 32'hc24e7b3a, 32'hc24a2514};
test_output[35928:35935] = '{32'h42715ca1, 32'h0, 32'h0, 32'h4213723f, 32'h0, 32'h4212b636, 32'h0, 32'h0};
test_input[35936:35943] = '{32'h425b5c52, 32'hc2a01327, 32'hc0c21c8c, 32'hc1a66e55, 32'hc20e3428, 32'h4239a9f7, 32'hc26cb701, 32'h42bd4e13};
test_output[35936:35943] = '{32'h425b5c52, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4239a9f7, 32'h0, 32'h42bd4e13};
test_input[35944:35951] = '{32'hbfdef03d, 32'h411b0cb8, 32'h42b69ed4, 32'h429919ae, 32'h42863662, 32'hc20af5a6, 32'hc24b48bf, 32'h4228ab38};
test_output[35944:35951] = '{32'h0, 32'h411b0cb8, 32'h42b69ed4, 32'h429919ae, 32'h42863662, 32'h0, 32'h0, 32'h4228ab38};
test_input[35952:35959] = '{32'h4204a2ce, 32'h4217f260, 32'hc2007541, 32'hc23896be, 32'hc22e31a4, 32'hc159992e, 32'hc1cf44c0, 32'hc28280f8};
test_output[35952:35959] = '{32'h4204a2ce, 32'h4217f260, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[35960:35967] = '{32'hc1cf7d0d, 32'hc2c77cc0, 32'h3fddcff1, 32'hc28676d5, 32'hc16156a7, 32'hc21ae185, 32'hc297ecfa, 32'h41edb139};
test_output[35960:35967] = '{32'h0, 32'h0, 32'h3fddcff1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41edb139};
test_input[35968:35975] = '{32'h42a3f47c, 32'hc1c26ffd, 32'h41c686d0, 32'hc2c74a81, 32'h42048ba3, 32'h42489e4f, 32'hc2896d0b, 32'h429dd063};
test_output[35968:35975] = '{32'h42a3f47c, 32'h0, 32'h41c686d0, 32'h0, 32'h42048ba3, 32'h42489e4f, 32'h0, 32'h429dd063};
test_input[35976:35983] = '{32'h429a7ba2, 32'h42ad5d71, 32'hc23469d9, 32'hc1d3f9ff, 32'hc237ba1c, 32'h425291e1, 32'hc1a62978, 32'hc1edb272};
test_output[35976:35983] = '{32'h429a7ba2, 32'h42ad5d71, 32'h0, 32'h0, 32'h0, 32'h425291e1, 32'h0, 32'h0};
test_input[35984:35991] = '{32'hc280f77e, 32'hc21f8937, 32'h42a7352c, 32'h3fcaab1e, 32'h41b038e0, 32'hc087c088, 32'h42286dbd, 32'h41783cdb};
test_output[35984:35991] = '{32'h0, 32'h0, 32'h42a7352c, 32'h3fcaab1e, 32'h41b038e0, 32'h0, 32'h42286dbd, 32'h41783cdb};
test_input[35992:35999] = '{32'hc2332e6f, 32'h42786af0, 32'h42625267, 32'hc287e0f7, 32'h42a65d22, 32'h4252f518, 32'hc1c377da, 32'h428f67a5};
test_output[35992:35999] = '{32'h0, 32'h42786af0, 32'h42625267, 32'h0, 32'h42a65d22, 32'h4252f518, 32'h0, 32'h428f67a5};
test_input[36000:36007] = '{32'h42696c9b, 32'hc1ba2734, 32'h426fc9b7, 32'hc22bc0cd, 32'h42975b3c, 32'h42865a04, 32'h42c6c8ba, 32'h42333758};
test_output[36000:36007] = '{32'h42696c9b, 32'h0, 32'h426fc9b7, 32'h0, 32'h42975b3c, 32'h42865a04, 32'h42c6c8ba, 32'h42333758};
test_input[36008:36015] = '{32'hc2197ace, 32'h41103896, 32'hc18b12a4, 32'h42951e80, 32'hc2971893, 32'hc253bc40, 32'hc269b895, 32'hc1721d73};
test_output[36008:36015] = '{32'h0, 32'h41103896, 32'h0, 32'h42951e80, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[36016:36023] = '{32'h41d764c6, 32'h41cfd8c7, 32'h42855681, 32'h428efc98, 32'hc0948cfc, 32'hc2552605, 32'hc2b436f0, 32'hc28b4bd0};
test_output[36016:36023] = '{32'h41d764c6, 32'h41cfd8c7, 32'h42855681, 32'h428efc98, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[36024:36031] = '{32'h41d77ca1, 32'hc2ac9fcf, 32'h422d8b4d, 32'h4162ee68, 32'h427cb3f4, 32'hc227d532, 32'hc1c2cc9a, 32'hc09b9299};
test_output[36024:36031] = '{32'h41d77ca1, 32'h0, 32'h422d8b4d, 32'h4162ee68, 32'h427cb3f4, 32'h0, 32'h0, 32'h0};
test_input[36032:36039] = '{32'h4095a238, 32'hc1407bef, 32'hc2c627f9, 32'hc2ab469b, 32'h42b91258, 32'hc2987357, 32'hc249fd88, 32'hc28f2dde};
test_output[36032:36039] = '{32'h4095a238, 32'h0, 32'h0, 32'h0, 32'h42b91258, 32'h0, 32'h0, 32'h0};
test_input[36040:36047] = '{32'hc1be0e10, 32'hc27dc51f, 32'h423afa93, 32'h4208dbf4, 32'h4254dc46, 32'h422faaa5, 32'hc2a79c05, 32'hc220f24c};
test_output[36040:36047] = '{32'h0, 32'h0, 32'h423afa93, 32'h4208dbf4, 32'h4254dc46, 32'h422faaa5, 32'h0, 32'h0};
test_input[36048:36055] = '{32'hc2279e17, 32'hc06e05ff, 32'hc2257ac4, 32'hc1e1bd00, 32'hc2be8366, 32'hc2330cd1, 32'h4287b493, 32'hc2a739eb};
test_output[36048:36055] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4287b493, 32'h0};
test_input[36056:36063] = '{32'hc0998d29, 32'hc0309518, 32'hc26df2d6, 32'h429c0e3b, 32'h4295c230, 32'hc21fda02, 32'h42c69c4d, 32'h4257cd95};
test_output[36056:36063] = '{32'h0, 32'h0, 32'h0, 32'h429c0e3b, 32'h4295c230, 32'h0, 32'h42c69c4d, 32'h4257cd95};
test_input[36064:36071] = '{32'h41ef9d16, 32'hc2aa4e8d, 32'hc1ac9f8f, 32'hc288d184, 32'h42b6bb6d, 32'h42a34686, 32'h429c302f, 32'hc1f9da02};
test_output[36064:36071] = '{32'h41ef9d16, 32'h0, 32'h0, 32'h0, 32'h42b6bb6d, 32'h42a34686, 32'h429c302f, 32'h0};
test_input[36072:36079] = '{32'h42bc7c9c, 32'hbfce0584, 32'h42c7bb11, 32'h42bb7830, 32'h405ee8bb, 32'h41e9e198, 32'h42a3c5f7, 32'h428017e7};
test_output[36072:36079] = '{32'h42bc7c9c, 32'h0, 32'h42c7bb11, 32'h42bb7830, 32'h405ee8bb, 32'h41e9e198, 32'h42a3c5f7, 32'h428017e7};
test_input[36080:36087] = '{32'hc21f7e84, 32'hc1ed4786, 32'h4242c6b3, 32'hc26ad376, 32'hc2a8d2f0, 32'h427be88e, 32'hc2aeeab6, 32'h407ca1eb};
test_output[36080:36087] = '{32'h0, 32'h0, 32'h4242c6b3, 32'h0, 32'h0, 32'h427be88e, 32'h0, 32'h407ca1eb};
test_input[36088:36095] = '{32'h428fa4d2, 32'h40b9bd25, 32'h408fbca0, 32'h42be7239, 32'h41f5a01e, 32'hc296e219, 32'hc17c1e12, 32'h4296e482};
test_output[36088:36095] = '{32'h428fa4d2, 32'h40b9bd25, 32'h408fbca0, 32'h42be7239, 32'h41f5a01e, 32'h0, 32'h0, 32'h4296e482};
test_input[36096:36103] = '{32'h428e0124, 32'hc1765cb3, 32'h41fe3728, 32'h4273c7c2, 32'hc0108d22, 32'h421905df, 32'hc207e683, 32'hc0415554};
test_output[36096:36103] = '{32'h428e0124, 32'h0, 32'h41fe3728, 32'h4273c7c2, 32'h0, 32'h421905df, 32'h0, 32'h0};
test_input[36104:36111] = '{32'hc29caf69, 32'hc2aadd14, 32'hc2b05912, 32'hc28fac35, 32'hc2ac11f0, 32'hc24086c2, 32'hc1112d3c, 32'h40b65393};
test_output[36104:36111] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40b65393};
test_input[36112:36119] = '{32'hc2acaa0b, 32'hc26df766, 32'h42bbfe0d, 32'hc223db51, 32'hc1a9cb08, 32'h41e1b495, 32'h421f260f, 32'hc10987dd};
test_output[36112:36119] = '{32'h0, 32'h0, 32'h42bbfe0d, 32'h0, 32'h0, 32'h41e1b495, 32'h421f260f, 32'h0};
test_input[36120:36127] = '{32'hc2833429, 32'h4169e402, 32'hc25990f1, 32'h4200d37d, 32'hc1548538, 32'h429d4215, 32'h42ac250d, 32'hc07cd9cb};
test_output[36120:36127] = '{32'h0, 32'h4169e402, 32'h0, 32'h4200d37d, 32'h0, 32'h429d4215, 32'h42ac250d, 32'h0};
test_input[36128:36135] = '{32'hc121ce44, 32'hc2852edf, 32'hc24d08ed, 32'hc2b71f2a, 32'h42c754e3, 32'hc1cf9728, 32'h414e205f, 32'hc293fb38};
test_output[36128:36135] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42c754e3, 32'h0, 32'h414e205f, 32'h0};
test_input[36136:36143] = '{32'h41435e4d, 32'hc234e3d7, 32'hc21279ae, 32'h4029fd4a, 32'h4106e3b6, 32'hc0b88afb, 32'hc29060d9, 32'h42a25fb0};
test_output[36136:36143] = '{32'h41435e4d, 32'h0, 32'h0, 32'h4029fd4a, 32'h4106e3b6, 32'h0, 32'h0, 32'h42a25fb0};
test_input[36144:36151] = '{32'h42845748, 32'hc23c2475, 32'hc2a215a1, 32'h42588ab8, 32'hc25c44fd, 32'hc2a112cd, 32'hc13ed82b, 32'h42264dea};
test_output[36144:36151] = '{32'h42845748, 32'h0, 32'h0, 32'h42588ab8, 32'h0, 32'h0, 32'h0, 32'h42264dea};
test_input[36152:36159] = '{32'hc26c7282, 32'hc1bcd016, 32'h42a34eda, 32'hc2577276, 32'hc1170f1a, 32'h421aefaf, 32'h4172c864, 32'h41b88ca5};
test_output[36152:36159] = '{32'h0, 32'h0, 32'h42a34eda, 32'h0, 32'h0, 32'h421aefaf, 32'h4172c864, 32'h41b88ca5};
test_input[36160:36167] = '{32'hc295bd5f, 32'hc28af730, 32'hc1b98ebb, 32'h427b5ae5, 32'hc1d0caa4, 32'h42556764, 32'hc225d640, 32'h423cfa8f};
test_output[36160:36167] = '{32'h0, 32'h0, 32'h0, 32'h427b5ae5, 32'h0, 32'h42556764, 32'h0, 32'h423cfa8f};
test_input[36168:36175] = '{32'h4295e43c, 32'h40fa344a, 32'hc0e46212, 32'hc105c7a6, 32'h414e1050, 32'h416785ce, 32'hc28a80f5, 32'h42c673b7};
test_output[36168:36175] = '{32'h4295e43c, 32'h40fa344a, 32'h0, 32'h0, 32'h414e1050, 32'h416785ce, 32'h0, 32'h42c673b7};
test_input[36176:36183] = '{32'hc293c5f3, 32'hc2b6ac67, 32'hc129c830, 32'h421114bc, 32'hc233d47d, 32'hc2c21227, 32'hc144dc97, 32'h429acb48};
test_output[36176:36183] = '{32'h0, 32'h0, 32'h0, 32'h421114bc, 32'h0, 32'h0, 32'h0, 32'h429acb48};
test_input[36184:36191] = '{32'hc2c0cf0f, 32'h40e89392, 32'h42a1fbbe, 32'h4290fd52, 32'hc28aa2f1, 32'h42975303, 32'hc28fbc45, 32'hc243bc56};
test_output[36184:36191] = '{32'h0, 32'h40e89392, 32'h42a1fbbe, 32'h4290fd52, 32'h0, 32'h42975303, 32'h0, 32'h0};
test_input[36192:36199] = '{32'hc2bd2644, 32'h4283ec9f, 32'h428c31e7, 32'h4219f991, 32'h424ed3f0, 32'h42479129, 32'hc0f902d7, 32'hc0a9003b};
test_output[36192:36199] = '{32'h0, 32'h4283ec9f, 32'h428c31e7, 32'h4219f991, 32'h424ed3f0, 32'h42479129, 32'h0, 32'h0};
test_input[36200:36207] = '{32'h426d46c8, 32'hc25c9103, 32'h42434578, 32'h4212f584, 32'hc10cfc2b, 32'hc200279a, 32'hbf4be9ed, 32'h41f9df20};
test_output[36200:36207] = '{32'h426d46c8, 32'h0, 32'h42434578, 32'h4212f584, 32'h0, 32'h0, 32'h0, 32'h41f9df20};
test_input[36208:36215] = '{32'hc2c6a25f, 32'h4298fbe0, 32'hc293031b, 32'hc2914ba7, 32'h421ce5a8, 32'h42779fdb, 32'h42332ea9, 32'h42537acf};
test_output[36208:36215] = '{32'h0, 32'h4298fbe0, 32'h0, 32'h0, 32'h421ce5a8, 32'h42779fdb, 32'h42332ea9, 32'h42537acf};
test_input[36216:36223] = '{32'h42b32437, 32'hc0ecf773, 32'h421ad3e1, 32'h42069dee, 32'hc223ddf7, 32'h415daa06, 32'hc2114b4e, 32'hc2a379ca};
test_output[36216:36223] = '{32'h42b32437, 32'h0, 32'h421ad3e1, 32'h42069dee, 32'h0, 32'h415daa06, 32'h0, 32'h0};
test_input[36224:36231] = '{32'hc298b3a6, 32'hc20bde62, 32'hc2b29a85, 32'hc2504afb, 32'hc2769857, 32'h428a5816, 32'h42240c32, 32'h429f22a2};
test_output[36224:36231] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h428a5816, 32'h42240c32, 32'h429f22a2};
test_input[36232:36239] = '{32'hc1e53347, 32'hc275d4c9, 32'hc29b4415, 32'h429d2a1b, 32'hc281e527, 32'h40b17b7f, 32'h429c8c21, 32'h429553e3};
test_output[36232:36239] = '{32'h0, 32'h0, 32'h0, 32'h429d2a1b, 32'h0, 32'h40b17b7f, 32'h429c8c21, 32'h429553e3};
test_input[36240:36247] = '{32'hc23b841c, 32'hc2a2c2eb, 32'h42463266, 32'hc29586e4, 32'hc2b83447, 32'hc2648cff, 32'h424a2df4, 32'hc04f9078};
test_output[36240:36247] = '{32'h0, 32'h0, 32'h42463266, 32'h0, 32'h0, 32'h0, 32'h424a2df4, 32'h0};
test_input[36248:36255] = '{32'hc0af854d, 32'h42c5f68b, 32'h40e014bd, 32'h42538e84, 32'h42081864, 32'hc181e449, 32'h4257c42f, 32'h42abbd0d};
test_output[36248:36255] = '{32'h0, 32'h42c5f68b, 32'h40e014bd, 32'h42538e84, 32'h42081864, 32'h0, 32'h4257c42f, 32'h42abbd0d};
test_input[36256:36263] = '{32'hc24e8245, 32'h42836d79, 32'h41ed54ac, 32'h42760df5, 32'h413eaee8, 32'hc22f3fd8, 32'h42aec597, 32'h42ad1dae};
test_output[36256:36263] = '{32'h0, 32'h42836d79, 32'h41ed54ac, 32'h42760df5, 32'h413eaee8, 32'h0, 32'h42aec597, 32'h42ad1dae};
test_input[36264:36271] = '{32'h426b815f, 32'hc2b3fef4, 32'hc2823ed0, 32'hc2b64531, 32'h42194caa, 32'h42afca2d, 32'hc2880a34, 32'h424cac87};
test_output[36264:36271] = '{32'h426b815f, 32'h0, 32'h0, 32'h0, 32'h42194caa, 32'h42afca2d, 32'h0, 32'h424cac87};
test_input[36272:36279] = '{32'h428464c7, 32'hc298f45b, 32'hc29a460b, 32'h42b0d1cd, 32'h420505c1, 32'h429e1316, 32'hc2a04fe4, 32'h422cbad4};
test_output[36272:36279] = '{32'h428464c7, 32'h0, 32'h0, 32'h42b0d1cd, 32'h420505c1, 32'h429e1316, 32'h0, 32'h422cbad4};
test_input[36280:36287] = '{32'h42b1f53b, 32'hc1e9b585, 32'hc2b827d4, 32'hc262d27b, 32'hc23f5c07, 32'h41185c12, 32'h42a6ba3a, 32'h42322a54};
test_output[36280:36287] = '{32'h42b1f53b, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41185c12, 32'h42a6ba3a, 32'h42322a54};
test_input[36288:36295] = '{32'hc1a83e9f, 32'h420b8186, 32'h42bdbe09, 32'h428105fd, 32'h423176e0, 32'h429d46f1, 32'hc284dbe2, 32'h4275b2b5};
test_output[36288:36295] = '{32'h0, 32'h420b8186, 32'h42bdbe09, 32'h428105fd, 32'h423176e0, 32'h429d46f1, 32'h0, 32'h4275b2b5};
test_input[36296:36303] = '{32'h42b6be73, 32'hc28d8233, 32'h4060c9a8, 32'h4202377a, 32'h41c5d4dc, 32'hc220e755, 32'h420f2d42, 32'h42b99204};
test_output[36296:36303] = '{32'h42b6be73, 32'h0, 32'h4060c9a8, 32'h4202377a, 32'h41c5d4dc, 32'h0, 32'h420f2d42, 32'h42b99204};
test_input[36304:36311] = '{32'hc2b1330d, 32'h428a8914, 32'h41d12e98, 32'h40680b16, 32'hc1a6200f, 32'h408af258, 32'hc20d1080, 32'h421e6541};
test_output[36304:36311] = '{32'h0, 32'h428a8914, 32'h41d12e98, 32'h40680b16, 32'h0, 32'h408af258, 32'h0, 32'h421e6541};
test_input[36312:36319] = '{32'h4240be3d, 32'h422e49aa, 32'hc05a47ac, 32'hc269ec2f, 32'hc2a07a1a, 32'h42700853, 32'hc2937da8, 32'hc1679c2e};
test_output[36312:36319] = '{32'h4240be3d, 32'h422e49aa, 32'h0, 32'h0, 32'h0, 32'h42700853, 32'h0, 32'h0};
test_input[36320:36327] = '{32'hc20b1398, 32'h4090bd54, 32'hc2c1965f, 32'h42ac9694, 32'h427aa16f, 32'hc09fe458, 32'hc1e33ff1, 32'hc2721f44};
test_output[36320:36327] = '{32'h0, 32'h4090bd54, 32'h0, 32'h42ac9694, 32'h427aa16f, 32'h0, 32'h0, 32'h0};
test_input[36328:36335] = '{32'h419cb50f, 32'h4281f22e, 32'h421b3485, 32'h4048ed4a, 32'h42189e10, 32'hc1bbfb3b, 32'hc20fbc19, 32'h3fd79e05};
test_output[36328:36335] = '{32'h419cb50f, 32'h4281f22e, 32'h421b3485, 32'h4048ed4a, 32'h42189e10, 32'h0, 32'h0, 32'h3fd79e05};
test_input[36336:36343] = '{32'h4271ba1d, 32'hc14461e4, 32'h421a3cb5, 32'hc02115de, 32'h42c23a18, 32'h4285581f, 32'hc281b3d7, 32'hc256c116};
test_output[36336:36343] = '{32'h4271ba1d, 32'h0, 32'h421a3cb5, 32'h0, 32'h42c23a18, 32'h4285581f, 32'h0, 32'h0};
test_input[36344:36351] = '{32'h412b628b, 32'hc12824a8, 32'h427fda64, 32'h41921147, 32'hc28bb881, 32'hc2a7c6a5, 32'h41b2a32a, 32'hc2a6856c};
test_output[36344:36351] = '{32'h412b628b, 32'h0, 32'h427fda64, 32'h41921147, 32'h0, 32'h0, 32'h41b2a32a, 32'h0};
test_input[36352:36359] = '{32'h41838e79, 32'hc2b172bb, 32'h417fb483, 32'h42bed9bb, 32'h427d0f38, 32'h428527a2, 32'h42257a4e, 32'h42b289f9};
test_output[36352:36359] = '{32'h41838e79, 32'h0, 32'h417fb483, 32'h42bed9bb, 32'h427d0f38, 32'h428527a2, 32'h42257a4e, 32'h42b289f9};
test_input[36360:36367] = '{32'h414ac241, 32'h42a23972, 32'hc191680b, 32'hc1c2d005, 32'h42012dad, 32'hc230f999, 32'h4284c384, 32'hc289024d};
test_output[36360:36367] = '{32'h414ac241, 32'h42a23972, 32'h0, 32'h0, 32'h42012dad, 32'h0, 32'h4284c384, 32'h0};
test_input[36368:36375] = '{32'hbe696b2d, 32'hc26a648b, 32'h424d2871, 32'hc2a7fdd7, 32'hc103ecb1, 32'h426b8f3a, 32'hc152e484, 32'h41e4d363};
test_output[36368:36375] = '{32'h0, 32'h0, 32'h424d2871, 32'h0, 32'h0, 32'h426b8f3a, 32'h0, 32'h41e4d363};
test_input[36376:36383] = '{32'h42812c4a, 32'h4269d9b6, 32'h42376201, 32'h42964736, 32'h42bf1bfe, 32'hc25b19c9, 32'hc1c58324, 32'hc2010db0};
test_output[36376:36383] = '{32'h42812c4a, 32'h4269d9b6, 32'h42376201, 32'h42964736, 32'h42bf1bfe, 32'h0, 32'h0, 32'h0};
test_input[36384:36391] = '{32'h42249a47, 32'hc2ab6783, 32'h410b78ba, 32'hc12fdb8b, 32'hc24d009c, 32'h42c7cead, 32'hc2363722, 32'h42b59ca2};
test_output[36384:36391] = '{32'h42249a47, 32'h0, 32'h410b78ba, 32'h0, 32'h0, 32'h42c7cead, 32'h0, 32'h42b59ca2};
test_input[36392:36399] = '{32'h428ff0fe, 32'hc2a17f97, 32'hc24170dd, 32'hc269ddb2, 32'h42484139, 32'hc2c0d7cd, 32'hc2b9504e, 32'hc28a98cd};
test_output[36392:36399] = '{32'h428ff0fe, 32'h0, 32'h0, 32'h0, 32'h42484139, 32'h0, 32'h0, 32'h0};
test_input[36400:36407] = '{32'h4279aeb6, 32'hc27cf354, 32'hc17b0509, 32'hc1e7b406, 32'hc018bb8c, 32'hc21a653e, 32'hc2ad64a9, 32'h4194a83e};
test_output[36400:36407] = '{32'h4279aeb6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4194a83e};
test_input[36408:36415] = '{32'h41d42c6b, 32'h425c6ff1, 32'h4049083b, 32'hc0db01f3, 32'h41a80abd, 32'hc227d260, 32'hc1e769b4, 32'hc295eef9};
test_output[36408:36415] = '{32'h41d42c6b, 32'h425c6ff1, 32'h4049083b, 32'h0, 32'h41a80abd, 32'h0, 32'h0, 32'h0};
test_input[36416:36423] = '{32'hc2322cf7, 32'h42a05c5c, 32'hc230fd85, 32'h41932c8b, 32'h42521c15, 32'hc28f2e08, 32'h424291c3, 32'h42109dee};
test_output[36416:36423] = '{32'h0, 32'h42a05c5c, 32'h0, 32'h41932c8b, 32'h42521c15, 32'h0, 32'h424291c3, 32'h42109dee};
test_input[36424:36431] = '{32'hc2a96380, 32'hc243b90c, 32'hc09019bf, 32'hc2805776, 32'hc1ae4984, 32'hc26bb094, 32'hc0f6d30a, 32'hc1c92d22};
test_output[36424:36431] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[36432:36439] = '{32'hc1fa2e21, 32'h427d8963, 32'hc15c8786, 32'hc2aa04c7, 32'h4139e4cc, 32'hbff9f163, 32'hc211b513, 32'h42c321ee};
test_output[36432:36439] = '{32'h0, 32'h427d8963, 32'h0, 32'h0, 32'h4139e4cc, 32'h0, 32'h0, 32'h42c321ee};
test_input[36440:36447] = '{32'hc2a98590, 32'h42754bb7, 32'h41e682c3, 32'hc2a64dc3, 32'h4211d2d4, 32'h422fc015, 32'h42c511c5, 32'h42ae5bae};
test_output[36440:36447] = '{32'h0, 32'h42754bb7, 32'h41e682c3, 32'h0, 32'h4211d2d4, 32'h422fc015, 32'h42c511c5, 32'h42ae5bae};
test_input[36448:36455] = '{32'h420fdf7d, 32'hc23c0cdc, 32'hc1934690, 32'hc2a43ab1, 32'h419a1ed7, 32'hc1ddd8f6, 32'h414354c1, 32'h41fcd228};
test_output[36448:36455] = '{32'h420fdf7d, 32'h0, 32'h0, 32'h0, 32'h419a1ed7, 32'h0, 32'h414354c1, 32'h41fcd228};
test_input[36456:36463] = '{32'h42adfc0b, 32'h42a62826, 32'hc2abfa18, 32'hc1e498c1, 32'hc272e1d8, 32'hc0f75c90, 32'h40133172, 32'h42c1a9b3};
test_output[36456:36463] = '{32'h42adfc0b, 32'h42a62826, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40133172, 32'h42c1a9b3};
test_input[36464:36471] = '{32'hc287b3a5, 32'hc1b8fdcd, 32'h424abaa0, 32'h427e4020, 32'hc14b3a0e, 32'hc23463c2, 32'h42904804, 32'hc255cb94};
test_output[36464:36471] = '{32'h0, 32'h0, 32'h424abaa0, 32'h427e4020, 32'h0, 32'h0, 32'h42904804, 32'h0};
test_input[36472:36479] = '{32'hc1679943, 32'hc1292022, 32'hc2b3a44a, 32'hc11efca4, 32'h418fe945, 32'h421eb6b6, 32'hc213143a, 32'h40009793};
test_output[36472:36479] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h418fe945, 32'h421eb6b6, 32'h0, 32'h40009793};
test_input[36480:36487] = '{32'hc21a8c32, 32'hc2922c7f, 32'hc2c22b7d, 32'hc270f340, 32'hc26ab7ff, 32'h421a9271, 32'hc26c0ac9, 32'hc2c2ff38};
test_output[36480:36487] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h421a9271, 32'h0, 32'h0};
test_input[36488:36495] = '{32'hc29bbe4b, 32'h4102c508, 32'h42a8fe1b, 32'hc1b9c2ad, 32'hc2757614, 32'h42160dbd, 32'hc25c0166, 32'h425fb257};
test_output[36488:36495] = '{32'h0, 32'h4102c508, 32'h42a8fe1b, 32'h0, 32'h0, 32'h42160dbd, 32'h0, 32'h425fb257};
test_input[36496:36503] = '{32'h429fcdec, 32'h42888aaf, 32'h42262af0, 32'hc287a4e0, 32'h426fd8ce, 32'h42202bf2, 32'h426a0a91, 32'hc26faf22};
test_output[36496:36503] = '{32'h429fcdec, 32'h42888aaf, 32'h42262af0, 32'h0, 32'h426fd8ce, 32'h42202bf2, 32'h426a0a91, 32'h0};
test_input[36504:36511] = '{32'hc2b985e1, 32'h40b0026b, 32'hc2b5054b, 32'hc2ad3275, 32'h428ebe45, 32'hc251298d, 32'h429f4210, 32'h4239828c};
test_output[36504:36511] = '{32'h0, 32'h40b0026b, 32'h0, 32'h0, 32'h428ebe45, 32'h0, 32'h429f4210, 32'h4239828c};
test_input[36512:36519] = '{32'h428a0eb0, 32'h42b4edcd, 32'h421b616e, 32'hc284ac32, 32'hc25279e8, 32'hc2109bbb, 32'h4040d747, 32'hc27a5f28};
test_output[36512:36519] = '{32'h428a0eb0, 32'h42b4edcd, 32'h421b616e, 32'h0, 32'h0, 32'h0, 32'h4040d747, 32'h0};
test_input[36520:36527] = '{32'hc24337ad, 32'h42b255ff, 32'hc2aeda34, 32'hc290f897, 32'h41c1eb65, 32'h42be6921, 32'h4299b198, 32'h42c66c51};
test_output[36520:36527] = '{32'h0, 32'h42b255ff, 32'h0, 32'h0, 32'h41c1eb65, 32'h42be6921, 32'h4299b198, 32'h42c66c51};
test_input[36528:36535] = '{32'hc20258ab, 32'h40e6fc29, 32'hc2856285, 32'hc29d35a9, 32'hc223181a, 32'h42c3972b, 32'h4220a2f1, 32'h425e176b};
test_output[36528:36535] = '{32'h0, 32'h40e6fc29, 32'h0, 32'h0, 32'h0, 32'h42c3972b, 32'h4220a2f1, 32'h425e176b};
test_input[36536:36543] = '{32'h41a38acc, 32'h41db3578, 32'h42255200, 32'h42af9a86, 32'h426d1335, 32'h4127625d, 32'hc08dc76c, 32'hc1d97768};
test_output[36536:36543] = '{32'h41a38acc, 32'h41db3578, 32'h42255200, 32'h42af9a86, 32'h426d1335, 32'h4127625d, 32'h0, 32'h0};
test_input[36544:36551] = '{32'h4287ef6c, 32'hc1cd16aa, 32'hc1cc2a4c, 32'h408c0024, 32'h40d63cdd, 32'hc2b1cd5d, 32'h421a1c69, 32'hc22384a2};
test_output[36544:36551] = '{32'h4287ef6c, 32'h0, 32'h0, 32'h408c0024, 32'h40d63cdd, 32'h0, 32'h421a1c69, 32'h0};
test_input[36552:36559] = '{32'h42769298, 32'h429eef0f, 32'hc225df8b, 32'hc2b5b089, 32'hc25150ff, 32'hc2b4960c, 32'hc287803f, 32'h42c44c4e};
test_output[36552:36559] = '{32'h42769298, 32'h429eef0f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42c44c4e};
test_input[36560:36567] = '{32'hc2097112, 32'hc2b78f6e, 32'h428ff219, 32'h42a2d06b, 32'hc2c36350, 32'hc260b857, 32'hc229b79b, 32'h42c596b5};
test_output[36560:36567] = '{32'h0, 32'h0, 32'h428ff219, 32'h42a2d06b, 32'h0, 32'h0, 32'h0, 32'h42c596b5};
test_input[36568:36575] = '{32'h4233703d, 32'h42a6cc06, 32'h428d4f1c, 32'h42966896, 32'h418b3dc8, 32'h42adc1cf, 32'hc0d692a4, 32'h424f8d35};
test_output[36568:36575] = '{32'h4233703d, 32'h42a6cc06, 32'h428d4f1c, 32'h42966896, 32'h418b3dc8, 32'h42adc1cf, 32'h0, 32'h424f8d35};
test_input[36576:36583] = '{32'hc2c5a14e, 32'hc1e9c8f2, 32'h4291e152, 32'hc29ee124, 32'h42a30e7b, 32'h42bde05a, 32'h426cae7b, 32'hc1ad052f};
test_output[36576:36583] = '{32'h0, 32'h0, 32'h4291e152, 32'h0, 32'h42a30e7b, 32'h42bde05a, 32'h426cae7b, 32'h0};
test_input[36584:36591] = '{32'hc296e447, 32'h42348ef8, 32'hc2b9dce6, 32'h4216da2e, 32'hc1fc8ed1, 32'h4290536f, 32'h4056ee89, 32'hc120fd82};
test_output[36584:36591] = '{32'h0, 32'h42348ef8, 32'h0, 32'h4216da2e, 32'h0, 32'h4290536f, 32'h4056ee89, 32'h0};
test_input[36592:36599] = '{32'hc2be9d30, 32'hc232b078, 32'h420373dc, 32'h4128f50f, 32'h4085d1b7, 32'hc2b5f0af, 32'h425575dd, 32'hc2bfeaf7};
test_output[36592:36599] = '{32'h0, 32'h0, 32'h420373dc, 32'h4128f50f, 32'h4085d1b7, 32'h0, 32'h425575dd, 32'h0};
test_input[36600:36607] = '{32'h428b6ca5, 32'h42a6dd85, 32'hc294b12f, 32'h41fd9e06, 32'hc263b896, 32'h42a6b7ef, 32'hc08d19f9, 32'h4177188d};
test_output[36600:36607] = '{32'h428b6ca5, 32'h42a6dd85, 32'h0, 32'h41fd9e06, 32'h0, 32'h42a6b7ef, 32'h0, 32'h4177188d};
test_input[36608:36615] = '{32'h42717e0b, 32'h4290969d, 32'h4231e05e, 32'hc10c3da7, 32'hc29f908a, 32'hc2b7fc31, 32'h4298c8d2, 32'hc25136ae};
test_output[36608:36615] = '{32'h42717e0b, 32'h4290969d, 32'h4231e05e, 32'h0, 32'h0, 32'h0, 32'h4298c8d2, 32'h0};
test_input[36616:36623] = '{32'hc26c113f, 32'hc2c2c453, 32'h4297d9d2, 32'h41f42974, 32'h42a6b186, 32'h41a58f3d, 32'h422308e1, 32'h41b70205};
test_output[36616:36623] = '{32'h0, 32'h0, 32'h4297d9d2, 32'h41f42974, 32'h42a6b186, 32'h41a58f3d, 32'h422308e1, 32'h41b70205};
test_input[36624:36631] = '{32'h41a985ef, 32'hc2c678c9, 32'h41f8aea9, 32'h424b4964, 32'h42897357, 32'h42ae2dd9, 32'h3fd678a3, 32'h42b58228};
test_output[36624:36631] = '{32'h41a985ef, 32'h0, 32'h41f8aea9, 32'h424b4964, 32'h42897357, 32'h42ae2dd9, 32'h3fd678a3, 32'h42b58228};
test_input[36632:36639] = '{32'h419b566c, 32'hc2239e54, 32'hc2bd6796, 32'h428d07bd, 32'h4283058a, 32'h425bc4e9, 32'h42262709, 32'h424780e6};
test_output[36632:36639] = '{32'h419b566c, 32'h0, 32'h0, 32'h428d07bd, 32'h4283058a, 32'h425bc4e9, 32'h42262709, 32'h424780e6};
test_input[36640:36647] = '{32'h42b98d83, 32'h41c34fff, 32'h4237669f, 32'hc184501d, 32'h415d19f5, 32'hc28071ff, 32'h42891837, 32'h42a1caa2};
test_output[36640:36647] = '{32'h42b98d83, 32'h41c34fff, 32'h4237669f, 32'h0, 32'h415d19f5, 32'h0, 32'h42891837, 32'h42a1caa2};
test_input[36648:36655] = '{32'h40cecbce, 32'h4285cfbe, 32'hc2bc50cc, 32'hc2a7a7d3, 32'h42993b60, 32'h4289bef0, 32'h42bb8fd2, 32'h420280ba};
test_output[36648:36655] = '{32'h40cecbce, 32'h4285cfbe, 32'h0, 32'h0, 32'h42993b60, 32'h4289bef0, 32'h42bb8fd2, 32'h420280ba};
test_input[36656:36663] = '{32'h419806f8, 32'h41a199e2, 32'hc29852de, 32'h41ecee11, 32'hc2c7ee12, 32'h420f0333, 32'hc218ec0e, 32'hc19a42ac};
test_output[36656:36663] = '{32'h419806f8, 32'h41a199e2, 32'h0, 32'h41ecee11, 32'h0, 32'h420f0333, 32'h0, 32'h0};
test_input[36664:36671] = '{32'h423089f6, 32'hc2841e55, 32'hc2344f48, 32'hc26bed0a, 32'h42c49203, 32'hc1fb7142, 32'h424cf3c7, 32'hc20f8c27};
test_output[36664:36671] = '{32'h423089f6, 32'h0, 32'h0, 32'h0, 32'h42c49203, 32'h0, 32'h424cf3c7, 32'h0};
test_input[36672:36679] = '{32'hc100bb2f, 32'h42b10c97, 32'h42267cfa, 32'h411699b4, 32'h41b9621a, 32'hc1e982b0, 32'hc24599b7, 32'h421f128f};
test_output[36672:36679] = '{32'h0, 32'h42b10c97, 32'h42267cfa, 32'h411699b4, 32'h41b9621a, 32'h0, 32'h0, 32'h421f128f};
test_input[36680:36687] = '{32'h42838268, 32'hc19ceb1d, 32'hc197bf6c, 32'h42942a10, 32'hc1629cf1, 32'hc21c2525, 32'hc15a3c57, 32'hc2a740df};
test_output[36680:36687] = '{32'h42838268, 32'h0, 32'h0, 32'h42942a10, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[36688:36695] = '{32'hc2428dca, 32'h408df77f, 32'hc299db31, 32'hc1d02399, 32'h427369c6, 32'h42000925, 32'hc1f68856, 32'hc091e586};
test_output[36688:36695] = '{32'h0, 32'h408df77f, 32'h0, 32'h0, 32'h427369c6, 32'h42000925, 32'h0, 32'h0};
test_input[36696:36703] = '{32'h41c1eea9, 32'hc286b9ce, 32'h4272ad87, 32'h409db695, 32'hc22a71cf, 32'h40b5f486, 32'hc29f97c3, 32'h42b13098};
test_output[36696:36703] = '{32'h41c1eea9, 32'h0, 32'h4272ad87, 32'h409db695, 32'h0, 32'h40b5f486, 32'h0, 32'h42b13098};
test_input[36704:36711] = '{32'hc251d6dd, 32'hc2220a7d, 32'hc285a92f, 32'h42997064, 32'h424a264e, 32'h427be672, 32'h429c13da, 32'hc28693a0};
test_output[36704:36711] = '{32'h0, 32'h0, 32'h0, 32'h42997064, 32'h424a264e, 32'h427be672, 32'h429c13da, 32'h0};
test_input[36712:36719] = '{32'hc28e476b, 32'hc26fe69c, 32'h42777f2b, 32'h42a2e531, 32'hc19a9071, 32'h4213edcf, 32'h428ed531, 32'hc2968af8};
test_output[36712:36719] = '{32'h0, 32'h0, 32'h42777f2b, 32'h42a2e531, 32'h0, 32'h4213edcf, 32'h428ed531, 32'h0};
test_input[36720:36727] = '{32'h42816f4f, 32'h426df045, 32'h42ae7982, 32'hc1af2d22, 32'hc246de36, 32'h41460e7b, 32'h425af64e, 32'h4281734e};
test_output[36720:36727] = '{32'h42816f4f, 32'h426df045, 32'h42ae7982, 32'h0, 32'h0, 32'h41460e7b, 32'h425af64e, 32'h4281734e};
test_input[36728:36735] = '{32'h425eb8ee, 32'hc26fde03, 32'h421c7aa0, 32'h419e99e4, 32'hc2471a5e, 32'h41e36661, 32'h419dc8a7, 32'hc27ff8ad};
test_output[36728:36735] = '{32'h425eb8ee, 32'h0, 32'h421c7aa0, 32'h419e99e4, 32'h0, 32'h41e36661, 32'h419dc8a7, 32'h0};
test_input[36736:36743] = '{32'hc1b7cb23, 32'h42bffe9c, 32'h4245e063, 32'h413a3ef2, 32'h42852556, 32'h428a7305, 32'h42af53ab, 32'hc2b510d6};
test_output[36736:36743] = '{32'h0, 32'h42bffe9c, 32'h4245e063, 32'h413a3ef2, 32'h42852556, 32'h428a7305, 32'h42af53ab, 32'h0};
test_input[36744:36751] = '{32'hc2bda610, 32'hc2070dfb, 32'hc2569277, 32'h41ee2a79, 32'hc2a63c03, 32'hc291dc66, 32'hc2989db5, 32'hc227a504};
test_output[36744:36751] = '{32'h0, 32'h0, 32'h0, 32'h41ee2a79, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[36752:36759] = '{32'hc2bd4f31, 32'h400a33cc, 32'hc2286d16, 32'h42b0af1f, 32'hbf01eb52, 32'hc29c6537, 32'hc2a34569, 32'hc1210b2a};
test_output[36752:36759] = '{32'h0, 32'h400a33cc, 32'h0, 32'h42b0af1f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[36760:36767] = '{32'h427627f7, 32'hc190be8d, 32'hc214ff77, 32'h422c1203, 32'h42895916, 32'h42b69b68, 32'h42823a7e, 32'hc28bc1c3};
test_output[36760:36767] = '{32'h427627f7, 32'h0, 32'h0, 32'h422c1203, 32'h42895916, 32'h42b69b68, 32'h42823a7e, 32'h0};
test_input[36768:36775] = '{32'h426bfb26, 32'hc1048f09, 32'hc2af1870, 32'h428b3b85, 32'hc180c96b, 32'h428c50ab, 32'hc018df84, 32'hc2810dec};
test_output[36768:36775] = '{32'h426bfb26, 32'h0, 32'h0, 32'h428b3b85, 32'h0, 32'h428c50ab, 32'h0, 32'h0};
test_input[36776:36783] = '{32'h41fbdb5e, 32'hc2932eef, 32'hc2af7089, 32'hc1ac49d7, 32'hc178fee1, 32'hc25018fc, 32'h4090652b, 32'h4246046b};
test_output[36776:36783] = '{32'h41fbdb5e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4090652b, 32'h4246046b};
test_input[36784:36791] = '{32'h42314d2a, 32'h42c15824, 32'hc26c043e, 32'hbf7f4683, 32'h41ae6f10, 32'hc22bcace, 32'hc24243a6, 32'hc1f9f598};
test_output[36784:36791] = '{32'h42314d2a, 32'h42c15824, 32'h0, 32'h0, 32'h41ae6f10, 32'h0, 32'h0, 32'h0};
test_input[36792:36799] = '{32'hc29b1fba, 32'hc2906196, 32'hc2c583f8, 32'hc1af2d98, 32'h42c19804, 32'hc1472855, 32'h424fc421, 32'hc263606c};
test_output[36792:36799] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42c19804, 32'h0, 32'h424fc421, 32'h0};
test_input[36800:36807] = '{32'h41ff3f8c, 32'hc2042a87, 32'hc27d0447, 32'hc10f555b, 32'hc22824c1, 32'hc2093f5e, 32'h40c38a15, 32'hc21fe79b};
test_output[36800:36807] = '{32'h41ff3f8c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40c38a15, 32'h0};
test_input[36808:36815] = '{32'h4282a1cb, 32'hc2ab558f, 32'hc230b873, 32'h416aad30, 32'h4289322e, 32'h429e77fd, 32'h429d3ed8, 32'h41cec457};
test_output[36808:36815] = '{32'h4282a1cb, 32'h0, 32'h0, 32'h416aad30, 32'h4289322e, 32'h429e77fd, 32'h429d3ed8, 32'h41cec457};
test_input[36816:36823] = '{32'hc225ad58, 32'h42802c23, 32'h4149c0e5, 32'h420714ed, 32'hc233491e, 32'hc17b8197, 32'h42ac31ea, 32'hc09499db};
test_output[36816:36823] = '{32'h0, 32'h42802c23, 32'h4149c0e5, 32'h420714ed, 32'h0, 32'h0, 32'h42ac31ea, 32'h0};
test_input[36824:36831] = '{32'hc26fb780, 32'hc0b1dbd0, 32'h42abf555, 32'hc20d8980, 32'h42be1f8d, 32'hc2ac3297, 32'hc241088c, 32'h4224137c};
test_output[36824:36831] = '{32'h0, 32'h0, 32'h42abf555, 32'h0, 32'h42be1f8d, 32'h0, 32'h0, 32'h4224137c};
test_input[36832:36839] = '{32'h41105daf, 32'h42aa1e25, 32'h41f6b069, 32'h4284a71e, 32'hc29aabb5, 32'hc25a77b0, 32'h4175e91a, 32'h42352f59};
test_output[36832:36839] = '{32'h41105daf, 32'h42aa1e25, 32'h41f6b069, 32'h4284a71e, 32'h0, 32'h0, 32'h4175e91a, 32'h42352f59};
test_input[36840:36847] = '{32'hc29d8a3b, 32'h411b5b94, 32'hbfff0e2b, 32'hc26b56db, 32'h421f325c, 32'hc2916afa, 32'h428e01f7, 32'h41ef8871};
test_output[36840:36847] = '{32'h0, 32'h411b5b94, 32'h0, 32'h0, 32'h421f325c, 32'h0, 32'h428e01f7, 32'h41ef8871};
test_input[36848:36855] = '{32'hc28cc12c, 32'h416761ea, 32'h422ac9a3, 32'h429f4cfc, 32'h42592c67, 32'hc28f070d, 32'hc1ce1047, 32'hc28d9a74};
test_output[36848:36855] = '{32'h0, 32'h416761ea, 32'h422ac9a3, 32'h429f4cfc, 32'h42592c67, 32'h0, 32'h0, 32'h0};
test_input[36856:36863] = '{32'h4291b95f, 32'hc069e664, 32'h429fe4bb, 32'hc2149fcc, 32'hc29cf48e, 32'h42adacee, 32'h429bc49d, 32'h42a89759};
test_output[36856:36863] = '{32'h4291b95f, 32'h0, 32'h429fe4bb, 32'h0, 32'h0, 32'h42adacee, 32'h429bc49d, 32'h42a89759};
test_input[36864:36871] = '{32'hc1d4249b, 32'hc2b2763e, 32'hc227d878, 32'h4266d5f6, 32'hc29d013a, 32'hc133a14e, 32'h42b87ddf, 32'h41569cd6};
test_output[36864:36871] = '{32'h0, 32'h0, 32'h0, 32'h4266d5f6, 32'h0, 32'h0, 32'h42b87ddf, 32'h41569cd6};
test_input[36872:36879] = '{32'hc1f7bdb8, 32'hc2a3de57, 32'h41aaceaa, 32'h424f6fc7, 32'hc27f5454, 32'h422b5c03, 32'h4274238c, 32'h4295b8db};
test_output[36872:36879] = '{32'h0, 32'h0, 32'h41aaceaa, 32'h424f6fc7, 32'h0, 32'h422b5c03, 32'h4274238c, 32'h4295b8db};
test_input[36880:36887] = '{32'h42965228, 32'h427d8da5, 32'h4216aa25, 32'hc24d17eb, 32'h40c256bd, 32'hc185dd5e, 32'h40f42723, 32'h427cd25b};
test_output[36880:36887] = '{32'h42965228, 32'h427d8da5, 32'h4216aa25, 32'h0, 32'h40c256bd, 32'h0, 32'h40f42723, 32'h427cd25b};
test_input[36888:36895] = '{32'hc2922697, 32'hc19127e6, 32'h423a2064, 32'hc1d6ca43, 32'hc2c3beac, 32'h41f04d24, 32'h4219b2b0, 32'hc2bbb7a0};
test_output[36888:36895] = '{32'h0, 32'h0, 32'h423a2064, 32'h0, 32'h0, 32'h41f04d24, 32'h4219b2b0, 32'h0};
test_input[36896:36903] = '{32'h4228c3a1, 32'h42a80625, 32'hc1d62bae, 32'h4241a55c, 32'h42be0b46, 32'h42950074, 32'h42ae5440, 32'h42c125e8};
test_output[36896:36903] = '{32'h4228c3a1, 32'h42a80625, 32'h0, 32'h4241a55c, 32'h42be0b46, 32'h42950074, 32'h42ae5440, 32'h42c125e8};
test_input[36904:36911] = '{32'hc294e8c2, 32'hc2288cac, 32'h41ba3bb8, 32'hc1ff47b9, 32'hc1edc8d5, 32'hc221bc90, 32'h428233f2, 32'hc0008c06};
test_output[36904:36911] = '{32'h0, 32'h0, 32'h41ba3bb8, 32'h0, 32'h0, 32'h0, 32'h428233f2, 32'h0};
test_input[36912:36919] = '{32'h42914f1d, 32'h4230d560, 32'h40b1e9b8, 32'h4283109b, 32'hc2c3e77b, 32'h426bda57, 32'h420b4964, 32'hc20724e7};
test_output[36912:36919] = '{32'h42914f1d, 32'h4230d560, 32'h40b1e9b8, 32'h4283109b, 32'h0, 32'h426bda57, 32'h420b4964, 32'h0};
test_input[36920:36927] = '{32'h428d9c3f, 32'hc2259b7e, 32'h4246c5a2, 32'h40e8a2fd, 32'hc2a615a7, 32'h42bf5b52, 32'hc2abbbd7, 32'h42095666};
test_output[36920:36927] = '{32'h428d9c3f, 32'h0, 32'h4246c5a2, 32'h40e8a2fd, 32'h0, 32'h42bf5b52, 32'h0, 32'h42095666};
test_input[36928:36935] = '{32'h4130550b, 32'h4255a424, 32'hc266d2d1, 32'h42bedd3a, 32'h424fbd7c, 32'hc24a8005, 32'h41361821, 32'h42c0be8e};
test_output[36928:36935] = '{32'h4130550b, 32'h4255a424, 32'h0, 32'h42bedd3a, 32'h424fbd7c, 32'h0, 32'h41361821, 32'h42c0be8e};
test_input[36936:36943] = '{32'h42c417c4, 32'h4242471b, 32'h420987f8, 32'hc285b92d, 32'hc29e59dd, 32'h4257163f, 32'hc2bd694e, 32'h41537fc2};
test_output[36936:36943] = '{32'h42c417c4, 32'h4242471b, 32'h420987f8, 32'h0, 32'h0, 32'h4257163f, 32'h0, 32'h41537fc2};
test_input[36944:36951] = '{32'hc28c95eb, 32'hc23e4f24, 32'hc1ade85f, 32'h40b3c285, 32'h423335a6, 32'hc24b8069, 32'hc24d8dc8, 32'hc2c2f687};
test_output[36944:36951] = '{32'h0, 32'h0, 32'h0, 32'h40b3c285, 32'h423335a6, 32'h0, 32'h0, 32'h0};
test_input[36952:36959] = '{32'h42c089bb, 32'hc260cce8, 32'h42977fc2, 32'h428ddb1c, 32'h4246ca4d, 32'hc1941f40, 32'hc2008dc9, 32'hc24b5170};
test_output[36952:36959] = '{32'h42c089bb, 32'h0, 32'h42977fc2, 32'h428ddb1c, 32'h4246ca4d, 32'h0, 32'h0, 32'h0};
test_input[36960:36967] = '{32'h42a01169, 32'h42855981, 32'hc29097ef, 32'h42916d41, 32'h426c7632, 32'h42c450ea, 32'hc180f1be, 32'h40ddf05e};
test_output[36960:36967] = '{32'h42a01169, 32'h42855981, 32'h0, 32'h42916d41, 32'h426c7632, 32'h42c450ea, 32'h0, 32'h40ddf05e};
test_input[36968:36975] = '{32'hc2b946e2, 32'h41ebc1d2, 32'hc2c4648a, 32'h4244d24d, 32'h42901783, 32'hc0c0185b, 32'hc240968b, 32'hc2ae1773};
test_output[36968:36975] = '{32'h0, 32'h41ebc1d2, 32'h0, 32'h4244d24d, 32'h42901783, 32'h0, 32'h0, 32'h0};
test_input[36976:36983] = '{32'hc174103c, 32'hc1e1c8e2, 32'hc24483da, 32'hc2b440a0, 32'h419dc88c, 32'hc23baff2, 32'hc290d643, 32'hc163058c};
test_output[36976:36983] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h419dc88c, 32'h0, 32'h0, 32'h0};
test_input[36984:36991] = '{32'h419bf338, 32'hc20933d1, 32'hc2a6b60e, 32'h42b47824, 32'h42c502a4, 32'hc24e855f, 32'h4086b45f, 32'h42c268d1};
test_output[36984:36991] = '{32'h419bf338, 32'h0, 32'h0, 32'h42b47824, 32'h42c502a4, 32'h0, 32'h4086b45f, 32'h42c268d1};
test_input[36992:36999] = '{32'hc29430f8, 32'h428012df, 32'hc2b4ac21, 32'h4290a31a, 32'hc22fc511, 32'hc2a283f7, 32'hbfa1faa5, 32'h42b4cc96};
test_output[36992:36999] = '{32'h0, 32'h428012df, 32'h0, 32'h4290a31a, 32'h0, 32'h0, 32'h0, 32'h42b4cc96};
test_input[37000:37007] = '{32'hc1fe2133, 32'h42668334, 32'hc22cb447, 32'hc1c0ea40, 32'hc235b64f, 32'hc0cf43d8, 32'h42920f7a, 32'h41989149};
test_output[37000:37007] = '{32'h0, 32'h42668334, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42920f7a, 32'h41989149};
test_input[37008:37015] = '{32'h42130b34, 32'h4292a129, 32'h41f44cd3, 32'h41117fcc, 32'h42589f8f, 32'h428d3f64, 32'h428bb6dd, 32'h42a34bf0};
test_output[37008:37015] = '{32'h42130b34, 32'h4292a129, 32'h41f44cd3, 32'h41117fcc, 32'h42589f8f, 32'h428d3f64, 32'h428bb6dd, 32'h42a34bf0};
test_input[37016:37023] = '{32'h42551cf6, 32'hc281154f, 32'h429b1e27, 32'hc21b9979, 32'h42b42f67, 32'hc2c2f91e, 32'hc1b1cec9, 32'hc21ae786};
test_output[37016:37023] = '{32'h42551cf6, 32'h0, 32'h429b1e27, 32'h0, 32'h42b42f67, 32'h0, 32'h0, 32'h0};
test_input[37024:37031] = '{32'hc26f0128, 32'h42734b55, 32'h40dc4fc2, 32'hc25be276, 32'hc23fe0c0, 32'hc221308a, 32'hc289a1fe, 32'hc1aa9efc};
test_output[37024:37031] = '{32'h0, 32'h42734b55, 32'h40dc4fc2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[37032:37039] = '{32'hc26e7566, 32'h428ef95b, 32'h423d35e5, 32'h42b2d48f, 32'hc2c1a4e6, 32'h3d66edf7, 32'h42b53bca, 32'hc2052faf};
test_output[37032:37039] = '{32'h0, 32'h428ef95b, 32'h423d35e5, 32'h42b2d48f, 32'h0, 32'h3d66edf7, 32'h42b53bca, 32'h0};
test_input[37040:37047] = '{32'h42a3ad11, 32'h42b51695, 32'h42921e25, 32'hc0d71074, 32'h42a60e56, 32'h40e4f2e8, 32'hc203485c, 32'hc1f4e1b6};
test_output[37040:37047] = '{32'h42a3ad11, 32'h42b51695, 32'h42921e25, 32'h0, 32'h42a60e56, 32'h40e4f2e8, 32'h0, 32'h0};
test_input[37048:37055] = '{32'h42a213e0, 32'hc282db88, 32'h41fe5f31, 32'h4212298f, 32'hc299bf88, 32'hc2a30215, 32'h4265cdca, 32'h411d079c};
test_output[37048:37055] = '{32'h42a213e0, 32'h0, 32'h41fe5f31, 32'h4212298f, 32'h0, 32'h0, 32'h4265cdca, 32'h411d079c};
test_input[37056:37063] = '{32'hbfa51e51, 32'hc282dcfd, 32'hc2c625d5, 32'h42500e08, 32'h42512714, 32'hc223f4bc, 32'hc21955da, 32'hc29e1c72};
test_output[37056:37063] = '{32'h0, 32'h0, 32'h0, 32'h42500e08, 32'h42512714, 32'h0, 32'h0, 32'h0};
test_input[37064:37071] = '{32'hc1b5d0d9, 32'h42a7cc0d, 32'h42bcaa9c, 32'h414bab20, 32'h4211ef36, 32'h42887f17, 32'h4202b6d9, 32'hc2ac8f9e};
test_output[37064:37071] = '{32'h0, 32'h42a7cc0d, 32'h42bcaa9c, 32'h414bab20, 32'h4211ef36, 32'h42887f17, 32'h4202b6d9, 32'h0};
test_input[37072:37079] = '{32'hc2529616, 32'hc225d1f6, 32'h401a19c1, 32'hc2bc7122, 32'hbfc15629, 32'hc2b8d51d, 32'h429dd6dc, 32'h421453b5};
test_output[37072:37079] = '{32'h0, 32'h0, 32'h401a19c1, 32'h0, 32'h0, 32'h0, 32'h429dd6dc, 32'h421453b5};
test_input[37080:37087] = '{32'hc29112ec, 32'h42654fec, 32'h4295a172, 32'hc289a8fe, 32'h424e7946, 32'hc2adb01f, 32'h422b8b89, 32'h42a4d093};
test_output[37080:37087] = '{32'h0, 32'h42654fec, 32'h4295a172, 32'h0, 32'h424e7946, 32'h0, 32'h422b8b89, 32'h42a4d093};
test_input[37088:37095] = '{32'h428b9c4b, 32'hc271f93e, 32'h423a546e, 32'hc296ff34, 32'hc1640c2b, 32'hc26c64f8, 32'hc1d523ae, 32'h4192efbf};
test_output[37088:37095] = '{32'h428b9c4b, 32'h0, 32'h423a546e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4192efbf};
test_input[37096:37103] = '{32'h41a8ed60, 32'h427134b6, 32'h413c1833, 32'hc269f06e, 32'h41dd2b6e, 32'h421592b5, 32'h42a05ee2, 32'hc28e0c28};
test_output[37096:37103] = '{32'h41a8ed60, 32'h427134b6, 32'h413c1833, 32'h0, 32'h41dd2b6e, 32'h421592b5, 32'h42a05ee2, 32'h0};
test_input[37104:37111] = '{32'h4211ad99, 32'h42c21e2a, 32'hc1f83f11, 32'h42c02b3c, 32'h3fd26d07, 32'h42c02e42, 32'hc2615b54, 32'h426c29fd};
test_output[37104:37111] = '{32'h4211ad99, 32'h42c21e2a, 32'h0, 32'h42c02b3c, 32'h3fd26d07, 32'h42c02e42, 32'h0, 32'h426c29fd};
test_input[37112:37119] = '{32'h42888f6e, 32'h425f0c37, 32'hc297be01, 32'h4198dc41, 32'h42320e30, 32'h420b6f44, 32'hc1b4a3cf, 32'h42aa3925};
test_output[37112:37119] = '{32'h42888f6e, 32'h425f0c37, 32'h0, 32'h4198dc41, 32'h42320e30, 32'h420b6f44, 32'h0, 32'h42aa3925};
test_input[37120:37127] = '{32'hc0a55d02, 32'h42b594b6, 32'hc2773328, 32'h427cc463, 32'h412d5528, 32'h41a72857, 32'h422a2eeb, 32'hc2164c32};
test_output[37120:37127] = '{32'h0, 32'h42b594b6, 32'h0, 32'h427cc463, 32'h412d5528, 32'h41a72857, 32'h422a2eeb, 32'h0};
test_input[37128:37135] = '{32'hc0c5df15, 32'hc12b46c7, 32'hc22ac803, 32'h4296eadf, 32'h428ecc4f, 32'h42039cf5, 32'hc29ccf52, 32'h41b13b5a};
test_output[37128:37135] = '{32'h0, 32'h0, 32'h0, 32'h4296eadf, 32'h428ecc4f, 32'h42039cf5, 32'h0, 32'h41b13b5a};
test_input[37136:37143] = '{32'hc2296972, 32'hc2a9e3e6, 32'h419011dc, 32'h40bad8ea, 32'h42aa4669, 32'hc208169f, 32'h424b6fd7, 32'h42934a55};
test_output[37136:37143] = '{32'h0, 32'h0, 32'h419011dc, 32'h40bad8ea, 32'h42aa4669, 32'h0, 32'h424b6fd7, 32'h42934a55};
test_input[37144:37151] = '{32'hc25344de, 32'hc19aa5cd, 32'h42a38267, 32'h4297bd09, 32'h42985e73, 32'h429f27a2, 32'h422a1d68, 32'h42be3e0c};
test_output[37144:37151] = '{32'h0, 32'h0, 32'h42a38267, 32'h4297bd09, 32'h42985e73, 32'h429f27a2, 32'h422a1d68, 32'h42be3e0c};
test_input[37152:37159] = '{32'hc2ac9b08, 32'h408af937, 32'h4220a6b5, 32'h427401ae, 32'hc2c702fa, 32'hc136da10, 32'h41b4b872, 32'hc095f8c0};
test_output[37152:37159] = '{32'h0, 32'h408af937, 32'h4220a6b5, 32'h427401ae, 32'h0, 32'h0, 32'h41b4b872, 32'h0};
test_input[37160:37167] = '{32'hc2af93fe, 32'hc21102bb, 32'h420492a0, 32'h424ac581, 32'hc1119686, 32'h4292a084, 32'h42147828, 32'h4264931a};
test_output[37160:37167] = '{32'h0, 32'h0, 32'h420492a0, 32'h424ac581, 32'h0, 32'h4292a084, 32'h42147828, 32'h4264931a};
test_input[37168:37175] = '{32'hc0c938b0, 32'hc230dd2d, 32'h42a36de3, 32'h412e8587, 32'hc2c7df02, 32'hc2be46e6, 32'hc0d248eb, 32'hc1dbe94d};
test_output[37168:37175] = '{32'h0, 32'h0, 32'h42a36de3, 32'h412e8587, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[37176:37183] = '{32'h42b300f8, 32'h42866be9, 32'h427fc245, 32'h41a7849e, 32'h42c78967, 32'hc141008f, 32'h424f0a18, 32'h42a05c63};
test_output[37176:37183] = '{32'h42b300f8, 32'h42866be9, 32'h427fc245, 32'h41a7849e, 32'h42c78967, 32'h0, 32'h424f0a18, 32'h42a05c63};
test_input[37184:37191] = '{32'h42b9210a, 32'h42887ffb, 32'h42826228, 32'h41e3ccd9, 32'h42223e25, 32'hc2887c4e, 32'hc2b2b02c, 32'hc211a7dc};
test_output[37184:37191] = '{32'h42b9210a, 32'h42887ffb, 32'h42826228, 32'h41e3ccd9, 32'h42223e25, 32'h0, 32'h0, 32'h0};
test_input[37192:37199] = '{32'h4205d967, 32'h425f8ab5, 32'h4291dbde, 32'h42016b81, 32'hc2b1d24c, 32'hbe394c47, 32'h42569635, 32'hc1f26890};
test_output[37192:37199] = '{32'h4205d967, 32'h425f8ab5, 32'h4291dbde, 32'h42016b81, 32'h0, 32'h0, 32'h42569635, 32'h0};
test_input[37200:37207] = '{32'h42c68a3f, 32'h41bf87cb, 32'h42418b79, 32'h41d7898c, 32'h42047148, 32'h42a1431d, 32'hc1c4c259, 32'hc10aea7b};
test_output[37200:37207] = '{32'h42c68a3f, 32'h41bf87cb, 32'h42418b79, 32'h41d7898c, 32'h42047148, 32'h42a1431d, 32'h0, 32'h0};
test_input[37208:37215] = '{32'hc2a59969, 32'hc28506d0, 32'hc2880b11, 32'hc12ff340, 32'hc07d3937, 32'hc0103b74, 32'hc1aa6403, 32'h409c558f};
test_output[37208:37215] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h409c558f};
test_input[37216:37223] = '{32'hc15a5975, 32'h4153c70a, 32'hc18de28b, 32'hc2ad5eb9, 32'h41b7e252, 32'h4244b8a0, 32'h42c5cf95, 32'h429fa296};
test_output[37216:37223] = '{32'h0, 32'h4153c70a, 32'h0, 32'h0, 32'h41b7e252, 32'h4244b8a0, 32'h42c5cf95, 32'h429fa296};
test_input[37224:37231] = '{32'hc1af8b1d, 32'hc18f0c40, 32'h4280204d, 32'hc235ea0f, 32'h4294983d, 32'hc29bce49, 32'hc1a79bc1, 32'hc169bb32};
test_output[37224:37231] = '{32'h0, 32'h0, 32'h4280204d, 32'h0, 32'h4294983d, 32'h0, 32'h0, 32'h0};
test_input[37232:37239] = '{32'h42463d2f, 32'h42066acf, 32'h409fd893, 32'hc1dd0350, 32'h42bac791, 32'hc0238aae, 32'hc199baff, 32'hc22c07e2};
test_output[37232:37239] = '{32'h42463d2f, 32'h42066acf, 32'h409fd893, 32'h0, 32'h42bac791, 32'h0, 32'h0, 32'h0};
test_input[37240:37247] = '{32'h427cb79f, 32'h422d7d59, 32'hc248f5d4, 32'hc0c5cb79, 32'hc24e8ab2, 32'hc28efd42, 32'h429fd39a, 32'hc1bbb37a};
test_output[37240:37247] = '{32'h427cb79f, 32'h422d7d59, 32'h0, 32'h0, 32'h0, 32'h0, 32'h429fd39a, 32'h0};
test_input[37248:37255] = '{32'hc25b1676, 32'h425be550, 32'h412db1ef, 32'h421e551e, 32'hc0a23d56, 32'hc0a4b0dd, 32'h42c0e71b, 32'h4250e246};
test_output[37248:37255] = '{32'h0, 32'h425be550, 32'h412db1ef, 32'h421e551e, 32'h0, 32'h0, 32'h42c0e71b, 32'h4250e246};
test_input[37256:37263] = '{32'hc23ffded, 32'hc2748656, 32'hc0d7d5fd, 32'h41a848f9, 32'hc235587c, 32'h4243fc62, 32'hc230c6b8, 32'h4212ae46};
test_output[37256:37263] = '{32'h0, 32'h0, 32'h0, 32'h41a848f9, 32'h0, 32'h4243fc62, 32'h0, 32'h4212ae46};
test_input[37264:37271] = '{32'h42a714ae, 32'h410f8ea4, 32'h4199362a, 32'h42462682, 32'hc1de5d48, 32'h41fbc28b, 32'hc1989780, 32'hc17063d3};
test_output[37264:37271] = '{32'h42a714ae, 32'h410f8ea4, 32'h4199362a, 32'h42462682, 32'h0, 32'h41fbc28b, 32'h0, 32'h0};
test_input[37272:37279] = '{32'h42596a21, 32'hc2a5aac7, 32'h3fc17c21, 32'hc2a7becc, 32'hc24e8c84, 32'h4268099c, 32'h42982655, 32'h428cc786};
test_output[37272:37279] = '{32'h42596a21, 32'h0, 32'h3fc17c21, 32'h0, 32'h0, 32'h4268099c, 32'h42982655, 32'h428cc786};
test_input[37280:37287] = '{32'h427ec1fc, 32'h40fa4059, 32'hc13c6d8b, 32'h41d8a65d, 32'hc2a899cb, 32'hc2b42c13, 32'h421d7ca6, 32'hc1ffa934};
test_output[37280:37287] = '{32'h427ec1fc, 32'h40fa4059, 32'h0, 32'h41d8a65d, 32'h0, 32'h0, 32'h421d7ca6, 32'h0};
test_input[37288:37295] = '{32'h404b1bcc, 32'hc22cf141, 32'hc27b4f87, 32'h41131da6, 32'hc296af97, 32'hc2b73657, 32'hc2a68f81, 32'h429bc901};
test_output[37288:37295] = '{32'h404b1bcc, 32'h0, 32'h0, 32'h41131da6, 32'h0, 32'h0, 32'h0, 32'h429bc901};
test_input[37296:37303] = '{32'hc29170b0, 32'h42b9bb77, 32'h428d89e6, 32'hc2bcab1d, 32'hc2a43488, 32'hc2944574, 32'h41b022ae, 32'hc2c46812};
test_output[37296:37303] = '{32'h0, 32'h42b9bb77, 32'h428d89e6, 32'h0, 32'h0, 32'h0, 32'h41b022ae, 32'h0};
test_input[37304:37311] = '{32'hc2266382, 32'h4103c937, 32'hc2accd0f, 32'hc2b5f6d5, 32'h417e3f4e, 32'hbfffcae1, 32'hc2856e97, 32'h40c06864};
test_output[37304:37311] = '{32'h0, 32'h4103c937, 32'h0, 32'h0, 32'h417e3f4e, 32'h0, 32'h0, 32'h40c06864};
test_input[37312:37319] = '{32'h410b516e, 32'h427d3e55, 32'h4240766f, 32'h419c12c7, 32'h42ae85c9, 32'h4274a255, 32'hbfa1a0a7, 32'hc2c29711};
test_output[37312:37319] = '{32'h410b516e, 32'h427d3e55, 32'h4240766f, 32'h419c12c7, 32'h42ae85c9, 32'h4274a255, 32'h0, 32'h0};
test_input[37320:37327] = '{32'hc175c4bb, 32'hc2467188, 32'hc147e252, 32'h42c28bae, 32'h414d7e91, 32'hc2a4bdce, 32'hc2a4e920, 32'hc2c676a1};
test_output[37320:37327] = '{32'h0, 32'h0, 32'h0, 32'h42c28bae, 32'h414d7e91, 32'h0, 32'h0, 32'h0};
test_input[37328:37335] = '{32'hc2aef2a8, 32'h422f2520, 32'h425bae98, 32'hc2bd72c8, 32'h4255786b, 32'h42203c9c, 32'hc2bc7e0b, 32'hc2152789};
test_output[37328:37335] = '{32'h0, 32'h422f2520, 32'h425bae98, 32'h0, 32'h4255786b, 32'h42203c9c, 32'h0, 32'h0};
test_input[37336:37343] = '{32'h40cca784, 32'hc24f2681, 32'hc1b346c3, 32'hc229846f, 32'hc2b507d8, 32'h4192b800, 32'h4226137e, 32'h42911ac0};
test_output[37336:37343] = '{32'h40cca784, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4192b800, 32'h4226137e, 32'h42911ac0};
test_input[37344:37351] = '{32'hc1339823, 32'hc17244fa, 32'h425d08ce, 32'h42994bf2, 32'h41f79e17, 32'h411d2534, 32'h42a68fad, 32'hc28ee3d6};
test_output[37344:37351] = '{32'h0, 32'h0, 32'h425d08ce, 32'h42994bf2, 32'h41f79e17, 32'h411d2534, 32'h42a68fad, 32'h0};
test_input[37352:37359] = '{32'h40949852, 32'h42b86e25, 32'h426a2394, 32'hc25d1c5d, 32'h4211c68c, 32'h42011ad5, 32'hc2b86cb8, 32'h419fd63f};
test_output[37352:37359] = '{32'h40949852, 32'h42b86e25, 32'h426a2394, 32'h0, 32'h4211c68c, 32'h42011ad5, 32'h0, 32'h419fd63f};
test_input[37360:37367] = '{32'h42317ed5, 32'hc280950e, 32'h416a65da, 32'h4279b867, 32'h424fe81e, 32'hc19d0e1a, 32'hc2925129, 32'hc24e431e};
test_output[37360:37367] = '{32'h42317ed5, 32'h0, 32'h416a65da, 32'h4279b867, 32'h424fe81e, 32'h0, 32'h0, 32'h0};
test_input[37368:37375] = '{32'hc101f806, 32'h420b6b7c, 32'h42378861, 32'h426c700e, 32'h422f1538, 32'hc263e2bc, 32'h41d074f5, 32'hc21cd269};
test_output[37368:37375] = '{32'h0, 32'h420b6b7c, 32'h42378861, 32'h426c700e, 32'h422f1538, 32'h0, 32'h41d074f5, 32'h0};
test_input[37376:37383] = '{32'hc2a4434f, 32'h41cc390e, 32'h41e6cab7, 32'hc2a9c6fc, 32'h41e5ec05, 32'h427c5e02, 32'hc2adea7f, 32'h4204bb13};
test_output[37376:37383] = '{32'h0, 32'h41cc390e, 32'h41e6cab7, 32'h0, 32'h41e5ec05, 32'h427c5e02, 32'h0, 32'h4204bb13};
test_input[37384:37391] = '{32'h42b38523, 32'hc2881d69, 32'h41c3b9f9, 32'h42584ca4, 32'h426147fe, 32'h4122f5b6, 32'hc2240c45, 32'hc293ea8c};
test_output[37384:37391] = '{32'h42b38523, 32'h0, 32'h41c3b9f9, 32'h42584ca4, 32'h426147fe, 32'h4122f5b6, 32'h0, 32'h0};
test_input[37392:37399] = '{32'hc2a022b0, 32'hc2a9653c, 32'hc28101b1, 32'hc27e5061, 32'hc2877094, 32'h42be84f0, 32'hc1eacc22, 32'hc0dab1a6};
test_output[37392:37399] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42be84f0, 32'h0, 32'h0};
test_input[37400:37407] = '{32'h42a85235, 32'hc158ed37, 32'hc1037b72, 32'h42a37ecb, 32'hc006a9a3, 32'hc1e02698, 32'h428ec1a6, 32'hc263052a};
test_output[37400:37407] = '{32'h42a85235, 32'h0, 32'h0, 32'h42a37ecb, 32'h0, 32'h0, 32'h428ec1a6, 32'h0};
test_input[37408:37415] = '{32'hc2782907, 32'h42c4c1f8, 32'h425fbcf2, 32'hc1d120f3, 32'h4103bad9, 32'h42316a8b, 32'hc2902fe0, 32'h42b90703};
test_output[37408:37415] = '{32'h0, 32'h42c4c1f8, 32'h425fbcf2, 32'h0, 32'h4103bad9, 32'h42316a8b, 32'h0, 32'h42b90703};
test_input[37416:37423] = '{32'hc2b45519, 32'h42b07c23, 32'hc2277d15, 32'h42b2796b, 32'h415aa76a, 32'h42c05796, 32'hc2c769a3, 32'hc12da7b2};
test_output[37416:37423] = '{32'h0, 32'h42b07c23, 32'h0, 32'h42b2796b, 32'h415aa76a, 32'h42c05796, 32'h0, 32'h0};
test_input[37424:37431] = '{32'hc2a41cde, 32'h42705219, 32'h4285b6c3, 32'hc2adc7d5, 32'h428cdcc9, 32'hc20983a7, 32'h41c1dc40, 32'hc292ebcd};
test_output[37424:37431] = '{32'h0, 32'h42705219, 32'h4285b6c3, 32'h0, 32'h428cdcc9, 32'h0, 32'h41c1dc40, 32'h0};
test_input[37432:37439] = '{32'h4260e1a9, 32'hc20634a2, 32'hc2bb323d, 32'hc2493f13, 32'hc2b71f8d, 32'h42a3475b, 32'h4229018d, 32'h41b65603};
test_output[37432:37439] = '{32'h4260e1a9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a3475b, 32'h4229018d, 32'h41b65603};
test_input[37440:37447] = '{32'h41b45318, 32'hc2969419, 32'hc24f61ab, 32'hc1b0f206, 32'h42afdd6d, 32'hc01057c1, 32'hc2a3e758, 32'h42679bde};
test_output[37440:37447] = '{32'h41b45318, 32'h0, 32'h0, 32'h0, 32'h42afdd6d, 32'h0, 32'h0, 32'h42679bde};
test_input[37448:37455] = '{32'h41fdfe58, 32'h40b72461, 32'h4225baef, 32'hc20d6d6d, 32'h427420be, 32'h425fd694, 32'h42bddd04, 32'h4293d351};
test_output[37448:37455] = '{32'h41fdfe58, 32'h40b72461, 32'h4225baef, 32'h0, 32'h427420be, 32'h425fd694, 32'h42bddd04, 32'h4293d351};
test_input[37456:37463] = '{32'hc2a33afa, 32'hc0e58881, 32'h42951d52, 32'hc2462c27, 32'hc22c52a5, 32'hc2913a46, 32'h42447ac5, 32'hc2493ed5};
test_output[37456:37463] = '{32'h0, 32'h0, 32'h42951d52, 32'h0, 32'h0, 32'h0, 32'h42447ac5, 32'h0};
test_input[37464:37471] = '{32'hc2690f0d, 32'h417b3f11, 32'hc29313b5, 32'hc2bd9c00, 32'hc2bea625, 32'h4286431a, 32'h42884242, 32'hc2bffa3e};
test_output[37464:37471] = '{32'h0, 32'h417b3f11, 32'h0, 32'h0, 32'h0, 32'h4286431a, 32'h42884242, 32'h0};
test_input[37472:37479] = '{32'hc060e572, 32'hc2a287f3, 32'h4154f176, 32'hc2b8852e, 32'h42b6a0c6, 32'h429e59e2, 32'h42b50235, 32'hc26cceb9};
test_output[37472:37479] = '{32'h0, 32'h0, 32'h4154f176, 32'h0, 32'h42b6a0c6, 32'h429e59e2, 32'h42b50235, 32'h0};
test_input[37480:37487] = '{32'hc21cd1cd, 32'hc2a28c8f, 32'hc171ece8, 32'hc1e4851f, 32'hc26bf03e, 32'h426ca2d4, 32'h426be319, 32'h428009b3};
test_output[37480:37487] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426ca2d4, 32'h426be319, 32'h428009b3};
test_input[37488:37495] = '{32'h41c7f859, 32'h42908378, 32'hc0ec93ef, 32'h418e973f, 32'h410511bd, 32'hc24991b8, 32'h4249d9f9, 32'hc279a77e};
test_output[37488:37495] = '{32'h41c7f859, 32'h42908378, 32'h0, 32'h418e973f, 32'h410511bd, 32'h0, 32'h4249d9f9, 32'h0};
test_input[37496:37503] = '{32'h41d75fe0, 32'hc1dc15a6, 32'hc23a5e9b, 32'hc2969cb7, 32'hc24a0240, 32'hc26afbe3, 32'h42518ea8, 32'hc0f3aa08};
test_output[37496:37503] = '{32'h41d75fe0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42518ea8, 32'h0};
test_input[37504:37511] = '{32'h4255fff2, 32'h417c7319, 32'h42c0482a, 32'hc1947b8f, 32'h42bb5810, 32'h421a549c, 32'hc24ae8fc, 32'h409047f9};
test_output[37504:37511] = '{32'h4255fff2, 32'h417c7319, 32'h42c0482a, 32'h0, 32'h42bb5810, 32'h421a549c, 32'h0, 32'h409047f9};
test_input[37512:37519] = '{32'h41de5c45, 32'h4297ec4a, 32'hc0d7c011, 32'hc1a21f1b, 32'hc250c945, 32'h4122fbff, 32'h42704303, 32'hc2c7c2fc};
test_output[37512:37519] = '{32'h41de5c45, 32'h4297ec4a, 32'h0, 32'h0, 32'h0, 32'h4122fbff, 32'h42704303, 32'h0};
test_input[37520:37527] = '{32'hc29feaf2, 32'hc2a696cc, 32'h422033de, 32'h41b7d598, 32'h41b01256, 32'h426c0da5, 32'h42a8fd98, 32'h4202e109};
test_output[37520:37527] = '{32'h0, 32'h0, 32'h422033de, 32'h41b7d598, 32'h41b01256, 32'h426c0da5, 32'h42a8fd98, 32'h4202e109};
test_input[37528:37535] = '{32'hc2b1e4cf, 32'h421b06f2, 32'h42b7ca06, 32'h4214276b, 32'h41a66bc5, 32'h41ab8e0d, 32'hc21386e4, 32'hc119a012};
test_output[37528:37535] = '{32'h0, 32'h421b06f2, 32'h42b7ca06, 32'h4214276b, 32'h41a66bc5, 32'h41ab8e0d, 32'h0, 32'h0};
test_input[37536:37543] = '{32'h42b6669e, 32'hc2952e42, 32'hc2921971, 32'h42599167, 32'hc1d4cc65, 32'h42491013, 32'hc16341e2, 32'h425a0bad};
test_output[37536:37543] = '{32'h42b6669e, 32'h0, 32'h0, 32'h42599167, 32'h0, 32'h42491013, 32'h0, 32'h425a0bad};
test_input[37544:37551] = '{32'hc236f61d, 32'hc2a8897b, 32'h41b19440, 32'hc2a223b8, 32'hc17463bc, 32'h416c1e11, 32'h4225cba1, 32'h41c6aa46};
test_output[37544:37551] = '{32'h0, 32'h0, 32'h41b19440, 32'h0, 32'h0, 32'h416c1e11, 32'h4225cba1, 32'h41c6aa46};
test_input[37552:37559] = '{32'h403ec07a, 32'hc20b7022, 32'hc2c3ce8a, 32'h42aa4ac9, 32'h4225cf87, 32'h42287a9d, 32'h4242b458, 32'hc2c649d1};
test_output[37552:37559] = '{32'h403ec07a, 32'h0, 32'h0, 32'h42aa4ac9, 32'h4225cf87, 32'h42287a9d, 32'h4242b458, 32'h0};
test_input[37560:37567] = '{32'h40a10fc5, 32'h41aec5d2, 32'h4291967a, 32'h42794bc5, 32'hc2315577, 32'h4242a5f7, 32'h429d55b9, 32'hc1b3548f};
test_output[37560:37567] = '{32'h40a10fc5, 32'h41aec5d2, 32'h4291967a, 32'h42794bc5, 32'h0, 32'h4242a5f7, 32'h429d55b9, 32'h0};
test_input[37568:37575] = '{32'hc28a5090, 32'h410376a8, 32'h41113511, 32'hc2b23cd8, 32'hc2456269, 32'hc181ee05, 32'h409e01aa, 32'h4283ae7a};
test_output[37568:37575] = '{32'h0, 32'h410376a8, 32'h41113511, 32'h0, 32'h0, 32'h0, 32'h409e01aa, 32'h4283ae7a};
test_input[37576:37583] = '{32'h41f8fb39, 32'h4284ee14, 32'hc260c480, 32'hc21d7c06, 32'h421f4486, 32'h4281456b, 32'hc143bf50, 32'h41f8caf4};
test_output[37576:37583] = '{32'h41f8fb39, 32'h4284ee14, 32'h0, 32'h0, 32'h421f4486, 32'h4281456b, 32'h0, 32'h41f8caf4};
test_input[37584:37591] = '{32'h42c373ab, 32'hc27de41d, 32'h42446d51, 32'hc22c2112, 32'hc1c96a5a, 32'h40c0e3f6, 32'hc1d5fb6e, 32'hc2266f9f};
test_output[37584:37591] = '{32'h42c373ab, 32'h0, 32'h42446d51, 32'h0, 32'h0, 32'h40c0e3f6, 32'h0, 32'h0};
test_input[37592:37599] = '{32'hc035d953, 32'hc019631d, 32'hc2bbb9ef, 32'h42b11f08, 32'h412942d9, 32'hc27ffb8d, 32'h423094ce, 32'hc2c08a97};
test_output[37592:37599] = '{32'h0, 32'h0, 32'h0, 32'h42b11f08, 32'h412942d9, 32'h0, 32'h423094ce, 32'h0};
test_input[37600:37607] = '{32'h408ba098, 32'h429cf598, 32'h41114db1, 32'h41151e35, 32'h42b35cd2, 32'hc11e952b, 32'hbfaf759c, 32'h41a24c20};
test_output[37600:37607] = '{32'h408ba098, 32'h429cf598, 32'h41114db1, 32'h41151e35, 32'h42b35cd2, 32'h0, 32'h0, 32'h41a24c20};
test_input[37608:37615] = '{32'hc1e15896, 32'h4290bc38, 32'h41cc769f, 32'h4232fecd, 32'h4283a6a1, 32'h42c78733, 32'h42a40eb7, 32'h42b2a410};
test_output[37608:37615] = '{32'h0, 32'h4290bc38, 32'h41cc769f, 32'h4232fecd, 32'h4283a6a1, 32'h42c78733, 32'h42a40eb7, 32'h42b2a410};
test_input[37616:37623] = '{32'h41b4c696, 32'h42827196, 32'h42b75cce, 32'hc1d9c70d, 32'hc0aa826f, 32'hc2aaacd9, 32'h41ab71fd, 32'h415e4144};
test_output[37616:37623] = '{32'h41b4c696, 32'h42827196, 32'h42b75cce, 32'h0, 32'h0, 32'h0, 32'h41ab71fd, 32'h415e4144};
test_input[37624:37631] = '{32'hc25a4a40, 32'h42443f32, 32'h42bee132, 32'hc15ce18b, 32'h425f9294, 32'h41d502b5, 32'h425e357b, 32'h42b6b523};
test_output[37624:37631] = '{32'h0, 32'h42443f32, 32'h42bee132, 32'h0, 32'h425f9294, 32'h41d502b5, 32'h425e357b, 32'h42b6b523};
test_input[37632:37639] = '{32'h41b2eefa, 32'h4196f5b0, 32'h427883c8, 32'hc24a4c14, 32'h41af6329, 32'h41c2d78c, 32'hc1549f98, 32'h4270ca7c};
test_output[37632:37639] = '{32'h41b2eefa, 32'h4196f5b0, 32'h427883c8, 32'h0, 32'h41af6329, 32'h41c2d78c, 32'h0, 32'h4270ca7c};
test_input[37640:37647] = '{32'h4017e1ab, 32'h42ae26fd, 32'h429a2727, 32'h429c68c2, 32'h42a2366d, 32'h426fc091, 32'hc2a9343c, 32'hc27472ab};
test_output[37640:37647] = '{32'h4017e1ab, 32'h42ae26fd, 32'h429a2727, 32'h429c68c2, 32'h42a2366d, 32'h426fc091, 32'h0, 32'h0};
test_input[37648:37655] = '{32'hc282b217, 32'h42896288, 32'h41a1a331, 32'hc2607ba2, 32'h42bb483a, 32'hc2802ea8, 32'hc1bae7b1, 32'hbf1980d6};
test_output[37648:37655] = '{32'h0, 32'h42896288, 32'h41a1a331, 32'h0, 32'h42bb483a, 32'h0, 32'h0, 32'h0};
test_input[37656:37663] = '{32'hc1865edd, 32'h41111281, 32'hc28a03fd, 32'h426c573d, 32'h42be6778, 32'h4298aab2, 32'hc2863405, 32'h421ba17b};
test_output[37656:37663] = '{32'h0, 32'h41111281, 32'h0, 32'h426c573d, 32'h42be6778, 32'h4298aab2, 32'h0, 32'h421ba17b};
test_input[37664:37671] = '{32'h425b72ec, 32'h4289884d, 32'hc19f0d57, 32'h415efc33, 32'hc2591645, 32'hc26f1e76, 32'hc150cd37, 32'h42c711d3};
test_output[37664:37671] = '{32'h425b72ec, 32'h4289884d, 32'h0, 32'h415efc33, 32'h0, 32'h0, 32'h0, 32'h42c711d3};
test_input[37672:37679] = '{32'h41b167e4, 32'hc284b247, 32'hc00d2ee6, 32'hc2ae4ce7, 32'h42b5c0b4, 32'h4024670a, 32'hc1a5e0d4, 32'hc1d1fa84};
test_output[37672:37679] = '{32'h41b167e4, 32'h0, 32'h0, 32'h0, 32'h42b5c0b4, 32'h4024670a, 32'h0, 32'h0};
test_input[37680:37687] = '{32'hc29ba555, 32'h4066ff61, 32'hc2344968, 32'h4288cfd5, 32'h42a67f84, 32'h42bd2016, 32'h428c4842, 32'hc1d465be};
test_output[37680:37687] = '{32'h0, 32'h4066ff61, 32'h0, 32'h4288cfd5, 32'h42a67f84, 32'h42bd2016, 32'h428c4842, 32'h0};
test_input[37688:37695] = '{32'h422f2c7a, 32'h4270d183, 32'hc2530086, 32'h42c52a3d, 32'h42c6836c, 32'h427d225c, 32'hc26b78f1, 32'h4297d45c};
test_output[37688:37695] = '{32'h422f2c7a, 32'h4270d183, 32'h0, 32'h42c52a3d, 32'h42c6836c, 32'h427d225c, 32'h0, 32'h4297d45c};
test_input[37696:37703] = '{32'hc05d4faa, 32'h42bed4d3, 32'h422dedab, 32'h418b2a63, 32'h42961af6, 32'h403f1fed, 32'h429760ef, 32'h429c6b88};
test_output[37696:37703] = '{32'h0, 32'h42bed4d3, 32'h422dedab, 32'h418b2a63, 32'h42961af6, 32'h403f1fed, 32'h429760ef, 32'h429c6b88};
test_input[37704:37711] = '{32'hc27759df, 32'hc29f1b8c, 32'h4110c573, 32'h4217b619, 32'hc2af5439, 32'hc290221e, 32'h4080d3c1, 32'hc2957924};
test_output[37704:37711] = '{32'h0, 32'h0, 32'h4110c573, 32'h4217b619, 32'h0, 32'h0, 32'h4080d3c1, 32'h0};
test_input[37712:37719] = '{32'h42b14040, 32'h420f0be0, 32'h41167b6b, 32'h429fe451, 32'hc19e1124, 32'hc067df1b, 32'hc2be82a3, 32'hc16e51aa};
test_output[37712:37719] = '{32'h42b14040, 32'h420f0be0, 32'h41167b6b, 32'h429fe451, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[37720:37727] = '{32'h420f48e9, 32'hc2246294, 32'hc2c6006d, 32'h41643df2, 32'hc1b76dac, 32'h4274e65b, 32'h4268db8f, 32'hc2642e7d};
test_output[37720:37727] = '{32'h420f48e9, 32'h0, 32'h0, 32'h41643df2, 32'h0, 32'h4274e65b, 32'h4268db8f, 32'h0};
test_input[37728:37735] = '{32'h3fac274a, 32'hc264e516, 32'h40864c7b, 32'hc22a3468, 32'hc280f4a3, 32'h41dfb07f, 32'h42aeb7b9, 32'h42be9b94};
test_output[37728:37735] = '{32'h3fac274a, 32'h0, 32'h40864c7b, 32'h0, 32'h0, 32'h41dfb07f, 32'h42aeb7b9, 32'h42be9b94};
test_input[37736:37743] = '{32'h41ffdc5e, 32'h42b38832, 32'h42517435, 32'hbf81c2c4, 32'h42aa39c7, 32'h428120f2, 32'h428997a2, 32'hc1e27cb2};
test_output[37736:37743] = '{32'h41ffdc5e, 32'h42b38832, 32'h42517435, 32'h0, 32'h42aa39c7, 32'h428120f2, 32'h428997a2, 32'h0};
test_input[37744:37751] = '{32'hc0d05829, 32'h4295e811, 32'h42a45e3f, 32'hc23ae73c, 32'hc2920303, 32'hc202fb6c, 32'h428f3c49, 32'h40d736f3};
test_output[37744:37751] = '{32'h0, 32'h4295e811, 32'h42a45e3f, 32'h0, 32'h0, 32'h0, 32'h428f3c49, 32'h40d736f3};
test_input[37752:37759] = '{32'hc20b6f0f, 32'hc26e0a8f, 32'h416e19ee, 32'h41bdd82a, 32'hc18fc49e, 32'hc26c2946, 32'hc2bf0bf4, 32'hc18fab76};
test_output[37752:37759] = '{32'h0, 32'h0, 32'h416e19ee, 32'h41bdd82a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[37760:37767] = '{32'hc1845117, 32'h4236ac7b, 32'h417ccb7b, 32'h41f3ee9f, 32'hc1eb4ebb, 32'h42950c53, 32'hc18ab64e, 32'h425c8619};
test_output[37760:37767] = '{32'h0, 32'h4236ac7b, 32'h417ccb7b, 32'h41f3ee9f, 32'h0, 32'h42950c53, 32'h0, 32'h425c8619};
test_input[37768:37775] = '{32'h42933d41, 32'h40a8b242, 32'hc28fcebd, 32'h41674205, 32'h4242978d, 32'hc23657d3, 32'h426a90e4, 32'h4277df98};
test_output[37768:37775] = '{32'h42933d41, 32'h40a8b242, 32'h0, 32'h41674205, 32'h4242978d, 32'h0, 32'h426a90e4, 32'h4277df98};
test_input[37776:37783] = '{32'h41d3d501, 32'h417e2416, 32'hc125b929, 32'hc2aa308c, 32'hbfdd9fb5, 32'h4185d5cb, 32'hc1e166ad, 32'hc22ae10b};
test_output[37776:37783] = '{32'h41d3d501, 32'h417e2416, 32'h0, 32'h0, 32'h0, 32'h4185d5cb, 32'h0, 32'h0};
test_input[37784:37791] = '{32'h429e3cf0, 32'hc203ead5, 32'h42938dfc, 32'h400c02d8, 32'hc2847bd8, 32'hc2b5dce0, 32'hc29f7f72, 32'hc2330cae};
test_output[37784:37791] = '{32'h429e3cf0, 32'h0, 32'h42938dfc, 32'h400c02d8, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[37792:37799] = '{32'hc1b0aac9, 32'h42a1fef6, 32'h422def94, 32'hc260ec19, 32'hc0b3eb47, 32'hc29778e8, 32'hc21aa10c, 32'h3fee1927};
test_output[37792:37799] = '{32'h0, 32'h42a1fef6, 32'h422def94, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3fee1927};
test_input[37800:37807] = '{32'h4292c72a, 32'h423d8577, 32'hc15b72e6, 32'hc05d0c6c, 32'h4268014e, 32'h4293f6ea, 32'hc29f8afa, 32'hc24f3739};
test_output[37800:37807] = '{32'h4292c72a, 32'h423d8577, 32'h0, 32'h0, 32'h4268014e, 32'h4293f6ea, 32'h0, 32'h0};
test_input[37808:37815] = '{32'hc070d466, 32'h4117fd4c, 32'h42443ac5, 32'h3facb691, 32'hc1412d25, 32'hc2441276, 32'hc2819fec, 32'h41811a49};
test_output[37808:37815] = '{32'h0, 32'h4117fd4c, 32'h42443ac5, 32'h3facb691, 32'h0, 32'h0, 32'h0, 32'h41811a49};
test_input[37816:37823] = '{32'hc21e8f7f, 32'h40779d68, 32'hc1ecae35, 32'h40b864f7, 32'hc20e93de, 32'h40c6e455, 32'h41bf954e, 32'h429ea6f7};
test_output[37816:37823] = '{32'h0, 32'h40779d68, 32'h0, 32'h40b864f7, 32'h0, 32'h40c6e455, 32'h41bf954e, 32'h429ea6f7};
test_input[37824:37831] = '{32'h4239e245, 32'h42b417ef, 32'h421afb95, 32'h42b3e37c, 32'hc1d2f5e3, 32'hc1ad00c3, 32'hc1d33f8f, 32'hc228e4f3};
test_output[37824:37831] = '{32'h4239e245, 32'h42b417ef, 32'h421afb95, 32'h42b3e37c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[37832:37839] = '{32'hc2114004, 32'h42221126, 32'hc0cc33ab, 32'h423e4e92, 32'hc2bd35f6, 32'hc136c65a, 32'h421b73f4, 32'hc2bbbd38};
test_output[37832:37839] = '{32'h0, 32'h42221126, 32'h0, 32'h423e4e92, 32'h0, 32'h0, 32'h421b73f4, 32'h0};
test_input[37840:37847] = '{32'hc24d7ae4, 32'h41fa50d3, 32'hbf2a6373, 32'h42b8bdb9, 32'hc2977245, 32'h41fcc8ec, 32'h42044f40, 32'h40a3a549};
test_output[37840:37847] = '{32'h0, 32'h41fa50d3, 32'h0, 32'h42b8bdb9, 32'h0, 32'h41fcc8ec, 32'h42044f40, 32'h40a3a549};
test_input[37848:37855] = '{32'hc21eeba3, 32'hc20fc4a9, 32'h427fe6cc, 32'h42aee352, 32'hc2490a20, 32'h42523936, 32'hc1f6c569, 32'h41c67aac};
test_output[37848:37855] = '{32'h0, 32'h0, 32'h427fe6cc, 32'h42aee352, 32'h0, 32'h42523936, 32'h0, 32'h41c67aac};
test_input[37856:37863] = '{32'hc28bd596, 32'hc103e10d, 32'h42a4a042, 32'h41f6f409, 32'hc096b293, 32'hc2ba6b15, 32'h42bfae9c, 32'h42aa25a8};
test_output[37856:37863] = '{32'h0, 32'h0, 32'h42a4a042, 32'h41f6f409, 32'h0, 32'h0, 32'h42bfae9c, 32'h42aa25a8};
test_input[37864:37871] = '{32'h42bc3d63, 32'hc2624179, 32'h411eeeba, 32'h4219df20, 32'h40915aca, 32'h42c0464d, 32'hc278d269, 32'hc2c47616};
test_output[37864:37871] = '{32'h42bc3d63, 32'h0, 32'h411eeeba, 32'h4219df20, 32'h40915aca, 32'h42c0464d, 32'h0, 32'h0};
test_input[37872:37879] = '{32'hc2466bd1, 32'hc2409d52, 32'hc19c4fb3, 32'hc088eb5b, 32'hc01ffa86, 32'hc060c87d, 32'h4277d61c, 32'hc290c568};
test_output[37872:37879] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4277d61c, 32'h0};
test_input[37880:37887] = '{32'h416eeddc, 32'hc26db626, 32'hc27cddc4, 32'hc2744b2d, 32'h42896d03, 32'h4258cfbe, 32'hc1d64246, 32'h4296eb71};
test_output[37880:37887] = '{32'h416eeddc, 32'h0, 32'h0, 32'h0, 32'h42896d03, 32'h4258cfbe, 32'h0, 32'h4296eb71};
test_input[37888:37895] = '{32'h4218958b, 32'h4219ad24, 32'h41c1e176, 32'hc277b469, 32'h42933167, 32'hc268191c, 32'hc28824ce, 32'hc29d8de8};
test_output[37888:37895] = '{32'h4218958b, 32'h4219ad24, 32'h41c1e176, 32'h0, 32'h42933167, 32'h0, 32'h0, 32'h0};
test_input[37896:37903] = '{32'hc09e7d59, 32'hc26238a0, 32'h42b7f6bf, 32'h42a3395e, 32'h42aca4f9, 32'h40dd630c, 32'hc2a63a23, 32'h42251257};
test_output[37896:37903] = '{32'h0, 32'h0, 32'h42b7f6bf, 32'h42a3395e, 32'h42aca4f9, 32'h40dd630c, 32'h0, 32'h42251257};
test_input[37904:37911] = '{32'h4188f3b6, 32'h42952256, 32'h429cab87, 32'h40e113b1, 32'h426fde91, 32'h41fba361, 32'h4207dbbe, 32'hc207f5df};
test_output[37904:37911] = '{32'h4188f3b6, 32'h42952256, 32'h429cab87, 32'h40e113b1, 32'h426fde91, 32'h41fba361, 32'h4207dbbe, 32'h0};
test_input[37912:37919] = '{32'h42520d13, 32'h4284d2fe, 32'hc219cd51, 32'h41a66b79, 32'h426d851b, 32'h422c0f88, 32'hc1af7b0c, 32'h40c24eab};
test_output[37912:37919] = '{32'h42520d13, 32'h4284d2fe, 32'h0, 32'h41a66b79, 32'h426d851b, 32'h422c0f88, 32'h0, 32'h40c24eab};
test_input[37920:37927] = '{32'h4034f524, 32'h420aab4f, 32'h42859d64, 32'hc1afc765, 32'h4048fad1, 32'h4218760f, 32'h422e9f29, 32'h41c9509b};
test_output[37920:37927] = '{32'h4034f524, 32'h420aab4f, 32'h42859d64, 32'h0, 32'h4048fad1, 32'h4218760f, 32'h422e9f29, 32'h41c9509b};
test_input[37928:37935] = '{32'hc270a634, 32'hc0f694a6, 32'h41d85e21, 32'h423f709d, 32'hc1b4719d, 32'h42a1e179, 32'h42b648be, 32'hc25288c5};
test_output[37928:37935] = '{32'h0, 32'h0, 32'h41d85e21, 32'h423f709d, 32'h0, 32'h42a1e179, 32'h42b648be, 32'h0};
test_input[37936:37943] = '{32'h42afffcd, 32'h423ddb50, 32'h42135d53, 32'h418515c8, 32'hc28f01ef, 32'hc1e8e92d, 32'h41f9ad24, 32'h41d705a3};
test_output[37936:37943] = '{32'h42afffcd, 32'h423ddb50, 32'h42135d53, 32'h418515c8, 32'h0, 32'h0, 32'h41f9ad24, 32'h41d705a3};
test_input[37944:37951] = '{32'h426d0fc3, 32'hc0bf5ab0, 32'hc2bf62fe, 32'h42b456d2, 32'hc2ad7074, 32'h42b44c55, 32'hc2c5c9ab, 32'h4200bd14};
test_output[37944:37951] = '{32'h426d0fc3, 32'h0, 32'h0, 32'h42b456d2, 32'h0, 32'h42b44c55, 32'h0, 32'h4200bd14};
test_input[37952:37959] = '{32'hc2435269, 32'h42984207, 32'h42991dca, 32'h41cef9ba, 32'hc14599f3, 32'hc19edcad, 32'h419a1832, 32'h427cd637};
test_output[37952:37959] = '{32'h0, 32'h42984207, 32'h42991dca, 32'h41cef9ba, 32'h0, 32'h0, 32'h419a1832, 32'h427cd637};
test_input[37960:37967] = '{32'hc04d88f0, 32'hc2aac46e, 32'h421ddabd, 32'h42a105d5, 32'h42a50855, 32'h3ebcd7d3, 32'hc2af9604, 32'hc1eef071};
test_output[37960:37967] = '{32'h0, 32'h0, 32'h421ddabd, 32'h42a105d5, 32'h42a50855, 32'h3ebcd7d3, 32'h0, 32'h0};
test_input[37968:37975] = '{32'h426a7767, 32'h41fbea3c, 32'h42a33772, 32'hc1454bfa, 32'h4083c782, 32'hc2b46630, 32'h42945a09, 32'hc205e9ad};
test_output[37968:37975] = '{32'h426a7767, 32'h41fbea3c, 32'h42a33772, 32'h0, 32'h4083c782, 32'h0, 32'h42945a09, 32'h0};
test_input[37976:37983] = '{32'h429f677d, 32'hc2a9bd97, 32'h40324513, 32'hc136ec88, 32'h4192e55e, 32'hc1a71e74, 32'h42b65423, 32'hc2a6e027};
test_output[37976:37983] = '{32'h429f677d, 32'h0, 32'h40324513, 32'h0, 32'h4192e55e, 32'h0, 32'h42b65423, 32'h0};
test_input[37984:37991] = '{32'h42c7acee, 32'h421e1841, 32'h4177eb72, 32'h426a40d6, 32'h4255a5ac, 32'hc2a3a80e, 32'h4100ae6c, 32'hc20c06c0};
test_output[37984:37991] = '{32'h42c7acee, 32'h421e1841, 32'h4177eb72, 32'h426a40d6, 32'h4255a5ac, 32'h0, 32'h4100ae6c, 32'h0};
test_input[37992:37999] = '{32'h4254938e, 32'hc23bc2f1, 32'h428a4e12, 32'h41ec8e4c, 32'hc126fb08, 32'hc22c020c, 32'h421b1579, 32'hc2a285bb};
test_output[37992:37999] = '{32'h4254938e, 32'h0, 32'h428a4e12, 32'h41ec8e4c, 32'h0, 32'h0, 32'h421b1579, 32'h0};
test_input[38000:38007] = '{32'h42b43d5c, 32'h418ff669, 32'h42b2041f, 32'hc2748da7, 32'h42a4154f, 32'hc179d2d0, 32'hc19a4cab, 32'h4231b4f0};
test_output[38000:38007] = '{32'h42b43d5c, 32'h418ff669, 32'h42b2041f, 32'h0, 32'h42a4154f, 32'h0, 32'h0, 32'h4231b4f0};
test_input[38008:38015] = '{32'h42148f66, 32'hc16d3e80, 32'h42c3dfa5, 32'h4287f304, 32'h42056732, 32'hc20f1a66, 32'h420e4eb5, 32'h4292db45};
test_output[38008:38015] = '{32'h42148f66, 32'h0, 32'h42c3dfa5, 32'h4287f304, 32'h42056732, 32'h0, 32'h420e4eb5, 32'h4292db45};
test_input[38016:38023] = '{32'h41fcf9d4, 32'hc26ea8ff, 32'hc25baa83, 32'hc1ca8e18, 32'h42163e06, 32'hc1b155cc, 32'h428084d7, 32'hc212702b};
test_output[38016:38023] = '{32'h41fcf9d4, 32'h0, 32'h0, 32'h0, 32'h42163e06, 32'h0, 32'h428084d7, 32'h0};
test_input[38024:38031] = '{32'h42b6a497, 32'hbf52ee19, 32'hc29afe4b, 32'hc2c1d179, 32'h419d1ba6, 32'h4280260b, 32'h427f6e72, 32'hc1ad0502};
test_output[38024:38031] = '{32'h42b6a497, 32'h0, 32'h0, 32'h0, 32'h419d1ba6, 32'h4280260b, 32'h427f6e72, 32'h0};
test_input[38032:38039] = '{32'h40f466ae, 32'hc276fe3e, 32'hc26b1bbb, 32'h42003826, 32'h41a9612d, 32'hc2019dde, 32'h411eb1cf, 32'h42bbae8f};
test_output[38032:38039] = '{32'h40f466ae, 32'h0, 32'h0, 32'h42003826, 32'h41a9612d, 32'h0, 32'h411eb1cf, 32'h42bbae8f};
test_input[38040:38047] = '{32'h41a6c09b, 32'hc29a708c, 32'hc1f77327, 32'h423f772f, 32'hc2869c56, 32'hc1f765ea, 32'h42b1788a, 32'h42c28560};
test_output[38040:38047] = '{32'h41a6c09b, 32'h0, 32'h0, 32'h423f772f, 32'h0, 32'h0, 32'h42b1788a, 32'h42c28560};
test_input[38048:38055] = '{32'h42bbc1df, 32'hc1cc7ea3, 32'h422295a8, 32'hc2c7e88c, 32'hc193e4ba, 32'hc134414c, 32'h421dc73f, 32'h426f6684};
test_output[38048:38055] = '{32'h42bbc1df, 32'h0, 32'h422295a8, 32'h0, 32'h0, 32'h0, 32'h421dc73f, 32'h426f6684};
test_input[38056:38063] = '{32'h42a7cd9d, 32'hc2c315d8, 32'hc21e1547, 32'h419f547a, 32'hc26665c2, 32'hc2ba696b, 32'hc1ebafcf, 32'hc2044a78};
test_output[38056:38063] = '{32'h42a7cd9d, 32'h0, 32'h0, 32'h419f547a, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[38064:38071] = '{32'hc23e17fd, 32'h425957a4, 32'h42a53746, 32'hc29973a5, 32'h429d6ec3, 32'hc1945302, 32'h42891405, 32'h429de97a};
test_output[38064:38071] = '{32'h0, 32'h425957a4, 32'h42a53746, 32'h0, 32'h429d6ec3, 32'h0, 32'h42891405, 32'h429de97a};
test_input[38072:38079] = '{32'hc1e784c0, 32'h421849c3, 32'h42bcd09f, 32'h4254c316, 32'h4266a743, 32'hc2a24237, 32'h4263c5b3, 32'h419370ff};
test_output[38072:38079] = '{32'h0, 32'h421849c3, 32'h42bcd09f, 32'h4254c316, 32'h4266a743, 32'h0, 32'h4263c5b3, 32'h419370ff};
test_input[38080:38087] = '{32'hc2823f9a, 32'h41eaf209, 32'hc2a6101e, 32'hc10a4e1b, 32'hc01d1485, 32'hc1c4f8e4, 32'h4252edcd, 32'h40fa02d1};
test_output[38080:38087] = '{32'h0, 32'h41eaf209, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4252edcd, 32'h40fa02d1};
test_input[38088:38095] = '{32'hc1079a6d, 32'hc23c85ff, 32'h41ed2e48, 32'hc290213a, 32'hc234f65c, 32'hc2be9aa5, 32'h410b3778, 32'hc1519c61};
test_output[38088:38095] = '{32'h0, 32'h0, 32'h41ed2e48, 32'h0, 32'h0, 32'h0, 32'h410b3778, 32'h0};
test_input[38096:38103] = '{32'h411035d8, 32'hc2b8d464, 32'hc2a8ad7d, 32'h42c55b7e, 32'h4281bc61, 32'h421c0d89, 32'hc28ac78d, 32'h4298424d};
test_output[38096:38103] = '{32'h411035d8, 32'h0, 32'h0, 32'h42c55b7e, 32'h4281bc61, 32'h421c0d89, 32'h0, 32'h4298424d};
test_input[38104:38111] = '{32'hc2aa0456, 32'hc208b1f5, 32'hc1a91bc1, 32'h420591bb, 32'h4199c489, 32'h428cfd3f, 32'h4283c270, 32'h42a60db4};
test_output[38104:38111] = '{32'h0, 32'h0, 32'h0, 32'h420591bb, 32'h4199c489, 32'h428cfd3f, 32'h4283c270, 32'h42a60db4};
test_input[38112:38119] = '{32'hc1ef6442, 32'h4289fa04, 32'h40658c38, 32'h42197a9f, 32'hbfdd7a47, 32'h41817301, 32'hc2432e5e, 32'hc2b753db};
test_output[38112:38119] = '{32'h0, 32'h4289fa04, 32'h40658c38, 32'h42197a9f, 32'h0, 32'h41817301, 32'h0, 32'h0};
test_input[38120:38127] = '{32'hc14c8f6b, 32'hc19aa812, 32'h42c23670, 32'hc1fc04b4, 32'hc2279cb7, 32'hc1e31b64, 32'hc290598b, 32'hc2606435};
test_output[38120:38127] = '{32'h0, 32'h0, 32'h42c23670, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[38128:38135] = '{32'hc1ff6bc2, 32'hc2825201, 32'h42c7372c, 32'h4238e02b, 32'hc2592248, 32'h42871852, 32'h429e5f89, 32'h4215d719};
test_output[38128:38135] = '{32'h0, 32'h0, 32'h42c7372c, 32'h4238e02b, 32'h0, 32'h42871852, 32'h429e5f89, 32'h4215d719};
test_input[38136:38143] = '{32'hc295855e, 32'hc287a743, 32'hc161164f, 32'h40ac8273, 32'hc0c30dae, 32'h42693921, 32'hc2ade2df, 32'hc2190ce8};
test_output[38136:38143] = '{32'h0, 32'h0, 32'h0, 32'h40ac8273, 32'h0, 32'h42693921, 32'h0, 32'h0};
test_input[38144:38151] = '{32'hbfa32caa, 32'h4294440a, 32'hbfa8044a, 32'h42a2ca87, 32'h4276dacb, 32'hc2b695af, 32'h42b47036, 32'h42298d36};
test_output[38144:38151] = '{32'h0, 32'h4294440a, 32'h0, 32'h42a2ca87, 32'h4276dacb, 32'h0, 32'h42b47036, 32'h42298d36};
test_input[38152:38159] = '{32'h426500b8, 32'h4122c5c2, 32'hc1532d94, 32'hc1b3cc58, 32'hc287099c, 32'hc2490911, 32'hc28e4b4e, 32'hc27436c6};
test_output[38152:38159] = '{32'h426500b8, 32'h4122c5c2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[38160:38167] = '{32'h4237ed49, 32'hc2bf6c85, 32'hc1e7a827, 32'h42b0938a, 32'h41dfef3c, 32'hc1f49c31, 32'hc283b8a1, 32'hc250d633};
test_output[38160:38167] = '{32'h4237ed49, 32'h0, 32'h0, 32'h42b0938a, 32'h41dfef3c, 32'h0, 32'h0, 32'h0};
test_input[38168:38175] = '{32'hc28ef5fe, 32'hc2abe537, 32'h4296a35b, 32'h42b8dd60, 32'h4116fddf, 32'hc27d1feb, 32'hc2c21fc6, 32'hc2b23e4a};
test_output[38168:38175] = '{32'h0, 32'h0, 32'h4296a35b, 32'h42b8dd60, 32'h4116fddf, 32'h0, 32'h0, 32'h0};
test_input[38176:38183] = '{32'hc10c1103, 32'h41ed8087, 32'h427711b7, 32'h41272d8c, 32'hc2b89dc7, 32'h42b3e855, 32'hc2beb436, 32'h42819d30};
test_output[38176:38183] = '{32'h0, 32'h41ed8087, 32'h427711b7, 32'h41272d8c, 32'h0, 32'h42b3e855, 32'h0, 32'h42819d30};
test_input[38184:38191] = '{32'hc2b02b5f, 32'hc2b4f6dc, 32'hc1a4aebb, 32'hc1216666, 32'hc27a2887, 32'h3f5f7272, 32'h42bf4686, 32'h421f9c77};
test_output[38184:38191] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3f5f7272, 32'h42bf4686, 32'h421f9c77};
test_input[38192:38199] = '{32'hc100dca8, 32'h41b90869, 32'h41eeadf5, 32'h41911740, 32'hbfbec9f8, 32'h41d885b2, 32'hc2099aa7, 32'hc1ddbd2d};
test_output[38192:38199] = '{32'h0, 32'h41b90869, 32'h41eeadf5, 32'h41911740, 32'h0, 32'h41d885b2, 32'h0, 32'h0};
test_input[38200:38207] = '{32'hc17b8094, 32'h422a3f6f, 32'hc28e2911, 32'hc26f9a65, 32'hc13f4acb, 32'hc284e067, 32'hc1f1c3d6, 32'hc22e2151};
test_output[38200:38207] = '{32'h0, 32'h422a3f6f, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[38208:38215] = '{32'hc26764b2, 32'h42145944, 32'hc222b8b5, 32'h41162c69, 32'h427de35a, 32'h424a5301, 32'h427e5b58, 32'h42c34c89};
test_output[38208:38215] = '{32'h0, 32'h42145944, 32'h0, 32'h41162c69, 32'h427de35a, 32'h424a5301, 32'h427e5b58, 32'h42c34c89};
test_input[38216:38223] = '{32'h4110449d, 32'hc2be83ff, 32'hc205d040, 32'h42c56088, 32'h40dba1de, 32'hc1d7f151, 32'hc218b81b, 32'h421d199a};
test_output[38216:38223] = '{32'h4110449d, 32'h0, 32'h0, 32'h42c56088, 32'h40dba1de, 32'h0, 32'h0, 32'h421d199a};
test_input[38224:38231] = '{32'hc23b8bb3, 32'h42ad05c7, 32'h4117ad76, 32'h4262086f, 32'hc10cce86, 32'h42a41d7a, 32'h4266a769, 32'hc2583d3b};
test_output[38224:38231] = '{32'h0, 32'h42ad05c7, 32'h4117ad76, 32'h4262086f, 32'h0, 32'h42a41d7a, 32'h4266a769, 32'h0};
test_input[38232:38239] = '{32'hc27fc7ad, 32'h42af7fb7, 32'h42a0778f, 32'h42c1a670, 32'h42a56b40, 32'h41e56e55, 32'hc27d5935, 32'h42bc10f1};
test_output[38232:38239] = '{32'h0, 32'h42af7fb7, 32'h42a0778f, 32'h42c1a670, 32'h42a56b40, 32'h41e56e55, 32'h0, 32'h42bc10f1};
test_input[38240:38247] = '{32'hc24dc9fb, 32'h41fdd8b9, 32'hc24f8759, 32'hc248465f, 32'hc2a7eb60, 32'hc234b234, 32'hc2b63ae5, 32'hc2c635ae};
test_output[38240:38247] = '{32'h0, 32'h41fdd8b9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[38248:38255] = '{32'h414dd684, 32'h4296500e, 32'hc0cc6e74, 32'h424a0b26, 32'hc277565a, 32'h428dda87, 32'h427846f6, 32'hc2bde65f};
test_output[38248:38255] = '{32'h414dd684, 32'h4296500e, 32'h0, 32'h424a0b26, 32'h0, 32'h428dda87, 32'h427846f6, 32'h0};
test_input[38256:38263] = '{32'hc1ec321d, 32'h413dce80, 32'hc29f97a6, 32'h42bab16a, 32'hc24c8c31, 32'h428e6cb5, 32'h4235d30a, 32'hc2bd0939};
test_output[38256:38263] = '{32'h0, 32'h413dce80, 32'h0, 32'h42bab16a, 32'h0, 32'h428e6cb5, 32'h4235d30a, 32'h0};
test_input[38264:38271] = '{32'hc1817a6d, 32'hc29a6dc7, 32'hc222d9fb, 32'hc287f0e2, 32'hc026cf73, 32'hc21d4a63, 32'h4200cae8, 32'hc20d99a1};
test_output[38264:38271] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4200cae8, 32'h0};
test_input[38272:38279] = '{32'hc2a80731, 32'h424d72fe, 32'hc28a7ccf, 32'hc1ee9423, 32'hc243e9cc, 32'h42a774ab, 32'hc2189f27, 32'hc19c7cca};
test_output[38272:38279] = '{32'h0, 32'h424d72fe, 32'h0, 32'h0, 32'h0, 32'h42a774ab, 32'h0, 32'h0};
test_input[38280:38287] = '{32'hc28ed5a7, 32'hc2b26150, 32'hc2b3c704, 32'hc2312827, 32'hc2b46c28, 32'h4182a9ac, 32'h418fbac6, 32'h42ab0988};
test_output[38280:38287] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4182a9ac, 32'h418fbac6, 32'h42ab0988};
test_input[38288:38295] = '{32'h429c0f73, 32'h4201424b, 32'hc294fedf, 32'hc2a8d057, 32'h4085082a, 32'h4282c7de, 32'h42a42a11, 32'hc1f8728c};
test_output[38288:38295] = '{32'h429c0f73, 32'h4201424b, 32'h0, 32'h0, 32'h4085082a, 32'h4282c7de, 32'h42a42a11, 32'h0};
test_input[38296:38303] = '{32'h42679e1d, 32'hc241bb46, 32'h40c0d114, 32'hc2af3138, 32'hc23e6cc2, 32'h41b48c87, 32'h42a93bad, 32'hc27d57f3};
test_output[38296:38303] = '{32'h42679e1d, 32'h0, 32'h40c0d114, 32'h0, 32'h0, 32'h41b48c87, 32'h42a93bad, 32'h0};
test_input[38304:38311] = '{32'hc1beb467, 32'hc14a828b, 32'hc2bc8f60, 32'h42c46d7e, 32'hc2c2729c, 32'h4132c54c, 32'h421a146c, 32'h40ba4e76};
test_output[38304:38311] = '{32'h0, 32'h0, 32'h0, 32'h42c46d7e, 32'h0, 32'h4132c54c, 32'h421a146c, 32'h40ba4e76};
test_input[38312:38319] = '{32'h42650150, 32'h42923604, 32'h41677b1a, 32'h41493833, 32'h41223d38, 32'h42903e1e, 32'h42ad50d0, 32'hbedaed5b};
test_output[38312:38319] = '{32'h42650150, 32'h42923604, 32'h41677b1a, 32'h41493833, 32'h41223d38, 32'h42903e1e, 32'h42ad50d0, 32'h0};
test_input[38320:38327] = '{32'h42014f0c, 32'h4253cb3b, 32'h42664acf, 32'h423854e0, 32'h41d8c65e, 32'hbf70ea5b, 32'h4244cf63, 32'h41e708bd};
test_output[38320:38327] = '{32'h42014f0c, 32'h4253cb3b, 32'h42664acf, 32'h423854e0, 32'h41d8c65e, 32'h0, 32'h4244cf63, 32'h41e708bd};
test_input[38328:38335] = '{32'h428d5cfc, 32'h42158a33, 32'h422c0011, 32'hc28abe11, 32'hc2b4fb5b, 32'h3fd3ac98, 32'hc1d6c823, 32'hc280afab};
test_output[38328:38335] = '{32'h428d5cfc, 32'h42158a33, 32'h422c0011, 32'h0, 32'h0, 32'h3fd3ac98, 32'h0, 32'h0};
test_input[38336:38343] = '{32'h41b899aa, 32'h42b05d3e, 32'hc2536c42, 32'h4291f363, 32'h408437c2, 32'hc25d17b3, 32'h41ee5429, 32'h42216f92};
test_output[38336:38343] = '{32'h41b899aa, 32'h42b05d3e, 32'h0, 32'h4291f363, 32'h408437c2, 32'h0, 32'h41ee5429, 32'h42216f92};
test_input[38344:38351] = '{32'h428c4ccc, 32'hc26f57ab, 32'hc2974f0b, 32'hc2bdfa0e, 32'hc2b28a25, 32'hc2121c93, 32'h426296f1, 32'hc22ecabe};
test_output[38344:38351] = '{32'h428c4ccc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426296f1, 32'h0};
test_input[38352:38359] = '{32'hc2748611, 32'hc2a045d3, 32'hc2ae83d8, 32'hc09bed13, 32'h4209fc1b, 32'hc26ff5e0, 32'hc180fe37, 32'h4237de72};
test_output[38352:38359] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4209fc1b, 32'h0, 32'h0, 32'h4237de72};
test_input[38360:38367] = '{32'hc17f4fe8, 32'hc282ca33, 32'hc2b2a04e, 32'hc2115882, 32'h4197cf8a, 32'hc239c606, 32'h42825ca2, 32'hc29eb20b};
test_output[38360:38367] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h4197cf8a, 32'h0, 32'h42825ca2, 32'h0};
test_input[38368:38375] = '{32'hc1b1a80f, 32'hc2b770b9, 32'h42b5f93e, 32'h4232846e, 32'h4013e5f4, 32'hc28bc643, 32'h42b2dcd7, 32'hc233ecc2};
test_output[38368:38375] = '{32'h0, 32'h0, 32'h42b5f93e, 32'h4232846e, 32'h4013e5f4, 32'h0, 32'h42b2dcd7, 32'h0};
test_input[38376:38383] = '{32'h42b6b280, 32'h42804786, 32'h422b934d, 32'hc28cfc8c, 32'hc2a49a89, 32'h42052550, 32'hc2ba8820, 32'hc296f619};
test_output[38376:38383] = '{32'h42b6b280, 32'h42804786, 32'h422b934d, 32'h0, 32'h0, 32'h42052550, 32'h0, 32'h0};
test_input[38384:38391] = '{32'hc234b966, 32'h425d9a20, 32'hc28b6045, 32'h4036cb79, 32'h4294de81, 32'hc249426a, 32'h42a4c240, 32'h420d7ff0};
test_output[38384:38391] = '{32'h0, 32'h425d9a20, 32'h0, 32'h4036cb79, 32'h4294de81, 32'h0, 32'h42a4c240, 32'h420d7ff0};
test_input[38392:38399] = '{32'hc2bd6070, 32'h42864979, 32'hc219054b, 32'hc2aafd21, 32'hc2202354, 32'hc2389f0b, 32'h40a87569, 32'hc268e1ad};
test_output[38392:38399] = '{32'h0, 32'h42864979, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40a87569, 32'h0};
test_input[38400:38407] = '{32'hc22bbffe, 32'h42c32869, 32'h42611d8a, 32'hc297e32a, 32'h4297c235, 32'hc28c2136, 32'hc1ce7b01, 32'h42be7d25};
test_output[38400:38407] = '{32'h0, 32'h42c32869, 32'h42611d8a, 32'h0, 32'h4297c235, 32'h0, 32'h0, 32'h42be7d25};
test_input[38408:38415] = '{32'hc2a40b51, 32'h40f19dca, 32'hc25b873a, 32'h424b3be6, 32'hc27bf36b, 32'h42b866b7, 32'h419ecb08, 32'h428521d1};
test_output[38408:38415] = '{32'h0, 32'h40f19dca, 32'h0, 32'h424b3be6, 32'h0, 32'h42b866b7, 32'h419ecb08, 32'h428521d1};
test_input[38416:38423] = '{32'h415e2204, 32'h428d8d5a, 32'h42353239, 32'h420e1c6f, 32'hc0fc20ad, 32'h41e0c419, 32'h423dfc4d, 32'h420a2b10};
test_output[38416:38423] = '{32'h415e2204, 32'h428d8d5a, 32'h42353239, 32'h420e1c6f, 32'h0, 32'h41e0c419, 32'h423dfc4d, 32'h420a2b10};
test_input[38424:38431] = '{32'hc26961f6, 32'hc14fe8ac, 32'h42b31d1a, 32'hc2824591, 32'h418634e9, 32'h42a7df06, 32'h4167eedc, 32'h42ad8a39};
test_output[38424:38431] = '{32'h0, 32'h0, 32'h42b31d1a, 32'h0, 32'h418634e9, 32'h42a7df06, 32'h4167eedc, 32'h42ad8a39};
test_input[38432:38439] = '{32'h40e9f0ea, 32'h42a41b9d, 32'hc217ef02, 32'h42b6d2e2, 32'hc1e3989f, 32'h42bd690b, 32'h42075558, 32'h425d6b5d};
test_output[38432:38439] = '{32'h40e9f0ea, 32'h42a41b9d, 32'h0, 32'h42b6d2e2, 32'h0, 32'h42bd690b, 32'h42075558, 32'h425d6b5d};
test_input[38440:38447] = '{32'h41d92b78, 32'hc2b10021, 32'h42434f76, 32'hc269fd96, 32'hc2c71587, 32'h428c08f5, 32'h4137683f, 32'hc04fcd41};
test_output[38440:38447] = '{32'h41d92b78, 32'h0, 32'h42434f76, 32'h0, 32'h0, 32'h428c08f5, 32'h4137683f, 32'h0};
test_input[38448:38455] = '{32'hc1e027fc, 32'hc2b4b17e, 32'hc2087a96, 32'h4027389d, 32'h41b4c747, 32'h426b9ca2, 32'hc2a84904, 32'h41a5c68a};
test_output[38448:38455] = '{32'h0, 32'h0, 32'h0, 32'h4027389d, 32'h41b4c747, 32'h426b9ca2, 32'h0, 32'h41a5c68a};
test_input[38456:38463] = '{32'hc26c94b1, 32'hc28249ab, 32'h41deb432, 32'hc2bed599, 32'h41fa68cc, 32'hc1c61a8c, 32'h42783732, 32'hc2021862};
test_output[38456:38463] = '{32'h0, 32'h0, 32'h41deb432, 32'h0, 32'h41fa68cc, 32'h0, 32'h42783732, 32'h0};
test_input[38464:38471] = '{32'h40f5e72b, 32'hc2a922b2, 32'hc2724447, 32'h420d129a, 32'hc19947be, 32'h42877be7, 32'h422b7a22, 32'hc1cf2d1d};
test_output[38464:38471] = '{32'h40f5e72b, 32'h0, 32'h0, 32'h420d129a, 32'h0, 32'h42877be7, 32'h422b7a22, 32'h0};
test_input[38472:38479] = '{32'h41f56d31, 32'hc2a6510e, 32'h41e59f04, 32'hc2818c0a, 32'h402d5d34, 32'hc2c7e6e1, 32'h422fffd4, 32'hc208b16b};
test_output[38472:38479] = '{32'h41f56d31, 32'h0, 32'h41e59f04, 32'h0, 32'h402d5d34, 32'h0, 32'h422fffd4, 32'h0};
test_input[38480:38487] = '{32'hc2970632, 32'h42b0249f, 32'hc2740c6e, 32'hc1c44965, 32'h41ec680e, 32'h42874374, 32'h42a5ee02, 32'h429d0c0a};
test_output[38480:38487] = '{32'h0, 32'h42b0249f, 32'h0, 32'h0, 32'h41ec680e, 32'h42874374, 32'h42a5ee02, 32'h429d0c0a};
test_input[38488:38495] = '{32'hc17a3c08, 32'h4111910d, 32'hc25faa8c, 32'hc29c711a, 32'hc265ead4, 32'hc294bcf0, 32'h42aef991, 32'hc101e661};
test_output[38488:38495] = '{32'h0, 32'h4111910d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42aef991, 32'h0};
test_input[38496:38503] = '{32'hc06642b6, 32'h41a410e4, 32'h41eb7b7c, 32'h405d7140, 32'h41edd0a6, 32'hc2559478, 32'h420ad350, 32'hc28a452a};
test_output[38496:38503] = '{32'h0, 32'h41a410e4, 32'h41eb7b7c, 32'h405d7140, 32'h41edd0a6, 32'h0, 32'h420ad350, 32'h0};
test_input[38504:38511] = '{32'hc29bc0c1, 32'hc1f40c9d, 32'h41dad097, 32'hc114e569, 32'hc1611066, 32'hc28fb19d, 32'h42a67c69, 32'h42ba30ef};
test_output[38504:38511] = '{32'h0, 32'h0, 32'h41dad097, 32'h0, 32'h0, 32'h0, 32'h42a67c69, 32'h42ba30ef};
test_input[38512:38519] = '{32'hc2535012, 32'hc2c5f034, 32'h409e7898, 32'hc2c4c98d, 32'h4229613c, 32'hc2a1d58d, 32'h42a84224, 32'h42bcf7ab};
test_output[38512:38519] = '{32'h0, 32'h0, 32'h409e7898, 32'h0, 32'h4229613c, 32'h0, 32'h42a84224, 32'h42bcf7ab};
test_input[38520:38527] = '{32'hc2929b2e, 32'hc27b6066, 32'hc2852683, 32'hc081b660, 32'h429de7c1, 32'hc255208d, 32'h4264573c, 32'hc23bf699};
test_output[38520:38527] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h429de7c1, 32'h0, 32'h4264573c, 32'h0};
test_input[38528:38535] = '{32'h41853f53, 32'h429c492a, 32'h428f5e03, 32'h4098dcb9, 32'h415d0492, 32'hc2b3b0e3, 32'h42c2876c, 32'hc1f9806e};
test_output[38528:38535] = '{32'h41853f53, 32'h429c492a, 32'h428f5e03, 32'h4098dcb9, 32'h415d0492, 32'h0, 32'h42c2876c, 32'h0};
test_input[38536:38543] = '{32'h42585d48, 32'h4137de3c, 32'h426f8e3a, 32'h41e976d0, 32'hc2861666, 32'h41add3a1, 32'h4271d3f2, 32'hc2a5efc7};
test_output[38536:38543] = '{32'h42585d48, 32'h4137de3c, 32'h426f8e3a, 32'h41e976d0, 32'h0, 32'h41add3a1, 32'h4271d3f2, 32'h0};
test_input[38544:38551] = '{32'hc1ae4f9f, 32'h420cc44c, 32'hc2c70d8c, 32'hc0a76536, 32'hc1f45207, 32'hc2886e5c, 32'h40fa333c, 32'hc1c120f9};
test_output[38544:38551] = '{32'h0, 32'h420cc44c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40fa333c, 32'h0};
test_input[38552:38559] = '{32'hc23d712b, 32'h42ac1e19, 32'hc257a97e, 32'h42b23d89, 32'h42a1170b, 32'h42c51eac, 32'hc069e5fd, 32'hc2a2629a};
test_output[38552:38559] = '{32'h0, 32'h42ac1e19, 32'h0, 32'h42b23d89, 32'h42a1170b, 32'h42c51eac, 32'h0, 32'h0};
test_input[38560:38567] = '{32'hc2a5cebb, 32'h42b62094, 32'hc2b559ac, 32'h424d9846, 32'hc236819a, 32'h4253a08e, 32'h4296687b, 32'h426d511c};
test_output[38560:38567] = '{32'h0, 32'h42b62094, 32'h0, 32'h424d9846, 32'h0, 32'h4253a08e, 32'h4296687b, 32'h426d511c};
test_input[38568:38575] = '{32'h40acd67c, 32'h42b66c5f, 32'h42c25842, 32'hc27819c0, 32'h41fa638a, 32'h42172a47, 32'hc2871429, 32'hc087e319};
test_output[38568:38575] = '{32'h40acd67c, 32'h42b66c5f, 32'h42c25842, 32'h0, 32'h41fa638a, 32'h42172a47, 32'h0, 32'h0};
test_input[38576:38583] = '{32'h4149fb8f, 32'hc2512964, 32'h42bd8360, 32'h422e8b96, 32'hc257b62d, 32'h42a3cad3, 32'hc2b2a408, 32'h40c5ce81};
test_output[38576:38583] = '{32'h4149fb8f, 32'h0, 32'h42bd8360, 32'h422e8b96, 32'h0, 32'h42a3cad3, 32'h0, 32'h40c5ce81};
test_input[38584:38591] = '{32'hc11e85ee, 32'h4234f75f, 32'h41b6f4e5, 32'h3f766f63, 32'hc2a3e993, 32'hbfaaaf2e, 32'h4176368f, 32'h41641540};
test_output[38584:38591] = '{32'h0, 32'h4234f75f, 32'h41b6f4e5, 32'h3f766f63, 32'h0, 32'h0, 32'h4176368f, 32'h41641540};
test_input[38592:38599] = '{32'hc1ebe5d4, 32'h424dc81d, 32'h42aa6a24, 32'h41efb45b, 32'h424a0a02, 32'h428d3b4b, 32'h4020f321, 32'hc19f2eb9};
test_output[38592:38599] = '{32'h0, 32'h424dc81d, 32'h42aa6a24, 32'h41efb45b, 32'h424a0a02, 32'h428d3b4b, 32'h4020f321, 32'h0};
test_input[38600:38607] = '{32'hc20bb033, 32'hc1ed5849, 32'h423cc61c, 32'h42acc9e5, 32'hc2b5de1a, 32'hc24fb800, 32'hc281ec07, 32'h4237373e};
test_output[38600:38607] = '{32'h0, 32'h0, 32'h423cc61c, 32'h42acc9e5, 32'h0, 32'h0, 32'h0, 32'h4237373e};
test_input[38608:38615] = '{32'hc2661f32, 32'hc2118abe, 32'hc200ac33, 32'hc2a53076, 32'hc29fa3c4, 32'h42b9fa38, 32'hc2995895, 32'hc243c9ba};
test_output[38608:38615] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b9fa38, 32'h0, 32'h0};
test_input[38616:38623] = '{32'hc205da74, 32'hc1fe94db, 32'h42b4497b, 32'h42b20ac2, 32'hc2ad7ca9, 32'h42c6d194, 32'h428fa05e, 32'h420cea3d};
test_output[38616:38623] = '{32'h0, 32'h0, 32'h42b4497b, 32'h42b20ac2, 32'h0, 32'h42c6d194, 32'h428fa05e, 32'h420cea3d};
test_input[38624:38631] = '{32'h42472619, 32'hc150219e, 32'hc25ff979, 32'h4223cac7, 32'h42664deb, 32'h41b5e63c, 32'hc28bd5b9, 32'hc252c33d};
test_output[38624:38631] = '{32'h42472619, 32'h0, 32'h0, 32'h4223cac7, 32'h42664deb, 32'h41b5e63c, 32'h0, 32'h0};
test_input[38632:38639] = '{32'hc2bd6ea8, 32'h419ee0a8, 32'h41c37aa0, 32'hc1a2be96, 32'hc0b13355, 32'hc281835a, 32'h424cd9c4, 32'hc2870272};
test_output[38632:38639] = '{32'h0, 32'h419ee0a8, 32'h41c37aa0, 32'h0, 32'h0, 32'h0, 32'h424cd9c4, 32'h0};
test_input[38640:38647] = '{32'h418e230c, 32'hc2bca83f, 32'hc2807731, 32'h42a2499d, 32'hc1a4df42, 32'hc28d2b04, 32'hc2c3d736, 32'h429b4543};
test_output[38640:38647] = '{32'h418e230c, 32'h0, 32'h0, 32'h42a2499d, 32'h0, 32'h0, 32'h0, 32'h429b4543};
test_input[38648:38655] = '{32'hc2c59b0b, 32'h41f2cc10, 32'h42561c17, 32'hc295abdd, 32'h4029f9af, 32'hc2b10238, 32'hc13b1db4, 32'h4191318a};
test_output[38648:38655] = '{32'h0, 32'h41f2cc10, 32'h42561c17, 32'h0, 32'h4029f9af, 32'h0, 32'h0, 32'h4191318a};
test_input[38656:38663] = '{32'hc25b7e29, 32'h42b94a2b, 32'h4218ab39, 32'hc18a5f1b, 32'hc13727b0, 32'h3fd36cba, 32'hc2c6d780, 32'hc2aec4cd};
test_output[38656:38663] = '{32'h0, 32'h42b94a2b, 32'h4218ab39, 32'h0, 32'h0, 32'h3fd36cba, 32'h0, 32'h0};
test_input[38664:38671] = '{32'h41f3c866, 32'hc2c45004, 32'hc2bbd7f7, 32'hc2c05740, 32'h42b89e0d, 32'h4214e841, 32'h42b164fb, 32'h4237d991};
test_output[38664:38671] = '{32'h41f3c866, 32'h0, 32'h0, 32'h0, 32'h42b89e0d, 32'h4214e841, 32'h42b164fb, 32'h4237d991};
test_input[38672:38679] = '{32'h42716277, 32'h425b250d, 32'hc165d52f, 32'h429dd309, 32'hc19d105c, 32'h42b96561, 32'hc0e5149b, 32'h4241382d};
test_output[38672:38679] = '{32'h42716277, 32'h425b250d, 32'h0, 32'h429dd309, 32'h0, 32'h42b96561, 32'h0, 32'h4241382d};
test_input[38680:38687] = '{32'hc1af4078, 32'h42a0c6e5, 32'h417f812f, 32'h41d99d9c, 32'hc20e28fb, 32'h429f31cc, 32'hc2755e8f, 32'h3e6d59e6};
test_output[38680:38687] = '{32'h0, 32'h42a0c6e5, 32'h417f812f, 32'h41d99d9c, 32'h0, 32'h429f31cc, 32'h0, 32'h3e6d59e6};
test_input[38688:38695] = '{32'h42301760, 32'h425e4c35, 32'hbf86b9f9, 32'h41e31a74, 32'hc0ceefeb, 32'hc0c6f35a, 32'hc23d0cc3, 32'h426c7e0f};
test_output[38688:38695] = '{32'h42301760, 32'h425e4c35, 32'h0, 32'h41e31a74, 32'h0, 32'h0, 32'h0, 32'h426c7e0f};
test_input[38696:38703] = '{32'h4283e150, 32'hc1fdd965, 32'hc2bf55ed, 32'h42ac02c0, 32'hc1094054, 32'h421559ed, 32'hc200583c, 32'h41fd189f};
test_output[38696:38703] = '{32'h4283e150, 32'h0, 32'h0, 32'h42ac02c0, 32'h0, 32'h421559ed, 32'h0, 32'h41fd189f};
test_input[38704:38711] = '{32'h4266b328, 32'h42a3cdb2, 32'h42a2117d, 32'hc2404e2f, 32'hc206bf5b, 32'hc1be6c1f, 32'hc230375b, 32'h413b526d};
test_output[38704:38711] = '{32'h4266b328, 32'h42a3cdb2, 32'h42a2117d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h413b526d};
test_input[38712:38719] = '{32'h42ada3a0, 32'hc10ec468, 32'hc2441adf, 32'hc1e07334, 32'h41e01e5e, 32'hc191117a, 32'hc27c6e89, 32'h42603e82};
test_output[38712:38719] = '{32'h42ada3a0, 32'h0, 32'h0, 32'h0, 32'h41e01e5e, 32'h0, 32'h0, 32'h42603e82};
test_input[38720:38727] = '{32'hc287cfc1, 32'h428e2a8b, 32'hc2aef2ba, 32'h42a9027d, 32'hc28c00af, 32'hc12b0f11, 32'h4121295c, 32'h41c85903};
test_output[38720:38727] = '{32'h0, 32'h428e2a8b, 32'h0, 32'h42a9027d, 32'h0, 32'h0, 32'h4121295c, 32'h41c85903};
test_input[38728:38735] = '{32'hc220dbe0, 32'hc299e92e, 32'h40a82604, 32'h429b4ba5, 32'h429e4af3, 32'h42bd6d8f, 32'hc2a81b14, 32'hc2a7eaaa};
test_output[38728:38735] = '{32'h0, 32'h0, 32'h40a82604, 32'h429b4ba5, 32'h429e4af3, 32'h42bd6d8f, 32'h0, 32'h0};
test_input[38736:38743] = '{32'h427c11f2, 32'h429df91b, 32'hc210248e, 32'hc2af3c17, 32'h41abedb1, 32'hc1d8f9d8, 32'h405ccd30, 32'hc28f44c2};
test_output[38736:38743] = '{32'h427c11f2, 32'h429df91b, 32'h0, 32'h0, 32'h41abedb1, 32'h0, 32'h405ccd30, 32'h0};
test_input[38744:38751] = '{32'hc25183ce, 32'hc2ae8e79, 32'hc1f73a11, 32'h4193406f, 32'h41996f99, 32'hc0ad4404, 32'hc2b708f2, 32'h411eddd9};
test_output[38744:38751] = '{32'h0, 32'h0, 32'h0, 32'h4193406f, 32'h41996f99, 32'h0, 32'h0, 32'h411eddd9};
test_input[38752:38759] = '{32'h41dfb929, 32'hc1a35bd3, 32'h41811b00, 32'h42bf5f8a, 32'h425a7d4e, 32'h42419339, 32'h4182c0fb, 32'hc1821bb2};
test_output[38752:38759] = '{32'h41dfb929, 32'h0, 32'h41811b00, 32'h42bf5f8a, 32'h425a7d4e, 32'h42419339, 32'h4182c0fb, 32'h0};
test_input[38760:38767] = '{32'hc2ae80de, 32'hc1efaeb2, 32'hc288f36c, 32'h40b9e6e1, 32'hc219a0d1, 32'h401b4fdf, 32'hc21b48ea, 32'h42574c09};
test_output[38760:38767] = '{32'h0, 32'h0, 32'h0, 32'h40b9e6e1, 32'h0, 32'h401b4fdf, 32'h0, 32'h42574c09};
test_input[38768:38775] = '{32'hbfa0d786, 32'h41b8d830, 32'h405aa5bc, 32'hc2c09532, 32'h41de910d, 32'hc1e927d2, 32'h42a15d76, 32'hc2552ed1};
test_output[38768:38775] = '{32'h0, 32'h41b8d830, 32'h405aa5bc, 32'h0, 32'h41de910d, 32'h0, 32'h42a15d76, 32'h0};
test_input[38776:38783] = '{32'h42be4cbb, 32'h42c27957, 32'h42911c2a, 32'h42846651, 32'hc2b06cd5, 32'hc22f1686, 32'hc2139ba6, 32'h42873910};
test_output[38776:38783] = '{32'h42be4cbb, 32'h42c27957, 32'h42911c2a, 32'h42846651, 32'h0, 32'h0, 32'h0, 32'h42873910};
test_input[38784:38791] = '{32'hc03aad0b, 32'h42c56420, 32'hc2c44e45, 32'hc2c10ee5, 32'hc2bccf2e, 32'hc1516186, 32'h4195bffb, 32'hc1dc559f};
test_output[38784:38791] = '{32'h0, 32'h42c56420, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4195bffb, 32'h0};
test_input[38792:38799] = '{32'h429260c7, 32'hc28aef7c, 32'h42c4ba68, 32'h41b3a285, 32'h426cd310, 32'hc215c0d4, 32'hc2a57075, 32'h41ef5f8d};
test_output[38792:38799] = '{32'h429260c7, 32'h0, 32'h42c4ba68, 32'h41b3a285, 32'h426cd310, 32'h0, 32'h0, 32'h41ef5f8d};
test_input[38800:38807] = '{32'h4232c231, 32'h424679cd, 32'hc10aa9ee, 32'h424a632b, 32'hc1b60eb3, 32'hc1ac2bc5, 32'hc2c35719, 32'h419f158f};
test_output[38800:38807] = '{32'h4232c231, 32'h424679cd, 32'h0, 32'h424a632b, 32'h0, 32'h0, 32'h0, 32'h419f158f};
test_input[38808:38815] = '{32'h41e6bed8, 32'h42568182, 32'hc284c48d, 32'hc2c0e2b2, 32'hc2a7d6d9, 32'h4244cff9, 32'hc173d142, 32'h42bc10a3};
test_output[38808:38815] = '{32'h41e6bed8, 32'h42568182, 32'h0, 32'h0, 32'h0, 32'h4244cff9, 32'h0, 32'h42bc10a3};
test_input[38816:38823] = '{32'hc2699850, 32'hc2c69a75, 32'h4191f65a, 32'h42996899, 32'h407b617d, 32'hc2c44743, 32'h41e8847a, 32'h411c5c5d};
test_output[38816:38823] = '{32'h0, 32'h0, 32'h4191f65a, 32'h42996899, 32'h407b617d, 32'h0, 32'h41e8847a, 32'h411c5c5d};
test_input[38824:38831] = '{32'h41afb8ec, 32'hc29600db, 32'h41547c1d, 32'hc19f88e4, 32'h41d3ddb9, 32'h4236d2a3, 32'h4215ef3e, 32'hc1540841};
test_output[38824:38831] = '{32'h41afb8ec, 32'h0, 32'h41547c1d, 32'h0, 32'h41d3ddb9, 32'h4236d2a3, 32'h4215ef3e, 32'h0};
test_input[38832:38839] = '{32'h42815bd8, 32'hc2640d98, 32'h42897a13, 32'hc2974bde, 32'hc23852d3, 32'h428118c2, 32'hc28969ef, 32'h42a69217};
test_output[38832:38839] = '{32'h42815bd8, 32'h0, 32'h42897a13, 32'h0, 32'h0, 32'h428118c2, 32'h0, 32'h42a69217};
test_input[38840:38847] = '{32'h42c564ce, 32'h4286013e, 32'hc20d0264, 32'h42996a60, 32'hc1abcf15, 32'hc2a93d5a, 32'h410754c0, 32'hc26c5809};
test_output[38840:38847] = '{32'h42c564ce, 32'h4286013e, 32'h0, 32'h42996a60, 32'h0, 32'h0, 32'h410754c0, 32'h0};
test_input[38848:38855] = '{32'h400df0a8, 32'h40141e3d, 32'hc1d3f03f, 32'hc142277a, 32'h41d6a0df, 32'hc2a5ca0a, 32'h42c352aa, 32'h4293800f};
test_output[38848:38855] = '{32'h400df0a8, 32'h40141e3d, 32'h0, 32'h0, 32'h41d6a0df, 32'h0, 32'h42c352aa, 32'h4293800f};
test_input[38856:38863] = '{32'h4210952a, 32'h42a513a3, 32'h4260bf5b, 32'hc28d3b26, 32'hc2a592da, 32'h42be03fa, 32'h42b8da84, 32'h423b038f};
test_output[38856:38863] = '{32'h4210952a, 32'h42a513a3, 32'h4260bf5b, 32'h0, 32'h0, 32'h42be03fa, 32'h42b8da84, 32'h423b038f};
test_input[38864:38871] = '{32'hc2369b41, 32'h42a638e0, 32'h42888383, 32'h42c0a126, 32'hc10c239a, 32'hc1b282a7, 32'h4148dd6c, 32'hc0b52f0f};
test_output[38864:38871] = '{32'h0, 32'h42a638e0, 32'h42888383, 32'h42c0a126, 32'h0, 32'h0, 32'h4148dd6c, 32'h0};
test_input[38872:38879] = '{32'hc298ddde, 32'h425e2949, 32'hc2bbbd78, 32'h42c16e35, 32'h41c93557, 32'hc20a3e5d, 32'h429575da, 32'h41b070fe};
test_output[38872:38879] = '{32'h0, 32'h425e2949, 32'h0, 32'h42c16e35, 32'h41c93557, 32'h0, 32'h429575da, 32'h41b070fe};
test_input[38880:38887] = '{32'hc1a564c4, 32'h40708dfb, 32'hc28cd01f, 32'hc030c768, 32'hc250ccfa, 32'h42aca455, 32'h42bbaacf, 32'hc29d4357};
test_output[38880:38887] = '{32'h0, 32'h40708dfb, 32'h0, 32'h0, 32'h0, 32'h42aca455, 32'h42bbaacf, 32'h0};
test_input[38888:38895] = '{32'h42695ab7, 32'h42259b28, 32'hc2b6e97a, 32'hc1fb0453, 32'h42600c23, 32'h422c2d57, 32'h42aebc32, 32'h42a00cfa};
test_output[38888:38895] = '{32'h42695ab7, 32'h42259b28, 32'h0, 32'h0, 32'h42600c23, 32'h422c2d57, 32'h42aebc32, 32'h42a00cfa};
test_input[38896:38903] = '{32'h4277446d, 32'hc21e8f7d, 32'h420e7b02, 32'h4273bdd3, 32'h422e164f, 32'hc20121c5, 32'hc28f386e, 32'h42bf527f};
test_output[38896:38903] = '{32'h4277446d, 32'h0, 32'h420e7b02, 32'h4273bdd3, 32'h422e164f, 32'h0, 32'h0, 32'h42bf527f};
test_input[38904:38911] = '{32'h42b63d95, 32'h426639db, 32'hc0841b52, 32'h42b73328, 32'h4120be67, 32'hc2156501, 32'h42b7d9ec, 32'h416a5b7a};
test_output[38904:38911] = '{32'h42b63d95, 32'h426639db, 32'h0, 32'h42b73328, 32'h4120be67, 32'h0, 32'h42b7d9ec, 32'h416a5b7a};
test_input[38912:38919] = '{32'h42c1c1f6, 32'h41bfd27f, 32'h421eb4f9, 32'h40cd5c19, 32'h426b180e, 32'h42c7ebe0, 32'h40a53e9a, 32'hc22a4624};
test_output[38912:38919] = '{32'h42c1c1f6, 32'h41bfd27f, 32'h421eb4f9, 32'h40cd5c19, 32'h426b180e, 32'h42c7ebe0, 32'h40a53e9a, 32'h0};
test_input[38920:38927] = '{32'h404bd612, 32'h42529458, 32'h41542a46, 32'h422a7311, 32'hc2b1cfc9, 32'h422e2aa1, 32'h42817ca3, 32'hc20e9fc8};
test_output[38920:38927] = '{32'h404bd612, 32'h42529458, 32'h41542a46, 32'h422a7311, 32'h0, 32'h422e2aa1, 32'h42817ca3, 32'h0};
test_input[38928:38935] = '{32'hc2b96dd3, 32'hc251d745, 32'h422b0357, 32'hc281f724, 32'h42ad9726, 32'hc189b273, 32'hc284ba4f, 32'hc26e325a};
test_output[38928:38935] = '{32'h0, 32'h0, 32'h422b0357, 32'h0, 32'h42ad9726, 32'h0, 32'h0, 32'h0};
test_input[38936:38943] = '{32'hc1d25b01, 32'h42048da1, 32'hc29ed8aa, 32'hc18dfc45, 32'h42368ed1, 32'h428b9895, 32'hc22efe71, 32'h4270fa0f};
test_output[38936:38943] = '{32'h0, 32'h42048da1, 32'h0, 32'h0, 32'h42368ed1, 32'h428b9895, 32'h0, 32'h4270fa0f};
test_input[38944:38951] = '{32'h41dd91b8, 32'hc1a702dc, 32'hc2baafcc, 32'hc0d8e62a, 32'hc230424f, 32'hbf58f527, 32'h421616cf, 32'hc1fa991b};
test_output[38944:38951] = '{32'h41dd91b8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h421616cf, 32'h0};
test_input[38952:38959] = '{32'h41b203f7, 32'h4201a136, 32'h42b3aa13, 32'hc289fb62, 32'hc207e360, 32'hc2be8118, 32'h42232a84, 32'h428f1e81};
test_output[38952:38959] = '{32'h41b203f7, 32'h4201a136, 32'h42b3aa13, 32'h0, 32'h0, 32'h0, 32'h42232a84, 32'h428f1e81};
test_input[38960:38967] = '{32'hc11f928a, 32'h41fdeae1, 32'hc296403c, 32'hc273445a, 32'hc2847144, 32'h41394dd7, 32'h421bb536, 32'h4246e0b3};
test_output[38960:38967] = '{32'h0, 32'h41fdeae1, 32'h0, 32'h0, 32'h0, 32'h41394dd7, 32'h421bb536, 32'h4246e0b3};
test_input[38968:38975] = '{32'hc2be6a9a, 32'hc1875e91, 32'hc21822d1, 32'hc2a409a4, 32'h41e08a0c, 32'h420da1ce, 32'h421b925e, 32'h4252aeaf};
test_output[38968:38975] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41e08a0c, 32'h420da1ce, 32'h421b925e, 32'h4252aeaf};
test_input[38976:38983] = '{32'hc22c10cc, 32'hc21caf75, 32'hc1cb8610, 32'hc24925cf, 32'h41852b7c, 32'hc2a478a5, 32'h41e6734d, 32'h42a7382e};
test_output[38976:38983] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41852b7c, 32'h0, 32'h41e6734d, 32'h42a7382e};
test_input[38984:38991] = '{32'h42b84a72, 32'h4110dd4b, 32'hc29aa81a, 32'h3f0f54a3, 32'h4091f10f, 32'h42606248, 32'h42b67cb5, 32'h40534278};
test_output[38984:38991] = '{32'h42b84a72, 32'h4110dd4b, 32'h0, 32'h3f0f54a3, 32'h4091f10f, 32'h42606248, 32'h42b67cb5, 32'h40534278};
test_input[38992:38999] = '{32'h421a4678, 32'hc23cf8bb, 32'hc1c98b29, 32'h424e8ef3, 32'h40be8479, 32'h42372635, 32'hc1a0453a, 32'hc1a184c2};
test_output[38992:38999] = '{32'h421a4678, 32'h0, 32'h0, 32'h424e8ef3, 32'h40be8479, 32'h42372635, 32'h0, 32'h0};
test_input[39000:39007] = '{32'h423bdf7a, 32'h41b7d55f, 32'h428bc106, 32'hc28fd5df, 32'h4248feed, 32'hc238589a, 32'h41c29fe0, 32'hc213ebab};
test_output[39000:39007] = '{32'h423bdf7a, 32'h41b7d55f, 32'h428bc106, 32'h0, 32'h4248feed, 32'h0, 32'h41c29fe0, 32'h0};
test_input[39008:39015] = '{32'h4297a9d5, 32'hc176971d, 32'hc26279b3, 32'hc25cee85, 32'hc21e25ec, 32'hc293d3b3, 32'h42b778dc, 32'h42a0059d};
test_output[39008:39015] = '{32'h4297a9d5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42b778dc, 32'h42a0059d};
test_input[39016:39023] = '{32'h4264d2d8, 32'hc284ff16, 32'hc19e6552, 32'h42b5d111, 32'hc28ea1bf, 32'hc20b13cb, 32'h4285824d, 32'h429f7c84};
test_output[39016:39023] = '{32'h4264d2d8, 32'h0, 32'h0, 32'h42b5d111, 32'h0, 32'h0, 32'h4285824d, 32'h429f7c84};
test_input[39024:39031] = '{32'h426d50fd, 32'hc23438c0, 32'hc2a8b7f5, 32'h41a146f6, 32'h421cd293, 32'h41ce5106, 32'hc1b588d0, 32'h4191033b};
test_output[39024:39031] = '{32'h426d50fd, 32'h0, 32'h0, 32'h41a146f6, 32'h421cd293, 32'h41ce5106, 32'h0, 32'h4191033b};
test_input[39032:39039] = '{32'h429784c0, 32'hc1d310ed, 32'h42c0be77, 32'hc28a4eaa, 32'h428bb549, 32'hc1d39273, 32'h42ba222d, 32'h4170232d};
test_output[39032:39039] = '{32'h429784c0, 32'h0, 32'h42c0be77, 32'h0, 32'h428bb549, 32'h0, 32'h42ba222d, 32'h4170232d};
test_input[39040:39047] = '{32'hc2ba37c1, 32'hc2a1aa72, 32'hc2a2fae3, 32'h416106ae, 32'h41ecb1ad, 32'hc1dc7986, 32'h41a820f8, 32'h41cd4b60};
test_output[39040:39047] = '{32'h0, 32'h0, 32'h0, 32'h416106ae, 32'h41ecb1ad, 32'h0, 32'h41a820f8, 32'h41cd4b60};
test_input[39048:39055] = '{32'h419f9b1c, 32'h427fff3f, 32'h42a2e1d0, 32'h40efd353, 32'hc25340d4, 32'h41217482, 32'hc25934a3, 32'h4240dd66};
test_output[39048:39055] = '{32'h419f9b1c, 32'h427fff3f, 32'h42a2e1d0, 32'h40efd353, 32'h0, 32'h41217482, 32'h0, 32'h4240dd66};
test_input[39056:39063] = '{32'h42aec007, 32'h42a3aa1a, 32'h427016b4, 32'hc29671b3, 32'hc0e27aba, 32'h42587d23, 32'h4209ab30, 32'h418d12b3};
test_output[39056:39063] = '{32'h42aec007, 32'h42a3aa1a, 32'h427016b4, 32'h0, 32'h0, 32'h42587d23, 32'h4209ab30, 32'h418d12b3};
test_input[39064:39071] = '{32'hc2ba833f, 32'h423e2b30, 32'hc2762ab7, 32'h42aa382c, 32'hc2935fbd, 32'hc29a001a, 32'h42674d8e, 32'hc264077a};
test_output[39064:39071] = '{32'h0, 32'h423e2b30, 32'h0, 32'h42aa382c, 32'h0, 32'h0, 32'h42674d8e, 32'h0};
test_input[39072:39079] = '{32'h41a2656e, 32'hc2494c82, 32'h42b4c908, 32'hc20e96b3, 32'hc1a06bc4, 32'h41850fdb, 32'h42c26624, 32'h41e91a6a};
test_output[39072:39079] = '{32'h41a2656e, 32'h0, 32'h42b4c908, 32'h0, 32'h0, 32'h41850fdb, 32'h42c26624, 32'h41e91a6a};
test_input[39080:39087] = '{32'hc232466e, 32'hc29ed49c, 32'h42abbbd0, 32'hc24c62f1, 32'h426412f8, 32'h42a0c303, 32'hc298b55b, 32'h4209d190};
test_output[39080:39087] = '{32'h0, 32'h0, 32'h42abbbd0, 32'h0, 32'h426412f8, 32'h42a0c303, 32'h0, 32'h4209d190};
test_input[39088:39095] = '{32'hc257a73e, 32'hc2577393, 32'h41106ca5, 32'hc295f763, 32'h41e1b630, 32'hc11da2d0, 32'hc288d600, 32'hc1e887bd};
test_output[39088:39095] = '{32'h0, 32'h0, 32'h41106ca5, 32'h0, 32'h41e1b630, 32'h0, 32'h0, 32'h0};
test_input[39096:39103] = '{32'h42244e77, 32'hc29c575c, 32'hc2528f72, 32'hc109e211, 32'hbfb617c0, 32'h423c8af7, 32'hc28ba89d, 32'hc26706ad};
test_output[39096:39103] = '{32'h42244e77, 32'h0, 32'h0, 32'h0, 32'h0, 32'h423c8af7, 32'h0, 32'h0};
test_input[39104:39111] = '{32'h42b6251b, 32'h42b2c59a, 32'h41e55be6, 32'h4287267f, 32'hc22929b4, 32'h4280e78a, 32'h4281a3c2, 32'hc25e74de};
test_output[39104:39111] = '{32'h42b6251b, 32'h42b2c59a, 32'h41e55be6, 32'h4287267f, 32'h0, 32'h4280e78a, 32'h4281a3c2, 32'h0};
test_input[39112:39119] = '{32'h4181bd6c, 32'h4252eedf, 32'h4129ba43, 32'hc28e273a, 32'h41890ff2, 32'hc28a98c8, 32'hc251e42a, 32'hc21189b3};
test_output[39112:39119] = '{32'h4181bd6c, 32'h4252eedf, 32'h4129ba43, 32'h0, 32'h41890ff2, 32'h0, 32'h0, 32'h0};
test_input[39120:39127] = '{32'hc2042551, 32'h4242393a, 32'hc251eb2f, 32'h423594a2, 32'hc2bacb5a, 32'hc19b9714, 32'h4156f6d2, 32'h4106f2b4};
test_output[39120:39127] = '{32'h0, 32'h4242393a, 32'h0, 32'h423594a2, 32'h0, 32'h0, 32'h4156f6d2, 32'h4106f2b4};
test_input[39128:39135] = '{32'hc116dafd, 32'h424d390e, 32'h418790e1, 32'h4216ba92, 32'h42359fa6, 32'hc1a519ed, 32'h42b9d64d, 32'hc0089689};
test_output[39128:39135] = '{32'h0, 32'h424d390e, 32'h418790e1, 32'h4216ba92, 32'h42359fa6, 32'h0, 32'h42b9d64d, 32'h0};
test_input[39136:39143] = '{32'hc25d5366, 32'h4265aad0, 32'h429d33fb, 32'hc1eaa58e, 32'h41ba7070, 32'h42919035, 32'hc1b15e2e, 32'hc2a54426};
test_output[39136:39143] = '{32'h0, 32'h4265aad0, 32'h429d33fb, 32'h0, 32'h41ba7070, 32'h42919035, 32'h0, 32'h0};
test_input[39144:39151] = '{32'h42c13943, 32'hc2a5c75d, 32'h41ade05b, 32'h418e7dd9, 32'hc2b01ae8, 32'h41f6c254, 32'hc28c05ff, 32'hc0af46b8};
test_output[39144:39151] = '{32'h42c13943, 32'h0, 32'h41ade05b, 32'h418e7dd9, 32'h0, 32'h41f6c254, 32'h0, 32'h0};
test_input[39152:39159] = '{32'h42bf63c4, 32'h41a4f265, 32'h41f12b8d, 32'hc250a39d, 32'h4291e0d1, 32'h41282d74, 32'h418f2f67, 32'hc2936a30};
test_output[39152:39159] = '{32'h42bf63c4, 32'h41a4f265, 32'h41f12b8d, 32'h0, 32'h4291e0d1, 32'h41282d74, 32'h418f2f67, 32'h0};
test_input[39160:39167] = '{32'h42045da0, 32'hc044f261, 32'h41d5235c, 32'h417b7063, 32'hc2c74a2e, 32'hc2b45172, 32'hc29e33bc, 32'h42adc1f6};
test_output[39160:39167] = '{32'h42045da0, 32'h0, 32'h41d5235c, 32'h417b7063, 32'h0, 32'h0, 32'h0, 32'h42adc1f6};
test_input[39168:39175] = '{32'h4111e6f4, 32'h410bb2de, 32'h4238f356, 32'h413d8164, 32'hc20477e1, 32'h4130deb7, 32'hc2afab42, 32'h41f61714};
test_output[39168:39175] = '{32'h4111e6f4, 32'h410bb2de, 32'h4238f356, 32'h413d8164, 32'h0, 32'h4130deb7, 32'h0, 32'h41f61714};
test_input[39176:39183] = '{32'h4273a1a0, 32'hc2c2377b, 32'hc2905626, 32'hc008fcca, 32'hc2846896, 32'h42bc9486, 32'hc244f541, 32'h41ecd23e};
test_output[39176:39183] = '{32'h4273a1a0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42bc9486, 32'h0, 32'h41ecd23e};
test_input[39184:39191] = '{32'hc2907ead, 32'hc212f516, 32'h4158168a, 32'h429c640a, 32'hc2a5816e, 32'h41b88b8e, 32'h4205f11d, 32'h41c995b4};
test_output[39184:39191] = '{32'h0, 32'h0, 32'h4158168a, 32'h429c640a, 32'h0, 32'h41b88b8e, 32'h4205f11d, 32'h41c995b4};
test_input[39192:39199] = '{32'h42612bc2, 32'hc13e0742, 32'h42b86628, 32'h416b4394, 32'hc19d352f, 32'hc195f6cd, 32'h42bc230f, 32'hc25695c4};
test_output[39192:39199] = '{32'h42612bc2, 32'h0, 32'h42b86628, 32'h416b4394, 32'h0, 32'h0, 32'h42bc230f, 32'h0};
test_input[39200:39207] = '{32'h4282cefa, 32'h409de56b, 32'hc22068c0, 32'h421663fe, 32'h4290ff43, 32'hc1657654, 32'hc28524a2, 32'hc275bdcc};
test_output[39200:39207] = '{32'h4282cefa, 32'h409de56b, 32'h0, 32'h421663fe, 32'h4290ff43, 32'h0, 32'h0, 32'h0};
test_input[39208:39215] = '{32'hc1428e61, 32'hc241de0d, 32'h41115f67, 32'hc2925e55, 32'hc259e960, 32'h42559544, 32'hc286af2d, 32'hc205a939};
test_output[39208:39215] = '{32'h0, 32'h0, 32'h41115f67, 32'h0, 32'h0, 32'h42559544, 32'h0, 32'h0};
test_input[39216:39223] = '{32'hc2013522, 32'hc2bf6c07, 32'h41f61ae9, 32'h41dbfa00, 32'h4259b39f, 32'hc2ae40f9, 32'hc2920f9c, 32'hc2246bb6};
test_output[39216:39223] = '{32'h0, 32'h0, 32'h41f61ae9, 32'h41dbfa00, 32'h4259b39f, 32'h0, 32'h0, 32'h0};
test_input[39224:39231] = '{32'h40f55112, 32'hc01f5c24, 32'hc2808064, 32'hc2c4ca5a, 32'hc24f9acb, 32'h41d5308c, 32'h4286d1e2, 32'h426280c1};
test_output[39224:39231] = '{32'h40f55112, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41d5308c, 32'h4286d1e2, 32'h426280c1};
test_input[39232:39239] = '{32'h4241fcee, 32'h428e33ad, 32'h4282ab7f, 32'hc10cff66, 32'h40354476, 32'hc2a4c451, 32'h429fab53, 32'hc28a54e7};
test_output[39232:39239] = '{32'h4241fcee, 32'h428e33ad, 32'h4282ab7f, 32'h0, 32'h40354476, 32'h0, 32'h429fab53, 32'h0};
test_input[39240:39247] = '{32'h428b3f3f, 32'h42b41083, 32'hc25b7145, 32'hc2563ff4, 32'h42a260fb, 32'h4297a391, 32'hc2c02ba6, 32'h4206b7df};
test_output[39240:39247] = '{32'h428b3f3f, 32'h42b41083, 32'h0, 32'h0, 32'h42a260fb, 32'h4297a391, 32'h0, 32'h4206b7df};
test_input[39248:39255] = '{32'h41e5b3f3, 32'hc17b934d, 32'h422cd008, 32'hc2a52c17, 32'h414533ff, 32'h41cb9298, 32'h41d1b552, 32'hc111486e};
test_output[39248:39255] = '{32'h41e5b3f3, 32'h0, 32'h422cd008, 32'h0, 32'h414533ff, 32'h41cb9298, 32'h41d1b552, 32'h0};
test_input[39256:39263] = '{32'h404376e0, 32'h4234ddce, 32'hc285191d, 32'h428214f0, 32'hc1dc3047, 32'hc2b5bc8b, 32'h42013edb, 32'hc2710479};
test_output[39256:39263] = '{32'h404376e0, 32'h4234ddce, 32'h0, 32'h428214f0, 32'h0, 32'h0, 32'h42013edb, 32'h0};
test_input[39264:39271] = '{32'h42975c05, 32'h40218aff, 32'hc2c2a179, 32'h41822d6b, 32'h40f5f9d3, 32'h425faf07, 32'h42b1e8c1, 32'h424a2c06};
test_output[39264:39271] = '{32'h42975c05, 32'h40218aff, 32'h0, 32'h41822d6b, 32'h40f5f9d3, 32'h425faf07, 32'h42b1e8c1, 32'h424a2c06};
test_input[39272:39279] = '{32'hc22fdfb9, 32'h412198c0, 32'h41802a92, 32'hc2606d87, 32'h4201976b, 32'h42b75faf, 32'hc21d8e7c, 32'hc2b10cc6};
test_output[39272:39279] = '{32'h0, 32'h412198c0, 32'h41802a92, 32'h0, 32'h4201976b, 32'h42b75faf, 32'h0, 32'h0};
test_input[39280:39287] = '{32'hc151857d, 32'hc2988815, 32'hc297b10f, 32'hc1ffa4fe, 32'h42a3693a, 32'hc1efea48, 32'hc2bc02ad, 32'hc1a98492};
test_output[39280:39287] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a3693a, 32'h0, 32'h0, 32'h0};
test_input[39288:39295] = '{32'h428a0d2d, 32'h41af21d9, 32'hc20d0575, 32'hc2ad0a0e, 32'h42116490, 32'hc2b7df0d, 32'h42087b36, 32'hc16749eb};
test_output[39288:39295] = '{32'h428a0d2d, 32'h41af21d9, 32'h0, 32'h0, 32'h42116490, 32'h0, 32'h42087b36, 32'h0};
test_input[39296:39303] = '{32'hc20395e5, 32'h429ed1e8, 32'h423a774a, 32'hc214816d, 32'hc2b1e0a9, 32'hc25108cd, 32'h426657e2, 32'h42b2f26f};
test_output[39296:39303] = '{32'h0, 32'h429ed1e8, 32'h423a774a, 32'h0, 32'h0, 32'h0, 32'h426657e2, 32'h42b2f26f};
test_input[39304:39311] = '{32'h42881791, 32'hc26495ed, 32'hc1749c0b, 32'h428a4a6a, 32'h421afdbb, 32'hc29587b6, 32'hc05d537a, 32'hc18c77dc};
test_output[39304:39311] = '{32'h42881791, 32'h0, 32'h0, 32'h428a4a6a, 32'h421afdbb, 32'h0, 32'h0, 32'h0};
test_input[39312:39319] = '{32'h42c69dd9, 32'hc2160dc3, 32'hc0fe2d5b, 32'h40fad3af, 32'h42c2a33b, 32'h40de3433, 32'h41a7e49c, 32'hc19e1639};
test_output[39312:39319] = '{32'h42c69dd9, 32'h0, 32'h0, 32'h40fad3af, 32'h42c2a33b, 32'h40de3433, 32'h41a7e49c, 32'h0};
test_input[39320:39327] = '{32'hc2ab1586, 32'hc21ee651, 32'h41349bf8, 32'h4291450c, 32'hc2a869cd, 32'hc19c384a, 32'hc2929c6b, 32'hc28b7548};
test_output[39320:39327] = '{32'h0, 32'h0, 32'h41349bf8, 32'h4291450c, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[39328:39335] = '{32'hc0782b20, 32'hc1e2bfab, 32'hc204dab7, 32'h4298d730, 32'h428871e5, 32'hc1dccd90, 32'h41ed40b5, 32'h421b582b};
test_output[39328:39335] = '{32'h0, 32'h0, 32'h0, 32'h4298d730, 32'h428871e5, 32'h0, 32'h41ed40b5, 32'h421b582b};
test_input[39336:39343] = '{32'h428ee13a, 32'hc22a4670, 32'hc2c08ea7, 32'hc23545b5, 32'h42b03eac, 32'hc2ae1329, 32'h4297c23c, 32'h41b09c55};
test_output[39336:39343] = '{32'h428ee13a, 32'h0, 32'h0, 32'h0, 32'h42b03eac, 32'h0, 32'h4297c23c, 32'h41b09c55};
test_input[39344:39351] = '{32'hc2247fc6, 32'h42ba3154, 32'hc2218ed0, 32'hc25ac1a4, 32'h423bb507, 32'h42064db4, 32'h426b49e3, 32'h420f5304};
test_output[39344:39351] = '{32'h0, 32'h42ba3154, 32'h0, 32'h0, 32'h423bb507, 32'h42064db4, 32'h426b49e3, 32'h420f5304};
test_input[39352:39359] = '{32'h421ee9ff, 32'hc05aa9b6, 32'hc2b87457, 32'h429440ac, 32'h42098acd, 32'hc22335ab, 32'h422c189b, 32'h4242da8f};
test_output[39352:39359] = '{32'h421ee9ff, 32'h0, 32'h0, 32'h429440ac, 32'h42098acd, 32'h0, 32'h422c189b, 32'h4242da8f};
test_input[39360:39367] = '{32'hc29964c0, 32'h42953190, 32'h425653f4, 32'hc1587b40, 32'hc2aa7431, 32'hbf5d7e1e, 32'hc28c0a80, 32'h4248c22a};
test_output[39360:39367] = '{32'h0, 32'h42953190, 32'h425653f4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4248c22a};
test_input[39368:39375] = '{32'hc1bc8958, 32'h40aaadcb, 32'h429b12ac, 32'hc1da651d, 32'hc25ef985, 32'h42383f54, 32'hc0b553e6, 32'hc1483a49};
test_output[39368:39375] = '{32'h0, 32'h40aaadcb, 32'h429b12ac, 32'h0, 32'h0, 32'h42383f54, 32'h0, 32'h0};
test_input[39376:39383] = '{32'hc2c51110, 32'hc215fa28, 32'h412e3081, 32'hc21deefc, 32'h4202d92c, 32'h4268946e, 32'h4201c30a, 32'hc19e89a0};
test_output[39376:39383] = '{32'h0, 32'h0, 32'h412e3081, 32'h0, 32'h4202d92c, 32'h4268946e, 32'h4201c30a, 32'h0};
test_input[39384:39391] = '{32'hc23f4a27, 32'h42906b18, 32'hc28698b2, 32'hc29e0483, 32'hc1a90368, 32'hc274f500, 32'hc27b6b32, 32'hc1ba80c0};
test_output[39384:39391] = '{32'h0, 32'h42906b18, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[39392:39399] = '{32'hc2563a58, 32'h402ef661, 32'hc2a7be27, 32'hc29f0179, 32'hc23b3f1c, 32'h41758b10, 32'h4299234f, 32'hc261c4c4};
test_output[39392:39399] = '{32'h0, 32'h402ef661, 32'h0, 32'h0, 32'h0, 32'h41758b10, 32'h4299234f, 32'h0};
test_input[39400:39407] = '{32'h425ed9cb, 32'hc200d053, 32'h4245d7c7, 32'hc29e7dc9, 32'h42aaed77, 32'h42c45bf5, 32'hc2010e65, 32'hc2b4e2bf};
test_output[39400:39407] = '{32'h425ed9cb, 32'h0, 32'h4245d7c7, 32'h0, 32'h42aaed77, 32'h42c45bf5, 32'h0, 32'h0};
test_input[39408:39415] = '{32'h423d9bef, 32'hc0c1ade2, 32'h4224dd55, 32'h41d1a8a3, 32'hc20321ba, 32'h41ac508e, 32'hc0c8c239, 32'hc2617e98};
test_output[39408:39415] = '{32'h423d9bef, 32'h0, 32'h4224dd55, 32'h41d1a8a3, 32'h0, 32'h41ac508e, 32'h0, 32'h0};
test_input[39416:39423] = '{32'h42198fc1, 32'hc263678d, 32'hc21feda1, 32'hc2aabe0e, 32'h42ad89e8, 32'hc1a1797a, 32'hc24c623e, 32'hc266ad7d};
test_output[39416:39423] = '{32'h42198fc1, 32'h0, 32'h0, 32'h0, 32'h42ad89e8, 32'h0, 32'h0, 32'h0};
test_input[39424:39431] = '{32'h42be2cd6, 32'hc2ba961c, 32'h42745c40, 32'h40ff1648, 32'hc2125efc, 32'hc148d733, 32'hc2123c84, 32'hc2481914};
test_output[39424:39431] = '{32'h42be2cd6, 32'h0, 32'h42745c40, 32'h40ff1648, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[39432:39439] = '{32'h42a69bdc, 32'h42b1c8d5, 32'hc265cbbc, 32'hc26772e7, 32'hc2a4f98e, 32'h4200ce90, 32'h418cd91b, 32'hc26b1820};
test_output[39432:39439] = '{32'h42a69bdc, 32'h42b1c8d5, 32'h0, 32'h0, 32'h0, 32'h4200ce90, 32'h418cd91b, 32'h0};
test_input[39440:39447] = '{32'h42b0bd53, 32'h428745b5, 32'h42a9a12a, 32'hc2945e4a, 32'hc2be1221, 32'h42baa869, 32'hc2a2e754, 32'hc255b301};
test_output[39440:39447] = '{32'h42b0bd53, 32'h428745b5, 32'h42a9a12a, 32'h0, 32'h0, 32'h42baa869, 32'h0, 32'h0};
test_input[39448:39455] = '{32'hc2730f6d, 32'hc282e6bd, 32'h42adf346, 32'hc270a8f0, 32'h41aa9b4d, 32'hc1c91c65, 32'h4217253e, 32'h41ef3cd1};
test_output[39448:39455] = '{32'h0, 32'h0, 32'h42adf346, 32'h0, 32'h41aa9b4d, 32'h0, 32'h4217253e, 32'h41ef3cd1};
test_input[39456:39463] = '{32'hc248f0f9, 32'h4287006d, 32'hc18ffc2a, 32'hc15ad4a6, 32'hc2994bd6, 32'h422214f1, 32'h429c57e2, 32'hc29d5680};
test_output[39456:39463] = '{32'h0, 32'h4287006d, 32'h0, 32'h0, 32'h0, 32'h422214f1, 32'h429c57e2, 32'h0};
test_input[39464:39471] = '{32'h41b7fd4d, 32'h4113673c, 32'hc2b8a187, 32'hc292b7c9, 32'h411e5643, 32'hc21151da, 32'h416710ba, 32'hc2326b0a};
test_output[39464:39471] = '{32'h41b7fd4d, 32'h4113673c, 32'h0, 32'h0, 32'h411e5643, 32'h0, 32'h416710ba, 32'h0};
test_input[39472:39479] = '{32'hc26052ed, 32'hc209b280, 32'hc296eef9, 32'hc28884bc, 32'h42901786, 32'h422193b3, 32'hc22ec283, 32'hc21bec60};
test_output[39472:39479] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42901786, 32'h422193b3, 32'h0, 32'h0};
test_input[39480:39487] = '{32'hc2a1321a, 32'h42afae7b, 32'hc2a0493b, 32'h42c4d9e1, 32'h42a229cf, 32'h42bb05d3, 32'h41fd396c, 32'h42ad505f};
test_output[39480:39487] = '{32'h0, 32'h42afae7b, 32'h0, 32'h42c4d9e1, 32'h42a229cf, 32'h42bb05d3, 32'h41fd396c, 32'h42ad505f};
test_input[39488:39495] = '{32'hc28453d8, 32'hc273f946, 32'hc1cc3487, 32'hc1a18029, 32'h42866e8e, 32'hc2a264ef, 32'hc2b90b68, 32'h429c7603};
test_output[39488:39495] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42866e8e, 32'h0, 32'h0, 32'h429c7603};
test_input[39496:39503] = '{32'hc1f382e0, 32'hc14dd3aa, 32'hc2ae9bbc, 32'h42977204, 32'hc26c6e59, 32'h419761a4, 32'hc2171f6e, 32'h42695882};
test_output[39496:39503] = '{32'h0, 32'h0, 32'h0, 32'h42977204, 32'h0, 32'h419761a4, 32'h0, 32'h42695882};
test_input[39504:39511] = '{32'h415f0686, 32'hc21486f8, 32'hc23a0b3f, 32'hc2b789cf, 32'h42ab3348, 32'hc254f74a, 32'h42a61c90, 32'hc0d756f9};
test_output[39504:39511] = '{32'h415f0686, 32'h0, 32'h0, 32'h0, 32'h42ab3348, 32'h0, 32'h42a61c90, 32'h0};
test_input[39512:39519] = '{32'h42682341, 32'hc28b4145, 32'h4289af1b, 32'hc1c096b6, 32'hc0aca497, 32'h42873d1c, 32'h42297671, 32'hc21050bf};
test_output[39512:39519] = '{32'h42682341, 32'h0, 32'h4289af1b, 32'h0, 32'h0, 32'h42873d1c, 32'h42297671, 32'h0};
test_input[39520:39527] = '{32'hc257c8d5, 32'h410431c3, 32'h420e7b05, 32'h41009f26, 32'hbfcb330e, 32'h42bf269b, 32'hc28fb6c4, 32'hc250b0be};
test_output[39520:39527] = '{32'h0, 32'h410431c3, 32'h420e7b05, 32'h41009f26, 32'h0, 32'h42bf269b, 32'h0, 32'h0};
test_input[39528:39535] = '{32'hc2a72a39, 32'hc27253a3, 32'h4246d640, 32'hc2954ecc, 32'hc24c9fb5, 32'hc27e6900, 32'hc1f1309e, 32'h42125486};
test_output[39528:39535] = '{32'h0, 32'h0, 32'h4246d640, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42125486};
test_input[39536:39543] = '{32'hc121f754, 32'h42b23f22, 32'hc1ba43fa, 32'hc2114052, 32'hc2c5851d, 32'hc266289b, 32'hc2b6b9ff, 32'h4298ef9a};
test_output[39536:39543] = '{32'h0, 32'h42b23f22, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4298ef9a};
test_input[39544:39551] = '{32'hc1f757cc, 32'h429ea21c, 32'hc27b32c4, 32'hc2228c54, 32'hc2614f7d, 32'h42c58f46, 32'hc1b53373, 32'h42c38e4b};
test_output[39544:39551] = '{32'h0, 32'h429ea21c, 32'h0, 32'h0, 32'h0, 32'h42c58f46, 32'h0, 32'h42c38e4b};
test_input[39552:39559] = '{32'hc2a20935, 32'hc145022a, 32'hc292062d, 32'h4296d961, 32'h420cc5a0, 32'hc29d44b8, 32'hc27b57d7, 32'h427fcbaa};
test_output[39552:39559] = '{32'h0, 32'h0, 32'h0, 32'h4296d961, 32'h420cc5a0, 32'h0, 32'h0, 32'h427fcbaa};
test_input[39560:39567] = '{32'hc18c01fa, 32'h40f754a9, 32'h426c2f48, 32'hc213d829, 32'hc238889d, 32'hc215782b, 32'hc2874985, 32'h41b24682};
test_output[39560:39567] = '{32'h0, 32'h40f754a9, 32'h426c2f48, 32'h0, 32'h0, 32'h0, 32'h0, 32'h41b24682};
test_input[39568:39575] = '{32'hc29bb71c, 32'hc2b7ff13, 32'h41b0664e, 32'hc05d20e7, 32'hc28ac1ae, 32'h42a4332f, 32'h4187485a, 32'hc21f68d0};
test_output[39568:39575] = '{32'h0, 32'h0, 32'h41b0664e, 32'h0, 32'h0, 32'h42a4332f, 32'h4187485a, 32'h0};
test_input[39576:39583] = '{32'h42062133, 32'h42153353, 32'hc23f6d25, 32'hc28b4acd, 32'hc20f724b, 32'hc2b659e3, 32'hc206e06f, 32'hc2911520};
test_output[39576:39583] = '{32'h42062133, 32'h42153353, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[39584:39591] = '{32'h42bacbd5, 32'hc07da510, 32'hc258606a, 32'h41df1b3b, 32'hc21d78f5, 32'h42c3e47e, 32'h42a2dbf4, 32'hc00ab64c};
test_output[39584:39591] = '{32'h42bacbd5, 32'h0, 32'h0, 32'h41df1b3b, 32'h0, 32'h42c3e47e, 32'h42a2dbf4, 32'h0};
test_input[39592:39599] = '{32'hc2ac3ac8, 32'h421c2c84, 32'h429dc555, 32'h42a6bcff, 32'hc2419eb5, 32'h4108d66c, 32'h425cf87a, 32'h402e5535};
test_output[39592:39599] = '{32'h0, 32'h421c2c84, 32'h429dc555, 32'h42a6bcff, 32'h0, 32'h4108d66c, 32'h425cf87a, 32'h402e5535};
test_input[39600:39607] = '{32'hc1c6319a, 32'hc21f1e59, 32'h4200acee, 32'hc29bea76, 32'h4217afd7, 32'h42959100, 32'hc2bea75a, 32'hc2c4f57d};
test_output[39600:39607] = '{32'h0, 32'h0, 32'h4200acee, 32'h0, 32'h4217afd7, 32'h42959100, 32'h0, 32'h0};
test_input[39608:39615] = '{32'h42afbfe2, 32'h41b0d862, 32'h42be8a1b, 32'hc1bb51f2, 32'h429659a3, 32'h40ad7440, 32'h425053fe, 32'h42b802cc};
test_output[39608:39615] = '{32'h42afbfe2, 32'h41b0d862, 32'h42be8a1b, 32'h0, 32'h429659a3, 32'h40ad7440, 32'h425053fe, 32'h42b802cc};
test_input[39616:39623] = '{32'hc01326e3, 32'hc2214eb3, 32'hc2c7c1c7, 32'hc2481b13, 32'h41afa066, 32'hc1fd5b2e, 32'h42662b96, 32'h42a1ce04};
test_output[39616:39623] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h41afa066, 32'h0, 32'h42662b96, 32'h42a1ce04};
test_input[39624:39631] = '{32'h428dba98, 32'hc2c49851, 32'hc28269cc, 32'hc27a0b1e, 32'h41fa8475, 32'hc229c33b, 32'h42a3a1d3, 32'h40976ea2};
test_output[39624:39631] = '{32'h428dba98, 32'h0, 32'h0, 32'h0, 32'h41fa8475, 32'h0, 32'h42a3a1d3, 32'h40976ea2};
test_input[39632:39639] = '{32'hc1f4a635, 32'h3fb09b9e, 32'hc2acb878, 32'h420c6603, 32'hc283839d, 32'hc2b39c5e, 32'hc29e87e9, 32'hc228105a};
test_output[39632:39639] = '{32'h0, 32'h3fb09b9e, 32'h0, 32'h420c6603, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[39640:39647] = '{32'hc0e7a78a, 32'h42c72864, 32'hc1dfb7bf, 32'h42bb8e2f, 32'h42987cc3, 32'h428bcff1, 32'h4280beef, 32'hc22b24f9};
test_output[39640:39647] = '{32'h0, 32'h42c72864, 32'h0, 32'h42bb8e2f, 32'h42987cc3, 32'h428bcff1, 32'h4280beef, 32'h0};
test_input[39648:39655] = '{32'h42696903, 32'hc167ffc8, 32'h41a871a3, 32'hc290245f, 32'hc28e9ebf, 32'hc1a1faf6, 32'hc1df7d5d, 32'hc2ac5b95};
test_output[39648:39655] = '{32'h42696903, 32'h0, 32'h41a871a3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[39656:39663] = '{32'hc0330382, 32'hc2902010, 32'h415c3f16, 32'hc2423006, 32'h424cb6db, 32'h423b592b, 32'hc2529a57, 32'hc11f59b5};
test_output[39656:39663] = '{32'h0, 32'h0, 32'h415c3f16, 32'h0, 32'h424cb6db, 32'h423b592b, 32'h0, 32'h0};
test_input[39664:39671] = '{32'h41a0247c, 32'hbffd19c2, 32'hc2989200, 32'hc2aa0a63, 32'hc28919b4, 32'h42a6218b, 32'h3fea51ce, 32'hc2bedfa4};
test_output[39664:39671] = '{32'h41a0247c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42a6218b, 32'h3fea51ce, 32'h0};
test_input[39672:39679] = '{32'hc2a83c05, 32'hc22ffdf5, 32'h42973f53, 32'hc118736a, 32'hc2b18f0c, 32'h420f204e, 32'hc173ca3f, 32'h419f3b0f};
test_output[39672:39679] = '{32'h0, 32'h0, 32'h42973f53, 32'h0, 32'h0, 32'h420f204e, 32'h0, 32'h419f3b0f};
test_input[39680:39687] = '{32'hc2a733dd, 32'h4255420d, 32'hc200c2f4, 32'h420c407a, 32'h4129d384, 32'hc1be2018, 32'h428cf843, 32'h42b595e1};
test_output[39680:39687] = '{32'h0, 32'h4255420d, 32'h0, 32'h420c407a, 32'h4129d384, 32'h0, 32'h428cf843, 32'h42b595e1};
test_input[39688:39695] = '{32'hc27fa268, 32'h42a0825a, 32'hc2345383, 32'hc2748e05, 32'h42737715, 32'hc18d9b6f, 32'hc1790819, 32'h429fe0a3};
test_output[39688:39695] = '{32'h0, 32'h42a0825a, 32'h0, 32'h0, 32'h42737715, 32'h0, 32'h0, 32'h429fe0a3};
test_input[39696:39703] = '{32'h41745e5d, 32'h41e9d4f7, 32'hc084424a, 32'h42a2b7f1, 32'hc2b32f07, 32'hc1af7ffd, 32'hc11ba1fe, 32'h42907792};
test_output[39696:39703] = '{32'h41745e5d, 32'h41e9d4f7, 32'h0, 32'h42a2b7f1, 32'h0, 32'h0, 32'h0, 32'h42907792};
test_input[39704:39711] = '{32'hc27c3636, 32'hc2947102, 32'h426703ef, 32'h4256a41d, 32'hc2c31e3c, 32'hc29066f4, 32'h42085a96, 32'hc1efb997};
test_output[39704:39711] = '{32'h0, 32'h0, 32'h426703ef, 32'h4256a41d, 32'h0, 32'h0, 32'h42085a96, 32'h0};
test_input[39712:39719] = '{32'h41c58600, 32'h429ef7fc, 32'h42c49d73, 32'h42677c79, 32'h4280768a, 32'hc2bcc0c9, 32'h4282833f, 32'hc2a10dff};
test_output[39712:39719] = '{32'h41c58600, 32'h429ef7fc, 32'h42c49d73, 32'h42677c79, 32'h4280768a, 32'h0, 32'h4282833f, 32'h0};
test_input[39720:39727] = '{32'hc2bc9fbd, 32'hc2872185, 32'h42198141, 32'h422cae81, 32'h41f7046c, 32'hc14f44c8, 32'h4221eee1, 32'h42a5350d};
test_output[39720:39727] = '{32'h0, 32'h0, 32'h42198141, 32'h422cae81, 32'h41f7046c, 32'h0, 32'h4221eee1, 32'h42a5350d};
test_input[39728:39735] = '{32'hc2259ccb, 32'hc24bf233, 32'hc28c84f8, 32'hc27b0e5e, 32'h42a4e0f9, 32'hc25d6b61, 32'h42ab9a07, 32'hc23476fa};
test_output[39728:39735] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h42a4e0f9, 32'h0, 32'h42ab9a07, 32'h0};
test_input[39736:39743] = '{32'hc2c72bec, 32'h42c52642, 32'hc284c0fd, 32'hc0219bf6, 32'h412489f7, 32'h408b93fb, 32'hc28c8aa6, 32'h41ae1a35};
test_output[39736:39743] = '{32'h0, 32'h42c52642, 32'h0, 32'h0, 32'h412489f7, 32'h408b93fb, 32'h0, 32'h41ae1a35};
test_input[39744:39751] = '{32'hc2898046, 32'hc167fb46, 32'hc2c72fd9, 32'h42a4656b, 32'h4231bf82, 32'hc29767f4, 32'hc296b2e9, 32'hc06525e0};
test_output[39744:39751] = '{32'h0, 32'h0, 32'h0, 32'h42a4656b, 32'h4231bf82, 32'h0, 32'h0, 32'h0};
test_input[39752:39759] = '{32'h41ecd353, 32'hc27f276c, 32'h42bfd6b4, 32'hc24f6964, 32'h42a682ec, 32'h42ad6706, 32'h42a13256, 32'hc2971022};
test_output[39752:39759] = '{32'h41ecd353, 32'h0, 32'h42bfd6b4, 32'h0, 32'h42a682ec, 32'h42ad6706, 32'h42a13256, 32'h0};
test_input[39760:39767] = '{32'h41f0cdf6, 32'h4090a6c6, 32'hc1c716e7, 32'hc2bd3f43, 32'hc066fde2, 32'h426596fe, 32'hc0ec3734, 32'h429f0f93};
test_output[39760:39767] = '{32'h41f0cdf6, 32'h4090a6c6, 32'h0, 32'h0, 32'h0, 32'h426596fe, 32'h0, 32'h429f0f93};
test_input[39768:39775] = '{32'hc27eef2c, 32'h42110537, 32'h42b90d12, 32'hc173a488, 32'hc1fc9309, 32'hc2386445, 32'hc2b8e7c1, 32'h4104eee7};
test_output[39768:39775] = '{32'h0, 32'h42110537, 32'h42b90d12, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4104eee7};
test_input[39776:39783] = '{32'h426f4a4c, 32'h40c4865c, 32'h4173d2e6, 32'hc22d5f07, 32'h42c6e18b, 32'h41deca29, 32'h423f84c0, 32'hc1ac4ad5};
test_output[39776:39783] = '{32'h426f4a4c, 32'h40c4865c, 32'h4173d2e6, 32'h0, 32'h42c6e18b, 32'h41deca29, 32'h423f84c0, 32'h0};
test_input[39784:39791] = '{32'h41eee728, 32'h429a34c0, 32'h42a671f0, 32'hc28192b0, 32'hc21357bd, 32'h423b6757, 32'h4230e51c, 32'h420fc79e};
test_output[39784:39791] = '{32'h41eee728, 32'h429a34c0, 32'h42a671f0, 32'h0, 32'h0, 32'h423b6757, 32'h4230e51c, 32'h420fc79e};
test_input[39792:39799] = '{32'hc0b9b21a, 32'h42a52343, 32'hc25e3e80, 32'h40996323, 32'h421756ac, 32'hc1e5f9ce, 32'hc228bdc5, 32'hc29a97f1};
test_output[39792:39799] = '{32'h0, 32'h42a52343, 32'h0, 32'h40996323, 32'h421756ac, 32'h0, 32'h0, 32'h0};
test_input[39800:39807] = '{32'hc2bc6f6b, 32'hc20362a3, 32'h41daa53c, 32'hc2a8785e, 32'h4038f530, 32'h41a8d87c, 32'hc14875f1, 32'hc112b575};
test_output[39800:39807] = '{32'h0, 32'h0, 32'h41daa53c, 32'h0, 32'h4038f530, 32'h41a8d87c, 32'h0, 32'h0};
test_input[39808:39815] = '{32'hc1902d5d, 32'hc24aae44, 32'hc1c86c4b, 32'h42a25d6c, 32'h42b62d85, 32'h42b4212e, 32'hc2065aa3, 32'h41abb744};
test_output[39808:39815] = '{32'h0, 32'h0, 32'h0, 32'h42a25d6c, 32'h42b62d85, 32'h42b4212e, 32'h0, 32'h41abb744};
test_input[39816:39823] = '{32'hc232a46b, 32'hc29acd8e, 32'h42921651, 32'h4218a78f, 32'hc19bf3d5, 32'h4225bfea, 32'h42c77f5d, 32'hc2402727};
test_output[39816:39823] = '{32'h0, 32'h0, 32'h42921651, 32'h4218a78f, 32'h0, 32'h4225bfea, 32'h42c77f5d, 32'h0};
test_input[39824:39831] = '{32'hc1d65567, 32'hc2b33599, 32'h42620bae, 32'hc2a0061d, 32'h4266312d, 32'h4087af39, 32'hbf5891a5, 32'h415d758a};
test_output[39824:39831] = '{32'h0, 32'h0, 32'h42620bae, 32'h0, 32'h4266312d, 32'h4087af39, 32'h0, 32'h415d758a};
test_input[39832:39839] = '{32'hc102cf53, 32'h4222da86, 32'h4280cc96, 32'hc158106d, 32'h42443670, 32'hc26f9ea8, 32'hc26ea8d0, 32'h42a3c32f};
test_output[39832:39839] = '{32'h0, 32'h4222da86, 32'h4280cc96, 32'h0, 32'h42443670, 32'h0, 32'h0, 32'h42a3c32f};
test_input[39840:39847] = '{32'h41d82304, 32'hc225fcd8, 32'hc2c3c1d9, 32'h40d4899f, 32'h4196d171, 32'h41b7f69f, 32'h4284088b, 32'h417235c6};
test_output[39840:39847] = '{32'h41d82304, 32'h0, 32'h0, 32'h40d4899f, 32'h4196d171, 32'h41b7f69f, 32'h4284088b, 32'h417235c6};
test_input[39848:39855] = '{32'h42593ebc, 32'hc2457ed9, 32'h421c479b, 32'h41a83563, 32'h410ff5fa, 32'h41470a9e, 32'h41b69328, 32'hc2a9cc51};
test_output[39848:39855] = '{32'h42593ebc, 32'h0, 32'h421c479b, 32'h41a83563, 32'h410ff5fa, 32'h41470a9e, 32'h41b69328, 32'h0};
test_input[39856:39863] = '{32'hc0dc4072, 32'hc29a9457, 32'hc09899da, 32'h41fea5b4, 32'hc2b25fa7, 32'h3fb0c3dc, 32'h42509d0b, 32'h420ee581};
test_output[39856:39863] = '{32'h0, 32'h0, 32'h0, 32'h41fea5b4, 32'h0, 32'h3fb0c3dc, 32'h42509d0b, 32'h420ee581};
test_input[39864:39871] = '{32'hc1b8dd3c, 32'hc2b2f2ee, 32'h42a7c9cc, 32'hc24a7f8f, 32'h410836d3, 32'h41866c9a, 32'h410e14e9, 32'h4221e09a};
test_output[39864:39871] = '{32'h0, 32'h0, 32'h42a7c9cc, 32'h0, 32'h410836d3, 32'h41866c9a, 32'h410e14e9, 32'h4221e09a};
test_input[39872:39879] = '{32'hc1bbcf4a, 32'hc2a86cef, 32'h41df82ba, 32'h42be5a7f, 32'h42a6066d, 32'h428d0eba, 32'h40bbad52, 32'h42b6c402};
test_output[39872:39879] = '{32'h0, 32'h0, 32'h41df82ba, 32'h42be5a7f, 32'h42a6066d, 32'h428d0eba, 32'h40bbad52, 32'h42b6c402};
test_input[39880:39887] = '{32'hc25e0820, 32'hc0e11de7, 32'hc2c526a9, 32'hc1667e7f, 32'h427e582f, 32'h42083ca6, 32'h41c9cc4c, 32'h4130f852};
test_output[39880:39887] = '{32'h0, 32'h0, 32'h0, 32'h0, 32'h427e582f, 32'h42083ca6, 32'h41c9cc4c, 32'h4130f852};
test_input[39888:39895] = '{32'h418a561a, 32'hc248e3e7, 32'h418b17a4, 32'h424ad2f4, 32'h42b2b90b, 32'h421f9976, 32'h42838732, 32'h3f88771d};
test_output[39888:39895] = '{32'h418a561a, 32'h0, 32'h418b17a4, 32'h424ad2f4, 32'h42b2b90b, 32'h421f9976, 32'h42838732, 32'h3f88771d};
test_input[39896:39903] = '{32'h41ef6a7f, 32'hc2be1a3a, 32'h41091cd1, 32'h421b8033, 32'h428d0e22, 32'hc17bb517, 32'h42242c0e, 32'h42aed7fc};
test_output[39896:39903] = '{32'h41ef6a7f, 32'h0, 32'h41091cd1, 32'h421b8033, 32'h428d0e22, 32'h0, 32'h42242c0e, 32'h42aed7fc};
test_input[39904:39911] = '{32'hc2590fcb, 32'h428fd998, 32'h42733b1e, 32'hc29c53cb, 32'hc183f548, 32'hc1b9b587, 32'hc2ab976c, 32'hc2a8bf49};
test_output[39904:39911] = '{32'h0, 32'h428fd998, 32'h42733b1e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[39912:39919] = '{32'hc27044be, 32'hc2989af4, 32'h429feb50, 32'h42a7d4af, 32'hc2369141, 32'h41e8b6fc, 32'h428ad1dc, 32'h414c343e};
test_output[39912:39919] = '{32'h0, 32'h0, 32'h429feb50, 32'h42a7d4af, 32'h0, 32'h41e8b6fc, 32'h428ad1dc, 32'h414c343e};
test_input[39920:39927] = '{32'hc166ac97, 32'h427dd83c, 32'h4197a347, 32'h41ce4b1e, 32'h4292bff8, 32'h428eba7e, 32'hc2bb5175, 32'h40962a3f};
test_output[39920:39927] = '{32'h0, 32'h427dd83c, 32'h4197a347, 32'h41ce4b1e, 32'h4292bff8, 32'h428eba7e, 32'h0, 32'h40962a3f};
test_input[39928:39935] = '{32'h41849f2f, 32'h41cc8fbd, 32'hc2aaa5bc, 32'h4231f15e, 32'h42a635c4, 32'hc26662de, 32'hc2117c4c, 32'hc200dc19};
test_output[39928:39935] = '{32'h41849f2f, 32'h41cc8fbd, 32'h0, 32'h4231f15e, 32'h42a635c4, 32'h0, 32'h0, 32'h0};
test_input[39936:39943] = '{32'hc2acb6a9, 32'h42480f0c, 32'hc2839f2e, 32'hc06a7ee0, 32'h4239976d, 32'h42595b42, 32'hc2a7a1e9, 32'hc1d68294};
test_output[39936:39943] = '{32'h0, 32'h42480f0c, 32'h0, 32'h0, 32'h4239976d, 32'h42595b42, 32'h0, 32'h0};
test_input[39944:39951] = '{32'h42763ed5, 32'h404b0c3e, 32'h4200a363, 32'hbf356f8f, 32'hc2b09656, 32'h4278a3f1, 32'hc22527d1, 32'h429a9bc0};
test_output[39944:39951] = '{32'h42763ed5, 32'h404b0c3e, 32'h4200a363, 32'h0, 32'h0, 32'h4278a3f1, 32'h0, 32'h429a9bc0};
test_input[39952:39959] = '{32'h42897b1d, 32'hc261f371, 32'hc1310a99, 32'hc19500d7, 32'h41803882, 32'h42b2f052, 32'hc2451b04, 32'hc0f1f547};
test_output[39952:39959] = '{32'h42897b1d, 32'h0, 32'h0, 32'h0, 32'h41803882, 32'h42b2f052, 32'h0, 32'h0};
test_input[39960:39967] = '{32'h429bc615, 32'hc1ab9dcf, 32'h42075aa1, 32'h4243708f, 32'hc255330a, 32'hc21f7b35, 32'hc1e033ea, 32'hc2a8d3b7};
test_output[39960:39967] = '{32'h429bc615, 32'h0, 32'h42075aa1, 32'h4243708f, 32'h0, 32'h0, 32'h0, 32'h0};
test_input[39968:39975] = '{32'hc189e257, 32'h42008349, 32'h4280d1ae, 32'h417c16bc, 32'hc2374294, 32'hc24cd194, 32'hc0e83ff1, 32'h4287f607};
test_output[39968:39975] = '{32'h0, 32'h42008349, 32'h4280d1ae, 32'h417c16bc, 32'h0, 32'h0, 32'h0, 32'h4287f607};
test_input[39976:39983] = '{32'h403310bd, 32'h427c5348, 32'h42485bab, 32'hc271dfab, 32'h41a4c2c7, 32'h41ae10f8, 32'h41000d1d, 32'h42a8aab2};
test_output[39976:39983] = '{32'h403310bd, 32'h427c5348, 32'h42485bab, 32'h0, 32'h41a4c2c7, 32'h41ae10f8, 32'h41000d1d, 32'h42a8aab2};
test_input[39984:39991] = '{32'h4136acd3, 32'hc28899b2, 32'hc204ff45, 32'hc2be00fb, 32'hc13742c9, 32'hc14e081e, 32'h426a5a2f, 32'h42b096c5};
test_output[39984:39991] = '{32'h4136acd3, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h426a5a2f, 32'h42b096c5};
test_input[39992:39999] = '{32'hc2c50650, 32'h42a92bff, 32'hc29834ce, 32'h42c46845, 32'hc25a0858, 32'h42c709f6, 32'hc185bacb, 32'hc2b7c579};
test_output[39992:39999] = '{32'h0, 32'h42a92bff, 32'h0, 32'h42c46845, 32'h0, 32'h42c709f6, 32'h0, 32'h0};
end
`endif
