`timescale 1ns/1ns

module conv_forward_layer_tb();

	parameter CYCLE			= 2;
	parameter MULT_DELAY		= 5;
	parameter ADD_DELAY		= 7;
	parameter WIDTH			= 8;
	
	parameter NUM_TESTS		= 10000;
	parameter NUM_COLS		= (WIDTH*2) +2;
	parameter MEM_SIZE		= NUM_TESTS*NUM_COLS; 

	reg clk, reset, enable;
	logic [31:0] in_vec [WIDTH-1:0];
	logic [31:0] weight_vec [WIDTH-1:0];
	logic [31:0] bias_term;
	logic [31:0] out;
	reg [31:0] mem [MEM_SIZE];
	int count;
	
	//forever cycle the clk
	
	
	
//	conv_forward_layer 	#(.WIDTH(WIDTH))
//						conv_forward_inst(
//							.clk(clk),
//							.reset(reset),
//							.enable(enable),
//							.in_data(in_vec),
//							.weights(weight_vec),
//							.out_data(out)
//						);
	float_add float_add_inst(
												.aclr(!enable),
												.clock(clk),
												.dataa(in_vec[0]),
												.datab(weight_vec[0]),
												.result(out)
												);					
	
	always @(posedge clk) begin
		count = count + 1;
	end
	
	int i, j;
	initial begin
		clk = 0;
		forever #(CYCLE) clk = ~clk;
		reset = 0;
		enable = 0;
		out = 0;
		#(CYCLE*2)
		enable = 1;
		#(CYCLE*2)
		
		#1 $display("clk1: %d\n", clk);
		$display("count: %d\n", count);
		#1 $display("clk2: %d\n", clk);
		$display("count: %d\n", count);
		#1 $display("clk3: %d\n", clk);
		$display("count: %d\n", count);
		#1 $display("clk4: %d\n", clk);
		$display("count: %d\n", count);
		#1 $display("clk5: %d\n", clk);
		$display("count: %d\n", count);
		#1 $display("clk6: %d\n", clk);
		#1 $display("clk7: %d\n", clk);
		#1 $display("clk8: %d\n", clk);
		//read the test data generated by Python into memory
		$readmemh("/home/b/FPGA-CNN/test/test_data/conv_forward_test_data.hex", mem);
		//for all test cases
		 for (i = 0; i < MEM_SIZE/1000; i=i+NUM_COLS) begin
			//copy input to register
			for (j = 0; j < WIDTH; j++) begin
				in_vec[j] = mem[i+j];
			end
			//copy weight vector to register
			for (j = 0; j < WIDTH; j++) begin
				weight_vec[j] = mem[i+WIDTH+j];
			end
			//read bias term 
			bias_term = mem[i+2*WIDTH+1];
			
			//wait for it...
			//#(CYCLE*(MULT_DELAY + ADD_DELAY*WIDTH)+100)
			#(CYCLE*20)
			//check output
//			$display("in_vec: %b", in_vec[0]);
//			$display("we_vec: %b", weight_vec[0]);
//			$display("out: %b", out);
//			$display("mem: %b", mem[i+2*WIDTH]);
			assert( out == mem[i+2*WIDTH] );
			//increment twice to skip output val and bias_term, once to move pointer
			//i = i + 3;
		end
		$display("############################################\n");
		$display("All tests passed!\n");
		$display("############################################\n");
	end

endmodule
