//====================================================================
//
// interfaces.sv
//
// Original Author : George Powley
// Original Date   : 2015/01/21
//
// Copyright (c) 2015 Intel Corporation
// Intel Proprietary
//
// Description:
//  - All interfaces must be included here
//====================================================================

`include "spl_iface.sv"
`include "afu_iface.sv"
`include "sw_iface.sv"
