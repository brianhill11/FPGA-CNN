`ifndef CONV_FORWARD_TEST_H
`define CONV_FORWARD_TEST_H
reg [31:0] test_input [80000];
reg [31:0] test_output [10000];
reg [31:0] test_index [10000];
initial begin
test_input[0:7] = '{32'h4228e6a9, 32'hc1efaffd, 32'hc23e2aee, 32'hc11d9607, 32'hc220aeec, 32'h42a6336e, 32'hc2a80d82, 32'h4201f10f};
test_output[0] = '{32'h42a6336e};
test_index[0] = '{5};
test_input[8:15] = '{32'h425d5f52, 32'hc2be8707, 32'h4192547a, 32'h42bf2cf1, 32'hc212a717, 32'h42bd9cbb, 32'hc204c6f0, 32'h42ad4885};
test_output[1] = '{32'h42bf2cf1};
test_index[1] = '{3};
test_input[16:23] = '{32'h425d2cea, 32'h42a0ad9d, 32'hc29fe83a, 32'hc2b27e38, 32'h4233be3d, 32'h42aaf55d, 32'hc1357b90, 32'hbec4b965};
test_output[2] = '{32'h42aaf55d};
test_index[2] = '{5};
test_input[24:31] = '{32'h42a7a487, 32'h42204756, 32'h4279fd75, 32'hc23540c2, 32'h42bca100, 32'hc28c0ddd, 32'h42be037a, 32'hc16e243c};
test_output[3] = '{32'h42be037a};
test_index[3] = '{6};
test_input[32:39] = '{32'hc2a58d4e, 32'hc1923fd4, 32'hbfa462e4, 32'hc2767b89, 32'h429d1732, 32'hc15df575, 32'hc0e16091, 32'h429c06d6};
test_output[4] = '{32'h429d1732};
test_index[4] = '{4};
test_input[40:47] = '{32'hc1235be0, 32'h426336bd, 32'hc0b86901, 32'h42c11d1c, 32'hc23a9dc9, 32'h425c8a6c, 32'h4232a4cc, 32'h418ff52d};
test_output[5] = '{32'h42c11d1c};
test_index[5] = '{3};
test_input[48:55] = '{32'hc2827123, 32'hc28a9be2, 32'hc287e9ca, 32'hc291b029, 32'hc2b0bc44, 32'h4220516a, 32'h426b7bb9, 32'hc2b26735};
test_output[6] = '{32'h426b7bb9};
test_index[6] = '{6};
test_input[56:63] = '{32'h408f70bb, 32'hc26325c1, 32'hc2c12fc3, 32'hc293e80b, 32'h4191b51a, 32'h4244b9e7, 32'h42bc4ba8, 32'h42b525f3};
test_output[7] = '{32'h42bc4ba8};
test_index[7] = '{6};
test_input[64:71] = '{32'h428288af, 32'hc2b92f0a, 32'hc18ea877, 32'hc2869ad8, 32'h41e6c7a6, 32'hc26e90ef, 32'hc24034be, 32'h41e37d3f};
test_output[8] = '{32'h428288af};
test_index[8] = '{0};
test_input[72:79] = '{32'h41dfd351, 32'hc274eb08, 32'hc2a5c3ba, 32'h42b5c8b0, 32'hc12ec700, 32'h420e1a91, 32'h42703662, 32'hc208e6af};
test_output[9] = '{32'h42b5c8b0};
test_index[9] = '{3};
test_input[80:87] = '{32'hc28a2b04, 32'hc28dd6cf, 32'h42098c74, 32'h4240eccf, 32'hc17befe6, 32'h4258d950, 32'hc2598e35, 32'hc13ba7fb};
test_output[10] = '{32'h4258d950};
test_index[10] = '{5};
test_input[88:95] = '{32'h42a0c2c6, 32'h429d20ff, 32'hc1c406e5, 32'hc25ec1a8, 32'hc28eab94, 32'hc284d1d5, 32'hc1889be6, 32'hc1b3f9db};
test_output[11] = '{32'h42a0c2c6};
test_index[11] = '{0};
test_input[96:103] = '{32'h42622922, 32'hc2adeb5d, 32'hc2572866, 32'h424e6303, 32'h42a8e39b, 32'hc29cd4f0, 32'h40011e39, 32'hc04c46ff};
test_output[12] = '{32'h42a8e39b};
test_index[12] = '{4};
test_input[104:111] = '{32'h4226c2a2, 32'hc283e2b9, 32'h409c4737, 32'h41c119f1, 32'hc25129e6, 32'h42c4f232, 32'h423d42d9, 32'hc2be6bf5};
test_output[13] = '{32'h42c4f232};
test_index[13] = '{5};
test_input[112:119] = '{32'h42905f4a, 32'hc29720c4, 32'hc1f382a6, 32'h42c72984, 32'hc270c102, 32'h41237a7f, 32'h416e1d07, 32'h4172a536};
test_output[14] = '{32'h42c72984};
test_index[14] = '{3};
test_input[120:127] = '{32'h424394f7, 32'hc10b19cd, 32'h42a9a387, 32'h42a0062c, 32'h42c11f84, 32'hc21d0568, 32'hc23a54d4, 32'h4123d06f};
test_output[15] = '{32'h42c11f84};
test_index[15] = '{4};
test_input[128:135] = '{32'hc1afc650, 32'hc2c6f290, 32'hc1b58758, 32'hc1fde1c8, 32'hc2ae79dd, 32'hc1edb884, 32'h42897555, 32'hc1d29dfe};
test_output[16] = '{32'h42897555};
test_index[16] = '{6};
test_input[136:143] = '{32'hc190bc2a, 32'hc2399da6, 32'h420be6db, 32'hc187562a, 32'hc2876838, 32'hc282e7b7, 32'h41876d03, 32'h4242c0f3};
test_output[17] = '{32'h4242c0f3};
test_index[17] = '{7};
test_input[144:151] = '{32'hc165f623, 32'hc188f0d7, 32'h419bd3b9, 32'hc0ef6a6e, 32'h42395eb8, 32'hc179ea45, 32'h41328507, 32'hc09d6e06};
test_output[18] = '{32'h42395eb8};
test_index[18] = '{4};
test_input[152:159] = '{32'h429b4383, 32'h42102e43, 32'h42aefd52, 32'hc28fe3a3, 32'h42856cfb, 32'h42115524, 32'hbf3e8328, 32'h42b0a5a0};
test_output[19] = '{32'h42b0a5a0};
test_index[19] = '{7};
test_input[160:167] = '{32'h41c2b5d4, 32'hc20701f2, 32'hc28f30df, 32'h41cf3f4a, 32'hc1cfc320, 32'h42c182ad, 32'hc2bdc642, 32'h42a4f583};
test_output[20] = '{32'h42c182ad};
test_index[20] = '{5};
test_input[168:175] = '{32'hc1cf9edc, 32'h42873713, 32'hc203c2a0, 32'hbff4e2db, 32'hc1b2e709, 32'h42a2faf3, 32'hc22c578f, 32'h422633a1};
test_output[21] = '{32'h42a2faf3};
test_index[21] = '{5};
test_input[176:183] = '{32'hc29e1e6a, 32'h41d991e1, 32'h42a6e4c8, 32'hc11c30ac, 32'h42491cdf, 32'h4237605a, 32'h4205b883, 32'hc20c96f8};
test_output[22] = '{32'h42a6e4c8};
test_index[22] = '{2};
test_input[184:191] = '{32'hc1ee5f4f, 32'h425acb4e, 32'hc2865e26, 32'hc287c854, 32'hc1b486f7, 32'hc2bd0992, 32'hc12021db, 32'hc209fb7d};
test_output[23] = '{32'h425acb4e};
test_index[23] = '{1};
test_input[192:199] = '{32'hc2765435, 32'hc25ef254, 32'h41a87837, 32'h420f4435, 32'hc29b5086, 32'hc202b1b9, 32'hc1ef805d, 32'h428b96fe};
test_output[24] = '{32'h428b96fe};
test_index[24] = '{7};
test_input[200:207] = '{32'h42632fba, 32'hc24e7962, 32'h42b449ee, 32'hc25b6f18, 32'h42a4b1a3, 32'hc26da7cd, 32'h42a86980, 32'h42390088};
test_output[25] = '{32'h42b449ee};
test_index[25] = '{2};
test_input[208:215] = '{32'h42266fd7, 32'h4222d5be, 32'hc288dda7, 32'hc2a086bc, 32'hc2a54e8a, 32'hc28981df, 32'hc14a4fbc, 32'h41bed64a};
test_output[26] = '{32'h42266fd7};
test_index[26] = '{0};
test_input[216:223] = '{32'hc1f9e069, 32'hc22a7ad3, 32'h426ebccf, 32'hc2a9bf16, 32'h42149264, 32'h42bb8c6c, 32'h407e4f5a, 32'h4203a56c};
test_output[27] = '{32'h42bb8c6c};
test_index[27] = '{5};
test_input[224:231] = '{32'h41ffdcff, 32'h41b91c06, 32'h42999ed5, 32'h4281b2f7, 32'hc1fcde4e, 32'h41e1a892, 32'h42622fcc, 32'hc207ebaa};
test_output[28] = '{32'h42999ed5};
test_index[28] = '{2};
test_input[232:239] = '{32'h42aadf86, 32'h41f11fcc, 32'hc2a48a11, 32'hc12510e4, 32'h412ca339, 32'hc2a79abe, 32'hc18177d0, 32'h427c9823};
test_output[29] = '{32'h42aadf86};
test_index[29] = '{0};
test_input[240:247] = '{32'h403b8c63, 32'hc2b60f31, 32'hc2648f10, 32'h422b9c30, 32'h42a6e336, 32'hc2b58fbd, 32'hc10a2e47, 32'hc2ab95c6};
test_output[30] = '{32'h42a6e336};
test_index[30] = '{4};
test_input[248:255] = '{32'h429b45e0, 32'hc0ddeea7, 32'hc1682d13, 32'hc25fdbcb, 32'hc2107e99, 32'hc28982da, 32'hc27e2a1a, 32'hc0b58aab};
test_output[31] = '{32'h429b45e0};
test_index[31] = '{0};
test_input[256:263] = '{32'h4280a1f6, 32'h4262466d, 32'hc2a3f0ed, 32'hc2533371, 32'h427dea40, 32'hc2aeda89, 32'hc2b98c37, 32'h410d501f};
test_output[32] = '{32'h4280a1f6};
test_index[32] = '{0};
test_input[264:271] = '{32'hc2873609, 32'h42b9479c, 32'hc2345275, 32'hc28f463d, 32'h42b8cafe, 32'h428235bc, 32'h41ceba48, 32'hc20d6ba0};
test_output[33] = '{32'h42b9479c};
test_index[33] = '{1};
test_input[272:279] = '{32'hc2ade0d5, 32'h42029e5a, 32'hc21d7817, 32'hc267eb6b, 32'hc29526b5, 32'hbea5821e, 32'hc2172c09, 32'hc2c6c885};
test_output[34] = '{32'h42029e5a};
test_index[34] = '{1};
test_input[280:287] = '{32'hc2576990, 32'h423a6815, 32'h4299be0f, 32'hc2140cd9, 32'hc032d2ca, 32'hc2c04ad2, 32'hc2954eff, 32'h4082cac1};
test_output[35] = '{32'h4299be0f};
test_index[35] = '{2};
test_input[288:295] = '{32'hc21aaeff, 32'hc2a5a948, 32'h3f1c1dd5, 32'h428772f7, 32'h425aeb72, 32'h42596e0a, 32'h41a5b003, 32'h429a79a8};
test_output[36] = '{32'h429a79a8};
test_index[36] = '{7};
test_input[296:303] = '{32'hc27457aa, 32'h42a83171, 32'hc1b506d6, 32'h42c5642f, 32'h4229a6af, 32'h42b5fce6, 32'hc2b48af9, 32'h42c2470f};
test_output[37] = '{32'h42c5642f};
test_index[37] = '{3};
test_input[304:311] = '{32'h42bed08b, 32'h41a80290, 32'hc2b75534, 32'h42859f7f, 32'h4239701b, 32'h420b79fa, 32'h41c1cc1c, 32'hc1f9a0f4};
test_output[38] = '{32'h42bed08b};
test_index[38] = '{0};
test_input[312:319] = '{32'hc2239dc5, 32'hc216cbf0, 32'h4017c8e2, 32'h4145de8c, 32'hc2308dae, 32'h41a35e00, 32'hc28a1ecc, 32'hc143a96e};
test_output[39] = '{32'h41a35e00};
test_index[39] = '{5};
test_input[320:327] = '{32'hc1dcc22a, 32'h42b16c33, 32'hc2060d77, 32'h4284225a, 32'h41c7d184, 32'hc2ae855c, 32'hc1a5f780, 32'h4280b6cf};
test_output[40] = '{32'h42b16c33};
test_index[40] = '{1};
test_input[328:335] = '{32'h41a1d162, 32'h41d4a715, 32'h4041fd96, 32'hc2b21584, 32'hc2871767, 32'hc169874c, 32'h428bfb3f, 32'h41096063};
test_output[41] = '{32'h428bfb3f};
test_index[41] = '{6};
test_input[336:343] = '{32'hc28a8eed, 32'h42852288, 32'h42255700, 32'hc2b8ea05, 32'hc2bab548, 32'h4292ecda, 32'h4235b830, 32'h426af937};
test_output[42] = '{32'h4292ecda};
test_index[42] = '{5};
test_input[344:351] = '{32'h41bdae12, 32'h4228e628, 32'h42890002, 32'hc2b7fc59, 32'h425331bd, 32'h42180854, 32'h422d13c4, 32'h42b32e95};
test_output[43] = '{32'h42b32e95};
test_index[43] = '{7};
test_input[352:359] = '{32'h42094cc4, 32'h42b1a238, 32'hc26f5644, 32'h42685559, 32'hc0892e58, 32'h4283d24e, 32'h419219f2, 32'h425f07df};
test_output[44] = '{32'h42b1a238};
test_index[44] = '{1};
test_input[360:367] = '{32'h420a351e, 32'hc20d9a09, 32'h417ad7d3, 32'h428c4a0b, 32'hc20674e0, 32'h415c0610, 32'h404e0e17, 32'h409bc0c8};
test_output[45] = '{32'h428c4a0b};
test_index[45] = '{3};
test_input[368:375] = '{32'h429de55b, 32'h426a629a, 32'hc2b2db26, 32'hc2bb4850, 32'h41e0f832, 32'hc2407125, 32'h4210dd83, 32'hc2be51b7};
test_output[46] = '{32'h429de55b};
test_index[46] = '{0};
test_input[376:383] = '{32'h421ccbdc, 32'hc29cedf5, 32'h42b2155f, 32'h42ab5b60, 32'h41034174, 32'h4288d1bd, 32'hc2b851ed, 32'h4231be18};
test_output[47] = '{32'h42b2155f};
test_index[47] = '{2};
test_input[384:391] = '{32'hc26f3af2, 32'hc29c7eb0, 32'h4280d964, 32'hc0ca9493, 32'h41843dcb, 32'h41a48788, 32'h42017cd4, 32'h42b92b09};
test_output[48] = '{32'h42b92b09};
test_index[48] = '{7};
test_input[392:399] = '{32'hc2904b3e, 32'h42070632, 32'hc171a427, 32'hc2355a30, 32'hc2c4418d, 32'h42a63956, 32'h42773f3c, 32'hc257bf12};
test_output[49] = '{32'h42a63956};
test_index[49] = '{5};
test_input[400:407] = '{32'hc1fbcea6, 32'hc22c1d8d, 32'hc209b1df, 32'h41cbae6d, 32'h3ecc1963, 32'h428af20d, 32'h4250d3f7, 32'hc1fdc526};
test_output[50] = '{32'h428af20d};
test_index[50] = '{5};
test_input[408:415] = '{32'h42aed8bd, 32'hc29d6d88, 32'h42c2586e, 32'h42b86290, 32'hc28b52e2, 32'h41eed5dc, 32'hc1d8e8c0, 32'hc2460a8c};
test_output[51] = '{32'h42c2586e};
test_index[51] = '{2};
test_input[416:423] = '{32'h41c2fd5b, 32'hc0a10448, 32'h41e2db26, 32'h41801ba6, 32'hc2b49ebc, 32'h41ff75e0, 32'h42aaa5e0, 32'hc245fdd3};
test_output[52] = '{32'h42aaa5e0};
test_index[52] = '{6};
test_input[424:431] = '{32'h4290de9c, 32'h428bd848, 32'hc280debb, 32'h41fa8a04, 32'hc24f437b, 32'hc0f5cdd7, 32'hc03e8318, 32'hc2821826};
test_output[53] = '{32'h4290de9c};
test_index[53] = '{0};
test_input[432:439] = '{32'h42b5f838, 32'hc0dc5b49, 32'hc2829ec1, 32'hc29d3a47, 32'hc24ab51f, 32'h4299d8d2, 32'h407f1c1f, 32'hc26eafa9};
test_output[54] = '{32'h42b5f838};
test_index[54] = '{0};
test_input[440:447] = '{32'hbf74a5c3, 32'hc18c3981, 32'h4268fc6d, 32'h42452bb0, 32'h4283c18b, 32'hc2080e43, 32'h41e6d556, 32'h41c0d5dd};
test_output[55] = '{32'h4283c18b};
test_index[55] = '{4};
test_input[448:455] = '{32'hc2bcbed1, 32'h418f4638, 32'hc2a932ef, 32'h42b9050b, 32'h42a7da43, 32'hc2baa396, 32'h42565060, 32'h419ea698};
test_output[56] = '{32'h42b9050b};
test_index[56] = '{3};
test_input[456:463] = '{32'h422825c3, 32'h40cfc1b3, 32'hc2b55871, 32'h42a2d072, 32'h4258e9a5, 32'hc1f87ba5, 32'hc1ad18e0, 32'hc1686498};
test_output[57] = '{32'h42a2d072};
test_index[57] = '{3};
test_input[464:471] = '{32'hc1fb4b37, 32'hc28272df, 32'h42a991b1, 32'h428d831a, 32'hc21c49ab, 32'hc283c428, 32'h424efad1, 32'hc291a586};
test_output[58] = '{32'h42a991b1};
test_index[58] = '{2};
test_input[472:479] = '{32'hc2940b1c, 32'hc2997688, 32'h401c91d0, 32'hc298d2ac, 32'hc14777ff, 32'hc2864425, 32'hc1c02163, 32'h42878b53};
test_output[59] = '{32'h42878b53};
test_index[59] = '{7};
test_input[480:487] = '{32'h4083941b, 32'hc2aaa30d, 32'h417740b1, 32'hc2c11007, 32'h425c221a, 32'hc2a8235a, 32'hc28775f7, 32'hc2a6f8a6};
test_output[60] = '{32'h425c221a};
test_index[60] = '{4};
test_input[488:495] = '{32'h4262a72e, 32'hc17cad44, 32'h4003a59b, 32'h42ba8089, 32'hc2b9ae18, 32'h41defe1d, 32'h414d9a6b, 32'hc25f4a00};
test_output[61] = '{32'h42ba8089};
test_index[61] = '{3};
test_input[496:503] = '{32'hc264aa83, 32'h428f3707, 32'hc2616c9c, 32'h42ac00a8, 32'hc1f7abe1, 32'hc221e92c, 32'h416c059f, 32'hc29c91fb};
test_output[62] = '{32'h42ac00a8};
test_index[62] = '{3};
test_input[504:511] = '{32'hc2a9a7fe, 32'h4199cf1a, 32'hc28c8a7c, 32'hc201deff, 32'hc2740163, 32'h4196ecff, 32'h429e6dca, 32'hc085c9cd};
test_output[63] = '{32'h429e6dca};
test_index[63] = '{6};
test_input[512:519] = '{32'hc2a1eeb8, 32'h429316da, 32'h42b6fec6, 32'hc1c9cf65, 32'h42b02150, 32'hc2434d80, 32'hc2806b46, 32'hc2bc85e6};
test_output[64] = '{32'h42b6fec6};
test_index[64] = '{2};
test_input[520:527] = '{32'h4192dfba, 32'h418bb9d6, 32'hc07b9969, 32'hc10d75ed, 32'hc2c2bdb4, 32'hc1cc916e, 32'h4253dca5, 32'h422a5827};
test_output[65] = '{32'h4253dca5};
test_index[65] = '{6};
test_input[528:535] = '{32'h41810bd8, 32'h3fdf5d39, 32'hc233368f, 32'hc2ac58c4, 32'h415e3342, 32'hc269ee42, 32'h42a3d1e4, 32'h427158f2};
test_output[66] = '{32'h42a3d1e4};
test_index[66] = '{6};
test_input[536:543] = '{32'hc1f247a7, 32'h4182175f, 32'hc202d2e4, 32'h42a7205f, 32'h42bed7b1, 32'hc275a4a5, 32'hc26fb8ac, 32'hc2010478};
test_output[67] = '{32'h42bed7b1};
test_index[67] = '{4};
test_input[544:551] = '{32'h42bc37e7, 32'h4276332a, 32'h42727a96, 32'hc1bdc86b, 32'hc1eef8a1, 32'hbf910d7f, 32'hc28b4c7a, 32'hc2c7ff5a};
test_output[68] = '{32'h42bc37e7};
test_index[68] = '{0};
test_input[552:559] = '{32'hc2b1750b, 32'hc226f088, 32'h42b569a2, 32'h42bb198c, 32'hbef088ce, 32'h42b1ca42, 32'h41e6f54f, 32'h424e1fce};
test_output[69] = '{32'h42bb198c};
test_index[69] = '{3};
test_input[560:567] = '{32'hc2b3c08a, 32'h416c152d, 32'h428bd366, 32'h42c785e6, 32'h42310a00, 32'h41083db9, 32'h40026c30, 32'hc220722b};
test_output[70] = '{32'h42c785e6};
test_index[70] = '{3};
test_input[568:575] = '{32'hc2b3d7c9, 32'hc2518a82, 32'h400f8d59, 32'h425aac88, 32'hc0ce5264, 32'h42255dfc, 32'h41eb9190, 32'hc1fb15fa};
test_output[71] = '{32'h425aac88};
test_index[71] = '{3};
test_input[576:583] = '{32'hc2a7043f, 32'hc2b1a9d8, 32'hc28b2b88, 32'h424d020a, 32'hc26f8466, 32'h42371f31, 32'hc1f67e26, 32'hc28b5eb2};
test_output[72] = '{32'h424d020a};
test_index[72] = '{3};
test_input[584:591] = '{32'hc2910082, 32'hc275f14f, 32'hc2720260, 32'hc292aa00, 32'h4211a6a4, 32'hc2bb40cc, 32'hc19a4320, 32'h4221d741};
test_output[73] = '{32'h4221d741};
test_index[73] = '{7};
test_input[592:599] = '{32'h42a58440, 32'h41b89c07, 32'hc2272efe, 32'hc213af17, 32'hc20a81ca, 32'hc2b3ace8, 32'hc282d263, 32'hc13d0336};
test_output[74] = '{32'h42a58440};
test_index[74] = '{0};
test_input[600:607] = '{32'h42bb6e53, 32'hc290f01b, 32'h4249548d, 32'h428eb2b2, 32'h423aaf5c, 32'h427c83ad, 32'h40d88e01, 32'hc2b222de};
test_output[75] = '{32'h42bb6e53};
test_index[75] = '{0};
test_input[608:615] = '{32'h42468066, 32'h421d6d0c, 32'hc1ef3fa4, 32'hc2beadf8, 32'h420686c2, 32'hc240c044, 32'h41f584a5, 32'h40ed18be};
test_output[76] = '{32'h42468066};
test_index[76] = '{0};
test_input[616:623] = '{32'hc29cfb76, 32'hc24bff4b, 32'h4281ac29, 32'hc2c11e60, 32'h42a3d429, 32'h42c01b05, 32'hc01a1164, 32'hbf9d3fb5};
test_output[77] = '{32'h42c01b05};
test_index[77] = '{5};
test_input[624:631] = '{32'h424255b0, 32'hc281f4ff, 32'h42540e48, 32'h41d90ebc, 32'h429b8852, 32'hc2b4db7f, 32'hc23dd3ca, 32'h42a76198};
test_output[78] = '{32'h42a76198};
test_index[78] = '{7};
test_input[632:639] = '{32'hc24b11dd, 32'hc2a96d0e, 32'hc21d575b, 32'hc2bbb426, 32'h41c1c5db, 32'hc1ee0751, 32'hc1ffadb9, 32'hc0f4ad1b};
test_output[79] = '{32'h41c1c5db};
test_index[79] = '{4};
test_input[640:647] = '{32'hc23017e1, 32'hc2833a88, 32'hc2a87f64, 32'hc2ad3f7b, 32'h41a89bbf, 32'hc22cf363, 32'hc2a5ef7c, 32'h41c1ac8a};
test_output[80] = '{32'h41c1ac8a};
test_index[80] = '{7};
test_input[648:655] = '{32'hc2b01e4b, 32'hc2c02170, 32'hc2ad6835, 32'hc1326860, 32'h3fb4e0f9, 32'h42561dec, 32'hc24840ad, 32'hc1efc1b2};
test_output[81] = '{32'h42561dec};
test_index[81] = '{5};
test_input[656:663] = '{32'hc09efab0, 32'h42b36c4e, 32'hc0a7d84e, 32'h420bb9c4, 32'hc04be7ef, 32'hc1dca01d, 32'h4208076b, 32'h41a880a4};
test_output[82] = '{32'h42b36c4e};
test_index[82] = '{1};
test_input[664:671] = '{32'h421daba9, 32'hbcdc9aad, 32'h42c78f8a, 32'h4299db75, 32'h42c0531e, 32'h411d29bb, 32'h42a9102e, 32'h41ce768e};
test_output[83] = '{32'h42c78f8a};
test_index[83] = '{2};
test_input[672:679] = '{32'hc2b3285b, 32'hc291f110, 32'hc12d9344, 32'hc0cf05ef, 32'hc22b5552, 32'h3ee4be52, 32'h42a79247, 32'hc28a80b3};
test_output[84] = '{32'h42a79247};
test_index[84] = '{6};
test_input[680:687] = '{32'h42b44c80, 32'hc1bca00d, 32'hc22752be, 32'h41225922, 32'hc2c1dcb1, 32'hc1fa3471, 32'hc292c3df, 32'h418db84a};
test_output[85] = '{32'h42b44c80};
test_index[85] = '{0};
test_input[688:695] = '{32'h40a3af07, 32'hc2008d3a, 32'hc26c88de, 32'hc25e4109, 32'h42be8d57, 32'h42bbb6af, 32'h40bd327a, 32'hc2a0ec18};
test_output[86] = '{32'h42be8d57};
test_index[86] = '{4};
test_input[696:703] = '{32'hc2b198fc, 32'h424fa934, 32'h421e86bc, 32'h4280164a, 32'hc2866add, 32'h423e1028, 32'hc2556104, 32'hc2178286};
test_output[87] = '{32'h4280164a};
test_index[87] = '{3};
test_input[704:711] = '{32'hc29005e6, 32'hc2769499, 32'h42168f40, 32'h42b33754, 32'h422dd93c, 32'h4295424b, 32'h40afb0a9, 32'hc1c32a8d};
test_output[88] = '{32'h42b33754};
test_index[88] = '{3};
test_input[712:719] = '{32'hc28877f6, 32'hc253140a, 32'h4233ccb2, 32'hc2397306, 32'h3e0d32a2, 32'hbf137bf7, 32'h421ebcd9, 32'h3fb5966c};
test_output[89] = '{32'h4233ccb2};
test_index[89] = '{2};
test_input[720:727] = '{32'h42133ac1, 32'hc2145656, 32'h42c746fc, 32'hc2a5568b, 32'hc2b9b1d7, 32'h42b5f8c6, 32'hc2928f62, 32'hc25ea78c};
test_output[90] = '{32'h42c746fc};
test_index[90] = '{2};
test_input[728:735] = '{32'hc2843261, 32'h41ce4582, 32'h429bf8c6, 32'hc215ae9a, 32'h41f48469, 32'h3e914405, 32'h42a0efae, 32'h42825475};
test_output[91] = '{32'h42a0efae};
test_index[91] = '{6};
test_input[736:743] = '{32'h42a02473, 32'hc2abffaa, 32'h426b083f, 32'h423184d8, 32'h42b052bf, 32'h417cd9a2, 32'hc2383bc3, 32'hc12d43d7};
test_output[92] = '{32'h42b052bf};
test_index[92] = '{4};
test_input[744:751] = '{32'hc021354f, 32'hc246532e, 32'h42c5a0c0, 32'h42a9763b, 32'hc1997cab, 32'hc1e9e545, 32'h42242d55, 32'h41e9afe8};
test_output[93] = '{32'h42c5a0c0};
test_index[93] = '{2};
test_input[752:759] = '{32'h415d54e1, 32'hc2557d6b, 32'h42b70e57, 32'h42916f56, 32'hc2183d0d, 32'hc2a2d717, 32'h429f2704, 32'h427b2520};
test_output[94] = '{32'h42b70e57};
test_index[94] = '{2};
test_input[760:767] = '{32'h4291440a, 32'h427508b6, 32'h426a1e64, 32'h41ab73a0, 32'h4217949e, 32'hc24d7abc, 32'hc29a6b86, 32'hc1e2b9f0};
test_output[95] = '{32'h4291440a};
test_index[95] = '{0};
test_input[768:775] = '{32'hc2baa4b2, 32'h4110e2ef, 32'hc24cbbbe, 32'h421dbbc8, 32'h42433b26, 32'hc2a6f2cf, 32'hc286dee6, 32'h4240d083};
test_output[96] = '{32'h42433b26};
test_index[96] = '{4};
test_input[776:783] = '{32'hc235dea1, 32'h4121c702, 32'hc20b136c, 32'hc27189b9, 32'hc20a57f1, 32'hc2c0f710, 32'hc2aab357, 32'h42743376};
test_output[97] = '{32'h42743376};
test_index[97] = '{7};
test_input[784:791] = '{32'h42bd0b6f, 32'h40b88287, 32'h421b256a, 32'hc274629f, 32'h42c44a1f, 32'hc069987f, 32'h41911aac, 32'h40f3fb87};
test_output[98] = '{32'h42c44a1f};
test_index[98] = '{4};
test_input[792:799] = '{32'hc1c2e017, 32'h41fbd884, 32'hc0a3e14d, 32'hc288913e, 32'h423f9086, 32'hc2521d31, 32'h41a8b74b, 32'hc0c7017f};
test_output[99] = '{32'h423f9086};
test_index[99] = '{4};
test_input[800:807] = '{32'hc12a73a8, 32'h41e9bab8, 32'h4181f2d4, 32'hc25c84d1, 32'h4271c7d4, 32'h428747a8, 32'hc2ad42fa, 32'hc2a7a382};
test_output[100] = '{32'h428747a8};
test_index[100] = '{5};
test_input[808:815] = '{32'h42913938, 32'h42834b18, 32'hc2803e24, 32'hc226d38e, 32'h417d337a, 32'h429a420b, 32'h4291e0d6, 32'hc1879a1e};
test_output[101] = '{32'h429a420b};
test_index[101] = '{5};
test_input[816:823] = '{32'hc240823c, 32'hc28dd9e0, 32'hc2972759, 32'hc14594ad, 32'h426ba751, 32'hc27451f7, 32'hc2c09660, 32'hc1a55faf};
test_output[102] = '{32'h426ba751};
test_index[102] = '{4};
test_input[824:831] = '{32'h4224df8d, 32'h42505931, 32'h42292116, 32'h42818f06, 32'h42959046, 32'h42a0a70d, 32'hc0f1cb14, 32'hc29786a3};
test_output[103] = '{32'h42a0a70d};
test_index[103] = '{5};
test_input[832:839] = '{32'h4286f45a, 32'hc20385ee, 32'h40b587d4, 32'hc1cfbd31, 32'hc2509595, 32'h41bc573e, 32'hc1a03fb1, 32'hc2597adb};
test_output[104] = '{32'h4286f45a};
test_index[104] = '{0};
test_input[840:847] = '{32'hc29c3038, 32'h42a06d85, 32'h422b2e51, 32'hc2811e47, 32'hc241d7c3, 32'hc2b84aeb, 32'hc2ad4846, 32'h42a7aaa4};
test_output[105] = '{32'h42a7aaa4};
test_index[105] = '{7};
test_input[848:855] = '{32'hc2071660, 32'hc28c8765, 32'h42b85ebe, 32'h4249d36d, 32'hc2b820db, 32'hc15a786e, 32'hc251a32c, 32'h419af3d7};
test_output[106] = '{32'h42b85ebe};
test_index[106] = '{2};
test_input[856:863] = '{32'hc2ad3bf3, 32'hc253783f, 32'h42b82300, 32'h42bf80bc, 32'hc2a0acbd, 32'h42641151, 32'hc28cd5e0, 32'h4254d352};
test_output[107] = '{32'h42bf80bc};
test_index[107] = '{3};
test_input[864:871] = '{32'hc1ca0e11, 32'hc050bdef, 32'h42b4162f, 32'h4207449b, 32'hc29eeffa, 32'h42b150e0, 32'h4260f487, 32'hc2bee018};
test_output[108] = '{32'h42b4162f};
test_index[108] = '{2};
test_input[872:879] = '{32'hc1712061, 32'hc2c09c52, 32'h42b2793a, 32'h429c03cf, 32'h4197f37b, 32'hc287246d, 32'hc2b32d42, 32'h421fccab};
test_output[109] = '{32'h42b2793a};
test_index[109] = '{2};
test_input[880:887] = '{32'h421dd0b0, 32'hc29484d5, 32'h41c2fe9b, 32'h41378bcb, 32'hc1ead5ac, 32'h4244f7a0, 32'hbfcddd1d, 32'h4236b07a};
test_output[110] = '{32'h4244f7a0};
test_index[110] = '{5};
test_input[888:895] = '{32'h41d0742a, 32'h4261e1aa, 32'hc10827b3, 32'hc2691278, 32'h416d88c1, 32'hc2a96d65, 32'h4202f165, 32'h42c5cd25};
test_output[111] = '{32'h42c5cd25};
test_index[111] = '{7};
test_input[896:903] = '{32'hc01b66b5, 32'hc1fd18cb, 32'hc292580a, 32'hc29ccb6a, 32'hc23bcbf4, 32'h426939e8, 32'hc2c3ccd4, 32'h414edd40};
test_output[112] = '{32'h426939e8};
test_index[112] = '{5};
test_input[904:911] = '{32'h42998c7b, 32'h411c83e1, 32'h4144fab4, 32'hc2c3c398, 32'hc2c136b5, 32'h41762e51, 32'hc2a5f833, 32'h42406e94};
test_output[113] = '{32'h42998c7b};
test_index[113] = '{0};
test_input[912:919] = '{32'hc092c404, 32'hc27e447f, 32'hc2aae00a, 32'h42045227, 32'hc203c052, 32'h429a845e, 32'h42886679, 32'h427d62bd};
test_output[114] = '{32'h429a845e};
test_index[114] = '{5};
test_input[920:927] = '{32'hc29c5138, 32'hc2abfffc, 32'hc0dd7861, 32'hc1e5564b, 32'hc1cc4bc7, 32'hc2ad0db0, 32'h42a45d0d, 32'hc263d1c0};
test_output[115] = '{32'h42a45d0d};
test_index[115] = '{6};
test_input[928:935] = '{32'h42828488, 32'h418cb407, 32'hc285e3eb, 32'h42bc40d9, 32'hc2abd679, 32'hc29f14ee, 32'h426c7dac, 32'h4208a7e7};
test_output[116] = '{32'h42bc40d9};
test_index[116] = '{3};
test_input[936:943] = '{32'h429f82a2, 32'h41c16425, 32'hc1813376, 32'hc2380b5d, 32'hc2bb585c, 32'hc2672dbb, 32'h41815fe8, 32'hc2960541};
test_output[117] = '{32'h429f82a2};
test_index[117] = '{0};
test_input[944:951] = '{32'h423afcb4, 32'hbfb01c06, 32'h4222607a, 32'hc1a87fe0, 32'hc266ab1d, 32'hc1868fad, 32'h428f28e0, 32'h427dbbdc};
test_output[118] = '{32'h428f28e0};
test_index[118] = '{6};
test_input[952:959] = '{32'h42c377de, 32'hc24f3da1, 32'h4229bdb6, 32'h428a0376, 32'h408f913a, 32'hc1c93424, 32'h4282106b, 32'hc25ec11b};
test_output[119] = '{32'h42c377de};
test_index[119] = '{0};
test_input[960:967] = '{32'hc2b82b50, 32'h4133612a, 32'hc28c2dca, 32'hc214d800, 32'h42a7e671, 32'hc27aaf3b, 32'hc2ace1d5, 32'hc209b15f};
test_output[120] = '{32'h42a7e671};
test_index[120] = '{4};
test_input[968:975] = '{32'h42523165, 32'hc2bff94a, 32'hc19d0714, 32'h4289937b, 32'hc28c50a9, 32'h41dff8b2, 32'hc27820de, 32'h4089ed7a};
test_output[121] = '{32'h4289937b};
test_index[121] = '{3};
test_input[976:983] = '{32'h429163e3, 32'h42865516, 32'hc1ce8302, 32'h4273a8b0, 32'hc247bfcb, 32'h423c39b2, 32'h4281f187, 32'h41662849};
test_output[122] = '{32'h429163e3};
test_index[122] = '{0};
test_input[984:991] = '{32'h4256326a, 32'h41242fcc, 32'h403348f0, 32'hc1eb69f4, 32'h424e104e, 32'hc25ca9fb, 32'hc2c781ff, 32'hc2443752};
test_output[123] = '{32'h4256326a};
test_index[123] = '{0};
test_input[992:999] = '{32'h4296dd61, 32'h428a864e, 32'h417d42ed, 32'hc1f3f2be, 32'h4113b1e5, 32'hc263dc62, 32'hc1638116, 32'h3fab8bf6};
test_output[124] = '{32'h4296dd61};
test_index[124] = '{0};
test_input[1000:1007] = '{32'hc12fddc5, 32'h41b1fbb3, 32'hc206731c, 32'hc2a0d32e, 32'h4290aa33, 32'hc28d7de7, 32'h424b3424, 32'hc0941474};
test_output[125] = '{32'h4290aa33};
test_index[125] = '{4};
test_input[1008:1015] = '{32'h42a62877, 32'h421b170f, 32'hc25a5dad, 32'h418a6b92, 32'h429b7b15, 32'h42a0d9b9, 32'h41c4254f, 32'hc291e0d3};
test_output[126] = '{32'h42a62877};
test_index[126] = '{0};
test_input[1016:1023] = '{32'h42871a74, 32'hc2895103, 32'hc27f6c6f, 32'h4249d4e9, 32'hc2359639, 32'hc0d758e1, 32'h40b1d924, 32'h421477f0};
test_output[127] = '{32'h42871a74};
test_index[127] = '{0};
test_input[1024:1031] = '{32'h42ae78ed, 32'hc1a0a534, 32'h4184fec4, 32'h427699a9, 32'hc15fb650, 32'hc2ba575a, 32'hc034236c, 32'hc18eb866};
test_output[128] = '{32'h42ae78ed};
test_index[128] = '{0};
test_input[1032:1039] = '{32'hc2b5f9fe, 32'h42446d57, 32'hc2929893, 32'hc26118ea, 32'hc2c57cfc, 32'h41d76995, 32'h424453fc, 32'h4284ac49};
test_output[129] = '{32'h4284ac49};
test_index[129] = '{7};
test_input[1040:1047] = '{32'h42714930, 32'h4287566a, 32'h422143f4, 32'h4236be46, 32'hc2268dc0, 32'h41da2645, 32'hc2756450, 32'h4297e2b5};
test_output[130] = '{32'h4297e2b5};
test_index[130] = '{7};
test_input[1048:1055] = '{32'hc22b6ab7, 32'h42bb2433, 32'hc290cb0a, 32'hc1cf8b7f, 32'hc254786d, 32'hc2affbed, 32'h422003e0, 32'h42220359};
test_output[131] = '{32'h42bb2433};
test_index[131] = '{1};
test_input[1056:1063] = '{32'h422a6125, 32'hc1ffe7d6, 32'h4250097a, 32'hc1812333, 32'h428bbc31, 32'hc1fb5958, 32'h42bbd043, 32'hc27777a5};
test_output[132] = '{32'h42bbd043};
test_index[132] = '{6};
test_input[1064:1071] = '{32'hc20c23af, 32'h4231bf73, 32'hc21128ee, 32'h41dc4b58, 32'h429bc2f7, 32'hc2027e77, 32'h429eda8e, 32'hc1e57a2c};
test_output[133] = '{32'h429eda8e};
test_index[133] = '{6};
test_input[1072:1079] = '{32'h41b3d892, 32'hc24419d8, 32'hc1c70fa9, 32'hc290644f, 32'hc13fcc78, 32'hc2264b3c, 32'hc22971b4, 32'h422bab5d};
test_output[134] = '{32'h422bab5d};
test_index[134] = '{7};
test_input[1080:1087] = '{32'hc2c2378a, 32'hc24125bf, 32'h41e151f4, 32'hc29990b7, 32'h428f85d4, 32'hc22d7659, 32'h410ac4ed, 32'h41f9cda2};
test_output[135] = '{32'h428f85d4};
test_index[135] = '{4};
test_input[1088:1095] = '{32'h41d5e1d9, 32'hc294ed51, 32'hc296618b, 32'h42acbac8, 32'h42121f67, 32'h4243e9f7, 32'hc1463084, 32'h40cdb417};
test_output[136] = '{32'h42acbac8};
test_index[136] = '{3};
test_input[1096:1103] = '{32'h423e4c9c, 32'h42b94991, 32'hc29514e8, 32'hc17b572b, 32'h412b8849, 32'h4226e787, 32'h40c73236, 32'hc1346420};
test_output[137] = '{32'h42b94991};
test_index[137] = '{1};
test_input[1104:1111] = '{32'h41dcc6f3, 32'h420e17b6, 32'hc1abc201, 32'hc2026761, 32'hc1e23dbe, 32'hc2c708f7, 32'h428e13ed, 32'h4147298d};
test_output[138] = '{32'h428e13ed};
test_index[138] = '{6};
test_input[1112:1119] = '{32'h42a94de0, 32'h41d2739b, 32'hc262ad2d, 32'hc1dbf78b, 32'h41a0d7ae, 32'h3fd2dc5d, 32'h42bcf13b, 32'h42c42b8c};
test_output[139] = '{32'h42c42b8c};
test_index[139] = '{7};
test_input[1120:1127] = '{32'hc29fadb4, 32'hc21b8bac, 32'h42800b91, 32'hc103eecd, 32'hc283ed28, 32'hc284005c, 32'h42a707da, 32'h429d4418};
test_output[140] = '{32'h42a707da};
test_index[140] = '{6};
test_input[1128:1135] = '{32'h4297be0a, 32'hc2a68fda, 32'h41d8804b, 32'hc2170998, 32'h4206f0b5, 32'hc23910cc, 32'hc248ee41, 32'hc2ad4595};
test_output[141] = '{32'h4297be0a};
test_index[141] = '{0};
test_input[1136:1143] = '{32'h41494c95, 32'h41cfcb65, 32'h42c147f2, 32'hc0afeaf0, 32'hc20eac07, 32'hc185fdc8, 32'hc13f830a, 32'hbf1528ff};
test_output[142] = '{32'h42c147f2};
test_index[142] = '{2};
test_input[1144:1151] = '{32'h4143087c, 32'h41fa493e, 32'h42766471, 32'h4253555f, 32'h42312a44, 32'hc242e1c1, 32'hc2a473a0, 32'hc216e852};
test_output[143] = '{32'h42766471};
test_index[143] = '{2};
test_input[1152:1159] = '{32'hc1637401, 32'h429f0815, 32'hc284c467, 32'hc225630b, 32'hc21db9f8, 32'h413b7507, 32'hc21ace43, 32'hc18c2de7};
test_output[144] = '{32'h429f0815};
test_index[144] = '{1};
test_input[1160:1167] = '{32'hc237d82b, 32'h426632e9, 32'hc28b44af, 32'hc2b45d26, 32'h42aa1e3b, 32'h422f7aec, 32'h40c827c5, 32'hc257f0cf};
test_output[145] = '{32'h42aa1e3b};
test_index[145] = '{4};
test_input[1168:1175] = '{32'h4048f04b, 32'h416d79e8, 32'hc189eac5, 32'hc17a2914, 32'h4233c416, 32'hc2bf54c5, 32'h3f1cf0d1, 32'hc00ae045};
test_output[146] = '{32'h4233c416};
test_index[146] = '{4};
test_input[1176:1183] = '{32'h41922116, 32'h42b2b1f2, 32'hc1e9d462, 32'hc1a52b40, 32'hc28d8b27, 32'h41d9487d, 32'h4219f18c, 32'h4201b165};
test_output[147] = '{32'h42b2b1f2};
test_index[147] = '{1};
test_input[1184:1191] = '{32'h42afbda9, 32'hc2a4d8b9, 32'hc10a0c48, 32'hc284ad4a, 32'h41a3dc61, 32'h414d17c0, 32'hc1f427e1, 32'h422cc166};
test_output[148] = '{32'h42afbda9};
test_index[148] = '{0};
test_input[1192:1199] = '{32'hc12a1f7b, 32'hc29eb4d8, 32'h42022827, 32'h4266ee28, 32'hc141e986, 32'hc2951d05, 32'hc0957340, 32'hc2b7b867};
test_output[149] = '{32'h4266ee28};
test_index[149] = '{3};
test_input[1200:1207] = '{32'h429e6131, 32'hc298f814, 32'hc2a72aca, 32'h42b6175e, 32'hc2afa34b, 32'h4136baad, 32'hc2405552, 32'h42a37694};
test_output[150] = '{32'h42b6175e};
test_index[150] = '{3};
test_input[1208:1215] = '{32'h4298dbdb, 32'hc17b89fc, 32'hc2a54234, 32'hc2b8f5ed, 32'hc2c7b4a3, 32'h427e061f, 32'hc1b4d311, 32'h41a8afd4};
test_output[151] = '{32'h4298dbdb};
test_index[151] = '{0};
test_input[1216:1223] = '{32'h40aba6b9, 32'h424038d7, 32'h428bde76, 32'hc28dfa88, 32'h42b412f6, 32'hc1121545, 32'hc1a5b956, 32'h429f299d};
test_output[152] = '{32'h42b412f6};
test_index[152] = '{4};
test_input[1224:1231] = '{32'h422cabf3, 32'h429a08ab, 32'hc2616e4b, 32'hc298add3, 32'hc2c1e8c1, 32'h41ba03ea, 32'hc22293e7, 32'h4204d49c};
test_output[153] = '{32'h429a08ab};
test_index[153] = '{1};
test_input[1232:1239] = '{32'hc2ae349d, 32'hc21ebb01, 32'h41c90e80, 32'hc2bf39ed, 32'hc218bf5a, 32'h40b0a456, 32'h4240eadc, 32'h41f408cb};
test_output[154] = '{32'h4240eadc};
test_index[154] = '{6};
test_input[1240:1247] = '{32'hc284a847, 32'hc2360b39, 32'hc1921f65, 32'hc25806fa, 32'hc23314a6, 32'h403111c9, 32'h429e7292, 32'hc291bb05};
test_output[155] = '{32'h429e7292};
test_index[155] = '{6};
test_input[1248:1255] = '{32'hc12dc1a6, 32'h42ade992, 32'h425377e6, 32'h42647fa7, 32'hc26cf8f9, 32'hc16e2499, 32'h42b44d87, 32'h416e5534};
test_output[156] = '{32'h42b44d87};
test_index[156] = '{6};
test_input[1256:1263] = '{32'h4239817e, 32'h4268185e, 32'h41a81a39, 32'h42527686, 32'h42550cf4, 32'h4290493f, 32'hc1e35b95, 32'hc2c32c65};
test_output[157] = '{32'h4290493f};
test_index[157] = '{5};
test_input[1264:1271] = '{32'hc26db27b, 32'hc1c83c30, 32'hc196975d, 32'hc20e20f9, 32'h428e707c, 32'hc29c3275, 32'hbfef6803, 32'h413f765e};
test_output[158] = '{32'h428e707c};
test_index[158] = '{4};
test_input[1272:1279] = '{32'h42b7030a, 32'hc209aad2, 32'hc202d7f4, 32'h419bc795, 32'h41f0a61b, 32'hc2069f22, 32'hc2a6ccbf, 32'hc1bb2886};
test_output[159] = '{32'h42b7030a};
test_index[159] = '{0};
test_input[1280:1287] = '{32'h428c1b52, 32'h420e01d0, 32'h41047669, 32'h423b97d6, 32'h42ac300c, 32'h42acf996, 32'h428c8726, 32'h42a1cd56};
test_output[160] = '{32'h42acf996};
test_index[160] = '{5};
test_input[1288:1295] = '{32'hc1a758fc, 32'h42711bd4, 32'h42b9ec0f, 32'h422e0db3, 32'h4294ded0, 32'h42bd8710, 32'h42ba5f95, 32'h4268650c};
test_output[161] = '{32'h42bd8710};
test_index[161] = '{5};
test_input[1296:1303] = '{32'h4170ab68, 32'hc10d340d, 32'h4196a887, 32'hc1dcc2ec, 32'h425f5049, 32'h3fd12729, 32'hc2a36554, 32'h406c2500};
test_output[162] = '{32'h425f5049};
test_index[162] = '{4};
test_input[1304:1311] = '{32'hc202cd9e, 32'hc2123ba4, 32'hc27f425a, 32'h411972fc, 32'hc25266db, 32'hc299dd9b, 32'hc272d9db, 32'h42504494};
test_output[163] = '{32'h42504494};
test_index[163] = '{7};
test_input[1312:1319] = '{32'h41a8805b, 32'h40db9f31, 32'h422b8f95, 32'h42b5a60e, 32'h41fc7634, 32'hc0925a90, 32'hc22fcd74, 32'h42a38878};
test_output[164] = '{32'h42b5a60e};
test_index[164] = '{3};
test_input[1320:1327] = '{32'h3ed7fc0a, 32'h42984c33, 32'h41b03437, 32'h42174073, 32'h40bfbb0c, 32'hc2818b3a, 32'hc26516ca, 32'hc2ae0b50};
test_output[165] = '{32'h42984c33};
test_index[165] = '{1};
test_input[1328:1335] = '{32'h4107f3f9, 32'hc157f766, 32'h42b3c0db, 32'hc25829fe, 32'hc2850ea2, 32'hc115762c, 32'hc297e555, 32'h427d3bea};
test_output[166] = '{32'h42b3c0db};
test_index[166] = '{2};
test_input[1336:1343] = '{32'hc124f047, 32'hc18ce0aa, 32'h42ad4f02, 32'h41cdc227, 32'h42b6976a, 32'h3f989ce7, 32'hc0aeeca4, 32'hc2485562};
test_output[167] = '{32'h42b6976a};
test_index[167] = '{4};
test_input[1344:1351] = '{32'hc0a5760a, 32'hc11bc2a2, 32'hc284eabc, 32'hc2075709, 32'h429a9850, 32'h42c3a85f, 32'hc281828f, 32'h42322547};
test_output[168] = '{32'h42c3a85f};
test_index[168] = '{5};
test_input[1352:1359] = '{32'hc15cac79, 32'h42c6f093, 32'h4262e05b, 32'hc2a16c86, 32'h42111f3a, 32'h4205c334, 32'h41d0640e, 32'hc21522cd};
test_output[169] = '{32'h42c6f093};
test_index[169] = '{1};
test_input[1360:1367] = '{32'h42b95e84, 32'h42397b21, 32'h429d1d99, 32'h41b20b4d, 32'hc28e4404, 32'hc1f1767f, 32'h41ddae27, 32'h4296fde9};
test_output[170] = '{32'h42b95e84};
test_index[170] = '{0};
test_input[1368:1375] = '{32'hc2607864, 32'h428a498d, 32'h42b5a6e6, 32'h42368cf2, 32'hc29dc647, 32'h4150f465, 32'h427040b3, 32'h40ebffb9};
test_output[171] = '{32'h42b5a6e6};
test_index[171] = '{2};
test_input[1376:1383] = '{32'h42c2080f, 32'h4168a38d, 32'h42699540, 32'h4230ac25, 32'hc2a65144, 32'h42b2061f, 32'h420e896e, 32'hc2b75522};
test_output[172] = '{32'h42c2080f};
test_index[172] = '{0};
test_input[1384:1391] = '{32'h42aaa407, 32'h42314140, 32'h420199ba, 32'h419eece9, 32'hc28ad8e8, 32'h427fb2e8, 32'hc2bf2cd0, 32'hc21c7cb1};
test_output[173] = '{32'h42aaa407};
test_index[173] = '{0};
test_input[1392:1399] = '{32'h4244461b, 32'h420a7d57, 32'hc2bc031c, 32'hc29690b4, 32'h41e2f796, 32'hc21614f7, 32'h4274b6e6, 32'hc2061ba8};
test_output[174] = '{32'h4274b6e6};
test_index[174] = '{6};
test_input[1400:1407] = '{32'hc2bccf21, 32'h3f993f67, 32'hc1bed259, 32'h4125881d, 32'hc1c53f9e, 32'h41867266, 32'hc2896baf, 32'h425fbdcf};
test_output[175] = '{32'h425fbdcf};
test_index[175] = '{7};
test_input[1408:1415] = '{32'h42b7d741, 32'h427fd8c9, 32'h420e8d23, 32'h41ff67e2, 32'hc2a6fdc4, 32'hc22128cf, 32'hc20e134d, 32'h42b5f860};
test_output[176] = '{32'h42b7d741};
test_index[176] = '{0};
test_input[1416:1423] = '{32'h428a2d6f, 32'h41decb2a, 32'h424aadf9, 32'h42b8bf84, 32'hc287300e, 32'hc28bdae1, 32'hc281efbc, 32'hc2a43719};
test_output[177] = '{32'h42b8bf84};
test_index[177] = '{3};
test_input[1424:1431] = '{32'h4297fc60, 32'h42b88517, 32'h41df78a7, 32'hc0b1987a, 32'h42420230, 32'hc185d827, 32'h41b68c02, 32'hc211a941};
test_output[178] = '{32'h42b88517};
test_index[178] = '{1};
test_input[1432:1439] = '{32'h42abcdb8, 32'hc2b22662, 32'h4295f68e, 32'hc1ca50ba, 32'hc115d431, 32'hc22a4f3f, 32'hc2390d88, 32'h425c2e38};
test_output[179] = '{32'h42abcdb8};
test_index[179] = '{0};
test_input[1440:1447] = '{32'h429940ae, 32'h42bf4bb1, 32'h418c71c4, 32'hc23c7648, 32'h424e49af, 32'h42ba49bb, 32'hc1e0fbd3, 32'hc2426208};
test_output[180] = '{32'h42bf4bb1};
test_index[180] = '{1};
test_input[1448:1455] = '{32'hc247c2e3, 32'h425d36bb, 32'h42c45a6c, 32'h4299c568, 32'hc24cbac6, 32'hc2a9e9c3, 32'h41904cb1, 32'hc14cb206};
test_output[181] = '{32'h42c45a6c};
test_index[181] = '{2};
test_input[1456:1463] = '{32'hc23ad929, 32'hc21f278e, 32'h42bd5a13, 32'h42a9cb7e, 32'h42888e6e, 32'hc20de797, 32'h42a8dee9, 32'hc1ac9ecb};
test_output[182] = '{32'h42bd5a13};
test_index[182] = '{2};
test_input[1464:1471] = '{32'hc2790a4b, 32'hc15eaeff, 32'hc1f1dd00, 32'hc1140c24, 32'h42b792f6, 32'hc292a0f5, 32'hc2a83bdf, 32'h418eae45};
test_output[183] = '{32'h42b792f6};
test_index[183] = '{4};
test_input[1472:1479] = '{32'hc1cf8f4b, 32'hc109edb1, 32'h42a51172, 32'h423a6934, 32'hc2a602ab, 32'hc2944532, 32'h42262d35, 32'h4201215d};
test_output[184] = '{32'h42a51172};
test_index[184] = '{2};
test_input[1480:1487] = '{32'hc2b07d9f, 32'hc201581f, 32'hc2a3a55b, 32'h424e50ff, 32'h41164e19, 32'hc237e190, 32'hc2ab8b3d, 32'h4206a0a8};
test_output[185] = '{32'h424e50ff};
test_index[185] = '{3};
test_input[1488:1495] = '{32'h41fa505c, 32'hc1c67985, 32'h4251e003, 32'hc25c5a42, 32'h4081e580, 32'h4284778e, 32'h41eb368e, 32'hc2c14929};
test_output[186] = '{32'h4284778e};
test_index[186] = '{5};
test_input[1496:1503] = '{32'hc1daa09c, 32'hc29e884b, 32'hc2585e75, 32'h4292cd0d, 32'h415faa6b, 32'h42ab64ba, 32'hc2805b0b, 32'h41620266};
test_output[187] = '{32'h42ab64ba};
test_index[187] = '{5};
test_input[1504:1511] = '{32'h40bb309c, 32'h423b9c71, 32'hc2b18a6c, 32'h41069bfd, 32'h424b5e10, 32'hc060fe6f, 32'h42ad02ae, 32'h42a319b8};
test_output[188] = '{32'h42ad02ae};
test_index[188] = '{6};
test_input[1512:1519] = '{32'hc2b777f3, 32'hc2b3cc17, 32'h421165e3, 32'h418ef7f5, 32'h42c1c70e, 32'h422ffefb, 32'h410f65a2, 32'hc249fc59};
test_output[189] = '{32'h42c1c70e};
test_index[189] = '{4};
test_input[1520:1527] = '{32'h426a7269, 32'hc28fd057, 32'hc16ae1da, 32'hc2431fa7, 32'h42aa86a7, 32'hc2c3dcdf, 32'hc1e0aa68, 32'h417aacfe};
test_output[190] = '{32'h42aa86a7};
test_index[190] = '{4};
test_input[1528:1535] = '{32'h3f57262a, 32'h423d6abe, 32'h418a0b54, 32'h424a7b4d, 32'hc2b1ba7d, 32'hc218c52c, 32'h408cd0c2, 32'hc24ff5ba};
test_output[191] = '{32'h424a7b4d};
test_index[191] = '{3};
test_input[1536:1543] = '{32'h420e224e, 32'h42b424a0, 32'h42c61b16, 32'hc2889c42, 32'h4167711e, 32'h42b77c3a, 32'hc16c3e58, 32'h42bbf8f0};
test_output[192] = '{32'h42c61b16};
test_index[192] = '{2};
test_input[1544:1551] = '{32'h41f54103, 32'h4172e4e2, 32'hc24a8a4f, 32'hc2799667, 32'hc26b4daa, 32'h428d704b, 32'hc09f5564, 32'hc2471923};
test_output[193] = '{32'h428d704b};
test_index[193] = '{5};
test_input[1552:1559] = '{32'h41a7201d, 32'h4297feda, 32'h41c325a6, 32'hc0eb8e52, 32'hc2671a37, 32'hc293c5d9, 32'h42b74fd3, 32'hc29ded5c};
test_output[194] = '{32'h42b74fd3};
test_index[194] = '{6};
test_input[1560:1567] = '{32'h4286a773, 32'hc1dd44a8, 32'hc2bca815, 32'hc1c64561, 32'hc1a39c1d, 32'h42c2cbd0, 32'h4093caf3, 32'h41b5b612};
test_output[195] = '{32'h42c2cbd0};
test_index[195] = '{5};
test_input[1568:1575] = '{32'h41748d64, 32'hc216645a, 32'hc2c1afca, 32'hc276c6d1, 32'h42c12f03, 32'h42387ec9, 32'h428271bb, 32'hc25256e0};
test_output[196] = '{32'h42c12f03};
test_index[196] = '{4};
test_input[1576:1583] = '{32'hc26c78a1, 32'h42a47fa6, 32'hc0c89b3a, 32'h42c43843, 32'h426840f2, 32'h4213762a, 32'h42a552be, 32'hc206ba11};
test_output[197] = '{32'h42c43843};
test_index[197] = '{3};
test_input[1584:1591] = '{32'h42368b13, 32'h421740cf, 32'h41c7e5b3, 32'h42b569db, 32'h42b0df2d, 32'h42648307, 32'h42b15eeb, 32'hc261948e};
test_output[198] = '{32'h42b569db};
test_index[198] = '{3};
test_input[1592:1599] = '{32'hc210d653, 32'h42c2e7d2, 32'hc2ac9c50, 32'hc281c294, 32'hc0c614c1, 32'h41d4fd99, 32'h4111be14, 32'h424c4733};
test_output[199] = '{32'h42c2e7d2};
test_index[199] = '{1};
test_input[1600:1607] = '{32'hc20aacc6, 32'hc0ce41a1, 32'hc2956192, 32'hc1dce6df, 32'hc21b4046, 32'h42bdf1b5, 32'hc1b876f0, 32'h4206fa50};
test_output[200] = '{32'h42bdf1b5};
test_index[200] = '{5};
test_input[1608:1615] = '{32'hc1a1b0f1, 32'hc240ec0a, 32'h429d3163, 32'h42beeedf, 32'h412a974c, 32'hbf8b511e, 32'hc2bfd3c7, 32'h429623b4};
test_output[201] = '{32'h42beeedf};
test_index[201] = '{3};
test_input[1616:1623] = '{32'h425be194, 32'h41ee8132, 32'h4209f16b, 32'hc1fbef39, 32'h41c4e8f6, 32'hc1261a6f, 32'hbec2fe40, 32'h42594851};
test_output[202] = '{32'h425be194};
test_index[202] = '{0};
test_input[1624:1631] = '{32'h42346359, 32'h42468a5b, 32'h42098462, 32'hc20d441a, 32'hc249f017, 32'hc26814a2, 32'hc1f916dd, 32'h428c074c};
test_output[203] = '{32'h428c074c};
test_index[203] = '{7};
test_input[1632:1639] = '{32'hc2ae3bac, 32'h41e68472, 32'hc28bab1d, 32'hc2054650, 32'h4086628e, 32'h4216f102, 32'h428b1420, 32'hc2b38c82};
test_output[204] = '{32'h428b1420};
test_index[204] = '{6};
test_input[1640:1647] = '{32'h4166715a, 32'h42a4a777, 32'h40c495ea, 32'h42a57c55, 32'h42978d59, 32'hc28d3b97, 32'hc24b2744, 32'hc1951790};
test_output[205] = '{32'h42a57c55};
test_index[205] = '{3};
test_input[1648:1655] = '{32'h402a56af, 32'hc29cadcb, 32'h42be8e8a, 32'h42328bd6, 32'hc1a5219b, 32'hc1eca916, 32'hc2b9c651, 32'h42c3da0b};
test_output[206] = '{32'h42c3da0b};
test_index[206] = '{7};
test_input[1656:1663] = '{32'h42b92056, 32'h41e6e648, 32'hc279aec0, 32'h4282e9e2, 32'hc2a47e36, 32'hc268db55, 32'hc2b7e81d, 32'hc20f3b26};
test_output[207] = '{32'h42b92056};
test_index[207] = '{0};
test_input[1664:1671] = '{32'hc28b5044, 32'h42ba4e74, 32'h426ee3e2, 32'h42afbcb4, 32'hc2b32915, 32'hc2872d99, 32'hc0513934, 32'h422f4cfd};
test_output[208] = '{32'h42ba4e74};
test_index[208] = '{1};
test_input[1672:1679] = '{32'hc1d0ea13, 32'hc1bda63e, 32'h42569d26, 32'hc2c53644, 32'hc2318ddb, 32'h420f9227, 32'h4277c9be, 32'h426ec651};
test_output[209] = '{32'h4277c9be};
test_index[209] = '{6};
test_input[1680:1687] = '{32'hc27e1625, 32'hc2c1d477, 32'h4209fbb9, 32'h42c0d61b, 32'hc1c189a3, 32'h40a61c41, 32'h40d6153b, 32'h42306dfc};
test_output[210] = '{32'h42c0d61b};
test_index[210] = '{3};
test_input[1688:1695] = '{32'h418dcb15, 32'hc107598c, 32'hc1952715, 32'h42c1ce0a, 32'h42a11d1f, 32'h428c6900, 32'hc29f0cc4, 32'hc25be6c1};
test_output[211] = '{32'h42c1ce0a};
test_index[211] = '{3};
test_input[1696:1703] = '{32'h429c4175, 32'h420a1736, 32'h42ba9c63, 32'hc1b42252, 32'hc173a102, 32'hc27764ef, 32'hc181e9de, 32'hc260c9cb};
test_output[212] = '{32'h42ba9c63};
test_index[212] = '{2};
test_input[1704:1711] = '{32'h42b2d7fc, 32'hc239bacc, 32'h414d061f, 32'hc27bcc5e, 32'h424246bf, 32'h41b062bd, 32'hc17b7a84, 32'hc1df95ce};
test_output[213] = '{32'h42b2d7fc};
test_index[213] = '{0};
test_input[1712:1719] = '{32'h426d29cc, 32'h420bd976, 32'hc20f2061, 32'h428b3aad, 32'h42a953a9, 32'h42c5135e, 32'hc162c2a4, 32'hc10affbe};
test_output[214] = '{32'h42c5135e};
test_index[214] = '{5};
test_input[1720:1727] = '{32'hc1e4e7a3, 32'hc232f3e5, 32'h42bd1a90, 32'h42768dff, 32'hc27b42c0, 32'h41a83d08, 32'h420d0eb7, 32'h429d9740};
test_output[215] = '{32'h42bd1a90};
test_index[215] = '{2};
test_input[1728:1735] = '{32'h429a418f, 32'h42833c69, 32'hc2918637, 32'h421896bc, 32'h42855225, 32'hc2c72366, 32'h41e02b0b, 32'h42419b41};
test_output[216] = '{32'h429a418f};
test_index[216] = '{0};
test_input[1736:1743] = '{32'hc10ae044, 32'h41f79d0c, 32'hc2a1a215, 32'hc232dfcf, 32'hc2845706, 32'h4295bbbb, 32'h42ac5e52, 32'h42b97f97};
test_output[217] = '{32'h42b97f97};
test_index[217] = '{7};
test_input[1744:1751] = '{32'hc2970c58, 32'hc2a88b2c, 32'hc253970c, 32'hc05bad4c, 32'hc1d5aaad, 32'h41a1022f, 32'h41b25a82, 32'hc1a3b181};
test_output[218] = '{32'h41b25a82};
test_index[218] = '{6};
test_input[1752:1759] = '{32'hc21c420d, 32'hc221de35, 32'hc2407837, 32'h40178f52, 32'h42b37fae, 32'h3fe42ef1, 32'h3fbe4711, 32'hc262fc47};
test_output[219] = '{32'h42b37fae};
test_index[219] = '{4};
test_input[1760:1767] = '{32'h421291d6, 32'h41bfac28, 32'hc26daed6, 32'hc24003a6, 32'hc210b294, 32'hc2407e7c, 32'h420c5fcc, 32'h42851a85};
test_output[220] = '{32'h42851a85};
test_index[220] = '{7};
test_input[1768:1775] = '{32'h42a4e826, 32'h41d7ffa4, 32'hc26cc3aa, 32'hc219ae31, 32'hc1b9de53, 32'hc139fa55, 32'h42bcffad, 32'h42972e32};
test_output[221] = '{32'h42bcffad};
test_index[221] = '{6};
test_input[1776:1783] = '{32'h425c7220, 32'h41bf2214, 32'h42a00d40, 32'hc28ec39d, 32'hc2a61f96, 32'hc26544a6, 32'hc1503436, 32'hc250c8ec};
test_output[222] = '{32'h42a00d40};
test_index[222] = '{2};
test_input[1784:1791] = '{32'hc2ba870b, 32'hc25814a3, 32'hc2a77664, 32'hc232f68f, 32'hc274b38b, 32'h4257035a, 32'hc2485b3a, 32'hc2938e3e};
test_output[223] = '{32'h4257035a};
test_index[223] = '{5};
test_input[1792:1799] = '{32'h42a64367, 32'h42552746, 32'h41939ea0, 32'hc2ad5f68, 32'hc26c3e7b, 32'hc2815219, 32'h4282d32d, 32'h42b0e9c8};
test_output[224] = '{32'h42b0e9c8};
test_index[224] = '{7};
test_input[1800:1807] = '{32'h41812422, 32'h42813cb7, 32'h416b5211, 32'h4292ddb4, 32'hc277ffaf, 32'h42726697, 32'h4250966a, 32'h41cae8d9};
test_output[225] = '{32'h4292ddb4};
test_index[225] = '{3};
test_input[1808:1815] = '{32'hc2c3deea, 32'hc2599547, 32'hc1f3abd4, 32'hc2972a9a, 32'h41873773, 32'hc1e22937, 32'hc23851f4, 32'hc2594d16};
test_output[226] = '{32'h41873773};
test_index[226] = '{4};
test_input[1816:1823] = '{32'h42c69332, 32'h4252777c, 32'h41ba0d8d, 32'hc1392484, 32'h42835b62, 32'hc0a74011, 32'hc25a1b0a, 32'hc2a96722};
test_output[227] = '{32'h42c69332};
test_index[227] = '{0};
test_input[1824:1831] = '{32'hc29a9c13, 32'h424f4c15, 32'hc2a5fa44, 32'h4237ad10, 32'hc21afdb3, 32'h428d0239, 32'hc1ef485c, 32'h429a6629};
test_output[228] = '{32'h429a6629};
test_index[228] = '{7};
test_input[1832:1839] = '{32'hc28fd76c, 32'hc16eb776, 32'h41df7c40, 32'h40105b24, 32'hc12b21ab, 32'hc204a0cc, 32'hc18a5246, 32'h42a74086};
test_output[229] = '{32'h42a74086};
test_index[229] = '{7};
test_input[1840:1847] = '{32'hc24c4b50, 32'h4222d1f8, 32'h42bd5b83, 32'hc2032314, 32'hc2bd876a, 32'hc2c0b64c, 32'hc2acf673, 32'hc295ca64};
test_output[230] = '{32'h42bd5b83};
test_index[230] = '{2};
test_input[1848:1855] = '{32'h42b3c2b2, 32'h42aa4100, 32'h428dbdba, 32'h4288ce5d, 32'h417170aa, 32'hc29d38ec, 32'hc197bf37, 32'hc1dfec4e};
test_output[231] = '{32'h42b3c2b2};
test_index[231] = '{0};
test_input[1856:1863] = '{32'h4281a246, 32'hc22a6cb3, 32'h41fc3c28, 32'h42af1da8, 32'hc284adcf, 32'hc0098791, 32'h421dfad4, 32'hc29dbd57};
test_output[232] = '{32'h42af1da8};
test_index[232] = '{3};
test_input[1864:1871] = '{32'h4209d054, 32'hc2b13cbb, 32'hc2795b80, 32'h41b1d52e, 32'hc1adc170, 32'h41ac64d6, 32'hc275207c, 32'hc2b6a44f};
test_output[233] = '{32'h4209d054};
test_index[233] = '{0};
test_input[1872:1879] = '{32'hc254f03b, 32'hc1c90b40, 32'hc2b147d9, 32'hc27b1112, 32'h42adb187, 32'h4246f7cf, 32'h411c9e8b, 32'hc177395a};
test_output[234] = '{32'h42adb187};
test_index[234] = '{4};
test_input[1880:1887] = '{32'h407f56b7, 32'h41ed97ba, 32'hc0bedfc8, 32'h428d05f8, 32'hc2b7935a, 32'hc2bad630, 32'hc1f5776d, 32'h41ff51c0};
test_output[235] = '{32'h428d05f8};
test_index[235] = '{3};
test_input[1888:1895] = '{32'h41facf51, 32'h428bcfad, 32'hc2921053, 32'hc1766232, 32'hc1d7523a, 32'hc29b3260, 32'h406b4659, 32'hc2b7955c};
test_output[236] = '{32'h428bcfad};
test_index[236] = '{1};
test_input[1896:1903] = '{32'hc21ad32e, 32'hc25de600, 32'hc20831c7, 32'h42a648ed, 32'hc0ece842, 32'hc2556523, 32'h42a89aed, 32'h419b50bf};
test_output[237] = '{32'h42a89aed};
test_index[237] = '{6};
test_input[1904:1911] = '{32'h4290380c, 32'hc2b3059b, 32'h4241ac7b, 32'h424bda1a, 32'h41a8a582, 32'h41200cf0, 32'hc2accea5, 32'hc2c74f36};
test_output[238] = '{32'h4290380c};
test_index[238] = '{0};
test_input[1912:1919] = '{32'h40ddc299, 32'h4224bb8c, 32'h42a957a0, 32'hc2a03211, 32'h4286b581, 32'hc2236794, 32'h423d7f38, 32'hc276992a};
test_output[239] = '{32'h42a957a0};
test_index[239] = '{2};
test_input[1920:1927] = '{32'h4238c839, 32'hc23c860e, 32'hc1fae521, 32'hc276706c, 32'hc2a0358e, 32'hc227a0bd, 32'hc2b096bc, 32'hc226c670};
test_output[240] = '{32'h4238c839};
test_index[240] = '{0};
test_input[1928:1935] = '{32'hc27252fe, 32'hc1a44137, 32'hc1447906, 32'hc1e15b76, 32'hc29ebbb9, 32'hc2111435, 32'hc0597b87, 32'h42b1aa6b};
test_output[241] = '{32'h42b1aa6b};
test_index[241] = '{7};
test_input[1936:1943] = '{32'hc1baa1c7, 32'h42bcced4, 32'h429c044e, 32'hc20f90ad, 32'hc1e38090, 32'h42918e78, 32'hc2abb0ec, 32'hc268a9fa};
test_output[242] = '{32'h42bcced4};
test_index[242] = '{1};
test_input[1944:1951] = '{32'hc18c2f2a, 32'h42a75094, 32'h4153b849, 32'hc202f0e5, 32'h42c4980a, 32'h413b2bd4, 32'hc2a24484, 32'hc11d17b9};
test_output[243] = '{32'h42c4980a};
test_index[243] = '{4};
test_input[1952:1959] = '{32'hc14118ce, 32'h421811d6, 32'hc283b0e9, 32'hc2ac8f39, 32'hc2b42891, 32'h428297dd, 32'hc28b7daf, 32'hc26c8894};
test_output[244] = '{32'h428297dd};
test_index[244] = '{5};
test_input[1960:1967] = '{32'h427cb40c, 32'h42b30061, 32'h41fcab93, 32'h42bf7625, 32'hc0a493dd, 32'hc2b2ffdc, 32'h42881484, 32'h42124b72};
test_output[245] = '{32'h42bf7625};
test_index[245] = '{3};
test_input[1968:1975] = '{32'hc2239ed8, 32'hc2903564, 32'h423c547d, 32'hc148cc41, 32'h41c36347, 32'hc2254827, 32'hc2583935, 32'h429e56fc};
test_output[246] = '{32'h429e56fc};
test_index[246] = '{7};
test_input[1976:1983] = '{32'hc1727daf, 32'h42c078ea, 32'h421fe0c7, 32'h421c3e12, 32'h416cde95, 32'h410805b5, 32'h425eac3b, 32'h4160ca24};
test_output[247] = '{32'h42c078ea};
test_index[247] = '{1};
test_input[1984:1991] = '{32'h3faa9c9b, 32'hc26e7606, 32'hc246140a, 32'h42614b7e, 32'hc0f71fc8, 32'hc28fe364, 32'h4195b2dc, 32'h426c3efa};
test_output[248] = '{32'h426c3efa};
test_index[248] = '{7};
test_input[1992:1999] = '{32'h42a5f0ce, 32'hc160037a, 32'hc29a05b1, 32'h42b209d6, 32'hc214430e, 32'hc27059f6, 32'h41b115c7, 32'h420dddae};
test_output[249] = '{32'h42b209d6};
test_index[249] = '{3};
test_input[2000:2007] = '{32'h42ab5127, 32'hc199ded8, 32'h40ae4370, 32'h4256a22b, 32'hc28c8398, 32'h42bf7883, 32'h41d02b45, 32'h41f11146};
test_output[250] = '{32'h42bf7883};
test_index[250] = '{5};
test_input[2008:2015] = '{32'hc28ca8aa, 32'hc27d0861, 32'h42c511cd, 32'hc25e3fe4, 32'h427e6672, 32'h4229e8a3, 32'h4122ad26, 32'h424f6ea2};
test_output[251] = '{32'h42c511cd};
test_index[251] = '{2};
test_input[2016:2023] = '{32'hc26ff754, 32'hc2c6a3e7, 32'h41fc8281, 32'h42470e44, 32'h42a7741b, 32'h42ac2681, 32'h40fbfb59, 32'h428a6263};
test_output[252] = '{32'h42ac2681};
test_index[252] = '{5};
test_input[2024:2031] = '{32'hc1b5336c, 32'hc2b51acf, 32'hc18b7706, 32'hc2b85d26, 32'h4297ab1f, 32'hc2afa3b9, 32'hc12b91de, 32'h4185825a};
test_output[253] = '{32'h4297ab1f};
test_index[253] = '{4};
test_input[2032:2039] = '{32'h429ea048, 32'hc29a62cf, 32'hc2215961, 32'hc265a350, 32'hc294077f, 32'hc1e6f6bd, 32'hc1d638d1, 32'hc2b5d8da};
test_output[254] = '{32'h429ea048};
test_index[254] = '{0};
test_input[2040:2047] = '{32'h41d424a5, 32'hc0d6cac9, 32'h421b4640, 32'hc2183d10, 32'h42a0d567, 32'hc0903071, 32'hc2974576, 32'hc29efd9c};
test_output[255] = '{32'h42a0d567};
test_index[255] = '{4};
test_input[2048:2055] = '{32'hc2be90ed, 32'hc1dc3b51, 32'h42b511dc, 32'h426e2562, 32'h42b33097, 32'h42765cf1, 32'h42527cc7, 32'hc286739b};
test_output[256] = '{32'h42b511dc};
test_index[256] = '{2};
test_input[2056:2063] = '{32'hc01dcafe, 32'hc2af712e, 32'hc28ede37, 32'h4278b770, 32'h419126ad, 32'h41a64353, 32'h416c3535, 32'hc097bfaf};
test_output[257] = '{32'h4278b770};
test_index[257] = '{3};
test_input[2064:2071] = '{32'hc2a20771, 32'h41504e90, 32'hc221b1ed, 32'hc288aa5b, 32'h42308f27, 32'hc297fcf5, 32'hc24cdb79, 32'hc2586513};
test_output[258] = '{32'h42308f27};
test_index[258] = '{4};
test_input[2072:2079] = '{32'hc2a157fe, 32'hc238267e, 32'hc2ba4f56, 32'h41ef94de, 32'hc2c7eb40, 32'hc1f7db01, 32'hc235bdab, 32'h420c06d0};
test_output[259] = '{32'h420c06d0};
test_index[259] = '{7};
test_input[2080:2087] = '{32'h429c5caf, 32'hc291d412, 32'hc2574b42, 32'h42922409, 32'hc1c629a3, 32'h42a644b3, 32'hc1a49c73, 32'hc2c073d6};
test_output[260] = '{32'h42a644b3};
test_index[260] = '{5};
test_input[2088:2095] = '{32'h422c912d, 32'hc2aefb41, 32'h4194aaff, 32'h4119c645, 32'h41dcbdbb, 32'hc039d126, 32'h4294684b, 32'h42803d78};
test_output[261] = '{32'h4294684b};
test_index[261] = '{6};
test_input[2096:2103] = '{32'hc2b5cb3e, 32'h420c09f0, 32'hc29fbc82, 32'hc2a1f299, 32'hc1f9ddb0, 32'hc226ebaf, 32'hc1e69687, 32'h42aacab1};
test_output[262] = '{32'h42aacab1};
test_index[262] = '{7};
test_input[2104:2111] = '{32'hc15ead8f, 32'h413715df, 32'hc17a34e8, 32'hc1b724ae, 32'hc2c69b08, 32'h42a06f43, 32'hc232c97e, 32'hc2bac159};
test_output[263] = '{32'h42a06f43};
test_index[263] = '{5};
test_input[2112:2119] = '{32'hc11eb19c, 32'h41f23f52, 32'hc2589c59, 32'hc2513ccc, 32'hc2089980, 32'hc13b8a44, 32'h42bbb63a, 32'hc25f6636};
test_output[264] = '{32'h42bbb63a};
test_index[264] = '{6};
test_input[2120:2127] = '{32'h4085f94c, 32'h4252933f, 32'h42c54cea, 32'hc1977b2a, 32'h414caf0b, 32'h40c19722, 32'h42027956, 32'hc2c7be81};
test_output[265] = '{32'h42c54cea};
test_index[265] = '{2};
test_input[2128:2135] = '{32'h4021ea5c, 32'hc22f734f, 32'hc2a29ddd, 32'h423ad253, 32'hc2b73574, 32'hc2991409, 32'h42aec9d0, 32'hc29f774f};
test_output[266] = '{32'h42aec9d0};
test_index[266] = '{6};
test_input[2136:2143] = '{32'h4073098e, 32'hc0145e19, 32'h4286b5ec, 32'hc192db08, 32'hc1f957d3, 32'h422c9816, 32'hc0920fa0, 32'hbfd228ea};
test_output[267] = '{32'h4286b5ec};
test_index[267] = '{2};
test_input[2144:2151] = '{32'h426d2069, 32'hc2aad8a7, 32'hc291f311, 32'h428d8459, 32'hc2378853, 32'h419dd6ca, 32'hc291ce04, 32'h42956793};
test_output[268] = '{32'h42956793};
test_index[268] = '{7};
test_input[2152:2159] = '{32'hc24d6870, 32'h4232b981, 32'hc28d6851, 32'hc20ec19f, 32'hbf9f655c, 32'h410f7b03, 32'h42b6ced9, 32'hc294d386};
test_output[269] = '{32'h42b6ced9};
test_index[269] = '{6};
test_input[2160:2167] = '{32'h4295fccc, 32'hc1776800, 32'hc288cdac, 32'hc229414a, 32'h42a3b511, 32'hc2351e2d, 32'hc26eaf77, 32'h42c4ba49};
test_output[270] = '{32'h42c4ba49};
test_index[270] = '{7};
test_input[2168:2175] = '{32'hc0c0b02b, 32'hc19dbe6c, 32'h425538d1, 32'h40e7407a, 32'hc2b8a3f9, 32'hc28897c1, 32'h41c5ce36, 32'hc207ebd2};
test_output[271] = '{32'h425538d1};
test_index[271] = '{2};
test_input[2176:2183] = '{32'h4220c640, 32'hc10671af, 32'hc27823fa, 32'hc2693a59, 32'h40339ff7, 32'hc11190e0, 32'hc249a8a8, 32'h42145fb7};
test_output[272] = '{32'h4220c640};
test_index[272] = '{0};
test_input[2184:2191] = '{32'h41c8745e, 32'h42c5ed4b, 32'h418b9967, 32'h4255d1d5, 32'hc1784241, 32'h42c20677, 32'hc1a5e5f2, 32'hc1ee0b7c};
test_output[273] = '{32'h42c5ed4b};
test_index[273] = '{1};
test_input[2192:2199] = '{32'hc2536682, 32'h42a17f14, 32'h422d04b4, 32'hc22f5477, 32'h40ec35b8, 32'hc20d0f24, 32'hc291df8b, 32'h41a16234};
test_output[274] = '{32'h42a17f14};
test_index[274] = '{1};
test_input[2200:2207] = '{32'h425b707d, 32'hc2b12d54, 32'hc0cd8575, 32'h4284e42a, 32'hc238aab4, 32'h42a10fa4, 32'h4153bd10, 32'h410623f9};
test_output[275] = '{32'h42a10fa4};
test_index[275] = '{5};
test_input[2208:2215] = '{32'hc262d4ed, 32'hc24d2131, 32'h42c15452, 32'hc2632cde, 32'hc229c50e, 32'hc24f82fe, 32'h423e6129, 32'h41a51164};
test_output[276] = '{32'h42c15452};
test_index[276] = '{2};
test_input[2216:2223] = '{32'hc2055df9, 32'hc15dc2ef, 32'hc26cd1f0, 32'h419af84a, 32'hc1ea091d, 32'h42869060, 32'h41d995e9, 32'h42c3092a};
test_output[277] = '{32'h42c3092a};
test_index[277] = '{7};
test_input[2224:2231] = '{32'h42946f70, 32'h42b4c9e5, 32'hc2283821, 32'hc2a4d9d9, 32'hc26bb1d1, 32'hc299fd77, 32'hc2788305, 32'hc2b2270c};
test_output[278] = '{32'h42b4c9e5};
test_index[278] = '{1};
test_input[2232:2239] = '{32'hc1df1320, 32'h422afced, 32'h42a496d5, 32'hc2a3bb94, 32'h42ae922c, 32'hc2a6f917, 32'h427f86e6, 32'hc25d3927};
test_output[279] = '{32'h42ae922c};
test_index[279] = '{4};
test_input[2240:2247] = '{32'h4275fd2d, 32'h42c21de1, 32'hc1872a5e, 32'h42200148, 32'hc2a883ba, 32'h3fa6cc04, 32'hc0ac01c2, 32'h42292500};
test_output[280] = '{32'h42c21de1};
test_index[280] = '{1};
test_input[2248:2255] = '{32'hc2a15486, 32'hc29ace3b, 32'h41302242, 32'h429b0846, 32'h423de7ba, 32'h40fe2a87, 32'h419ee480, 32'h42c64a0f};
test_output[281] = '{32'h42c64a0f};
test_index[281] = '{7};
test_input[2256:2263] = '{32'h42a0231f, 32'hc1e982ae, 32'hc2541551, 32'h41969f85, 32'h41fcb2c2, 32'h421d2f1e, 32'hc28f83ee, 32'h4031a4e8};
test_output[282] = '{32'h42a0231f};
test_index[282] = '{0};
test_input[2264:2271] = '{32'h407003dc, 32'hc26c939a, 32'h411cc6ef, 32'hc18a6a5b, 32'h4234fc9a, 32'h4294988a, 32'hc2c49d7d, 32'hc23ed41e};
test_output[283] = '{32'h4294988a};
test_index[283] = '{5};
test_input[2272:2279] = '{32'hc142c1b8, 32'hc296404f, 32'hc0aee615, 32'hc2890ad4, 32'hc14a6f8a, 32'h4175da62, 32'hc25e262c, 32'hc27e3a77};
test_output[284] = '{32'h4175da62};
test_index[284] = '{5};
test_input[2280:2287] = '{32'hc22ef804, 32'h4293d3d3, 32'h41384ee3, 32'h4253788d, 32'hc2bfe048, 32'h420859a6, 32'h42a394cd, 32'hc2bf5b3f};
test_output[285] = '{32'h42a394cd};
test_index[285] = '{6};
test_input[2288:2295] = '{32'hc11e7760, 32'hc2aaa1d6, 32'hc2097f58, 32'hc22268c1, 32'h429ee87a, 32'hc23e1964, 32'hc23cf2d7, 32'hc2279be0};
test_output[286] = '{32'h429ee87a};
test_index[286] = '{4};
test_input[2296:2303] = '{32'hc1960ba1, 32'h42509baa, 32'hc22c76a1, 32'h42c7ecc6, 32'h425675dc, 32'hc2497b69, 32'h4228471f, 32'h423b807c};
test_output[287] = '{32'h42c7ecc6};
test_index[287] = '{3};
test_input[2304:2311] = '{32'h42a9de12, 32'h428ef2f1, 32'h42c62744, 32'h41d23910, 32'hc243ef0e, 32'hc22d9885, 32'h4266ab8a, 32'h40179e63};
test_output[288] = '{32'h42c62744};
test_index[288] = '{2};
test_input[2312:2319] = '{32'hc22c0ddf, 32'h42c555a3, 32'hc1b470d5, 32'hc2aa40cd, 32'hc1c7f3d7, 32'h41091285, 32'hc29e06ee, 32'hc282257e};
test_output[289] = '{32'h42c555a3};
test_index[289] = '{1};
test_input[2320:2327] = '{32'hc2790d70, 32'hc2a4eaef, 32'h425c1dbe, 32'h428a7830, 32'h4247ff27, 32'h42945b53, 32'hc25c4397, 32'h412a3383};
test_output[290] = '{32'h42945b53};
test_index[290] = '{5};
test_input[2328:2335] = '{32'hc231436a, 32'hc2c66582, 32'h42a78570, 32'h426cfc70, 32'hc27cf29b, 32'hc2ac4f04, 32'hc1d82df2, 32'h4006335f};
test_output[291] = '{32'h42a78570};
test_index[291] = '{2};
test_input[2336:2343] = '{32'h42c45aeb, 32'h425f721f, 32'h41e2b35b, 32'hc2271c53, 32'h414e0213, 32'h4265a297, 32'hc1cdb99d, 32'hc2b618bd};
test_output[292] = '{32'h42c45aeb};
test_index[292] = '{0};
test_input[2344:2351] = '{32'hc26f216b, 32'hc2c62cfd, 32'hbf70c00f, 32'h42280ebd, 32'h419574ff, 32'hc2910cc5, 32'hc24c2902, 32'h42bdc790};
test_output[293] = '{32'h42bdc790};
test_index[293] = '{7};
test_input[2352:2359] = '{32'h4273251e, 32'h425ba5a4, 32'h428ae514, 32'hc2552f04, 32'h41961b8d, 32'h40d21383, 32'h41b6b083, 32'hc2b8884c};
test_output[294] = '{32'h428ae514};
test_index[294] = '{2};
test_input[2360:2367] = '{32'hc265ea01, 32'hc2857812, 32'h418fd915, 32'h42bc3105, 32'h41adcba7, 32'h42a811d9, 32'h42709f9f, 32'hc1c0f6aa};
test_output[295] = '{32'h42bc3105};
test_index[295] = '{3};
test_input[2368:2375] = '{32'h425fc9ea, 32'h4287fa45, 32'hc21f7522, 32'hc2868374, 32'hc2780863, 32'hc23acbd6, 32'h40ab990f, 32'h42948d87};
test_output[296] = '{32'h42948d87};
test_index[296] = '{7};
test_input[2376:2383] = '{32'h412425c2, 32'h42c413bc, 32'h417a0134, 32'h428c6ce0, 32'hc2c246ef, 32'h4299e195, 32'h40fedd93, 32'hc1fdd4a6};
test_output[297] = '{32'h42c413bc};
test_index[297] = '{1};
test_input[2384:2391] = '{32'hc118fbe7, 32'h4295cd46, 32'hc2a24e57, 32'hc2a0c988, 32'hc2c690db, 32'h42b0dca5, 32'h42671897, 32'hc1a47d85};
test_output[298] = '{32'h42b0dca5};
test_index[298] = '{5};
test_input[2392:2399] = '{32'hc1f2ead6, 32'h4295fb16, 32'hc14262a9, 32'hc12a3424, 32'hc1b57356, 32'hc11f127d, 32'hc0ad1321, 32'hc207026c};
test_output[299] = '{32'h4295fb16};
test_index[299] = '{1};
test_input[2400:2407] = '{32'h418f1b34, 32'h428cc298, 32'h41a5d6ed, 32'hc26dae96, 32'h42ad5e57, 32'hc10f1f0b, 32'h42211be9, 32'hc28e76a8};
test_output[300] = '{32'h42ad5e57};
test_index[300] = '{4};
test_input[2408:2415] = '{32'h41ff3217, 32'h420c3a05, 32'h42bfe821, 32'h426f49fe, 32'h428be2ca, 32'hc258f96c, 32'h4253a2f8, 32'hbf06f1d4};
test_output[301] = '{32'h42bfe821};
test_index[301] = '{2};
test_input[2416:2423] = '{32'hc1c35ee9, 32'h4238f18b, 32'h428b7635, 32'h4207f3eb, 32'h42ab7751, 32'hc234277e, 32'hc28f9f54, 32'h4281eb3a};
test_output[302] = '{32'h42ab7751};
test_index[302] = '{4};
test_input[2424:2431] = '{32'h4220d044, 32'h428732b1, 32'h411b839e, 32'h41dbcf0e, 32'hc2398ae9, 32'hc2c603fc, 32'hc0527b41, 32'h42bef4ea};
test_output[303] = '{32'h42bef4ea};
test_index[303] = '{7};
test_input[2432:2439] = '{32'h42095723, 32'hc1b63cbc, 32'h424a0f5e, 32'hc2c59375, 32'hc28fbc5c, 32'hc0e5f047, 32'hc2c135e9, 32'hc0b236f0};
test_output[304] = '{32'h424a0f5e};
test_index[304] = '{2};
test_input[2440:2447] = '{32'hc241fe1c, 32'hc098be7e, 32'hc13ae6d4, 32'h4207b426, 32'hc18c216b, 32'hc28c2ca6, 32'hc2a478c7, 32'hc2abf1ef};
test_output[305] = '{32'h4207b426};
test_index[305] = '{3};
test_input[2448:2455] = '{32'hc1c43971, 32'hc23d941f, 32'h42bbf5be, 32'h421b188f, 32'h421a2791, 32'hc29bd01f, 32'h427b443a, 32'hc205e70f};
test_output[306] = '{32'h42bbf5be};
test_index[306] = '{2};
test_input[2456:2463] = '{32'h429480aa, 32'hc1c562cd, 32'h41a22f56, 32'hc296744a, 32'hc2a89d5e, 32'hc1f6b93a, 32'h41bbf2a6, 32'h4161d9b1};
test_output[307] = '{32'h429480aa};
test_index[307] = '{0};
test_input[2464:2471] = '{32'h42c292a3, 32'h427f0c43, 32'hc1ce5046, 32'hc2395fab, 32'hc2131c2e, 32'h3fa74978, 32'h41112464, 32'hc09f3d7c};
test_output[308] = '{32'h42c292a3};
test_index[308] = '{0};
test_input[2472:2479] = '{32'hc227799f, 32'h40a2bd70, 32'h42b1fa31, 32'hbf3433af, 32'hc0bb5db8, 32'hc29fadb0, 32'h422e8d25, 32'hc2218a49};
test_output[309] = '{32'h42b1fa31};
test_index[309] = '{2};
test_input[2480:2487] = '{32'hc27e8a01, 32'hc1eddcdd, 32'hc249bb0f, 32'hc2a8dbc1, 32'h42b2ec98, 32'hc17bf27b, 32'h42b90085, 32'h41d0d42d};
test_output[310] = '{32'h42b90085};
test_index[310] = '{6};
test_input[2488:2495] = '{32'hc1b6bdac, 32'hc2bcaeae, 32'h4276017c, 32'h42362063, 32'h42bf8e0f, 32'hc13213e3, 32'h42c3aeaf, 32'h41f7b45f};
test_output[311] = '{32'h42c3aeaf};
test_index[311] = '{6};
test_input[2496:2503] = '{32'h4238336a, 32'h4287701d, 32'hc161d8fe, 32'hc24c8110, 32'hc26103d6, 32'h42ae6f19, 32'hc2b7a462, 32'hc2479e1a};
test_output[312] = '{32'h42ae6f19};
test_index[312] = '{5};
test_input[2504:2511] = '{32'hc276e612, 32'h423b5f30, 32'hc11077ae, 32'h412c57ea, 32'hc2599d3c, 32'h421bf134, 32'h41736916, 32'h4201ae5f};
test_output[313] = '{32'h423b5f30};
test_index[313] = '{1};
test_input[2512:2519] = '{32'hc1f81c8c, 32'hc284c8c5, 32'hc2035b9f, 32'h42501c3d, 32'hc184582a, 32'hc288363f, 32'h42c2565e, 32'h42ade65a};
test_output[314] = '{32'h42c2565e};
test_index[314] = '{6};
test_input[2520:2527] = '{32'hc1e55995, 32'hc20589f1, 32'hc103ab7f, 32'hc131d8cc, 32'hc1893217, 32'h428d6209, 32'hc11f2ee4, 32'hc1d32aac};
test_output[315] = '{32'h428d6209};
test_index[315] = '{5};
test_input[2528:2535] = '{32'hc1a2042f, 32'hc206c184, 32'h42906826, 32'hc1cd0889, 32'hc19a81e9, 32'hc29343d6, 32'hc1effcdf, 32'h4255d898};
test_output[316] = '{32'h42906826};
test_index[316] = '{2};
test_input[2536:2543] = '{32'h42be16a9, 32'hc270d107, 32'hc20edb0b, 32'hc29bece2, 32'hc18b9633, 32'hc21b5ebe, 32'hc2981694, 32'h42c1a336};
test_output[317] = '{32'h42c1a336};
test_index[317] = '{7};
test_input[2544:2551] = '{32'hc0ac60ab, 32'hc242da6d, 32'hc290f44f, 32'hc2832304, 32'hc2a2ea37, 32'hc29638bc, 32'h428e4a86, 32'h42b60612};
test_output[318] = '{32'h42b60612};
test_index[318] = '{7};
test_input[2552:2559] = '{32'h42398e6d, 32'h41a4059f, 32'h414b770e, 32'hc2162484, 32'hc1f25e10, 32'h42602a72, 32'h424e211b, 32'hc212c8c1};
test_output[319] = '{32'h42602a72};
test_index[319] = '{5};
test_input[2560:2567] = '{32'h42b1ca97, 32'hc121fcc6, 32'h422e3dc9, 32'hc2b31928, 32'hc2c1211e, 32'hc2c7c4d6, 32'h41464d04, 32'hc2c15319};
test_output[320] = '{32'h42b1ca97};
test_index[320] = '{0};
test_input[2568:2575] = '{32'h42a61cb9, 32'hbfe3036e, 32'hc255c703, 32'h421e9b1c, 32'hc28d6366, 32'hc24d73e7, 32'h42bd10c4, 32'h42552470};
test_output[321] = '{32'h42bd10c4};
test_index[321] = '{6};
test_input[2576:2583] = '{32'h42b72090, 32'hc26dd336, 32'h4270e7e6, 32'hc2081127, 32'h4239cecd, 32'hc202c8f8, 32'hc22f9f9f, 32'hc1fa4772};
test_output[322] = '{32'h42b72090};
test_index[322] = '{0};
test_input[2584:2591] = '{32'hc291a621, 32'hc2ae0c35, 32'h42bf83c7, 32'h421f4163, 32'h422cc883, 32'h4299b8c9, 32'hc183b8bd, 32'h418a1d97};
test_output[323] = '{32'h42bf83c7};
test_index[323] = '{2};
test_input[2592:2599] = '{32'h4293e7e7, 32'h424296fc, 32'h42a0b6f1, 32'h417217f8, 32'h42537a72, 32'h42716a22, 32'hc28892c4, 32'h4162801c};
test_output[324] = '{32'h42a0b6f1};
test_index[324] = '{2};
test_input[2600:2607] = '{32'hc299f92b, 32'hc1666522, 32'h42851b52, 32'h429cc763, 32'hc2b4e67c, 32'hc1f016dd, 32'h41ecf171, 32'h424c7dde};
test_output[325] = '{32'h429cc763};
test_index[325] = '{3};
test_input[2608:2615] = '{32'h420c117d, 32'hc018b40b, 32'h425d809b, 32'hc045386d, 32'h41e71331, 32'h42b130f6, 32'hc1fc4842, 32'hc27e36da};
test_output[326] = '{32'h42b130f6};
test_index[326] = '{5};
test_input[2616:2623] = '{32'h42a313d1, 32'hc286a92e, 32'hc094f6bf, 32'hc256b563, 32'hc2367cba, 32'h409ba6bb, 32'hc21644bf, 32'hc284a0e7};
test_output[327] = '{32'h42a313d1};
test_index[327] = '{0};
test_input[2624:2631] = '{32'hc1437d16, 32'h41014c62, 32'hc1076aa6, 32'h42a013e6, 32'hc0baffc9, 32'hc284b6f0, 32'hc22bf7e0, 32'hc2c5dca5};
test_output[328] = '{32'h42a013e6};
test_index[328] = '{3};
test_input[2632:2639] = '{32'h4292b181, 32'hc1a4fa08, 32'h42c05bf9, 32'hc26bc236, 32'h42b17669, 32'h42b10aee, 32'h4204ad90, 32'hc1aeb745};
test_output[329] = '{32'h42c05bf9};
test_index[329] = '{2};
test_input[2640:2647] = '{32'hc216e196, 32'hc29cb268, 32'hc2be7b53, 32'hc2346929, 32'h4294face, 32'h42577292, 32'h427821c0, 32'hc1fa343e};
test_output[330] = '{32'h4294face};
test_index[330] = '{4};
test_input[2648:2655] = '{32'hc1facebb, 32'h408663f5, 32'hc1de02b1, 32'hc226997e, 32'h40ad4c7f, 32'h4100ac3b, 32'hc1b77d0a, 32'hc2ac8c29};
test_output[331] = '{32'h4100ac3b};
test_index[331] = '{5};
test_input[2656:2663] = '{32'hc1b5e166, 32'hc283c710, 32'hc27c425c, 32'hc1995d02, 32'h3eb544bb, 32'hc26c38ae, 32'hc2ab0b1f, 32'h41749035};
test_output[332] = '{32'h41749035};
test_index[332] = '{7};
test_input[2664:2671] = '{32'h41bbd8c2, 32'hc2aaa2e3, 32'h42bd3033, 32'hc2291748, 32'h426997a7, 32'h4242d361, 32'hc2aa5e63, 32'h429f76b4};
test_output[333] = '{32'h42bd3033};
test_index[333] = '{2};
test_input[2672:2679] = '{32'h40f67a6c, 32'hc28e289d, 32'h41e89974, 32'h421691a0, 32'h426c7cea, 32'hc2c359f4, 32'h419f63ef, 32'hc2905116};
test_output[334] = '{32'h426c7cea};
test_index[334] = '{4};
test_input[2680:2687] = '{32'hc1a677bb, 32'hc25223cf, 32'hc0bcea38, 32'hc2116a3b, 32'h424d206d, 32'hc1947d67, 32'h41caf431, 32'h42c70753};
test_output[335] = '{32'h42c70753};
test_index[335] = '{7};
test_input[2688:2695] = '{32'hc276e0de, 32'hc23bc0d0, 32'hc2638a61, 32'hc23a53f2, 32'h4233dd82, 32'h4204d5d3, 32'hc1672c51, 32'h423d0c18};
test_output[336] = '{32'h423d0c18};
test_index[336] = '{7};
test_input[2696:2703] = '{32'h4184d9bb, 32'hbe105c78, 32'h425116d0, 32'h42ba0efe, 32'h41b1be1f, 32'hc20391fa, 32'hc28e3081, 32'h427ccc0b};
test_output[337] = '{32'h42ba0efe};
test_index[337] = '{3};
test_input[2704:2711] = '{32'hc25bf2e6, 32'h422b2035, 32'hc2a79a3e, 32'h42c04c3b, 32'h414a8148, 32'h42bc8b29, 32'h42a8191d, 32'hc14b0406};
test_output[338] = '{32'h42c04c3b};
test_index[338] = '{3};
test_input[2712:2719] = '{32'hc1c48e88, 32'h42c634e8, 32'hc2a75eb6, 32'hc2675be8, 32'h42aaa15b, 32'h4031b152, 32'h42694fcf, 32'hc277248d};
test_output[339] = '{32'h42c634e8};
test_index[339] = '{1};
test_input[2720:2727] = '{32'h4263d97e, 32'h421678e2, 32'h412b96c1, 32'hc2be9890, 32'hc2a6c837, 32'hc21e2a0e, 32'hc27c698d, 32'hc07bec7b};
test_output[340] = '{32'h4263d97e};
test_index[340] = '{0};
test_input[2728:2735] = '{32'hc1bb0a31, 32'h41638d4f, 32'h423aa5ca, 32'h41035201, 32'h42a2181d, 32'hc2c19c16, 32'hc28045a6, 32'h428366dc};
test_output[341] = '{32'h42a2181d};
test_index[341] = '{4};
test_input[2736:2743] = '{32'h42579ba7, 32'hc23cf05b, 32'hc103ee21, 32'hc18ec624, 32'h427cd600, 32'h4254b00f, 32'hc2c52edf, 32'hc28eb44b};
test_output[342] = '{32'h427cd600};
test_index[342] = '{4};
test_input[2744:2751] = '{32'h42426dde, 32'hc1981372, 32'h41977ebd, 32'hc05eebc4, 32'hc25f9e4e, 32'h42b96060, 32'hc2b63e47, 32'h41dda4b7};
test_output[343] = '{32'h42b96060};
test_index[343] = '{5};
test_input[2752:2759] = '{32'h420cd361, 32'h42b98c46, 32'hc1d3891a, 32'hc23b3e1a, 32'hc22cc1fa, 32'hc2c21dc4, 32'h421cce04, 32'h414e962e};
test_output[344] = '{32'h42b98c46};
test_index[344] = '{1};
test_input[2760:2767] = '{32'h42811416, 32'h428256ea, 32'hc196108a, 32'h4106724a, 32'h42ad5c1f, 32'hc0aa8538, 32'h4250e124, 32'h40858b5d};
test_output[345] = '{32'h42ad5c1f};
test_index[345] = '{4};
test_input[2768:2775] = '{32'hc26c76b3, 32'hc2878f4e, 32'h425a3770, 32'h427ae657, 32'h42adc817, 32'hc21bf304, 32'hc2926f72, 32'h410f8598};
test_output[346] = '{32'h42adc817};
test_index[346] = '{4};
test_input[2776:2783] = '{32'hc1dbec21, 32'hc25c239f, 32'hc0fe47f9, 32'h428d8b67, 32'h427d9e23, 32'hc22e9973, 32'h423944df, 32'hc21ff128};
test_output[347] = '{32'h428d8b67};
test_index[347] = '{3};
test_input[2784:2791] = '{32'hc2c24508, 32'h41877089, 32'hc1c489cf, 32'hc26365bb, 32'hc29c115e, 32'hc27e2bbd, 32'hc2bf2c63, 32'hc1c89266};
test_output[348] = '{32'h41877089};
test_index[348] = '{1};
test_input[2792:2799] = '{32'hc28884fa, 32'h42713e8c, 32'h41d497e6, 32'h42c453cf, 32'h41bbb9ec, 32'h423b563c, 32'h41f316b1, 32'h41f75318};
test_output[349] = '{32'h42c453cf};
test_index[349] = '{3};
test_input[2800:2807] = '{32'h41ef6e7b, 32'hc2428189, 32'h41a8b30a, 32'h41f4f948, 32'h4182e3dd, 32'h4219d0de, 32'hc24df28d, 32'h3eeed3f1};
test_output[350] = '{32'h4219d0de};
test_index[350] = '{5};
test_input[2808:2815] = '{32'h42877bf0, 32'h41f8c3dc, 32'hc2855339, 32'hc2af50be, 32'h415cfec5, 32'h42c35565, 32'h41a5abaa, 32'hc2c0cf37};
test_output[351] = '{32'h42c35565};
test_index[351] = '{5};
test_input[2816:2823] = '{32'h429c5f0f, 32'hc1ae9d00, 32'h41bfb065, 32'h429c9236, 32'h42a3eef5, 32'hc115be51, 32'hc1fca7cf, 32'hc2821c9d};
test_output[352] = '{32'h42a3eef5};
test_index[352] = '{4};
test_input[2824:2831] = '{32'h42135fe1, 32'hc2b213d7, 32'h423a61a2, 32'hbf20e3d4, 32'hc22468c6, 32'h422c8404, 32'hc2b051c2, 32'hc2c2ff92};
test_output[353] = '{32'h423a61a2};
test_index[353] = '{2};
test_input[2832:2839] = '{32'h429581c4, 32'h4211e5e2, 32'h41f8e3e4, 32'h4278b8a6, 32'h42991932, 32'hc205be62, 32'h418d55e4, 32'h42c367ba};
test_output[354] = '{32'h42c367ba};
test_index[354] = '{7};
test_input[2840:2847] = '{32'hc2a5e041, 32'hc281cb77, 32'hc22d4166, 32'hc2c7c9fa, 32'h42adc2b8, 32'h4257be48, 32'h42808f67, 32'h42995134};
test_output[355] = '{32'h42adc2b8};
test_index[355] = '{4};
test_input[2848:2855] = '{32'h427a6782, 32'hc22ff2b6, 32'h409a0016, 32'hc136879f, 32'hc2c6cef4, 32'hc2c583a6, 32'h424a3de0, 32'h42527501};
test_output[356] = '{32'h427a6782};
test_index[356] = '{0};
test_input[2856:2863] = '{32'hc189ed39, 32'hc2a36075, 32'h41070aef, 32'h411a918c, 32'h415abe86, 32'h42ae5810, 32'h41ba0dfb, 32'hc2496e0d};
test_output[357] = '{32'h42ae5810};
test_index[357] = '{5};
test_input[2864:2871] = '{32'h421cfdca, 32'hc272b13b, 32'h42a38610, 32'hc2581565, 32'h42140b27, 32'hc2856e07, 32'h4274af15, 32'hc28a10ea};
test_output[358] = '{32'h42a38610};
test_index[358] = '{2};
test_input[2872:2879] = '{32'hc2b6fb6c, 32'h4053a952, 32'hc1a87753, 32'hc14a2d9c, 32'hc144710b, 32'h4010d837, 32'h42a13c7e, 32'hc25089c8};
test_output[359] = '{32'h42a13c7e};
test_index[359] = '{6};
test_input[2880:2887] = '{32'h413573ca, 32'hc18eac67, 32'h4289e72d, 32'h424d4838, 32'hc28f17bb, 32'h412fcc6c, 32'hc1fe037b, 32'h42a77391};
test_output[360] = '{32'h42a77391};
test_index[360] = '{7};
test_input[2888:2895] = '{32'h41fde906, 32'hc2b10125, 32'hc2b55349, 32'hc1d1b434, 32'hc21c6c86, 32'hc285ae18, 32'hc1e19ef9, 32'hc2329c25};
test_output[361] = '{32'h41fde906};
test_index[361] = '{0};
test_input[2896:2903] = '{32'h42a49391, 32'hc24f3793, 32'h4287ef6f, 32'h42a8a5c4, 32'h40ac7dda, 32'h42973276, 32'h423c568d, 32'h4117a14f};
test_output[362] = '{32'h42a8a5c4};
test_index[362] = '{3};
test_input[2904:2911] = '{32'h41d0550f, 32'h42b7e3f0, 32'h428e5872, 32'h419f7175, 32'h420afb01, 32'hc2940eaf, 32'h42aa89a7, 32'h42b82b06};
test_output[363] = '{32'h42b82b06};
test_index[363] = '{7};
test_input[2912:2919] = '{32'hc1535b43, 32'h419bc2d3, 32'h42342184, 32'hc2840912, 32'h4108f5de, 32'h42b51059, 32'hc29ab945, 32'hc294fd19};
test_output[364] = '{32'h42b51059};
test_index[364] = '{5};
test_input[2920:2927] = '{32'hc2ac4855, 32'h411b6625, 32'hc2664378, 32'h410f4532, 32'hc1e3c5a0, 32'h42905939, 32'h410e08e2, 32'h42577dd6};
test_output[365] = '{32'h42905939};
test_index[365] = '{5};
test_input[2928:2935] = '{32'hc0a37513, 32'h4280566e, 32'hc138a554, 32'h3e6fcf44, 32'hc03db24d, 32'hc2393c3c, 32'h4153513f, 32'h40323d89};
test_output[366] = '{32'h4280566e};
test_index[366] = '{1};
test_input[2936:2943] = '{32'hc25f8c98, 32'h41da7c94, 32'hc2b4c425, 32'h422014b0, 32'hc20c14ee, 32'h4260a1c1, 32'hc284a200, 32'h42189f82};
test_output[367] = '{32'h4260a1c1};
test_index[367] = '{5};
test_input[2944:2951] = '{32'h41c4adce, 32'hc2830a1a, 32'hc2b06720, 32'hc260b393, 32'h41d49358, 32'hc2048ac9, 32'hc29e387e, 32'h4239d233};
test_output[368] = '{32'h4239d233};
test_index[368] = '{7};
test_input[2952:2959] = '{32'hc2b98478, 32'h42b11146, 32'h42308815, 32'hc20eceaf, 32'h3f2e849b, 32'h422e570a, 32'h4225ea32, 32'h4180f78f};
test_output[369] = '{32'h42b11146};
test_index[369] = '{1};
test_input[2960:2967] = '{32'h42b71b3c, 32'h4287391e, 32'h428c52d6, 32'h42014c58, 32'h42a40b25, 32'h42573435, 32'h413f5392, 32'h4288b61c};
test_output[370] = '{32'h42b71b3c};
test_index[370] = '{0};
test_input[2968:2975] = '{32'h41e2d556, 32'h41ba037e, 32'hc2b26c87, 32'h4206a5e9, 32'h42aea64f, 32'hc2a38089, 32'h424d18f9, 32'hc243f437};
test_output[371] = '{32'h42aea64f};
test_index[371] = '{4};
test_input[2976:2983] = '{32'hc27076cb, 32'hc2b4e0c1, 32'h42955c37, 32'hc23206b0, 32'h41f0bbe2, 32'hc298b5e7, 32'h42bcb531, 32'h42b5f3b4};
test_output[372] = '{32'h42bcb531};
test_index[372] = '{6};
test_input[2984:2991] = '{32'hc25c3d43, 32'hc1c0e49e, 32'h42288e86, 32'h42a80631, 32'hc2075904, 32'h42c4933c, 32'hc293345d, 32'hc28c98c9};
test_output[373] = '{32'h42c4933c};
test_index[373] = '{5};
test_input[2992:2999] = '{32'h3fad907a, 32'hc20ad531, 32'h4225a541, 32'hc2828303, 32'hc13fe0d0, 32'hc29c9275, 32'hc2a74a4c, 32'hc2b7aad3};
test_output[374] = '{32'h4225a541};
test_index[374] = '{2};
test_input[3000:3007] = '{32'hbf5fabf6, 32'hbd153535, 32'h42819381, 32'h4216fe67, 32'h4254ea06, 32'hc2959e55, 32'h42a94580, 32'hc2bc820b};
test_output[375] = '{32'h42a94580};
test_index[375] = '{6};
test_input[3008:3015] = '{32'h41b3e71d, 32'h41577e6d, 32'h42848258, 32'h41c235d4, 32'hc28e65fa, 32'hc222ec42, 32'hc2b031c3, 32'hc1ce5bdd};
test_output[376] = '{32'h42848258};
test_index[376] = '{2};
test_input[3016:3023] = '{32'hbf299d9c, 32'hc2182cc6, 32'hc2b1d168, 32'h40184ab1, 32'h408b19ed, 32'h41b933ba, 32'h42c7d911, 32'h420f637b};
test_output[377] = '{32'h42c7d911};
test_index[377] = '{6};
test_input[3024:3031] = '{32'hc29899f0, 32'hc137b128, 32'hc2c0f6a4, 32'hc2a0bd6f, 32'hc18e0347, 32'hc25771a1, 32'hc2024ea6, 32'hc196a53c};
test_output[378] = '{32'hc137b128};
test_index[378] = '{1};
test_input[3032:3039] = '{32'hc20f3f63, 32'hc2c0d9e6, 32'hc16e856a, 32'hc279537c, 32'h424aaf6e, 32'h42adb1de, 32'hc20335b7, 32'hc2971a13};
test_output[379] = '{32'h42adb1de};
test_index[379] = '{5};
test_input[3040:3047] = '{32'h41dd268a, 32'h414f9e70, 32'h424e5e38, 32'hc1093d6b, 32'h429be13f, 32'hc1d65637, 32'h4146fe7a, 32'h42895ace};
test_output[380] = '{32'h429be13f};
test_index[380] = '{4};
test_input[3048:3055] = '{32'h42bf1eb0, 32'hc25bd04f, 32'hc1fa596c, 32'h42a80911, 32'h42b9ecb9, 32'hc193b9f0, 32'hc21a2954, 32'hc2181841};
test_output[381] = '{32'h42bf1eb0};
test_index[381] = '{0};
test_input[3056:3063] = '{32'hc26400ea, 32'h428d473c, 32'h4214130f, 32'h428fe1ee, 32'h427c1154, 32'hc2143715, 32'h428cd2c1, 32'hc11e390a};
test_output[382] = '{32'h428fe1ee};
test_index[382] = '{3};
test_input[3064:3071] = '{32'hc1efd96a, 32'h42506476, 32'h40ce2fc0, 32'hc228840c, 32'h427fe940, 32'hc299b2c0, 32'hc179074b, 32'hc2afbe51};
test_output[383] = '{32'h427fe940};
test_index[383] = '{4};
test_input[3072:3079] = '{32'hc2b0cef7, 32'h41054dc2, 32'h41444961, 32'hc1dddd13, 32'h4222e10d, 32'h42be29ce, 32'hc2834caf, 32'hbf99b5db};
test_output[384] = '{32'h42be29ce};
test_index[384] = '{5};
test_input[3080:3087] = '{32'h427c7962, 32'hc293457d, 32'h42afb60a, 32'h424c3140, 32'h4186033f, 32'hc21c7a4e, 32'h428a6bb7, 32'hc229a1d3};
test_output[385] = '{32'h42afb60a};
test_index[385] = '{2};
test_input[3088:3095] = '{32'h41dc783a, 32'h41b7f926, 32'hc2814342, 32'hc2a771be, 32'h42894b50, 32'h40cf154f, 32'hc28da1ef, 32'h41442cae};
test_output[386] = '{32'h42894b50};
test_index[386] = '{4};
test_input[3096:3103] = '{32'hc16441b8, 32'h42af9894, 32'hc26da170, 32'h428598e7, 32'h42910115, 32'hc1b948e1, 32'hc1f73c16, 32'h4262b425};
test_output[387] = '{32'h42af9894};
test_index[387] = '{1};
test_input[3104:3111] = '{32'hc17bb2ca, 32'h42615735, 32'h4295a67f, 32'hc11d8927, 32'hc2af01d5, 32'h418456f9, 32'h3fc91967, 32'hc275602d};
test_output[388] = '{32'h4295a67f};
test_index[388] = '{2};
test_input[3112:3119] = '{32'h4259ae9b, 32'hc2b69580, 32'hc263fa85, 32'h42ae5d03, 32'hc23ac7cd, 32'hc258aaef, 32'h3fdc42be, 32'h42a1e191};
test_output[389] = '{32'h42ae5d03};
test_index[389] = '{3};
test_input[3120:3127] = '{32'h42998a1e, 32'hc29a1b3e, 32'hc115ab22, 32'hc268f12e, 32'h4244f717, 32'h42c4bab7, 32'hc2c615f8, 32'hc0a12a1a};
test_output[390] = '{32'h42c4bab7};
test_index[390] = '{5};
test_input[3128:3135] = '{32'h428eabc7, 32'h428d92d0, 32'hc273c981, 32'h429b51dd, 32'h41afbcea, 32'h4252448d, 32'hc1f247e0, 32'h42b2fbf0};
test_output[391] = '{32'h42b2fbf0};
test_index[391] = '{7};
test_input[3136:3143] = '{32'hc2a94e4c, 32'hc1f5b51a, 32'h42aeaa20, 32'hc0091138, 32'h41a5629c, 32'h40612739, 32'h4290bf27, 32'hc269f07c};
test_output[392] = '{32'h42aeaa20};
test_index[392] = '{2};
test_input[3144:3151] = '{32'hc1967540, 32'hc1c89e9c, 32'h426af1f4, 32'hc26e4529, 32'h4205c3f3, 32'hc196b877, 32'hbf33bc75, 32'h42b00854};
test_output[393] = '{32'h42b00854};
test_index[393] = '{7};
test_input[3152:3159] = '{32'hc1fc7b8c, 32'h42452ae3, 32'hc29ef430, 32'hc1637572, 32'h418c7da1, 32'hc286bd67, 32'h428c9df1, 32'h41913991};
test_output[394] = '{32'h428c9df1};
test_index[394] = '{6};
test_input[3160:3167] = '{32'h42c40b64, 32'h425610e0, 32'h42826c04, 32'h4174f61b, 32'h42a34c23, 32'h42b9b208, 32'hc24d9581, 32'h408bcc5a};
test_output[395] = '{32'h42c40b64};
test_index[395] = '{0};
test_input[3168:3175] = '{32'hc27a79b2, 32'hc2b17904, 32'h41094f36, 32'h42a6ecab, 32'h419a3701, 32'h4178e6a4, 32'h42a9bd08, 32'h415f0e2e};
test_output[396] = '{32'h42a9bd08};
test_index[396] = '{6};
test_input[3176:3183] = '{32'h4144fd68, 32'h41430a2f, 32'h425255bd, 32'hc00ed833, 32'h41dce7e5, 32'h42904bb3, 32'h42bba332, 32'h42933d94};
test_output[397] = '{32'h42bba332};
test_index[397] = '{6};
test_input[3184:3191] = '{32'h428efc3c, 32'hc27d281a, 32'h4270dfa0, 32'h420296c8, 32'hc21d70d7, 32'hc0e15169, 32'h42b9860f, 32'h426ad173};
test_output[398] = '{32'h42b9860f};
test_index[398] = '{6};
test_input[3192:3199] = '{32'hc1e8e227, 32'hc10f2a4f, 32'h42b95a47, 32'h4084e832, 32'hc093a9b9, 32'h429a967e, 32'h427a7749, 32'hc2c7019b};
test_output[399] = '{32'h42b95a47};
test_index[399] = '{2};
test_input[3200:3207] = '{32'hc246af32, 32'h41f7302e, 32'h417d431b, 32'h41c88b9c, 32'hc2b0d84c, 32'hc2be2d92, 32'h429a5b04, 32'hc2995148};
test_output[400] = '{32'h429a5b04};
test_index[400] = '{6};
test_input[3208:3215] = '{32'h4296e292, 32'h428f8cd5, 32'h42125aa3, 32'hc269951d, 32'hc2806b72, 32'hc2bdd052, 32'hc23b9151, 32'h412f4bd0};
test_output[401] = '{32'h4296e292};
test_index[401] = '{0};
test_input[3216:3223] = '{32'h41b0369b, 32'h42c49165, 32'h42bd0611, 32'hc2348faf, 32'hc294e4ee, 32'hc26a1b53, 32'hc1e5cefc, 32'h4024417a};
test_output[402] = '{32'h42c49165};
test_index[402] = '{1};
test_input[3224:3231] = '{32'h42a4c78b, 32'hc0e942d4, 32'hc28e9cd0, 32'h42a35565, 32'h408730f8, 32'hc1c67549, 32'hc20cce51, 32'h42a700b4};
test_output[403] = '{32'h42a700b4};
test_index[403] = '{7};
test_input[3232:3239] = '{32'hc231a871, 32'hc22cc57e, 32'h40b87eed, 32'hc2c1e94e, 32'hc257afb2, 32'hc2b202a7, 32'h405345de, 32'hc23e903e};
test_output[404] = '{32'h40b87eed};
test_index[404] = '{2};
test_input[3240:3247] = '{32'h3fae174b, 32'h42b29ec0, 32'h42c062b3, 32'h4293b40a, 32'h41768324, 32'hc2bbd968, 32'h4290bcfb, 32'h42c7ebab};
test_output[405] = '{32'h42c7ebab};
test_index[405] = '{7};
test_input[3248:3255] = '{32'hc28d6f3c, 32'h4200d852, 32'h4268a1db, 32'h428aeeaa, 32'hc2ae3d7b, 32'hc2869fe1, 32'hc293e540, 32'h42bb1a97};
test_output[406] = '{32'h42bb1a97};
test_index[406] = '{7};
test_input[3256:3263] = '{32'hc269e7f0, 32'h42b01f43, 32'h4187d5fc, 32'hc23e5466, 32'h42abd3e7, 32'h41f7e06f, 32'h4198f3be, 32'h427bd738};
test_output[407] = '{32'h42b01f43};
test_index[407] = '{1};
test_input[3264:3271] = '{32'h42200a55, 32'h42556331, 32'hc201e0e7, 32'hc209683e, 32'hc184bee7, 32'hc2a97a5c, 32'h411e9c31, 32'hc1ad19f6};
test_output[408] = '{32'h42556331};
test_index[408] = '{1};
test_input[3272:3279] = '{32'h40dce4bc, 32'h418f7cae, 32'h409dbbbe, 32'hc2084e2e, 32'hc1d69f38, 32'h421e99df, 32'hc25b21ec, 32'h4217b563};
test_output[409] = '{32'h421e99df};
test_index[409] = '{5};
test_input[3280:3287] = '{32'hc1e40caf, 32'h42b8a524, 32'h42ad206e, 32'h420dbf90, 32'h40935b72, 32'h418957ee, 32'h420e0889, 32'hc29f0e9c};
test_output[410] = '{32'h42b8a524};
test_index[410] = '{1};
test_input[3288:3295] = '{32'h42aa04d6, 32'h426bcdc9, 32'hc1e40092, 32'h41b9190d, 32'h4220da39, 32'hc28ad476, 32'h42c29dd9, 32'hc0932c38};
test_output[411] = '{32'h42c29dd9};
test_index[411] = '{6};
test_input[3296:3303] = '{32'h4231fdba, 32'hc2b6be0a, 32'hc2a7bd50, 32'hc1f18aa6, 32'h4131317d, 32'hc035d833, 32'hc1dca2df, 32'h41843a3f};
test_output[412] = '{32'h4231fdba};
test_index[412] = '{0};
test_input[3304:3311] = '{32'h42acb36e, 32'hc1b34216, 32'hc24459d7, 32'h424080d0, 32'h40b5f17d, 32'h424653d4, 32'h42131eb7, 32'h424f6cec};
test_output[413] = '{32'h42acb36e};
test_index[413] = '{0};
test_input[3312:3319] = '{32'h428d0954, 32'h4215675f, 32'h42870d29, 32'hc2782adc, 32'hc2ac38a9, 32'h420ceb28, 32'h42b7a9eb, 32'hc2a4169e};
test_output[414] = '{32'h42b7a9eb};
test_index[414] = '{6};
test_input[3320:3327] = '{32'h4231fb06, 32'h42a808c5, 32'h41c983e1, 32'h423f9c08, 32'hc234d461, 32'h421798f1, 32'h425c07b0, 32'hc245f282};
test_output[415] = '{32'h42a808c5};
test_index[415] = '{1};
test_input[3328:3335] = '{32'hc29d4872, 32'hc2ae8eb6, 32'hc12590b5, 32'h41f874f3, 32'hc2ad2326, 32'hc291d3f9, 32'hc2987312, 32'hc208d579};
test_output[416] = '{32'h41f874f3};
test_index[416] = '{3};
test_input[3336:3343] = '{32'hc2a41817, 32'hc1f62fad, 32'hc21268ea, 32'h42bce576, 32'hc2897fde, 32'hc2aaae73, 32'hc2bfd0a5, 32'hc287eaa8};
test_output[417] = '{32'h42bce576};
test_index[417] = '{3};
test_input[3344:3351] = '{32'hc27e6b89, 32'h428ce34f, 32'hc1edeb5f, 32'hc2bd8dac, 32'hc2385cef, 32'hbfb763c7, 32'h414e6f1b, 32'h42aacdf9};
test_output[418] = '{32'h42aacdf9};
test_index[418] = '{7};
test_input[3352:3359] = '{32'hc223e26a, 32'hc2105db0, 32'h414dd97c, 32'h4289025a, 32'hc23edadf, 32'hc243425a, 32'hc27bae43, 32'hc2ad58f8};
test_output[419] = '{32'h4289025a};
test_index[419] = '{3};
test_input[3360:3367] = '{32'hc279815f, 32'hc23250af, 32'hc01be36d, 32'hc2c49839, 32'h42612b62, 32'hc2c10be2, 32'h424d2895, 32'h42a6d25a};
test_output[420] = '{32'h42a6d25a};
test_index[420] = '{7};
test_input[3368:3375] = '{32'hbee419d2, 32'h4106bb2b, 32'hc12a849d, 32'h427d5933, 32'hc2b1beba, 32'hc243d258, 32'h4279ae75, 32'h42465259};
test_output[421] = '{32'h427d5933};
test_index[421] = '{3};
test_input[3376:3383] = '{32'h412bf679, 32'h42ba568b, 32'h42894f64, 32'h419e0e8a, 32'hc25ad203, 32'hc1981a93, 32'hc1cd2e3e, 32'h4267b265};
test_output[422] = '{32'h42ba568b};
test_index[422] = '{1};
test_input[3384:3391] = '{32'hc1c50226, 32'h41312557, 32'hc26f1f9f, 32'hc2042d30, 32'hc2c7ae4c, 32'h40e4f5fd, 32'hc05fb08f, 32'hc1ec2f07};
test_output[423] = '{32'h41312557};
test_index[423] = '{1};
test_input[3392:3399] = '{32'hc1dbc4b1, 32'h42aae14b, 32'h4289e77f, 32'hc28c83da, 32'h41e4e089, 32'hc20d7ba6, 32'h41faa3b0, 32'hc24560eb};
test_output[424] = '{32'h42aae14b};
test_index[424] = '{1};
test_input[3400:3407] = '{32'h42b58e5f, 32'hc147e973, 32'hc2b8e99f, 32'hc289055a, 32'h4255605c, 32'hc231dd5f, 32'h425b15ef, 32'hc179f830};
test_output[425] = '{32'h42b58e5f};
test_index[425] = '{0};
test_input[3408:3415] = '{32'hc0af9d59, 32'h41a47268, 32'hc2a9f3da, 32'hc0657475, 32'hc297de89, 32'hc240e54d, 32'hc0583f87, 32'hc120273f};
test_output[426] = '{32'h41a47268};
test_index[426] = '{1};
test_input[3416:3423] = '{32'h41f9bc6d, 32'h42784a07, 32'hc0a65e2f, 32'h42bb5ae2, 32'h426d4c13, 32'hc08f8e5f, 32'hc19ced48, 32'h41a6abcf};
test_output[427] = '{32'h42bb5ae2};
test_index[427] = '{3};
test_input[3424:3431] = '{32'hc20c209c, 32'h41c0ba41, 32'hc125d16d, 32'hc275345d, 32'hc16bb0f8, 32'h42bd4d8f, 32'hc298ec40, 32'hc2a9b53f};
test_output[428] = '{32'h42bd4d8f};
test_index[428] = '{5};
test_input[3432:3439] = '{32'h425205fa, 32'h42a6e25f, 32'h42b5d1cd, 32'h42859539, 32'hc2a4e559, 32'hc2319bf8, 32'h42a7f129, 32'hc2bf9549};
test_output[429] = '{32'h42b5d1cd};
test_index[429] = '{2};
test_input[3440:3447] = '{32'h42afea9f, 32'hc2a35faa, 32'hc2ab13a5, 32'hc1939dc0, 32'h41ad30f4, 32'hc22cd060, 32'h40a687be, 32'h404aa259};
test_output[430] = '{32'h42afea9f};
test_index[430] = '{0};
test_input[3448:3455] = '{32'h41d38440, 32'h429e2a70, 32'h42c7ce60, 32'h42ba8a01, 32'h42388cde, 32'hc26e5ecb, 32'h42c6dfca, 32'hc2bc9b64};
test_output[431] = '{32'h42c7ce60};
test_index[431] = '{2};
test_input[3456:3463] = '{32'hc2822134, 32'hc1a89246, 32'h42905ed0, 32'h424233e1, 32'hc19c2c06, 32'h4266d94d, 32'hc1d84820, 32'h42b8a241};
test_output[432] = '{32'h42b8a241};
test_index[432] = '{7};
test_input[3464:3471] = '{32'h42a8cc60, 32'hc0136af2, 32'h41f17508, 32'h427f217b, 32'hc27b6fdd, 32'hc14f0a46, 32'h423fae4f, 32'hc1fedde3};
test_output[433] = '{32'h42a8cc60};
test_index[433] = '{0};
test_input[3472:3479] = '{32'h42231288, 32'hc0b4d04d, 32'h423b456d, 32'h42149a2b, 32'hc2523ea6, 32'h424c7193, 32'hbdbf44af, 32'hc19f279b};
test_output[434] = '{32'h424c7193};
test_index[434] = '{5};
test_input[3480:3487] = '{32'hc20597f5, 32'hc2776280, 32'hc2c15f56, 32'hc0e73e6e, 32'hc1be5f73, 32'h42abf303, 32'h424259b5, 32'h42adba97};
test_output[435] = '{32'h42adba97};
test_index[435] = '{7};
test_input[3488:3495] = '{32'h4261110b, 32'hc2546734, 32'hc2567dae, 32'h42b4b28b, 32'hc2729674, 32'hc24e7acb, 32'hc1c9812f, 32'h42c3c354};
test_output[436] = '{32'h42c3c354};
test_index[436] = '{7};
test_input[3496:3503] = '{32'h42a1ea47, 32'h4197b663, 32'hc2bbeff8, 32'h42aaf4f0, 32'hc29326c2, 32'hc2be71a1, 32'hc236ec3f, 32'hc1ae8a3d};
test_output[437] = '{32'h42aaf4f0};
test_index[437] = '{3};
test_input[3504:3511] = '{32'h4236dfd2, 32'h4284bc22, 32'hc1bd9b8b, 32'hc21d2b4f, 32'h4240e47c, 32'h42c3b83a, 32'h42316592, 32'hc1b2616c};
test_output[438] = '{32'h42c3b83a};
test_index[438] = '{5};
test_input[3512:3519] = '{32'hc294dee6, 32'hc1a584b3, 32'h429ca8b3, 32'hc262f827, 32'hc20295a0, 32'h429d99d3, 32'hc226e831, 32'hc243a91f};
test_output[439] = '{32'h429d99d3};
test_index[439] = '{5};
test_input[3520:3527] = '{32'h42731f6c, 32'h42af25f7, 32'h420a6d13, 32'h429a5e6f, 32'h425b273d, 32'h42bae1ef, 32'h41041eba, 32'h42707cca};
test_output[440] = '{32'h42bae1ef};
test_index[440] = '{5};
test_input[3528:3535] = '{32'hc17c7a59, 32'hc2107c2c, 32'h41deb923, 32'h42531697, 32'hc161b6ef, 32'hc1ddc81f, 32'h42129772, 32'h4286bf69};
test_output[441] = '{32'h4286bf69};
test_index[441] = '{7};
test_input[3536:3543] = '{32'hc1f57f3c, 32'h428ed9b7, 32'h4291c865, 32'h413ee22c, 32'hc1c731da, 32'hc2b15d1c, 32'hc28a1530, 32'h42bcd08a};
test_output[442] = '{32'h42bcd08a};
test_index[442] = '{7};
test_input[3544:3551] = '{32'h42c216eb, 32'hc29a9d60, 32'hc2c15d6b, 32'hc21b8db3, 32'hc000757c, 32'h42bdae0b, 32'hc2b4dfcf, 32'h420e3417};
test_output[443] = '{32'h42c216eb};
test_index[443] = '{0};
test_input[3552:3559] = '{32'h405b38b2, 32'h42526c13, 32'hc261fe55, 32'h42b469b0, 32'hc295535a, 32'hc0b0813f, 32'hc2c4c996, 32'h42992df7};
test_output[444] = '{32'h42b469b0};
test_index[444] = '{3};
test_input[3560:3567] = '{32'hc2a0e3b8, 32'hc1a81439, 32'hc1c7a438, 32'hc228f539, 32'h422c713c, 32'h4291bc0d, 32'h423d6a5a, 32'h4195b9b1};
test_output[445] = '{32'h4291bc0d};
test_index[445] = '{5};
test_input[3568:3575] = '{32'hc29b0188, 32'hc22cdd88, 32'h42a49474, 32'hc2b5ce4b, 32'hc1523deb, 32'h41c41fc6, 32'hc23e572f, 32'h41bf1e70};
test_output[446] = '{32'h42a49474};
test_index[446] = '{2};
test_input[3576:3583] = '{32'h41d5725b, 32'hc2c0ccb1, 32'hc182b838, 32'h427f139d, 32'h42c0a9ae, 32'hc1bdb726, 32'hc25dea47, 32'h42a57bd9};
test_output[447] = '{32'h42c0a9ae};
test_index[447] = '{4};
test_input[3584:3591] = '{32'h41a9efa0, 32'hc28e298d, 32'hc2b3d332, 32'h42b53f4c, 32'hc1314769, 32'hc2668501, 32'hc269dba4, 32'hc23d5007};
test_output[448] = '{32'h42b53f4c};
test_index[448] = '{3};
test_input[3592:3599] = '{32'hc27fc8f1, 32'h40d6fea0, 32'hc24074c5, 32'h419f331e, 32'h41f85ae8, 32'hc2b9b90c, 32'hc14522db, 32'h420d6aee};
test_output[449] = '{32'h420d6aee};
test_index[449] = '{7};
test_input[3600:3607] = '{32'hc1853db9, 32'hc28c7490, 32'h426c534b, 32'h40d776f1, 32'hc2a1f263, 32'hc1ee43c0, 32'h4068091e, 32'h428b7e0b};
test_output[450] = '{32'h428b7e0b};
test_index[450] = '{7};
test_input[3608:3615] = '{32'h419ac530, 32'hc2738f85, 32'hc290b9c8, 32'h42bf7968, 32'hbf1d515f, 32'hc245337a, 32'h41503509, 32'hc2a17017};
test_output[451] = '{32'h42bf7968};
test_index[451] = '{3};
test_input[3616:3623] = '{32'hc2676570, 32'hc20a8032, 32'hc19eb416, 32'hc1905421, 32'hbf1bcf95, 32'h41abf58c, 32'hc2117d8c, 32'h42c7ea64};
test_output[452] = '{32'h42c7ea64};
test_index[452] = '{7};
test_input[3624:3631] = '{32'h42065c33, 32'h41696408, 32'hc2ac085b, 32'h429f81ad, 32'h4267c1fc, 32'h42c4f97d, 32'hc21a419a, 32'hc1b1d4cf};
test_output[453] = '{32'h42c4f97d};
test_index[453] = '{5};
test_input[3632:3639] = '{32'h428f06ae, 32'h40cca98a, 32'hc296b8da, 32'hc22e7aaf, 32'hc2848d2e, 32'h422c2f36, 32'h426eca5b, 32'h42a97793};
test_output[454] = '{32'h42a97793};
test_index[454] = '{7};
test_input[3640:3647] = '{32'hc1c71405, 32'hc2b7be84, 32'h416fdf0f, 32'h42bbbf2c, 32'hc1d7fb9b, 32'h41529061, 32'h41df2490, 32'h41ee46e2};
test_output[455] = '{32'h42bbbf2c};
test_index[455] = '{3};
test_input[3648:3655] = '{32'h421ea1f3, 32'hc29c4787, 32'h42ae8240, 32'h429fe3ec, 32'h42c16dd1, 32'h421700b9, 32'hc1cfce84, 32'h4269b8be};
test_output[456] = '{32'h42c16dd1};
test_index[456] = '{4};
test_input[3656:3663] = '{32'h42c718a5, 32'hc21e37c9, 32'hc1b4c8f1, 32'hc0c47577, 32'hc184e47f, 32'h41b6d653, 32'h42a7cd4c, 32'h4250bf70};
test_output[457] = '{32'h42c718a5};
test_index[457] = '{0};
test_input[3664:3671] = '{32'h40a9478d, 32'h42ba2458, 32'hc2244434, 32'hc29ed868, 32'h420c5d14, 32'hc22e3dfe, 32'hc295aa32, 32'h414731b3};
test_output[458] = '{32'h42ba2458};
test_index[458] = '{1};
test_input[3672:3679] = '{32'h4227d5d4, 32'h42a65b50, 32'hc284937e, 32'h42916f0b, 32'hc1ecface, 32'h42962511, 32'h428702ae, 32'h42722046};
test_output[459] = '{32'h42a65b50};
test_index[459] = '{1};
test_input[3680:3687] = '{32'hc28be9b3, 32'hc1cbf648, 32'h41d98bd0, 32'h41a61826, 32'hc279f43e, 32'h42953bd3, 32'hc29fa171, 32'hc20cffe0};
test_output[460] = '{32'h42953bd3};
test_index[460] = '{5};
test_input[3688:3695] = '{32'hc2b42085, 32'h408550f8, 32'hc237073a, 32'h4285b138, 32'hc2bf7b40, 32'hc250213e, 32'h4202be77, 32'hc0b183f2};
test_output[461] = '{32'h4285b138};
test_index[461] = '{3};
test_input[3696:3703] = '{32'h421fbd61, 32'h421737eb, 32'h428fd3a5, 32'h429a0bc5, 32'h41f7fcbf, 32'hc282dfdb, 32'h4220fc8e, 32'h422e6972};
test_output[462] = '{32'h429a0bc5};
test_index[462] = '{3};
test_input[3704:3711] = '{32'hc29ef006, 32'hc2007819, 32'h4210663e, 32'hc22fb399, 32'hc2aaf04f, 32'h428d74af, 32'h42af08b0, 32'h426a0ad6};
test_output[463] = '{32'h42af08b0};
test_index[463] = '{6};
test_input[3712:3719] = '{32'h42aee39c, 32'h41821c7b, 32'hc2941ecf, 32'hc2b5cbb2, 32'hc19dddc6, 32'hc1f06ee1, 32'h422a01f8, 32'h4092ffa2};
test_output[464] = '{32'h42aee39c};
test_index[464] = '{0};
test_input[3720:3727] = '{32'h42c254cb, 32'h4123705b, 32'h42c0a69c, 32'h425d8f77, 32'hc2bca3e5, 32'h41a98fb8, 32'hc2aab6f5, 32'hc2b5820d};
test_output[465] = '{32'h42c254cb};
test_index[465] = '{0};
test_input[3728:3735] = '{32'h42c10261, 32'h423935c9, 32'hc1ac4a5e, 32'h4268eeec, 32'h40a89f6e, 32'hc0bfdd65, 32'hc288aee7, 32'hc247ec3a};
test_output[466] = '{32'h42c10261};
test_index[466] = '{0};
test_input[3736:3743] = '{32'hc22a4cc7, 32'h42ae88c7, 32'hc29d512f, 32'hc206d314, 32'hc223f037, 32'h42391a72, 32'hc2698796, 32'h40b55c1c};
test_output[467] = '{32'h42ae88c7};
test_index[467] = '{1};
test_input[3744:3751] = '{32'h428fd46c, 32'h42b97f52, 32'h42862afc, 32'h42899c2a, 32'h40d347f7, 32'hc1fb0a71, 32'hc22ee215, 32'hc0f9dcb0};
test_output[468] = '{32'h42b97f52};
test_index[468] = '{1};
test_input[3752:3759] = '{32'h41a50ba2, 32'hc1d51918, 32'h42073c63, 32'hc25ceaa1, 32'hc20a7ff0, 32'h42ab1407, 32'hc18fb054, 32'h42bf2b30};
test_output[469] = '{32'h42bf2b30};
test_index[469] = '{7};
test_input[3760:3767] = '{32'h42bbb71e, 32'hc2518e29, 32'h3e9cb97a, 32'h4120541f, 32'hc2c396a3, 32'h42695e7a, 32'hc2c5fd73, 32'h421f515a};
test_output[470] = '{32'h42bbb71e};
test_index[470] = '{0};
test_input[3768:3775] = '{32'hc291d8f0, 32'hc20ed4f2, 32'hc2be7aa3, 32'hc0a1644b, 32'h429360a9, 32'h4223daeb, 32'h42c55cda, 32'hc2c5b78b};
test_output[471] = '{32'h42c55cda};
test_index[471] = '{6};
test_input[3776:3783] = '{32'h42267663, 32'h413312f7, 32'hc2924999, 32'hc2a188d2, 32'h4294cdd7, 32'h4234cfa7, 32'hc291bd27, 32'hc13eb46e};
test_output[472] = '{32'h4294cdd7};
test_index[472] = '{4};
test_input[3784:3791] = '{32'h413cf58b, 32'hc29a7ec1, 32'hc1a59890, 32'h428b0924, 32'hc2adf4f5, 32'hc0f48516, 32'h4270a9e9, 32'hc2b8df95};
test_output[473] = '{32'h428b0924};
test_index[473] = '{3};
test_input[3792:3799] = '{32'h42897a3e, 32'hbe6355b6, 32'h42b58494, 32'h4296f4f2, 32'hc2c6ad8d, 32'hc2782fc6, 32'hc29bda92, 32'h418c7de0};
test_output[474] = '{32'h42b58494};
test_index[474] = '{2};
test_input[3800:3807] = '{32'h40dac38e, 32'hc28593ca, 32'hc18b00ba, 32'h4155d24d, 32'h428f8f55, 32'h42b68fc9, 32'h4226a472, 32'hc0b4c017};
test_output[475] = '{32'h42b68fc9};
test_index[475] = '{5};
test_input[3808:3815] = '{32'h420a75d4, 32'h42bc93d1, 32'h42ba345b, 32'h406f15e4, 32'h4183c160, 32'hc090ee91, 32'hc27f462b, 32'h41a0ff1f};
test_output[476] = '{32'h42bc93d1};
test_index[476] = '{1};
test_input[3816:3823] = '{32'hc233e484, 32'hc2a5a820, 32'hc134a222, 32'h41516dff, 32'h4291961e, 32'hc2b042be, 32'h41e8415c, 32'h42beb53e};
test_output[477] = '{32'h42beb53e};
test_index[477] = '{7};
test_input[3824:3831] = '{32'hc251ebd5, 32'h42190dec, 32'h425f39f0, 32'h4200a21d, 32'h420f8465, 32'h4261eca4, 32'h41d3fbcd, 32'h42a088fe};
test_output[478] = '{32'h42a088fe};
test_index[478] = '{7};
test_input[3832:3839] = '{32'hc299d41d, 32'h41bd2ad5, 32'h415e2954, 32'h42c3489a, 32'h4164528e, 32'hc21950a1, 32'hc0e86f76, 32'h41c9949d};
test_output[479] = '{32'h42c3489a};
test_index[479] = '{3};
test_input[3840:3847] = '{32'hc1fcb46e, 32'h41bee961, 32'hc15d7db3, 32'h42b5b4b8, 32'h4293eb55, 32'hc2a2b264, 32'hc26f3e74, 32'hc2a9bc28};
test_output[480] = '{32'h42b5b4b8};
test_index[480] = '{3};
test_input[3848:3855] = '{32'h4275edc2, 32'hbe644ed5, 32'hc246a094, 32'h42b5b4e3, 32'h42c48716, 32'hc2181b30, 32'hc129c82f, 32'h41f6ded0};
test_output[481] = '{32'h42c48716};
test_index[481] = '{4};
test_input[3856:3863] = '{32'hc26c49b9, 32'hc0c87a48, 32'h41569a6c, 32'hc20c31e5, 32'h42c67e80, 32'h41d130f3, 32'hc255a9fb, 32'hc2b88607};
test_output[482] = '{32'h42c67e80};
test_index[482] = '{4};
test_input[3864:3871] = '{32'hc24c718c, 32'h4220909b, 32'h3ffb153a, 32'hc276d79c, 32'h3fd050d5, 32'hc278f567, 32'hc0a01168, 32'hc292bba6};
test_output[483] = '{32'h4220909b};
test_index[483] = '{1};
test_input[3872:3879] = '{32'h417f771c, 32'h42a71634, 32'hc28bed16, 32'h42a003ed, 32'hc2b91d7b, 32'h41144c22, 32'hc1d96039, 32'h42a374d3};
test_output[484] = '{32'h42a71634};
test_index[484] = '{1};
test_input[3880:3887] = '{32'h42939097, 32'hc2820009, 32'hc24d71b7, 32'hc18f1bdc, 32'hc27fdaf3, 32'hc268f4be, 32'hc0fe8cb4, 32'hc2438067};
test_output[485] = '{32'h42939097};
test_index[485] = '{0};
test_input[3888:3895] = '{32'h42bd82cc, 32'hc2b14bd1, 32'hc1fa6d54, 32'h41f1e72c, 32'hc12e6aad, 32'hc2b432ca, 32'hc28527e4, 32'h417ffdf4};
test_output[486] = '{32'h42bd82cc};
test_index[486] = '{0};
test_input[3896:3903] = '{32'h42c22385, 32'h428ba93b, 32'h41d07c1c, 32'h4249d26a, 32'h41fb246e, 32'h422a80d7, 32'h42bc8038, 32'hc2c52c8c};
test_output[487] = '{32'h42c22385};
test_index[487] = '{0};
test_input[3904:3911] = '{32'h42c72fbb, 32'h42a04d9f, 32'hc2881065, 32'hc24db7ba, 32'h41615951, 32'h4097c1d9, 32'h40a6b8cf, 32'hc2997fd5};
test_output[488] = '{32'h42c72fbb};
test_index[488] = '{0};
test_input[3912:3919] = '{32'hc2c6eb68, 32'hc1f01e25, 32'hc1cf2332, 32'hc1f4f5a2, 32'hc2465ce4, 32'h41a9d203, 32'h4126880f, 32'hc2ac9cb6};
test_output[489] = '{32'h41a9d203};
test_index[489] = '{5};
test_input[3920:3927] = '{32'hc28d771a, 32'h42b92f4f, 32'h421f59cb, 32'hc209e407, 32'h4200fffc, 32'hbebb5356, 32'h416ec71d, 32'h42918dd2};
test_output[490] = '{32'h42b92f4f};
test_index[490] = '{1};
test_input[3928:3935] = '{32'hc02db271, 32'hc2a52605, 32'h427a4c81, 32'hc1a9884a, 32'hc1cc8918, 32'hc2a14175, 32'h42084f3f, 32'h42ae0fc7};
test_output[491] = '{32'h42ae0fc7};
test_index[491] = '{7};
test_input[3936:3943] = '{32'h428c6ae8, 32'hc26211fd, 32'h413aef16, 32'h4283fde1, 32'h428ec35a, 32'hc26ea062, 32'hc196fc3d, 32'h41b6989b};
test_output[492] = '{32'h428ec35a};
test_index[492] = '{4};
test_input[3944:3951] = '{32'h3cf046a1, 32'hc2bf48ef, 32'h41c032d0, 32'h4284e118, 32'hc1929413, 32'h413702ba, 32'h429990df, 32'hc1b602a9};
test_output[493] = '{32'h429990df};
test_index[493] = '{6};
test_input[3952:3959] = '{32'h419043fe, 32'h421ac7fd, 32'hc1ea28bc, 32'hc21ee8e9, 32'hc2acd432, 32'h41ff2fa9, 32'h41e3c262, 32'h42a6de78};
test_output[494] = '{32'h42a6de78};
test_index[494] = '{7};
test_input[3960:3967] = '{32'hc1b5b316, 32'hbfb8d644, 32'hc2a5808c, 32'h42440cdf, 32'h4258cea0, 32'h419cd80a, 32'h41dc86f0, 32'hc26ea593};
test_output[495] = '{32'h4258cea0};
test_index[495] = '{4};
test_input[3968:3975] = '{32'hc09a3219, 32'hc2ac699c, 32'hc1dd7b61, 32'hc28b42c6, 32'h4233a3c8, 32'hc25454cc, 32'h42693e9d, 32'h420da672};
test_output[496] = '{32'h42693e9d};
test_index[496] = '{6};
test_input[3976:3983] = '{32'hc2b20fb6, 32'h41796e8b, 32'h4289a7d4, 32'h42a86edd, 32'h3f110a90, 32'h41d58530, 32'h4138d73b, 32'hc1c2bf70};
test_output[497] = '{32'h42a86edd};
test_index[497] = '{3};
test_input[3984:3991] = '{32'hc25373e7, 32'hc18a632b, 32'h40bbfb20, 32'h4260ec74, 32'hc1da34f3, 32'hc0f053b6, 32'hc2c45d31, 32'h41838f1c};
test_output[498] = '{32'h4260ec74};
test_index[498] = '{3};
test_input[3992:3999] = '{32'hc263145d, 32'hc2862c83, 32'hc28a8172, 32'hc186946b, 32'h4286d230, 32'hc2361770, 32'h42402064, 32'hc2973c5b};
test_output[499] = '{32'h4286d230};
test_index[499] = '{4};
test_input[4000:4007] = '{32'h3ef0ee80, 32'h41f467e2, 32'h418c980e, 32'hc1c977c2, 32'hc1fd2ccc, 32'h40dd147d, 32'h42c4a9f9, 32'hc20ebe95};
test_output[500] = '{32'h42c4a9f9};
test_index[500] = '{6};
test_input[4008:4015] = '{32'hc2652804, 32'h422ebcf7, 32'h42718623, 32'h42b4b397, 32'hc23aa497, 32'hc2bbfc0f, 32'hc279f640, 32'h40d375d0};
test_output[501] = '{32'h42b4b397};
test_index[501] = '{3};
test_input[4016:4023] = '{32'hc1113868, 32'h425a40a2, 32'hc28b3dfe, 32'h417561e2, 32'h41e9261e, 32'hc276a5ff, 32'hc2190185, 32'hc14d5a78};
test_output[502] = '{32'h425a40a2};
test_index[502] = '{1};
test_input[4024:4031] = '{32'h4295c5ec, 32'h42bfe414, 32'h41dc5858, 32'h41cfb44e, 32'hc28f6696, 32'h429eb7bd, 32'h416e3e0a, 32'hc19b7740};
test_output[503] = '{32'h42bfe414};
test_index[503] = '{1};
test_input[4032:4039] = '{32'hc21bbc2b, 32'hc2b444ba, 32'hc2038180, 32'hc26ed0c8, 32'h4257af61, 32'h421102c9, 32'h41b7b2d3, 32'hc2960b32};
test_output[504] = '{32'h4257af61};
test_index[504] = '{4};
test_input[4040:4047] = '{32'hc1e6c724, 32'h428280b2, 32'hc16105a7, 32'h408fcdf1, 32'h424945f8, 32'hc20efcd7, 32'h42adf07f, 32'h412dde8e};
test_output[505] = '{32'h42adf07f};
test_index[505] = '{6};
test_input[4048:4055] = '{32'hc23155c3, 32'h42597197, 32'h42b5a77a, 32'h428d9dc1, 32'hc28eb89d, 32'hc2c40919, 32'h41c07c70, 32'hc28cb637};
test_output[506] = '{32'h42b5a77a};
test_index[506] = '{2};
test_input[4056:4063] = '{32'hc18e5d2c, 32'h41a45ff1, 32'h4254d641, 32'h425ab526, 32'hc2b2dd83, 32'h42a2861c, 32'h424a7cfe, 32'hc2a0d70e};
test_output[507] = '{32'h42a2861c};
test_index[507] = '{5};
test_input[4064:4071] = '{32'hc2933626, 32'h4291ed26, 32'h4259cddf, 32'hc28b25b6, 32'hc2711998, 32'h41754985, 32'hc0da8c61, 32'h41dd62e5};
test_output[508] = '{32'h4291ed26};
test_index[508] = '{1};
test_input[4072:4079] = '{32'h429044fc, 32'h421b82f2, 32'hc1814938, 32'hc1d929bf, 32'hc15152c1, 32'hc2c47b27, 32'hc2c758cf, 32'h420eeda5};
test_output[509] = '{32'h429044fc};
test_index[509] = '{0};
test_input[4080:4087] = '{32'hc27044f2, 32'h413850d1, 32'h423faead, 32'hc2a801b7, 32'h4272a34c, 32'h42a1c2a5, 32'hc28a4b34, 32'h42ac03e7};
test_output[510] = '{32'h42ac03e7};
test_index[510] = '{7};
test_input[4088:4095] = '{32'h40c23a1d, 32'hc1a090c2, 32'hc2bb3e81, 32'hc27dbb79, 32'hc23d4085, 32'h40fe1aed, 32'hc1f8d081, 32'h42739af4};
test_output[511] = '{32'h42739af4};
test_index[511] = '{7};
test_input[4096:4103] = '{32'h4227a776, 32'h425524ea, 32'h42c65877, 32'hc1acd3e6, 32'h422e7f0c, 32'hc2433da5, 32'h414c8106, 32'hc09acc15};
test_output[512] = '{32'h42c65877};
test_index[512] = '{2};
test_input[4104:4111] = '{32'h41735ad0, 32'hc1df7826, 32'h41407aa7, 32'h422859b1, 32'h428b9bc5, 32'hc2673a35, 32'h4104e729, 32'h41a208e0};
test_output[513] = '{32'h428b9bc5};
test_index[513] = '{4};
test_input[4112:4119] = '{32'h426b835a, 32'hc1b2c71e, 32'h41a0923f, 32'hc2a00a27, 32'hc2b5af47, 32'hc2b86635, 32'hc1ca6424, 32'hc220de24};
test_output[514] = '{32'h426b835a};
test_index[514] = '{0};
test_input[4120:4127] = '{32'h41f2a051, 32'h427cb6b5, 32'h41be7c24, 32'hc17ca47b, 32'hc1de517a, 32'hc000cd68, 32'hc01f5174, 32'hc19e667e};
test_output[515] = '{32'h427cb6b5};
test_index[515] = '{1};
test_input[4128:4135] = '{32'hc23a49d8, 32'h428cfb7a, 32'h42101c5b, 32'h421fb6cb, 32'h421b3925, 32'hc2923394, 32'hc2ad2f43, 32'h4169c5cf};
test_output[516] = '{32'h428cfb7a};
test_index[516] = '{1};
test_input[4136:4143] = '{32'hc24730de, 32'h428ab287, 32'h4219f9f2, 32'hc1057ca8, 32'hc2a35eeb, 32'hc21ba695, 32'h40fd2ec9, 32'hc28ee82d};
test_output[517] = '{32'h428ab287};
test_index[517] = '{1};
test_input[4144:4151] = '{32'hc1f0cae0, 32'hbfaae2cd, 32'hc270d12f, 32'h42c47ddb, 32'h41815905, 32'h427fd591, 32'h42c2c64e, 32'hc27b9c77};
test_output[518] = '{32'h42c47ddb};
test_index[518] = '{3};
test_input[4152:4159] = '{32'hc1847128, 32'hc134be30, 32'hbf42957b, 32'h42609c4f, 32'h42ad664b, 32'h410c7e4d, 32'h427ee6c1, 32'h4186cbff};
test_output[519] = '{32'h42ad664b};
test_index[519] = '{4};
test_input[4160:4167] = '{32'hc23958a3, 32'h3fe28a8d, 32'h4220e76f, 32'hc2a9d03e, 32'hc28e59dd, 32'h420b1f02, 32'hc224a228, 32'h42247153};
test_output[520] = '{32'h42247153};
test_index[520] = '{7};
test_input[4168:4175] = '{32'h4271be87, 32'hc24ab622, 32'h42a85092, 32'h425af912, 32'h412fe152, 32'hc2bbb472, 32'hc1817ac6, 32'h426496d7};
test_output[521] = '{32'h42a85092};
test_index[521] = '{2};
test_input[4176:4183] = '{32'h424a2c33, 32'h41dc454e, 32'h428b20e0, 32'hc2c5a4f4, 32'h420fd0cc, 32'h42b3d9aa, 32'hc281c5f3, 32'h42c5914c};
test_output[522] = '{32'h42c5914c};
test_index[522] = '{7};
test_input[4184:4191] = '{32'h42c708f0, 32'h428c2eff, 32'hc2221637, 32'h42b62fb3, 32'hc2c619f2, 32'hc26142e1, 32'hc272230d, 32'hc0bf35f8};
test_output[523] = '{32'h42c708f0};
test_index[523] = '{0};
test_input[4192:4199] = '{32'hc2bc9e89, 32'hc2a5446e, 32'h4285a752, 32'h427706de, 32'hc289ce25, 32'hc280881f, 32'h41985f2f, 32'h41e93d12};
test_output[524] = '{32'h4285a752};
test_index[524] = '{2};
test_input[4200:4207] = '{32'h420d8c1e, 32'hc201fff3, 32'hc1c62bbf, 32'hc2a0d5b7, 32'hc25c14c0, 32'hc2564a25, 32'h4133a676, 32'h42b69bbe};
test_output[525] = '{32'h42b69bbe};
test_index[525] = '{7};
test_input[4208:4215] = '{32'h42823628, 32'hc1dbf48d, 32'hc12cd617, 32'hc2a171a8, 32'h424e9e79, 32'h42b4d5fb, 32'hc286508d, 32'h41a6704c};
test_output[526] = '{32'h42b4d5fb};
test_index[526] = '{5};
test_input[4216:4223] = '{32'h42b7cebe, 32'hc227e5f5, 32'hc27d3556, 32'hc1ce8c24, 32'hc1af2405, 32'hbfafaaa5, 32'hc2a88e23, 32'hc2016768};
test_output[527] = '{32'h42b7cebe};
test_index[527] = '{0};
test_input[4224:4231] = '{32'h42ab3871, 32'h42434d69, 32'h42a9aafd, 32'hc2502176, 32'hc2bd4adc, 32'hc22722a0, 32'hc2681afd, 32'hc2188b0f};
test_output[528] = '{32'h42ab3871};
test_index[528] = '{0};
test_input[4232:4239] = '{32'hc296e26e, 32'h42ac4af8, 32'hc26d1a24, 32'h425b6ccb, 32'h42c1f1cd, 32'h42207116, 32'h41f23935, 32'hc2ba2024};
test_output[529] = '{32'h42c1f1cd};
test_index[529] = '{4};
test_input[4240:4247] = '{32'hc2b154af, 32'h427e3ca4, 32'hc2a14912, 32'hc1b19ad0, 32'h40e88958, 32'h410189c2, 32'hc2c64288, 32'hc1ed37c4};
test_output[530] = '{32'h427e3ca4};
test_index[530] = '{1};
test_input[4248:4255] = '{32'hc04d47f7, 32'hc0cc9a80, 32'hc28dd6bc, 32'hc1320019, 32'h42a1f4cf, 32'hc293fee0, 32'hc0c56a00, 32'hc2bc22e6};
test_output[531] = '{32'h42a1f4cf};
test_index[531] = '{4};
test_input[4256:4263] = '{32'hc2ac4c71, 32'hc26b807f, 32'hc27dec24, 32'hc2445a59, 32'hc26afe58, 32'h425ebb03, 32'h3dd7e730, 32'hc17b133f};
test_output[532] = '{32'h425ebb03};
test_index[532] = '{5};
test_input[4264:4271] = '{32'h424f54b3, 32'h42b0b888, 32'hc2c4f18a, 32'h4277f799, 32'hc215f486, 32'h42122592, 32'hc299b381, 32'h42b6c9c4};
test_output[533] = '{32'h42b6c9c4};
test_index[533] = '{7};
test_input[4272:4279] = '{32'hc2147426, 32'hc1ea4d8d, 32'hc29a2d88, 32'h423ae250, 32'h42043a7b, 32'hc1881073, 32'hc1b0b1e2, 32'hc2974778};
test_output[534] = '{32'h423ae250};
test_index[534] = '{3};
test_input[4280:4287] = '{32'hc1f98ad7, 32'h42c6eda3, 32'h428791d1, 32'h42b08e8a, 32'h42aceec2, 32'hc20c188b, 32'h4253f410, 32'h4122d2be};
test_output[535] = '{32'h42c6eda3};
test_index[535] = '{1};
test_input[4288:4295] = '{32'hc10c2905, 32'h4212135a, 32'h42862b28, 32'h421633e2, 32'hc020cbad, 32'hc29ed345, 32'h42a51591, 32'hc26a9339};
test_output[536] = '{32'h42a51591};
test_index[536] = '{6};
test_input[4296:4303] = '{32'hc219f994, 32'h4290f4ad, 32'hc2208dad, 32'h4252b3e2, 32'h41797235, 32'hc21f13c4, 32'hc197ee1c, 32'hc1f0ca90};
test_output[537] = '{32'h4290f4ad};
test_index[537] = '{1};
test_input[4304:4311] = '{32'hc0446564, 32'hc259e931, 32'h41d26ae3, 32'hc24ad3fa, 32'h426c2789, 32'hbfbf40b3, 32'hc21c7f07, 32'h42adec40};
test_output[538] = '{32'h42adec40};
test_index[538] = '{7};
test_input[4312:4319] = '{32'h4214c2ef, 32'h4273227a, 32'h42a03460, 32'h42837999, 32'h42af1e15, 32'hc1a55a96, 32'h42159b3c, 32'hc172f396};
test_output[539] = '{32'h42af1e15};
test_index[539] = '{4};
test_input[4320:4327] = '{32'hc295ed96, 32'h422613d4, 32'hc23552ca, 32'h42232e76, 32'hc2a94017, 32'h4277529e, 32'h42a72df9, 32'hc07ff786};
test_output[540] = '{32'h42a72df9};
test_index[540] = '{6};
test_input[4328:4335] = '{32'h42125b48, 32'h422a5dba, 32'h4165163a, 32'h424226c6, 32'h42772ca5, 32'hc2b2247b, 32'h42c6ab3f, 32'hc23b2bf8};
test_output[541] = '{32'h42c6ab3f};
test_index[541] = '{6};
test_input[4336:4343] = '{32'h42a9406d, 32'hbfe28e75, 32'hc2ba6dcd, 32'hc2af278b, 32'hc214a844, 32'hc19eb4ea, 32'hc2667550, 32'hc1324571};
test_output[542] = '{32'h42a9406d};
test_index[542] = '{0};
test_input[4344:4351] = '{32'h41a00bd7, 32'hc1f1f0a5, 32'hc2861fb8, 32'h421c86f2, 32'hc1e54c59, 32'h42351537, 32'hc222d71e, 32'h42b67e74};
test_output[543] = '{32'h42b67e74};
test_index[543] = '{7};
test_input[4352:4359] = '{32'hc1a000cc, 32'h428bb285, 32'h426db81d, 32'h42c730a5, 32'hc173ad58, 32'hc1e3e112, 32'hc25a337d, 32'hc12e8b9e};
test_output[544] = '{32'h42c730a5};
test_index[544] = '{3};
test_input[4360:4367] = '{32'hc23f1e26, 32'hc26391e4, 32'hc29cc32e, 32'h421fde2c, 32'hc28b686f, 32'hc2712d1a, 32'hc29fbe25, 32'hc214df78};
test_output[545] = '{32'h421fde2c};
test_index[545] = '{3};
test_input[4368:4375] = '{32'hc22a3288, 32'h42061c0e, 32'h42bc9304, 32'hc127164f, 32'h4295dea5, 32'hc2915214, 32'hc238bc9c, 32'h429cbd92};
test_output[546] = '{32'h42bc9304};
test_index[546] = '{2};
test_input[4376:4383] = '{32'h42a64735, 32'hc2c3df08, 32'hc2761dc9, 32'h42c0120a, 32'h3d94f7a3, 32'h41ff4a16, 32'h42beea43, 32'h42409b55};
test_output[547] = '{32'h42c0120a};
test_index[547] = '{3};
test_input[4384:4391] = '{32'h414974c3, 32'h41ec9968, 32'h42788801, 32'hc2a672e5, 32'hbfb23ed4, 32'hc2c260b5, 32'hc2a58753, 32'h4133f519};
test_output[548] = '{32'h42788801};
test_index[548] = '{2};
test_input[4392:4399] = '{32'h42c6211f, 32'h414bbb6b, 32'h410f7af0, 32'h4260485d, 32'h40ed16a6, 32'hc202a946, 32'h423c0c38, 32'h420691f3};
test_output[549] = '{32'h42c6211f};
test_index[549] = '{0};
test_input[4400:4407] = '{32'h42801ab7, 32'hc29fc4bc, 32'hc2c16692, 32'h41c39614, 32'hc1a62b21, 32'hc2b6744a, 32'hc26e01e2, 32'hc25d6543};
test_output[550] = '{32'h42801ab7};
test_index[550] = '{0};
test_input[4408:4415] = '{32'h41bbde33, 32'h42909eb4, 32'h3fb518c4, 32'h429cf55e, 32'hc1b65257, 32'h42b28183, 32'hc2b62d18, 32'hc084ed3f};
test_output[551] = '{32'h42b28183};
test_index[551] = '{5};
test_input[4416:4423] = '{32'hc2074f84, 32'hc261d69f, 32'hc2931265, 32'h41480e05, 32'h418b6680, 32'h4244772f, 32'h42b98207, 32'hc1ee869e};
test_output[552] = '{32'h42b98207};
test_index[552] = '{6};
test_input[4424:4431] = '{32'h41928c52, 32'h41b389ed, 32'hc2602e59, 32'h3f24cc73, 32'h423756e1, 32'h4224cc91, 32'h42a238d7, 32'hc296e38b};
test_output[553] = '{32'h42a238d7};
test_index[553] = '{6};
test_input[4432:4439] = '{32'h425a03a2, 32'hc2ac792f, 32'hc1edfee1, 32'hc294dd96, 32'hc2bff5af, 32'hc0b491dc, 32'h42809eee, 32'hc29cc1a7};
test_output[554] = '{32'h42809eee};
test_index[554] = '{6};
test_input[4440:4447] = '{32'hc23f8ff8, 32'h40b2db2f, 32'hc277b281, 32'h41b52cbe, 32'h411199f7, 32'h41f7652f, 32'hc2bce8fb, 32'h42279da3};
test_output[555] = '{32'h42279da3};
test_index[555] = '{7};
test_input[4448:4455] = '{32'hc1c6c0c3, 32'h4285e397, 32'hc1be81f2, 32'h414c4da2, 32'h42658b8f, 32'h429a9e2c, 32'h4235241c, 32'h421a31bb};
test_output[556] = '{32'h429a9e2c};
test_index[556] = '{5};
test_input[4456:4463] = '{32'h42a4da47, 32'h41ad0bbb, 32'h425ad543, 32'hc180dad3, 32'h429749a5, 32'h4294a7ec, 32'hc1a197f9, 32'h426055b2};
test_output[557] = '{32'h42a4da47};
test_index[557] = '{0};
test_input[4464:4471] = '{32'hc2b0b47a, 32'h41fe2522, 32'hc2aba62d, 32'h421ee6b3, 32'h41b6f235, 32'hc29da7e0, 32'hc2a871f9, 32'h42814683};
test_output[558] = '{32'h42814683};
test_index[558] = '{7};
test_input[4472:4479] = '{32'hc2c70ec0, 32'hbf14899c, 32'hc29342de, 32'h420e7fd4, 32'hc2b6f9a1, 32'h415c775a, 32'h4269ab91, 32'h415eb3bc};
test_output[559] = '{32'h4269ab91};
test_index[559] = '{6};
test_input[4480:4487] = '{32'hc2c28874, 32'hc2aec32d, 32'hc1b58ccb, 32'h4205f259, 32'h429e2550, 32'hc25d535a, 32'h42c7bd99, 32'h4296ba21};
test_output[560] = '{32'h42c7bd99};
test_index[560] = '{6};
test_input[4488:4495] = '{32'hc094b069, 32'h42b1659c, 32'hc22f6015, 32'hc2b14d1f, 32'hc26b1c34, 32'h42ab7561, 32'hc22ef0f4, 32'h424c509e};
test_output[561] = '{32'h42b1659c};
test_index[561] = '{1};
test_input[4496:4503] = '{32'h427ad229, 32'h3fe11ac9, 32'hc18853d4, 32'h414aefe0, 32'hc0667952, 32'h42a623ca, 32'hc24da69e, 32'hc2b7051d};
test_output[562] = '{32'h42a623ca};
test_index[562] = '{5};
test_input[4504:4511] = '{32'hc0d7ecaa, 32'hc1521704, 32'h42a30c5f, 32'hc277634c, 32'h420acb0e, 32'h42b215c8, 32'h42b23f85, 32'h42a71cfb};
test_output[563] = '{32'h42b23f85};
test_index[563] = '{6};
test_input[4512:4519] = '{32'hc28259fe, 32'hc239b7f2, 32'hc19e733c, 32'hc27fc627, 32'h419900e6, 32'h42bd9281, 32'hc2b20f7a, 32'hc27c1591};
test_output[564] = '{32'h42bd9281};
test_index[564] = '{5};
test_input[4520:4527] = '{32'hc2798906, 32'h423bcb43, 32'h41e5390b, 32'h420ebd5b, 32'hc295cbee, 32'hc28b7b3e, 32'h4287c18d, 32'hc28ec54e};
test_output[565] = '{32'h4287c18d};
test_index[565] = '{6};
test_input[4528:4535] = '{32'hbfa08e38, 32'hc26aa034, 32'h428be008, 32'hc28d4fee, 32'hc1119377, 32'hc1e03aa5, 32'hc28865bd, 32'h42b166e8};
test_output[566] = '{32'h42b166e8};
test_index[566] = '{7};
test_input[4536:4543] = '{32'hc1f3d592, 32'h41293d93, 32'hc25fd106, 32'h3ea810ce, 32'h4199f5ae, 32'h41f341f8, 32'h41f7e369, 32'hc295f7dc};
test_output[567] = '{32'h41f7e369};
test_index[567] = '{6};
test_input[4544:4551] = '{32'h41f20997, 32'h42023445, 32'h4251e4ef, 32'h42937a0b, 32'h4226435f, 32'hc2c161a9, 32'h42743e41, 32'hc294d52f};
test_output[568] = '{32'h42937a0b};
test_index[568] = '{3};
test_input[4552:4559] = '{32'h41f7a5e2, 32'h4193d812, 32'h42c3ff4d, 32'h42a8495c, 32'h4037f2c2, 32'h41dbacf6, 32'hc20db6b3, 32'h4282b062};
test_output[569] = '{32'h42c3ff4d};
test_index[569] = '{2};
test_input[4560:4567] = '{32'hc2c4b343, 32'hc2c13ea4, 32'hc23be6d8, 32'hc1c63420, 32'h42944bbe, 32'h42c2dc92, 32'h417e8467, 32'h3f89e340};
test_output[570] = '{32'h42c2dc92};
test_index[570] = '{5};
test_input[4568:4575] = '{32'hc282a9b5, 32'h42c59a36, 32'h42661fca, 32'h4112f882, 32'h42c54ef1, 32'h42c6be40, 32'hc2a0d1af, 32'h41cb15ae};
test_output[571] = '{32'h42c6be40};
test_index[571] = '{5};
test_input[4576:4583] = '{32'h429cc464, 32'hc2a8cfbf, 32'hc1810add, 32'hc0e97384, 32'h425b53b2, 32'h42b792c3, 32'h41cc8207, 32'h42b13250};
test_output[572] = '{32'h42b792c3};
test_index[572] = '{5};
test_input[4584:4591] = '{32'hc251e350, 32'hc24e939d, 32'h42a47765, 32'h4223e018, 32'hc22ffd84, 32'h429fa59f, 32'hc03ff82a, 32'h42a3b8ae};
test_output[573] = '{32'h42a47765};
test_index[573] = '{2};
test_input[4592:4599] = '{32'h42a61287, 32'hc19b9301, 32'hc246bb09, 32'hc25d3b30, 32'hc1874222, 32'hc283400a, 32'h415bed1a, 32'hc1cdded9};
test_output[574] = '{32'h42a61287};
test_index[574] = '{0};
test_input[4600:4607] = '{32'hc2965791, 32'hc2c639eb, 32'hc018a81b, 32'h428b75d5, 32'h4282966f, 32'hbfaae30f, 32'hc2b4524d, 32'h4129cea4};
test_output[575] = '{32'h428b75d5};
test_index[575] = '{3};
test_input[4608:4615] = '{32'h41feb6b0, 32'hc26ad9c6, 32'hc18de789, 32'hc1c74842, 32'hc1a0e5c2, 32'h426ed5b5, 32'hc283cb9f, 32'hc0ba98a3};
test_output[576] = '{32'h426ed5b5};
test_index[576] = '{5};
test_input[4616:4623] = '{32'hc2715d87, 32'h42ab8235, 32'hc1361037, 32'h42361a5a, 32'hc202b8ce, 32'h428396f7, 32'h42911194, 32'hc254907b};
test_output[577] = '{32'h42ab8235};
test_index[577] = '{1};
test_input[4624:4631] = '{32'hc25da8f6, 32'hc11cf77b, 32'h41a75bf2, 32'hc2474db4, 32'hc27c7d19, 32'h413e3f24, 32'h415a9c5d, 32'hc2aa21d2};
test_output[578] = '{32'h41a75bf2};
test_index[578] = '{2};
test_input[4632:4639] = '{32'hc298d661, 32'hbf9500e1, 32'hc2b8d454, 32'hc2ba79a3, 32'hc250d18f, 32'h41cb8c1f, 32'hc27379ec, 32'hc2be383e};
test_output[579] = '{32'h41cb8c1f};
test_index[579] = '{5};
test_input[4640:4647] = '{32'h412c211b, 32'hc2949268, 32'h42a1a513, 32'hc28dbebe, 32'h42753f9e, 32'h4286b766, 32'h40f40bda, 32'h424cccb1};
test_output[580] = '{32'h42a1a513};
test_index[580] = '{2};
test_input[4648:4655] = '{32'h425a2b3a, 32'h423cfd58, 32'hc1a51628, 32'h42c4cfb2, 32'hc2c52a92, 32'hc28245e8, 32'hc18d8d08, 32'h418ae291};
test_output[581] = '{32'h42c4cfb2};
test_index[581] = '{3};
test_input[4656:4663] = '{32'h417d06da, 32'hc23a65b0, 32'hc1c84f50, 32'hc20319be, 32'h42784b50, 32'h426a6e42, 32'hc2b34652, 32'hc28c6ad9};
test_output[582] = '{32'h42784b50};
test_index[582] = '{4};
test_input[4664:4671] = '{32'h422c1ce2, 32'h42664ad1, 32'hc10ef538, 32'hc2a748b2, 32'h4237f104, 32'hc2124fd0, 32'hc2bd301f, 32'hc27dd249};
test_output[583] = '{32'h42664ad1};
test_index[583] = '{1};
test_input[4672:4679] = '{32'h42b563d7, 32'h42819590, 32'h42876365, 32'hc21dfff5, 32'hc258c9c2, 32'hc14ba26d, 32'h42ac05a1, 32'h41e0b7e8};
test_output[584] = '{32'h42b563d7};
test_index[584] = '{0};
test_input[4680:4687] = '{32'hc279cdfe, 32'h421b21d6, 32'h42b68ab6, 32'h407f49fa, 32'hc2305fea, 32'h41bc3f75, 32'h42a28861, 32'h4267a119};
test_output[585] = '{32'h42b68ab6};
test_index[585] = '{2};
test_input[4688:4695] = '{32'hc2ac2258, 32'h4175866c, 32'hc29c6e7f, 32'hc1c6fee0, 32'hc2bd17ee, 32'h412e2a7b, 32'h428188b7, 32'hc22781e4};
test_output[586] = '{32'h428188b7};
test_index[586] = '{6};
test_input[4696:4703] = '{32'h4288a9d6, 32'h41875a5b, 32'h425bcc96, 32'h42c65be2, 32'h41b32b74, 32'h41a55cd1, 32'hc20b3191, 32'h428fedae};
test_output[587] = '{32'h42c65be2};
test_index[587] = '{3};
test_input[4704:4711] = '{32'h4292143d, 32'h40e9d48a, 32'hc29dc926, 32'hc13dca0d, 32'hc282d787, 32'h419a51c5, 32'h429d9ae7, 32'h41544d75};
test_output[588] = '{32'h429d9ae7};
test_index[588] = '{6};
test_input[4712:4719] = '{32'h41c24943, 32'hc29f4493, 32'h41240801, 32'hc1a0348f, 32'h42851a09, 32'h42aa80fc, 32'hc19df920, 32'hc19df358};
test_output[589] = '{32'h42aa80fc};
test_index[589] = '{5};
test_input[4720:4727] = '{32'hbffec3d1, 32'hc07a0632, 32'h4211b5dd, 32'h427d0210, 32'h42b79af4, 32'hc1e08f30, 32'hc1f35a7d, 32'h41405d64};
test_output[590] = '{32'h42b79af4};
test_index[590] = '{4};
test_input[4728:4735] = '{32'hc2bef38e, 32'hc21a797d, 32'hc2971ab1, 32'hc21e76bb, 32'hc103cfc2, 32'h4260a547, 32'hc22bc390, 32'hc24c41d0};
test_output[591] = '{32'h4260a547};
test_index[591] = '{5};
test_input[4736:4743] = '{32'hc296ae22, 32'hc211048b, 32'h42bff51b, 32'hc21eaf17, 32'hc21fa2ab, 32'hc281bf06, 32'h425e1bce, 32'h414c3b2a};
test_output[592] = '{32'h42bff51b};
test_index[592] = '{2};
test_input[4744:4751] = '{32'hc22d71ec, 32'h4211b645, 32'h422a2e94, 32'h4193fffa, 32'h420923ac, 32'h41391734, 32'h428352c1, 32'h4168f237};
test_output[593] = '{32'h428352c1};
test_index[593] = '{6};
test_input[4752:4759] = '{32'hc1684d8e, 32'h41329661, 32'h427255f6, 32'hc25fee69, 32'h428f96b9, 32'hc21bbfbb, 32'h4182a641, 32'h428146c9};
test_output[594] = '{32'h428f96b9};
test_index[594] = '{4};
test_input[4760:4767] = '{32'hc2843b7f, 32'hc2509019, 32'hc18b0d71, 32'h429e18a0, 32'h428f029e, 32'hc286e257, 32'hc286ede7, 32'h41dd9f44};
test_output[595] = '{32'h429e18a0};
test_index[595] = '{3};
test_input[4768:4775] = '{32'h42c22a16, 32'hc222bf9b, 32'hc27d7d41, 32'hc15bc793, 32'h41c470a1, 32'h421cd75e, 32'h42aa7410, 32'h420c77b3};
test_output[596] = '{32'h42c22a16};
test_index[596] = '{0};
test_input[4776:4783] = '{32'hc2c72d75, 32'h421191e0, 32'hc2c5448b, 32'h40f38fa7, 32'h42c27db2, 32'h40875b70, 32'h4212b07f, 32'hc21df1e8};
test_output[597] = '{32'h42c27db2};
test_index[597] = '{4};
test_input[4784:4791] = '{32'h42627fb4, 32'hc292c2af, 32'hc2c3ab38, 32'h42abd920, 32'hc13fc2ef, 32'hc065f753, 32'hc2c36823, 32'hc1a0ff77};
test_output[598] = '{32'h42abd920};
test_index[598] = '{3};
test_input[4792:4799] = '{32'hc270cb38, 32'hc2bd9328, 32'h42568fd4, 32'h41f1cc4a, 32'h41bffbaa, 32'hc29149be, 32'hc126000f, 32'h42a5b380};
test_output[599] = '{32'h42a5b380};
test_index[599] = '{7};
test_input[4800:4807] = '{32'hc239ac6b, 32'h42707a23, 32'h421c26f1, 32'hc2af3900, 32'h417247a9, 32'hc29b6b52, 32'h42988501, 32'h4162574d};
test_output[600] = '{32'h42988501};
test_index[600] = '{6};
test_input[4808:4815] = '{32'h42849c7d, 32'h40cc4d29, 32'h414dd125, 32'hc149eee2, 32'hc2a5cda2, 32'h42a72503, 32'h42365ccd, 32'h40b30550};
test_output[601] = '{32'h42a72503};
test_index[601] = '{5};
test_input[4816:4823] = '{32'h42c09116, 32'h425732e8, 32'hc29d5adf, 32'h40836300, 32'hc25e5fb2, 32'h414d6bc3, 32'hc1e410c2, 32'h41ec8640};
test_output[602] = '{32'h42c09116};
test_index[602] = '{0};
test_input[4824:4831] = '{32'hc1501b82, 32'h40d05eda, 32'hc1dd90da, 32'hc139c5f4, 32'h42c3cc1c, 32'hc256972d, 32'h42561fda, 32'hc22454ea};
test_output[603] = '{32'h42c3cc1c};
test_index[603] = '{4};
test_input[4832:4839] = '{32'h42804853, 32'hc231e4bc, 32'hc2b0d7b2, 32'h42bde4f3, 32'h421e3b99, 32'hc2841826, 32'hc25b6aac, 32'h42b624b2};
test_output[604] = '{32'h42bde4f3};
test_index[604] = '{3};
test_input[4840:4847] = '{32'h412f7cce, 32'h42307965, 32'h411f6a15, 32'h42ad12e8, 32'h425105e7, 32'h42b71014, 32'h4190ef63, 32'hc2b0be92};
test_output[605] = '{32'h42b71014};
test_index[605] = '{5};
test_input[4848:4855] = '{32'h42aca4bd, 32'h42b3d719, 32'h414688c0, 32'hc1cd7f59, 32'h4242f75d, 32'hc0f5a592, 32'hc218508c, 32'h42bec2cb};
test_output[606] = '{32'h42bec2cb};
test_index[606] = '{7};
test_input[4856:4863] = '{32'h42906866, 32'h429b4b92, 32'hc12e3482, 32'h42aa4274, 32'h41a64eac, 32'hc2aff40d, 32'h418e08ff, 32'h42912224};
test_output[607] = '{32'h42aa4274};
test_index[607] = '{3};
test_input[4864:4871] = '{32'h428b51bf, 32'h420565a1, 32'hc21aed0f, 32'hc1b168b0, 32'h42c3d182, 32'h429222dc, 32'hc24197da, 32'hc1180272};
test_output[608] = '{32'h42c3d182};
test_index[608] = '{4};
test_input[4872:4879] = '{32'hc1f4c8aa, 32'h423348e1, 32'hc28f63f3, 32'hc21ea0df, 32'h429f8e87, 32'hc2b748af, 32'hc15c5b23, 32'h410805f9};
test_output[609] = '{32'h429f8e87};
test_index[609] = '{4};
test_input[4880:4887] = '{32'h426b14b1, 32'h421a3331, 32'hc1c2bd25, 32'hc03d7e44, 32'h428551a7, 32'h41d1876a, 32'h428f72f8, 32'hc24e4eb9};
test_output[610] = '{32'h428f72f8};
test_index[610] = '{6};
test_input[4888:4895] = '{32'hc293c15a, 32'h42409de5, 32'hc21a72c5, 32'h420281bf, 32'h42947bd5, 32'hc10044f6, 32'h414ebdf1, 32'h426abaef};
test_output[611] = '{32'h42947bd5};
test_index[611] = '{4};
test_input[4896:4903] = '{32'hc26e2611, 32'hc2c2dfff, 32'hc2550191, 32'h42b87066, 32'h42c5edcc, 32'h42c7a368, 32'h42b60895, 32'hc2b9d98a};
test_output[612] = '{32'h42c7a368};
test_index[612] = '{5};
test_input[4904:4911] = '{32'h428ff7b1, 32'h4198d67c, 32'hc16e2b33, 32'hc26e422e, 32'hbf833e7c, 32'hc281386f, 32'hc228a152, 32'hc2053628};
test_output[613] = '{32'h428ff7b1};
test_index[613] = '{0};
test_input[4912:4919] = '{32'h4298e8b1, 32'hc2b7e6f2, 32'h42046fa5, 32'h4213388f, 32'hc1b1e559, 32'hc23bd0c1, 32'hc2295687, 32'h429f521f};
test_output[614] = '{32'h429f521f};
test_index[614] = '{7};
test_input[4920:4927] = '{32'h41702f8e, 32'h42b74a10, 32'hc1eb20b0, 32'hc2b20b69, 32'h3fb22566, 32'hc274612c, 32'h421b380f, 32'h4220439e};
test_output[615] = '{32'h42b74a10};
test_index[615] = '{1};
test_input[4928:4935] = '{32'hc2afc18e, 32'hc1f349c0, 32'h42110a64, 32'h4250378a, 32'hc2c4e29b, 32'h423314ec, 32'h42432f3b, 32'hc2bec51f};
test_output[616] = '{32'h4250378a};
test_index[616] = '{3};
test_input[4936:4943] = '{32'hc1367fcf, 32'h42262977, 32'h42b34b60, 32'h4166844f, 32'hc26359f6, 32'h41d08ca5, 32'h41bd0b83, 32'hc28ca7de};
test_output[617] = '{32'h42b34b60};
test_index[617] = '{2};
test_input[4944:4951] = '{32'h42905b1a, 32'h42bf4e92, 32'h427e0cdb, 32'h41b3507a, 32'h42a1920a, 32'hc2287f9e, 32'h42b03093, 32'hc2851d11};
test_output[618] = '{32'h42bf4e92};
test_index[618] = '{1};
test_input[4952:4959] = '{32'hc23f6c69, 32'h41db12c4, 32'hc2345515, 32'h4223bf9e, 32'hc1c332f9, 32'hc067c194, 32'h419a0039, 32'hc1ec4b57};
test_output[619] = '{32'h4223bf9e};
test_index[619] = '{3};
test_input[4960:4967] = '{32'h42405c6e, 32'hc2631ac1, 32'h4143f339, 32'h4246c9ed, 32'h429790df, 32'h40e8b509, 32'h42822e8b, 32'hc2b6329d};
test_output[620] = '{32'h429790df};
test_index[620] = '{4};
test_input[4968:4975] = '{32'hc1b1ec77, 32'hc290b203, 32'h41e6d1b1, 32'hc2b37ec1, 32'h42840c37, 32'h4244e260, 32'h425bdf27, 32'h42986097};
test_output[621] = '{32'h42986097};
test_index[621] = '{7};
test_input[4976:4983] = '{32'h42c6e394, 32'h426dcba6, 32'h42b823ba, 32'hc19332f0, 32'hc29adc1d, 32'h42b424eb, 32'hc2b0b3ca, 32'h421052a1};
test_output[622] = '{32'h42c6e394};
test_index[622] = '{0};
test_input[4984:4991] = '{32'h42531df8, 32'hc201afd5, 32'h412a4217, 32'h41860ca4, 32'h40804ca1, 32'hc2022a6a, 32'h42985fa9, 32'hc2c20596};
test_output[623] = '{32'h42985fa9};
test_index[623] = '{6};
test_input[4992:4999] = '{32'h42af375e, 32'h420c6fe5, 32'h42a131e1, 32'h40de7187, 32'hc112bc64, 32'h4226a1e9, 32'hc15e38cc, 32'hc2a88051};
test_output[624] = '{32'h42af375e};
test_index[624] = '{0};
test_input[5000:5007] = '{32'hc191cfba, 32'hc2329612, 32'hc1d784f8, 32'h42b00221, 32'hc2551ff4, 32'h42aaa370, 32'h417c6604, 32'hc10c8b09};
test_output[625] = '{32'h42b00221};
test_index[625] = '{3};
test_input[5008:5015] = '{32'h42ac1842, 32'hc1ac8d61, 32'h41eaa212, 32'hc2bb4623, 32'hc22e196f, 32'hc2308900, 32'h3fa6447a, 32'h41a79075};
test_output[626] = '{32'h42ac1842};
test_index[626] = '{0};
test_input[5016:5023] = '{32'hc29c9207, 32'hc29d8b99, 32'h42bf9c4d, 32'hc2c6a696, 32'h41da207f, 32'h42a1da1a, 32'h4270e3f4, 32'hc07a7d55};
test_output[627] = '{32'h42bf9c4d};
test_index[627] = '{2};
test_input[5024:5031] = '{32'h42933d88, 32'h424fa4fe, 32'hc25455b7, 32'hc1d09b20, 32'hc27feae7, 32'hc11d840d, 32'h42890547, 32'h42a987f2};
test_output[628] = '{32'h42a987f2};
test_index[628] = '{7};
test_input[5032:5039] = '{32'hc232211a, 32'h42b1a6c2, 32'hc1e39da4, 32'h42a77f79, 32'h42c62b05, 32'hc16502eb, 32'hc277cee2, 32'hc0ff5698};
test_output[629] = '{32'h42c62b05};
test_index[629] = '{4};
test_input[5040:5047] = '{32'hc2b349e4, 32'h428ce26d, 32'h42abcf17, 32'hc2840d2d, 32'h42acd10d, 32'hc250a11f, 32'hc288f0c1, 32'h4175f785};
test_output[630] = '{32'h42acd10d};
test_index[630] = '{4};
test_input[5048:5055] = '{32'hc2b9c619, 32'h42772dbc, 32'hc29653e2, 32'h421cfd4f, 32'hc2badee1, 32'h417892c6, 32'hc1fda976, 32'h424c21d9};
test_output[631] = '{32'h42772dbc};
test_index[631] = '{1};
test_input[5056:5063] = '{32'h4232571c, 32'hc2844f52, 32'hc231a3aa, 32'h42184a16, 32'hc1e78c73, 32'h3ff39da3, 32'hc2b8c27a, 32'h425a2925};
test_output[632] = '{32'h425a2925};
test_index[632] = '{7};
test_input[5064:5071] = '{32'hc297a6c1, 32'hc2844cac, 32'h419eeda5, 32'h42b52be0, 32'hc13ea9ac, 32'h4216623f, 32'h4162dc98, 32'hc29e5c2a};
test_output[633] = '{32'h42b52be0};
test_index[633] = '{3};
test_input[5072:5079] = '{32'h42126416, 32'h419cc8ee, 32'h41025a2c, 32'hc2c5feb2, 32'hc06a5fdc, 32'hc2acf809, 32'h4100d3a2, 32'hc238adda};
test_output[634] = '{32'h42126416};
test_index[634] = '{0};
test_input[5080:5087] = '{32'hc2187a65, 32'hc21a2b20, 32'hc0c03cda, 32'h425c1dba, 32'hc2312ced, 32'h4224a4da, 32'h42458dd8, 32'hc2999537};
test_output[635] = '{32'h425c1dba};
test_index[635] = '{3};
test_input[5088:5095] = '{32'hc1ac9bed, 32'hc23ae240, 32'hc261a9ef, 32'h4209e504, 32'hc0d8eb59, 32'hc2b66998, 32'h4239ff94, 32'hc2680407};
test_output[636] = '{32'h4239ff94};
test_index[636] = '{6};
test_input[5096:5103] = '{32'h4162c5ef, 32'hc292e735, 32'hc21e9a87, 32'hc2b25dd9, 32'hc185eaf5, 32'hc10e36c0, 32'h4241af5c, 32'hc2b3d4aa};
test_output[637] = '{32'h4241af5c};
test_index[637] = '{6};
test_input[5104:5111] = '{32'h42adc105, 32'h42c46124, 32'hc0e29b06, 32'hc28edd49, 32'hc29f76c9, 32'hc235eca3, 32'h425abf2b, 32'hc2c2dea6};
test_output[638] = '{32'h42c46124};
test_index[638] = '{1};
test_input[5112:5119] = '{32'h4077e639, 32'hc2a141de, 32'h41b5f108, 32'h4250ed77, 32'hc24bf41c, 32'h429e079c, 32'h426d2883, 32'h41de93e3};
test_output[639] = '{32'h429e079c};
test_index[639] = '{5};
test_input[5120:5127] = '{32'hc199262e, 32'hc180ae46, 32'hc178e76c, 32'h42712be6, 32'h428f6ccf, 32'hc29fe526, 32'h41d265db, 32'h42b4bdae};
test_output[640] = '{32'h42b4bdae};
test_index[640] = '{7};
test_input[5128:5135] = '{32'hc1f7ca27, 32'h415402e1, 32'h42acf686, 32'hc2c62a8e, 32'hc19c6d12, 32'h42bfcc52, 32'h41328ac0, 32'h4258fe91};
test_output[641] = '{32'h42bfcc52};
test_index[641] = '{5};
test_input[5136:5143] = '{32'h42ae10a4, 32'hc221bddc, 32'h42b13ebd, 32'hc286ec09, 32'hc1599f67, 32'h42af238f, 32'hc200ec41, 32'hc2b8495d};
test_output[642] = '{32'h42b13ebd};
test_index[642] = '{2};
test_input[5144:5151] = '{32'hc2134434, 32'h42b35d30, 32'hc2b8c926, 32'h4132eecf, 32'h41f50e82, 32'h42635cc1, 32'h428fe024, 32'h41d0709f};
test_output[643] = '{32'h42b35d30};
test_index[643] = '{1};
test_input[5152:5159] = '{32'hc13a60e3, 32'h4283779f, 32'h41a13849, 32'hc2c27109, 32'h4212c9c3, 32'hc2569a86, 32'h42bf0dec, 32'h42c28f83};
test_output[644] = '{32'h42c28f83};
test_index[644] = '{7};
test_input[5160:5167] = '{32'h419e0aee, 32'hc1545f3f, 32'h428e58e9, 32'h429a1cd8, 32'h410a0cca, 32'hc0902213, 32'h40a8f04d, 32'h42b4ed9c};
test_output[645] = '{32'h42b4ed9c};
test_index[645] = '{7};
test_input[5168:5175] = '{32'h41eda211, 32'hc279193b, 32'hc28cd31d, 32'hc2b98c0c, 32'hc238e4a6, 32'h42a9df24, 32'hc1bed986, 32'h41c146e2};
test_output[646] = '{32'h42a9df24};
test_index[646] = '{5};
test_input[5176:5183] = '{32'h3f37df7f, 32'h424b0494, 32'hc21cb0c5, 32'hc19c78f8, 32'h42b8484f, 32'hc0cff3a5, 32'hc28facef, 32'hc2bd0e59};
test_output[647] = '{32'h42b8484f};
test_index[647] = '{4};
test_input[5184:5191] = '{32'h4283416b, 32'h42290ba2, 32'h42c7e047, 32'h421a817d, 32'hc269d711, 32'h42b6c4a2, 32'hc02289b3, 32'hc15a2e69};
test_output[648] = '{32'h42c7e047};
test_index[648] = '{2};
test_input[5192:5199] = '{32'h4295697e, 32'hc0a8251d, 32'h42080a69, 32'hc2567381, 32'h427d0203, 32'hc17f079e, 32'h4254c5fc, 32'hc2a4f044};
test_output[649] = '{32'h4295697e};
test_index[649] = '{0};
test_input[5200:5207] = '{32'h425e1d90, 32'h429fc44b, 32'hc2022666, 32'h40328a43, 32'h41b9fb61, 32'hc2b871bd, 32'h422f08fd, 32'hc2481841};
test_output[650] = '{32'h429fc44b};
test_index[650] = '{1};
test_input[5208:5215] = '{32'h42a7478c, 32'hc29498ed, 32'hc2c3d0f8, 32'h42b18adb, 32'h41eeb48e, 32'hc2c104c4, 32'h42995263, 32'h41d221fe};
test_output[651] = '{32'h42b18adb};
test_index[651] = '{3};
test_input[5216:5223] = '{32'hc232555c, 32'hc1e42d17, 32'hc21ba6c0, 32'hc28e01fd, 32'hc1152144, 32'h425313db, 32'h41b668d3, 32'h421579c1};
test_output[652] = '{32'h425313db};
test_index[652] = '{5};
test_input[5224:5231] = '{32'hc27d15ca, 32'hc2993b14, 32'hc284d23f, 32'h41d75ae4, 32'hc1ab1338, 32'hc2b6eed6, 32'hc1ff4ae3, 32'h4285db6b};
test_output[653] = '{32'h4285db6b};
test_index[653] = '{7};
test_input[5232:5239] = '{32'h428647a2, 32'hc2013cde, 32'hc2a6ac88, 32'hc2b1f41f, 32'h4031babe, 32'h42135e81, 32'h411dcf05, 32'h4118be36};
test_output[654] = '{32'h428647a2};
test_index[654] = '{0};
test_input[5240:5247] = '{32'hc2036b85, 32'h42723ae7, 32'h421535de, 32'h423c6582, 32'hc18c5d67, 32'hc26b4aef, 32'h42b6e453, 32'hc20be0af};
test_output[655] = '{32'h42b6e453};
test_index[655] = '{6};
test_input[5248:5255] = '{32'h41d49cdd, 32'hc29aed3f, 32'hc26ef577, 32'h41b091fd, 32'h428e02a6, 32'hc1624dcd, 32'hc2517d45, 32'hc222f94a};
test_output[656] = '{32'h428e02a6};
test_index[656] = '{4};
test_input[5256:5263] = '{32'h42944b63, 32'hc1d848ef, 32'h41cb6e69, 32'hc1e5ba85, 32'hc2c274b1, 32'h42b761f4, 32'hc27985a7, 32'hc2970376};
test_output[657] = '{32'h42b761f4};
test_index[657] = '{5};
test_input[5264:5271] = '{32'hc28eb352, 32'h41ccb687, 32'h4241e87e, 32'hc1b4c044, 32'hc2b177f2, 32'hc1ad5079, 32'hc21a0b60, 32'hc105b7af};
test_output[658] = '{32'h4241e87e};
test_index[658] = '{2};
test_input[5272:5279] = '{32'h42b751a2, 32'hc16b896d, 32'hc256d087, 32'hc20d9c17, 32'hc2521d20, 32'hc1d230c9, 32'hc2622df7, 32'h42c38d56};
test_output[659] = '{32'h42c38d56};
test_index[659] = '{7};
test_input[5280:5287] = '{32'hc2a622a4, 32'hc0f254cc, 32'h42aa61bd, 32'hc2be3722, 32'h41f0e3ce, 32'hc282b3f2, 32'h418f0e13, 32'hc1435820};
test_output[660] = '{32'h42aa61bd};
test_index[660] = '{2};
test_input[5288:5295] = '{32'h422ab997, 32'hc07578bc, 32'h42b5b707, 32'hc2547f50, 32'h4299c8a9, 32'hc2b40ae4, 32'hc28e2a0d, 32'hc17c2ba6};
test_output[661] = '{32'h42b5b707};
test_index[661] = '{2};
test_input[5296:5303] = '{32'hc186e331, 32'hc249b9d0, 32'h42881851, 32'h42845799, 32'hc146cee1, 32'hc1d3e0c9, 32'hc2246fc8, 32'h41eef3c3};
test_output[662] = '{32'h42881851};
test_index[662] = '{2};
test_input[5304:5311] = '{32'h4286185d, 32'h42838449, 32'h421ea9f0, 32'h41b7349b, 32'h4251bd0d, 32'hc15619bd, 32'hc1e7619b, 32'h420e774c};
test_output[663] = '{32'h4286185d};
test_index[663] = '{0};
test_input[5312:5319] = '{32'h42bfeb98, 32'h4213e3db, 32'h42918333, 32'h4235ffd0, 32'h42104552, 32'hc2b90ab7, 32'h4164fd35, 32'hc03b3f3a};
test_output[664] = '{32'h42bfeb98};
test_index[664] = '{0};
test_input[5320:5327] = '{32'h41ef8e13, 32'h42c19e85, 32'hc267b5ca, 32'hc2aa443e, 32'h4246dd97, 32'hc2c62f30, 32'h421f0af8, 32'hc26af838};
test_output[665] = '{32'h42c19e85};
test_index[665] = '{1};
test_input[5328:5335] = '{32'h407fc33e, 32'h42c701af, 32'h412582b0, 32'h424e350a, 32'hc1db29e6, 32'h41a8c47c, 32'h41b4cb2b, 32'h421c0de6};
test_output[666] = '{32'h42c701af};
test_index[666] = '{1};
test_input[5336:5343] = '{32'hc26f00a1, 32'hc2129319, 32'h424c2e9b, 32'h4298e930, 32'h4255c8cd, 32'hc282a1e6, 32'h427fefcb, 32'h42c6e5cf};
test_output[667] = '{32'h42c6e5cf};
test_index[667] = '{7};
test_input[5344:5351] = '{32'hc28a5ca0, 32'hc285cbcb, 32'hc284faaa, 32'h413c7dbf, 32'h4290f500, 32'hc1cf28fc, 32'hc26d83e6, 32'hc2601f9d};
test_output[668] = '{32'h4290f500};
test_index[668] = '{4};
test_input[5352:5359] = '{32'hc2513f25, 32'h42285d4f, 32'hc01da764, 32'hc0c3c495, 32'h42b08ef5, 32'hc267264f, 32'hc2845514, 32'h42501c94};
test_output[669] = '{32'h42b08ef5};
test_index[669] = '{4};
test_input[5360:5367] = '{32'hc1ceecbf, 32'h4278c265, 32'h428011a9, 32'hc200ec5e, 32'h4173ab62, 32'h42045a1b, 32'hc019b0db, 32'hc23a8e71};
test_output[670] = '{32'h428011a9};
test_index[670] = '{2};
test_input[5368:5375] = '{32'h42458e14, 32'h40ff33a4, 32'hc2b46cae, 32'h42076de5, 32'h4250aa67, 32'h429d13bc, 32'hc2a65601, 32'h414bb05e};
test_output[671] = '{32'h429d13bc};
test_index[671] = '{5};
test_input[5376:5383] = '{32'hc2c07595, 32'h42b8c981, 32'hc204ac2e, 32'hc2a29635, 32'hc2300ac1, 32'h423fd7d8, 32'hc2658ca6, 32'h42aede43};
test_output[672] = '{32'h42b8c981};
test_index[672] = '{1};
test_input[5384:5391] = '{32'h411de5a5, 32'h42ac38cc, 32'h424fee0f, 32'hc29e4dea, 32'hc2b1073d, 32'h4287e80e, 32'hc214e7f1, 32'h421be11a};
test_output[673] = '{32'h42ac38cc};
test_index[673] = '{1};
test_input[5392:5399] = '{32'h4227a31e, 32'h4295de63, 32'h419464d7, 32'hc22566e2, 32'hc2ad20f4, 32'h41c4d5e5, 32'h408bbac0, 32'hc2078de0};
test_output[674] = '{32'h4295de63};
test_index[674] = '{1};
test_input[5400:5407] = '{32'h428cb14b, 32'h42a8c538, 32'hc291f608, 32'hc2be0d27, 32'h4203d4e7, 32'h42b56af6, 32'hc27e9d91, 32'h42a57d2d};
test_output[675] = '{32'h42b56af6};
test_index[675] = '{5};
test_input[5408:5415] = '{32'h42108cb6, 32'hc2ba050d, 32'h42bf788e, 32'h42b63369, 32'h42105fb3, 32'hc059a5ad, 32'h42a6966c, 32'hc2386d0f};
test_output[676] = '{32'h42bf788e};
test_index[676] = '{2};
test_input[5416:5423] = '{32'hc2867cc6, 32'hc296ccca, 32'h42aeeb72, 32'hc1f87b1f, 32'h40f919f5, 32'h41d4137c, 32'hc1e2ba75, 32'h41659834};
test_output[677] = '{32'h42aeeb72};
test_index[677] = '{2};
test_input[5424:5431] = '{32'h419830c9, 32'hc0ed6fef, 32'h4281e120, 32'h423a8338, 32'hc267dc2f, 32'h42bbe2f3, 32'h42398d5b, 32'h425c8621};
test_output[678] = '{32'h42bbe2f3};
test_index[678] = '{5};
test_input[5432:5439] = '{32'h42a409e7, 32'hc26b52ca, 32'hc2b81775, 32'h4224cf07, 32'h42a42344, 32'hc2601762, 32'hc262cacc, 32'hc2b41552};
test_output[679] = '{32'h42a42344};
test_index[679] = '{4};
test_input[5440:5447] = '{32'hc1897db8, 32'hc292c82d, 32'h41d9abbf, 32'hc0a19f31, 32'h41a0c931, 32'h3fb29157, 32'hc2346e33, 32'hc2753c0c};
test_output[680] = '{32'h41d9abbf};
test_index[680] = '{2};
test_input[5448:5455] = '{32'h42664eba, 32'h42997674, 32'h41f03f2f, 32'hc20897ae, 32'hc2433acd, 32'hc12a2ca1, 32'hc1ec58c9, 32'h41dafd4b};
test_output[681] = '{32'h42997674};
test_index[681] = '{1};
test_input[5456:5463] = '{32'h406c33b3, 32'h424f965b, 32'hc2c1d6f7, 32'hc28cca11, 32'h427e8157, 32'hc226d72f, 32'h424bc40d, 32'h422baca1};
test_output[682] = '{32'h427e8157};
test_index[682] = '{4};
test_input[5464:5471] = '{32'hc1e5cdc4, 32'hc24d2f5b, 32'hc1961b7b, 32'h408c7dc5, 32'hc28f786b, 32'h42b96ee7, 32'hc28fd0a3, 32'hc1a2ee77};
test_output[683] = '{32'h42b96ee7};
test_index[683] = '{5};
test_input[5472:5479] = '{32'hc258deaa, 32'h42275c49, 32'h41c5de82, 32'h42bd494b, 32'hc2adb85f, 32'h4223c501, 32'hc178d7c5, 32'h4235afd9};
test_output[684] = '{32'h42bd494b};
test_index[684] = '{3};
test_input[5480:5487] = '{32'h428e502e, 32'hc20df0ef, 32'h4239b8c9, 32'hc28d9cfe, 32'hc28118d3, 32'hc29f10e8, 32'h42b609fe, 32'h41806f6b};
test_output[685] = '{32'h42b609fe};
test_index[685] = '{6};
test_input[5488:5495] = '{32'hc2760974, 32'h42677575, 32'h42b018de, 32'h42928048, 32'hc2622495, 32'h419ae535, 32'hc28ace57, 32'h419a3026};
test_output[686] = '{32'h42b018de};
test_index[686] = '{2};
test_input[5496:5503] = '{32'h429df44d, 32'h4291b955, 32'hc29d0bfa, 32'h42883975, 32'hc2a84043, 32'hc210c858, 32'hc16ca6bb, 32'h4104dc36};
test_output[687] = '{32'h429df44d};
test_index[687] = '{0};
test_input[5504:5511] = '{32'hc2c550dd, 32'hc06a1c8c, 32'hc273f973, 32'h42911d8d, 32'h415898e0, 32'h42a7a588, 32'h42c4e880, 32'hc2b4920b};
test_output[688] = '{32'h42c4e880};
test_index[688] = '{6};
test_input[5512:5519] = '{32'h42afc41c, 32'hc260524f, 32'hc2a6c081, 32'hc1a597d0, 32'h42781a2a, 32'h4279766b, 32'h42a6b055, 32'h42a98a05};
test_output[689] = '{32'h42afc41c};
test_index[689] = '{0};
test_input[5520:5527] = '{32'hc264a13e, 32'hc1862845, 32'hc1e6e039, 32'hc24f884a, 32'hc1d13f86, 32'hc26ea9db, 32'h4227e1f3, 32'h42c205bb};
test_output[690] = '{32'h42c205bb};
test_index[690] = '{7};
test_input[5528:5535] = '{32'h41eb5101, 32'hc25ed367, 32'h42bdf638, 32'hc24e6b72, 32'h4279c40b, 32'hc2aa6bdf, 32'h42bd99a7, 32'h42a6c868};
test_output[691] = '{32'h42bdf638};
test_index[691] = '{2};
test_input[5536:5543] = '{32'hc2a5fd63, 32'h42b59e6c, 32'hc2b72549, 32'hc2399c0e, 32'h42bc32c9, 32'hc20536cd, 32'h40fd8f27, 32'h413285c7};
test_output[692] = '{32'h42bc32c9};
test_index[692] = '{4};
test_input[5544:5551] = '{32'hc256b1db, 32'hc1b0e402, 32'h4256b0d9, 32'h42324b92, 32'hc2419236, 32'hc29b2c47, 32'hc23f988c, 32'h42ab228e};
test_output[693] = '{32'h42ab228e};
test_index[693] = '{7};
test_input[5552:5559] = '{32'h428b3a1b, 32'hc2883e72, 32'hc250556a, 32'hc2191f87, 32'hc29f7b42, 32'h41f22b9a, 32'h4174b5d7, 32'h411b8fc7};
test_output[694] = '{32'h428b3a1b};
test_index[694] = '{0};
test_input[5560:5567] = '{32'h423e7889, 32'h40e33169, 32'hc2913c7d, 32'h418637e0, 32'hc2c63b3f, 32'hc231c8a2, 32'hc28e4988, 32'hc0e416f1};
test_output[695] = '{32'h423e7889};
test_index[695] = '{0};
test_input[5568:5575] = '{32'h420e7b68, 32'h42223898, 32'hc244e3f6, 32'h42614f36, 32'h42c413b5, 32'hc1d6ed62, 32'hc28b52a4, 32'hc2a6e3c8};
test_output[696] = '{32'h42c413b5};
test_index[696] = '{4};
test_input[5576:5583] = '{32'hc1bb8873, 32'hc26301ce, 32'h4252ff96, 32'h42bfee1a, 32'hc0924f2e, 32'h42930dd9, 32'h42ab8ea1, 32'hc2920cd7};
test_output[697] = '{32'h42bfee1a};
test_index[697] = '{3};
test_input[5584:5591] = '{32'h422c9f1f, 32'h42a2cab8, 32'h3f6663fa, 32'h40d468ae, 32'h41174099, 32'hc2c6e9db, 32'hc1eb9712, 32'hc0578965};
test_output[698] = '{32'h42a2cab8};
test_index[698] = '{1};
test_input[5592:5599] = '{32'hc26c71fa, 32'hc24bb46e, 32'h421e520f, 32'h42b93f3d, 32'hc21e683e, 32'hc2085d28, 32'hc0f3ff28, 32'h41d8e6af};
test_output[699] = '{32'h42b93f3d};
test_index[699] = '{3};
test_input[5600:5607] = '{32'h4274829e, 32'hc2aa5a1b, 32'h42921b73, 32'hc20a5b4d, 32'h4236fea2, 32'h41c7cae7, 32'h42b45c67, 32'hc29c1e3d};
test_output[700] = '{32'h42b45c67};
test_index[700] = '{6};
test_input[5608:5615] = '{32'h42503030, 32'hc2ab16f1, 32'h42405fb7, 32'hc1b72f95, 32'hbc8772e8, 32'h41831707, 32'hc293585a, 32'h42b050c6};
test_output[701] = '{32'h42b050c6};
test_index[701] = '{7};
test_input[5616:5623] = '{32'hc271be45, 32'hc22e559c, 32'h41cb622a, 32'h42abe510, 32'hc25ed250, 32'h42824ba1, 32'hc280341d, 32'hc2846c07};
test_output[702] = '{32'h42abe510};
test_index[702] = '{3};
test_input[5624:5631] = '{32'h4204a3fd, 32'hc2bce9b9, 32'hc24d9b6c, 32'hc29be795, 32'h425a7603, 32'h41ceedba, 32'h42aaa10e, 32'hc2999a3c};
test_output[703] = '{32'h42aaa10e};
test_index[703] = '{6};
test_input[5632:5639] = '{32'h4210ea43, 32'h42aa3dfb, 32'hc268f550, 32'hc295d10c, 32'h42440cda, 32'h41454d5b, 32'hc27b86d2, 32'h41e7840f};
test_output[704] = '{32'h42aa3dfb};
test_index[704] = '{1};
test_input[5640:5647] = '{32'h426104a2, 32'h425e3b05, 32'h40df170b, 32'h429b8d55, 32'hc2a936bf, 32'h41271618, 32'hc2257de2, 32'hc26864a4};
test_output[705] = '{32'h429b8d55};
test_index[705] = '{3};
test_input[5648:5655] = '{32'hc28f84e0, 32'hc10d027e, 32'h4296c2dd, 32'h42bda70e, 32'hc295df31, 32'h42609598, 32'hc1a594b2, 32'hc216116e};
test_output[706] = '{32'h42bda70e};
test_index[706] = '{3};
test_input[5656:5663] = '{32'h42a810c6, 32'hc28853aa, 32'hc26c28b4, 32'hc26e75c1, 32'hc11d9b4d, 32'h4263559c, 32'hbb90bd6a, 32'hc2500967};
test_output[707] = '{32'h42a810c6};
test_index[707] = '{0};
test_input[5664:5671] = '{32'hc19d12a0, 32'hc2aa826b, 32'h42794785, 32'hc1b67967, 32'hc287b577, 32'hc208f3e8, 32'h42618777, 32'h42364e39};
test_output[708] = '{32'h42794785};
test_index[708] = '{2};
test_input[5672:5679] = '{32'hc1ebf889, 32'hc2a49d22, 32'hc23be55b, 32'hc1969f63, 32'hc2927cbc, 32'hc1ae3b4a, 32'hc2a8d918, 32'h42bc8b9f};
test_output[709] = '{32'h42bc8b9f};
test_index[709] = '{7};
test_input[5680:5687] = '{32'h422aaa57, 32'h41a9988a, 32'h42880dfb, 32'hc28998e5, 32'h4194c5c2, 32'hc2af7ebc, 32'hc2b648e9, 32'h42688063};
test_output[710] = '{32'h42880dfb};
test_index[710] = '{2};
test_input[5688:5695] = '{32'h427fb2ef, 32'h4298810f, 32'h41879d80, 32'h42b4a36d, 32'hc210aa8f, 32'hc25db2ac, 32'hc2c30108, 32'hc0b0daff};
test_output[711] = '{32'h42b4a36d};
test_index[711] = '{3};
test_input[5696:5703] = '{32'hc222e595, 32'h3e21517b, 32'h42312d1e, 32'h4278efd2, 32'hc2bcf9c4, 32'hc1819fd0, 32'hc21e2fbb, 32'h421f4914};
test_output[712] = '{32'h4278efd2};
test_index[712] = '{3};
test_input[5704:5711] = '{32'hc2ab0773, 32'hc2c7166b, 32'hc1e257a1, 32'hc1a16490, 32'hc266593f, 32'hc1419cc0, 32'h41e878b4, 32'h4227a3ec};
test_output[713] = '{32'h4227a3ec};
test_index[713] = '{7};
test_input[5712:5719] = '{32'hc139a7c8, 32'hc25f6e35, 32'hc2c643b2, 32'h41b0b4ee, 32'hc2910f6d, 32'h41fcc9a1, 32'h41bfe189, 32'hc2a3fb92};
test_output[714] = '{32'h41fcc9a1};
test_index[714] = '{5};
test_input[5720:5727] = '{32'h41ae3360, 32'hc2b8975d, 32'hc1b952f0, 32'h4283b4d5, 32'hc1cf5d7f, 32'hc2a150b9, 32'hc24ecac5, 32'h418e864d};
test_output[715] = '{32'h4283b4d5};
test_index[715] = '{3};
test_input[5728:5735] = '{32'h426ccb57, 32'h41376e9e, 32'h42adc6a2, 32'h4154700e, 32'hc09fadcc, 32'h428ad3e6, 32'h42c2b61f, 32'hc2826aa4};
test_output[716] = '{32'h42c2b61f};
test_index[716] = '{6};
test_input[5736:5743] = '{32'hc2a7cfcd, 32'h42941471, 32'hc24aaff9, 32'hc22415a2, 32'h417e5679, 32'h4090f85b, 32'h401f7bec, 32'hc263460e};
test_output[717] = '{32'h42941471};
test_index[717] = '{1};
test_input[5744:5751] = '{32'h42a24bfd, 32'h41dadf56, 32'hc241e30e, 32'h42902adc, 32'h42be18b0, 32'hc1142211, 32'hc2b406a4, 32'hc299e0e7};
test_output[718] = '{32'h42be18b0};
test_index[718] = '{4};
test_input[5752:5759] = '{32'h41aedf26, 32'h42b9f560, 32'h42585f22, 32'h418e2f9a, 32'h429ccef4, 32'hc246d321, 32'h42000ac9, 32'hc1a6f710};
test_output[719] = '{32'h42b9f560};
test_index[719] = '{1};
test_input[5760:5767] = '{32'h40e29238, 32'hc2009fc2, 32'hc203be83, 32'h4256b823, 32'h42973d5b, 32'h427bdabf, 32'h429ba39d, 32'h42a9a8d8};
test_output[720] = '{32'h42a9a8d8};
test_index[720] = '{7};
test_input[5768:5775] = '{32'hc25295fd, 32'hc1dab848, 32'hc1cbd916, 32'hc1c49497, 32'h4280a29e, 32'hc18ac103, 32'h41ca5a4d, 32'h427114df};
test_output[721] = '{32'h4280a29e};
test_index[721] = '{4};
test_input[5776:5783] = '{32'h424b8b90, 32'hc24d0e53, 32'hc2a92c29, 32'h40660c15, 32'hc2a85a1d, 32'hc2b8f586, 32'h42b8a772, 32'hc268298c};
test_output[722] = '{32'h42b8a772};
test_index[722] = '{6};
test_input[5784:5791] = '{32'h41f32181, 32'h428ab411, 32'hc1ac1e8b, 32'h41f32d25, 32'h41ab6bc0, 32'h41c3ba20, 32'h413c8685, 32'hc2c71c23};
test_output[723] = '{32'h428ab411};
test_index[723] = '{1};
test_input[5792:5799] = '{32'h428dc081, 32'hc294720e, 32'h41ee75ab, 32'hc24df0a9, 32'h418590f1, 32'hc05c6858, 32'h411d1d1a, 32'hc25d9854};
test_output[724] = '{32'h428dc081};
test_index[724] = '{0};
test_input[5800:5807] = '{32'h421448b1, 32'h428750c9, 32'h4280c41f, 32'h423d52df, 32'hc2904d1b, 32'hc29a0ab2, 32'h427f43ef, 32'hc2b1b58a};
test_output[725] = '{32'h428750c9};
test_index[725] = '{1};
test_input[5808:5815] = '{32'hc26a1798, 32'h41f41ac8, 32'h41d677d8, 32'h41d61d28, 32'h42b9f952, 32'hc21e1020, 32'h426d9647, 32'hc2a56004};
test_output[726] = '{32'h42b9f952};
test_index[726] = '{4};
test_input[5816:5823] = '{32'h4202cc27, 32'hc2058ede, 32'h41b4a3c5, 32'hc2835f0b, 32'h4192afc7, 32'h40839440, 32'hc29dae77, 32'h401990cc};
test_output[727] = '{32'h4202cc27};
test_index[727] = '{0};
test_input[5824:5831] = '{32'hc2949a15, 32'hc2926116, 32'hc25cb283, 32'hc1044f38, 32'hc10ff2ec, 32'h429955a1, 32'h40cb1d68, 32'h42834d43};
test_output[728] = '{32'h429955a1};
test_index[728] = '{5};
test_input[5832:5839] = '{32'hc18addfc, 32'hc14ed0a4, 32'h428b76c4, 32'hc2b77d0d, 32'hc27a0cf5, 32'hc134bd97, 32'hc244b2cd, 32'h426e1ed3};
test_output[729] = '{32'h428b76c4};
test_index[729] = '{2};
test_input[5840:5847] = '{32'h4287ee7d, 32'h426f12b1, 32'hc2c4cc39, 32'hc21aeda4, 32'h4212c447, 32'h4223650b, 32'h42a65aaa, 32'hc20880b2};
test_output[730] = '{32'h42a65aaa};
test_index[730] = '{6};
test_input[5848:5855] = '{32'hc203a319, 32'h3f9c9c4e, 32'h42c6ac16, 32'hbef24890, 32'h421db0e8, 32'h4185bf2d, 32'h4284ad0f, 32'h41dd46ff};
test_output[731] = '{32'h42c6ac16};
test_index[731] = '{2};
test_input[5856:5863] = '{32'h413bf38c, 32'h4286fa4b, 32'hc1761378, 32'h41e4ffdb, 32'h413f5a14, 32'h41d4e613, 32'hc1a80868, 32'h42a29f0e};
test_output[732] = '{32'h42a29f0e};
test_index[732] = '{7};
test_input[5864:5871] = '{32'h40f70492, 32'h42c59059, 32'hc231e908, 32'hc2b7d327, 32'h42408867, 32'hc1bc0643, 32'h42236620, 32'h4231f53b};
test_output[733] = '{32'h42c59059};
test_index[733] = '{1};
test_input[5872:5879] = '{32'hc294bb1f, 32'hc022c0b2, 32'h41d3dec7, 32'hc284758c, 32'h429f11b3, 32'h42a65b8e, 32'h42415d6f, 32'h40ee1ace};
test_output[734] = '{32'h42a65b8e};
test_index[734] = '{5};
test_input[5880:5887] = '{32'h4275e409, 32'h428621f4, 32'h4234ca4a, 32'h427d00eb, 32'hc29f741a, 32'hc2a5b4af, 32'h4264a04d, 32'h4276a94f};
test_output[735] = '{32'h428621f4};
test_index[735] = '{1};
test_input[5888:5895] = '{32'hc2abb2f0, 32'h420efcf3, 32'h413b13aa, 32'hc24c1f94, 32'h42a09073, 32'h41ac31d1, 32'h40f71058, 32'h42b12d41};
test_output[736] = '{32'h42b12d41};
test_index[736] = '{7};
test_input[5896:5903] = '{32'hc2a96e84, 32'hc251642a, 32'h41cc2d9f, 32'h42a5a9cc, 32'hc23201fc, 32'h4141330b, 32'h42a04bab, 32'hc293e66f};
test_output[737] = '{32'h42a5a9cc};
test_index[737] = '{3};
test_input[5904:5911] = '{32'h4202d4bb, 32'hc1d2ebbb, 32'hc23ff89b, 32'h428223bf, 32'h42802edf, 32'hc1ddc2cd, 32'h4280f6c2, 32'h40212fbb};
test_output[738] = '{32'h428223bf};
test_index[738] = '{3};
test_input[5912:5919] = '{32'h410a7171, 32'h41c878aa, 32'h42afa058, 32'h42a30c77, 32'hc20f6eaa, 32'h427fa6c6, 32'h42198a14, 32'h42077c7b};
test_output[739] = '{32'h42afa058};
test_index[739] = '{2};
test_input[5920:5927] = '{32'hc2914401, 32'hc0cc90d4, 32'h427691f7, 32'h42602889, 32'h423cc856, 32'h418fcb15, 32'hc11dc5b0, 32'hc1949c6c};
test_output[740] = '{32'h427691f7};
test_index[740] = '{2};
test_input[5928:5935] = '{32'h408b9c35, 32'h42313ab2, 32'h42922c92, 32'h42745acd, 32'h42b830cb, 32'h42738d69, 32'h42b43e5c, 32'hc2ba2188};
test_output[741] = '{32'h42b830cb};
test_index[741] = '{4};
test_input[5936:5943] = '{32'hc0a50ea2, 32'hc1ebc8a9, 32'hc2c6e045, 32'h4224c869, 32'hc1edfd99, 32'h421ecc72, 32'hc0a8cadf, 32'hc2578838};
test_output[742] = '{32'h4224c869};
test_index[742] = '{3};
test_input[5944:5951] = '{32'hc281356c, 32'hc1119ae0, 32'hc185aaf5, 32'h424c9251, 32'hc234570c, 32'hc283b5eb, 32'h42282c98, 32'h42a94a5b};
test_output[743] = '{32'h42a94a5b};
test_index[743] = '{7};
test_input[5952:5959] = '{32'hc004dc3a, 32'h42457f8f, 32'hc2bc335b, 32'h42694d6b, 32'h420d16d6, 32'hc129913f, 32'h4273a192, 32'hc2b30db4};
test_output[744] = '{32'h4273a192};
test_index[744] = '{6};
test_input[5960:5967] = '{32'hc00c69de, 32'h422b93e4, 32'hc1981cfc, 32'hc238e5bd, 32'h428a4397, 32'h425e3e39, 32'h41df6ede, 32'hc223b6bc};
test_output[745] = '{32'h428a4397};
test_index[745] = '{4};
test_input[5968:5975] = '{32'h428ea355, 32'h42b3c815, 32'h41deb302, 32'h429dc96e, 32'h426d5c92, 32'h425c6e00, 32'hc21f2a78, 32'h41f1aba5};
test_output[746] = '{32'h42b3c815};
test_index[746] = '{1};
test_input[5976:5983] = '{32'h42982352, 32'h41874354, 32'hc1d613fc, 32'h417b6d7f, 32'hc2b0214c, 32'hc27c0ea1, 32'h41f2d5b6, 32'h42b8904c};
test_output[747] = '{32'h42b8904c};
test_index[747] = '{7};
test_input[5984:5991] = '{32'hc1a4c4f2, 32'h42ba079b, 32'hc27f2636, 32'hc286a66f, 32'h428ee8c0, 32'hc2bbb0b5, 32'hc286dd93, 32'h4257dccb};
test_output[748] = '{32'h42ba079b};
test_index[748] = '{1};
test_input[5992:5999] = '{32'hc255f2b9, 32'hc27c42df, 32'hc23ea690, 32'h42b09bd4, 32'h42a15901, 32'h41130e51, 32'h4216ef55, 32'hc2c01205};
test_output[749] = '{32'h42b09bd4};
test_index[749] = '{3};
test_input[6000:6007] = '{32'h42bf5ab5, 32'hc1602ce8, 32'hc208cd69, 32'hc26b69f9, 32'hc1d497d2, 32'hc15cb326, 32'hc1644926, 32'h42a9a66f};
test_output[750] = '{32'h42bf5ab5};
test_index[750] = '{0};
test_input[6008:6015] = '{32'hc228626f, 32'hc226786f, 32'hc266e50c, 32'h423bdd0b, 32'hc24c9117, 32'hc2781f2e, 32'hc25a5a17, 32'hc240ec64};
test_output[751] = '{32'h423bdd0b};
test_index[751] = '{3};
test_input[6016:6023] = '{32'h4244691b, 32'h42ab984f, 32'h42147ece, 32'hc291b359, 32'hc2272f61, 32'h42b15aba, 32'h418caa0e, 32'h41ec55f0};
test_output[752] = '{32'h42b15aba};
test_index[752] = '{5};
test_input[6024:6031] = '{32'hc2c7ce35, 32'h42583c8f, 32'h42b158a9, 32'hc28b4ee9, 32'hc09f8856, 32'hc2954dc0, 32'hc212f6d9, 32'hc2ad7ad9};
test_output[753] = '{32'h42b158a9};
test_index[753] = '{2};
test_input[6032:6039] = '{32'hc1f12a38, 32'hc25e3d9b, 32'h423899cd, 32'h424a898b, 32'h42991ae1, 32'hc031dbf6, 32'h428058d7, 32'h421dcd2a};
test_output[754] = '{32'h42991ae1};
test_index[754] = '{4};
test_input[6040:6047] = '{32'h421112d5, 32'h41e2a906, 32'h426c4c72, 32'h3fc03b08, 32'hbfc7f8d1, 32'hc19a29cb, 32'hc2c5aa83, 32'h42aa2ea5};
test_output[755] = '{32'h42aa2ea5};
test_index[755] = '{7};
test_input[6048:6055] = '{32'hc26103aa, 32'h42549219, 32'hc21450cd, 32'hc2163510, 32'h42920df5, 32'hc28f81ed, 32'hc204a993, 32'hc2a161d4};
test_output[756] = '{32'h42920df5};
test_index[756] = '{4};
test_input[6056:6063] = '{32'h41c75905, 32'hc1610243, 32'hc194dba3, 32'hc26efc4e, 32'h42aff377, 32'hc21ab009, 32'h42a4733c, 32'hc2663b82};
test_output[757] = '{32'h42aff377};
test_index[757] = '{4};
test_input[6064:6071] = '{32'h42597b2f, 32'hc197b4b9, 32'hc2ba19a8, 32'h42874463, 32'h42a5dac0, 32'h42696dfa, 32'hc294ed53, 32'hc2a5363a};
test_output[758] = '{32'h42a5dac0};
test_index[758] = '{4};
test_input[6072:6079] = '{32'hc24f67a7, 32'hc239fe4c, 32'h4297784e, 32'hbe9add73, 32'hc2ab3751, 32'hc09bfa7f, 32'h42c4c802, 32'hc1b24790};
test_output[759] = '{32'h42c4c802};
test_index[759] = '{6};
test_input[6080:6087] = '{32'h4272149e, 32'hc23af568, 32'hc29352ea, 32'hc21d6946, 32'h419ceee9, 32'hc12febfb, 32'h41e4e74d, 32'hc1c1423c};
test_output[760] = '{32'h4272149e};
test_index[760] = '{0};
test_input[6088:6095] = '{32'hc2a75cb6, 32'h42847e28, 32'hc15fb82a, 32'hc293f570, 32'h4269b8df, 32'hc241958c, 32'hc102186a, 32'h41d5b560};
test_output[761] = '{32'h42847e28};
test_index[761] = '{1};
test_input[6096:6103] = '{32'hc2040eca, 32'h42bdd123, 32'h4065ae70, 32'hc0363914, 32'h42badf82, 32'h421afc96, 32'h4219c47e, 32'h4272e1aa};
test_output[762] = '{32'h42bdd123};
test_index[762] = '{1};
test_input[6104:6111] = '{32'hc2452a5b, 32'hc1e9f588, 32'hc17f5821, 32'h4255b08b, 32'h42355c89, 32'hc1a8f535, 32'hc20c6d26, 32'hc20fdffe};
test_output[763] = '{32'h4255b08b};
test_index[763] = '{3};
test_input[6112:6119] = '{32'h4299804f, 32'h40237472, 32'h42b0243f, 32'hc2044414, 32'h422bc6a2, 32'hc21b5cb0, 32'hc263d28b, 32'hc2bdda02};
test_output[764] = '{32'h42b0243f};
test_index[764] = '{2};
test_input[6120:6127] = '{32'h41fe10ee, 32'h40e211c9, 32'hc1634adf, 32'hc299e79d, 32'hc283534c, 32'h42169b20, 32'hc078a97d, 32'h42c72eaf};
test_output[765] = '{32'h42c72eaf};
test_index[765] = '{7};
test_input[6128:6135] = '{32'h42416467, 32'h42c4fc69, 32'h42219f4e, 32'hc242c51c, 32'h428fb1b4, 32'hc209e13b, 32'hc292c844, 32'hc253fe1c};
test_output[766] = '{32'h42c4fc69};
test_index[766] = '{1};
test_input[6136:6143] = '{32'h4171001b, 32'hc21cd11e, 32'hc27c71d8, 32'h42c44670, 32'h42115d01, 32'hbfa9f867, 32'h4239345d, 32'hc28e277f};
test_output[767] = '{32'h42c44670};
test_index[767] = '{3};
test_input[6144:6151] = '{32'hc2774599, 32'hc29928f3, 32'h41c35abf, 32'hc0b0590d, 32'hc13dedce, 32'h42a3a339, 32'h42b0cbc0, 32'hc292c8e6};
test_output[768] = '{32'h42b0cbc0};
test_index[768] = '{6};
test_input[6152:6159] = '{32'hc2751686, 32'h410cfa33, 32'h42c22857, 32'h419ab774, 32'hc27ec632, 32'h41ca58f0, 32'hc2781b9e, 32'h428deaa0};
test_output[769] = '{32'h42c22857};
test_index[769] = '{2};
test_input[6160:6167] = '{32'hc28f281e, 32'hc282fe7e, 32'h423f1094, 32'hc147a519, 32'h429fbec7, 32'h42a7d22a, 32'h425398d4, 32'h41e22751};
test_output[770] = '{32'h42a7d22a};
test_index[770] = '{5};
test_input[6168:6175] = '{32'hc221e12f, 32'h427db03b, 32'hc2248ee9, 32'h42b85294, 32'hc2418170, 32'hc27d32e8, 32'h42966b3f, 32'h42c412b2};
test_output[771] = '{32'h42c412b2};
test_index[771] = '{7};
test_input[6176:6183] = '{32'hc2519a1e, 32'hc18dbcbf, 32'h42b809bd, 32'h422928ee, 32'hc29f5cf3, 32'h404823ea, 32'h42b1b057, 32'h40124b18};
test_output[772] = '{32'h42b809bd};
test_index[772] = '{2};
test_input[6184:6191] = '{32'h42471d23, 32'hc1a29494, 32'h4240a166, 32'h4214b5e5, 32'hc289a722, 32'hc2429e46, 32'h42b7a29a, 32'hc2c518e2};
test_output[773] = '{32'h42b7a29a};
test_index[773] = '{6};
test_input[6192:6199] = '{32'h4257b35b, 32'h42b9e694, 32'hc18124db, 32'h411881ca, 32'hc21dffef, 32'h42547240, 32'h411c4eca, 32'hc28e38fd};
test_output[774] = '{32'h42b9e694};
test_index[774] = '{1};
test_input[6200:6207] = '{32'h42bcbe9f, 32'hc233f890, 32'hc27fadb0, 32'hc2167f27, 32'h42943181, 32'h4255f25c, 32'h41aa0991, 32'h410432db};
test_output[775] = '{32'h42bcbe9f};
test_index[775] = '{0};
test_input[6208:6215] = '{32'h42c3bf43, 32'h42648abc, 32'hc180105d, 32'hc24ec993, 32'hc2af3e33, 32'hc1320163, 32'h41892a16, 32'hc2897d82};
test_output[776] = '{32'h42c3bf43};
test_index[776] = '{0};
test_input[6216:6223] = '{32'hc2ba3dbd, 32'hc2c5a062, 32'hc2a6c90f, 32'h4183cefe, 32'hc2984d4b, 32'hc2af4272, 32'hc184c864, 32'hc1aec586};
test_output[777] = '{32'h4183cefe};
test_index[777] = '{3};
test_input[6224:6231] = '{32'hc2a2c935, 32'hc2b1bdbe, 32'hc2ab5355, 32'h41aff8bb, 32'hc2b61663, 32'h4282b1e2, 32'h418f2f8f, 32'hc1c640cc};
test_output[778] = '{32'h4282b1e2};
test_index[778] = '{5};
test_input[6232:6239] = '{32'h42a947a3, 32'hc2272308, 32'h42a67ccf, 32'h412b0b05, 32'h42c210e6, 32'h41c55f3d, 32'h425a3bea, 32'h41d729dd};
test_output[779] = '{32'h42c210e6};
test_index[779] = '{4};
test_input[6240:6247] = '{32'hc22fe6b7, 32'hc2a91080, 32'hc20410bf, 32'hc1ce13d2, 32'h412ea46d, 32'hc25c7bb1, 32'hc28ae22a, 32'h41176a74};
test_output[780] = '{32'h412ea46d};
test_index[780] = '{4};
test_input[6248:6255] = '{32'h428f54e1, 32'h42bb467e, 32'hc0731b29, 32'h410b59ec, 32'hc24ec3cc, 32'h412c1edf, 32'h428c3e96, 32'h424e7a18};
test_output[781] = '{32'h42bb467e};
test_index[781] = '{1};
test_input[6256:6263] = '{32'h4264d103, 32'hc22a72b8, 32'hc2194bc0, 32'h42b0d35b, 32'hc22a9019, 32'h40fd3c09, 32'hc2800ba9, 32'h42ae6bd0};
test_output[782] = '{32'h42b0d35b};
test_index[782] = '{3};
test_input[6264:6271] = '{32'hc2ab07d6, 32'h41d618b8, 32'h42685b7b, 32'h42b6ff9e, 32'hc291aba0, 32'hc28901bb, 32'h423798e9, 32'h42c20f6a};
test_output[783] = '{32'h42c20f6a};
test_index[783] = '{7};
test_input[6272:6279] = '{32'hc1877feb, 32'hc185d96e, 32'hc253d9f1, 32'hc23e9178, 32'h42293525, 32'h414af0fb, 32'h429cef39, 32'h429dce50};
test_output[784] = '{32'h429dce50};
test_index[784] = '{7};
test_input[6280:6287] = '{32'hc1aaa037, 32'h4040d859, 32'hc200f23e, 32'hc167dcdd, 32'hc2b4f48d, 32'hc223cb42, 32'hc16a0661, 32'hc2be697f};
test_output[785] = '{32'h4040d859};
test_index[785] = '{1};
test_input[6288:6295] = '{32'hc253bdf9, 32'hc29533f6, 32'h42c78a34, 32'h4035bd53, 32'hc22a2aaa, 32'h41577d75, 32'h4176eb98, 32'h4250234a};
test_output[786] = '{32'h42c78a34};
test_index[786] = '{2};
test_input[6296:6303] = '{32'hc254f34d, 32'h41af9b20, 32'h4283340b, 32'h4178c698, 32'h4087d1a2, 32'h4052ed3c, 32'hc2c7d95e, 32'h42022105};
test_output[787] = '{32'h4283340b};
test_index[787] = '{2};
test_input[6304:6311] = '{32'hc2aa0053, 32'h42ac6e6c, 32'h4186a211, 32'h42b18ba8, 32'h42c509ec, 32'h422a4243, 32'hc2afc679, 32'h41ae1116};
test_output[788] = '{32'h42c509ec};
test_index[788] = '{4};
test_input[6312:6319] = '{32'h418f91f9, 32'hc1ad7d19, 32'h41ac5452, 32'hc2af6d55, 32'h41d10cf9, 32'hc27c7024, 32'hc29a3513, 32'h4199738e};
test_output[789] = '{32'h41d10cf9};
test_index[789] = '{4};
test_input[6320:6327] = '{32'h42c17e01, 32'hc010ec9f, 32'hc0c6cdb3, 32'h428c4ca1, 32'h423d9480, 32'h420c3cb0, 32'hc2814a70, 32'h42c4bab8};
test_output[790] = '{32'h42c4bab8};
test_index[790] = '{7};
test_input[6328:6335] = '{32'hc29474ce, 32'h42990ac2, 32'h4285e44f, 32'hc1d5dde6, 32'hc294e875, 32'hc2b628be, 32'hc19058e8, 32'h424f2a7d};
test_output[791] = '{32'h42990ac2};
test_index[791] = '{1};
test_input[6336:6343] = '{32'h423408ff, 32'h42c2c90d, 32'hc20de096, 32'h423fb084, 32'hc29c293a, 32'hc2be0b39, 32'hc28c247e, 32'h416068c0};
test_output[792] = '{32'h42c2c90d};
test_index[792] = '{1};
test_input[6344:6351] = '{32'hc270687b, 32'h4196bfcb, 32'hbff7d057, 32'h41d740ee, 32'h4243713e, 32'hc039c001, 32'h41ce19fd, 32'h428253cd};
test_output[793] = '{32'h428253cd};
test_index[793] = '{7};
test_input[6352:6359] = '{32'h4225312e, 32'h41e5ef7d, 32'h423a4b41, 32'hc208a18a, 32'hc28568cd, 32'hc1c28614, 32'hc2b3a113, 32'h4270f817};
test_output[794] = '{32'h4270f817};
test_index[794] = '{7};
test_input[6360:6367] = '{32'h42033c53, 32'h4218441e, 32'h41ada518, 32'hc28a46ee, 32'hc1ffe843, 32'hc1f24269, 32'h4222cbdd, 32'hc1eab300};
test_output[795] = '{32'h4222cbdd};
test_index[795] = '{6};
test_input[6368:6375] = '{32'hc25ff9b8, 32'h3f5f1d2b, 32'h42b414e6, 32'hc2c75e68, 32'h415744cb, 32'h42123b7e, 32'h425e4e25, 32'hc14b77e5};
test_output[796] = '{32'h42b414e6};
test_index[796] = '{2};
test_input[6376:6383] = '{32'h42814343, 32'hc2503e90, 32'hc29ea7a8, 32'h42acd0cb, 32'hbfcf99f4, 32'hc2817ed5, 32'hc09a25ac, 32'hc2c4a01c};
test_output[797] = '{32'h42acd0cb};
test_index[797] = '{3};
test_input[6384:6391] = '{32'h422b82f8, 32'h42991e14, 32'hc2357984, 32'hc230af81, 32'hc2b0bbae, 32'h41fb41b9, 32'h42921bb7, 32'hc0c2fa02};
test_output[798] = '{32'h42991e14};
test_index[798] = '{1};
test_input[6392:6399] = '{32'h42295c43, 32'h42891a8a, 32'hc236d69f, 32'hc15e9fbe, 32'h42897e7f, 32'hc2b2107d, 32'h40e51903, 32'hc2afef0c};
test_output[799] = '{32'h42897e7f};
test_index[799] = '{4};
test_input[6400:6407] = '{32'hc201cf19, 32'h429400b3, 32'hc2440b6d, 32'hc2a83328, 32'hc25496c6, 32'h42259c07, 32'h429d8c82, 32'h42be89f7};
test_output[800] = '{32'h42be89f7};
test_index[800] = '{7};
test_input[6408:6415] = '{32'hc258f231, 32'hc19b67d3, 32'hc22265fa, 32'h41e042dd, 32'hc127a8f4, 32'h4296e562, 32'hc2bcce9f, 32'hc2bf1d44};
test_output[801] = '{32'h4296e562};
test_index[801] = '{5};
test_input[6416:6423] = '{32'hc29ca432, 32'h4287249e, 32'hc194885f, 32'h419b4361, 32'hc2020306, 32'h424dfa02, 32'hc06c2db3, 32'h4174f054};
test_output[802] = '{32'h4287249e};
test_index[802] = '{1};
test_input[6424:6431] = '{32'h3f5c5018, 32'hc2ab4fbf, 32'h426aa2bc, 32'h41ecd2f9, 32'hc2a1374a, 32'h429168f6, 32'h41111442, 32'hc24ee2ca};
test_output[803] = '{32'h429168f6};
test_index[803] = '{5};
test_input[6432:6439] = '{32'h424395ee, 32'hc2a89af2, 32'h42addcf3, 32'h42320681, 32'h417b2488, 32'hc2546551, 32'hc23d4a6d, 32'h41795a5e};
test_output[804] = '{32'h42addcf3};
test_index[804] = '{2};
test_input[6440:6447] = '{32'hc26417f3, 32'h411943a8, 32'h417ee78a, 32'h42637e9b, 32'hc1143dba, 32'hc21ac38a, 32'hc1d85f69, 32'hc244587e};
test_output[805] = '{32'h42637e9b};
test_index[805] = '{3};
test_input[6448:6455] = '{32'hc27ea93c, 32'hc2b61701, 32'hc2117781, 32'hc2aec66d, 32'h423a6001, 32'hc2aa5918, 32'hc2b92570, 32'hbfc52872};
test_output[806] = '{32'h423a6001};
test_index[806] = '{4};
test_input[6456:6463] = '{32'hc1d524c9, 32'h42b8f8d9, 32'h420d39bd, 32'hc044f81f, 32'h4105ece8, 32'h422ca74a, 32'hc2b81c99, 32'h415cf72f};
test_output[807] = '{32'h42b8f8d9};
test_index[807] = '{1};
test_input[6464:6471] = '{32'h41b8580c, 32'h425276f5, 32'hc29c76bf, 32'hc1dc82b3, 32'h42a93356, 32'h429fa7a6, 32'h40cc9f3f, 32'h4141038f};
test_output[808] = '{32'h42a93356};
test_index[808] = '{4};
test_input[6472:6479] = '{32'h41e8e2dc, 32'hc288c733, 32'h422b52cf, 32'hc232a563, 32'h422f18de, 32'h41df1abb, 32'h40b99ed2, 32'h41d9778c};
test_output[809] = '{32'h422f18de};
test_index[809] = '{4};
test_input[6480:6487] = '{32'h422ca2f9, 32'hc13e8cf8, 32'hc2b74271, 32'h42be8f58, 32'hc236e799, 32'hc2906c14, 32'h4234a2f3, 32'hc2b476e1};
test_output[810] = '{32'h42be8f58};
test_index[810] = '{3};
test_input[6488:6495] = '{32'h42c02cae, 32'h41ed6d70, 32'hc2775bec, 32'hc235abce, 32'hc07e4e24, 32'h420ea260, 32'h424a7a33, 32'h429c36b7};
test_output[811] = '{32'h42c02cae};
test_index[811] = '{0};
test_input[6496:6503] = '{32'hc2a572dd, 32'h417f6c72, 32'h428816ff, 32'h41d15155, 32'hc28b12f9, 32'hc1821a66, 32'h428f8200, 32'hc1a4c501};
test_output[812] = '{32'h428f8200};
test_index[812] = '{6};
test_input[6504:6511] = '{32'hc27fd0e0, 32'hc04a560c, 32'hc200a0b4, 32'h42c4c57b, 32'h4283c781, 32'h4293b0ff, 32'hc29b5d31, 32'h42419247};
test_output[813] = '{32'h42c4c57b};
test_index[813] = '{3};
test_input[6512:6519] = '{32'hc28fa560, 32'hc1b59dee, 32'h42a674e6, 32'h429c95f4, 32'hc26be1bc, 32'hc296a5fc, 32'h41b47ae3, 32'hc29c0959};
test_output[814] = '{32'h42a674e6};
test_index[814] = '{2};
test_input[6520:6527] = '{32'hc21d6e71, 32'hc2a9beef, 32'hc2c6fd59, 32'hc20e783c, 32'hc20b6a86, 32'h4157be21, 32'h4196f7f4, 32'h40e7642d};
test_output[815] = '{32'h4196f7f4};
test_index[815] = '{6};
test_input[6528:6535] = '{32'hc2c09671, 32'hc29c3936, 32'hc1f3aea2, 32'h4261ec87, 32'hc217b5a0, 32'hc2318f89, 32'hc28f88a7, 32'h42c7511e};
test_output[816] = '{32'h42c7511e};
test_index[816] = '{7};
test_input[6536:6543] = '{32'hc23fbd53, 32'h42bd3c1b, 32'hc24f512b, 32'h41f53c9b, 32'hc2bee566, 32'hc1ddd489, 32'hc1a070e6, 32'h42c081d2};
test_output[817] = '{32'h42c081d2};
test_index[817] = '{7};
test_input[6544:6551] = '{32'h428f9b83, 32'h42c5548f, 32'h40e48668, 32'hc24ef337, 32'hc2824dc1, 32'hc1d18c27, 32'hc2070f11, 32'hc200a2be};
test_output[818] = '{32'h42c5548f};
test_index[818] = '{1};
test_input[6552:6559] = '{32'h42acc29f, 32'h429550cc, 32'h418328f3, 32'hc14d7738, 32'hc21f4709, 32'h42b9004a, 32'h427322ac, 32'hc209172f};
test_output[819] = '{32'h42b9004a};
test_index[819] = '{5};
test_input[6560:6567] = '{32'h421cefbc, 32'h40c14ec2, 32'hc2c0698f, 32'h42936b19, 32'hc0e91dfe, 32'hc2a3d98e, 32'hc2b1a968, 32'hc29e024c};
test_output[820] = '{32'h42936b19};
test_index[820] = '{3};
test_input[6568:6575] = '{32'h41726b6f, 32'h42bd165a, 32'hc1d29163, 32'hc179a6ee, 32'h4224ceae, 32'h428bf830, 32'hc20cd8ff, 32'h42c7b916};
test_output[821] = '{32'h42c7b916};
test_index[821] = '{7};
test_input[6576:6583] = '{32'h41c903c5, 32'hc1ed4128, 32'hc1b8eced, 32'hc28d8e06, 32'hc2687943, 32'hc2b253df, 32'hc1d31a24, 32'hc209ec02};
test_output[822] = '{32'h41c903c5};
test_index[822] = '{0};
test_input[6584:6591] = '{32'h42a936e0, 32'h4286c5e2, 32'hc18e64fa, 32'h42494aa2, 32'hc192d66f, 32'h41c321a8, 32'h40ef847f, 32'hc14ea504};
test_output[823] = '{32'h42a936e0};
test_index[823] = '{0};
test_input[6592:6599] = '{32'h415a51a2, 32'hc2413c97, 32'hc298e68e, 32'hc2751f75, 32'h41606eb3, 32'h42be57db, 32'hc28a89eb, 32'h4154f897};
test_output[824] = '{32'h42be57db};
test_index[824] = '{5};
test_input[6600:6607] = '{32'h4296202f, 32'hc29e6e6d, 32'hc26f5b4a, 32'hc2a4e35e, 32'hc20290bf, 32'hc27dc89e, 32'hc2122092, 32'hc29e4cd5};
test_output[825] = '{32'h4296202f};
test_index[825] = '{0};
test_input[6608:6615] = '{32'h42342967, 32'hc1ac2df5, 32'hc1ede8a3, 32'hc1aec8b4, 32'h4282a2d8, 32'h42b9222b, 32'hc28e48c8, 32'h42a7bce1};
test_output[826] = '{32'h42b9222b};
test_index[826] = '{5};
test_input[6616:6623] = '{32'h4227656d, 32'h42ad457e, 32'h422e7951, 32'h429f9980, 32'h4232f20d, 32'h4279cf7a, 32'h41a0b9f0, 32'hc20bd157};
test_output[827] = '{32'h42ad457e};
test_index[827] = '{1};
test_input[6624:6631] = '{32'hc18049ba, 32'h42b7e98d, 32'h415690f6, 32'hc227e5b8, 32'h41df28ba, 32'h425477ba, 32'h416e1aaf, 32'hc2537c9d};
test_output[828] = '{32'h42b7e98d};
test_index[828] = '{1};
test_input[6632:6639] = '{32'h42a5e735, 32'hc24581d7, 32'hc2b5f55e, 32'hc2b33edb, 32'h428f3837, 32'h42c730fa, 32'h42b9f21c, 32'hc27996e3};
test_output[829] = '{32'h42c730fa};
test_index[829] = '{5};
test_input[6640:6647] = '{32'h4152167c, 32'h41b732ca, 32'h426ba4d7, 32'h3f7e2c11, 32'h423bd592, 32'hc21cca97, 32'hc278f76e, 32'hc2933454};
test_output[830] = '{32'h426ba4d7};
test_index[830] = '{2};
test_input[6648:6655] = '{32'hc2ba634b, 32'hc2a946b3, 32'hc29307af, 32'hc06fc0f7, 32'h4130085d, 32'hc145fadc, 32'h41094199, 32'hc28e4f36};
test_output[831] = '{32'h4130085d};
test_index[831] = '{4};
test_input[6656:6663] = '{32'hc2ab709d, 32'h41c06fc3, 32'h42b33925, 32'h428ae5d1, 32'h4284d59a, 32'hc22dbe06, 32'h427620f2, 32'h4258720e};
test_output[832] = '{32'h42b33925};
test_index[832] = '{2};
test_input[6664:6671] = '{32'hc239ea71, 32'hc18fe28c, 32'h42136933, 32'hc2b786b4, 32'hc264b873, 32'h41e2cad5, 32'h42c20bc6, 32'hc2aae7b3};
test_output[833] = '{32'h42c20bc6};
test_index[833] = '{6};
test_input[6672:6679] = '{32'hc16c24eb, 32'h42171424, 32'h41deba11, 32'hc2814344, 32'h3fa058a5, 32'h409ee778, 32'h429d0c3b, 32'h41083ebb};
test_output[834] = '{32'h429d0c3b};
test_index[834] = '{6};
test_input[6680:6687] = '{32'hc227ad95, 32'hc2802375, 32'h420ae982, 32'hc2a9d3b6, 32'h422e3d65, 32'h41a440a2, 32'hc21e3ebb, 32'h40da45f1};
test_output[835] = '{32'h422e3d65};
test_index[835] = '{4};
test_input[6688:6695] = '{32'h41b4384d, 32'h42984051, 32'h4260cc9e, 32'hc2514a3e, 32'h42762c0e, 32'hc2984983, 32'h41c0e4b4, 32'h401e5ce1};
test_output[836] = '{32'h42984051};
test_index[836] = '{1};
test_input[6696:6703] = '{32'hc0939d54, 32'hc0c310c6, 32'h429a0e63, 32'h41c48d10, 32'h422fdefa, 32'hc2473614, 32'h42b19ff1, 32'hc23e5637};
test_output[837] = '{32'h42b19ff1};
test_index[837] = '{6};
test_input[6704:6711] = '{32'hc2bfa187, 32'h42c1ffd6, 32'h42ad922b, 32'h42bb8b14, 32'hc29f161b, 32'h424909f5, 32'hc1623ed5, 32'hc1c1247c};
test_output[838] = '{32'h42c1ffd6};
test_index[838] = '{1};
test_input[6712:6719] = '{32'h42c35b05, 32'h42325678, 32'h429797eb, 32'h41e201e8, 32'hc2b02171, 32'h42917b1e, 32'h42a3d9cc, 32'h429916d6};
test_output[839] = '{32'h42c35b05};
test_index[839] = '{0};
test_input[6720:6727] = '{32'h4223ca57, 32'hc13e8d54, 32'hc18836d1, 32'h42b0ffc3, 32'h40a55ecd, 32'hc28aa8a3, 32'hc294a355, 32'hc2c428c9};
test_output[840] = '{32'h42b0ffc3};
test_index[840] = '{3};
test_input[6728:6735] = '{32'hc142184a, 32'h4047ede9, 32'hc2827a4b, 32'hc2adfbd3, 32'h41bea7c6, 32'h415eb9f3, 32'hc21cfb5f, 32'hc1bb5df4};
test_output[841] = '{32'h41bea7c6};
test_index[841] = '{4};
test_input[6736:6743] = '{32'hc266a914, 32'h40a8a759, 32'hc2be2a5e, 32'h423c9f99, 32'h42630e7f, 32'h429aeee3, 32'h414d8a90, 32'hc1e48e1c};
test_output[842] = '{32'h429aeee3};
test_index[842] = '{5};
test_input[6744:6751] = '{32'hc2b77be9, 32'hbefe1c70, 32'h41f691f5, 32'h42c5df61, 32'hc2a81dff, 32'hc1ae4c90, 32'h428a8cec, 32'hc2c61b46};
test_output[843] = '{32'h42c5df61};
test_index[843] = '{3};
test_input[6752:6759] = '{32'h424f3f56, 32'h41bcae64, 32'h412f2243, 32'hc082adcf, 32'hc2c7a8ac, 32'hc299645a, 32'hc2b07340, 32'h42bf88d0};
test_output[844] = '{32'h42bf88d0};
test_index[844] = '{7};
test_input[6760:6767] = '{32'hc22e3a39, 32'hc20f7e23, 32'hc2aa2cba, 32'h4279a42b, 32'h41d79d52, 32'hc1044069, 32'h4292d874, 32'hc24e453a};
test_output[845] = '{32'h4292d874};
test_index[845] = '{6};
test_input[6768:6775] = '{32'hc26492a5, 32'hc238731b, 32'hc270b06e, 32'hc2039130, 32'h4281f01c, 32'h422eb16f, 32'h419aa4fb, 32'h4195136f};
test_output[846] = '{32'h4281f01c};
test_index[846] = '{4};
test_input[6776:6783] = '{32'hc2ba930c, 32'h4222dd96, 32'h42bd7622, 32'h42c6d83d, 32'h424327c4, 32'h4290829a, 32'h42a6f5fd, 32'hc212be83};
test_output[847] = '{32'h42c6d83d};
test_index[847] = '{3};
test_input[6784:6791] = '{32'h427d0c29, 32'hc2b9a48a, 32'hc1853eca, 32'h42563ef9, 32'hc2522847, 32'hc10eb0ab, 32'hc027e039, 32'hc2a264dd};
test_output[848] = '{32'h427d0c29};
test_index[848] = '{0};
test_input[6792:6799] = '{32'hc126c75b, 32'h425fb0f7, 32'h42c6e961, 32'h4292a781, 32'hc2a5f1e3, 32'hc280cb65, 32'hc162b516, 32'h41abd882};
test_output[849] = '{32'h42c6e961};
test_index[849] = '{2};
test_input[6800:6807] = '{32'hbeea2480, 32'h42484502, 32'h41d9bfae, 32'hc1d948de, 32'hc29a669d, 32'h42950b52, 32'h422a71cf, 32'h424803b0};
test_output[850] = '{32'h42950b52};
test_index[850] = '{5};
test_input[6808:6815] = '{32'hc1bf765b, 32'hc29779f4, 32'hc137f9ec, 32'h42c31bef, 32'hc27a9185, 32'hc2857f02, 32'h40438d0d, 32'hc20ff03d};
test_output[851] = '{32'h42c31bef};
test_index[851] = '{3};
test_input[6816:6823] = '{32'h410a252f, 32'hc1a6962f, 32'h428afaa8, 32'h40c0edd2, 32'hc2ba297c, 32'hc21b4788, 32'hc2c44d05, 32'hc2b1655e};
test_output[852] = '{32'h428afaa8};
test_index[852] = '{2};
test_input[6824:6831] = '{32'h4228652e, 32'h41bd999c, 32'hc2a1f59c, 32'h41b65cd4, 32'h428aa588, 32'h41c33b9c, 32'h4261f3da, 32'h42c3a587};
test_output[853] = '{32'h42c3a587};
test_index[853] = '{7};
test_input[6832:6839] = '{32'hc1c74aa1, 32'hc252fcaa, 32'h42aaeeae, 32'hc108b504, 32'hc22de5b2, 32'hc29d38c6, 32'hc08c3626, 32'h42341864};
test_output[854] = '{32'h42aaeeae};
test_index[854] = '{2};
test_input[6840:6847] = '{32'hc2b0a951, 32'h42736b3d, 32'hc23afe78, 32'h4132ca60, 32'hc1cc5622, 32'h429e436f, 32'h4085ac60, 32'hc231c16c};
test_output[855] = '{32'h429e436f};
test_index[855] = '{5};
test_input[6848:6855] = '{32'h4132f552, 32'h426c4870, 32'h41044c61, 32'hc2180a29, 32'hc2881fee, 32'h42352f6a, 32'h41e29cf7, 32'h41c9aede};
test_output[856] = '{32'h426c4870};
test_index[856] = '{1};
test_input[6856:6863] = '{32'h42b24f59, 32'h426ed028, 32'h42aeffc4, 32'hc282219c, 32'hc2835736, 32'h4260eb87, 32'h42b743ca, 32'hc29a7b4a};
test_output[857] = '{32'h42b743ca};
test_index[857] = '{6};
test_input[6864:6871] = '{32'h429b1747, 32'h4284af30, 32'hc1dc6483, 32'hc0808814, 32'hc2697e86, 32'h4258887d, 32'h42262964, 32'h4295bab1};
test_output[858] = '{32'h429b1747};
test_index[858] = '{0};
test_input[6872:6879] = '{32'h41938c1a, 32'hc1be6ae8, 32'hc2c31d64, 32'hc287af1b, 32'hc298a15a, 32'h402bbd4c, 32'h41e8f36b, 32'h42c2160d};
test_output[859] = '{32'h42c2160d};
test_index[859] = '{7};
test_input[6880:6887] = '{32'h42beee33, 32'hc24defba, 32'h41d46b38, 32'h41b9dfe1, 32'hc28dcc54, 32'hc1758a89, 32'hc23e1e5f, 32'h420ee7f9};
test_output[860] = '{32'h42beee33};
test_index[860] = '{0};
test_input[6888:6895] = '{32'h42acf6c0, 32'h40b09abd, 32'hc2b37ca9, 32'hc24e9a59, 32'hc2c3f6a4, 32'hc25cdf6d, 32'h42a1fff2, 32'h42811850};
test_output[861] = '{32'h42acf6c0};
test_index[861] = '{0};
test_input[6896:6903] = '{32'h40d4da43, 32'h427fb67d, 32'h423a5ae5, 32'hc2343ade, 32'h42925ed8, 32'hc2beb6e8, 32'hc220b7dd, 32'h42979bf5};
test_output[862] = '{32'h42979bf5};
test_index[862] = '{7};
test_input[6904:6911] = '{32'hc2811719, 32'h3fc8339f, 32'h4243b1f8, 32'h4285e2dd, 32'hc255d68e, 32'h41be244f, 32'h429e15b0, 32'hc22f2c83};
test_output[863] = '{32'h429e15b0};
test_index[863] = '{6};
test_input[6912:6919] = '{32'hc25cbf5a, 32'h42776a7a, 32'hc1b6b24e, 32'h4203eac0, 32'h42184ec5, 32'hc288036e, 32'hc21e72f4, 32'hc2005f12};
test_output[864] = '{32'h42776a7a};
test_index[864] = '{1};
test_input[6920:6927] = '{32'hc25e1396, 32'h42b22b50, 32'hc1fc3065, 32'hc1d48f2e, 32'hc1b73aaa, 32'h42202344, 32'h42aaf474, 32'h41cf913e};
test_output[865] = '{32'h42b22b50};
test_index[865] = '{1};
test_input[6928:6935] = '{32'h429e3124, 32'h425809f8, 32'h4293f9f7, 32'hc2afd4e2, 32'h42ab7661, 32'h4206b0f0, 32'hc09b8975, 32'hc2c0d356};
test_output[866] = '{32'h42ab7661};
test_index[866] = '{4};
test_input[6936:6943] = '{32'hbfcd2113, 32'h3e457719, 32'h41cc4c39, 32'h42beba14, 32'hc20030fa, 32'h428503c2, 32'hc263fc6b, 32'h42a155bc};
test_output[867] = '{32'h42beba14};
test_index[867] = '{3};
test_input[6944:6951] = '{32'hc22d62aa, 32'hc2553190, 32'hc286e53e, 32'hc2428ed7, 32'hc0e8434b, 32'h4218b5ae, 32'h3f771b0d, 32'hc20a2e84};
test_output[868] = '{32'h4218b5ae};
test_index[868] = '{5};
test_input[6952:6959] = '{32'h41b252b8, 32'hc214e5b2, 32'h419ed5d0, 32'h422c44c1, 32'h403b64bf, 32'h422e7204, 32'hc1048d4a, 32'h42ac6bbe};
test_output[869] = '{32'h42ac6bbe};
test_index[869] = '{7};
test_input[6960:6967] = '{32'hc23978bd, 32'hc2969217, 32'h42483b81, 32'h40897a03, 32'h42b4fa1e, 32'h4275e2c9, 32'hc2031371, 32'h3f200250};
test_output[870] = '{32'h42b4fa1e};
test_index[870] = '{4};
test_input[6968:6975] = '{32'h42ad9f74, 32'h42a45f62, 32'hc0c54eb2, 32'h416ce5b5, 32'h413b80b8, 32'h4134a029, 32'hc1408dc0, 32'hc2457206};
test_output[871] = '{32'h42ad9f74};
test_index[871] = '{0};
test_input[6976:6983] = '{32'h423aaf96, 32'hc290a5cc, 32'hc2aeb19e, 32'hc25c6f1f, 32'h4177c06d, 32'hc27dce4f, 32'hc24c81ad, 32'h420c89e8};
test_output[872] = '{32'h423aaf96};
test_index[872] = '{0};
test_input[6984:6991] = '{32'hc2c3572e, 32'hc26a4431, 32'hc2564c79, 32'h42a1550a, 32'hc2990d9a, 32'hc256e11d, 32'hc2067e62, 32'hc21ca963};
test_output[873] = '{32'h42a1550a};
test_index[873] = '{3};
test_input[6992:6999] = '{32'hc1a6d65a, 32'hc2bf7309, 32'h4262c425, 32'hc28e627c, 32'hc29caa01, 32'hc2b85397, 32'hc287416c, 32'hc21001e5};
test_output[874] = '{32'h4262c425};
test_index[874] = '{2};
test_input[7000:7007] = '{32'hbf85c21e, 32'h40c53325, 32'hc26e18c3, 32'h42053ad8, 32'hc10c4e64, 32'h418b6a5e, 32'hc1aa62c7, 32'h4259198f};
test_output[875] = '{32'h4259198f};
test_index[875] = '{7};
test_input[7008:7015] = '{32'hc01bf1dd, 32'hc241addf, 32'hc21cb6bc, 32'hc19ddc06, 32'hc197b6a2, 32'h41988665, 32'hc18182da, 32'hc25d0f84};
test_output[876] = '{32'h41988665};
test_index[876] = '{5};
test_input[7016:7023] = '{32'hc2322734, 32'hc297e8df, 32'hc09ea5fd, 32'hc2c4d37b, 32'h429b12b9, 32'h42b08386, 32'h41b53d28, 32'h42964af5};
test_output[877] = '{32'h42b08386};
test_index[877] = '{5};
test_input[7024:7031] = '{32'h3fb2116a, 32'h42a62ef1, 32'hc199a861, 32'h42873323, 32'hc296cbb8, 32'h41e29fae, 32'hc218a4a1, 32'h42a33c19};
test_output[878] = '{32'h42a62ef1};
test_index[878] = '{1};
test_input[7032:7039] = '{32'hc0b2781f, 32'hc16dacaf, 32'h429e2292, 32'hc27911c9, 32'h3f6a6514, 32'h42c723f4, 32'h40cb03d5, 32'h42a26058};
test_output[879] = '{32'h42c723f4};
test_index[879] = '{5};
test_input[7040:7047] = '{32'h42490d3d, 32'hc250f88a, 32'h42a7a754, 32'hc23ec705, 32'hc23dda81, 32'hc264a400, 32'hc27a474f, 32'hc275fdc5};
test_output[880] = '{32'h42a7a754};
test_index[880] = '{2};
test_input[7048:7055] = '{32'hc2014fd7, 32'hc21fbcd0, 32'h41a044e2, 32'hc21f2482, 32'h42a6f989, 32'hbe50943e, 32'h417d2f80, 32'h42b7f6f5};
test_output[881] = '{32'h42b7f6f5};
test_index[881] = '{7};
test_input[7056:7063] = '{32'h4204c2d4, 32'hc2a8e2b9, 32'hc20d178d, 32'hc29ba32e, 32'h42aecf05, 32'hc248bcab, 32'hc222c6ed, 32'h427e8088};
test_output[882] = '{32'h42aecf05};
test_index[882] = '{4};
test_input[7064:7071] = '{32'h4273e43a, 32'hc2ab5da3, 32'hc2bf0a73, 32'h41d33764, 32'hc2c6d6ed, 32'hc2bb5727, 32'hc200b285, 32'hc2904f04};
test_output[883] = '{32'h4273e43a};
test_index[883] = '{0};
test_input[7072:7079] = '{32'hc26a2f4d, 32'hc29ba3e1, 32'hc25419b4, 32'hc1f6d1df, 32'hc2315460, 32'h4219471d, 32'h423735bd, 32'hc1ee38c6};
test_output[884] = '{32'h423735bd};
test_index[884] = '{6};
test_input[7080:7087] = '{32'h42beb8c1, 32'hc0195340, 32'h41d2b095, 32'hc1fbf350, 32'h40d98036, 32'hc286319e, 32'hc23b527f, 32'h423db87c};
test_output[885] = '{32'h42beb8c1};
test_index[885] = '{0};
test_input[7088:7095] = '{32'hc27afe61, 32'h413f6db6, 32'hc200a3a6, 32'h421175f1, 32'h421e2bfd, 32'h4048c9c5, 32'h42701c0c, 32'hc124bcff};
test_output[886] = '{32'h42701c0c};
test_index[886] = '{6};
test_input[7096:7103] = '{32'hc28c711d, 32'h42bb76a4, 32'h429503a1, 32'h429988a0, 32'h4230416f, 32'h42740d20, 32'h4250a059, 32'h421c750e};
test_output[887] = '{32'h42bb76a4};
test_index[887] = '{1};
test_input[7104:7111] = '{32'h42acec39, 32'hc286024e, 32'h41673e62, 32'hc2949678, 32'hc15a61f6, 32'hc29a5e71, 32'hc20ed68c, 32'h409fd6f0};
test_output[888] = '{32'h42acec39};
test_index[888] = '{0};
test_input[7112:7119] = '{32'h4220c41d, 32'h4285c434, 32'h42253fb8, 32'h4245b287, 32'h3ea4111e, 32'h422068f5, 32'hc1ae9ce5, 32'hc2a17d6d};
test_output[889] = '{32'h4285c434};
test_index[889] = '{1};
test_input[7120:7127] = '{32'h426c28b4, 32'hc11f0deb, 32'h42198809, 32'hc2b9cce8, 32'h42b0443a, 32'h424039c5, 32'h42980322, 32'h42ae8c93};
test_output[890] = '{32'h42b0443a};
test_index[890] = '{4};
test_input[7128:7135] = '{32'hc2a45f4c, 32'hc252b3b0, 32'h41efa445, 32'hc2c675dc, 32'hc17a1b6d, 32'hc2c7550a, 32'h4267420b, 32'h41e738e4};
test_output[891] = '{32'h4267420b};
test_index[891] = '{6};
test_input[7136:7143] = '{32'hc2b37e22, 32'hc263df69, 32'h42a3ddfc, 32'h426da0dd, 32'hc28f327e, 32'hc26dca0c, 32'hc22a5197, 32'h429d331b};
test_output[892] = '{32'h42a3ddfc};
test_index[892] = '{2};
test_input[7144:7151] = '{32'h4224a3d8, 32'h425197bf, 32'hc254e75b, 32'h42a38b52, 32'hc2a65068, 32'hc28eee5e, 32'hc2b8fdc5, 32'h41a3d3b4};
test_output[893] = '{32'h42a38b52};
test_index[893] = '{3};
test_input[7152:7159] = '{32'h41d44c2f, 32'h42971755, 32'hc214e149, 32'hc1650e86, 32'hc07ce16b, 32'h42bddfad, 32'h415a0c7b, 32'hc2683f11};
test_output[894] = '{32'h42bddfad};
test_index[894] = '{5};
test_input[7160:7167] = '{32'hc220e429, 32'hc24a07ea, 32'hc29e488c, 32'h3f002d0e, 32'hc296bab8, 32'hc17a7dbd, 32'h411fd660, 32'h4260d9cd};
test_output[895] = '{32'h4260d9cd};
test_index[895] = '{7};
test_input[7168:7175] = '{32'hc2539e86, 32'h4096b12e, 32'hc291f4bc, 32'h414cf6bf, 32'h42a44c07, 32'hc28cb873, 32'h42277c4d, 32'hc287636f};
test_output[896] = '{32'h42a44c07};
test_index[896] = '{4};
test_input[7176:7183] = '{32'hc2016942, 32'h418fa42d, 32'h3fb68eab, 32'hc1a98f3e, 32'hc2095a85, 32'h4210f96b, 32'h42758321, 32'hbdf9e793};
test_output[897] = '{32'h42758321};
test_index[897] = '{6};
test_input[7184:7191] = '{32'hc1f2d415, 32'h429b5021, 32'h42b2eb20, 32'h421088b6, 32'h42b9de2a, 32'hc2912430, 32'h4251f820, 32'hc1702e6c};
test_output[898] = '{32'h42b9de2a};
test_index[898] = '{4};
test_input[7192:7199] = '{32'h429a2aae, 32'h42463f2c, 32'h42a8956f, 32'hc296e6de, 32'h428fbc12, 32'h428fb18d, 32'h4139c15a, 32'hc202cb57};
test_output[899] = '{32'h42a8956f};
test_index[899] = '{2};
test_input[7200:7207] = '{32'hc2b70a07, 32'h414eda81, 32'h429d4d56, 32'hc2afee3c, 32'hc2696ffd, 32'hc1a98f03, 32'hc1cfd47c, 32'hc2679290};
test_output[900] = '{32'h429d4d56};
test_index[900] = '{2};
test_input[7208:7215] = '{32'hc2801edc, 32'hc2a2d99f, 32'hc26b5bab, 32'hc2969904, 32'h423a88d0, 32'h426da613, 32'hc1892f32, 32'h42ab8cc4};
test_output[901] = '{32'h42ab8cc4};
test_index[901] = '{7};
test_input[7216:7223] = '{32'h42026e93, 32'hc1ee3798, 32'hc21cf654, 32'hc1e395c3, 32'h4220463d, 32'h41db2413, 32'h42aa8320, 32'hc1b7b3b2};
test_output[902] = '{32'h42aa8320};
test_index[902] = '{6};
test_input[7224:7231] = '{32'hc29dec0f, 32'h426be366, 32'h41d7a26b, 32'hc25d0147, 32'h4256aea1, 32'hc0c5224b, 32'hc2c203ed, 32'h42a7cf6c};
test_output[903] = '{32'h42a7cf6c};
test_index[903] = '{7};
test_input[7232:7239] = '{32'h42890ffa, 32'h410b42f0, 32'h427ec65d, 32'h4208c1fa, 32'hc28ea0d6, 32'h42b43082, 32'hc2c2ebed, 32'hc23578d7};
test_output[904] = '{32'h42b43082};
test_index[904] = '{5};
test_input[7240:7247] = '{32'hc11416a6, 32'hc2a0c6dc, 32'h425504ab, 32'hc2a7bec5, 32'hc2c1d307, 32'h427b25d4, 32'hc2162a95, 32'h428152f3};
test_output[905] = '{32'h428152f3};
test_index[905] = '{7};
test_input[7248:7255] = '{32'h428ec5ad, 32'hc2876628, 32'h41a8adc0, 32'hc2a8a350, 32'hc1663646, 32'h4162e881, 32'h4180880a, 32'h410263a5};
test_output[906] = '{32'h428ec5ad};
test_index[906] = '{0};
test_input[7256:7263] = '{32'hc185a042, 32'h418f617f, 32'h427ffbaf, 32'hc29c5149, 32'hc296eb70, 32'hc1f25a79, 32'h42c79d0d, 32'hc2908530};
test_output[907] = '{32'h42c79d0d};
test_index[907] = '{6};
test_input[7264:7271] = '{32'h42b54b65, 32'h429fdaee, 32'h4246b16d, 32'h42a00b67, 32'hc29b69f1, 32'h4235e0d0, 32'hc149f32d, 32'hc20b263d};
test_output[908] = '{32'h42b54b65};
test_index[908] = '{0};
test_input[7272:7279] = '{32'hc2674cce, 32'h42249b7f, 32'h42c20026, 32'h42681290, 32'h3ed601e6, 32'hc2b2a6d8, 32'h4263d1b8, 32'h42453d5e};
test_output[909] = '{32'h42c20026};
test_index[909] = '{2};
test_input[7280:7287] = '{32'h407aa112, 32'hc149814f, 32'hc265d4c6, 32'hbf388794, 32'h42b32fd1, 32'h41b58de2, 32'hc21e82cc, 32'h41c5c2e3};
test_output[910] = '{32'h42b32fd1};
test_index[910] = '{4};
test_input[7288:7295] = '{32'hc18f30fe, 32'hc25e6461, 32'h42abf4e3, 32'hc2a369a5, 32'h424d401f, 32'hc1fd006b, 32'hc2824c09, 32'hc22f96a5};
test_output[911] = '{32'h42abf4e3};
test_index[911] = '{2};
test_input[7296:7303] = '{32'h42c5deb7, 32'h42a6e7bc, 32'hc266a6b0, 32'h426bcd97, 32'h41265cb5, 32'hc1f620ad, 32'hc27d5ffe, 32'hc2926465};
test_output[912] = '{32'h42c5deb7};
test_index[912] = '{0};
test_input[7304:7311] = '{32'hc2bcbf00, 32'hc190cdd1, 32'hc2b6cbf6, 32'hc294c250, 32'hc281a73f, 32'h42ba7825, 32'h4292c28b, 32'hc1d700c3};
test_output[913] = '{32'h42ba7825};
test_index[913] = '{5};
test_input[7312:7319] = '{32'hc24e9e50, 32'h4272df08, 32'hc128cca2, 32'h42061b30, 32'h4292d3c3, 32'hc249c925, 32'h41ee33c7, 32'hc201aefe};
test_output[914] = '{32'h4292d3c3};
test_index[914] = '{4};
test_input[7320:7327] = '{32'hc29035dc, 32'hc2a842e9, 32'h42c0d1fd, 32'h42942f0d, 32'h404009e1, 32'h419d207b, 32'h40f90766, 32'hc1df0c9e};
test_output[915] = '{32'h42c0d1fd};
test_index[915] = '{2};
test_input[7328:7335] = '{32'hc25bbb08, 32'h42a47d0f, 32'hc23d5964, 32'h41785fb8, 32'h424b8988, 32'h4295cdc2, 32'hc11f6ba9, 32'h41586402};
test_output[916] = '{32'h42a47d0f};
test_index[916] = '{1};
test_input[7336:7343] = '{32'hc1702a92, 32'h42657999, 32'hc29b60b1, 32'hc2736a59, 32'h4297ad96, 32'hc293f0fa, 32'hc2be6d04, 32'h423e4601};
test_output[917] = '{32'h4297ad96};
test_index[917] = '{4};
test_input[7344:7351] = '{32'hc26e41ef, 32'hc203520c, 32'hc2a7adba, 32'hc238966a, 32'h41c758ad, 32'hc235bbb7, 32'h4122452a, 32'h414f80b8};
test_output[918] = '{32'h41c758ad};
test_index[918] = '{4};
test_input[7352:7359] = '{32'h41578bad, 32'hbf45bb16, 32'hc29d12f4, 32'hc19a614b, 32'h41cdbaba, 32'hc2a7abc6, 32'hc1b03905, 32'h4265c98e};
test_output[919] = '{32'h4265c98e};
test_index[919] = '{7};
test_input[7360:7367] = '{32'h42825434, 32'h419059fc, 32'h427b4153, 32'h4289cb2b, 32'h42567c99, 32'hc28c68c4, 32'hc1dbfd92, 32'h42829a04};
test_output[920] = '{32'h4289cb2b};
test_index[920] = '{3};
test_input[7368:7375] = '{32'hc236fe9a, 32'hc222617e, 32'hc29f66b3, 32'h427bad62, 32'h41ecd418, 32'h3e53dc34, 32'hc25837c5, 32'hc00616d6};
test_output[921] = '{32'h427bad62};
test_index[921] = '{3};
test_input[7376:7383] = '{32'hc24a0577, 32'h424c5fe4, 32'h4271dad0, 32'h4278ed48, 32'h42ac5729, 32'hc166c6e5, 32'hc1cbf6fb, 32'h413af8f7};
test_output[922] = '{32'h42ac5729};
test_index[922] = '{4};
test_input[7384:7391] = '{32'h4119b498, 32'h424835fa, 32'h42a22c63, 32'h4264c05b, 32'hc26f7be3, 32'hc1ca68a1, 32'h4290cade, 32'hc2a760f4};
test_output[923] = '{32'h42a22c63};
test_index[923] = '{2};
test_input[7392:7399] = '{32'h411d7b22, 32'h423459b7, 32'hc2143657, 32'hc1f2a42b, 32'hc29a171e, 32'h429880e4, 32'h41172da3, 32'h424c9bc9};
test_output[924] = '{32'h429880e4};
test_index[924] = '{5};
test_input[7400:7407] = '{32'hc1f622f4, 32'h412cc936, 32'hc24aeea5, 32'hc28061a4, 32'h4200357d, 32'h41ad1b22, 32'h42742721, 32'hc25e5428};
test_output[925] = '{32'h42742721};
test_index[925] = '{6};
test_input[7408:7415] = '{32'h42736eef, 32'hc2663e49, 32'hc201462a, 32'hc208476f, 32'hc1a81796, 32'h42aff86b, 32'hc288430e, 32'h4250bc24};
test_output[926] = '{32'h42aff86b};
test_index[926] = '{5};
test_input[7416:7423] = '{32'h426e0f43, 32'h427072ee, 32'hc2928768, 32'h41d958b9, 32'hc2a3c1b8, 32'hc293c61c, 32'h428e4181, 32'h42189c7a};
test_output[927] = '{32'h428e4181};
test_index[927] = '{6};
test_input[7424:7431] = '{32'hc2c2e839, 32'h418329b9, 32'h425b2702, 32'hc2697128, 32'hc2b82fa0, 32'h418f77ce, 32'h4293b08a, 32'h42a7a6db};
test_output[928] = '{32'h42a7a6db};
test_index[928] = '{7};
test_input[7432:7439] = '{32'hc1e93485, 32'hc289ed9c, 32'hc245ccdc, 32'h42b16ed1, 32'h402e73c2, 32'h42824d9c, 32'hc2599b24, 32'hc1b80550};
test_output[929] = '{32'h42b16ed1};
test_index[929] = '{3};
test_input[7440:7447] = '{32'h407ad7f7, 32'h4282026c, 32'h42b752e7, 32'hc0cdcd5b, 32'h41d81157, 32'hc1e63892, 32'h4121eecf, 32'hc1abe1a9};
test_output[930] = '{32'h42b752e7};
test_index[930] = '{2};
test_input[7448:7455] = '{32'h42475c38, 32'hc2816d46, 32'h41625c08, 32'hc14a7acf, 32'h4112c52f, 32'h4291d2c4, 32'h41776992, 32'h422b8882};
test_output[931] = '{32'h4291d2c4};
test_index[931] = '{5};
test_input[7456:7463] = '{32'hc2b62d2a, 32'h42691e46, 32'h42adf3a6, 32'hc211b5bb, 32'hc224b610, 32'h420cc18c, 32'h421eb7c5, 32'hc272b4db};
test_output[932] = '{32'h42adf3a6};
test_index[932] = '{2};
test_input[7464:7471] = '{32'hc008c873, 32'h42baf97f, 32'h420b4db8, 32'h41a89ca8, 32'hc256d1ca, 32'hc1dd27cc, 32'hc0098d94, 32'hc25aa2fc};
test_output[933] = '{32'h42baf97f};
test_index[933] = '{1};
test_input[7472:7479] = '{32'h4215a97b, 32'hc2b4e804, 32'hc2ac6e52, 32'hc1b88f86, 32'h4098b914, 32'h41c12a9d, 32'h3fb512c5, 32'h420876f2};
test_output[934] = '{32'h4215a97b};
test_index[934] = '{0};
test_input[7480:7487] = '{32'h42231371, 32'h41e1f58f, 32'h42bc742b, 32'hc2a1508b, 32'hc2b2cf42, 32'hc29098a6, 32'h42bd0b8c, 32'h42ae87ec};
test_output[935] = '{32'h42bd0b8c};
test_index[935] = '{6};
test_input[7488:7495] = '{32'hc2973f4b, 32'h419ef153, 32'hc2c00729, 32'h416d1997, 32'hbf898db5, 32'h41eb251c, 32'h42a696a0, 32'hc264878b};
test_output[936] = '{32'h42a696a0};
test_index[936] = '{6};
test_input[7496:7503] = '{32'hc2393fd7, 32'h4234cce0, 32'hc286a622, 32'h429a06e4, 32'h421a5a7c, 32'hc2a71f83, 32'h413978e2, 32'hc21a3547};
test_output[937] = '{32'h429a06e4};
test_index[937] = '{3};
test_input[7504:7511] = '{32'hc1629b09, 32'hc1f591bb, 32'hc1d4e3dc, 32'h422004ee, 32'h42bfc6f0, 32'h429d363e, 32'hc177dea5, 32'h427f69e5};
test_output[938] = '{32'h42bfc6f0};
test_index[938] = '{4};
test_input[7512:7519] = '{32'h41c78ac5, 32'h424c4b5d, 32'h410f0168, 32'h42a007b8, 32'h4187aeee, 32'hc1f0bb18, 32'hc26bdaac, 32'hc23dc2cb};
test_output[939] = '{32'h42a007b8};
test_index[939] = '{3};
test_input[7520:7527] = '{32'hc28b728e, 32'hc1626beb, 32'h418a4b70, 32'h400f83da, 32'h422d8d18, 32'h42975b65, 32'hc2a6db6d, 32'hc254e791};
test_output[940] = '{32'h42975b65};
test_index[940] = '{5};
test_input[7528:7535] = '{32'hc2427d3f, 32'h4293d616, 32'hc2390e95, 32'h426f6991, 32'hc0b55cad, 32'hc1839dce, 32'hc237e3f1, 32'hc2a31011};
test_output[941] = '{32'h4293d616};
test_index[941] = '{1};
test_input[7536:7543] = '{32'hc2990bf8, 32'hc2973fa3, 32'h42a89474, 32'h428d51b1, 32'h42219183, 32'h3f95b03e, 32'h41e35376, 32'h42855dc2};
test_output[942] = '{32'h42a89474};
test_index[942] = '{2};
test_input[7544:7551] = '{32'h42ba5a08, 32'h42c13263, 32'hc29d7400, 32'hc199a032, 32'hc2ba9659, 32'hc1e6afc8, 32'hc2b0bb29, 32'hc0bf097f};
test_output[943] = '{32'h42c13263};
test_index[943] = '{1};
test_input[7552:7559] = '{32'hc1cc57a7, 32'hc29bb4bb, 32'hc2015e6b, 32'h41141bf1, 32'h41a15570, 32'hc1007da5, 32'h4245b521, 32'hc2aa8e6b};
test_output[944] = '{32'h4245b521};
test_index[944] = '{6};
test_input[7560:7567] = '{32'hc1b76ce6, 32'hc29937ce, 32'hc1f4777d, 32'h4236d215, 32'h41277b0e, 32'h41ce550c, 32'h429744a1, 32'h421bd244};
test_output[945] = '{32'h429744a1};
test_index[945] = '{6};
test_input[7568:7575] = '{32'h428fa866, 32'hc0ae0533, 32'hc22e7a8a, 32'h42bc8d69, 32'h416e1e16, 32'h42af42a6, 32'h4253e916, 32'hc2808053};
test_output[946] = '{32'h42bc8d69};
test_index[946] = '{3};
test_input[7576:7583] = '{32'h42974f33, 32'hc1877bb7, 32'hc1dd79bf, 32'h42ade3b5, 32'hc20c8b70, 32'h41d126c4, 32'h40f4939b, 32'h420ae9a8};
test_output[947] = '{32'h42ade3b5};
test_index[947] = '{3};
test_input[7584:7591] = '{32'hc149456f, 32'h41e08491, 32'hc2b21efd, 32'h42bbc075, 32'h4291b5f4, 32'hc2c218d2, 32'hc2aba3ce, 32'hc20110c9};
test_output[948] = '{32'h42bbc075};
test_index[948] = '{3};
test_input[7592:7599] = '{32'hc2b62569, 32'h427b48bb, 32'h4138c2bb, 32'h40d24aa7, 32'h42a087eb, 32'hc2b1eaa1, 32'h42408ca8, 32'h42bc7d6f};
test_output[949] = '{32'h42bc7d6f};
test_index[949] = '{7};
test_input[7600:7607] = '{32'hc24caf03, 32'h42606bbb, 32'h42694bb1, 32'h42bd0dff, 32'h423ba96f, 32'hc2a399cc, 32'hc1aad433, 32'hc2367668};
test_output[950] = '{32'h42bd0dff};
test_index[950] = '{3};
test_input[7608:7615] = '{32'hc2c1b17f, 32'h429d2ce5, 32'hc2b954f5, 32'h410725b2, 32'hc1f5a794, 32'hc0f6735a, 32'hc240d6ac, 32'h41921cc0};
test_output[951] = '{32'h429d2ce5};
test_index[951] = '{1};
test_input[7616:7623] = '{32'h4283218b, 32'hc2a5d963, 32'h42b783fe, 32'hc1079224, 32'hc2c6d37e, 32'h42853578, 32'h425c86ae, 32'hc2466cf4};
test_output[952] = '{32'h42b783fe};
test_index[952] = '{2};
test_input[7624:7631] = '{32'h426ad11d, 32'h42897fd6, 32'hc1bcc233, 32'h4261d9aa, 32'h420ee69a, 32'h40b54d8a, 32'h4210cd32, 32'hc27ad800};
test_output[953] = '{32'h42897fd6};
test_index[953] = '{1};
test_input[7632:7639] = '{32'h41b74277, 32'h42335d70, 32'hc2b97ef7, 32'hc2702b96, 32'hc289eb76, 32'hc25d6e90, 32'hc2aabd2a, 32'h425ef448};
test_output[954] = '{32'h425ef448};
test_index[954] = '{7};
test_input[7640:7647] = '{32'h41dc15f2, 32'h4207026c, 32'h418efccb, 32'hc2883719, 32'hc2b94555, 32'hc2ac7a8a, 32'hc29fb8f3, 32'hc18e9ddd};
test_output[955] = '{32'h4207026c};
test_index[955] = '{1};
test_input[7648:7655] = '{32'h41668875, 32'hc2b07300, 32'h4195d56f, 32'h427da89b, 32'h427a85c6, 32'hc2becd87, 32'hbfc2bb5b, 32'hc177e3bc};
test_output[956] = '{32'h427da89b};
test_index[956] = '{3};
test_input[7656:7663] = '{32'h42ad5c00, 32'h42b37ee5, 32'h40a95cc2, 32'hc1acd2f7, 32'hc1747830, 32'hc2630913, 32'hc29e7fa4, 32'hc0734e05};
test_output[957] = '{32'h42b37ee5};
test_index[957] = '{1};
test_input[7664:7671] = '{32'h41bb1634, 32'h4286e599, 32'hc26fb670, 32'hc282e527, 32'hc2c0580a, 32'hc2c1777f, 32'hc24bdd75, 32'h42318638};
test_output[958] = '{32'h4286e599};
test_index[958] = '{1};
test_input[7672:7679] = '{32'h42a4db90, 32'h41aae4e8, 32'h42b59e90, 32'h42c0b59b, 32'hc2b871b8, 32'h41eae3a9, 32'hc28b5c08, 32'hc29254d1};
test_output[959] = '{32'h42c0b59b};
test_index[959] = '{3};
test_input[7680:7687] = '{32'hc20f5452, 32'hc293f935, 32'h428aa9c0, 32'h4122664b, 32'h422513cc, 32'h42685976, 32'h420fe087, 32'hc2a8c5ed};
test_output[960] = '{32'h428aa9c0};
test_index[960] = '{2};
test_input[7688:7695] = '{32'hbf0b00d3, 32'hc2a5f1b5, 32'hc1b08b70, 32'hc28be61e, 32'hc2ba0313, 32'h41fde217, 32'hc1823ee0, 32'h4211840b};
test_output[961] = '{32'h4211840b};
test_index[961] = '{7};
test_input[7696:7703] = '{32'hc2936e7a, 32'h42009b32, 32'hc26d3104, 32'h425ca8a1, 32'h42b7c03e, 32'hc12907bc, 32'h421c16c0, 32'hc23cecda};
test_output[962] = '{32'h42b7c03e};
test_index[962] = '{4};
test_input[7704:7711] = '{32'hc29f409c, 32'hc2ac2a37, 32'hc2afe2d5, 32'h42a754fa, 32'h41e970ca, 32'h4144d2e3, 32'hc08d538d, 32'h42ac3150};
test_output[963] = '{32'h42ac3150};
test_index[963] = '{7};
test_input[7712:7719] = '{32'hc29d9a54, 32'h42a6ba8a, 32'h42b88884, 32'hc2b81632, 32'h423ccc27, 32'h41d2d9df, 32'h418a6aee, 32'h42a86991};
test_output[964] = '{32'h42b88884};
test_index[964] = '{2};
test_input[7720:7727] = '{32'h421cc9d2, 32'hc2969b84, 32'hc240ebc3, 32'hc2b16ff9, 32'h428e7b01, 32'h42451860, 32'hc1095326, 32'hc2067239};
test_output[965] = '{32'h428e7b01};
test_index[965] = '{4};
test_input[7728:7735] = '{32'h42259ce6, 32'hc2a753bc, 32'h42242e59, 32'h42b3cea4, 32'h428fa857, 32'h42321173, 32'hc2b56a12, 32'h40eb8ad2};
test_output[966] = '{32'h42b3cea4};
test_index[966] = '{3};
test_input[7736:7743] = '{32'hc292ea2f, 32'h3fbbfea6, 32'h42156a75, 32'hc28fa043, 32'hc268b631, 32'h4290f2f0, 32'h4289a86e, 32'hc1230fde};
test_output[967] = '{32'h4290f2f0};
test_index[967] = '{5};
test_input[7744:7751] = '{32'h41ace316, 32'h42418a9d, 32'hc29efc63, 32'h419f63ff, 32'hc291802d, 32'h42c2979f, 32'h4200dc72, 32'h42a493ae};
test_output[968] = '{32'h42c2979f};
test_index[968] = '{5};
test_input[7752:7759] = '{32'hc2bf24d4, 32'hc2b7025f, 32'h41b418af, 32'hc2a204d8, 32'hc20a9548, 32'h42960d1c, 32'h42887cbf, 32'hc1d7c613};
test_output[969] = '{32'h42960d1c};
test_index[969] = '{5};
test_input[7760:7767] = '{32'h42c3f7e2, 32'h428d406c, 32'h41a3ec69, 32'hc226d7f6, 32'h42c1076c, 32'h410fdbe1, 32'h4114cb35, 32'h42040191};
test_output[970] = '{32'h42c3f7e2};
test_index[970] = '{0};
test_input[7768:7775] = '{32'hc1bb1aca, 32'h423bd5dd, 32'hc2319318, 32'hc2179e46, 32'hc17287a1, 32'h423b1b57, 32'hc215f890, 32'h42b40802};
test_output[971] = '{32'h42b40802};
test_index[971] = '{7};
test_input[7776:7783] = '{32'hc23ad07f, 32'h40ae699d, 32'h425e13bb, 32'h42b51640, 32'hc1aa6a6e, 32'hc25329e7, 32'h42ab20aa, 32'h424ea65f};
test_output[972] = '{32'h42b51640};
test_index[972] = '{3};
test_input[7784:7791] = '{32'hc21277ab, 32'hc2514026, 32'h414031d2, 32'h42af6d2b, 32'hc2a35309, 32'h4161e448, 32'h42846a89, 32'h4167f90c};
test_output[973] = '{32'h42af6d2b};
test_index[973] = '{3};
test_input[7792:7799] = '{32'h40aff509, 32'h425b59ab, 32'hc2c61327, 32'h42b6874e, 32'h429d3f06, 32'h4283d942, 32'hc18c16c3, 32'h4280854d};
test_output[974] = '{32'h42b6874e};
test_index[974] = '{3};
test_input[7800:7807] = '{32'h4292a0d5, 32'hc2aca706, 32'hc1e762ab, 32'hc2b85238, 32'h41aa9d98, 32'hc2216783, 32'h4283b732, 32'h42548ccf};
test_output[975] = '{32'h4292a0d5};
test_index[975] = '{0};
test_input[7808:7815] = '{32'hc29701d4, 32'hc1ea817a, 32'h42827666, 32'hc28fdbbb, 32'h41ed20b1, 32'h42a110c1, 32'h4142960e, 32'h408195a6};
test_output[976] = '{32'h42a110c1};
test_index[976] = '{5};
test_input[7816:7823] = '{32'hc24c80b0, 32'h418b889c, 32'h42a51564, 32'hc273e1ea, 32'hc194be45, 32'hc2bce9ee, 32'hc2ab936b, 32'hc13d1799};
test_output[977] = '{32'h42a51564};
test_index[977] = '{2};
test_input[7824:7831] = '{32'hc235b2ff, 32'h42c20ae5, 32'h42c390a5, 32'hc24f3011, 32'hc116dd06, 32'hc228fc5c, 32'h417032fb, 32'hc21d78e4};
test_output[978] = '{32'h42c390a5};
test_index[978] = '{2};
test_input[7832:7839] = '{32'h429b82d9, 32'hc2a0e0c4, 32'h42adb416, 32'h4282d32c, 32'h42bb08e7, 32'h428761b1, 32'hc29f14d7, 32'hc261062f};
test_output[979] = '{32'h42bb08e7};
test_index[979] = '{4};
test_input[7840:7847] = '{32'h4273b063, 32'h4225562c, 32'hc2bfc95b, 32'h42bf3fa1, 32'h419a64e4, 32'hc2ad2526, 32'h42c514e2, 32'hbfe532cf};
test_output[980] = '{32'h42c514e2};
test_index[980] = '{6};
test_input[7848:7855] = '{32'h42a49809, 32'h3ca74c0a, 32'hbf10051d, 32'hc1cd71cd, 32'h429ddf2a, 32'hc21dd855, 32'h42b13a39, 32'h420aab31};
test_output[981] = '{32'h42b13a39};
test_index[981] = '{6};
test_input[7856:7863] = '{32'h401cb427, 32'h42b44bcb, 32'h3e1faa5f, 32'h4140a57f, 32'h42a5f84e, 32'hc18ad44f, 32'h4291df61, 32'hc21c4e6c};
test_output[982] = '{32'h42b44bcb};
test_index[982] = '{1};
test_input[7864:7871] = '{32'h429b6664, 32'hc19101fe, 32'hc1e63990, 32'h42bfa490, 32'h42b1c171, 32'hbbb2f705, 32'hc2c59a57, 32'h425e39c6};
test_output[983] = '{32'h42bfa490};
test_index[983] = '{3};
test_input[7872:7879] = '{32'hc14d1bdc, 32'h3fba6a4a, 32'hc2944123, 32'h42145be8, 32'h417bc79a, 32'hc226c153, 32'h41f89086, 32'hc240a50c};
test_output[984] = '{32'h42145be8};
test_index[984] = '{3};
test_input[7880:7887] = '{32'hc1ef5cd8, 32'hc2a836f1, 32'hc194eddb, 32'h41f1c37b, 32'hc29b203a, 32'hc18e052d, 32'h4285ac8d, 32'hc2a90893};
test_output[985] = '{32'h4285ac8d};
test_index[985] = '{6};
test_input[7888:7895] = '{32'h42bcd8b2, 32'hc22be826, 32'hc181b3d9, 32'h4242b755, 32'hc1156b03, 32'hc29b9c60, 32'h42ad924d, 32'hc060c282};
test_output[986] = '{32'h42bcd8b2};
test_index[986] = '{0};
test_input[7896:7903] = '{32'h4256cff9, 32'hc28477f3, 32'h4239a76b, 32'hc2c7808b, 32'h41e07cbd, 32'h429c67d3, 32'h416a1451, 32'hc26c9e4d};
test_output[987] = '{32'h429c67d3};
test_index[987] = '{5};
test_input[7904:7911] = '{32'hc1678b54, 32'h4077ee8d, 32'h429958c3, 32'h42544ff5, 32'h4221ccde, 32'h428387ce, 32'hc2873e2b, 32'hc296141d};
test_output[988] = '{32'h429958c3};
test_index[988] = '{2};
test_input[7912:7919] = '{32'h42c5b466, 32'hc2a42d32, 32'hc1d05e4b, 32'hc20ac735, 32'hc2077d3a, 32'h429346c7, 32'h4270007c, 32'hc16e5389};
test_output[989] = '{32'h42c5b466};
test_index[989] = '{0};
test_input[7920:7927] = '{32'hc2adb4f8, 32'h42aa9b8a, 32'hc236b829, 32'h41948eab, 32'h413da365, 32'h40f5e905, 32'hc20ef1c8, 32'h420b9628};
test_output[990] = '{32'h42aa9b8a};
test_index[990] = '{1};
test_input[7928:7935] = '{32'hc19c2d7e, 32'hc258ba9a, 32'h421d57f7, 32'hc27b8233, 32'h42a18cfc, 32'h411995e4, 32'hc28dc227, 32'h418f4955};
test_output[991] = '{32'h42a18cfc};
test_index[991] = '{4};
test_input[7936:7943] = '{32'h424b50da, 32'hc1e24a1a, 32'h42ad7bf8, 32'hc2b9afcf, 32'h412c43d3, 32'hc22b21b8, 32'h42368059, 32'hc2c1e4b4};
test_output[992] = '{32'h42ad7bf8};
test_index[992] = '{2};
test_input[7944:7951] = '{32'hc2a4aa86, 32'h41ee2e7f, 32'h42bf7351, 32'h42b22517, 32'hc2c17a61, 32'hc1c60cad, 32'hc1ee4f32, 32'h42219a4e};
test_output[993] = '{32'h42bf7351};
test_index[993] = '{2};
test_input[7952:7959] = '{32'h424e8f63, 32'hc2b4ded6, 32'h429413b3, 32'h424db02e, 32'h421731f6, 32'h42bb782b, 32'hc203b5a2, 32'hc255445c};
test_output[994] = '{32'h42bb782b};
test_index[994] = '{5};
test_input[7960:7967] = '{32'h42a08d6c, 32'h42862956, 32'hc22fb5b9, 32'h41a71eb4, 32'hc2beb097, 32'hc2b575eb, 32'hc2a94311, 32'h41831c74};
test_output[995] = '{32'h42a08d6c};
test_index[995] = '{0};
test_input[7968:7975] = '{32'h40eed4f4, 32'h41e678cd, 32'hc2b23fe3, 32'h42a1e73d, 32'hc2810649, 32'hc2c1e0a2, 32'h42c138db, 32'hc29b9002};
test_output[996] = '{32'h42c138db};
test_index[996] = '{6};
test_input[7976:7983] = '{32'h4124e231, 32'h41c2eeca, 32'hc16e8b51, 32'hc2128f50, 32'h40ce28f0, 32'hc2aab9fb, 32'h41961525, 32'h4201e2c7};
test_output[997] = '{32'h4201e2c7};
test_index[997] = '{7};
test_input[7984:7991] = '{32'h4259faba, 32'h411e8496, 32'h42995c2d, 32'h41f297b4, 32'h42a91dba, 32'h4298fbaf, 32'hc28e8da2, 32'hc186da15};
test_output[998] = '{32'h42a91dba};
test_index[998] = '{4};
test_input[7992:7999] = '{32'h4170694a, 32'hc260f756, 32'h41e11403, 32'h4110f3c4, 32'h42900e89, 32'h40d7dc07, 32'h4299d37e, 32'hc2c6834e};
test_output[999] = '{32'h4299d37e};
test_index[999] = '{6};
test_input[8000:8007] = '{32'h4172b15f, 32'hc2472f34, 32'hc1c1052d, 32'hc1aa0241, 32'hc11f150f, 32'hc22a8a8c, 32'hc28e4fac, 32'hc23ae256};
test_output[1000] = '{32'h4172b15f};
test_index[1000] = '{0};
test_input[8008:8015] = '{32'hc2b3a150, 32'hc247e299, 32'h42abd221, 32'hc25c293b, 32'hc2826b85, 32'hc2a244c8, 32'hc2914b9c, 32'h414adfed};
test_output[1001] = '{32'h42abd221};
test_index[1001] = '{2};
test_input[8016:8023] = '{32'hc29a4d47, 32'hc231d3bb, 32'hc2c2ddbc, 32'hc2020cee, 32'h4284a7a7, 32'h42b4fbd4, 32'h408f719f, 32'hc13017f9};
test_output[1002] = '{32'h42b4fbd4};
test_index[1002] = '{5};
test_input[8024:8031] = '{32'h418f37b1, 32'h42c7a1d5, 32'hc2ba8581, 32'h422f776e, 32'hc267e659, 32'hc2778b2f, 32'hc25df5e4, 32'hc206f124};
test_output[1003] = '{32'h42c7a1d5};
test_index[1003] = '{1};
test_input[8032:8039] = '{32'hc11b51f9, 32'h41a3f98a, 32'h421206ed, 32'h42bfd677, 32'hc1861161, 32'h427476e3, 32'h425619c4, 32'h42b0ad45};
test_output[1004] = '{32'h42bfd677};
test_index[1004] = '{3};
test_input[8040:8047] = '{32'hc2ab1de4, 32'hc2aafc1d, 32'hc2075717, 32'h42865b5b, 32'hc2b0d1f8, 32'hc288e755, 32'h4215db06, 32'h41c3328f};
test_output[1005] = '{32'h42865b5b};
test_index[1005] = '{3};
test_input[8048:8055] = '{32'h427d00b3, 32'h4284363a, 32'h429d762c, 32'hc22afdf7, 32'h42897d91, 32'hc280a4ed, 32'hc2195d06, 32'h42464c2d};
test_output[1006] = '{32'h429d762c};
test_index[1006] = '{2};
test_input[8056:8063] = '{32'h40a6c9d3, 32'hc10b13ad, 32'hc2b2a91d, 32'hc02aa410, 32'hc2197a39, 32'hc198d7f3, 32'hc219aabb, 32'h423a5425};
test_output[1007] = '{32'h423a5425};
test_index[1007] = '{7};
test_input[8064:8071] = '{32'hc0a99ad8, 32'h42c48c30, 32'hc2a25f3b, 32'hc1ceb3ae, 32'h414ccb6a, 32'h42b4f0c7, 32'h41ffe910, 32'h42b91fe0};
test_output[1008] = '{32'h42c48c30};
test_index[1008] = '{1};
test_input[8072:8079] = '{32'hc25a41e2, 32'hc22fd67e, 32'hc2015ce1, 32'h42a9e474, 32'h420827a8, 32'h4259848b, 32'hc1a58414, 32'hc1fcdaf1};
test_output[1009] = '{32'h42a9e474};
test_index[1009] = '{3};
test_input[8080:8087] = '{32'h41e3862e, 32'h4263c9b1, 32'hc28221f5, 32'hc244677c, 32'h429b093b, 32'h42b7feca, 32'h4282ea05, 32'hc29376fe};
test_output[1010] = '{32'h42b7feca};
test_index[1010] = '{5};
test_input[8088:8095] = '{32'h3e0e3a79, 32'h3f9fd857, 32'hc2bd02be, 32'hc2a8a76f, 32'h418c925f, 32'h40c34925, 32'h4194ab8a, 32'hc07fbcd0};
test_output[1011] = '{32'h4194ab8a};
test_index[1011] = '{6};
test_input[8096:8103] = '{32'h42a4297a, 32'h41f7d301, 32'h42b90089, 32'h429739c0, 32'hc21cfc26, 32'hc0dede36, 32'h4135e3a0, 32'hc1167b7f};
test_output[1012] = '{32'h42b90089};
test_index[1012] = '{2};
test_input[8104:8111] = '{32'hc0dc9521, 32'h41df6df1, 32'h428c83b2, 32'hc1365f3a, 32'hc2c18c21, 32'hc2ba5652, 32'hc20b10c6, 32'h4074d174};
test_output[1013] = '{32'h428c83b2};
test_index[1013] = '{2};
test_input[8112:8119] = '{32'h42170238, 32'hc159b205, 32'h428b50a1, 32'h4141c922, 32'hc279397d, 32'hc11355f2, 32'hc2402316, 32'hc1252dc3};
test_output[1014] = '{32'h428b50a1};
test_index[1014] = '{2};
test_input[8120:8127] = '{32'hc0bf64c8, 32'hc275e2b9, 32'h3d18c914, 32'hc28c0262, 32'h41a3b76f, 32'hc28d37fc, 32'h413573e4, 32'h41fd273d};
test_output[1015] = '{32'h41fd273d};
test_index[1015] = '{7};
test_input[8128:8135] = '{32'h42a210f7, 32'hc11de228, 32'h41fbb03c, 32'h42263d87, 32'hc26bdc87, 32'h415d19e9, 32'h4286aeb6, 32'h426c4c23};
test_output[1016] = '{32'h42a210f7};
test_index[1016] = '{0};
test_input[8136:8143] = '{32'hc1f4d215, 32'h42a82560, 32'hc2602fb6, 32'h408f90e2, 32'h4294f8ce, 32'h42806258, 32'hc28c110e, 32'h41c296fb};
test_output[1017] = '{32'h42a82560};
test_index[1017] = '{1};
test_input[8144:8151] = '{32'hc27df77b, 32'h4261807e, 32'hc10d0254, 32'hc244082c, 32'hc1f9020c, 32'hc2c0be4d, 32'hc1b896ca, 32'h4284068c};
test_output[1018] = '{32'h4284068c};
test_index[1018] = '{7};
test_input[8152:8159] = '{32'hc25b8f61, 32'hc275a3ed, 32'hc2921e69, 32'hc2449816, 32'hc28d3288, 32'hc1458bce, 32'hc12da407, 32'hc2ae2c06};
test_output[1019] = '{32'hc12da407};
test_index[1019] = '{6};
test_input[8160:8167] = '{32'hc28c428b, 32'h42994487, 32'hc06fbee9, 32'hc20f040c, 32'h42a3806d, 32'h425d8473, 32'h41886c37, 32'hc2193080};
test_output[1020] = '{32'h42a3806d};
test_index[1020] = '{4};
test_input[8168:8175] = '{32'hc1904035, 32'hc1e188e6, 32'h42c57ca1, 32'h4152b59d, 32'h41588fdf, 32'h42a7129b, 32'hc2769fbb, 32'hc216dcfd};
test_output[1021] = '{32'h42c57ca1};
test_index[1021] = '{2};
test_input[8176:8183] = '{32'h423ce37e, 32'hc21df242, 32'hc231ec67, 32'h4281cdb0, 32'h424ee7e3, 32'hc2b57894, 32'hc28ac156, 32'hc143f281};
test_output[1022] = '{32'h4281cdb0};
test_index[1022] = '{3};
test_input[8184:8191] = '{32'hc2a57772, 32'hc21110c6, 32'hc2077cea, 32'hc287340b, 32'hc1f95cb7, 32'hc1b65fc4, 32'h429a7a1c, 32'hc0b40053};
test_output[1023] = '{32'h429a7a1c};
test_index[1023] = '{6};
test_input[8192:8199] = '{32'h4286270b, 32'h42c143ce, 32'hc28d631c, 32'hc2b9efa4, 32'hc2836606, 32'h412afc92, 32'hc2465b9b, 32'hc0f34bd9};
test_output[1024] = '{32'h42c143ce};
test_index[1024] = '{1};
test_input[8200:8207] = '{32'h429877bd, 32'h4285ec77, 32'h4104efac, 32'h42a9545a, 32'hc2b667b9, 32'h429d5c9e, 32'h41afa11b, 32'hc117b4b8};
test_output[1025] = '{32'h42a9545a};
test_index[1025] = '{3};
test_input[8208:8215] = '{32'h426a5175, 32'hc27eac6f, 32'hc0eb6b93, 32'hc2a5f620, 32'hc29ef934, 32'h42c1b292, 32'h40a190fc, 32'hc209de35};
test_output[1026] = '{32'h42c1b292};
test_index[1026] = '{5};
test_input[8216:8223] = '{32'hc21df04a, 32'h42652b70, 32'h42655987, 32'h4154d553, 32'hc25cfd65, 32'h4130eb47, 32'h4288b31b, 32'h40e87380};
test_output[1027] = '{32'h4288b31b};
test_index[1027] = '{6};
test_input[8224:8231] = '{32'h42826d1a, 32'h4227e991, 32'h4254a6d9, 32'h426ebf02, 32'h428f1df5, 32'h42907dd0, 32'hc24dfd5f, 32'h42917023};
test_output[1028] = '{32'h42917023};
test_index[1028] = '{7};
test_input[8232:8239] = '{32'hc284ddcd, 32'h4212d3b1, 32'h42104a25, 32'h4135b8dc, 32'h4262503d, 32'hc20d43dd, 32'h4277b680, 32'h429d3586};
test_output[1029] = '{32'h429d3586};
test_index[1029] = '{7};
test_input[8240:8247] = '{32'hc21a38d9, 32'hc23f0f6a, 32'h42808d9d, 32'hc229acd1, 32'hc2029555, 32'hc1a978b2, 32'h424a800b, 32'hc21b7afc};
test_output[1030] = '{32'h42808d9d};
test_index[1030] = '{2};
test_input[8248:8255] = '{32'h41d1c70f, 32'h4264d246, 32'hc26c9ab2, 32'h41911a1c, 32'h4271dafb, 32'hc1f0e58e, 32'h41ba8c5b, 32'h41bcbfb1};
test_output[1031] = '{32'h4271dafb};
test_index[1031] = '{4};
test_input[8256:8263] = '{32'h42afc210, 32'hc159b993, 32'hc2525795, 32'hc2a4d1af, 32'h409f278d, 32'h425da0fd, 32'h417ceac0, 32'h41d58b7d};
test_output[1032] = '{32'h42afc210};
test_index[1032] = '{0};
test_input[8264:8271] = '{32'h42bc7b6c, 32'hc267ec54, 32'hc2b846e9, 32'hc23285b3, 32'hc1c4f3a3, 32'hc1eec8b9, 32'h42ae349d, 32'hc24eaeae};
test_output[1033] = '{32'h42bc7b6c};
test_index[1033] = '{0};
test_input[8272:8279] = '{32'h428533db, 32'hc2aa167c, 32'h42a53361, 32'h429189d8, 32'hc29e016d, 32'hc2b08799, 32'h4109472e, 32'h408da501};
test_output[1034] = '{32'h42a53361};
test_index[1034] = '{2};
test_input[8280:8287] = '{32'h4267d9b9, 32'hc1c5e698, 32'h42a23bd6, 32'h4246722c, 32'hc21e44bf, 32'h4201bf53, 32'h411b4532, 32'h41fdf673};
test_output[1035] = '{32'h42a23bd6};
test_index[1035] = '{2};
test_input[8288:8295] = '{32'hc1385dc7, 32'hc2ad19ba, 32'h41b054c0, 32'h42a503d9, 32'h41df6a7b, 32'hc27b7a81, 32'hc1f5a3ac, 32'hc2924d59};
test_output[1036] = '{32'h42a503d9};
test_index[1036] = '{3};
test_input[8296:8303] = '{32'h42708ace, 32'hc2915938, 32'h42c1e17a, 32'h4294a606, 32'hc29e7714, 32'hc1661cbe, 32'h42c09b59, 32'h42c1bd0b};
test_output[1037] = '{32'h42c1e17a};
test_index[1037] = '{2};
test_input[8304:8311] = '{32'hc212d086, 32'h422e4b72, 32'hc21f0285, 32'h42b024f0, 32'hc20ad9ca, 32'h427317cc, 32'hc0b39428, 32'hc28c63de};
test_output[1038] = '{32'h42b024f0};
test_index[1038] = '{3};
test_input[8312:8319] = '{32'h4257a871, 32'hc2534b74, 32'hc24c7cc6, 32'h4239104b, 32'hc2977420, 32'hc1fa4d0c, 32'h41525b9d, 32'hc263b0d1};
test_output[1039] = '{32'h4257a871};
test_index[1039] = '{0};
test_input[8320:8327] = '{32'h42b9b2a5, 32'hc2b502ce, 32'h42aa208e, 32'h40e218ec, 32'h42a79cd7, 32'hc00cdea8, 32'h428a04eb, 32'h421e8473};
test_output[1040] = '{32'h42b9b2a5};
test_index[1040] = '{0};
test_input[8328:8335] = '{32'h418952fe, 32'hc2b5caf9, 32'h40ed3c37, 32'hc2219490, 32'h4158e544, 32'hc235dd23, 32'h4204143c, 32'h428f5056};
test_output[1041] = '{32'h428f5056};
test_index[1041] = '{7};
test_input[8336:8343] = '{32'hc1927c29, 32'h42c7ebbf, 32'hc2070c60, 32'hc2c50d2a, 32'hc0d926ae, 32'hc2a04e43, 32'hc1f7bb24, 32'hc218e389};
test_output[1042] = '{32'h42c7ebbf};
test_index[1042] = '{1};
test_input[8344:8351] = '{32'h425d6454, 32'hc2503d31, 32'hc2006d4e, 32'hc22b39a5, 32'h428e28d8, 32'h42b20731, 32'h422b8f98, 32'hc246e87b};
test_output[1043] = '{32'h42b20731};
test_index[1043] = '{5};
test_input[8352:8359] = '{32'hc196f406, 32'hc27d2028, 32'hc17d9119, 32'h42b7905c, 32'hc2451d99, 32'hc26c04b9, 32'h40d5c7d8, 32'h41782930};
test_output[1044] = '{32'h42b7905c};
test_index[1044] = '{3};
test_input[8360:8367] = '{32'h42a3af7d, 32'hc29265f2, 32'hc1fd4a1a, 32'h427e9fc1, 32'h428a029b, 32'h41ae9280, 32'hc191954a, 32'hc24ad38a};
test_output[1045] = '{32'h42a3af7d};
test_index[1045] = '{0};
test_input[8368:8375] = '{32'h41730de8, 32'hc127f16c, 32'hc29693be, 32'hc23b9da7, 32'h42b2b88c, 32'hc1ca8dbc, 32'hc21a9453, 32'h4231e3cc};
test_output[1046] = '{32'h42b2b88c};
test_index[1046] = '{4};
test_input[8376:8383] = '{32'hc268578d, 32'h4240c421, 32'hc2a420b4, 32'hc29ce306, 32'h42b601e6, 32'h4033286a, 32'h4253fc1b, 32'h4295d5e7};
test_output[1047] = '{32'h42b601e6};
test_index[1047] = '{4};
test_input[8384:8391] = '{32'hc0b11bb2, 32'h41c1fca5, 32'h41e0566a, 32'hc218eaea, 32'hc2130560, 32'h421190c2, 32'hc2083cf8, 32'h42bd94d8};
test_output[1048] = '{32'h42bd94d8};
test_index[1048] = '{7};
test_input[8392:8399] = '{32'h42311bab, 32'hc2687262, 32'hbfcc6595, 32'hc188c40a, 32'h41097128, 32'hc1d21b14, 32'hc16c7ca9, 32'hc2a16e13};
test_output[1049] = '{32'h42311bab};
test_index[1049] = '{0};
test_input[8400:8407] = '{32'h425e82de, 32'hc11c7f11, 32'hc29eb589, 32'h425b0c6a, 32'hc2008638, 32'hc1a24e53, 32'h3d9dd594, 32'hc1a74a80};
test_output[1050] = '{32'h425e82de};
test_index[1050] = '{0};
test_input[8408:8415] = '{32'h42449705, 32'hc2379f01, 32'hc265fdca, 32'hc2b34999, 32'hc2836583, 32'h4296a515, 32'h42c409f7, 32'hc29d4548};
test_output[1051] = '{32'h42c409f7};
test_index[1051] = '{6};
test_input[8416:8423] = '{32'hc2220f15, 32'h42463cbf, 32'h429f0608, 32'h42bbb079, 32'hc27e0a64, 32'hc26f1a07, 32'hbfc685bb, 32'h42251ee9};
test_output[1052] = '{32'h42bbb079};
test_index[1052] = '{3};
test_input[8424:8431] = '{32'hc273c498, 32'h3fc0bebe, 32'h42ad63b8, 32'hc1d8d3ff, 32'h4213d781, 32'hc2ad1690, 32'hc2bdf6c8, 32'h4201e066};
test_output[1053] = '{32'h42ad63b8};
test_index[1053] = '{2};
test_input[8432:8439] = '{32'hc1ffd7e5, 32'hc25118ab, 32'hc19cc5b3, 32'hc02e33fd, 32'hc299619a, 32'hc2bd1123, 32'h42766844, 32'hc2974424};
test_output[1054] = '{32'h42766844};
test_index[1054] = '{6};
test_input[8440:8447] = '{32'h42a49056, 32'h42b352a1, 32'h3ff4e3b9, 32'h426d22a3, 32'hc206ae67, 32'h42b9ed6a, 32'h41fa3286, 32'hc085d632};
test_output[1055] = '{32'h42b9ed6a};
test_index[1055] = '{5};
test_input[8448:8455] = '{32'h4285cc3d, 32'h421f73a4, 32'hc28c3883, 32'h42acc8d2, 32'h4239932e, 32'hc235e987, 32'hc284cd8b, 32'h41c12690};
test_output[1056] = '{32'h42acc8d2};
test_index[1056] = '{3};
test_input[8456:8463] = '{32'h426c486f, 32'hc1ac2ff8, 32'h413cc68a, 32'hc28f3ef6, 32'hc293fe9f, 32'h42918ce4, 32'hc278ce7a, 32'h4235507f};
test_output[1057] = '{32'h42918ce4};
test_index[1057] = '{5};
test_input[8464:8471] = '{32'h42b4a788, 32'h4270480a, 32'h4289a683, 32'hc2c1961a, 32'h42ac8cc7, 32'h42bf3ba1, 32'hc2b65326, 32'h41e6a078};
test_output[1058] = '{32'h42bf3ba1};
test_index[1058] = '{5};
test_input[8472:8479] = '{32'h4236433b, 32'h4260d824, 32'hc2a555e0, 32'h42ac992a, 32'h4290e4f8, 32'h42490024, 32'hc203801f, 32'h40dbc321};
test_output[1059] = '{32'h42ac992a};
test_index[1059] = '{3};
test_input[8480:8487] = '{32'hc24b7169, 32'hc1b83c59, 32'h42211f7a, 32'h42b258bf, 32'hc27e2b1c, 32'h42a6eb67, 32'h4198d446, 32'hc28f8842};
test_output[1060] = '{32'h42b258bf};
test_index[1060] = '{3};
test_input[8488:8495] = '{32'h42757d56, 32'hc15f44a3, 32'hc1dffa92, 32'hc18efbf3, 32'h4218b3eb, 32'h4226f03d, 32'h42a11509, 32'hc25697bb};
test_output[1061] = '{32'h42a11509};
test_index[1061] = '{6};
test_input[8496:8503] = '{32'hc2aa88c9, 32'h414c4e92, 32'h421e7ff1, 32'h4288a9db, 32'h42b80de1, 32'h41e6e52b, 32'h42839d42, 32'h41856e7e};
test_output[1062] = '{32'h42b80de1};
test_index[1062] = '{4};
test_input[8504:8511] = '{32'h428c21cb, 32'h42737919, 32'hc28ed98f, 32'hbffc3d8d, 32'h42be02f4, 32'h429d9013, 32'hc1278b7b, 32'h421a960d};
test_output[1063] = '{32'h42be02f4};
test_index[1063] = '{4};
test_input[8512:8519] = '{32'h420b2f2c, 32'hc25ba8ba, 32'h41d979c0, 32'h41d52382, 32'hc051dcdb, 32'hc186fa97, 32'hc260f886, 32'hc27bdffc};
test_output[1064] = '{32'h420b2f2c};
test_index[1064] = '{0};
test_input[8520:8527] = '{32'h427ff8fb, 32'h4298de91, 32'h4183c50e, 32'hc234efc3, 32'h42979f6f, 32'hc2083446, 32'h42392361, 32'h41c456b9};
test_output[1065] = '{32'h4298de91};
test_index[1065] = '{1};
test_input[8528:8535] = '{32'h42a4a31f, 32'h42133c25, 32'h412a2c39, 32'h4281361b, 32'hc2741e0d, 32'h4298afc4, 32'hc1dd9c28, 32'hc193d60b};
test_output[1066] = '{32'h42a4a31f};
test_index[1066] = '{0};
test_input[8536:8543] = '{32'h4261d1c7, 32'hc2bf8c4c, 32'hc2a101fb, 32'h41e6cb6b, 32'hc29cf531, 32'h4292ccca, 32'h4148fcc6, 32'hc274d3ef};
test_output[1067] = '{32'h4292ccca};
test_index[1067] = '{5};
test_input[8544:8551] = '{32'h4295e909, 32'h4025ad85, 32'h42a26653, 32'hc2196e80, 32'h41f12bb6, 32'hc1db7bc5, 32'h420f9460, 32'h428d63e4};
test_output[1068] = '{32'h42a26653};
test_index[1068] = '{2};
test_input[8552:8559] = '{32'hc27f8b41, 32'hc2b78dba, 32'hbff036e0, 32'hc25e4fd6, 32'h41896b7f, 32'h41621a35, 32'hc299ab56, 32'h42129cbb};
test_output[1069] = '{32'h42129cbb};
test_index[1069] = '{7};
test_input[8560:8567] = '{32'hc15f8054, 32'h420aa923, 32'h4281914b, 32'hc11c9d4b, 32'h41a243df, 32'hc2908cb6, 32'hc1c61ac7, 32'h42b56eaf};
test_output[1070] = '{32'h42b56eaf};
test_index[1070] = '{7};
test_input[8568:8575] = '{32'hc10c4586, 32'h402bf9fb, 32'hc1f7886e, 32'h427d55fb, 32'hc002a3b4, 32'h4249bb45, 32'hc2195df4, 32'h4181ca4b};
test_output[1071] = '{32'h427d55fb};
test_index[1071] = '{3};
test_input[8576:8583] = '{32'hc2b087f6, 32'hc1ad3161, 32'hc297861a, 32'hc0d351a7, 32'h426e0ee4, 32'hc20053eb, 32'hc2b6ad4c, 32'h42417233};
test_output[1072] = '{32'h426e0ee4};
test_index[1072] = '{4};
test_input[8584:8591] = '{32'hc15565c4, 32'hc1d83c2a, 32'hc220c60f, 32'hc1c2b19b, 32'h426e84b3, 32'hc1fdfb99, 32'hc2bbba01, 32'hc26a58ef};
test_output[1073] = '{32'h426e84b3};
test_index[1073] = '{4};
test_input[8592:8599] = '{32'hc161694d, 32'hc180f71d, 32'hc1f77fc7, 32'h414ed4a3, 32'h4236e987, 32'hc17a1b5b, 32'hc29bc70c, 32'h3f037e1c};
test_output[1074] = '{32'h4236e987};
test_index[1074] = '{4};
test_input[8600:8607] = '{32'hc1b3514e, 32'h402f7156, 32'h42a181b5, 32'h42a3d994, 32'hc0c7a75d, 32'h420fc77e, 32'hc24a95bc, 32'hc0cb7b89};
test_output[1075] = '{32'h42a3d994};
test_index[1075] = '{3};
test_input[8608:8615] = '{32'h42c5b8ef, 32'h4209ca0b, 32'h425cca69, 32'hc2c574cb, 32'hc2b9f47c, 32'h41798cfd, 32'hc259e62d, 32'h426298c4};
test_output[1076] = '{32'h42c5b8ef};
test_index[1076] = '{0};
test_input[8616:8623] = '{32'hc11790a1, 32'h42b84934, 32'h4242dcec, 32'hc27d825a, 32'hc0fd209f, 32'hc21c38da, 32'hc2aee95d, 32'h421c4b50};
test_output[1077] = '{32'h42b84934};
test_index[1077] = '{1};
test_input[8624:8631] = '{32'hc29d268e, 32'h41f6b3ef, 32'h41abca1e, 32'h4289d1ef, 32'h426c80de, 32'hc234d5d6, 32'hc19a3d5f, 32'h40645956};
test_output[1078] = '{32'h4289d1ef};
test_index[1078] = '{3};
test_input[8632:8639] = '{32'hc247da01, 32'h426226d9, 32'hc1e92d68, 32'hc28097b1, 32'h40d84fc3, 32'hc168666e, 32'hc0280539, 32'h40cb84fc};
test_output[1079] = '{32'h426226d9};
test_index[1079] = '{1};
test_input[8640:8647] = '{32'h42b10c77, 32'hc2b4e18b, 32'h4106016f, 32'h3f88f318, 32'hc09d2970, 32'hc2be9afe, 32'hc20ad76f, 32'h42bc362e};
test_output[1080] = '{32'h42bc362e};
test_index[1080] = '{7};
test_input[8648:8655] = '{32'hc272d395, 32'h429fb006, 32'hc23e7ca1, 32'h421f1a7c, 32'h4197de0d, 32'hc23c5edc, 32'h4282747b, 32'h41c7d59b};
test_output[1081] = '{32'h429fb006};
test_index[1081] = '{1};
test_input[8656:8663] = '{32'hc1ac2d17, 32'hc2c3625d, 32'hc2c0be5c, 32'hbf19d7b9, 32'h4291a6e4, 32'hc2b16fc6, 32'hc0b23fdb, 32'hc2a42d90};
test_output[1082] = '{32'h4291a6e4};
test_index[1082] = '{4};
test_input[8664:8671] = '{32'h424b731e, 32'h41aae02e, 32'h42b9f5bd, 32'hc298a1db, 32'h4284933b, 32'hc19b6659, 32'hc1920569, 32'hc2635283};
test_output[1083] = '{32'h42b9f5bd};
test_index[1083] = '{2};
test_input[8672:8679] = '{32'hc2968ae0, 32'h42abade0, 32'hc16680c1, 32'hc2892e48, 32'h42916758, 32'hc1de3057, 32'h40f5150b, 32'hc29ee929};
test_output[1084] = '{32'h42abade0};
test_index[1084] = '{1};
test_input[8680:8687] = '{32'hc2b664c1, 32'hc1a1fe39, 32'h42c7007e, 32'h42234fe5, 32'h42162f9c, 32'hc247d193, 32'hc207262f, 32'h42a8d24e};
test_output[1085] = '{32'h42c7007e};
test_index[1085] = '{2};
test_input[8688:8695] = '{32'hc210d9c7, 32'hc263b084, 32'hc26af094, 32'h42b66426, 32'h42510d4b, 32'hc29adb57, 32'hc281826d, 32'h429180e3};
test_output[1086] = '{32'h42b66426};
test_index[1086] = '{3};
test_input[8696:8703] = '{32'hc26680ba, 32'h427e32b7, 32'h420c0432, 32'h42ae117f, 32'h42829ea4, 32'h42a50a8b, 32'hc2492cf0, 32'h41b7b334};
test_output[1087] = '{32'h42ae117f};
test_index[1087] = '{3};
test_input[8704:8711] = '{32'h42a3b7b3, 32'hc2881099, 32'hc2578493, 32'h42327c30, 32'h426f161c, 32'h42ba3279, 32'hc231dcd2, 32'h42a79728};
test_output[1088] = '{32'h42ba3279};
test_index[1088] = '{5};
test_input[8712:8719] = '{32'hc23ceec6, 32'hc25c64d4, 32'hc0ef806e, 32'h421afd4b, 32'hc29a6797, 32'h41e1960c, 32'hc1849194, 32'h42ac63ee};
test_output[1089] = '{32'h42ac63ee};
test_index[1089] = '{7};
test_input[8720:8727] = '{32'hc284614b, 32'h41eab7cc, 32'h428edd1f, 32'h412123af, 32'hc1001aba, 32'hc2874da7, 32'hc285e1ab, 32'h42a85dd2};
test_output[1090] = '{32'h42a85dd2};
test_index[1090] = '{7};
test_input[8728:8735] = '{32'hc259536d, 32'hc29a483e, 32'hc289ac8c, 32'hc1bea723, 32'h41006724, 32'h4222d7fc, 32'hc1065eed, 32'h41ea0f70};
test_output[1091] = '{32'h4222d7fc};
test_index[1091] = '{5};
test_input[8736:8743] = '{32'h4274e89c, 32'h4201bff1, 32'h42c67ee0, 32'hc2ae269d, 32'h41b88c6a, 32'h42a598c1, 32'hc2a46b4b, 32'h41b53677};
test_output[1092] = '{32'h42c67ee0};
test_index[1092] = '{2};
test_input[8744:8751] = '{32'hc261aef3, 32'h421cfd4f, 32'h42a1563a, 32'hc18ffe28, 32'h40ffdff2, 32'hc282f522, 32'hc042fe24, 32'hc1b59fd0};
test_output[1093] = '{32'h42a1563a};
test_index[1093] = '{2};
test_input[8752:8759] = '{32'h408287a6, 32'h41b4918e, 32'h420dbb17, 32'hc2b82941, 32'h42894f11, 32'h429a4d80, 32'hc29b0d4f, 32'h429e4666};
test_output[1094] = '{32'h429e4666};
test_index[1094] = '{7};
test_input[8760:8767] = '{32'hc2548ae1, 32'hc25063a9, 32'hc288999b, 32'hc2918cb8, 32'hc1e360cf, 32'hc081c33f, 32'hc2914e24, 32'hc23195a8};
test_output[1095] = '{32'hc081c33f};
test_index[1095] = '{5};
test_input[8768:8775] = '{32'hc221b96a, 32'hc21023db, 32'hc29d3e6b, 32'hc1cb5b13, 32'hc22331d8, 32'h429ec297, 32'hc1cfbc65, 32'hc220599f};
test_output[1096] = '{32'h429ec297};
test_index[1096] = '{5};
test_input[8776:8783] = '{32'h421607e0, 32'h4227f22b, 32'hc1f634d9, 32'hc2be466f, 32'h41a4aa3a, 32'hc2c5bd29, 32'h429f379f, 32'h42b359c4};
test_output[1097] = '{32'h42b359c4};
test_index[1097] = '{7};
test_input[8784:8791] = '{32'hc2aa0f3d, 32'h425ba766, 32'h429913de, 32'hc2a6fe2b, 32'hc2a2d512, 32'h41873c1b, 32'h418d2354, 32'hc2829de0};
test_output[1098] = '{32'h429913de};
test_index[1098] = '{2};
test_input[8792:8799] = '{32'hc2656158, 32'hc280d6fa, 32'hc214db02, 32'h420e7330, 32'hc2b712de, 32'hc2a37132, 32'hbfc4664d, 32'h41a4ac03};
test_output[1099] = '{32'h420e7330};
test_index[1099] = '{3};
test_input[8800:8807] = '{32'hc2b73408, 32'hc1d69f43, 32'hc2c4da8f, 32'hc2b6240f, 32'hc0680045, 32'hc2a47001, 32'h428333ae, 32'h4219724d};
test_output[1100] = '{32'h428333ae};
test_index[1100] = '{6};
test_input[8808:8815] = '{32'hc2ba64ce, 32'h41ff46cb, 32'h42b84082, 32'h3fc63d62, 32'hc0f55244, 32'hc12e72d8, 32'h41a1a3f0, 32'hc1ee982e};
test_output[1101] = '{32'h42b84082};
test_index[1101] = '{2};
test_input[8816:8823] = '{32'h41cb3362, 32'hc2472897, 32'h429f35be, 32'hc1f935a5, 32'hc2603e4f, 32'h42491132, 32'h42918779, 32'hc27f3483};
test_output[1102] = '{32'h429f35be};
test_index[1102] = '{2};
test_input[8824:8831] = '{32'hc2b06d19, 32'h4295e171, 32'h4138c5f4, 32'h425c5f81, 32'hc1bba0f9, 32'h427957d9, 32'h41ed3c4f, 32'hc274aba3};
test_output[1103] = '{32'h4295e171};
test_index[1103] = '{1};
test_input[8832:8839] = '{32'h42b45969, 32'hc264b79a, 32'hc1986e6b, 32'hc2a575b4, 32'h42c2f53e, 32'h4226ee4f, 32'h42a88509, 32'h423ed2b8};
test_output[1104] = '{32'h42c2f53e};
test_index[1104] = '{4};
test_input[8840:8847] = '{32'h417218c2, 32'h423943af, 32'h426dad0b, 32'hc24fe5d7, 32'hc2379a24, 32'hc16e1aa5, 32'hc2b2455b, 32'h4228b60b};
test_output[1105] = '{32'h426dad0b};
test_index[1105] = '{2};
test_input[8848:8855] = '{32'h425ccda9, 32'hc29bc1e7, 32'hc21ddbe6, 32'h41d2b048, 32'h428e6a0a, 32'h42143519, 32'h42313534, 32'hc239c766};
test_output[1106] = '{32'h428e6a0a};
test_index[1106] = '{4};
test_input[8856:8863] = '{32'h42a44d77, 32'hc2542ff0, 32'h42134a80, 32'h42c1eeaf, 32'hc25adede, 32'hc10d8270, 32'hc091af7a, 32'h42c0fa0c};
test_output[1107] = '{32'h42c1eeaf};
test_index[1107] = '{3};
test_input[8864:8871] = '{32'hc233b28a, 32'hc2c28cd4, 32'h4111b505, 32'h40511a66, 32'hc27d828d, 32'hc169470d, 32'hc2053a44, 32'h416e6f00};
test_output[1108] = '{32'h416e6f00};
test_index[1108] = '{7};
test_input[8872:8879] = '{32'h42aa1a2e, 32'h42b09da8, 32'h42a7226c, 32'h4290740a, 32'h429ec0be, 32'h422366f8, 32'h40c1ce84, 32'h424a6365};
test_output[1109] = '{32'h42b09da8};
test_index[1109] = '{1};
test_input[8880:8887] = '{32'h425ccf3a, 32'h426c4497, 32'h3fb1bafc, 32'hc298ea6e, 32'h4233da27, 32'hc2a93da0, 32'hc2b08340, 32'hc2165034};
test_output[1110] = '{32'h426c4497};
test_index[1110] = '{1};
test_input[8888:8895] = '{32'hc2227950, 32'h425dfdba, 32'hc2ba2ce1, 32'hc29ee104, 32'hc239724d, 32'hc1a1f3b4, 32'h3dbe5f76, 32'hc2925857};
test_output[1111] = '{32'h425dfdba};
test_index[1111] = '{1};
test_input[8896:8903] = '{32'hc2a74ef0, 32'h42c43445, 32'h4296ca8b, 32'hc28719e8, 32'hc20e0aeb, 32'h428ff75d, 32'hbde41f13, 32'hc2a37dd2};
test_output[1112] = '{32'h42c43445};
test_index[1112] = '{1};
test_input[8904:8911] = '{32'hc28f3ef5, 32'hc27cc6bf, 32'hc2b70359, 32'h42014e28, 32'hc23e2707, 32'hc2b45a6b, 32'hc2b952f9, 32'h428c1b0c};
test_output[1113] = '{32'h428c1b0c};
test_index[1113] = '{7};
test_input[8912:8919] = '{32'hc2765df4, 32'h424a03a8, 32'hc28c2eee, 32'h41e895a2, 32'hc2b1e353, 32'h418d3c25, 32'hc1c55099, 32'h401dd4e1};
test_output[1114] = '{32'h424a03a8};
test_index[1114] = '{1};
test_input[8920:8927] = '{32'h41a6f0e9, 32'hc2addb85, 32'h4129fa2a, 32'h41fd4a42, 32'hc1ecdd0f, 32'h41a97d7b, 32'hc1c2f56b, 32'hc21174d4};
test_output[1115] = '{32'h41fd4a42};
test_index[1115] = '{3};
test_input[8928:8935] = '{32'hc2af9bf0, 32'hc2bacd5b, 32'hc25ae67f, 32'h42a61b55, 32'hc1e87489, 32'hc27f7be3, 32'h4117bfb6, 32'h404c4cff};
test_output[1116] = '{32'h42a61b55};
test_index[1116] = '{3};
test_input[8936:8943] = '{32'h427b842a, 32'h4251236b, 32'h40ca8404, 32'h423f3e46, 32'h3d28cbfa, 32'hc0a5bcbc, 32'hc2af02c1, 32'h42b64d8b};
test_output[1117] = '{32'h42b64d8b};
test_index[1117] = '{7};
test_input[8944:8951] = '{32'h4288e253, 32'h420f45f6, 32'hc25a17e9, 32'hbe63590b, 32'h4111cc70, 32'h42a9d13d, 32'hc26d5944, 32'h4156ca3b};
test_output[1118] = '{32'h42a9d13d};
test_index[1118] = '{5};
test_input[8952:8959] = '{32'h4259e241, 32'hc28eecee, 32'h4286b521, 32'h41c6dfb5, 32'hc28cd453, 32'h425143ce, 32'h418ded97, 32'h424c0f14};
test_output[1119] = '{32'h4286b521};
test_index[1119] = '{2};
test_input[8960:8967] = '{32'hc28a6ac1, 32'hc2a6b879, 32'h41f75a6b, 32'hc1509de2, 32'h3fdc2dd2, 32'h42b29d5e, 32'h42b32263, 32'h42c4bfbe};
test_output[1120] = '{32'h42c4bfbe};
test_index[1120] = '{7};
test_input[8968:8975] = '{32'h41750f5d, 32'hc2a3d72c, 32'h413978f5, 32'h42856f5f, 32'h425a86ff, 32'h428d6a8a, 32'h42012653, 32'h4121614e};
test_output[1121] = '{32'h428d6a8a};
test_index[1121] = '{5};
test_input[8976:8983] = '{32'hc28d871c, 32'h42acdfc4, 32'h42bdfeb4, 32'hc206e612, 32'hc26a42a5, 32'hc2b1ce0b, 32'h429dcbfc, 32'hc2b37c49};
test_output[1122] = '{32'h42bdfeb4};
test_index[1122] = '{2};
test_input[8984:8991] = '{32'hc2b27a98, 32'h42a1095c, 32'hc2c4c952, 32'hc2007ade, 32'hc1b98fc4, 32'h422c7b27, 32'h427b2cf6, 32'h41ac98d7};
test_output[1123] = '{32'h42a1095c};
test_index[1123] = '{1};
test_input[8992:8999] = '{32'hc1c90764, 32'h42b0cf4e, 32'hc290e7d1, 32'hc2a79594, 32'hc2c2d738, 32'hc1c8d15b, 32'h42c44a8a, 32'hc0435e6f};
test_output[1124] = '{32'h42c44a8a};
test_index[1124] = '{6};
test_input[9000:9007] = '{32'hc2907b89, 32'hc24a38c7, 32'h41c5a3a9, 32'h424aefa6, 32'hc288519b, 32'hc23aac03, 32'h425fcb52, 32'h42941486};
test_output[1125] = '{32'h42941486};
test_index[1125] = '{7};
test_input[9008:9015] = '{32'hc2ae4f0a, 32'hc150b789, 32'hc29146dd, 32'hc19d8376, 32'hc1f9a875, 32'h41d13753, 32'h42841e07, 32'hc23a5725};
test_output[1126] = '{32'h42841e07};
test_index[1126] = '{6};
test_input[9016:9023] = '{32'h42977959, 32'h428eea87, 32'h42158cf6, 32'hc21bacd6, 32'hc28e4026, 32'hc2c4a0cb, 32'hc2bfbc81, 32'hc24da4dd};
test_output[1127] = '{32'h42977959};
test_index[1127] = '{0};
test_input[9024:9031] = '{32'hc2525db4, 32'hc21119b3, 32'h42b2229d, 32'h42a19248, 32'hc1e2ca01, 32'hc288b824, 32'hc2c24558, 32'hc204face};
test_output[1128] = '{32'h42b2229d};
test_index[1128] = '{2};
test_input[9032:9039] = '{32'h42470fbd, 32'h42aa44d7, 32'h423d9ab4, 32'hc1bba67c, 32'hc2c1c091, 32'hc1dd0d24, 32'hc29d5a0d, 32'hc219a347};
test_output[1129] = '{32'h42aa44d7};
test_index[1129] = '{1};
test_input[9040:9047] = '{32'h420dee97, 32'h41de4c95, 32'h42c462be, 32'hc29b69e3, 32'h41d21807, 32'hc22958af, 32'h42c21c24, 32'h42c45b2f};
test_output[1130] = '{32'h42c462be};
test_index[1130] = '{2};
test_input[9048:9055] = '{32'hc2a90454, 32'h42927a3a, 32'hc2ae8a93, 32'hc16d5034, 32'h42354850, 32'hc2aff678, 32'h42b789e0, 32'hc0855276};
test_output[1131] = '{32'h42b789e0};
test_index[1131] = '{6};
test_input[9056:9063] = '{32'hc28311a4, 32'hc10f3692, 32'h42351728, 32'hc24088c3, 32'h42b2bd8a, 32'h4127428e, 32'h42b9b7de, 32'hc1a583ac};
test_output[1132] = '{32'h42b9b7de};
test_index[1132] = '{6};
test_input[9064:9071] = '{32'hc1c69532, 32'hc17a272e, 32'h423f5c3f, 32'hc27e7e3c, 32'hc2930ee0, 32'hc12cccfe, 32'hbee6f832, 32'hbff4b583};
test_output[1133] = '{32'h423f5c3f};
test_index[1133] = '{2};
test_input[9072:9079] = '{32'h41972358, 32'h4193278f, 32'h42b16695, 32'hc2a3206c, 32'hc2b54cc0, 32'h42c781a6, 32'h427041ba, 32'h40eb0c20};
test_output[1134] = '{32'h42c781a6};
test_index[1134] = '{5};
test_input[9080:9087] = '{32'h42ab1222, 32'hc1da3b82, 32'hc04da711, 32'hc24cdd27, 32'hc278a9e7, 32'hc2b2263c, 32'h4285ee52, 32'hc27ea275};
test_output[1135] = '{32'h42ab1222};
test_index[1135] = '{0};
test_input[9088:9095] = '{32'h4258d160, 32'hc2c301c9, 32'h428bda33, 32'hc2c04d3e, 32'hc21c574c, 32'hc28d9e1a, 32'h4234f614, 32'hc11a76c5};
test_output[1136] = '{32'h428bda33};
test_index[1136] = '{2};
test_input[9096:9103] = '{32'hc20bd5dc, 32'h42a51d48, 32'h42554ed8, 32'h42bb5c5f, 32'hc27e725f, 32'h41f4b3e7, 32'h422d25c4, 32'h42a55d02};
test_output[1137] = '{32'h42bb5c5f};
test_index[1137] = '{3};
test_input[9104:9111] = '{32'hc1d2a251, 32'hc23ecdaf, 32'h41cca60a, 32'h42a8989d, 32'hc102144b, 32'h41ba9614, 32'h423ca6e9, 32'h427f06c8};
test_output[1138] = '{32'h42a8989d};
test_index[1138] = '{3};
test_input[9112:9119] = '{32'hc2836d8e, 32'hc2905fbb, 32'h42a8ece5, 32'h41990f4c, 32'hc215c2ad, 32'hc25f0399, 32'hc1100542, 32'hc1f3d8fd};
test_output[1139] = '{32'h42a8ece5};
test_index[1139] = '{2};
test_input[9120:9127] = '{32'h42937f81, 32'h41a0e912, 32'hc1d5c8c5, 32'hc2ac4b9c, 32'h410511d4, 32'h4199dda5, 32'h42695c47, 32'h4144a99d};
test_output[1140] = '{32'h42937f81};
test_index[1140] = '{0};
test_input[9128:9135] = '{32'h42c51ce8, 32'hc28f0cfb, 32'hc2150fce, 32'hc28b6e77, 32'h42526ee8, 32'hc1ba4c30, 32'h42c14bc3, 32'h424b550d};
test_output[1141] = '{32'h42c51ce8};
test_index[1141] = '{0};
test_input[9136:9143] = '{32'h4222b5d6, 32'hc2a97e8b, 32'h4276c48a, 32'h419a2387, 32'h4239524f, 32'hc2941ef5, 32'hc1f5a233, 32'h429fb7cf};
test_output[1142] = '{32'h429fb7cf};
test_index[1142] = '{7};
test_input[9144:9151] = '{32'hc23a4bd2, 32'h42b09218, 32'hc22cd686, 32'hc2bfdbac, 32'h42bad9a6, 32'hc287173f, 32'hc2067787, 32'hc1afe052};
test_output[1143] = '{32'h42bad9a6};
test_index[1143] = '{4};
test_input[9152:9159] = '{32'hc1babfeb, 32'hc285e2a3, 32'h41f52288, 32'h4259e2b4, 32'hc2730a5f, 32'hc28894b7, 32'hc273f6c5, 32'hc211b44d};
test_output[1144] = '{32'h4259e2b4};
test_index[1144] = '{3};
test_input[9160:9167] = '{32'hc2044de4, 32'hc26f1d66, 32'hc20ef471, 32'h422a3c3d, 32'h41df041a, 32'hc23fc39a, 32'h4266f3a1, 32'hbfa765a0};
test_output[1145] = '{32'h4266f3a1};
test_index[1145] = '{6};
test_input[9168:9175] = '{32'hc1363bf4, 32'hc2b8e083, 32'hc0054acc, 32'h423bb873, 32'hc0f9aef6, 32'hc1ebe501, 32'hc292110e, 32'hc0a6508d};
test_output[1146] = '{32'h423bb873};
test_index[1146] = '{3};
test_input[9176:9183] = '{32'h42687c28, 32'hc1d9077c, 32'hc28ce329, 32'hc28d7fd0, 32'hc25f8ec1, 32'hc18d2eec, 32'hc1c2117f, 32'h41fcf328};
test_output[1147] = '{32'h42687c28};
test_index[1147] = '{0};
test_input[9184:9191] = '{32'h41446618, 32'hc28f68a9, 32'hc2571df9, 32'hc27852cb, 32'h421e1944, 32'h42b79ce5, 32'hc2609eac, 32'h429c4a0e};
test_output[1148] = '{32'h42b79ce5};
test_index[1148] = '{5};
test_input[9192:9199] = '{32'hc208c09f, 32'h40ac010c, 32'h4204e09f, 32'h42678cde, 32'hc225c5b1, 32'hc2a8b559, 32'h420058b9, 32'hc14a30d4};
test_output[1149] = '{32'h42678cde};
test_index[1149] = '{3};
test_input[9200:9207] = '{32'hc10c9554, 32'h41f0cb23, 32'h42998aad, 32'hc102b3d1, 32'h4270ad19, 32'hc2b2b876, 32'h422ebe26, 32'hc1ac0ba2};
test_output[1150] = '{32'h42998aad};
test_index[1150] = '{2};
test_input[9208:9215] = '{32'h429fd622, 32'hc268e032, 32'h420ef701, 32'hc294498e, 32'h42977dbe, 32'h429a9457, 32'hc2bce5f2, 32'hc2877d8a};
test_output[1151] = '{32'h429fd622};
test_index[1151] = '{0};
test_input[9216:9223] = '{32'h416de7cc, 32'h4287f14a, 32'hc2379030, 32'hc02ca4ad, 32'h42285bb5, 32'hc22cd589, 32'h419611e6, 32'hc2b46c30};
test_output[1152] = '{32'h4287f14a};
test_index[1152] = '{1};
test_input[9224:9231] = '{32'hc1976ed2, 32'h422b47d0, 32'hc24cf1bd, 32'hc1322560, 32'h4217902b, 32'hc1c5c01e, 32'hc20e7a60, 32'hc1b218ee};
test_output[1153] = '{32'h422b47d0};
test_index[1153] = '{1};
test_input[9232:9239] = '{32'hc27c910e, 32'hc2a27739, 32'h424caa03, 32'h41b3f762, 32'hc2bee583, 32'h42328cca, 32'h413b6305, 32'hc26eedae};
test_output[1154] = '{32'h424caa03};
test_index[1154] = '{2};
test_input[9240:9247] = '{32'h428e89bc, 32'h41bfca94, 32'h420e8118, 32'hc24643e2, 32'hc0f629ef, 32'h42916ffc, 32'hc12ba526, 32'h41f847e1};
test_output[1155] = '{32'h42916ffc};
test_index[1155] = '{5};
test_input[9248:9255] = '{32'h4255f859, 32'h401dd1a4, 32'h426e386b, 32'h4292b02f, 32'hc2bea0a6, 32'hc22b0046, 32'hc28a3a1b, 32'hc2a26211};
test_output[1156] = '{32'h4292b02f};
test_index[1156] = '{3};
test_input[9256:9263] = '{32'hc1298f62, 32'h427d9a12, 32'hbed2def3, 32'hc2248f61, 32'h415f545e, 32'h428926a6, 32'hc0aebf3b, 32'hc2be911f};
test_output[1157] = '{32'h428926a6};
test_index[1157] = '{5};
test_input[9264:9271] = '{32'h4214ede2, 32'hc28810ee, 32'hc23a9af8, 32'h42a53ab5, 32'hc2c6b412, 32'h4278d83d, 32'hc2312e32, 32'hc2c15a88};
test_output[1158] = '{32'h42a53ab5};
test_index[1158] = '{3};
test_input[9272:9279] = '{32'h41a9ef8b, 32'hc250a10a, 32'hc0635c85, 32'hc27d62f3, 32'h41fac73a, 32'hc1f9973f, 32'hc2ae0a3d, 32'hc2215fc6};
test_output[1159] = '{32'h41fac73a};
test_index[1159] = '{4};
test_input[9280:9287] = '{32'hc18c518e, 32'h41f6c14a, 32'h4280f7fb, 32'h429f78d7, 32'hc1a7eca2, 32'h427d6598, 32'h42c3053a, 32'hc230122e};
test_output[1160] = '{32'h42c3053a};
test_index[1160] = '{6};
test_input[9288:9295] = '{32'h4207a266, 32'h423dd0b8, 32'h414a3c11, 32'hc01a476d, 32'hc2877963, 32'hc124780e, 32'hc26f4ca3, 32'hc27df8c4};
test_output[1161] = '{32'h423dd0b8};
test_index[1161] = '{1};
test_input[9296:9303] = '{32'hc27abd3c, 32'hc2666096, 32'hc24cc32d, 32'h429bfc58, 32'hc217acc7, 32'h41aa2a47, 32'h422f86d8, 32'hc21f80f4};
test_output[1162] = '{32'h429bfc58};
test_index[1162] = '{3};
test_input[9304:9311] = '{32'hc21a7b05, 32'h40b25875, 32'h40819edf, 32'hc1d447b6, 32'hc18d6a9d, 32'hc2c16205, 32'hc2220e1f, 32'hc2025ddf};
test_output[1163] = '{32'h40b25875};
test_index[1163] = '{1};
test_input[9312:9319] = '{32'h428da30c, 32'hc2992787, 32'hc29a305c, 32'h4290d4ad, 32'hc1df2652, 32'hc26531f3, 32'hc2ad0156, 32'hc1fb0900};
test_output[1164] = '{32'h4290d4ad};
test_index[1164] = '{3};
test_input[9320:9327] = '{32'h428aaf47, 32'h3f8011a9, 32'hc21e740b, 32'hc29fff95, 32'h42118af0, 32'h428d0be8, 32'h42b96c2a, 32'hc1c95870};
test_output[1165] = '{32'h42b96c2a};
test_index[1165] = '{6};
test_input[9328:9335] = '{32'h40391ea8, 32'h42a2f78b, 32'hc2289ea0, 32'h410d282d, 32'hbf06c18a, 32'h429e1b33, 32'hc1bc0669, 32'h418006c1};
test_output[1166] = '{32'h42a2f78b};
test_index[1166] = '{1};
test_input[9336:9343] = '{32'h41a2cd06, 32'hc2b4fd1c, 32'h428aabe2, 32'h404e0dd6, 32'hc2967964, 32'hbfa07390, 32'hc23a7c19, 32'hc151b152};
test_output[1167] = '{32'h428aabe2};
test_index[1167] = '{2};
test_input[9344:9351] = '{32'hc2797c10, 32'h426f3857, 32'hc2619e92, 32'hc117133e, 32'hc23d7a89, 32'h42c15612, 32'hc24f0d0d, 32'h42791d20};
test_output[1168] = '{32'h42c15612};
test_index[1168] = '{5};
test_input[9352:9359] = '{32'h41a4ac8e, 32'hc1be7d05, 32'h427ea308, 32'hc2961fc9, 32'hc1efdb08, 32'hc2813ace, 32'h426b952f, 32'hc26174cb};
test_output[1169] = '{32'h427ea308};
test_index[1169] = '{2};
test_input[9360:9367] = '{32'hc2c52c08, 32'h3f0dbb61, 32'hc2c1c0b4, 32'h425cf4b0, 32'h3f5ef744, 32'h41ac6822, 32'h4295b458, 32'hc0ccd605};
test_output[1170] = '{32'h4295b458};
test_index[1170] = '{6};
test_input[9368:9375] = '{32'hc209bacc, 32'hc23f0712, 32'h42313ba3, 32'hc20c6f46, 32'hc2c075e1, 32'h423ae4dd, 32'hc251cac5, 32'h4267c56e};
test_output[1171] = '{32'h4267c56e};
test_index[1171] = '{7};
test_input[9376:9383] = '{32'hc12f00f0, 32'h404333d8, 32'h4269bf81, 32'h42675fe3, 32'h40b19ff2, 32'hc18d1c52, 32'h42ad9d70, 32'hc286dcad};
test_output[1172] = '{32'h42ad9d70};
test_index[1172] = '{6};
test_input[9384:9391] = '{32'h4277bee8, 32'h4148cedb, 32'hc2b92947, 32'hc1b6af27, 32'hc2adbcaf, 32'h42b2ac6a, 32'h42134fb6, 32'hc0f55191};
test_output[1173] = '{32'h42b2ac6a};
test_index[1173] = '{5};
test_input[9392:9399] = '{32'h4288616d, 32'h40d1ac6c, 32'hc217c015, 32'h423b6db2, 32'h427b5560, 32'hc2bfe9f0, 32'hc23e81e9, 32'hc1aa6bf8};
test_output[1174] = '{32'h4288616d};
test_index[1174] = '{0};
test_input[9400:9407] = '{32'h4145fe05, 32'hc1b9bf9d, 32'h4104092e, 32'hc228a1d1, 32'hc2968d83, 32'hc2056d6e, 32'h4121bf54, 32'hc23dc7a2};
test_output[1175] = '{32'h4145fe05};
test_index[1175] = '{0};
test_input[9408:9415] = '{32'hc2b46101, 32'hc1f661dd, 32'hc29a1dd5, 32'hc2c75497, 32'hc1f0608d, 32'hc2c54c68, 32'hc28f0dac, 32'h424c5238};
test_output[1176] = '{32'h424c5238};
test_index[1176] = '{7};
test_input[9416:9423] = '{32'hc1a839ff, 32'hc26d0688, 32'hc2501997, 32'hc2c0118a, 32'h41f1a300, 32'hc14bcf05, 32'hc24b32a7, 32'hc2059404};
test_output[1177] = '{32'h41f1a300};
test_index[1177] = '{4};
test_input[9424:9431] = '{32'h425b96d5, 32'h41af8c63, 32'h3f4a9f93, 32'h410984eb, 32'h429c47d4, 32'hc29179e2, 32'hc085eaca, 32'h427f628a};
test_output[1178] = '{32'h429c47d4};
test_index[1178] = '{4};
test_input[9432:9439] = '{32'h42a26bb1, 32'h426167ff, 32'hc08bc97b, 32'h42bf751a, 32'h42a2ae00, 32'hc295c45a, 32'h42ad1eff, 32'hc246420b};
test_output[1179] = '{32'h42bf751a};
test_index[1179] = '{3};
test_input[9440:9447] = '{32'hc2a727cb, 32'h422f3b03, 32'hc1c76325, 32'h41ec7a7a, 32'h4280c0aa, 32'h429804e9, 32'h424151e7, 32'hc24dd4eb};
test_output[1180] = '{32'h429804e9};
test_index[1180] = '{5};
test_input[9448:9455] = '{32'hc2a88723, 32'hc28cafa5, 32'hc235c5d2, 32'hc2474f95, 32'hc217bda0, 32'hc0f23840, 32'h42030e30, 32'hc1fbe4cd};
test_output[1181] = '{32'h42030e30};
test_index[1181] = '{6};
test_input[9456:9463] = '{32'h42c01cea, 32'hc2c4b5ef, 32'h42413845, 32'h418f40e4, 32'h426a5aad, 32'h4149df84, 32'h4282e73c, 32'h42a1e6d8};
test_output[1182] = '{32'h42c01cea};
test_index[1182] = '{0};
test_input[9464:9471] = '{32'h4297a2a4, 32'hc1772696, 32'hc27518be, 32'hc274d483, 32'h42880890, 32'hbea3846b, 32'h4221941d, 32'hc27eb9cf};
test_output[1183] = '{32'h4297a2a4};
test_index[1183] = '{0};
test_input[9472:9479] = '{32'h4281511a, 32'h421adc0c, 32'hc270e9da, 32'hc1859029, 32'hc2a60f72, 32'h421b6fd6, 32'hc2bc5f70, 32'hc2a4625f};
test_output[1184] = '{32'h4281511a};
test_index[1184] = '{0};
test_input[9480:9487] = '{32'hc2a336e4, 32'hc1ba15ed, 32'h428941d9, 32'h420d94ca, 32'h42a82b13, 32'h40f7adca, 32'hc0b83c3c, 32'h4281a908};
test_output[1185] = '{32'h42a82b13};
test_index[1185] = '{4};
test_input[9488:9495] = '{32'h41642b99, 32'hc2b11978, 32'hc24207fe, 32'h422e9cdc, 32'hc21137ee, 32'h41956f63, 32'h426b7a8c, 32'h42c46915};
test_output[1186] = '{32'h42c46915};
test_index[1186] = '{7};
test_input[9496:9503] = '{32'hc287c6d7, 32'hc2a93298, 32'h421336f9, 32'hc1904572, 32'h418fa74c, 32'h409c4997, 32'h418548b2, 32'h3ed3c727};
test_output[1187] = '{32'h421336f9};
test_index[1187] = '{2};
test_input[9504:9511] = '{32'hc2b38f27, 32'h426eb33e, 32'h4197858a, 32'hc09ffaa9, 32'hc281100b, 32'h423be2f1, 32'h4281ee61, 32'hc298ee3a};
test_output[1188] = '{32'h4281ee61};
test_index[1188] = '{6};
test_input[9512:9519] = '{32'hbfd2d6c2, 32'h423c2bc4, 32'h422abeb4, 32'h42270010, 32'hc2630f1b, 32'hc10124e0, 32'h4240c936, 32'hc1886914};
test_output[1189] = '{32'h4240c936};
test_index[1189] = '{6};
test_input[9520:9527] = '{32'hc2bab81a, 32'h425db69a, 32'h42a04d4c, 32'hc2284da2, 32'h429ae21a, 32'hc270431f, 32'h3f12bbc4, 32'h422c4348};
test_output[1190] = '{32'h42a04d4c};
test_index[1190] = '{2};
test_input[9528:9535] = '{32'h422fd8a6, 32'hc244a3b6, 32'hc1c1cc2b, 32'hc19912fe, 32'h41e384ad, 32'h424d2d3a, 32'h41ef9261, 32'h42b950a0};
test_output[1191] = '{32'h42b950a0};
test_index[1191] = '{7};
test_input[9536:9543] = '{32'h426fa013, 32'h42973ced, 32'h42b2a1b5, 32'hc0c6bf30, 32'h41e2146f, 32'h400e10ee, 32'hc1a16c0f, 32'h41266601};
test_output[1192] = '{32'h42b2a1b5};
test_index[1192] = '{2};
test_input[9544:9551] = '{32'hc1a31f0a, 32'hc2132d51, 32'h4284e670, 32'h42941e0c, 32'h428b9221, 32'h418b6851, 32'h4201a7fd, 32'hc1955f7e};
test_output[1193] = '{32'h42941e0c};
test_index[1193] = '{3};
test_input[9552:9559] = '{32'hc19b07b2, 32'hc2b46547, 32'h429e49b1, 32'hc1816166, 32'h42414507, 32'h40c4d80d, 32'hc2aaf188, 32'hc1bff936};
test_output[1194] = '{32'h429e49b1};
test_index[1194] = '{2};
test_input[9560:9567] = '{32'hc1bd27f5, 32'h40b2a84b, 32'hc2c56cb4, 32'hc1f8edd3, 32'h42afd481, 32'h4214cff1, 32'h413808cb, 32'hc2588992};
test_output[1195] = '{32'h42afd481};
test_index[1195] = '{4};
test_input[9568:9575] = '{32'h425fdddc, 32'hc192fd77, 32'hc01a2b89, 32'h42488d13, 32'h42a3a18b, 32'h429d234d, 32'h41b770dc, 32'hbff88dfd};
test_output[1196] = '{32'h42a3a18b};
test_index[1196] = '{4};
test_input[9576:9583] = '{32'hc2b4fba1, 32'h428a3f31, 32'h41f702f9, 32'h42915231, 32'h40f87cfe, 32'hc24f0377, 32'hc29ff2d3, 32'hc10cdcd1};
test_output[1197] = '{32'h42915231};
test_index[1197] = '{3};
test_input[9584:9591] = '{32'hbfa21989, 32'h429a8402, 32'hc15b817d, 32'h4265fe44, 32'hc2c17ef6, 32'hc245db6e, 32'hc2c4326e, 32'h42062b17};
test_output[1198] = '{32'h429a8402};
test_index[1198] = '{1};
test_input[9592:9599] = '{32'hc2bd5fcb, 32'h404c3fa7, 32'hc21df160, 32'h41e9eb9c, 32'hc1bae23f, 32'hc2835d0d, 32'hc2065444, 32'hc1c7d9d8};
test_output[1199] = '{32'h41e9eb9c};
test_index[1199] = '{3};
test_input[9600:9607] = '{32'hc252a36e, 32'h4171e292, 32'h429c3f8e, 32'hc2bf31d7, 32'h422f5818, 32'h40b54483, 32'h42b508d3, 32'hc0c199d1};
test_output[1200] = '{32'h42b508d3};
test_index[1200] = '{6};
test_input[9608:9615] = '{32'hc23e0cfc, 32'hc2118b32, 32'h42aaa6ae, 32'hc20775b5, 32'hc16c7f86, 32'hc28ad712, 32'h4198fcd4, 32'hc1fb7972};
test_output[1201] = '{32'h42aaa6ae};
test_index[1201] = '{2};
test_input[9616:9623] = '{32'hc0ac72f5, 32'h427eced6, 32'hc279e249, 32'hc1cfefe9, 32'h3e8f48ae, 32'h400828cd, 32'hc231218f, 32'h428773dd};
test_output[1202] = '{32'h428773dd};
test_index[1202] = '{7};
test_input[9624:9631] = '{32'hc28047f1, 32'h4283827b, 32'hc188994f, 32'hc2b4a10c, 32'h42c1ae57, 32'hc2a06963, 32'h42271afd, 32'hc255935b};
test_output[1203] = '{32'h42c1ae57};
test_index[1203] = '{4};
test_input[9632:9639] = '{32'hc1be224e, 32'hc261da69, 32'h42176949, 32'h42528615, 32'hc2a2776a, 32'hc1982d97, 32'hc2952134, 32'h41bab46d};
test_output[1204] = '{32'h42528615};
test_index[1204] = '{3};
test_input[9640:9647] = '{32'h41b17bbe, 32'hc2b6e260, 32'hc1728a77, 32'hc128363c, 32'hc24cb0a2, 32'hc25218f0, 32'hc2726b1d, 32'hc2231ec5};
test_output[1205] = '{32'h41b17bbe};
test_index[1205] = '{0};
test_input[9648:9655] = '{32'hc22e4fba, 32'h42910140, 32'h42a668f5, 32'hc29ce419, 32'hc24e8ef3, 32'hc2920b68, 32'hc25c4d4d, 32'hc22f8a71};
test_output[1206] = '{32'h42a668f5};
test_index[1206] = '{2};
test_input[9656:9663] = '{32'h42891221, 32'h41b5292a, 32'h42390da3, 32'h42612c70, 32'hc29f904f, 32'h42059dfc, 32'h42bbf0fc, 32'hc23f6ebe};
test_output[1207] = '{32'h42bbf0fc};
test_index[1207] = '{6};
test_input[9664:9671] = '{32'hc21a9a63, 32'h401c98a6, 32'h42193f58, 32'h42bb0796, 32'h4287fba9, 32'h424003d7, 32'hc262e849, 32'h421620d9};
test_output[1208] = '{32'h42bb0796};
test_index[1208] = '{3};
test_input[9672:9679] = '{32'hc2748403, 32'h428e29e9, 32'h422cc6c8, 32'h4210a719, 32'hc29d6399, 32'hc2b645a0, 32'hc20bba3d, 32'h42c6b5e2};
test_output[1209] = '{32'h42c6b5e2};
test_index[1209] = '{7};
test_input[9680:9687] = '{32'hc0e1b44c, 32'hc2b36999, 32'h41ec5679, 32'hc00d6ed4, 32'hc2bf0660, 32'hc20b7e37, 32'hc2c1a212, 32'hc03f6dcc};
test_output[1210] = '{32'h41ec5679};
test_index[1210] = '{2};
test_input[9688:9695] = '{32'hc213b4ec, 32'h42c5bea7, 32'hc2345c2f, 32'hc1b4c498, 32'hc2526327, 32'h42306b73, 32'h428533b4, 32'hc10e0dc0};
test_output[1211] = '{32'h42c5bea7};
test_index[1211] = '{1};
test_input[9696:9703] = '{32'h41ba598b, 32'hc134c340, 32'hbfbc8e7b, 32'hc1b75d82, 32'h425b6b21, 32'hc22bf780, 32'hc28a7da2, 32'h4244cb24};
test_output[1212] = '{32'h425b6b21};
test_index[1212] = '{4};
test_input[9704:9711] = '{32'hc0350949, 32'h41f5999a, 32'h42af5c9f, 32'h42296a61, 32'h40bb6310, 32'h42b0dcd0, 32'hc2709a8e, 32'h422b61ca};
test_output[1213] = '{32'h42b0dcd0};
test_index[1213] = '{5};
test_input[9712:9719] = '{32'hc1671c9b, 32'h41bc5168, 32'h426245fa, 32'h425df786, 32'h4293cc3f, 32'h420d0db9, 32'h42a10cd0, 32'h4248dcbc};
test_output[1214] = '{32'h42a10cd0};
test_index[1214] = '{6};
test_input[9720:9727] = '{32'hc2098ffb, 32'hc2228304, 32'h42b9885a, 32'h428b1542, 32'hc2a08d9d, 32'hbf57e7c5, 32'h42a944f8, 32'h4168c4ed};
test_output[1215] = '{32'h42b9885a};
test_index[1215] = '{2};
test_input[9728:9735] = '{32'h41a1ade7, 32'h42aa9fc9, 32'hc2b85cbb, 32'hc233719f, 32'hc1ddcb9f, 32'h42c16564, 32'hc1bf6674, 32'h4251d9fb};
test_output[1216] = '{32'h42c16564};
test_index[1216] = '{5};
test_input[9736:9743] = '{32'hc1af38a6, 32'hc1bddb90, 32'h42a69036, 32'hc2315b59, 32'h42a926e3, 32'hc1748af7, 32'hc23e623a, 32'hc2951ae9};
test_output[1217] = '{32'h42a926e3};
test_index[1217] = '{4};
test_input[9744:9751] = '{32'h426d05db, 32'h42378a46, 32'h418b75a1, 32'h418f229b, 32'h42780ded, 32'hc29455ad, 32'h4261ded5, 32'h41a2b7f0};
test_output[1218] = '{32'h42780ded};
test_index[1218] = '{4};
test_input[9752:9759] = '{32'h41df086b, 32'hbf9fd956, 32'h42be05aa, 32'h4229e591, 32'hc266d29a, 32'hc2bafa06, 32'h42bbdef0, 32'h41a4ebde};
test_output[1219] = '{32'h42be05aa};
test_index[1219] = '{2};
test_input[9760:9767] = '{32'hc1756768, 32'h4286b784, 32'hc20426eb, 32'h4222fa95, 32'hc0028f22, 32'h418d41f0, 32'hc28fbfe9, 32'hc25b2723};
test_output[1220] = '{32'h4286b784};
test_index[1220] = '{1};
test_input[9768:9775] = '{32'hc2137b24, 32'hc26c3129, 32'hc260d025, 32'h41832a86, 32'h427e2041, 32'hc23d54c3, 32'h412276a5, 32'hc2be7acf};
test_output[1221] = '{32'h427e2041};
test_index[1221] = '{4};
test_input[9776:9783] = '{32'h425d516f, 32'h42711222, 32'h42760ef3, 32'hc10c77e0, 32'h42a2d2a5, 32'h41a5c215, 32'hc2b07b7a, 32'h423edded};
test_output[1222] = '{32'h42a2d2a5};
test_index[1222] = '{4};
test_input[9784:9791] = '{32'h425f33e6, 32'hc221fca4, 32'hbfa04c59, 32'hc239c29f, 32'h40b91e5d, 32'hbfe6a429, 32'hc29b2890, 32'h42703f93};
test_output[1223] = '{32'h42703f93};
test_index[1223] = '{7};
test_input[9792:9799] = '{32'hc1fc19e1, 32'h410d2e39, 32'h41d81316, 32'h424a8ab9, 32'hc1850437, 32'hc2b84275, 32'hc1bb9c6b, 32'hc2ae525a};
test_output[1224] = '{32'h424a8ab9};
test_index[1224] = '{3};
test_input[9800:9807] = '{32'hc2891488, 32'hc2c6781e, 32'h4280f215, 32'hc24de157, 32'hc221eb21, 32'h42ab4b07, 32'hc2c218d8, 32'hc1845366};
test_output[1225] = '{32'h42ab4b07};
test_index[1225] = '{5};
test_input[9808:9815] = '{32'hc2162793, 32'hc202b432, 32'h4255c0a3, 32'h4275fd40, 32'hc23d8882, 32'hc2a48516, 32'hc2b7f0b3, 32'h42960b4c};
test_output[1226] = '{32'h42960b4c};
test_index[1226] = '{7};
test_input[9816:9823] = '{32'hc24cc374, 32'h421fab97, 32'hc269636c, 32'h41932785, 32'hc2b7834a, 32'h420c483a, 32'h41d82193, 32'hc2b6b1c9};
test_output[1227] = '{32'h421fab97};
test_index[1227] = '{1};
test_input[9824:9831] = '{32'h418ca5c5, 32'hc2a860ff, 32'hc2148afa, 32'hc1838dc6, 32'h423ac4d9, 32'hc2af413d, 32'h42854de8, 32'hc2b397db};
test_output[1228] = '{32'h42854de8};
test_index[1228] = '{6};
test_input[9832:9839] = '{32'h4189465e, 32'hc2b1c12e, 32'h427da73c, 32'hc26e6bea, 32'h41afed5b, 32'h42182010, 32'hc28c4bbd, 32'h42bd6e80};
test_output[1229] = '{32'h42bd6e80};
test_index[1229] = '{7};
test_input[9840:9847] = '{32'h42113487, 32'h42390b13, 32'hc0b1c055, 32'hc2aa9277, 32'h4200e793, 32'hc12b795d, 32'hc2c30cc7, 32'hc2aba93d};
test_output[1230] = '{32'h42390b13};
test_index[1230] = '{1};
test_input[9848:9855] = '{32'h3fd88dfe, 32'hc245f6a9, 32'hc227524d, 32'hc2619f9c, 32'h429fdd1c, 32'hc1514eaf, 32'hc2044a7e, 32'h4291947c};
test_output[1231] = '{32'h429fdd1c};
test_index[1231] = '{4};
test_input[9856:9863] = '{32'hc2b90d56, 32'h416ff5ac, 32'h421f3071, 32'hc15a07ab, 32'hc2aa1448, 32'h42bed300, 32'h41fbfb50, 32'h41f5d6ca};
test_output[1232] = '{32'h42bed300};
test_index[1232] = '{5};
test_input[9864:9871] = '{32'h41ad4cb1, 32'h42a38881, 32'h423fba05, 32'h429aead7, 32'h42b6add0, 32'h42b116e6, 32'hc2a4a730, 32'hc115e352};
test_output[1233] = '{32'h42b6add0};
test_index[1233] = '{4};
test_input[9872:9879] = '{32'hc27bc99c, 32'hc227383f, 32'h422a3810, 32'h4219ade3, 32'h4204e4c4, 32'h41aed38d, 32'h423a8b02, 32'h42299eed};
test_output[1234] = '{32'h423a8b02};
test_index[1234] = '{6};
test_input[9880:9887] = '{32'hc21ac5d9, 32'hc299f343, 32'hc1cc5c3f, 32'hc25b1ebe, 32'hc219a861, 32'h42565873, 32'h4098b62a, 32'h41aaccc6};
test_output[1235] = '{32'h42565873};
test_index[1235] = '{5};
test_input[9888:9895] = '{32'h4087a165, 32'h42b15674, 32'hc219f9c2, 32'hc1c39575, 32'h4167ae75, 32'h409c7ed2, 32'hbd936487, 32'h42963e82};
test_output[1236] = '{32'h42b15674};
test_index[1236] = '{1};
test_input[9896:9903] = '{32'hc224cf98, 32'h42a388cf, 32'h424c99e2, 32'hc2a2fb2f, 32'h4178be17, 32'h4292ce23, 32'hc1c98b37, 32'h4182cdd8};
test_output[1237] = '{32'h42a388cf};
test_index[1237] = '{1};
test_input[9904:9911] = '{32'hc2688bde, 32'hc1d1887b, 32'h42880524, 32'h411c30f2, 32'h42687f72, 32'h429cb768, 32'hc2163b3f, 32'hbfe2803e};
test_output[1238] = '{32'h429cb768};
test_index[1238] = '{5};
test_input[9912:9919] = '{32'hc1c4143c, 32'hc18bcf6b, 32'h41cdce92, 32'hc2476e0b, 32'hc26ef4c4, 32'h42ab7f1f, 32'h42c1754c, 32'h4218c7a1};
test_output[1239] = '{32'h42c1754c};
test_index[1239] = '{6};
test_input[9920:9927] = '{32'hc0952d1d, 32'h420cfa52, 32'hc1d2d390, 32'h424cc245, 32'hc294c653, 32'h421a2941, 32'hc246ca93, 32'hc21b5594};
test_output[1240] = '{32'h424cc245};
test_index[1240] = '{3};
test_input[9928:9935] = '{32'h427797c9, 32'h41c77cdb, 32'h428281eb, 32'h42b706b3, 32'hc282e7ca, 32'hc08b95b9, 32'h420dceb4, 32'h42bceebb};
test_output[1241] = '{32'h42bceebb};
test_index[1241] = '{7};
test_input[9936:9943] = '{32'hc184c4a5, 32'h4190e690, 32'hc24058e0, 32'hc226ba4b, 32'hc28d8a7f, 32'hc296f1ff, 32'hc2a09e4d, 32'h4242dd03};
test_output[1242] = '{32'h4242dd03};
test_index[1242] = '{7};
test_input[9944:9951] = '{32'hc2c6b182, 32'h42987ff0, 32'hc29f0fa2, 32'hc2a1264a, 32'h42641afa, 32'h42805998, 32'h40077da4, 32'h42638b5e};
test_output[1243] = '{32'h42987ff0};
test_index[1243] = '{1};
test_input[9952:9959] = '{32'h42c5106f, 32'hc1c25144, 32'hc127f7e9, 32'h421892e3, 32'hc26a273d, 32'h42bcda7a, 32'hc2a64c90, 32'h4298d732};
test_output[1244] = '{32'h42c5106f};
test_index[1244] = '{0};
test_input[9960:9967] = '{32'hc2a44bf8, 32'hc0753e2c, 32'hc278ce7c, 32'h42991b0a, 32'hc19a7863, 32'h42a6fc04, 32'h413ffc42, 32'hc2479227};
test_output[1245] = '{32'h42a6fc04};
test_index[1245] = '{5};
test_input[9968:9975] = '{32'h42c3218f, 32'hc15679f6, 32'h4287cc8b, 32'h42c50284, 32'hc281fddf, 32'hc2bf5ba5, 32'hc2b5551f, 32'h426c7052};
test_output[1246] = '{32'h42c50284};
test_index[1246] = '{3};
test_input[9976:9983] = '{32'h4137edc4, 32'h4248407f, 32'h4179de58, 32'hc1142f02, 32'hc214b14a, 32'hc29e7425, 32'hc2a40dcf, 32'hc2587522};
test_output[1247] = '{32'h4248407f};
test_index[1247] = '{1};
test_input[9984:9991] = '{32'hc0cad734, 32'h42673a7a, 32'hc1be059c, 32'h429c48a4, 32'h41b608ef, 32'hc286c2db, 32'hc053fd0c, 32'h42a5414a};
test_output[1248] = '{32'h42a5414a};
test_index[1248] = '{7};
test_input[9992:9999] = '{32'h4114e883, 32'hc28872e1, 32'h4178f933, 32'hc283a965, 32'h40520f5d, 32'hc0ff025c, 32'h422ceebf, 32'hc2850a31};
test_output[1249] = '{32'h422ceebf};
test_index[1249] = '{6};
test_input[10000:10007] = '{32'h421a0f1f, 32'h423a347f, 32'hc0aad89e, 32'hc23b402f, 32'h42a00b9c, 32'h424f5d46, 32'hc2c741ec, 32'hc141901b};
test_output[1250] = '{32'h42a00b9c};
test_index[1250] = '{4};
test_input[10008:10015] = '{32'h40e185c7, 32'hc2b14748, 32'h42942195, 32'hc181fab1, 32'hc2499d7e, 32'h42218393, 32'h4192c610, 32'hc18280e2};
test_output[1251] = '{32'h42942195};
test_index[1251] = '{2};
test_input[10016:10023] = '{32'hc28d1ff1, 32'hc1b36a4f, 32'h42696b37, 32'h42396076, 32'hc25340b4, 32'h429df8a3, 32'hc2b19c6c, 32'h42be9bb0};
test_output[1252] = '{32'h42be9bb0};
test_index[1252] = '{7};
test_input[10024:10031] = '{32'h41c5b2ee, 32'h40c0b4c8, 32'hc2a36207, 32'h413a27c3, 32'h42b3dd5b, 32'hc10e0adc, 32'hbfd761e5, 32'hc1d5c5cb};
test_output[1253] = '{32'h42b3dd5b};
test_index[1253] = '{4};
test_input[10032:10039] = '{32'hc244f27b, 32'h418d89bc, 32'h4216eac6, 32'h4257b374, 32'hc251174c, 32'hc2be204a, 32'h41187dcd, 32'hc0484d23};
test_output[1254] = '{32'h4257b374};
test_index[1254] = '{3};
test_input[10040:10047] = '{32'hc2a53906, 32'hc24814a3, 32'hc28f7e34, 32'h421fb5c4, 32'hc153a244, 32'hc25fdad3, 32'h42bed00c, 32'hc22c93b9};
test_output[1255] = '{32'h42bed00c};
test_index[1255] = '{6};
test_input[10048:10055] = '{32'hc1b3d6ff, 32'hc051cd00, 32'hc22eb8a8, 32'hc0d17c9d, 32'h426fce80, 32'h41dbca1b, 32'hc276741a, 32'h40d3b4b4};
test_output[1256] = '{32'h426fce80};
test_index[1256] = '{4};
test_input[10056:10063] = '{32'hc18b16fb, 32'hc20bafe2, 32'hc1dc7192, 32'hc2942f5a, 32'h414f6fc4, 32'h42bbbe4a, 32'h42b605cd, 32'hc1c14f29};
test_output[1257] = '{32'h42bbbe4a};
test_index[1257] = '{5};
test_input[10064:10071] = '{32'h42b9a6e5, 32'hc284e79e, 32'h42990b91, 32'h41c0c604, 32'h4266e331, 32'h4257073d, 32'hc1a5493d, 32'hc227a3e5};
test_output[1258] = '{32'h42b9a6e5};
test_index[1258] = '{0};
test_input[10072:10079] = '{32'hc2b1a74a, 32'hc2bfbdd6, 32'h429e4c88, 32'h41de163d, 32'h41eb05aa, 32'h420534a8, 32'hc1cf0e51, 32'h41647cf8};
test_output[1259] = '{32'h429e4c88};
test_index[1259] = '{2};
test_input[10080:10087] = '{32'h42800acf, 32'hc20ab061, 32'h410ef77f, 32'hc2b70df5, 32'h42c6a229, 32'hc1e3d0f1, 32'hc29dd5d3, 32'h429cf090};
test_output[1260] = '{32'h42c6a229};
test_index[1260] = '{4};
test_input[10088:10095] = '{32'h41ffff65, 32'h42a85d45, 32'hc276c94e, 32'hc29ffdb0, 32'h42828cdf, 32'hc24dc574, 32'hc250dea5, 32'h42708a63};
test_output[1261] = '{32'h42a85d45};
test_index[1261] = '{1};
test_input[10096:10103] = '{32'h4123ef1c, 32'hc115e731, 32'hc251b341, 32'h4283ef6a, 32'hc2394d41, 32'h420ace24, 32'h42ad5749, 32'h41dcd1c3};
test_output[1262] = '{32'h42ad5749};
test_index[1262] = '{6};
test_input[10104:10111] = '{32'hc10237ba, 32'hc1dd66de, 32'hc20e3823, 32'hc19dd6da, 32'hc270eaf3, 32'h41811114, 32'hc2085f74, 32'hc28bf4fb};
test_output[1263] = '{32'h41811114};
test_index[1263] = '{5};
test_input[10112:10119] = '{32'h41d2151f, 32'hc24745c4, 32'h416a0818, 32'h420187c4, 32'h4193482b, 32'h428f4460, 32'hc1629524, 32'h41d6d0b7};
test_output[1264] = '{32'h428f4460};
test_index[1264] = '{5};
test_input[10120:10127] = '{32'h41a57a5c, 32'h422a57cf, 32'h40edc1f2, 32'h40eee512, 32'hc1b7ea0c, 32'h41ee1408, 32'h4215ba53, 32'h42390a18};
test_output[1265] = '{32'h42390a18};
test_index[1265] = '{7};
test_input[10128:10135] = '{32'hc1f19f4f, 32'hc1993554, 32'hc22e1b7b, 32'hc2b4c107, 32'h423e65a1, 32'h42977616, 32'hc126f397, 32'hc2677fd8};
test_output[1266] = '{32'h42977616};
test_index[1266] = '{5};
test_input[10136:10143] = '{32'h405fd562, 32'h429f6f88, 32'hc2617030, 32'h4224610d, 32'h41a3ce34, 32'h4292e21f, 32'hc1849c38, 32'h429f0caf};
test_output[1267] = '{32'h429f6f88};
test_index[1267] = '{1};
test_input[10144:10151] = '{32'h41992fe6, 32'h42a7641f, 32'hc2b2c15b, 32'hc29b4d2c, 32'hc0ead935, 32'hc2beb66d, 32'hc129266e, 32'h42987861};
test_output[1268] = '{32'h42a7641f};
test_index[1268] = '{1};
test_input[10152:10159] = '{32'h417f8cb5, 32'h42375274, 32'hc228c618, 32'h423dfcc8, 32'h42c6ae93, 32'h423fd16d, 32'h41b3ef27, 32'hc2c598ce};
test_output[1269] = '{32'h42c6ae93};
test_index[1269] = '{4};
test_input[10160:10167] = '{32'hbb6152ad, 32'hc23d58f3, 32'hc1f9381f, 32'hc1c65c9e, 32'hc28086ee, 32'h42b0d143, 32'hc284322b, 32'hc2a20f12};
test_output[1270] = '{32'h42b0d143};
test_index[1270] = '{5};
test_input[10168:10175] = '{32'h426ed38f, 32'hc24a7c8f, 32'hc107773f, 32'h42be7a04, 32'hc248b577, 32'hc007cf0c, 32'hc227dccd, 32'h41b7300c};
test_output[1271] = '{32'h42be7a04};
test_index[1271] = '{3};
test_input[10176:10183] = '{32'hc2242995, 32'hc212b17e, 32'hc18ea8cb, 32'hc285881b, 32'hc2c76880, 32'h42269fa2, 32'h4181f5c6, 32'h42892248};
test_output[1272] = '{32'h42892248};
test_index[1272] = '{7};
test_input[10184:10191] = '{32'h40998db9, 32'h42c71ae0, 32'hc1d837f4, 32'hc2a2d323, 32'h40f0d44e, 32'h42932f88, 32'h42b5ab9b, 32'h42402f84};
test_output[1273] = '{32'h42c71ae0};
test_index[1273] = '{1};
test_input[10192:10199] = '{32'hc2b828d5, 32'h4169b0b4, 32'h41df911e, 32'hc29bbd90, 32'hc260109c, 32'hc168f4ed, 32'h3fc76802, 32'hc20611a6};
test_output[1274] = '{32'h41df911e};
test_index[1274] = '{2};
test_input[10200:10207] = '{32'hc20509d6, 32'hc2b530c1, 32'hc2984cd9, 32'hc1612d8d, 32'hc1c3116d, 32'hc1ea4f60, 32'hc2c4c665, 32'h41e2802c};
test_output[1275] = '{32'h41e2802c};
test_index[1275] = '{7};
test_input[10208:10215] = '{32'h429fe9d4, 32'hc24c2bbb, 32'h423409b5, 32'h42af1767, 32'h42af6bdf, 32'h4289b7e1, 32'h42a0b06d, 32'hc1d3a0c2};
test_output[1276] = '{32'h42af6bdf};
test_index[1276] = '{4};
test_input[10216:10223] = '{32'h42c36420, 32'hc155e6cf, 32'hc21ac7f5, 32'h424777d4, 32'h42a59191, 32'hc2a91d77, 32'h4292e170, 32'h4154bb50};
test_output[1277] = '{32'h42c36420};
test_index[1277] = '{0};
test_input[10224:10231] = '{32'h42bc15d2, 32'h4251899e, 32'hc28c66b4, 32'h42775246, 32'h42075d04, 32'h42be30b8, 32'h4201a1db, 32'h4268b814};
test_output[1278] = '{32'h42be30b8};
test_index[1278] = '{5};
test_input[10232:10239] = '{32'hc281cb87, 32'hc2a6bf2f, 32'h42453b18, 32'hc2511034, 32'h429ab1ab, 32'h42a23978, 32'hc11bc3a5, 32'hc2ab7f86};
test_output[1279] = '{32'h42a23978};
test_index[1279] = '{5};
test_input[10240:10247] = '{32'hc055e290, 32'hc13b2a77, 32'hc285dd92, 32'h426053af, 32'h417f172f, 32'hc2288c64, 32'hc2c5ca43, 32'hc2c30658};
test_output[1280] = '{32'h426053af};
test_index[1280] = '{3};
test_input[10248:10255] = '{32'h42881ed3, 32'hc2bc1dc9, 32'h425d7f32, 32'h42078aa7, 32'hc1e17a70, 32'h42b9e8c7, 32'hc23a9c30, 32'hc23dcfb8};
test_output[1281] = '{32'h42b9e8c7};
test_index[1281] = '{5};
test_input[10256:10263] = '{32'hc2aff29d, 32'h4260e2a9, 32'hc2c6b705, 32'hc21716b6, 32'h3fdbbff1, 32'hc286b42b, 32'hc26c9def, 32'hc136834f};
test_output[1282] = '{32'h4260e2a9};
test_index[1282] = '{1};
test_input[10264:10271] = '{32'h4211537e, 32'h42ac5722, 32'h42244953, 32'hc1e6f98c, 32'hc145237d, 32'hc2c4b15d, 32'hc287bb7a, 32'h42979660};
test_output[1283] = '{32'h42ac5722};
test_index[1283] = '{1};
test_input[10272:10279] = '{32'h42864458, 32'hc28ef95d, 32'h42bddd59, 32'hc1841864, 32'h428f88e1, 32'h42b9aa8e, 32'hc1eed233, 32'hc1443b6f};
test_output[1284] = '{32'h42bddd59};
test_index[1284] = '{2};
test_input[10280:10287] = '{32'h42916cb0, 32'hc1d2915e, 32'h41c577a7, 32'hc253cb91, 32'hc2c48885, 32'hc16561f0, 32'h4290110e, 32'hc21cf1ea};
test_output[1285] = '{32'h42916cb0};
test_index[1285] = '{0};
test_input[10288:10295] = '{32'h40157f7c, 32'h41c81614, 32'hc20a9639, 32'h429725a3, 32'hc26ad420, 32'h42ad33f4, 32'h42a4b701, 32'hc21382dd};
test_output[1286] = '{32'h42ad33f4};
test_index[1286] = '{5};
test_input[10296:10303] = '{32'hc0913293, 32'h4205bdf0, 32'hc2103786, 32'h4297139c, 32'h3f7e53ff, 32'hc247d7b7, 32'h418fa8e7, 32'h426faaa2};
test_output[1287] = '{32'h4297139c};
test_index[1287] = '{3};
test_input[10304:10311] = '{32'hc2b07872, 32'hc0cf8049, 32'h42c26883, 32'hc28d7581, 32'hc29cccb0, 32'hc2c6e6b7, 32'hc1037060, 32'hc252dceb};
test_output[1288] = '{32'h42c26883};
test_index[1288] = '{2};
test_input[10312:10319] = '{32'h42c2b493, 32'h42a135b8, 32'hc21b1bd7, 32'h41f6bef1, 32'hc261b591, 32'h411f2e5e, 32'h424e12cb, 32'hc2c02685};
test_output[1289] = '{32'h42c2b493};
test_index[1289] = '{0};
test_input[10320:10327] = '{32'h415491b7, 32'h42983e64, 32'h42136123, 32'h41c83dda, 32'hc288bd9d, 32'hc294f36d, 32'h420a37ab, 32'h40af5748};
test_output[1290] = '{32'h42983e64};
test_index[1290] = '{1};
test_input[10328:10335] = '{32'h4263b924, 32'h42934577, 32'hc285d77d, 32'h40fe2cba, 32'h42272c36, 32'hc1d87238, 32'h4223dc19, 32'h42b7e49a};
test_output[1291] = '{32'h42b7e49a};
test_index[1291] = '{7};
test_input[10336:10343] = '{32'hc2841dcc, 32'h42a7c6be, 32'h42b035c1, 32'h42781ea1, 32'h41e77c30, 32'h42aecb8f, 32'hc28768dc, 32'hc1229f96};
test_output[1292] = '{32'h42b035c1};
test_index[1292] = '{2};
test_input[10344:10351] = '{32'h41561c24, 32'hc2706109, 32'hc11cef8d, 32'hc28032ea, 32'h428be1e1, 32'h428b3a06, 32'hc2bc569d, 32'hc2c4f0ca};
test_output[1293] = '{32'h428be1e1};
test_index[1293] = '{4};
test_input[10352:10359] = '{32'hc2006f54, 32'h4226b927, 32'h42a8188e, 32'hc1f98627, 32'h412ed3f7, 32'hc2292d88, 32'hc1d96c4d, 32'hc1c9b9b1};
test_output[1294] = '{32'h42a8188e};
test_index[1294] = '{2};
test_input[10360:10367] = '{32'hc2a748d0, 32'hc1c88ed9, 32'hc2aba1a7, 32'hc2bd0b83, 32'h41cfc282, 32'hc0fa6447, 32'h42bebcea, 32'hc2838a68};
test_output[1295] = '{32'h42bebcea};
test_index[1295] = '{6};
test_input[10368:10375] = '{32'hc2518dc4, 32'hc2865c64, 32'hc2c0bc5f, 32'hc2baaa35, 32'hbfc06fe3, 32'hc221cca9, 32'h42729093, 32'hc0f03691};
test_output[1296] = '{32'h42729093};
test_index[1296] = '{6};
test_input[10376:10383] = '{32'hc212dd87, 32'hc1d6f6c8, 32'hc048297a, 32'hbf4e3a76, 32'hc22403b3, 32'hc24cfb15, 32'hc0c36971, 32'hc2ab649a};
test_output[1297] = '{32'hbf4e3a76};
test_index[1297] = '{3};
test_input[10384:10391] = '{32'h42aa894c, 32'h42387081, 32'h42485d3a, 32'h421a30c9, 32'hc2a7e6b9, 32'h425a2a0e, 32'hc2b62d34, 32'h41fdd028};
test_output[1298] = '{32'h42aa894c};
test_index[1298] = '{0};
test_input[10392:10399] = '{32'hc23defab, 32'h3f52bca7, 32'h41dce175, 32'hc281dc16, 32'hc2a33f09, 32'h4251f0c6, 32'hc2a5e731, 32'h42596f60};
test_output[1299] = '{32'h42596f60};
test_index[1299] = '{7};
test_input[10400:10407] = '{32'hc16ed713, 32'h42944594, 32'hc2ae3553, 32'hc27d7530, 32'h42859fd0, 32'h42bf737b, 32'hc2b41e7a, 32'h420915a2};
test_output[1300] = '{32'h42bf737b};
test_index[1300] = '{5};
test_input[10408:10415] = '{32'hc28bdd22, 32'h423230b8, 32'hc10c25dd, 32'hc0e41bc3, 32'h4293a139, 32'h425b10fa, 32'h41e8e746, 32'hc26f9deb};
test_output[1301] = '{32'h4293a139};
test_index[1301] = '{4};
test_input[10416:10423] = '{32'h413807b2, 32'hc2449c2d, 32'h429fa53b, 32'hc228872a, 32'hc2b1e97b, 32'hc091e79a, 32'hc0bca7bf, 32'hc22d3195};
test_output[1302] = '{32'h429fa53b};
test_index[1302] = '{2};
test_input[10424:10431] = '{32'hc295689c, 32'h42ae6a9f, 32'h42827c94, 32'h42876fbe, 32'hc1012715, 32'hc194f71a, 32'h420dd271, 32'hc139eeec};
test_output[1303] = '{32'h42ae6a9f};
test_index[1303] = '{1};
test_input[10432:10439] = '{32'hc15113d6, 32'hc2b4405a, 32'hc2b6fe77, 32'h421f4547, 32'h40aaeaa2, 32'h42c4cd19, 32'h425a8f6c, 32'hc1d515c5};
test_output[1304] = '{32'h42c4cd19};
test_index[1304] = '{5};
test_input[10440:10447] = '{32'h40508cbf, 32'h4109219e, 32'hc1a1e897, 32'h42bb1bed, 32'h41bcac66, 32'hc29a98f5, 32'hc28217d8, 32'hc268bc1e};
test_output[1305] = '{32'h42bb1bed};
test_index[1305] = '{3};
test_input[10448:10455] = '{32'h41c49f94, 32'hc1cc78c6, 32'h4125fc12, 32'hc2687206, 32'h4209b2e5, 32'h41ef5ddf, 32'hc2c22f14, 32'hc08adf9b};
test_output[1306] = '{32'h4209b2e5};
test_index[1306] = '{4};
test_input[10456:10463] = '{32'hc080f46b, 32'hc299223f, 32'h417e0070, 32'h42148b25, 32'h4217e951, 32'h4280b15d, 32'hc2b2a19c, 32'hc11197e9};
test_output[1307] = '{32'h4280b15d};
test_index[1307] = '{5};
test_input[10464:10471] = '{32'h4193baa2, 32'h401ffe02, 32'h423747e2, 32'hc26df0e8, 32'hc273dbf5, 32'hc245a36f, 32'h42685174, 32'hc2a984a3};
test_output[1308] = '{32'h42685174};
test_index[1308] = '{6};
test_input[10472:10479] = '{32'h41eb803e, 32'h40df8e60, 32'h4287dd89, 32'hbf0051d1, 32'h4293a320, 32'h42a8ab23, 32'hc1da0581, 32'hc29183b5};
test_output[1309] = '{32'h42a8ab23};
test_index[1309] = '{5};
test_input[10480:10487] = '{32'h429de9bc, 32'hc2a8c047, 32'hc2836d4b, 32'h42c3ef29, 32'h41b424c6, 32'hc2088cbc, 32'h41694823, 32'h41979d27};
test_output[1310] = '{32'h42c3ef29};
test_index[1310] = '{3};
test_input[10488:10495] = '{32'hc2107883, 32'h42816a4d, 32'hc150f7e1, 32'h4294344a, 32'h41be3ea8, 32'h40bd9536, 32'hc1f6e58a, 32'h420f3052};
test_output[1311] = '{32'h4294344a};
test_index[1311] = '{3};
test_input[10496:10503] = '{32'h42583ccf, 32'hc24bafac, 32'h423f316b, 32'hc254796d, 32'hc2178501, 32'h424f76f0, 32'hc18093a7, 32'h423a9d6f};
test_output[1312] = '{32'h42583ccf};
test_index[1312] = '{0};
test_input[10504:10511] = '{32'h42896df7, 32'h422a9342, 32'h41ae4a07, 32'h4285072c, 32'h42c07a04, 32'h42b7cf0c, 32'hc2445659, 32'h4293e739};
test_output[1313] = '{32'h42c07a04};
test_index[1313] = '{4};
test_input[10512:10519] = '{32'hc18e5a45, 32'hc1536c8f, 32'hc1d9610b, 32'hc2acecf2, 32'hc2161341, 32'hc29f296e, 32'h42a913f1, 32'h42c1a2d8};
test_output[1314] = '{32'h42c1a2d8};
test_index[1314] = '{7};
test_input[10520:10527] = '{32'h404b892d, 32'h42c3ef08, 32'hc29b5365, 32'hc28f8a9f, 32'h40eea73b, 32'h42b43884, 32'h41a0299f, 32'hc1822935};
test_output[1315] = '{32'h42c3ef08};
test_index[1315] = '{1};
test_input[10528:10535] = '{32'h411a2ba5, 32'h42a358a9, 32'hc2a05f33, 32'hc21966eb, 32'hc1df71ad, 32'hc1f85f92, 32'h429af639, 32'hc2be3b81};
test_output[1316] = '{32'h42a358a9};
test_index[1316] = '{1};
test_input[10536:10543] = '{32'h41ff1821, 32'h42b9fb96, 32'h42271339, 32'hc192c6ab, 32'h427495c6, 32'h4108a921, 32'hc2269599, 32'hc26a8274};
test_output[1317] = '{32'h42b9fb96};
test_index[1317] = '{1};
test_input[10544:10551] = '{32'hc2829862, 32'h424a27fd, 32'h42bc669c, 32'h42acb42b, 32'hc283ce8c, 32'h42227c32, 32'h429c84fd, 32'hc2a4c5e3};
test_output[1318] = '{32'h42bc669c};
test_index[1318] = '{2};
test_input[10552:10559] = '{32'hc290e965, 32'h42b425c2, 32'hc27ef3f3, 32'hc25b682b, 32'hc25e6a94, 32'h425d56b2, 32'hc2ab443e, 32'h428d27c4};
test_output[1319] = '{32'h42b425c2};
test_index[1319] = '{1};
test_input[10560:10567] = '{32'h42b5e6be, 32'h4225a412, 32'hc19c877c, 32'h410042aa, 32'h41a5fd8a, 32'hc1e77006, 32'hc286c947, 32'h42846ea1};
test_output[1320] = '{32'h42b5e6be};
test_index[1320] = '{0};
test_input[10568:10575] = '{32'hc22cdef5, 32'h428b3fd1, 32'hc2c4e197, 32'h4184e3d4, 32'h42c4e1d6, 32'h4299a272, 32'hc08dc060, 32'hc26ca5ba};
test_output[1321] = '{32'h42c4e1d6};
test_index[1321] = '{4};
test_input[10576:10583] = '{32'h426ae13a, 32'h425f1960, 32'hc0943e93, 32'hc222db51, 32'hc2658bab, 32'hc2b45d59, 32'h4291564c, 32'h41d3d64f};
test_output[1322] = '{32'h4291564c};
test_index[1322] = '{6};
test_input[10584:10591] = '{32'hc2a9287b, 32'h4276a8da, 32'h4146d19b, 32'hc2095615, 32'h42799a12, 32'hc2a3a622, 32'hc245a25e, 32'hc246b2bc};
test_output[1323] = '{32'h42799a12};
test_index[1323] = '{4};
test_input[10592:10599] = '{32'h42c56204, 32'h429db3a1, 32'hc01b17fc, 32'h42c4af77, 32'hc2c131e7, 32'h42ab9b64, 32'h428ea38d, 32'h40bf1d67};
test_output[1324] = '{32'h42c56204};
test_index[1324] = '{0};
test_input[10600:10607] = '{32'hc28e8f43, 32'h42b3bcce, 32'h421bcf05, 32'h42b7de44, 32'h428c5e21, 32'hc2b8a787, 32'h4244a57d, 32'hc11d3ec2};
test_output[1325] = '{32'h42b7de44};
test_index[1325] = '{3};
test_input[10608:10615] = '{32'hc1a03976, 32'hc1c09716, 32'hc2629386, 32'hc2bf7450, 32'h41d1bb81, 32'hc2378b2b, 32'hc2aa1778, 32'hc202c418};
test_output[1326] = '{32'h41d1bb81};
test_index[1326] = '{4};
test_input[10616:10623] = '{32'hc2033cfc, 32'h42a512dc, 32'hc1fb1942, 32'hc25bbd1c, 32'h422e27e0, 32'h41af7f8e, 32'hc2908552, 32'h4110680b};
test_output[1327] = '{32'h42a512dc};
test_index[1327] = '{1};
test_input[10624:10631] = '{32'h42829a38, 32'h40fc7667, 32'h41c2db55, 32'h40c33d53, 32'h41831fb0, 32'h4113b633, 32'hc2c4fd30, 32'hc2afd0b0};
test_output[1328] = '{32'h42829a38};
test_index[1328] = '{0};
test_input[10632:10639] = '{32'hc224d3d7, 32'h410d8834, 32'h42bb129a, 32'h41b39980, 32'hc299ef19, 32'hc1157d3d, 32'h42b2aa93, 32'hc0d22b41};
test_output[1329] = '{32'h42bb129a};
test_index[1329] = '{2};
test_input[10640:10647] = '{32'h42882429, 32'h42aaa923, 32'hc2b775f1, 32'hc26bb863, 32'hc21149f2, 32'hc11276d5, 32'h4287b83b, 32'hc2622cc3};
test_output[1330] = '{32'h42aaa923};
test_index[1330] = '{1};
test_input[10648:10655] = '{32'h42b239ef, 32'hc2929cf7, 32'h42151d9a, 32'h41c8b607, 32'h427f9861, 32'hc29ebaeb, 32'hc20b63d6, 32'h40944ae8};
test_output[1331] = '{32'h42b239ef};
test_index[1331] = '{0};
test_input[10656:10663] = '{32'hc28c15d2, 32'h424521f9, 32'hc2b905ea, 32'hc2a6f361, 32'h411b05c3, 32'h41a2b1bb, 32'hc138395a, 32'hc2290b2e};
test_output[1332] = '{32'h424521f9};
test_index[1332] = '{1};
test_input[10664:10671] = '{32'hc29db9aa, 32'hc293d1bc, 32'h42c7eeb5, 32'h41a737c4, 32'hc16b95f7, 32'hc2c605a9, 32'hc216462b, 32'hc2855782};
test_output[1333] = '{32'h42c7eeb5};
test_index[1333] = '{2};
test_input[10672:10679] = '{32'h4294eff4, 32'hc2aa6e46, 32'h429cf4fd, 32'hc2bb9faa, 32'h42708658, 32'hc2557538, 32'hc0f4ee20, 32'h42b18354};
test_output[1334] = '{32'h42b18354};
test_index[1334] = '{7};
test_input[10680:10687] = '{32'hc2bdff84, 32'hc2610b7a, 32'h41fa3416, 32'hbfe28fb7, 32'hc275127f, 32'h425995a3, 32'hc2a4706b, 32'hc1df0036};
test_output[1335] = '{32'h425995a3};
test_index[1335] = '{5};
test_input[10688:10695] = '{32'hc2b2beeb, 32'hc24fe642, 32'hc1f6ced3, 32'h4282b331, 32'h4292c0f7, 32'hc1153fd4, 32'hc267cb4a, 32'hc085d43e};
test_output[1336] = '{32'h4292c0f7};
test_index[1336] = '{4};
test_input[10696:10703] = '{32'h42b0cbcf, 32'h415f2e11, 32'h4227ca54, 32'hc1ba1c98, 32'h42c4c054, 32'h42c3f686, 32'hc2c59dcd, 32'h4282c018};
test_output[1337] = '{32'h42c4c054};
test_index[1337] = '{4};
test_input[10704:10711] = '{32'h428d1dd0, 32'h42a29e9f, 32'h40b0e35d, 32'hc27accab, 32'hc287dbc9, 32'h419c8c3e, 32'hc288eb6e, 32'hc1bc8706};
test_output[1338] = '{32'h42a29e9f};
test_index[1338] = '{1};
test_input[10712:10719] = '{32'hc18301b4, 32'h42b56351, 32'h4255f34c, 32'h42879178, 32'h4224eb41, 32'hc0a31a9b, 32'hc20d5be3, 32'h415cfdb0};
test_output[1339] = '{32'h42b56351};
test_index[1339] = '{1};
test_input[10720:10727] = '{32'hc242e717, 32'h41e032e0, 32'h41f8c916, 32'h42a54f64, 32'hc1878e0d, 32'hc09096b1, 32'hc20c2a1f, 32'hc2837f80};
test_output[1340] = '{32'h42a54f64};
test_index[1340] = '{3};
test_input[10728:10735] = '{32'h42254f09, 32'hc0ebb39f, 32'h418ddd61, 32'hc2b7ff59, 32'h4222bcef, 32'h42aa8566, 32'h4225e5aa, 32'hc1d96abd};
test_output[1341] = '{32'h42aa8566};
test_index[1341] = '{5};
test_input[10736:10743] = '{32'h41fb6769, 32'h426ddd3b, 32'h41e54847, 32'h428f158b, 32'h429be916, 32'hc2a63963, 32'h426393d8, 32'hc1bc0ece};
test_output[1342] = '{32'h429be916};
test_index[1342] = '{4};
test_input[10744:10751] = '{32'h425f1032, 32'h429894a0, 32'h420f28bc, 32'h3fe66fdf, 32'h42aeb91b, 32'h41de6972, 32'h41c1f29c, 32'hc2a7a684};
test_output[1343] = '{32'h42aeb91b};
test_index[1343] = '{4};
test_input[10752:10759] = '{32'hc1fd906d, 32'hc19d4ea0, 32'hc0202f08, 32'hc214e1e2, 32'h42ba8a3a, 32'hc1d9d82d, 32'hc2901f70, 32'hc1fe5dba};
test_output[1344] = '{32'h42ba8a3a};
test_index[1344] = '{4};
test_input[10760:10767] = '{32'h424940e5, 32'hc208076c, 32'hc238c5ba, 32'hc2a77bae, 32'hc2812d58, 32'h42071335, 32'hc1602990, 32'h42c3bf05};
test_output[1345] = '{32'h42c3bf05};
test_index[1345] = '{7};
test_input[10768:10775] = '{32'hc266bb6d, 32'hc1ddedba, 32'hc28b1790, 32'hc0ec707b, 32'hc0fe7385, 32'h42b430e0, 32'h42459a90, 32'hc1acbfe5};
test_output[1346] = '{32'h42b430e0};
test_index[1346] = '{5};
test_input[10776:10783] = '{32'h419a933d, 32'hc1c8e1f3, 32'h42a83d56, 32'h42978b74, 32'hc141c31c, 32'h4264f2bb, 32'h422a9486, 32'h42226cdd};
test_output[1347] = '{32'h42a83d56};
test_index[1347] = '{2};
test_input[10784:10791] = '{32'hc2526af2, 32'h41bc2bab, 32'h41fe3125, 32'h41cfce68, 32'h41b4caaf, 32'hc2a0d629, 32'h4256aa48, 32'hc1ffd49e};
test_output[1348] = '{32'h4256aa48};
test_index[1348] = '{6};
test_input[10792:10799] = '{32'hc245625e, 32'hc2bfd334, 32'hc2a7071e, 32'hc2707b18, 32'h423c74f6, 32'hc1dd0e2f, 32'h4274c62a, 32'hc294a3b7};
test_output[1349] = '{32'h4274c62a};
test_index[1349] = '{6};
test_input[10800:10807] = '{32'hc1a6a3f0, 32'hc2694764, 32'hc1ecab0f, 32'h415bc20d, 32'h42b1e7a9, 32'h414e9885, 32'h42aff40c, 32'h42b9c65d};
test_output[1350] = '{32'h42b9c65d};
test_index[1350] = '{7};
test_input[10808:10815] = '{32'hc19ebeaf, 32'hc2553db7, 32'hc1f2fabf, 32'h42915138, 32'hc2c0468c, 32'h424def43, 32'hc1864ce2, 32'h418cf247};
test_output[1351] = '{32'h42915138};
test_index[1351] = '{3};
test_input[10816:10823] = '{32'h41ea7915, 32'hc1d770b6, 32'h41612cf6, 32'h42954309, 32'hc289978b, 32'hc2ad4a33, 32'h426fe6a5, 32'hc2867cf4};
test_output[1352] = '{32'h42954309};
test_index[1352] = '{3};
test_input[10824:10831] = '{32'hc216824d, 32'hc24bceb6, 32'h40c771ca, 32'hc2277c3f, 32'h419b5d90, 32'hc27f460c, 32'hc2b4000b, 32'h4280159a};
test_output[1353] = '{32'h4280159a};
test_index[1353] = '{7};
test_input[10832:10839] = '{32'h41be3790, 32'hc24b4cff, 32'hc2c4ea4f, 32'hc232be00, 32'h4272157b, 32'hc2b51f1f, 32'h42c012c5, 32'h40c42ddc};
test_output[1354] = '{32'h42c012c5};
test_index[1354] = '{6};
test_input[10840:10847] = '{32'hc25c95f0, 32'h3fd8eed8, 32'hc282a80d, 32'hc2730aa2, 32'hc27ac7f0, 32'hc1f1ff57, 32'h42c5acd8, 32'h429de485};
test_output[1355] = '{32'h42c5acd8};
test_index[1355] = '{6};
test_input[10848:10855] = '{32'h4204bf6c, 32'hc2497131, 32'hc1bb8349, 32'h42c695e9, 32'h42073acb, 32'hc2a78030, 32'hc2b526b7, 32'h42a84691};
test_output[1356] = '{32'h42c695e9};
test_index[1356] = '{3};
test_input[10856:10863] = '{32'h427732c8, 32'hc17f8a8a, 32'h427437f0, 32'hc24eb677, 32'hc1b7fb4c, 32'hc1347c2b, 32'h42920ec4, 32'hc28eaadf};
test_output[1357] = '{32'h42920ec4};
test_index[1357] = '{6};
test_input[10864:10871] = '{32'hc0831373, 32'hc292791c, 32'h42271191, 32'h424ae906, 32'h42c37f27, 32'h420455c2, 32'hc293df71, 32'h41e48214};
test_output[1358] = '{32'h42c37f27};
test_index[1358] = '{4};
test_input[10872:10879] = '{32'hc12bae99, 32'hc28cb659, 32'hc2a33e00, 32'hc29d9837, 32'hc2af7dd7, 32'hc2885e5f, 32'h40958c73, 32'h421f799b};
test_output[1359] = '{32'h421f799b};
test_index[1359] = '{7};
test_input[10880:10887] = '{32'h4260885a, 32'hc260c5e6, 32'h42a69543, 32'hc2a99068, 32'hc174e749, 32'hc2b8b715, 32'hc1244a5c, 32'h427a88d3};
test_output[1360] = '{32'h42a69543};
test_index[1360] = '{2};
test_input[10888:10895] = '{32'h425b27c8, 32'hc240b85e, 32'h42b207f8, 32'hc1fe7b29, 32'h4123481d, 32'h41894e6b, 32'hc196b1b2, 32'h42903876};
test_output[1361] = '{32'h42b207f8};
test_index[1361] = '{2};
test_input[10896:10903] = '{32'hbf26cb55, 32'h407a235b, 32'h42ac6c87, 32'hc2569e30, 32'hc23ff857, 32'hc224b4d7, 32'h420bdf31, 32'h42a9a576};
test_output[1362] = '{32'h42ac6c87};
test_index[1362] = '{2};
test_input[10904:10911] = '{32'hc2a00c81, 32'h428b4c48, 32'hc1feaa1c, 32'h4144d24a, 32'hc2c04c61, 32'h41d7642e, 32'hc2b427df, 32'h41b0d7e5};
test_output[1363] = '{32'h428b4c48};
test_index[1363] = '{1};
test_input[10912:10919] = '{32'h4290645f, 32'h42802b58, 32'hc0d4e730, 32'h42833656, 32'h416b84cc, 32'h41a09688, 32'h420446cd, 32'h41da1065};
test_output[1364] = '{32'h4290645f};
test_index[1364] = '{0};
test_input[10920:10927] = '{32'hc1935c74, 32'hc014a86a, 32'h4190da5e, 32'h426ee4f1, 32'hc1375cbf, 32'h421a9ac9, 32'h42769643, 32'h417649fd};
test_output[1365] = '{32'h42769643};
test_index[1365] = '{6};
test_input[10928:10935] = '{32'h421809f5, 32'h41b1a1bf, 32'hc2b18280, 32'hc1953f7b, 32'hc24c13fe, 32'hc2a5bf06, 32'hc2ac4e0f, 32'hc2adf389};
test_output[1366] = '{32'h421809f5};
test_index[1366] = '{0};
test_input[10936:10943] = '{32'h42434528, 32'hc212171d, 32'h420b5f70, 32'hc2013c5a, 32'hc270bd09, 32'hc1fe2036, 32'h426f6e00, 32'hc252f398};
test_output[1367] = '{32'h426f6e00};
test_index[1367] = '{6};
test_input[10944:10951] = '{32'h419fc275, 32'h40d7ff8c, 32'h428c4eee, 32'h416256ff, 32'hc2a19e57, 32'h42b02acb, 32'h422c3730, 32'hc1cea48a};
test_output[1368] = '{32'h42b02acb};
test_index[1368] = '{5};
test_input[10952:10959] = '{32'h411b9a55, 32'hc2597d93, 32'hc2ab457d, 32'hc278752d, 32'h41577b2b, 32'hc1d63440, 32'hc27443b5, 32'h4288bcf1};
test_output[1369] = '{32'h4288bcf1};
test_index[1369] = '{7};
test_input[10960:10967] = '{32'hc2bc0823, 32'h4280cae1, 32'h420441fd, 32'hc226b44d, 32'hc21c82c9, 32'h4285556e, 32'hc23a1158, 32'hc2421435};
test_output[1370] = '{32'h4285556e};
test_index[1370] = '{5};
test_input[10968:10975] = '{32'hc2a9876b, 32'h42a67c64, 32'hc04d04c6, 32'hc1e4750e, 32'hc2b1c2f3, 32'hc20eb952, 32'h421b2045, 32'h41e2dd4b};
test_output[1371] = '{32'h42a67c64};
test_index[1371] = '{1};
test_input[10976:10983] = '{32'h429a8458, 32'h418d8722, 32'h42a38bbe, 32'hc048cebf, 32'h4212fb46, 32'hc1b49d68, 32'h42a48700, 32'h42850708};
test_output[1372] = '{32'h42a48700};
test_index[1372] = '{6};
test_input[10984:10991] = '{32'h41f141db, 32'h42b5b5e0, 32'h4212d5c5, 32'hc180e50f, 32'h429a6066, 32'hc1123097, 32'hc2348ffd, 32'hc29dfba2};
test_output[1373] = '{32'h42b5b5e0};
test_index[1373] = '{1};
test_input[10992:10999] = '{32'h4253f379, 32'hc0e6c46b, 32'hc29fc2b2, 32'hc2aabd09, 32'h41bd962b, 32'hc26da965, 32'hbff59a81, 32'h42b5fc84};
test_output[1374] = '{32'h42b5fc84};
test_index[1374] = '{7};
test_input[11000:11007] = '{32'h42a2ee04, 32'h414abbc3, 32'h41fb4a5b, 32'hc2960abc, 32'h4242516b, 32'hc27aeebf, 32'h41761aeb, 32'h42bf8384};
test_output[1375] = '{32'h42bf8384};
test_index[1375] = '{7};
test_input[11008:11015] = '{32'hc15c52e8, 32'hc25f6096, 32'hc2899ad9, 32'hc1871820, 32'hc0f29e52, 32'h41b1aa2f, 32'hc1729609, 32'hc1943db0};
test_output[1376] = '{32'h41b1aa2f};
test_index[1376] = '{5};
test_input[11016:11023] = '{32'hc26e18a3, 32'h41fb7f12, 32'hc22dfa46, 32'h426c72af, 32'hc23a5c1a, 32'hc197a329, 32'hc2353da1, 32'h4290227e};
test_output[1377] = '{32'h4290227e};
test_index[1377] = '{7};
test_input[11024:11031] = '{32'hc2af1b81, 32'hc2056eaf, 32'h4004e2e6, 32'h42ad7ee6, 32'hc29ffaf5, 32'hc289f30d, 32'hc2523cad, 32'h4270299b};
test_output[1378] = '{32'h42ad7ee6};
test_index[1378] = '{3};
test_input[11032:11039] = '{32'hc2546973, 32'hc28f1c14, 32'h4255f5b1, 32'h427ab006, 32'hc2289f6a, 32'hc287d84a, 32'h41de00c8, 32'hc2c06293};
test_output[1379] = '{32'h427ab006};
test_index[1379] = '{3};
test_input[11040:11047] = '{32'hc23bbe92, 32'hc14cd4f2, 32'h410ad372, 32'h42a6600d, 32'h423152de, 32'h41c35cd3, 32'h41eba9b0, 32'hc22b3ad3};
test_output[1380] = '{32'h42a6600d};
test_index[1380] = '{3};
test_input[11048:11055] = '{32'hc29c890c, 32'h420e57e0, 32'h41c08bf9, 32'h4250e279, 32'hc245f9d6, 32'h41fb580b, 32'hc28128c3, 32'h4223aac6};
test_output[1381] = '{32'h4250e279};
test_index[1381] = '{3};
test_input[11056:11063] = '{32'hc20cc880, 32'hc285863f, 32'hc230f05c, 32'hc1938ddb, 32'h42195522, 32'hc0e74e9d, 32'h429cb2e1, 32'hc0dcb9ff};
test_output[1382] = '{32'h429cb2e1};
test_index[1382] = '{6};
test_input[11064:11071] = '{32'hc2ab6f6d, 32'hc2c0ea16, 32'hc1a19e60, 32'hc298552d, 32'hc2c37773, 32'h42255ed0, 32'hc2aa1866, 32'hc2bea900};
test_output[1383] = '{32'h42255ed0};
test_index[1383] = '{5};
test_input[11072:11079] = '{32'h414049c5, 32'hc1dcb608, 32'hc1f79e81, 32'h40202edd, 32'h42bfba42, 32'hc2c3e706, 32'hc2078fdc, 32'h42464813};
test_output[1384] = '{32'h42bfba42};
test_index[1384] = '{4};
test_input[11080:11087] = '{32'hc20a23e5, 32'hc1b6ba12, 32'h42387a50, 32'hc22dc558, 32'h42078eec, 32'hc25b1979, 32'hc2103a6e, 32'hc2154705};
test_output[1385] = '{32'h42387a50};
test_index[1385] = '{2};
test_input[11088:11095] = '{32'hc261a91e, 32'hc0c7fac2, 32'hc19988d1, 32'hc2b16b24, 32'hc2a5bbb7, 32'hc2c74ddf, 32'hc2b64c56, 32'h413ed0f2};
test_output[1386] = '{32'h413ed0f2};
test_index[1386] = '{7};
test_input[11096:11103] = '{32'hc2402ccc, 32'h3d95fd4f, 32'hc23c6e6e, 32'h42033a7f, 32'h429705f6, 32'hc26d799c, 32'hc27cc522, 32'h420fb6e3};
test_output[1387] = '{32'h429705f6};
test_index[1387] = '{4};
test_input[11104:11111] = '{32'hc2a16805, 32'hc13b602a, 32'hc16e7500, 32'hc18a453f, 32'h429870bb, 32'h42be0114, 32'hc155aac1, 32'h42c2004b};
test_output[1388] = '{32'h42c2004b};
test_index[1388] = '{7};
test_input[11112:11119] = '{32'hc207a725, 32'hc29021da, 32'hc232b9da, 32'hc05b79d9, 32'hc117fd5a, 32'hc29bf977, 32'hc2acee1b, 32'hc1790d5a};
test_output[1389] = '{32'hc05b79d9};
test_index[1389] = '{3};
test_input[11120:11127] = '{32'hbfce166b, 32'h4261d262, 32'hc2175500, 32'h42bb8199, 32'h41c717a1, 32'hc25d14cd, 32'hc281a85e, 32'hc1c45ada};
test_output[1390] = '{32'h42bb8199};
test_index[1390] = '{3};
test_input[11128:11135] = '{32'hc1abc7be, 32'h4228478e, 32'hc1b1025e, 32'hc1f92833, 32'h4221e72c, 32'h4184faa4, 32'hc205d41c, 32'h42acb01d};
test_output[1391] = '{32'h42acb01d};
test_index[1391] = '{7};
test_input[11136:11143] = '{32'hc286cad7, 32'hc289a61e, 32'hc2417bbe, 32'hc143799c, 32'hbc426b96, 32'h41b06f9b, 32'hc2672f24, 32'hbf907f61};
test_output[1392] = '{32'h41b06f9b};
test_index[1392] = '{5};
test_input[11144:11151] = '{32'hc2891261, 32'h42960cef, 32'h42b58f2f, 32'hc2bee7ac, 32'hc21ad3d6, 32'hc29d7ca3, 32'h428ec6d4, 32'hc00cee81};
test_output[1393] = '{32'h42b58f2f};
test_index[1393] = '{2};
test_input[11152:11159] = '{32'hc22ba9b0, 32'h42b88dde, 32'hc2c6d763, 32'h42837c0d, 32'hc29a4a4c, 32'h42440d33, 32'h42647111, 32'hc2b05d32};
test_output[1394] = '{32'h42b88dde};
test_index[1394] = '{1};
test_input[11160:11167] = '{32'hc282a76c, 32'hc256946b, 32'hc2bd5af2, 32'hc03b99f4, 32'hc2bd9217, 32'h42b38c58, 32'h41bb131e, 32'h4296421f};
test_output[1395] = '{32'h42b38c58};
test_index[1395] = '{5};
test_input[11168:11175] = '{32'h41fc6ceb, 32'h424b06f9, 32'hc0c4d014, 32'hc27fe43e, 32'hc28a1127, 32'h4247dcfe, 32'h40dba17c, 32'h4282695a};
test_output[1396] = '{32'h4282695a};
test_index[1396] = '{7};
test_input[11176:11183] = '{32'h427e751d, 32'hc28386ab, 32'hc2b19e5b, 32'h426d1c20, 32'h42184b0f, 32'h4281bcb7, 32'hc2ab87db, 32'h42b807fe};
test_output[1397] = '{32'h42b807fe};
test_index[1397] = '{7};
test_input[11184:11191] = '{32'h42910256, 32'h42a15547, 32'h428a963a, 32'h41d7acd0, 32'hc1c4bf72, 32'h42bad22b, 32'hc224a7b9, 32'hc1184ca7};
test_output[1398] = '{32'h42bad22b};
test_index[1398] = '{5};
test_input[11192:11199] = '{32'hc27817dc, 32'hc192cdb1, 32'hc02b6a9e, 32'h42750ba8, 32'hc0f27022, 32'hc2ab1591, 32'h426a8564, 32'h42064ea9};
test_output[1399] = '{32'h42750ba8};
test_index[1399] = '{3};
test_input[11200:11207] = '{32'h42289e1b, 32'h414078f3, 32'h41ee7681, 32'hc0ce62fb, 32'h429e7d4b, 32'h41201862, 32'hc187b4a2, 32'h412108af};
test_output[1400] = '{32'h429e7d4b};
test_index[1400] = '{4};
test_input[11208:11215] = '{32'h41862179, 32'h4201be36, 32'hc2b0c7ae, 32'h42ae81cd, 32'h42c6f999, 32'h42a6e7ee, 32'h42b338b9, 32'h4265df02};
test_output[1401] = '{32'h42c6f999};
test_index[1401] = '{4};
test_input[11216:11223] = '{32'h4195be8f, 32'h429c177c, 32'hc2930dcc, 32'h41f85e5c, 32'h4287b833, 32'hc28c5068, 32'h425988a7, 32'h423a7bd6};
test_output[1402] = '{32'h429c177c};
test_index[1402] = '{1};
test_input[11224:11231] = '{32'h419f2c60, 32'h42a979af, 32'hc1ef6f60, 32'h4178282f, 32'h424e3f29, 32'hc214f452, 32'hc2c58199, 32'h424f0cea};
test_output[1403] = '{32'h42a979af};
test_index[1403] = '{1};
test_input[11232:11239] = '{32'hbf400a0a, 32'hc200153c, 32'hc2b2fae7, 32'h42c5e771, 32'h4082f7ba, 32'h421d2e3c, 32'h418f8d1d, 32'hc1a97f43};
test_output[1404] = '{32'h42c5e771};
test_index[1404] = '{3};
test_input[11240:11247] = '{32'hc286741c, 32'h4286c4f0, 32'h41d4cbe4, 32'h410a37f0, 32'hc2b798ca, 32'h423c5249, 32'h4191ff27, 32'hc11f9dec};
test_output[1405] = '{32'h4286c4f0};
test_index[1405] = '{1};
test_input[11248:11255] = '{32'hc28d768f, 32'hc2808ee9, 32'hc2847c97, 32'h424f4567, 32'hc2ab96b6, 32'hc29de0af, 32'h42ab2447, 32'hc1db8c0b};
test_output[1406] = '{32'h42ab2447};
test_index[1406] = '{6};
test_input[11256:11263] = '{32'hc223fd8a, 32'h3e92bfda, 32'h42b898b9, 32'hc22ca691, 32'hc2b0c153, 32'hc2151b82, 32'hc29ed983, 32'h41a77d24};
test_output[1407] = '{32'h42b898b9};
test_index[1407] = '{2};
test_input[11264:11271] = '{32'h4247e8b1, 32'h42070cf0, 32'hc2923613, 32'h411dad94, 32'h42a3efef, 32'h40e38d6e, 32'hc1a4ed15, 32'hc26fdd3e};
test_output[1408] = '{32'h42a3efef};
test_index[1408] = '{4};
test_input[11272:11279] = '{32'hc2562260, 32'h41ea7adf, 32'h42c0daab, 32'hc295e729, 32'h42b5d0cb, 32'h4207489d, 32'hc2bee0b2, 32'hc2b1b401};
test_output[1409] = '{32'h42c0daab};
test_index[1409] = '{2};
test_input[11280:11287] = '{32'hc1b09b90, 32'h41a4a2ee, 32'hc18167a7, 32'h41f506ac, 32'hc25b7622, 32'hc1db594b, 32'h42410c2b, 32'h42bce39d};
test_output[1410] = '{32'h42bce39d};
test_index[1410] = '{7};
test_input[11288:11295] = '{32'hc2b2c1cd, 32'h42016297, 32'hc1c81537, 32'hc28d438e, 32'h41d16e71, 32'h4044caa8, 32'hc1fe933f, 32'hc2b386a0};
test_output[1411] = '{32'h42016297};
test_index[1411] = '{1};
test_input[11296:11303] = '{32'h4278d0eb, 32'h4282a56a, 32'h4132604b, 32'hc29f861e, 32'hc245a26c, 32'hc1431c38, 32'hc27980e5, 32'h41d56021};
test_output[1412] = '{32'h4282a56a};
test_index[1412] = '{1};
test_input[11304:11311] = '{32'hc2aeb875, 32'hc2181fbf, 32'hc2ae176c, 32'hc2527a5c, 32'h41a0df83, 32'h42b78602, 32'h4034cd16, 32'hc1d79326};
test_output[1413] = '{32'h42b78602};
test_index[1413] = '{5};
test_input[11312:11319] = '{32'h42038a77, 32'hc25aa5d1, 32'hc2109806, 32'h429c2518, 32'hc27030a0, 32'h426b4b3b, 32'hc28844e3, 32'h3f88aba4};
test_output[1414] = '{32'h429c2518};
test_index[1414] = '{3};
test_input[11320:11327] = '{32'hc169a1f7, 32'hc169e511, 32'hc009dc6f, 32'hc280d5ce, 32'hc29a56f3, 32'hc2829e7c, 32'hc2bc3766, 32'hc26d60c6};
test_output[1415] = '{32'hc009dc6f};
test_index[1415] = '{2};
test_input[11328:11335] = '{32'h4264f02e, 32'h4202da4d, 32'hc194f0ea, 32'hc1b86a85, 32'h41a5931b, 32'hc1553c06, 32'h40d6a594, 32'h4241da88};
test_output[1416] = '{32'h4264f02e};
test_index[1416] = '{0};
test_input[11336:11343] = '{32'hc2a6ffd1, 32'hc2996eec, 32'h4299a9a7, 32'hc2c6097b, 32'h42a7fb2c, 32'h420b543e, 32'h42242cf6, 32'hc2343d9e};
test_output[1417] = '{32'h42a7fb2c};
test_index[1417] = '{4};
test_input[11344:11351] = '{32'hc1b38373, 32'hc2125c26, 32'h41beaaf1, 32'h4270b6a7, 32'h428e2132, 32'h410f1a25, 32'h40571952, 32'hc27f6012};
test_output[1418] = '{32'h428e2132};
test_index[1418] = '{4};
test_input[11352:11359] = '{32'hc1065515, 32'hc285c206, 32'h4237a4cd, 32'h425f5822, 32'h422a665d, 32'h41822433, 32'hc2212c39, 32'hc295a985};
test_output[1419] = '{32'h425f5822};
test_index[1419] = '{3};
test_input[11360:11367] = '{32'h42bdfb07, 32'hc2943fd1, 32'h42868ca3, 32'hc1d6a55a, 32'h428fbaf8, 32'h425dd4d0, 32'hc23dd28c, 32'hc1a093bc};
test_output[1420] = '{32'h42bdfb07};
test_index[1420] = '{0};
test_input[11368:11375] = '{32'h428970ac, 32'hc1ec85e2, 32'hc2c6ddd1, 32'hc2032ad4, 32'hc29dc293, 32'h4297e2ba, 32'hc1f74a97, 32'hc05bf391};
test_output[1421] = '{32'h4297e2ba};
test_index[1421] = '{5};
test_input[11376:11383] = '{32'hc1bd2c61, 32'hc242c25c, 32'h42bfad75, 32'hc2b7e397, 32'h40cbc964, 32'h42144797, 32'hc2a498ed, 32'hc117d2d0};
test_output[1422] = '{32'h42bfad75};
test_index[1422] = '{2};
test_input[11384:11391] = '{32'h40fcd972, 32'hc18d886f, 32'hbfb7a326, 32'h4249abc5, 32'hc22a2d11, 32'hbf65ad8b, 32'hc23f8ea3, 32'hc2833006};
test_output[1423] = '{32'h4249abc5};
test_index[1423] = '{3};
test_input[11392:11399] = '{32'h421d8601, 32'h41a27b90, 32'hc297ea20, 32'hc26ca0b5, 32'hc22dfb04, 32'h42a3980e, 32'h42343d2c, 32'h42ae8b04};
test_output[1424] = '{32'h42ae8b04};
test_index[1424] = '{7};
test_input[11400:11407] = '{32'h42b6d4e6, 32'hc2726c6a, 32'h4299fa9c, 32'h42a50db2, 32'hc1d6da90, 32'hc071a1a4, 32'h3f0071e8, 32'hc2b29051};
test_output[1425] = '{32'h42b6d4e6};
test_index[1425] = '{0};
test_input[11408:11415] = '{32'hc2471ab6, 32'hc1d405ec, 32'hc0418230, 32'hc1aab2b8, 32'hc28517b5, 32'h422fb72b, 32'hc1690c12, 32'hc0fc6603};
test_output[1426] = '{32'h422fb72b};
test_index[1426] = '{5};
test_input[11416:11423] = '{32'h42c418c6, 32'hc01abe80, 32'hc2b8d51f, 32'hc0e30eda, 32'hc225fce5, 32'hc28cfdc7, 32'hc293956f, 32'hc2341f20};
test_output[1427] = '{32'h42c418c6};
test_index[1427] = '{0};
test_input[11424:11431] = '{32'h429df289, 32'hc2a80a96, 32'hc24da0b2, 32'hc20b6229, 32'hc288abe8, 32'hc2c7db83, 32'h426a4dee, 32'hc298dfbb};
test_output[1428] = '{32'h429df289};
test_index[1428] = '{0};
test_input[11432:11439] = '{32'h429edebd, 32'hc1e4c3b6, 32'h41b979c6, 32'hc26c7c29, 32'hc28ed552, 32'h428c799c, 32'h423d324d, 32'hc03399bf};
test_output[1429] = '{32'h429edebd};
test_index[1429] = '{0};
test_input[11440:11447] = '{32'hbf19aace, 32'h419af81d, 32'hc2ae1ec2, 32'h424ad586, 32'hc27b4839, 32'hc2638d07, 32'hc105d1ee, 32'h41e2f452};
test_output[1430] = '{32'h424ad586};
test_index[1430] = '{3};
test_input[11448:11455] = '{32'hc27da39c, 32'h429580a9, 32'h41ed54ea, 32'h4293943e, 32'hc0bd394a, 32'h41e44039, 32'h429fb217, 32'hc286e584};
test_output[1431] = '{32'h429fb217};
test_index[1431] = '{6};
test_input[11456:11463] = '{32'h4285771e, 32'h412e07cc, 32'hc29561f5, 32'h41ea216a, 32'h42778055, 32'h4204dc99, 32'h426876a3, 32'hc1ecf961};
test_output[1432] = '{32'h4285771e};
test_index[1432] = '{0};
test_input[11464:11471] = '{32'h42071dd5, 32'hc223677e, 32'hc1a74021, 32'hc28046c9, 32'hc1741fa5, 32'hc19044b3, 32'h4241f97e, 32'h42b6bb8f};
test_output[1433] = '{32'h42b6bb8f};
test_index[1433] = '{7};
test_input[11472:11479] = '{32'h4288ff13, 32'h429edcc6, 32'hc2bd7382, 32'hc1c31870, 32'h42888cd3, 32'hc20f92d3, 32'h41a009a0, 32'hc213f96a};
test_output[1434] = '{32'h429edcc6};
test_index[1434] = '{1};
test_input[11480:11487] = '{32'h422ee0f2, 32'h4192c8d2, 32'h42630db9, 32'h4297c7e2, 32'hc11432f5, 32'hc2256bce, 32'h426bece4, 32'h42b5ba3e};
test_output[1435] = '{32'h42b5ba3e};
test_index[1435] = '{7};
test_input[11488:11495] = '{32'h4285b366, 32'h424b0d36, 32'hc20ac932, 32'h42bbeb8b, 32'hc2103692, 32'hc224cf87, 32'hbf5b350c, 32'hc0af7965};
test_output[1436] = '{32'h42bbeb8b};
test_index[1436] = '{3};
test_input[11496:11503] = '{32'hc258b043, 32'hc2b94d8c, 32'h417b4280, 32'hc290b98b, 32'h4187d751, 32'h4253ad96, 32'hc25bdf07, 32'h4257db85};
test_output[1437] = '{32'h4257db85};
test_index[1437] = '{7};
test_input[11504:11511] = '{32'h426a40fa, 32'h418e836c, 32'h41893843, 32'h42641f5d, 32'h41c3e397, 32'h42a984d7, 32'h4205a6c9, 32'h42baad2e};
test_output[1438] = '{32'h42baad2e};
test_index[1438] = '{7};
test_input[11512:11519] = '{32'h425c284f, 32'h41ee8d5f, 32'h423c08c9, 32'h42910525, 32'h41215994, 32'hc2ac8885, 32'hc2b55c76, 32'hc1e59069};
test_output[1439] = '{32'h42910525};
test_index[1439] = '{3};
test_input[11520:11527] = '{32'h41697b4a, 32'hc2ae4d8b, 32'hc1e0b726, 32'hc176f783, 32'hc239a82d, 32'hc0a0af24, 32'h42a1ca16, 32'h41828524};
test_output[1440] = '{32'h42a1ca16};
test_index[1440] = '{6};
test_input[11528:11535] = '{32'h422abafc, 32'h42247bb2, 32'h427a11a9, 32'h42a9e520, 32'h41edfdea, 32'h4226ad78, 32'h429ccdba, 32'h42425642};
test_output[1441] = '{32'h42a9e520};
test_index[1441] = '{3};
test_input[11536:11543] = '{32'hc2990a0d, 32'hc281be33, 32'hc1862fb8, 32'h4023d6ca, 32'h428532b9, 32'h40fca72b, 32'h42c0028c, 32'hc2c04854};
test_output[1442] = '{32'h42c0028c};
test_index[1442] = '{6};
test_input[11544:11551] = '{32'hc296da48, 32'hc1fa1373, 32'h423ae1d4, 32'h41282cba, 32'hc284e76d, 32'hc2c7f6aa, 32'h41c2d48d, 32'h42a2c27a};
test_output[1443] = '{32'h42a2c27a};
test_index[1443] = '{7};
test_input[11552:11559] = '{32'h4223f357, 32'h412b2e89, 32'h42592a68, 32'hc292da0a, 32'hc282b0db, 32'h42ad0f8a, 32'h426ecd9f, 32'hc2ada92c};
test_output[1444] = '{32'h42ad0f8a};
test_index[1444] = '{5};
test_input[11560:11567] = '{32'h41e10ec2, 32'h429b43e0, 32'h4230bba2, 32'h42b5eb93, 32'hc19ecebc, 32'hc059d5ad, 32'h42310404, 32'h4085d3d6};
test_output[1445] = '{32'h42b5eb93};
test_index[1445] = '{3};
test_input[11568:11575] = '{32'h427e610a, 32'hc1b395a0, 32'hc2935c69, 32'hc2632b95, 32'hc04b5f63, 32'hc1b1cb05, 32'hc171cd47, 32'h42325436};
test_output[1446] = '{32'h427e610a};
test_index[1446] = '{0};
test_input[11576:11583] = '{32'hc2acacf4, 32'hc29d7e51, 32'hc280948f, 32'h41568ea1, 32'h422536f6, 32'h42b01210, 32'hc2775f98, 32'hc2c05f6f};
test_output[1447] = '{32'h42b01210};
test_index[1447] = '{5};
test_input[11584:11591] = '{32'h42b8834f, 32'h4181c11a, 32'hc2aeddd1, 32'h423b60ea, 32'hc2964ccf, 32'hc2b797ce, 32'h4222639f, 32'h40d70b1f};
test_output[1448] = '{32'h42b8834f};
test_index[1448] = '{0};
test_input[11592:11599] = '{32'h4286a0c9, 32'hc277ca9b, 32'hc2a2ab36, 32'h421bd7ab, 32'h428f68c8, 32'h40a0c22b, 32'h42beddfc, 32'hc28a3bc3};
test_output[1449] = '{32'h42beddfc};
test_index[1449] = '{6};
test_input[11600:11607] = '{32'hc287e3f6, 32'hc1a92911, 32'hc161f412, 32'h42c2e93b, 32'h42195388, 32'h41be80a3, 32'hc17f7dfd, 32'hbff1c9f3};
test_output[1450] = '{32'h42c2e93b};
test_index[1450] = '{3};
test_input[11608:11615] = '{32'h4240aa16, 32'hc2ab1ed6, 32'hc2988ba6, 32'hc25faa97, 32'hc2657531, 32'hc239548a, 32'h42924417, 32'h42b23efd};
test_output[1451] = '{32'h42b23efd};
test_index[1451] = '{7};
test_input[11616:11623] = '{32'h425dca62, 32'h4214f331, 32'h4283cb40, 32'hc2892193, 32'hc2955075, 32'hc2aca667, 32'h42c3c7cf, 32'h417fafad};
test_output[1452] = '{32'h42c3c7cf};
test_index[1452] = '{6};
test_input[11624:11631] = '{32'hc222a057, 32'h42b83211, 32'h42bb3296, 32'hc23b3c48, 32'hc040c22e, 32'hc1a33c88, 32'h3fe4f4a1, 32'h41c4221c};
test_output[1453] = '{32'h42bb3296};
test_index[1453] = '{2};
test_input[11632:11639] = '{32'h42320e2a, 32'hc2b3ab54, 32'h42a23e22, 32'h42bd15f9, 32'h42c7cacf, 32'h42ac4370, 32'hbeab99f4, 32'h42885009};
test_output[1454] = '{32'h42c7cacf};
test_index[1454] = '{4};
test_input[11640:11647] = '{32'h428b5402, 32'h4271c344, 32'h42708dbf, 32'h42abaea8, 32'hc2850360, 32'hc16022b8, 32'hbe0cb4a5, 32'hc2149c7f};
test_output[1455] = '{32'h42abaea8};
test_index[1455] = '{3};
test_input[11648:11655] = '{32'hc1e92ce7, 32'hc214c3d5, 32'h41dd1f45, 32'h424490e4, 32'h40d10618, 32'hc26d9e88, 32'hc054a8f9, 32'hc2bc9f4d};
test_output[1456] = '{32'h424490e4};
test_index[1456] = '{3};
test_input[11656:11663] = '{32'h427d9a11, 32'hc29b52fc, 32'hc15b926f, 32'hc1334c9a, 32'hc1b39327, 32'h4238ac07, 32'h420799c9, 32'hc15d368e};
test_output[1457] = '{32'h427d9a11};
test_index[1457] = '{0};
test_input[11664:11671] = '{32'h4240922b, 32'hc26fef2f, 32'h4243ffaf, 32'h42867fda, 32'h42387ab5, 32'h40f8fe3b, 32'hc1568b17, 32'hc1f4d219};
test_output[1458] = '{32'h42867fda};
test_index[1458] = '{3};
test_input[11672:11679] = '{32'h429f1bd0, 32'h40ca1445, 32'h4294ea22, 32'h428b9d3f, 32'hc1271a72, 32'hc210df6e, 32'h42730841, 32'h4053c257};
test_output[1459] = '{32'h429f1bd0};
test_index[1459] = '{0};
test_input[11680:11687] = '{32'h41f12a89, 32'hc2bc8e76, 32'hc2673d4d, 32'hc2208576, 32'hc2472672, 32'h428e0a78, 32'hc1b5de3f, 32'hc2039c34};
test_output[1460] = '{32'h428e0a78};
test_index[1460] = '{5};
test_input[11688:11695] = '{32'hc29a9a6a, 32'h420253d1, 32'h416128dd, 32'hc216cf40, 32'hc2731838, 32'hc295191b, 32'hc0ebe4a3, 32'h42c4cbe5};
test_output[1461] = '{32'h42c4cbe5};
test_index[1461] = '{7};
test_input[11696:11703] = '{32'hc1af519b, 32'hc1dc9e4e, 32'h42a7cb05, 32'h42b9ee27, 32'h42b51717, 32'hc2c21164, 32'hc2baa567, 32'h42989cb4};
test_output[1462] = '{32'h42b9ee27};
test_index[1462] = '{3};
test_input[11704:11711] = '{32'h427ee7eb, 32'hc130ed8c, 32'h426dc23b, 32'hc24134b3, 32'hc2970c73, 32'h41cd55be, 32'h4211fb6a, 32'hc21aedb5};
test_output[1463] = '{32'h427ee7eb};
test_index[1463] = '{0};
test_input[11712:11719] = '{32'h42ba75c3, 32'h4138b471, 32'hc217f4e3, 32'hc27004a6, 32'hc2840641, 32'hc20a0037, 32'hc23a7d18, 32'h423e406e};
test_output[1464] = '{32'h42ba75c3};
test_index[1464] = '{0};
test_input[11720:11727] = '{32'hc0653f6b, 32'hc2bc1b01, 32'hc1d5cd1d, 32'h4235e27e, 32'hc28063b6, 32'hc2910709, 32'hc238f2a8, 32'h42c6189f};
test_output[1465] = '{32'h42c6189f};
test_index[1465] = '{7};
test_input[11728:11735] = '{32'h42a374a7, 32'h41154284, 32'h42b1f386, 32'hc2ad4e59, 32'hc24c290a, 32'h412cb57f, 32'hc272a0b0, 32'hc11baa50};
test_output[1466] = '{32'h42b1f386};
test_index[1466] = '{2};
test_input[11736:11743] = '{32'h4195a6e8, 32'h429a39ae, 32'hc0e3d543, 32'h42abd916, 32'h4102c3a2, 32'h42a7965b, 32'hc1e184d8, 32'h42352f3c};
test_output[1467] = '{32'h42abd916};
test_index[1467] = '{3};
test_input[11744:11751] = '{32'hc1f6dc17, 32'hc280af0c, 32'hc1ee802f, 32'hc09dba05, 32'h42828b30, 32'h428f8610, 32'h41e315ec, 32'hc27ffb26};
test_output[1468] = '{32'h428f8610};
test_index[1468] = '{5};
test_input[11752:11759] = '{32'hc2a58367, 32'hc284929b, 32'h42992f0e, 32'h4206f5db, 32'hc26983f2, 32'h41ed9e4b, 32'hc274f819, 32'h421de7cb};
test_output[1469] = '{32'h42992f0e};
test_index[1469] = '{2};
test_input[11760:11767] = '{32'hc09075f9, 32'h42aa22c0, 32'hc2474101, 32'h42ae351f, 32'hc252f6cb, 32'h421b92e1, 32'hc205b9b7, 32'h421d35c1};
test_output[1470] = '{32'h42ae351f};
test_index[1470] = '{3};
test_input[11768:11775] = '{32'hc1a904b3, 32'h42908422, 32'h42c16394, 32'h41503755, 32'hbf0dcd4b, 32'h429d2d86, 32'hc29b41af, 32'hc0fc3c37};
test_output[1471] = '{32'h42c16394};
test_index[1471] = '{2};
test_input[11776:11783] = '{32'h426f7a51, 32'hc275ba59, 32'h421ce8cd, 32'hc1ab72ef, 32'h42a41aef, 32'h4200269e, 32'h427bac4c, 32'hc2ae3d85};
test_output[1472] = '{32'h42a41aef};
test_index[1472] = '{4};
test_input[11784:11791] = '{32'h41917b4e, 32'h41b87682, 32'hc2ab6620, 32'h3f6b882c, 32'hc1829599, 32'h42bc8d91, 32'hc160f7e4, 32'hc120e761};
test_output[1473] = '{32'h42bc8d91};
test_index[1473] = '{5};
test_input[11792:11799] = '{32'h40463ac5, 32'h41b2101d, 32'hc0a72871, 32'h42a5da93, 32'hc24dd591, 32'hc1212ca9, 32'h421b1de9, 32'hc290ec79};
test_output[1474] = '{32'h42a5da93};
test_index[1474] = '{3};
test_input[11800:11807] = '{32'h421e8871, 32'hc230acd6, 32'hc1a8aecc, 32'h425f2daa, 32'hc1fd01e0, 32'h4202cd41, 32'hc25c409e, 32'h423a5d60};
test_output[1475] = '{32'h425f2daa};
test_index[1475] = '{3};
test_input[11808:11815] = '{32'h41af43e2, 32'hc27e22c4, 32'hc24f4503, 32'hc29f9beb, 32'h42bdbd2b, 32'h42b70151, 32'hc296f01b, 32'hc28e4ad3};
test_output[1476] = '{32'h42bdbd2b};
test_index[1476] = '{4};
test_input[11816:11823] = '{32'hc2baf078, 32'h42972f7b, 32'h423711a1, 32'hc205b1b4, 32'h42b6bda3, 32'hc2a4c566, 32'h42045cb7, 32'h42bac5fa};
test_output[1477] = '{32'h42bac5fa};
test_index[1477] = '{7};
test_input[11824:11831] = '{32'hc2c7009a, 32'hc2998b53, 32'h42c2f845, 32'hc253e3af, 32'h42c78474, 32'hc21c0590, 32'h4254a0f6, 32'hc2643543};
test_output[1478] = '{32'h42c78474};
test_index[1478] = '{4};
test_input[11832:11839] = '{32'hc2ad0f41, 32'hc21fa23b, 32'h4280757f, 32'hc11d6c59, 32'h421fc551, 32'hc1dbf4a4, 32'h422dbbac, 32'hc23eb7b2};
test_output[1479] = '{32'h4280757f};
test_index[1479] = '{2};
test_input[11840:11847] = '{32'hc16ca55d, 32'hc1d68eb8, 32'hc29f08b1, 32'h4167218f, 32'hc2c14892, 32'h42c4c0c6, 32'hc1eaf3dc, 32'hc1e61a79};
test_output[1480] = '{32'h42c4c0c6};
test_index[1480] = '{5};
test_input[11848:11855] = '{32'hc192bf5a, 32'h41efb11e, 32'h426ec8b1, 32'h4295f93e, 32'hc2c5cea4, 32'hc1ff6d59, 32'h41ce0abc, 32'hc2b44904};
test_output[1481] = '{32'h4295f93e};
test_index[1481] = '{3};
test_input[11856:11863] = '{32'hc2b0ca2f, 32'h4063435a, 32'hc2503e18, 32'h42a2a1a3, 32'h424d8e02, 32'h426110f2, 32'h42685b12, 32'hc2656262};
test_output[1482] = '{32'h42a2a1a3};
test_index[1482] = '{3};
test_input[11864:11871] = '{32'hc2531cc4, 32'h3e2ab28b, 32'h428b4466, 32'h41f93553, 32'h41fc94c5, 32'hc1d0af3e, 32'hc2bda12c, 32'h42941f2d};
test_output[1483] = '{32'h42941f2d};
test_index[1483] = '{7};
test_input[11872:11879] = '{32'hc2be73f2, 32'h429a1368, 32'h42bb1132, 32'hc2567e28, 32'hc1c3ee13, 32'hc22f6c21, 32'hc03ad80b, 32'h42ab98a8};
test_output[1484] = '{32'h42bb1132};
test_index[1484] = '{2};
test_input[11880:11887] = '{32'hc26033e5, 32'h4218a70f, 32'h426af616, 32'h42933c53, 32'hc293a058, 32'hc29b94ac, 32'h4296164a, 32'h41e27d7c};
test_output[1485] = '{32'h4296164a};
test_index[1485] = '{6};
test_input[11888:11895] = '{32'hc20d09ba, 32'h42c65db7, 32'hc1cf8028, 32'hc246391b, 32'hc23caf02, 32'hc2b04c86, 32'h42998fff, 32'h41a70cc1};
test_output[1486] = '{32'h42c65db7};
test_index[1486] = '{1};
test_input[11896:11903] = '{32'hc22bbb3c, 32'h42864afb, 32'h429acdee, 32'hbf3027aa, 32'h42425262, 32'h41c87277, 32'h42b1c0ac, 32'h4207a84f};
test_output[1487] = '{32'h42b1c0ac};
test_index[1487] = '{6};
test_input[11904:11911] = '{32'h41eb814b, 32'hc2896253, 32'h422c752a, 32'hc2c3df02, 32'hc2a4f0ac, 32'h42b0b2bb, 32'h4253c410, 32'h424c68db};
test_output[1488] = '{32'h42b0b2bb};
test_index[1488] = '{5};
test_input[11912:11919] = '{32'h42b8380d, 32'hc2138958, 32'hc158e31a, 32'hc20522c7, 32'hc2bf8bab, 32'hc2989c50, 32'h428254ed, 32'h41a9db63};
test_output[1489] = '{32'h42b8380d};
test_index[1489] = '{0};
test_input[11920:11927] = '{32'h41311012, 32'hc2821306, 32'hc090521a, 32'hc2a286df, 32'hc2829314, 32'hc0d115bf, 32'h4230e73e, 32'h41e517b3};
test_output[1490] = '{32'h4230e73e};
test_index[1490] = '{6};
test_input[11928:11935] = '{32'h41973304, 32'hc2aa60b5, 32'hc275534c, 32'hc281d618, 32'h4175fb0a, 32'h41e22663, 32'h42ad28cf, 32'hc1865b1d};
test_output[1491] = '{32'h42ad28cf};
test_index[1491] = '{6};
test_input[11936:11943] = '{32'h420bd434, 32'h42a2d7d8, 32'hc26d106b, 32'h41e2c1b4, 32'h428bac52, 32'h42adbad3, 32'h412adf07, 32'h417d56ba};
test_output[1492] = '{32'h42adbad3};
test_index[1492] = '{5};
test_input[11944:11951] = '{32'h4299f6b7, 32'h41c4a5ee, 32'h42baffff, 32'h42beab83, 32'hc291ae1e, 32'hc2349344, 32'hc2a2b790, 32'hc25beeed};
test_output[1493] = '{32'h42beab83};
test_index[1493] = '{3};
test_input[11952:11959] = '{32'h42965591, 32'h41da0d1e, 32'hc21600d0, 32'hc24a0aa0, 32'hc1232520, 32'h4195665f, 32'hc22d2dfe, 32'h4291281c};
test_output[1494] = '{32'h42965591};
test_index[1494] = '{0};
test_input[11960:11967] = '{32'hc2b388f4, 32'hc061b468, 32'hc24ebcfe, 32'hc209b283, 32'hc080d255, 32'hc28ecfed, 32'h42a493e8, 32'h4237c006};
test_output[1495] = '{32'h42a493e8};
test_index[1495] = '{6};
test_input[11968:11975] = '{32'hc285e719, 32'h41c8be78, 32'hc2a1950e, 32'h40dedf95, 32'h420dfc35, 32'h429648f3, 32'h42655791, 32'h428ca30e};
test_output[1496] = '{32'h429648f3};
test_index[1496] = '{5};
test_input[11976:11983] = '{32'h42329516, 32'h41c6d6e1, 32'hc1e5fa55, 32'h4287ffd9, 32'hc1733d2b, 32'h41552c8a, 32'hc0d3d0c4, 32'hc2b780f6};
test_output[1497] = '{32'h4287ffd9};
test_index[1497] = '{3};
test_input[11984:11991] = '{32'hc2a7435e, 32'h423a8123, 32'h41cb2eab, 32'hc2645346, 32'hc2036265, 32'hc1197e38, 32'h419bc842, 32'h42b54819};
test_output[1498] = '{32'h42b54819};
test_index[1498] = '{7};
test_input[11992:11999] = '{32'h41999b73, 32'hc0fd835d, 32'h42a8814d, 32'hc23df2b4, 32'hc265d233, 32'h42842335, 32'h410ba8f4, 32'h42b22f4b};
test_output[1499] = '{32'h42b22f4b};
test_index[1499] = '{7};
test_input[12000:12007] = '{32'h42078ea2, 32'h42544b53, 32'hc201eac6, 32'hc2a8f56a, 32'hc2a6f829, 32'hc29909e9, 32'hc28b0c00, 32'hc1d8f75a};
test_output[1500] = '{32'h42544b53};
test_index[1500] = '{1};
test_input[12008:12015] = '{32'h42b09ac5, 32'hc2b88370, 32'hc16a1380, 32'hc22a7154, 32'hc1448eee, 32'hc0511b60, 32'h4217234a, 32'h42bd1f84};
test_output[1501] = '{32'h42bd1f84};
test_index[1501] = '{7};
test_input[12016:12023] = '{32'h41a9c3cc, 32'hc21854fb, 32'hc2546ca8, 32'hc2b94b91, 32'h420bdfb8, 32'hc2b60783, 32'hc2afe096, 32'h424badd6};
test_output[1502] = '{32'h424badd6};
test_index[1502] = '{7};
test_input[12024:12031] = '{32'hc2a12e1b, 32'h426a15fa, 32'hc1806216, 32'h41c3896a, 32'h42896512, 32'h428c8f2f, 32'hc2c49b53, 32'h3fa4a3b5};
test_output[1503] = '{32'h428c8f2f};
test_index[1503] = '{5};
test_input[12032:12039] = '{32'hc267e57b, 32'h418b2318, 32'h424814ee, 32'hc17edc59, 32'h40a33463, 32'hc29e17fb, 32'hc2c1332a, 32'h42a7b0b1};
test_output[1504] = '{32'h42a7b0b1};
test_index[1504] = '{7};
test_input[12040:12047] = '{32'h42a7243f, 32'hc28b7ec5, 32'hc28c15b8, 32'hc2084055, 32'h42ab1ead, 32'hc2a292b0, 32'hc28d4580, 32'hbf49e8e9};
test_output[1505] = '{32'h42ab1ead};
test_index[1505] = '{4};
test_input[12048:12055] = '{32'hc234cec8, 32'h41423c83, 32'h41f17503, 32'h41bb87ca, 32'hc28fbb82, 32'h42c1055d, 32'h42c2451f, 32'hc2559230};
test_output[1506] = '{32'h42c2451f};
test_index[1506] = '{6};
test_input[12056:12063] = '{32'h42b8a4be, 32'h424991d8, 32'h42c75a6c, 32'h40484103, 32'hc2514937, 32'hc2a5d02c, 32'hc2b24f44, 32'hc20a0f67};
test_output[1507] = '{32'h42c75a6c};
test_index[1507] = '{2};
test_input[12064:12071] = '{32'hc2a87065, 32'h41da8f4d, 32'hc1d77f3e, 32'h41b7ddb8, 32'hc2b909fa, 32'hc253366d, 32'hc2690939, 32'hc20881c3};
test_output[1508] = '{32'h41da8f4d};
test_index[1508] = '{1};
test_input[12072:12079] = '{32'h4119afbd, 32'hc2204f7b, 32'h417c7509, 32'h4228057c, 32'hc2709637, 32'hc29fca09, 32'h41e6e43f, 32'h42c40df1};
test_output[1509] = '{32'h42c40df1};
test_index[1509] = '{7};
test_input[12080:12087] = '{32'hc2126897, 32'hc2516f5a, 32'hc283f5bf, 32'h41f6787b, 32'h421c8cb1, 32'hc2c66d34, 32'hc29dad1f, 32'h42304d53};
test_output[1510] = '{32'h42304d53};
test_index[1510] = '{7};
test_input[12088:12095] = '{32'hc14551ce, 32'hc184bda8, 32'hc281555d, 32'hc21d4619, 32'h41ad6976, 32'hc1442285, 32'hc262784b, 32'hc29096d0};
test_output[1511] = '{32'h41ad6976};
test_index[1511] = '{4};
test_input[12096:12103] = '{32'h423871b0, 32'hc28bd780, 32'h421fdf48, 32'hc026547f, 32'h4124a693, 32'h424c8c52, 32'h4299ee54, 32'h4269b5d0};
test_output[1512] = '{32'h4299ee54};
test_index[1512] = '{6};
test_input[12104:12111] = '{32'hc232f1a8, 32'h415f6c60, 32'h41f4685b, 32'h428db940, 32'h42c6dc28, 32'hc285dc7f, 32'h4258c057, 32'h420a2550};
test_output[1513] = '{32'h42c6dc28};
test_index[1513] = '{4};
test_input[12112:12119] = '{32'hc186d81d, 32'h41ec3f71, 32'h41ade6b4, 32'hc2092712, 32'hc232d13f, 32'hc1e9d2df, 32'hc28668ca, 32'h429cbb0c};
test_output[1514] = '{32'h429cbb0c};
test_index[1514] = '{7};
test_input[12120:12127] = '{32'hc15c39d3, 32'h42b29088, 32'hc196f28e, 32'h42bc2e13, 32'hc291f2c5, 32'h42683f2e, 32'h4242e414, 32'hc282a55d};
test_output[1515] = '{32'h42bc2e13};
test_index[1515] = '{3};
test_input[12128:12135] = '{32'h420f1914, 32'h41fce6bb, 32'hc2190dee, 32'h42844f4f, 32'hc2906b54, 32'h4265bf28, 32'hc299b48c, 32'h42c22ab5};
test_output[1516] = '{32'h42c22ab5};
test_index[1516] = '{7};
test_input[12136:12143] = '{32'hc22488d3, 32'h41d81671, 32'h4298cbf9, 32'hc29ee148, 32'hc1ebfee9, 32'hc05dff4d, 32'h4246c0f3, 32'hc2acd1ac};
test_output[1517] = '{32'h4298cbf9};
test_index[1517] = '{2};
test_input[12144:12151] = '{32'hc225b34d, 32'hbf31b6a4, 32'hc2803078, 32'hc222d2e4, 32'h410c4eb4, 32'hc2a4a6a9, 32'hc1ca30cd, 32'hc26f5720};
test_output[1518] = '{32'h410c4eb4};
test_index[1518] = '{4};
test_input[12152:12159] = '{32'h42937c49, 32'h427b91bb, 32'h427b83c8, 32'h422b7a96, 32'h4164328f, 32'h425f121d, 32'h42b29a83, 32'hc2b44b67};
test_output[1519] = '{32'h42b29a83};
test_index[1519] = '{6};
test_input[12160:12167] = '{32'h4263c75e, 32'h41ced349, 32'hc27904a9, 32'hc23c9e15, 32'h422a756c, 32'hc2a24495, 32'h41839bcc, 32'h424a9871};
test_output[1520] = '{32'h4263c75e};
test_index[1520] = '{0};
test_input[12168:12175] = '{32'hc29b7767, 32'h42c5688e, 32'h4186a0f4, 32'hc230fdd4, 32'h4264730c, 32'h41b46763, 32'h412d2dd9, 32'h429e893d};
test_output[1521] = '{32'h42c5688e};
test_index[1521] = '{1};
test_input[12176:12183] = '{32'hc160a96f, 32'h429cf629, 32'h42c6b2d2, 32'hc0e3f883, 32'hc297b2f7, 32'h4208b71e, 32'h42671ccc, 32'hc27613de};
test_output[1522] = '{32'h42c6b2d2};
test_index[1522] = '{2};
test_input[12184:12191] = '{32'hc254186e, 32'h42b72bda, 32'hc1c9138b, 32'h429ec873, 32'h4222d7e7, 32'h3f70fca2, 32'hc23ab0f7, 32'h42256a69};
test_output[1523] = '{32'h42b72bda};
test_index[1523] = '{1};
test_input[12192:12199] = '{32'hc2bc0040, 32'hc18ad0c9, 32'h42acc9b1, 32'h4298288c, 32'h4289a9d6, 32'hc216429d, 32'hc1a2fd04, 32'h42b8bb17};
test_output[1524] = '{32'h42b8bb17};
test_index[1524] = '{7};
test_input[12200:12207] = '{32'h425f2bf1, 32'hc2101756, 32'hc2b56e14, 32'h42aeb618, 32'h41cd26a0, 32'hc223ef24, 32'h410f1877, 32'hc118e7b1};
test_output[1525] = '{32'h42aeb618};
test_index[1525] = '{3};
test_input[12208:12215] = '{32'hc20e066b, 32'hbf3097fe, 32'h41d63f91, 32'h4244a5ca, 32'h41c1de93, 32'hc2c7a09c, 32'h42708ded, 32'h41512301};
test_output[1526] = '{32'h42708ded};
test_index[1526] = '{6};
test_input[12216:12223] = '{32'hc2659793, 32'hbfe075d2, 32'hc232ab44, 32'h4005cedd, 32'h40f85c81, 32'hc26b2a0f, 32'h419ce3f3, 32'h429c8664};
test_output[1527] = '{32'h429c8664};
test_index[1527] = '{7};
test_input[12224:12231] = '{32'h42453a7f, 32'h41759d2d, 32'h427c9539, 32'h41f0fe55, 32'h4261451a, 32'hc160e016, 32'h40802c4e, 32'hc205b121};
test_output[1528] = '{32'h427c9539};
test_index[1528] = '{2};
test_input[12232:12239] = '{32'h422aafdf, 32'h41b3a9f5, 32'h3f6cd174, 32'hc294eabb, 32'h42947920, 32'hc1e6f76d, 32'hc2c70bf2, 32'hc28699de};
test_output[1529] = '{32'h42947920};
test_index[1529] = '{4};
test_input[12240:12247] = '{32'hc25b02c9, 32'h4202f41a, 32'hc2a858cb, 32'hc2b0a7e2, 32'hc1db713c, 32'h429e39cd, 32'hc20994a4, 32'hc2b79373};
test_output[1530] = '{32'h429e39cd};
test_index[1530] = '{5};
test_input[12248:12255] = '{32'h42a757dc, 32'hc287ab8c, 32'h41418b28, 32'h41403e6c, 32'h420d3f2f, 32'hc205fb51, 32'hc1f36bef, 32'hc2852365};
test_output[1531] = '{32'h42a757dc};
test_index[1531] = '{0};
test_input[12256:12263] = '{32'hc1984a5c, 32'hc2813d26, 32'h42bc869a, 32'h421e67cf, 32'hc0a4c242, 32'hc28b1f93, 32'h421eac51, 32'hc2ba69ec};
test_output[1532] = '{32'h42bc869a};
test_index[1532] = '{2};
test_input[12264:12271] = '{32'h41c91b2e, 32'h410fd9e4, 32'h417960b3, 32'h429c9ff4, 32'h4203923c, 32'hc24a6d14, 32'h41fe5292, 32'hc22e3538};
test_output[1533] = '{32'h429c9ff4};
test_index[1533] = '{3};
test_input[12272:12279] = '{32'h42143b7e, 32'hc1585b18, 32'hc21a9721, 32'hc295fd08, 32'hc1a24a87, 32'h42c41b85, 32'hc14aab75, 32'h42a55aac};
test_output[1534] = '{32'h42c41b85};
test_index[1534] = '{5};
test_input[12280:12287] = '{32'hc1df1541, 32'h42b53a5c, 32'hc2477e95, 32'h42c25e4f, 32'h41cb90ec, 32'hc24c4aa0, 32'h41bead9a, 32'h420ee426};
test_output[1535] = '{32'h42c25e4f};
test_index[1535] = '{3};
test_input[12288:12295] = '{32'hc2104565, 32'hc287f4c5, 32'hc2a618ee, 32'hc06813de, 32'h42b65c16, 32'h41445119, 32'h42bfdeba, 32'h4298d62f};
test_output[1536] = '{32'h42bfdeba};
test_index[1536] = '{6};
test_input[12296:12303] = '{32'h42c2ef4e, 32'hc205db47, 32'h40f40a8f, 32'h42b9367d, 32'h421598aa, 32'hc241ef0a, 32'h4219a412, 32'h4228af24};
test_output[1537] = '{32'h42c2ef4e};
test_index[1537] = '{0};
test_input[12304:12311] = '{32'hc1b601a0, 32'hc2a61f4a, 32'h421f2363, 32'h403db03a, 32'hc2bdc108, 32'h42813299, 32'h42b26557, 32'h42417e09};
test_output[1538] = '{32'h42b26557};
test_index[1538] = '{6};
test_input[12312:12319] = '{32'hc29810ca, 32'h41ac5e43, 32'h4160b93d, 32'hc2b54948, 32'hc09761a2, 32'h42951705, 32'h42bccce1, 32'hc2a7733d};
test_output[1539] = '{32'h42bccce1};
test_index[1539] = '{6};
test_input[12320:12327] = '{32'h419234e2, 32'hc220cd65, 32'hc2345503, 32'hc288c76e, 32'h411d53ac, 32'h41dfad37, 32'hc1d16f47, 32'hc2b37109};
test_output[1540] = '{32'h41dfad37};
test_index[1540] = '{5};
test_input[12328:12335] = '{32'h426ddbdf, 32'h3f360a18, 32'h41a9897d, 32'h4260f51d, 32'hc1c31b54, 32'h42a30d89, 32'h421c0a5f, 32'hc23c33de};
test_output[1541] = '{32'h42a30d89};
test_index[1541] = '{5};
test_input[12336:12343] = '{32'h426e2b9f, 32'hc242f517, 32'hc1beb624, 32'hc2378850, 32'hc05d2a6c, 32'hc2a102d1, 32'hc24df3c3, 32'h41d76266};
test_output[1542] = '{32'h426e2b9f};
test_index[1542] = '{0};
test_input[12344:12351] = '{32'hc24e52c4, 32'h429d4755, 32'h41ac24b3, 32'h41d41aa8, 32'h41f8da2b, 32'h424d51c0, 32'h41f31ed8, 32'h42c4adc2};
test_output[1543] = '{32'h42c4adc2};
test_index[1543] = '{7};
test_input[12352:12359] = '{32'hc25765ad, 32'h42961ede, 32'hc1d6a9e9, 32'hc2870c64, 32'h407a28bb, 32'hc1b3a56e, 32'hc28c7e19, 32'h42900a39};
test_output[1544] = '{32'h42961ede};
test_index[1544] = '{1};
test_input[12360:12367] = '{32'h40c30651, 32'h42c122f1, 32'h42b90778, 32'h41ed840c, 32'hc220aa7e, 32'hc293c1d7, 32'h429cc34d, 32'h4287d4d9};
test_output[1545] = '{32'h42c122f1};
test_index[1545] = '{1};
test_input[12368:12375] = '{32'h42950448, 32'h41bfcec8, 32'hc2c4bfc5, 32'h41ca686d, 32'h428dfaa6, 32'hc284c088, 32'h3f50192d, 32'hc1bdb1f9};
test_output[1546] = '{32'h42950448};
test_index[1546] = '{0};
test_input[12376:12383] = '{32'h41c7d53e, 32'h42b52526, 32'hbfb99bf4, 32'hc28c3912, 32'h41d8f47b, 32'h419f0a1c, 32'h42a13259, 32'hc29e2279};
test_output[1547] = '{32'h42b52526};
test_index[1547] = '{1};
test_input[12384:12391] = '{32'hc1603ace, 32'hc0d13dd6, 32'hc29dc3da, 32'hbfd54ab2, 32'h428b348c, 32'hc2b8ee56, 32'h423750a8, 32'hc2947169};
test_output[1548] = '{32'h428b348c};
test_index[1548] = '{4};
test_input[12392:12399] = '{32'h42c007cc, 32'h42a4b94d, 32'h426817bd, 32'hc178b5d3, 32'h4299e348, 32'h41615b3f, 32'hc243271b, 32'h415646a2};
test_output[1549] = '{32'h42c007cc};
test_index[1549] = '{0};
test_input[12400:12407] = '{32'h4276aada, 32'hc2118126, 32'hc27eb11b, 32'h41da2086, 32'hc10c71dd, 32'hc1bc75f2, 32'h42018fa6, 32'h40aaedfb};
test_output[1550] = '{32'h4276aada};
test_index[1550] = '{0};
test_input[12408:12415] = '{32'h428d84f8, 32'h424bfd67, 32'h41cf41a7, 32'hc2aee794, 32'hc2812525, 32'h42021e10, 32'h40ecf42b, 32'h41f5e044};
test_output[1551] = '{32'h428d84f8};
test_index[1551] = '{0};
test_input[12416:12423] = '{32'hc18ed8a7, 32'h42435529, 32'h42725d9e, 32'h429d31de, 32'hc2c21646, 32'h4285f89f, 32'hc1bb9b48, 32'h40f86b34};
test_output[1552] = '{32'h429d31de};
test_index[1552] = '{3};
test_input[12424:12431] = '{32'h41e63c79, 32'h4203c70a, 32'h3facbe1d, 32'hc22e5b77, 32'hc255a3d9, 32'h41cb4461, 32'h421bd913, 32'h42c48144};
test_output[1553] = '{32'h42c48144};
test_index[1553] = '{7};
test_input[12432:12439] = '{32'h42b1caa7, 32'h40c7a95e, 32'hc283220f, 32'hc1fc8d3a, 32'hc1b092e7, 32'h40bf0c5d, 32'h4292fa7c, 32'hc0a24a32};
test_output[1554] = '{32'h42b1caa7};
test_index[1554] = '{0};
test_input[12440:12447] = '{32'hc2c65879, 32'hc29f8d40, 32'hc0bde3c7, 32'h41f09dbc, 32'hc289e9da, 32'h416145d4, 32'hc1e0362c, 32'h429189b9};
test_output[1555] = '{32'h429189b9};
test_index[1555] = '{7};
test_input[12448:12455] = '{32'h42135808, 32'hc25a32da, 32'hc1c1401a, 32'h42c6ecb8, 32'hc29c7206, 32'hc2497543, 32'h42bb49b5, 32'hc287d362};
test_output[1556] = '{32'h42c6ecb8};
test_index[1556] = '{3};
test_input[12456:12463] = '{32'hc255e9c8, 32'hc25a671c, 32'hc13993ec, 32'hc112c3d3, 32'h4287628f, 32'hc2648953, 32'hc15be3d3, 32'hc26b2685};
test_output[1557] = '{32'h4287628f};
test_index[1557] = '{4};
test_input[12464:12471] = '{32'h429687b4, 32'h42afb7ef, 32'hc2715914, 32'h425b034f, 32'hc0a6eef6, 32'hc1aa1a92, 32'h4286fc23, 32'hc0af2e04};
test_output[1558] = '{32'h42afb7ef};
test_index[1558] = '{1};
test_input[12472:12479] = '{32'h41a66a03, 32'h41ef96d2, 32'h428b8264, 32'hc2263021, 32'h4214df24, 32'hc1eeb896, 32'h427568c0, 32'h416ab29b};
test_output[1559] = '{32'h428b8264};
test_index[1559] = '{2};
test_input[12480:12487] = '{32'h41a89529, 32'hc22d28da, 32'h4282e3bc, 32'hc28b31ad, 32'hbebb55da, 32'h42b3a5ca, 32'hc1e2daaa, 32'h42af64de};
test_output[1560] = '{32'h42b3a5ca};
test_index[1560] = '{5};
test_input[12488:12495] = '{32'hc264ece8, 32'hc1f7cd2a, 32'hc2611ce3, 32'hc1d781ad, 32'hc2142f33, 32'hc278f468, 32'hc27f46b6, 32'h420d5b92};
test_output[1561] = '{32'h420d5b92};
test_index[1561] = '{7};
test_input[12496:12503] = '{32'h42acf0b0, 32'hc27e46db, 32'hc2af081e, 32'hc2bdc0b3, 32'hc29079d1, 32'hc2684cd0, 32'hc253b5c1, 32'hc2956e94};
test_output[1562] = '{32'h42acf0b0};
test_index[1562] = '{0};
test_input[12504:12511] = '{32'h42a635cc, 32'h40b20ce6, 32'hc1c9a411, 32'h429106fe, 32'h42843004, 32'hc1f78f5f, 32'hc1e12935, 32'h427d0a6a};
test_output[1563] = '{32'h42a635cc};
test_index[1563] = '{0};
test_input[12512:12519] = '{32'h42be33da, 32'hc2be1af0, 32'h42b9a3e2, 32'hc28c78d7, 32'h423c3fa6, 32'hc26211c8, 32'h42a1cb5b, 32'h42a67d0f};
test_output[1564] = '{32'h42be33da};
test_index[1564] = '{0};
test_input[12520:12527] = '{32'hc24fda0d, 32'hc2ae88da, 32'h42867000, 32'h41af732f, 32'hc28dd57b, 32'hc26f6e07, 32'hc2a41e80, 32'hc2208186};
test_output[1565] = '{32'h42867000};
test_index[1565] = '{2};
test_input[12528:12535] = '{32'hc1bb6853, 32'h426f7f56, 32'hc1ba116d, 32'h41205f17, 32'h42147a22, 32'h41dc7d49, 32'hc1a17dac, 32'h407e0498};
test_output[1566] = '{32'h426f7f56};
test_index[1566] = '{1};
test_input[12536:12543] = '{32'h42976bbb, 32'h4229ea40, 32'h42a56fb4, 32'hc29aaa69, 32'h4221d3dd, 32'h40ed89ff, 32'h41dbc47c, 32'h42746302};
test_output[1567] = '{32'h42a56fb4};
test_index[1567] = '{2};
test_input[12544:12551] = '{32'hc2abd6b9, 32'hc2ad1759, 32'hc2a024af, 32'hc2a571be, 32'h42701123, 32'h41d5e841, 32'h42829340, 32'h41f4a5e0};
test_output[1568] = '{32'h42829340};
test_index[1568] = '{6};
test_input[12552:12559] = '{32'hc1dd6217, 32'hc205c4d2, 32'h42bb2646, 32'h412875b2, 32'hc2a26715, 32'h42be9ea3, 32'hc2b06f70, 32'hc2a2eb40};
test_output[1569] = '{32'h42be9ea3};
test_index[1569] = '{5};
test_input[12560:12567] = '{32'h42adac53, 32'hc1855a6c, 32'h4247bbf8, 32'h416031a7, 32'h41b1170d, 32'hc286b52d, 32'hc1073657, 32'h41fc9549};
test_output[1570] = '{32'h42adac53};
test_index[1570] = '{0};
test_input[12568:12575] = '{32'h418ccecc, 32'h417541c3, 32'hc184fa1a, 32'h42ba0a0b, 32'h425f847b, 32'hc2be42f8, 32'h4289b924, 32'h419f3940};
test_output[1571] = '{32'h42ba0a0b};
test_index[1571] = '{3};
test_input[12576:12583] = '{32'hc2b12d24, 32'hc17708ff, 32'hc2055864, 32'h4296224d, 32'h41606809, 32'hc0de30ea, 32'hc2b45372, 32'h42408272};
test_output[1572] = '{32'h4296224d};
test_index[1572] = '{3};
test_input[12584:12591] = '{32'h42c10d89, 32'hc228289d, 32'h4188af6e, 32'hc1b47b02, 32'h41d847a1, 32'hc241d4c4, 32'hc1a9cb78, 32'hc27e8c65};
test_output[1573] = '{32'h42c10d89};
test_index[1573] = '{0};
test_input[12592:12599] = '{32'hc20aac02, 32'hc1c60a73, 32'h42c497ca, 32'hc2950e8a, 32'h42b0bcae, 32'hc2b639eb, 32'h4206b55f, 32'h42a3bd94};
test_output[1574] = '{32'h42c497ca};
test_index[1574] = '{2};
test_input[12600:12607] = '{32'h42aa5aa2, 32'h4201fd81, 32'h3f81da2e, 32'h418094d4, 32'hc23766a4, 32'h4188b8f8, 32'hc2c50fa0, 32'h4271fa2f};
test_output[1575] = '{32'h42aa5aa2};
test_index[1575] = '{0};
test_input[12608:12615] = '{32'h40cfb9d1, 32'h4271f2d5, 32'h429de830, 32'hc1bd2809, 32'hc2238f09, 32'hc1bc6654, 32'h41d8096d, 32'h419e64b0};
test_output[1576] = '{32'h429de830};
test_index[1576] = '{2};
test_input[12616:12623] = '{32'hc202d129, 32'h42216b91, 32'h429348ad, 32'h428f532a, 32'hc1897559, 32'h4166c3fb, 32'hc276981d, 32'h429ed5e9};
test_output[1577] = '{32'h429ed5e9};
test_index[1577] = '{7};
test_input[12624:12631] = '{32'h41e526bd, 32'hc2126824, 32'h4200598a, 32'h41f03c3b, 32'hc1cabe9e, 32'hc28f6b21, 32'hc19556cd, 32'h42af20a9};
test_output[1578] = '{32'h42af20a9};
test_index[1578] = '{7};
test_input[12632:12639] = '{32'h41a81320, 32'hc2bc802b, 32'h41f86a3c, 32'h42750c2e, 32'h41efcaac, 32'h41dfda38, 32'h42c1cc14, 32'h40b245ba};
test_output[1579] = '{32'h42c1cc14};
test_index[1579] = '{6};
test_input[12640:12647] = '{32'h427429c6, 32'hc298eca9, 32'h409501a0, 32'h421398d2, 32'hc1c2b628, 32'hc28d11d1, 32'h4297e7ec, 32'hc2a3935c};
test_output[1580] = '{32'h4297e7ec};
test_index[1580] = '{6};
test_input[12648:12655] = '{32'h412fb57e, 32'h420f9e92, 32'h40bdfeb3, 32'h42c7d1b6, 32'hc2177b67, 32'h4297bee9, 32'h425cde45, 32'hc25bb781};
test_output[1581] = '{32'h42c7d1b6};
test_index[1581] = '{3};
test_input[12656:12663] = '{32'hc27c1d9c, 32'hc1f99d53, 32'hc2967868, 32'hc2aba743, 32'hc180b752, 32'hc22a5f15, 32'h42419d17, 32'hc2a727b2};
test_output[1582] = '{32'h42419d17};
test_index[1582] = '{6};
test_input[12664:12671] = '{32'hc2a21a8a, 32'hc1efd2c1, 32'h41c94117, 32'hc2347990, 32'hc29781d2, 32'h421d75f8, 32'hc2a6f52b, 32'hc1ddd50e};
test_output[1583] = '{32'h421d75f8};
test_index[1583] = '{5};
test_input[12672:12679] = '{32'h422a67e6, 32'hc268c5c4, 32'hc1751379, 32'h41ca6654, 32'h414d4b5a, 32'h42c17cd6, 32'h4286ff28, 32'hc274a4cd};
test_output[1584] = '{32'h42c17cd6};
test_index[1584] = '{5};
test_input[12680:12687] = '{32'h41ef88fb, 32'h412e835a, 32'hc26be995, 32'hc165b030, 32'hc278ae9b, 32'h4265ff20, 32'hc168071f, 32'h422f396a};
test_output[1585] = '{32'h4265ff20};
test_index[1585] = '{5};
test_input[12688:12695] = '{32'hc19be054, 32'h429ec061, 32'h42832189, 32'h41a29abf, 32'h42b5896e, 32'hc2813ccb, 32'h429ad5b0, 32'hc1e147b7};
test_output[1586] = '{32'h42b5896e};
test_index[1586] = '{4};
test_input[12696:12703] = '{32'h42a4ff6f, 32'h4265f569, 32'h41dfe260, 32'h42bc73d5, 32'h40c156b4, 32'h41afb1a9, 32'h41aa964e, 32'hc1adc91d};
test_output[1587] = '{32'h42bc73d5};
test_index[1587] = '{3};
test_input[12704:12711] = '{32'h41b36548, 32'h424d809f, 32'h422d476a, 32'h40820866, 32'hc19b7246, 32'h41c82e69, 32'h42a836d5, 32'h429c47f6};
test_output[1588] = '{32'h42a836d5};
test_index[1588] = '{6};
test_input[12712:12719] = '{32'h42537ff6, 32'hc297eee0, 32'hc20e9057, 32'hc0601cdf, 32'hc2363798, 32'h42c6d231, 32'hc2210df0, 32'hc2b7d087};
test_output[1589] = '{32'h42c6d231};
test_index[1589] = '{5};
test_input[12720:12727] = '{32'hc20a90b5, 32'h42824609, 32'hc285b322, 32'h40925def, 32'hc183365d, 32'hc19f950e, 32'h417ebf58, 32'h4239703d};
test_output[1590] = '{32'h42824609};
test_index[1590] = '{1};
test_input[12728:12735] = '{32'h4292dd85, 32'hc2c36f11, 32'hc20a4d31, 32'h41cba20f, 32'hc1a79682, 32'h41bb26d8, 32'h422473dd, 32'hc29610cb};
test_output[1591] = '{32'h4292dd85};
test_index[1591] = '{0};
test_input[12736:12743] = '{32'h421513c1, 32'hc2988bdf, 32'hc2994415, 32'h4269089b, 32'hc2b37604, 32'hc24693fb, 32'h4288ea82, 32'h423b9e34};
test_output[1592] = '{32'h4288ea82};
test_index[1592] = '{6};
test_input[12744:12751] = '{32'hc2c19e12, 32'h42b6ebad, 32'hc29bb738, 32'hc1e01311, 32'hc132eb3f, 32'hbfdcf67a, 32'hc0c16efa, 32'hc2760507};
test_output[1593] = '{32'h42b6ebad};
test_index[1593] = '{1};
test_input[12752:12759] = '{32'hc289855c, 32'hc22bb1e6, 32'h424e8a72, 32'h4191dc6c, 32'hc19abb3f, 32'h42874267, 32'hc28993ba, 32'h42566839};
test_output[1594] = '{32'h42874267};
test_index[1594] = '{5};
test_input[12760:12767] = '{32'h41522855, 32'hc2a7ded3, 32'hc24e74b5, 32'h42c406b4, 32'hc0dfa54f, 32'h421ddc7c, 32'hc27e7f88, 32'h4206400b};
test_output[1595] = '{32'h42c406b4};
test_index[1595] = '{3};
test_input[12768:12775] = '{32'hc12fce63, 32'h42974b89, 32'hc15f94d1, 32'h421a5ba3, 32'hc22404e4, 32'h40882178, 32'hc1308052, 32'hc2b3921e};
test_output[1596] = '{32'h42974b89};
test_index[1596] = '{1};
test_input[12776:12783] = '{32'h4217c532, 32'hc28c4287, 32'hc2601ee4, 32'h41f4b78c, 32'h426e75cc, 32'hc214e2ec, 32'h42a88435, 32'hc202e9b6};
test_output[1597] = '{32'h42a88435};
test_index[1597] = '{6};
test_input[12784:12791] = '{32'h42b563b6, 32'hc27882b5, 32'h41e2526e, 32'hc1effd2f, 32'hc1e4de99, 32'h409585fd, 32'hc1bfed6f, 32'h42bffbce};
test_output[1598] = '{32'h42bffbce};
test_index[1598] = '{7};
test_input[12792:12799] = '{32'hc27da777, 32'hc02a7ebe, 32'hc2b9baba, 32'h41b03893, 32'h41d5e333, 32'hc2352b1d, 32'hc21a4f2a, 32'h42c3c88a};
test_output[1599] = '{32'h42c3c88a};
test_index[1599] = '{7};
test_input[12800:12807] = '{32'h429eda8e, 32'hc2b48148, 32'hc20433ac, 32'h42882313, 32'hc14076b2, 32'h416a5e70, 32'h42ab09c6, 32'hc2901676};
test_output[1600] = '{32'h42ab09c6};
test_index[1600] = '{6};
test_input[12808:12815] = '{32'h42383eb3, 32'hc267f1dc, 32'h42944167, 32'h4283828e, 32'hc1d3c818, 32'h42bc1c25, 32'hc13970e2, 32'hc25c3db3};
test_output[1601] = '{32'h42bc1c25};
test_index[1601] = '{5};
test_input[12816:12823] = '{32'hc2824fab, 32'hc25d9fc1, 32'h426fd336, 32'hc2c09569, 32'hc21c1fab, 32'hc2a31a1d, 32'h42c369ae, 32'h41ba4503};
test_output[1602] = '{32'h42c369ae};
test_index[1602] = '{6};
test_input[12824:12831] = '{32'h407da444, 32'hc22cce25, 32'h41931c5f, 32'hc2903d52, 32'h41597d17, 32'hc2be59d2, 32'hc2bc0ca6, 32'hc28927ef};
test_output[1603] = '{32'h41931c5f};
test_index[1603] = '{2};
test_input[12832:12839] = '{32'h41b24c7e, 32'hc0c0e641, 32'h4221d6d9, 32'hc2a0451f, 32'h42bd1696, 32'h41615fe6, 32'h42c64ceb, 32'hc1fcd215};
test_output[1604] = '{32'h42c64ceb};
test_index[1604] = '{6};
test_input[12840:12847] = '{32'h4283bb73, 32'h425a9a83, 32'hc170f5cc, 32'hc22e63dd, 32'hc2819c44, 32'hc2284a78, 32'hc295dfba, 32'hc24da90f};
test_output[1605] = '{32'h4283bb73};
test_index[1605] = '{0};
test_input[12848:12855] = '{32'h41f784ae, 32'h41a37555, 32'h41b255ae, 32'h42c2d95f, 32'h4239a386, 32'hc23a4a46, 32'hc1ceed64, 32'hc0ff872e};
test_output[1606] = '{32'h42c2d95f};
test_index[1606] = '{3};
test_input[12856:12863] = '{32'h40f79f89, 32'h429eb07d, 32'hc20cf749, 32'hc2a428d6, 32'h40582dcb, 32'h4223effd, 32'h41ccbef3, 32'hc2192e05};
test_output[1607] = '{32'h429eb07d};
test_index[1607] = '{1};
test_input[12864:12871] = '{32'hc2c7f075, 32'hc09ed664, 32'hc2907601, 32'h418eb16e, 32'h426d6ef7, 32'hc0fe010c, 32'hc23dc715, 32'h418e58af};
test_output[1608] = '{32'h426d6ef7};
test_index[1608] = '{4};
test_input[12872:12879] = '{32'h42a64f41, 32'hc291968b, 32'hc185cfaf, 32'h42c37b93, 32'hc2841110, 32'h41ceaafa, 32'hc26c3148, 32'h426fcb64};
test_output[1609] = '{32'h42c37b93};
test_index[1609] = '{3};
test_input[12880:12887] = '{32'h4167c4f6, 32'h424e2e51, 32'h3f555b5d, 32'hc294466b, 32'hc20fb4f6, 32'h42a410b3, 32'hc1ce47e4, 32'hc2a55e4b};
test_output[1610] = '{32'h42a410b3};
test_index[1610] = '{5};
test_input[12888:12895] = '{32'hc28920bf, 32'hc2a9b619, 32'h42829c44, 32'h4269d9d7, 32'hc2c36b8b, 32'h42a2a45a, 32'hc14f3a4f, 32'hc1715475};
test_output[1611] = '{32'h42a2a45a};
test_index[1611] = '{5};
test_input[12896:12903] = '{32'hc2a1162d, 32'h421590d1, 32'h429368dd, 32'hc0c744e4, 32'hc2bd543b, 32'hc295f95a, 32'h42c4e947, 32'h428d21b1};
test_output[1612] = '{32'h42c4e947};
test_index[1612] = '{6};
test_input[12904:12911] = '{32'h4273cb25, 32'h42c02905, 32'h428b933d, 32'h4281bfcf, 32'h41f90636, 32'hc2aebeab, 32'h42a42190, 32'h42c59f26};
test_output[1613] = '{32'h42c59f26};
test_index[1613] = '{7};
test_input[12912:12919] = '{32'hc0ce4a2b, 32'hc1553f87, 32'hc29cffa8, 32'h4161f3ff, 32'hc22aa5b7, 32'h42226adf, 32'h421e3478, 32'hc1c501ad};
test_output[1614] = '{32'h42226adf};
test_index[1614] = '{5};
test_input[12920:12927] = '{32'h41caee17, 32'h42bcf113, 32'hc2a2b43d, 32'h419a4aab, 32'h4295f716, 32'hbe75b355, 32'h423a69af, 32'hc1c0d111};
test_output[1615] = '{32'h42bcf113};
test_index[1615] = '{1};
test_input[12928:12935] = '{32'h3fb1bf2b, 32'hc2b29c64, 32'hc2b04705, 32'hc18439ae, 32'h42a24fcb, 32'h42c34656, 32'h411d8477, 32'hc0f2808a};
test_output[1616] = '{32'h42c34656};
test_index[1616] = '{5};
test_input[12936:12943] = '{32'h428faec5, 32'hc251aa29, 32'hc28f7834, 32'hc2932052, 32'h42891387, 32'h422f2ca3, 32'hc204e83b, 32'h4289371d};
test_output[1617] = '{32'h428faec5};
test_index[1617] = '{0};
test_input[12944:12951] = '{32'hbf81e3a7, 32'hc16bf3c1, 32'hc2ad5437, 32'hc27d2bd5, 32'hc2b0badc, 32'hc1bed82b, 32'hc2a79e35, 32'hc215a230};
test_output[1618] = '{32'hbf81e3a7};
test_index[1618] = '{0};
test_input[12952:12959] = '{32'hc26eb22e, 32'hc20b4363, 32'hc29a5686, 32'hc20ba033, 32'h42b369c0, 32'hc1e22969, 32'h42adbaad, 32'hc28e935e};
test_output[1619] = '{32'h42b369c0};
test_index[1619] = '{4};
test_input[12960:12967] = '{32'h41091dc2, 32'hc22cbb79, 32'hc09dc18e, 32'h40080ddb, 32'hc29110bd, 32'hc251da3c, 32'h4273098a, 32'h42a8857f};
test_output[1620] = '{32'h42a8857f};
test_index[1620] = '{7};
test_input[12968:12975] = '{32'hc20c2236, 32'hc23644ef, 32'h4219e9cc, 32'hc2bb5fd5, 32'h417e8abd, 32'hc296626f, 32'h4290706f, 32'hbfb5588c};
test_output[1621] = '{32'h4290706f};
test_index[1621] = '{6};
test_input[12976:12983] = '{32'hc2ad3442, 32'hc2abbeda, 32'hc238e986, 32'h41573028, 32'hc2a9dc14, 32'h4271448b, 32'h42668aef, 32'h4120191c};
test_output[1622] = '{32'h4271448b};
test_index[1622] = '{5};
test_input[12984:12991] = '{32'h429be4cb, 32'h422c49e9, 32'h41f24994, 32'hc294d8b9, 32'hc29a5945, 32'hc20f3143, 32'h418ff0aa, 32'hc25da19b};
test_output[1623] = '{32'h429be4cb};
test_index[1623] = '{0};
test_input[12992:12999] = '{32'h41b69a9b, 32'hc1eed4e7, 32'h422a8f38, 32'h41690409, 32'h420db63d, 32'h42652fc4, 32'h428d416b, 32'hc19f8ebf};
test_output[1624] = '{32'h428d416b};
test_index[1624] = '{6};
test_input[13000:13007] = '{32'hc27b5312, 32'hc1fa2f08, 32'hc239a41f, 32'hc2c2794f, 32'hc117d033, 32'h403859d1, 32'h416a8c60, 32'h42b99fb4};
test_output[1625] = '{32'h42b99fb4};
test_index[1625] = '{7};
test_input[13008:13015] = '{32'hc25f0dbd, 32'hc14ba34a, 32'h40a6822b, 32'hc289c47b, 32'h41840595, 32'hc1b04ddf, 32'h429b9c2c, 32'h42c1b28c};
test_output[1626] = '{32'h42c1b28c};
test_index[1626] = '{7};
test_input[13016:13023] = '{32'h42b2bf22, 32'hc2543612, 32'h4227db6b, 32'h421c972c, 32'h42be6bf5, 32'hc2b653b2, 32'hc2043b04, 32'h41bd415f};
test_output[1627] = '{32'h42be6bf5};
test_index[1627] = '{4};
test_input[13024:13031] = '{32'h428e1902, 32'hc16ecad3, 32'h42c241ff, 32'hc2ba79c9, 32'h42c16977, 32'h41ee6798, 32'hc162b577, 32'h42ac559b};
test_output[1628] = '{32'h42c241ff};
test_index[1628] = '{2};
test_input[13032:13039] = '{32'hc268f577, 32'hc0b4c004, 32'h400bc703, 32'hc1f44fab, 32'hc14539e9, 32'h420c3fcd, 32'h429c67eb, 32'h4230490a};
test_output[1629] = '{32'h429c67eb};
test_index[1629] = '{6};
test_input[13040:13047] = '{32'h42518332, 32'h42555cb9, 32'h4268046a, 32'h42c0f50f, 32'hc2bac564, 32'hc117fb2d, 32'h42a0ee9a, 32'hc2248917};
test_output[1630] = '{32'h42c0f50f};
test_index[1630] = '{3};
test_input[13048:13055] = '{32'h42a848c4, 32'hc036e7bf, 32'h421bb28c, 32'hc29c7d16, 32'hc2381f66, 32'hc1a50185, 32'h428a8be6, 32'h428a57f3};
test_output[1631] = '{32'h42a848c4};
test_index[1631] = '{0};
test_input[13056:13063] = '{32'h423f5f35, 32'hc2906c44, 32'h42ae20e7, 32'hbfbc0b47, 32'h42b2cff6, 32'hc24d275e, 32'h4254a235, 32'h42925f77};
test_output[1632] = '{32'h42b2cff6};
test_index[1632] = '{4};
test_input[13064:13071] = '{32'h42c78c5b, 32'hc228da7f, 32'hc2b30f71, 32'h42528139, 32'h4198ab9e, 32'h42910519, 32'hc2ad8a22, 32'h42a91b88};
test_output[1633] = '{32'h42c78c5b};
test_index[1633] = '{0};
test_input[13072:13079] = '{32'hc29c8690, 32'h4288b994, 32'h429853b5, 32'h41f6ca15, 32'h4168e236, 32'hc15fce9a, 32'hc196e30d, 32'h4238bbc8};
test_output[1634] = '{32'h429853b5};
test_index[1634] = '{2};
test_input[13080:13087] = '{32'h423f0d14, 32'h3f7baff9, 32'h42586681, 32'hc2b023b7, 32'hc2aa835f, 32'hc2a21375, 32'h424f95eb, 32'hc1ed0928};
test_output[1635] = '{32'h42586681};
test_index[1635] = '{2};
test_input[13088:13095] = '{32'hc2859b7d, 32'hc2bb691e, 32'h42b514bb, 32'hc24d0a69, 32'hc1ded8b0, 32'h42a18ca6, 32'h42c604ca, 32'h40fcfcc8};
test_output[1636] = '{32'h42c604ca};
test_index[1636] = '{6};
test_input[13096:13103] = '{32'h4294d176, 32'h428bd7b4, 32'hc280913d, 32'h42852799, 32'hc1d67c6a, 32'h42a24e7b, 32'hc2420ca2, 32'hc2a75148};
test_output[1637] = '{32'h42a24e7b};
test_index[1637] = '{5};
test_input[13104:13111] = '{32'h42c2d1ce, 32'h42a65a6c, 32'h42bf8017, 32'hc1fbc2cb, 32'hc29ed11f, 32'hc1849364, 32'h40b6b2c5, 32'hc204f241};
test_output[1638] = '{32'h42c2d1ce};
test_index[1638] = '{0};
test_input[13112:13119] = '{32'h4169ba3b, 32'h42b6cc18, 32'h42b0a3b7, 32'h4296a05f, 32'h427629bf, 32'hc242de4d, 32'h42124876, 32'hc2b6cf60};
test_output[1639] = '{32'h42b6cc18};
test_index[1639] = '{1};
test_input[13120:13127] = '{32'hc2508127, 32'hc246f3dd, 32'h42c7bfb8, 32'h41500116, 32'hc1c8b765, 32'h423bfa46, 32'h429ae3ff, 32'hc2199c86};
test_output[1640] = '{32'h42c7bfb8};
test_index[1640] = '{2};
test_input[13128:13135] = '{32'h41cdbc32, 32'hc1245b50, 32'hc2a0c8bc, 32'hc201545f, 32'hc292d237, 32'h41d94232, 32'h42963866, 32'hc194afa1};
test_output[1641] = '{32'h42963866};
test_index[1641] = '{6};
test_input[13136:13143] = '{32'h42a976b0, 32'h42406fd8, 32'h42a4da70, 32'h4288efd4, 32'h4169d139, 32'h429da28f, 32'hc2a5f72a, 32'hc2395e01};
test_output[1642] = '{32'h42a976b0};
test_index[1642] = '{0};
test_input[13144:13151] = '{32'hc13baad1, 32'hc215972e, 32'hc2637ee0, 32'h423327e3, 32'hc11256ec, 32'hc1d3690c, 32'h427e9bc3, 32'h4260f818};
test_output[1643] = '{32'h427e9bc3};
test_index[1643] = '{6};
test_input[13152:13159] = '{32'h42a0f4a0, 32'hc2b10365, 32'h42ba5403, 32'hc22fd9f8, 32'hc2abbbb9, 32'h4243fdae, 32'hc288615c, 32'hc2af2d18};
test_output[1644] = '{32'h42ba5403};
test_index[1644] = '{2};
test_input[13160:13167] = '{32'h426baa98, 32'h42bc8b15, 32'h427dac15, 32'hc28ca009, 32'h421496e8, 32'hc29e5a39, 32'h42ae190b, 32'h42156469};
test_output[1645] = '{32'h42bc8b15};
test_index[1645] = '{1};
test_input[13168:13175] = '{32'hc2c4e227, 32'h4200f7bf, 32'h41929fbf, 32'hc27df959, 32'hc25f059d, 32'hc1a42a56, 32'h42884b54, 32'h41107e73};
test_output[1646] = '{32'h42884b54};
test_index[1646] = '{6};
test_input[13176:13183] = '{32'hc2aa56ba, 32'hc2707052, 32'hc192a8a9, 32'hc2b4daf0, 32'h41cba005, 32'h4241b390, 32'h423df25c, 32'hc25bb087};
test_output[1647] = '{32'h4241b390};
test_index[1647] = '{5};
test_input[13184:13191] = '{32'hc189e856, 32'hc282aed8, 32'h41ac4920, 32'h4243fb6a, 32'h41816f3e, 32'hc2c7463b, 32'hc2a666ca, 32'h419c273e};
test_output[1648] = '{32'h4243fb6a};
test_index[1648] = '{3};
test_input[13192:13199] = '{32'hc2822196, 32'hc2c1e08a, 32'h42252d99, 32'h41b68d42, 32'h4223dd5a, 32'hc2a312cf, 32'hc29020a1, 32'h429cf3d8};
test_output[1649] = '{32'h429cf3d8};
test_index[1649] = '{7};
test_input[13200:13207] = '{32'h4251f4c9, 32'hc297fa86, 32'h42ab417e, 32'hc24f0b09, 32'h41827faf, 32'h4204f72e, 32'h42c46ba2, 32'h4296945b};
test_output[1650] = '{32'h42c46ba2};
test_index[1650] = '{6};
test_input[13208:13215] = '{32'hc1225a3b, 32'hc2424541, 32'hc0b5bcf6, 32'hc293e1de, 32'hc17a0b7c, 32'hc289fc5c, 32'hc141572e, 32'h4128aaee};
test_output[1651] = '{32'h4128aaee};
test_index[1651] = '{7};
test_input[13216:13223] = '{32'h4186362d, 32'h405aa698, 32'h42a1180b, 32'hc052b22d, 32'h413d8d23, 32'h426783e9, 32'h4283c7ed, 32'hc180b221};
test_output[1652] = '{32'h42a1180b};
test_index[1652] = '{2};
test_input[13224:13231] = '{32'h42a700c9, 32'h427639e3, 32'hc2592a23, 32'h42b12a8c, 32'h4231e8b8, 32'hc0894906, 32'hc2b23578, 32'h42ad15bb};
test_output[1653] = '{32'h42b12a8c};
test_index[1653] = '{3};
test_input[13232:13239] = '{32'hc28a0d5b, 32'h42a8f409, 32'hc1fb0d32, 32'hc24d848b, 32'hc14c61f9, 32'h41ea2d5a, 32'hbfad973b, 32'hc2c6a2d3};
test_output[1654] = '{32'h42a8f409};
test_index[1654] = '{1};
test_input[13240:13247] = '{32'hc150ba78, 32'h42283c4d, 32'h42bf92f1, 32'h4279c2e8, 32'h42421d0a, 32'hc1223f7e, 32'h429c237c, 32'hc18f797f};
test_output[1655] = '{32'h42bf92f1};
test_index[1655] = '{2};
test_input[13248:13255] = '{32'hc174a3ba, 32'h42b4dbc2, 32'h4284787e, 32'hc23bcd4f, 32'hc19fd78d, 32'h41a75fcc, 32'hc105a4fd, 32'h429c0b5f};
test_output[1656] = '{32'h42b4dbc2};
test_index[1656] = '{1};
test_input[13256:13263] = '{32'hc296096e, 32'hc2867c05, 32'h42a53c06, 32'hc28ec106, 32'h428e8337, 32'h42b72925, 32'h42a637ab, 32'hc1f538e8};
test_output[1657] = '{32'h42b72925};
test_index[1657] = '{5};
test_input[13264:13271] = '{32'hbdb3f14b, 32'hc2b69483, 32'hc295fdb8, 32'hc1ec93c5, 32'hc21854a7, 32'hc25148e9, 32'hc20b6512, 32'hc2a77d35};
test_output[1658] = '{32'hbdb3f14b};
test_index[1658] = '{0};
test_input[13272:13279] = '{32'h42a104d1, 32'h4045e10d, 32'hc12bef75, 32'h4223cd33, 32'h42469dbe, 32'hc279bde2, 32'hc24ab0ae, 32'h401e8a6a};
test_output[1659] = '{32'h42a104d1};
test_index[1659] = '{0};
test_input[13280:13287] = '{32'h408c35d9, 32'hc0f82093, 32'h42085c6d, 32'hc2ac853f, 32'hc28cb5a5, 32'h428d385f, 32'h425c506d, 32'h425fb70f};
test_output[1660] = '{32'h428d385f};
test_index[1660] = '{5};
test_input[13288:13295] = '{32'hc28e83c5, 32'h421f3e25, 32'hc198a378, 32'h42685750, 32'h4116b490, 32'h428bdf9c, 32'hc29549f8, 32'h42058333};
test_output[1661] = '{32'h428bdf9c};
test_index[1661] = '{5};
test_input[13296:13303] = '{32'hc206d0d5, 32'hc29476be, 32'h42483af9, 32'hc1845c4e, 32'hc28f6629, 32'hc2277257, 32'h42969ea0, 32'hc1b70ab8};
test_output[1662] = '{32'h42969ea0};
test_index[1662] = '{6};
test_input[13304:13311] = '{32'hc28951f2, 32'hc0d11082, 32'h42670143, 32'h40bed87f, 32'hc1a97c97, 32'h41a7b4f3, 32'hc16bf92d, 32'h4248c946};
test_output[1663] = '{32'h42670143};
test_index[1663] = '{2};
test_input[13312:13319] = '{32'h42b18d18, 32'hc1c6fa42, 32'h4287be46, 32'hc2bedcae, 32'h411bc60b, 32'h4280d567, 32'h41b0edf6, 32'hc2404135};
test_output[1664] = '{32'h42b18d18};
test_index[1664] = '{0};
test_input[13320:13327] = '{32'h425e5adf, 32'hc2738447, 32'h42ab6058, 32'h423e9771, 32'hc2be61e6, 32'hc2a339cc, 32'h421d1036, 32'hc2a2ba59};
test_output[1665] = '{32'h42ab6058};
test_index[1665] = '{2};
test_input[13328:13335] = '{32'h429f0600, 32'hc2a63c53, 32'h42900b3a, 32'h41c8f8be, 32'hc2a5afba, 32'h40b5ee4e, 32'hc2ab4800, 32'h41e06d70};
test_output[1666] = '{32'h429f0600};
test_index[1666] = '{0};
test_input[13336:13343] = '{32'h42675e0a, 32'h4277121a, 32'hc27b31a3, 32'h4231e953, 32'hc10f6ecb, 32'h42866fce, 32'h40311203, 32'h4188849f};
test_output[1667] = '{32'h42866fce};
test_index[1667] = '{5};
test_input[13344:13351] = '{32'h42bafb48, 32'hc01cdc93, 32'hc2a74898, 32'hc2b968fa, 32'hc2a43bea, 32'hc24ea668, 32'hbf113ef7, 32'hc26708dd};
test_output[1668] = '{32'h42bafb48};
test_index[1668] = '{0};
test_input[13352:13359] = '{32'hc210b681, 32'hc1e6a11a, 32'h413ab691, 32'h418b922b, 32'h42836aec, 32'hc2284c54, 32'hc2591e01, 32'h427ab452};
test_output[1669] = '{32'h42836aec};
test_index[1669] = '{4};
test_input[13360:13367] = '{32'h40efd22d, 32'hc280ef01, 32'h42760bfc, 32'hc063ba19, 32'h4182d0b2, 32'h429c5e28, 32'h42a1774f, 32'h42951a20};
test_output[1670] = '{32'h42a1774f};
test_index[1670] = '{6};
test_input[13368:13375] = '{32'h41bbb56e, 32'hc132f99b, 32'hc2427905, 32'h4107b89b, 32'h42422af0, 32'h42904250, 32'hc28a19e0, 32'h4228bca3};
test_output[1671] = '{32'h42904250};
test_index[1671] = '{5};
test_input[13376:13383] = '{32'hc2abeecf, 32'h4122b1f6, 32'hc18f8d4d, 32'hc2246985, 32'h429c8565, 32'hc06a7e7b, 32'hc1e16f2f, 32'h42496f55};
test_output[1672] = '{32'h429c8565};
test_index[1672] = '{4};
test_input[13384:13391] = '{32'hc2273709, 32'h4222dea2, 32'h4256a1cf, 32'h41aa110f, 32'hc2af133c, 32'hc1f0935d, 32'h4190abc8, 32'hc1cdb16e};
test_output[1673] = '{32'h4256a1cf};
test_index[1673] = '{2};
test_input[13392:13399] = '{32'hc2766a78, 32'hc15cb31d, 32'hc2c50b95, 32'h41b7f954, 32'hc20fdb31, 32'h409cda04, 32'h41e15365, 32'hc28e8bb0};
test_output[1674] = '{32'h41e15365};
test_index[1674] = '{6};
test_input[13400:13407] = '{32'h42ae8ee7, 32'hc2976614, 32'h42a557c7, 32'hc273c390, 32'h42051a2b, 32'hbf8a4cbf, 32'h42c12bd4, 32'hc18d7306};
test_output[1675] = '{32'h42c12bd4};
test_index[1675] = '{6};
test_input[13408:13415] = '{32'h4180a3e8, 32'hc28c30f6, 32'hc1844185, 32'hc1c2eb0a, 32'hc2b19494, 32'hc2a4e6cc, 32'h425030a7, 32'h428f82d1};
test_output[1676] = '{32'h428f82d1};
test_index[1676] = '{7};
test_input[13416:13423] = '{32'h421ad347, 32'h42bacfc8, 32'hc1f650c2, 32'h42a31fe9, 32'hc2bb2038, 32'hc285c0ad, 32'hc26cd9c0, 32'hc276a1f5};
test_output[1677] = '{32'h42bacfc8};
test_index[1677] = '{1};
test_input[13424:13431] = '{32'hc2932fa0, 32'h42b74cc6, 32'h42c4b6d6, 32'h417537a1, 32'hc1fb4d61, 32'h42704521, 32'h4152c180, 32'h418eaaf0};
test_output[1678] = '{32'h42c4b6d6};
test_index[1678] = '{2};
test_input[13432:13439] = '{32'hc179233c, 32'hc254ebfb, 32'hc2177a24, 32'h42b3b058, 32'hc10c55eb, 32'h4133b935, 32'hc1d24719, 32'hc2104395};
test_output[1679] = '{32'h42b3b058};
test_index[1679] = '{3};
test_input[13440:13447] = '{32'h42ba6a18, 32'h429fc48b, 32'h4254a59e, 32'h42b2a53c, 32'h426d9be9, 32'h42a8ee4d, 32'h428e630e, 32'hc2520b95};
test_output[1680] = '{32'h42ba6a18};
test_index[1680] = '{0};
test_input[13448:13455] = '{32'hc2b10a48, 32'hc28d360c, 32'h42739911, 32'hc274f3fb, 32'h41b79a67, 32'hc240b9f5, 32'hc2690046, 32'h42bf7ba7};
test_output[1681] = '{32'h42bf7ba7};
test_index[1681] = '{7};
test_input[13456:13463] = '{32'h41e83ca8, 32'h427dcf33, 32'hc2b14412, 32'hc1683098, 32'hc2a99156, 32'hc23e7f0b, 32'h42c6a0f6, 32'hc289c7ea};
test_output[1682] = '{32'h42c6a0f6};
test_index[1682] = '{6};
test_input[13464:13471] = '{32'h420a630a, 32'hc2ad6c12, 32'h42885117, 32'h4210817a, 32'h4242a61a, 32'h42c1d013, 32'h42afa404, 32'h42a38eca};
test_output[1683] = '{32'h42c1d013};
test_index[1683] = '{5};
test_input[13472:13479] = '{32'hc1064816, 32'h42a103c0, 32'h42ac6208, 32'h423910b9, 32'h426e597c, 32'h41c3c5f9, 32'hc1e338b7, 32'hc25d8672};
test_output[1684] = '{32'h42ac6208};
test_index[1684] = '{2};
test_input[13480:13487] = '{32'hc284aa9f, 32'hc2bb344c, 32'h4208cc6f, 32'hc26f72f2, 32'hc259b504, 32'hc2c3d40e, 32'hc1402e94, 32'h42a63588};
test_output[1685] = '{32'h42a63588};
test_index[1685] = '{7};
test_input[13488:13495] = '{32'hc1e46295, 32'h42273e93, 32'h41ca0de4, 32'hc2a6d7a3, 32'h42ac9ae8, 32'hc22dec68, 32'hc2055442, 32'hc134b57a};
test_output[1686] = '{32'h42ac9ae8};
test_index[1686] = '{4};
test_input[13496:13503] = '{32'h42b680a0, 32'hc29a0e81, 32'h429bf7d8, 32'h41e6fa56, 32'hc1062408, 32'hc0b03066, 32'hc29ac2f5, 32'h42bbe7f0};
test_output[1687] = '{32'h42bbe7f0};
test_index[1687] = '{7};
test_input[13504:13511] = '{32'h42681e10, 32'h4158a63f, 32'h42b5f1bd, 32'h42ba1c7a, 32'hc280c2a1, 32'hc28a896e, 32'h424f010d, 32'h41432424};
test_output[1688] = '{32'h42ba1c7a};
test_index[1688] = '{3};
test_input[13512:13519] = '{32'hc21109e8, 32'hc2ba94bd, 32'hc2ab2f08, 32'hc2420733, 32'h42b64e90, 32'h41e36ec4, 32'h41db4e32, 32'h42a488b8};
test_output[1689] = '{32'h42b64e90};
test_index[1689] = '{4};
test_input[13520:13527] = '{32'hc2bb2ff3, 32'hc2656c15, 32'hc17b89c8, 32'h42927e25, 32'hc2a7290c, 32'hc2af432f, 32'hc23b1974, 32'h42a9031b};
test_output[1690] = '{32'h42a9031b};
test_index[1690] = '{7};
test_input[13528:13535] = '{32'hc2b4b7bc, 32'hc282bf75, 32'hc28d7bc7, 32'hc27c3d9f, 32'hc09da201, 32'h41092eba, 32'h42aabbe5, 32'h4298744c};
test_output[1691] = '{32'h42aabbe5};
test_index[1691] = '{6};
test_input[13536:13543] = '{32'hc141dbe4, 32'hc244125b, 32'h42a8b07b, 32'hc1c26e02, 32'hc2afc28c, 32'hc25c4f2f, 32'hc27d484d, 32'h420d2700};
test_output[1692] = '{32'h42a8b07b};
test_index[1692] = '{2};
test_input[13544:13551] = '{32'h40a64f34, 32'hc04c9307, 32'hc114ca3a, 32'hc0b8bed2, 32'h41dd6a2e, 32'hc107bd2d, 32'hc2aab604, 32'h4294644d};
test_output[1693] = '{32'h4294644d};
test_index[1693] = '{7};
test_input[13552:13559] = '{32'hc27f8ea7, 32'h418d7b09, 32'h4181dc68, 32'h42388b5d, 32'hc25cbc48, 32'h401d3139, 32'h42a9f41e, 32'h422b6b3e};
test_output[1694] = '{32'h42a9f41e};
test_index[1694] = '{6};
test_input[13560:13567] = '{32'h41654584, 32'h427b82cb, 32'h4278eda5, 32'hc1cb086c, 32'h41d20f47, 32'hc27027f8, 32'hc265d1aa, 32'hc240ab76};
test_output[1695] = '{32'h427b82cb};
test_index[1695] = '{1};
test_input[13568:13575] = '{32'h424e1a32, 32'h42a06657, 32'hc13ac1f7, 32'h41d880a9, 32'h424c96ec, 32'h426a0391, 32'h4100047f, 32'h4230f5bc};
test_output[1696] = '{32'h42a06657};
test_index[1696] = '{1};
test_input[13576:13583] = '{32'h422fa72d, 32'h40f703c4, 32'h429cfe99, 32'hc1e3af45, 32'hc061e20e, 32'hc282accf, 32'hc2740994, 32'h428fc0c0};
test_output[1697] = '{32'h429cfe99};
test_index[1697] = '{2};
test_input[13584:13591] = '{32'hc2832792, 32'hc29ceb9c, 32'hc18ae673, 32'hc1c513bc, 32'hc2b84897, 32'h416f52c7, 32'hc2b8165b, 32'hc2a3a54b};
test_output[1698] = '{32'h416f52c7};
test_index[1698] = '{5};
test_input[13592:13599] = '{32'h423635d1, 32'h42544246, 32'hc2b7f006, 32'hc2b52a4e, 32'hc28667ba, 32'hc2a6216c, 32'h4281973e, 32'hc29d021b};
test_output[1699] = '{32'h4281973e};
test_index[1699] = '{6};
test_input[13600:13607] = '{32'h40bee89d, 32'h415dd0d8, 32'h400ea9e6, 32'hc1a12e6d, 32'hc2ba80b4, 32'h42b6bcb0, 32'h41d4689b, 32'h421a2428};
test_output[1700] = '{32'h42b6bcb0};
test_index[1700] = '{5};
test_input[13608:13615] = '{32'hc1e81bae, 32'hc2af9682, 32'hc27c69af, 32'hc22427d8, 32'hc2b2e1b0, 32'hc19cf3f1, 32'h420177e3, 32'h4229f583};
test_output[1701] = '{32'h4229f583};
test_index[1701] = '{7};
test_input[13616:13623] = '{32'h41a678f2, 32'h42bda7ca, 32'h42c65e07, 32'hc1522a82, 32'h4264082b, 32'h41aaffe1, 32'hc2b25b30, 32'hc23849ef};
test_output[1702] = '{32'h42c65e07};
test_index[1702] = '{2};
test_input[13624:13631] = '{32'hc2b4e541, 32'h42ba6ac9, 32'h420dc595, 32'hc23abb0b, 32'h426f66cb, 32'hc1c01e74, 32'hc28afda6, 32'h42acbd5e};
test_output[1703] = '{32'h42ba6ac9};
test_index[1703] = '{1};
test_input[13632:13639] = '{32'hc246df18, 32'h427e46f9, 32'h42915aa5, 32'hc24be488, 32'hc2023fdc, 32'hc26d8d0b, 32'h4104b10c, 32'h419f6104};
test_output[1704] = '{32'h42915aa5};
test_index[1704] = '{2};
test_input[13640:13647] = '{32'h4093ab16, 32'hc2b6712f, 32'hc1de52d9, 32'h428398ee, 32'h40af532d, 32'hc205ec49, 32'hc10b5d60, 32'hc294682a};
test_output[1705] = '{32'h428398ee};
test_index[1705] = '{3};
test_input[13648:13655] = '{32'h3f8da6a9, 32'hc23f3e29, 32'h423fe6e1, 32'h4235c036, 32'hc064395e, 32'hc1d3155b, 32'hc0a0b394, 32'hc20abd82};
test_output[1706] = '{32'h423fe6e1};
test_index[1706] = '{2};
test_input[13656:13663] = '{32'h4253d0da, 32'hc254d5a4, 32'hc26f2f0d, 32'h413d57d1, 32'hc200a672, 32'hc20517ae, 32'h41afd771, 32'h41b9cf9d};
test_output[1707] = '{32'h4253d0da};
test_index[1707] = '{0};
test_input[13664:13671] = '{32'h42bd7922, 32'h40ca930d, 32'h4282ab91, 32'h429c46f6, 32'h41f6c8a6, 32'h428071b0, 32'h40a4f303, 32'h4211b273};
test_output[1708] = '{32'h42bd7922};
test_index[1708] = '{0};
test_input[13672:13679] = '{32'h425be47d, 32'hc1999a69, 32'h3f3f16f4, 32'h425065ca, 32'hc2b83d69, 32'h41db0d30, 32'hc0340abc, 32'hc2c4139a};
test_output[1709] = '{32'h425be47d};
test_index[1709] = '{0};
test_input[13680:13687] = '{32'h3fd48719, 32'hc1ecdd80, 32'h429c7450, 32'h405473f9, 32'h416f89d3, 32'h42c13181, 32'h41dfe736, 32'h4011ab25};
test_output[1710] = '{32'h42c13181};
test_index[1710] = '{5};
test_input[13688:13695] = '{32'hc23f011a, 32'h418d0058, 32'h42ae3ee3, 32'hc2b045fe, 32'h426a5be0, 32'h4225eab1, 32'h424638e9, 32'hc2862079};
test_output[1711] = '{32'h42ae3ee3};
test_index[1711] = '{2};
test_input[13696:13703] = '{32'hc0c97e8e, 32'hc183a9a8, 32'hc2aa19b9, 32'hbf186189, 32'hc21982f6, 32'hc2bd80b0, 32'hc2a9c1d9, 32'h42c6f05d};
test_output[1712] = '{32'h42c6f05d};
test_index[1712] = '{7};
test_input[13704:13711] = '{32'h41e533d7, 32'h428c112c, 32'hbf53faed, 32'hc1fb2c30, 32'h429d08ef, 32'hc24102f7, 32'h41fd91ed, 32'hc1f3bfbd};
test_output[1713] = '{32'h429d08ef};
test_index[1713] = '{4};
test_input[13712:13719] = '{32'hc1ad27ce, 32'hc27a485a, 32'hc29c71d3, 32'hc2797f7f, 32'hc1928d22, 32'hc0bcab67, 32'hc29ba623, 32'hc2bc40ab};
test_output[1714] = '{32'hc0bcab67};
test_index[1714] = '{5};
test_input[13720:13727] = '{32'h42af32bd, 32'h428c58cc, 32'h422d2bd3, 32'h42c2e05a, 32'h4175b362, 32'hc2b0b08b, 32'hc1eac884, 32'h4284384b};
test_output[1715] = '{32'h42c2e05a};
test_index[1715] = '{3};
test_input[13728:13735] = '{32'h42042ef3, 32'h4285506a, 32'h4206c96b, 32'h424e331b, 32'h42bcf898, 32'h425c2a7f, 32'h4235609b, 32'hc2aa0d0a};
test_output[1716] = '{32'h42bcf898};
test_index[1716] = '{4};
test_input[13736:13743] = '{32'hc28827f1, 32'hc275376f, 32'h42c70ea2, 32'hc2abeacc, 32'h42ab77a6, 32'h42683bc4, 32'hc0b2ab35, 32'hc297edbe};
test_output[1717] = '{32'h42c70ea2};
test_index[1717] = '{2};
test_input[13744:13751] = '{32'h41fe50d4, 32'h42a3a23c, 32'hc2a1d6c5, 32'hc2747fe7, 32'h42370b8a, 32'hc20469ba, 32'hc1ae4627, 32'h429d9dfa};
test_output[1718] = '{32'h42a3a23c};
test_index[1718] = '{1};
test_input[13752:13759] = '{32'h4289132e, 32'hc226ec8a, 32'h41fc759d, 32'hc14c3205, 32'h426cbaaf, 32'h419909cc, 32'h428e2b89, 32'h4143ff71};
test_output[1719] = '{32'h428e2b89};
test_index[1719] = '{6};
test_input[13760:13767] = '{32'hc241780a, 32'h421a7c16, 32'hc1b3b5d7, 32'hc0289acf, 32'hc2b31759, 32'h42677b8a, 32'h42936634, 32'h42ab3c2c};
test_output[1720] = '{32'h42ab3c2c};
test_index[1720] = '{7};
test_input[13768:13775] = '{32'h42a5e593, 32'h4268126c, 32'hc150213c, 32'hc25caa99, 32'hc23b85da, 32'hc1efbfbd, 32'hc1033185, 32'h42108da6};
test_output[1721] = '{32'h42a5e593};
test_index[1721] = '{0};
test_input[13776:13783] = '{32'h428e8266, 32'hc06dfe37, 32'hc234661f, 32'hc1a01816, 32'h42590e11, 32'h41b22a24, 32'hc1c4e938, 32'h424718d3};
test_output[1722] = '{32'h428e8266};
test_index[1722] = '{0};
test_input[13784:13791] = '{32'h4276235e, 32'h42121847, 32'hc256f07d, 32'hc1aecdbf, 32'h428c0cfb, 32'hc28afe66, 32'hc0fc756e, 32'hc2c4e24a};
test_output[1723] = '{32'h428c0cfb};
test_index[1723] = '{4};
test_input[13792:13799] = '{32'h4273eefe, 32'hc15885d1, 32'h4123b086, 32'hc203fe72, 32'h428b19ce, 32'h427d84d7, 32'h424febc0, 32'h41a3a1a7};
test_output[1724] = '{32'h428b19ce};
test_index[1724] = '{4};
test_input[13800:13807] = '{32'hc2b90c39, 32'hc240b3b4, 32'h42b5d0e6, 32'hc297e1de, 32'h425e01fd, 32'h42a9af0d, 32'hc1d52a31, 32'hc28bb8cf};
test_output[1725] = '{32'h42b5d0e6};
test_index[1725] = '{2};
test_input[13808:13815] = '{32'h42a423c6, 32'hc24995e0, 32'hc2b90a00, 32'h429b2daf, 32'h42a3633a, 32'hc1b26d83, 32'h4293f11b, 32'hc1a4b101};
test_output[1726] = '{32'h42a423c6};
test_index[1726] = '{0};
test_input[13816:13823] = '{32'hc2300aae, 32'h42204120, 32'hc1dbd299, 32'h421d7d4c, 32'h3ed2e516, 32'h42384a4c, 32'h42216925, 32'h420ec722};
test_output[1727] = '{32'h42384a4c};
test_index[1727] = '{5};
test_input[13824:13831] = '{32'h429f65c2, 32'hc29ae7f6, 32'hc23328bb, 32'hc2bd6f50, 32'h42a5bf15, 32'h42a7b5c5, 32'h426f5274, 32'h40dab3fb};
test_output[1728] = '{32'h42a7b5c5};
test_index[1728] = '{5};
test_input[13832:13839] = '{32'h42514a94, 32'hc0f5b068, 32'h4286cbcd, 32'h3f94c8ae, 32'h41c1d607, 32'hc2108c59, 32'h420aa3fd, 32'h41c77f7b};
test_output[1729] = '{32'h4286cbcd};
test_index[1729] = '{2};
test_input[13840:13847] = '{32'h41e437d4, 32'h4288bcf1, 32'h42848a7d, 32'hc2b3d006, 32'h42c77252, 32'h428e2afd, 32'hc20c263a, 32'h42934aa3};
test_output[1730] = '{32'h42c77252};
test_index[1730] = '{4};
test_input[13848:13855] = '{32'h41b13fa2, 32'hc2762c9b, 32'hc274f563, 32'h42ac8208, 32'hc0005269, 32'h429e6e15, 32'h4248f761, 32'hc111c2aa};
test_output[1731] = '{32'h42ac8208};
test_index[1731] = '{3};
test_input[13856:13863] = '{32'h4241ed47, 32'hc1b36439, 32'h427ad3d6, 32'h40fc8bd9, 32'hc23c9b00, 32'h41e834b9, 32'h421d55fc, 32'h428a9435};
test_output[1732] = '{32'h428a9435};
test_index[1732] = '{7};
test_input[13864:13871] = '{32'h4210e440, 32'h42393163, 32'hc2c6b0ba, 32'h428fcdfc, 32'h42add7eb, 32'h424d1fc7, 32'h42634e6c, 32'hc2123724};
test_output[1733] = '{32'h42add7eb};
test_index[1733] = '{4};
test_input[13872:13879] = '{32'hc26019c7, 32'h417fc994, 32'hc286949b, 32'hc1686095, 32'h4260a85f, 32'hc2bacdbb, 32'hc2c569fd, 32'h41eadb4c};
test_output[1734] = '{32'h4260a85f};
test_index[1734] = '{4};
test_input[13880:13887] = '{32'h4205a38e, 32'hc1b7bfd7, 32'h42abfa94, 32'h42a186c6, 32'h41e8d771, 32'h429018e1, 32'h420d08c4, 32'h42b02c8d};
test_output[1735] = '{32'h42b02c8d};
test_index[1735] = '{7};
test_input[13888:13895] = '{32'h4272907d, 32'h422b82f2, 32'h415b6488, 32'h4295e662, 32'hc1babedd, 32'hc2a03023, 32'hc224eadc, 32'h42abfdcf};
test_output[1736] = '{32'h42abfdcf};
test_index[1736] = '{7};
test_input[13896:13903] = '{32'h42c77b5c, 32'hc13e8072, 32'h420a03ab, 32'h428e7b41, 32'h42ba793a, 32'hc266adc8, 32'h42973db6, 32'h42b7a0f8};
test_output[1737] = '{32'h42c77b5c};
test_index[1737] = '{0};
test_input[13904:13911] = '{32'hc2769157, 32'h41ad38cf, 32'h420196ca, 32'hc23ea36c, 32'hc23153a3, 32'hc261a540, 32'h4296c216, 32'h40464973};
test_output[1738] = '{32'h4296c216};
test_index[1738] = '{6};
test_input[13912:13919] = '{32'h42a330a0, 32'hc0d627bc, 32'hc28adc29, 32'hc11ef616, 32'h413b1a3c, 32'h41ba962d, 32'h41a9faf8, 32'h40d77458};
test_output[1739] = '{32'h42a330a0};
test_index[1739] = '{0};
test_input[13920:13927] = '{32'h425cc884, 32'h42a66863, 32'h3f482891, 32'hc1f3df51, 32'hc2bd24bd, 32'h41dd8a0f, 32'h42948308, 32'hc1d09907};
test_output[1740] = '{32'h42a66863};
test_index[1740] = '{1};
test_input[13928:13935] = '{32'h413b3efd, 32'hc2beac66, 32'h41ae1819, 32'hc15bd068, 32'h426aecb6, 32'hc1162eee, 32'h42a5ed20, 32'h42770496};
test_output[1741] = '{32'h42a5ed20};
test_index[1741] = '{6};
test_input[13936:13943] = '{32'hc1edbca7, 32'hc27e0bb4, 32'h421dc757, 32'hc299ce88, 32'h41765f19, 32'h4202dd7d, 32'h428c278d, 32'h40b1c051};
test_output[1742] = '{32'h428c278d};
test_index[1742] = '{6};
test_input[13944:13951] = '{32'hc1fe457d, 32'hc15ff7d2, 32'hc2800770, 32'hc1da2146, 32'h4298fd9d, 32'hc292562f, 32'h4240db8c, 32'hc2b7317e};
test_output[1743] = '{32'h4298fd9d};
test_index[1743] = '{4};
test_input[13952:13959] = '{32'h3f3cd7bd, 32'hc1459a00, 32'h42a4f681, 32'hc28d9c0d, 32'h42c29171, 32'h42806c1d, 32'h42940688, 32'hc0904729};
test_output[1744] = '{32'h42c29171};
test_index[1744] = '{4};
test_input[13960:13967] = '{32'hc17e8d73, 32'hc1d0b82b, 32'h41d53bc5, 32'hc29d3244, 32'hc24a2465, 32'hc2122758, 32'h412c5d58, 32'hc21e29a5};
test_output[1745] = '{32'h41d53bc5};
test_index[1745] = '{2};
test_input[13968:13975] = '{32'hc26b31f0, 32'hc242d7ba, 32'hc20cc932, 32'h42aa737b, 32'hc2bfaa5a, 32'h42857196, 32'h4258b026, 32'hc22613ec};
test_output[1746] = '{32'h42aa737b};
test_index[1746] = '{3};
test_input[13976:13983] = '{32'h3f21629b, 32'h41d2a793, 32'hc1c87d33, 32'hc148cef2, 32'hc22d1f4a, 32'h42acf64f, 32'h4283fe62, 32'h42259fd5};
test_output[1747] = '{32'h42acf64f};
test_index[1747] = '{5};
test_input[13984:13991] = '{32'h42272f89, 32'h405bac38, 32'h42b09c8b, 32'hc23d91a9, 32'h42a57eca, 32'h42b7741c, 32'hc0f503e3, 32'hc234fe3d};
test_output[1748] = '{32'h42b7741c};
test_index[1748] = '{5};
test_input[13992:13999] = '{32'hc2c36894, 32'hc189b87d, 32'hc278c849, 32'hc23388f5, 32'h4290fc86, 32'h42ada860, 32'hc2abfd02, 32'h42238314};
test_output[1749] = '{32'h42ada860};
test_index[1749] = '{5};
test_input[14000:14007] = '{32'hc2afeaff, 32'h42906a02, 32'h4222e279, 32'h4204960b, 32'hc230416f, 32'hc24e4bd9, 32'h4188ce88, 32'hc29a426b};
test_output[1750] = '{32'h42906a02};
test_index[1750] = '{1};
test_input[14008:14015] = '{32'hc2bc43bf, 32'h42ab6174, 32'hc2c0b7db, 32'hc2218729, 32'hc1809411, 32'hc2b82ec2, 32'h41cf4579, 32'hc24d9d8e};
test_output[1751] = '{32'h42ab6174};
test_index[1751] = '{1};
test_input[14016:14023] = '{32'h42694847, 32'h428c585c, 32'hc27bc6ec, 32'h41c8880b, 32'hc27dcdf5, 32'h42830019, 32'h41808e96, 32'hc25e72b3};
test_output[1752] = '{32'h428c585c};
test_index[1752] = '{1};
test_input[14024:14031] = '{32'h414496f5, 32'h424569d6, 32'h40a9a0d6, 32'h42b7f589, 32'h428d5379, 32'hc1500b40, 32'hc1f4dbd2, 32'hc27085dd};
test_output[1753] = '{32'h42b7f589};
test_index[1753] = '{3};
test_input[14032:14039] = '{32'h42925c3e, 32'h4080423e, 32'h42167c47, 32'h42682a3b, 32'hc259a48e, 32'h427ffc04, 32'h41879dc9, 32'hc181603e};
test_output[1754] = '{32'h42925c3e};
test_index[1754] = '{0};
test_input[14040:14047] = '{32'hc281ed86, 32'hc1cdf644, 32'hc26cc48b, 32'h427fde90, 32'h4215c49f, 32'h42b4c79d, 32'h42b27688, 32'h42b01b92};
test_output[1755] = '{32'h42b4c79d};
test_index[1755] = '{5};
test_input[14048:14055] = '{32'hc28c16d4, 32'hc1cd48c7, 32'hc28cbc90, 32'hc2158a62, 32'hc15854e0, 32'hc1aae562, 32'h41cfde51, 32'hc22feabc};
test_output[1756] = '{32'h41cfde51};
test_index[1756] = '{6};
test_input[14056:14063] = '{32'h41913a39, 32'hc186bbec, 32'hc204131d, 32'h421fe7fe, 32'h42c1d99a, 32'h420e08b1, 32'hc2a38af9, 32'hc2b92ad1};
test_output[1757] = '{32'h42c1d99a};
test_index[1757] = '{4};
test_input[14064:14071] = '{32'h415aee20, 32'hc213ea5a, 32'hc1901561, 32'hc29ddc6f, 32'hc2ade094, 32'hc170249c, 32'hc0f00da8, 32'h42a287be};
test_output[1758] = '{32'h42a287be};
test_index[1758] = '{7};
test_input[14072:14079] = '{32'h4286aee0, 32'hc2445e16, 32'hc29ce2d9, 32'hc1a23ed2, 32'h4256645b, 32'h421abf5a, 32'h41c647d1, 32'h4167659a};
test_output[1759] = '{32'h4286aee0};
test_index[1759] = '{0};
test_input[14080:14087] = '{32'h4288c859, 32'h41fa6c52, 32'h414efc6a, 32'hc19d5b9b, 32'h42b2f67e, 32'h418d1712, 32'hc2a424aa, 32'hc2878678};
test_output[1760] = '{32'h42b2f67e};
test_index[1760] = '{4};
test_input[14088:14095] = '{32'h420bc730, 32'h426e488e, 32'hc26e0d1a, 32'h41dfd4fc, 32'hc0f32a8c, 32'h428d6376, 32'hc21c5cd9, 32'h419cbfaa};
test_output[1761] = '{32'h428d6376};
test_index[1761] = '{5};
test_input[14096:14103] = '{32'hc12441e4, 32'hc2a57a5b, 32'hc2b74987, 32'hc252142f, 32'hc284b816, 32'h4281308b, 32'h4206b51c, 32'h4271e122};
test_output[1762] = '{32'h4281308b};
test_index[1762] = '{5};
test_input[14104:14111] = '{32'h424dec58, 32'hc1067252, 32'h40d11270, 32'hc21fec8d, 32'h42429ba2, 32'h428717ba, 32'hc28f8f59, 32'h422f52cc};
test_output[1763] = '{32'h428717ba};
test_index[1763] = '{5};
test_input[14112:14119] = '{32'h41e6dfe1, 32'h427a09a4, 32'h422f59d0, 32'hc24f50da, 32'h424eb5bb, 32'hc1c3f606, 32'h41abcf08, 32'h42bdcf7e};
test_output[1764] = '{32'h42bdcf7e};
test_index[1764] = '{7};
test_input[14120:14127] = '{32'h42a42f95, 32'h42820d98, 32'h41da7c7c, 32'h42287d6e, 32'hc1621416, 32'hc2af27f0, 32'h42a37a7f, 32'h42b6ff0e};
test_output[1765] = '{32'h42b6ff0e};
test_index[1765] = '{7};
test_input[14128:14135] = '{32'h428f1a09, 32'hc1e26a64, 32'hc2c54f4c, 32'hc2453a71, 32'h41cfaa37, 32'h4139af96, 32'hc2a3f2de, 32'hc2c62c2a};
test_output[1766] = '{32'h428f1a09};
test_index[1766] = '{0};
test_input[14136:14143] = '{32'hc231974d, 32'hc27896ac, 32'h42c10337, 32'hbe2f5047, 32'h41bc59b9, 32'hc275747b, 32'hc2bab2b5, 32'h3f89e468};
test_output[1767] = '{32'h42c10337};
test_index[1767] = '{2};
test_input[14144:14151] = '{32'h41fe459f, 32'h428ddd04, 32'hc232e458, 32'h419bef0e, 32'hc0405f97, 32'hc29b8f9a, 32'h426a0e8e, 32'h42bdea88};
test_output[1768] = '{32'h42bdea88};
test_index[1768] = '{7};
test_input[14152:14159] = '{32'h41fc57de, 32'hc10c546d, 32'h42ac230c, 32'hc1bea8ef, 32'hc2808068, 32'h4129396d, 32'h3f384672, 32'h41a60864};
test_output[1769] = '{32'h42ac230c};
test_index[1769] = '{2};
test_input[14160:14167] = '{32'hc2449ef4, 32'hc2bad619, 32'hc28b9407, 32'h42a1f3b8, 32'hc29bfe40, 32'h3fb2de0a, 32'h420be43f, 32'h42c61d66};
test_output[1770] = '{32'h42c61d66};
test_index[1770] = '{7};
test_input[14168:14175] = '{32'h40d11585, 32'hc00d1dd8, 32'hc24d7e04, 32'h41a63224, 32'hc222c43f, 32'h41f7834e, 32'h40cdb61e, 32'hc1a42167};
test_output[1771] = '{32'h41f7834e};
test_index[1771] = '{5};
test_input[14176:14183] = '{32'hc2b50da0, 32'hc2401c74, 32'h42bc7820, 32'h41eddeb5, 32'hc2bc2b3b, 32'h404c5ba7, 32'h42860d94, 32'hc269b482};
test_output[1772] = '{32'h42bc7820};
test_index[1772] = '{2};
test_input[14184:14191] = '{32'h4251924e, 32'h42a46c1d, 32'h42b8c60b, 32'h424d3792, 32'h42ab8f7d, 32'hc0434627, 32'hc283ca07, 32'h42aef340};
test_output[1773] = '{32'h42b8c60b};
test_index[1773] = '{2};
test_input[14192:14199] = '{32'h427225ea, 32'h426e9812, 32'h422be429, 32'hc2b0b72e, 32'h429425ed, 32'h423313d4, 32'hc28cb031, 32'hc29bee5a};
test_output[1774] = '{32'h429425ed};
test_index[1774] = '{4};
test_input[14200:14207] = '{32'hc2b09370, 32'hc24f9cf2, 32'hc2a460eb, 32'h427cfec7, 32'hc26d188b, 32'h40c2271a, 32'hc29b9e49, 32'h402044e6};
test_output[1775] = '{32'h427cfec7};
test_index[1775] = '{3};
test_input[14208:14215] = '{32'h419e649e, 32'hbf52d9e2, 32'hc093ef08, 32'hc270a6a9, 32'hc2859d4d, 32'h42c5f4a7, 32'hc2367d94, 32'hc0c4e81f};
test_output[1776] = '{32'h42c5f4a7};
test_index[1776] = '{5};
test_input[14216:14223] = '{32'hbf1bb3b7, 32'hc071aa47, 32'h40eaa731, 32'h411a739e, 32'hc23e9b63, 32'hc240e92b, 32'h42b63cf3, 32'hc2a018b3};
test_output[1777] = '{32'h42b63cf3};
test_index[1777] = '{6};
test_input[14224:14231] = '{32'hc28019a6, 32'h429055cb, 32'h428bd729, 32'hbf5f60f6, 32'hc0bf4dbc, 32'hc244aeef, 32'h4229a8c5, 32'hc2053c82};
test_output[1778] = '{32'h429055cb};
test_index[1778] = '{1};
test_input[14232:14239] = '{32'hbe48c5ed, 32'h4113a1fc, 32'h41bf8b1a, 32'h42955e72, 32'h42ba5465, 32'h40e8644b, 32'h429e672f, 32'h41d47c28};
test_output[1779] = '{32'h42ba5465};
test_index[1779] = '{4};
test_input[14240:14247] = '{32'h42164b9e, 32'hc20c5dd0, 32'h42990e62, 32'hc28e6ff6, 32'h42973fd8, 32'h42b02a1a, 32'hc1d81ea4, 32'h4252e1c5};
test_output[1780] = '{32'h42b02a1a};
test_index[1780] = '{5};
test_input[14248:14255] = '{32'hc1c0ba98, 32'h42b07000, 32'h4261a653, 32'h42124cb3, 32'h420f3ba7, 32'h419d08a2, 32'hc08e2d67, 32'h415e7d3a};
test_output[1781] = '{32'h42b07000};
test_index[1781] = '{1};
test_input[14256:14263] = '{32'hc28356fb, 32'h4220964a, 32'h41f1f5a0, 32'h425642df, 32'hc1ed1cd6, 32'h429abb47, 32'h41c12352, 32'hc27932b6};
test_output[1782] = '{32'h429abb47};
test_index[1782] = '{5};
test_input[14264:14271] = '{32'h4293d31f, 32'hc1905d99, 32'h42912851, 32'hc209d829, 32'hc214889f, 32'h429c1adf, 32'hc2564843, 32'h42ab9310};
test_output[1783] = '{32'h42ab9310};
test_index[1783] = '{7};
test_input[14272:14279] = '{32'hc23d1e7d, 32'hc2a2a101, 32'h41c31465, 32'h42bdf869, 32'hc13f0c59, 32'h4296ea1e, 32'h424140cd, 32'h428a9bbb};
test_output[1784] = '{32'h42bdf869};
test_index[1784] = '{3};
test_input[14280:14287] = '{32'hc2b85a4b, 32'hc22397e8, 32'h405432da, 32'hc2ae48ff, 32'h429d4010, 32'hc23e030d, 32'h40f96fa8, 32'hc1d5d3ff};
test_output[1785] = '{32'h429d4010};
test_index[1785] = '{4};
test_input[14288:14295] = '{32'hc1c0dbb2, 32'hc195a46d, 32'hc2376568, 32'h421e0ef0, 32'h42b8dc21, 32'h4186bef6, 32'h41f90e29, 32'hc2ae76c1};
test_output[1786] = '{32'h42b8dc21};
test_index[1786] = '{4};
test_input[14296:14303] = '{32'hc2594770, 32'hc2a15fc5, 32'h41b31261, 32'h420e419f, 32'hc23e3d3c, 32'hc0eabd30, 32'hc1f7c508, 32'hc2b8bbc8};
test_output[1787] = '{32'h420e419f};
test_index[1787] = '{3};
test_input[14304:14311] = '{32'h42615430, 32'h429e5aca, 32'hc205028a, 32'hc2bc6514, 32'hc225814a, 32'h41b7c299, 32'h4285c95f, 32'hc2a3ab34};
test_output[1788] = '{32'h429e5aca};
test_index[1788] = '{1};
test_input[14312:14319] = '{32'h42c74aec, 32'hc1e6bc73, 32'h410a1e94, 32'hc232535f, 32'hc2777de9, 32'hc2a24eaf, 32'h427725b9, 32'h42a86c9e};
test_output[1789] = '{32'h42c74aec};
test_index[1789] = '{0};
test_input[14320:14327] = '{32'h41340ef4, 32'hc28b3abb, 32'h42750aa8, 32'h41623225, 32'h4225988a, 32'h429051f8, 32'hc2bc753e, 32'h4230ea9b};
test_output[1790] = '{32'h429051f8};
test_index[1790] = '{5};
test_input[14328:14335] = '{32'hc2044dd6, 32'h3fdba274, 32'h42833173, 32'hc289ee52, 32'hc22bb679, 32'h427d7e4a, 32'hc18b192f, 32'hc28e7e7c};
test_output[1791] = '{32'h42833173};
test_index[1791] = '{2};
test_input[14336:14343] = '{32'hc1bf5b29, 32'hc2974587, 32'h4292b3aa, 32'hc211aa33, 32'h42947906, 32'h4139d9a1, 32'hc2743b64, 32'hc184b4e6};
test_output[1792] = '{32'h42947906};
test_index[1792] = '{4};
test_input[14344:14351] = '{32'h4123a8f9, 32'hc266960e, 32'h428e0c4e, 32'hc184dfe4, 32'hc16b8f17, 32'hc1f53ca3, 32'hc2824e50, 32'h41867c6c};
test_output[1793] = '{32'h428e0c4e};
test_index[1793] = '{2};
test_input[14352:14359] = '{32'h42836be7, 32'hc2a199e3, 32'h422124eb, 32'h42ae1101, 32'h40fa1a60, 32'h4178b082, 32'h4106135e, 32'hc2070ef3};
test_output[1794] = '{32'h42ae1101};
test_index[1794] = '{3};
test_input[14360:14367] = '{32'h423fed62, 32'h42b35bdc, 32'h421b20ac, 32'h4287a972, 32'hc28b1474, 32'h4118612d, 32'h41a9101c, 32'hc27a95b3};
test_output[1795] = '{32'h42b35bdc};
test_index[1795] = '{1};
test_input[14368:14375] = '{32'hc212b7a2, 32'h42b1831f, 32'h427f68ff, 32'h427279ee, 32'h428da63b, 32'h42900afd, 32'hc2c0a63a, 32'h42751b90};
test_output[1796] = '{32'h42b1831f};
test_index[1796] = '{1};
test_input[14376:14383] = '{32'h4298ce90, 32'hc2077e1b, 32'h42792303, 32'hc23e8d56, 32'hc2b6b3bd, 32'hc212940f, 32'hbf886a72, 32'h423c79f2};
test_output[1797] = '{32'h4298ce90};
test_index[1797] = '{0};
test_input[14384:14391] = '{32'h42904e1b, 32'hc28f39d2, 32'hc212e5a1, 32'h421789e9, 32'h4079f6ab, 32'hc26c896c, 32'h428ce117, 32'h41fdd2cd};
test_output[1798] = '{32'h42904e1b};
test_index[1798] = '{0};
test_input[14392:14399] = '{32'h42037cd5, 32'hc26a56e0, 32'hc1d4a089, 32'hc0aca86b, 32'h4287178b, 32'hc102671f, 32'hc2c457d0, 32'hc1da7cb7};
test_output[1799] = '{32'h4287178b};
test_index[1799] = '{4};
test_input[14400:14407] = '{32'hc283daea, 32'h42afc883, 32'h41cb617b, 32'hc040afb6, 32'hc1e5ddf4, 32'h4295e49e, 32'h42c2cb82, 32'hc2183e1a};
test_output[1800] = '{32'h42c2cb82};
test_index[1800] = '{6};
test_input[14408:14415] = '{32'h428b9a12, 32'hc26ffeb9, 32'hc0b54191, 32'h4100cdfd, 32'hc289b2ff, 32'h41bbae38, 32'h3f4e8a59, 32'hc1bca1f2};
test_output[1801] = '{32'h428b9a12};
test_index[1801] = '{0};
test_input[14416:14423] = '{32'h426b441e, 32'hc2ab8339, 32'h428e8406, 32'hc0f871de, 32'hc2ac64ec, 32'hc2c79b73, 32'h4249021d, 32'h42b52499};
test_output[1802] = '{32'h42b52499};
test_index[1802] = '{7};
test_input[14424:14431] = '{32'h412942af, 32'hc14feebd, 32'hc1dfcded, 32'hc21ccd70, 32'h42aeaf2d, 32'h4215de08, 32'h4234b649, 32'h42c39077};
test_output[1803] = '{32'h42c39077};
test_index[1803] = '{7};
test_input[14432:14439] = '{32'h40d811ca, 32'h424f69dc, 32'h42c27c76, 32'hc1db517a, 32'h42c7762e, 32'h42827aa4, 32'hc055e4de, 32'hc2594170};
test_output[1804] = '{32'h42c7762e};
test_index[1804] = '{4};
test_input[14440:14447] = '{32'h411e37d7, 32'hc19d33b0, 32'hc284535a, 32'h4223bb40, 32'hc28b9806, 32'hc16b11fb, 32'h40cb6f53, 32'hc2bd7bbb};
test_output[1805] = '{32'h4223bb40};
test_index[1805] = '{3};
test_input[14448:14455] = '{32'hc24b33cf, 32'h3fcda04a, 32'h428aedfb, 32'hc284d3ac, 32'h41f46b49, 32'hc28599f1, 32'h428242f2, 32'hc1869ca5};
test_output[1806] = '{32'h428aedfb};
test_index[1806] = '{2};
test_input[14456:14463] = '{32'hc26de436, 32'hc2c5d6fa, 32'h42975073, 32'h414cdfce, 32'hc2355bf6, 32'h42bb2263, 32'h429551f7, 32'h42ae7ac4};
test_output[1807] = '{32'h42bb2263};
test_index[1807] = '{5};
test_input[14464:14471] = '{32'h42559d9a, 32'hbfd64f0e, 32'hc2a89d04, 32'hc21fe1b0, 32'h40f4100b, 32'h427bef7e, 32'hc0e4516f, 32'h42980cfc};
test_output[1808] = '{32'h42980cfc};
test_index[1808] = '{7};
test_input[14472:14479] = '{32'h425b49e2, 32'h41de0354, 32'h420fb6d3, 32'hc2a838df, 32'h420e5d98, 32'h4258eb3a, 32'h42559925, 32'hc2688cc4};
test_output[1809] = '{32'h425b49e2};
test_index[1809] = '{0};
test_input[14480:14487] = '{32'h425bee5c, 32'hc284b0d4, 32'h41128fa1, 32'h42adfaa6, 32'h421d05dd, 32'hc29bae6f, 32'hc2aee54d, 32'hc23c30d6};
test_output[1810] = '{32'h42adfaa6};
test_index[1810] = '{3};
test_input[14488:14495] = '{32'hc248bf53, 32'h42c5ec67, 32'hc2aa0cb5, 32'h41e6e7ff, 32'h426cd2cb, 32'h40b1571d, 32'h4154bb57, 32'h406fce97};
test_output[1811] = '{32'h42c5ec67};
test_index[1811] = '{1};
test_input[14496:14503] = '{32'h3c0c34b2, 32'h405724a9, 32'hc1effbce, 32'h42bed8a9, 32'h40b92434, 32'h4296fda1, 32'hc234ea48, 32'hc2024979};
test_output[1812] = '{32'h42bed8a9};
test_index[1812] = '{3};
test_input[14504:14511] = '{32'hc26edf5e, 32'h4290fd5d, 32'hc23bb0a8, 32'hc1694acf, 32'hbe800add, 32'hc26b8b8c, 32'hc2ad00a4, 32'h428e4e9c};
test_output[1813] = '{32'h4290fd5d};
test_index[1813] = '{1};
test_input[14512:14519] = '{32'hc19f13e7, 32'h4239dad7, 32'hc2a45788, 32'hc2848ee4, 32'h4243dc7f, 32'hc1c35ade, 32'h4223097a, 32'hc28c0fb1};
test_output[1814] = '{32'h4243dc7f};
test_index[1814] = '{4};
test_input[14520:14527] = '{32'hc1bc5c9c, 32'hc29a2a74, 32'hc269993b, 32'hc274f575, 32'hc1baf943, 32'h42932e85, 32'h428b633b, 32'h42070ead};
test_output[1815] = '{32'h42932e85};
test_index[1815] = '{5};
test_input[14528:14535] = '{32'hc2c07500, 32'hc247c0dd, 32'hc28be436, 32'h42c4112d, 32'hc2432175, 32'hc2a8916c, 32'h41f80b31, 32'h41c6d53b};
test_output[1816] = '{32'h42c4112d};
test_index[1816] = '{3};
test_input[14536:14543] = '{32'h428b9d35, 32'hc21a7575, 32'hc293b863, 32'h420d0644, 32'h42b63a0b, 32'h420bf1b3, 32'hc2421730, 32'h4203ea33};
test_output[1817] = '{32'h42b63a0b};
test_index[1817] = '{4};
test_input[14544:14551] = '{32'hc27f13a9, 32'h41fce64f, 32'hc2a17681, 32'hc2c42f09, 32'hc2b12437, 32'hc293dfef, 32'h42a1b5b6, 32'hc11fa49e};
test_output[1818] = '{32'h42a1b5b6};
test_index[1818] = '{6};
test_input[14552:14559] = '{32'hc07a9cf8, 32'hc221e6e4, 32'h428a4e9b, 32'hc1a23418, 32'h4249bb4e, 32'hc23a4729, 32'h42b50c49, 32'h42be20ea};
test_output[1819] = '{32'h42be20ea};
test_index[1819] = '{7};
test_input[14560:14567] = '{32'h42765748, 32'h41451800, 32'hc28035cd, 32'hc2096a61, 32'h415525f8, 32'hc2909e48, 32'hc2ac000b, 32'h42b07b07};
test_output[1820] = '{32'h42b07b07};
test_index[1820] = '{7};
test_input[14568:14575] = '{32'h410d2300, 32'h4293d3e2, 32'h429cfab6, 32'h423cd6ad, 32'h429c5608, 32'h4281900b, 32'h42bc6f66, 32'hc256008c};
test_output[1821] = '{32'h42bc6f66};
test_index[1821] = '{6};
test_input[14576:14583] = '{32'h42063e14, 32'hc20d87e9, 32'hc2a8a2fe, 32'h429a5332, 32'hc1fe71c6, 32'hc286aec7, 32'hc287a34e, 32'h40683429};
test_output[1822] = '{32'h429a5332};
test_index[1822] = '{3};
test_input[14584:14591] = '{32'h41cf1614, 32'h4232f4cd, 32'hc2a2a732, 32'hc171396d, 32'h412e7327, 32'hc283abd9, 32'h42a1d49e, 32'h42bf98bc};
test_output[1823] = '{32'h42bf98bc};
test_index[1823] = '{7};
test_input[14592:14599] = '{32'h424d4429, 32'h429b031f, 32'h4290f89f, 32'h42b520b8, 32'hc23e5842, 32'hc0597730, 32'h41ca7957, 32'hc2424d37};
test_output[1824] = '{32'h42b520b8};
test_index[1824] = '{3};
test_input[14600:14607] = '{32'h420e932e, 32'hc24846ac, 32'h41791743, 32'h42a4a0ff, 32'hc2bf14e8, 32'hc216de96, 32'hc152ad6c, 32'hc2a5407c};
test_output[1825] = '{32'h42a4a0ff};
test_index[1825] = '{3};
test_input[14608:14615] = '{32'h42abc6cc, 32'h41256136, 32'h42c7de25, 32'h42c51c90, 32'h42a18a5c, 32'h4251e5b9, 32'hc2b6eb5a, 32'h4230fced};
test_output[1826] = '{32'h42c7de25};
test_index[1826] = '{2};
test_input[14616:14623] = '{32'hc28f03f6, 32'h42721041, 32'hc2a718aa, 32'h42ae8455, 32'h422ae6ca, 32'hc274c4b4, 32'hc2a01d06, 32'h420bf2ba};
test_output[1827] = '{32'h42ae8455};
test_index[1827] = '{3};
test_input[14624:14631] = '{32'h42bae559, 32'hc1c406c7, 32'h416df9d6, 32'hc222ed5d, 32'h42985056, 32'h41364a7f, 32'h42591895, 32'h42701416};
test_output[1828] = '{32'h42bae559};
test_index[1828] = '{0};
test_input[14632:14639] = '{32'h42bf8e8a, 32'hc2b8e5ec, 32'hc0b441f1, 32'hc296ef33, 32'h4174aae1, 32'hc29c0bfe, 32'h4242120d, 32'hc2534a66};
test_output[1829] = '{32'h42bf8e8a};
test_index[1829] = '{0};
test_input[14640:14647] = '{32'hc2990ac1, 32'h42713090, 32'h424398d1, 32'hc28bfd11, 32'hc2afb954, 32'h4187fd88, 32'h4291f54b, 32'h428b62fd};
test_output[1830] = '{32'h4291f54b};
test_index[1830] = '{6};
test_input[14648:14655] = '{32'h426bb497, 32'h42285596, 32'h4205b82e, 32'hc291915b, 32'h41050e53, 32'h4271c10c, 32'hc0193e05, 32'hc2c16539};
test_output[1831] = '{32'h4271c10c};
test_index[1831] = '{5};
test_input[14656:14663] = '{32'hc286d585, 32'hc12196ae, 32'h41cedbc0, 32'hc26eea29, 32'h401b7d01, 32'hc2af15ae, 32'hbf18b783, 32'h416fae97};
test_output[1832] = '{32'h41cedbc0};
test_index[1832] = '{2};
test_input[14664:14671] = '{32'h42bb3076, 32'hc038de39, 32'hc1ee5a07, 32'h41349f1a, 32'h42a5fe94, 32'hc26ea0bc, 32'hc24b0a06, 32'hc21e6f59};
test_output[1833] = '{32'h42bb3076};
test_index[1833] = '{0};
test_input[14672:14679] = '{32'hc28892f0, 32'h4031ff1b, 32'hc2b8bd16, 32'hc28c1bd9, 32'h42237a74, 32'h4240236a, 32'h42b3222d, 32'hc2a93609};
test_output[1834] = '{32'h42b3222d};
test_index[1834] = '{6};
test_input[14680:14687] = '{32'hc24c833c, 32'hc25c9b42, 32'h42c14198, 32'h40cdd5f4, 32'hc2896d51, 32'h428c1c03, 32'h421191f8, 32'hc26f15da};
test_output[1835] = '{32'h42c14198};
test_index[1835] = '{2};
test_input[14688:14695] = '{32'hc1d933f8, 32'h42009d11, 32'hc221b33b, 32'hc2651417, 32'h42b852bb, 32'hc28e5f3b, 32'hc2ae8122, 32'h42b05427};
test_output[1836] = '{32'h42b852bb};
test_index[1836] = '{4};
test_input[14696:14703] = '{32'h428fce64, 32'hc20ab7b9, 32'h429034b1, 32'hc1d0ec46, 32'h3e1baa75, 32'h42139b55, 32'h420c3cd8, 32'h42350749};
test_output[1837] = '{32'h429034b1};
test_index[1837] = '{2};
test_input[14704:14711] = '{32'h42c68769, 32'hc23fe023, 32'hc1d7a200, 32'hc2b08c25, 32'h414e9583, 32'h4299f1b2, 32'hc1f52327, 32'hc035652b};
test_output[1838] = '{32'h42c68769};
test_index[1838] = '{0};
test_input[14712:14719] = '{32'h3fca8e83, 32'hc2ac742b, 32'h423f212d, 32'hc1d624dd, 32'h4103f93a, 32'h40d462ec, 32'hc20479f8, 32'hbf67ab49};
test_output[1839] = '{32'h423f212d};
test_index[1839] = '{2};
test_input[14720:14727] = '{32'hc1a7506b, 32'h428e55ca, 32'h42a385d8, 32'h408b3698, 32'h423385f4, 32'hc253aab1, 32'hc2ad7f95, 32'h4233af39};
test_output[1840] = '{32'h42a385d8};
test_index[1840] = '{2};
test_input[14728:14735] = '{32'h42aa2a14, 32'hc28c0f4a, 32'hc27fed88, 32'h42624648, 32'hc266f8a5, 32'h413e48ab, 32'h42877e16, 32'hc1ad0c0b};
test_output[1841] = '{32'h42aa2a14};
test_index[1841] = '{0};
test_input[14736:14743] = '{32'hc233eaed, 32'hc00ec6f4, 32'h424fa8b4, 32'h4210c93d, 32'hc27f71c0, 32'hc24c8c3c, 32'hc14755c8, 32'h41f8bf32};
test_output[1842] = '{32'h424fa8b4};
test_index[1842] = '{2};
test_input[14744:14751] = '{32'hc17faa69, 32'hc253fc8e, 32'hc28f1ebf, 32'hc243ae69, 32'hc24d2e02, 32'h42a8b247, 32'h419b3531, 32'hc28db245};
test_output[1843] = '{32'h42a8b247};
test_index[1843] = '{5};
test_input[14752:14759] = '{32'h419fda75, 32'h42b7d728, 32'h42a8b5c5, 32'h407b6105, 32'hc289841c, 32'h424049b0, 32'h4291167b, 32'h4211afb9};
test_output[1844] = '{32'h42b7d728};
test_index[1844] = '{1};
test_input[14760:14767] = '{32'h4244704b, 32'hc26b502f, 32'hc2b145ce, 32'hc2262ee1, 32'h41861412, 32'hc0be22bc, 32'hc26b43e0, 32'h4266ff01};
test_output[1845] = '{32'h4266ff01};
test_index[1845] = '{7};
test_input[14768:14775] = '{32'hc28abd41, 32'h3f1e339a, 32'hc2946d8d, 32'hc257bd86, 32'hc21fde7d, 32'hc224d6f8, 32'hc234c300, 32'hc1fe7f6f};
test_output[1846] = '{32'h3f1e339a};
test_index[1846] = '{1};
test_input[14776:14783] = '{32'hc2b3b2c2, 32'h423bc931, 32'hc2690c55, 32'hc1408cbb, 32'h4221dc65, 32'hc2c6e15b, 32'h427227d9, 32'hc27a2a0c};
test_output[1847] = '{32'h427227d9};
test_index[1847] = '{6};
test_input[14784:14791] = '{32'hc0e0e9d1, 32'h41f28ad8, 32'hc08cb206, 32'hc24ec916, 32'hc2918d83, 32'hc227c798, 32'hc2bbed6b, 32'hc2883230};
test_output[1848] = '{32'h41f28ad8};
test_index[1848] = '{1};
test_input[14792:14799] = '{32'h42a6f121, 32'h4182e91f, 32'hc215ab1c, 32'h41b30848, 32'hc213ca96, 32'h407fa5c1, 32'h412ce58c, 32'h429a2055};
test_output[1849] = '{32'h42a6f121};
test_index[1849] = '{0};
test_input[14800:14807] = '{32'h42b55094, 32'h42b3cb62, 32'h40936a89, 32'hc29b56b0, 32'hc2489a61, 32'h42b765de, 32'hc2c16efa, 32'hc1c7c1e3};
test_output[1850] = '{32'h42b765de};
test_index[1850] = '{5};
test_input[14808:14815] = '{32'h425df6db, 32'h41fe0843, 32'h42525779, 32'hc2bfdce6, 32'h42affb2d, 32'h422bc9ca, 32'h42b59051, 32'h42a9a363};
test_output[1851] = '{32'h42b59051};
test_index[1851] = '{6};
test_input[14816:14823] = '{32'hc0fc8f56, 32'hc086ad51, 32'hc2a21d42, 32'hc1de2b00, 32'hc1c26cc5, 32'h4048c683, 32'hc288c8be, 32'hc28d3ee1};
test_output[1852] = '{32'h4048c683};
test_index[1852] = '{5};
test_input[14824:14831] = '{32'h4271b379, 32'hc2967cca, 32'h42c2076b, 32'h409266fa, 32'h428c4246, 32'hc2400635, 32'h426be4da, 32'hc2a2b747};
test_output[1853] = '{32'h42c2076b};
test_index[1853] = '{2};
test_input[14832:14839] = '{32'hc21e1eab, 32'hc2b31b0d, 32'hc1dc5c54, 32'hc2966af7, 32'h42b1b41b, 32'hc2795cf5, 32'h423a3d4e, 32'h4217f25b};
test_output[1854] = '{32'h42b1b41b};
test_index[1854] = '{4};
test_input[14840:14847] = '{32'hc117a584, 32'h425aa6b5, 32'hc2864cfd, 32'h41a8dcff, 32'hc23c24b6, 32'h412df1e3, 32'hc260c694, 32'hc26f72b3};
test_output[1855] = '{32'h425aa6b5};
test_index[1855] = '{1};
test_input[14848:14855] = '{32'h421c4971, 32'h4281a81c, 32'hc0b5bef1, 32'hc2194bfa, 32'hc0b58019, 32'h427961e4, 32'h4148447a, 32'hc273b1c4};
test_output[1856] = '{32'h4281a81c};
test_index[1856] = '{1};
test_input[14856:14863] = '{32'h41aed8a3, 32'hc28af23b, 32'hc2ac67b3, 32'hc2a29500, 32'h41ddc0e1, 32'hc0ec2596, 32'hc2bf556a, 32'h4289afd4};
test_output[1857] = '{32'h4289afd4};
test_index[1857] = '{7};
test_input[14864:14871] = '{32'hc2a17e1f, 32'hc2a01147, 32'hc2573c84, 32'h3eae5121, 32'h42a1bbcb, 32'hc2ab0835, 32'hc2b717d1, 32'h42b428fe};
test_output[1858] = '{32'h42b428fe};
test_index[1858] = '{7};
test_input[14872:14879] = '{32'h4216469a, 32'h42c3b9a1, 32'h42b6ecc5, 32'h428f2640, 32'hc2699a3c, 32'hc2556767, 32'h413f25e9, 32'h40bebe3c};
test_output[1859] = '{32'h42c3b9a1};
test_index[1859] = '{1};
test_input[14880:14887] = '{32'hc2b310e2, 32'h41da317c, 32'hc1dfe79b, 32'h41aae65c, 32'h42c50a3f, 32'h42a44cf8, 32'hc1291799, 32'hc0c1bffc};
test_output[1860] = '{32'h42c50a3f};
test_index[1860] = '{4};
test_input[14888:14895] = '{32'h40fb2ed9, 32'h4288fe60, 32'hc080bf4a, 32'h428a04e2, 32'h41b1d829, 32'hc20a69a5, 32'hc28f3059, 32'hc28899ef};
test_output[1861] = '{32'h428a04e2};
test_index[1861] = '{3};
test_input[14896:14903] = '{32'hc185bad6, 32'hc0bb7ff9, 32'h42b66e7b, 32'h4117df38, 32'hc25cb156, 32'h410ab25f, 32'h41682229, 32'h42399cab};
test_output[1862] = '{32'h42b66e7b};
test_index[1862] = '{2};
test_input[14904:14911] = '{32'h4162ce0e, 32'h42a81586, 32'hc0e1edc5, 32'h42a22196, 32'h42b3375b, 32'hc1d44387, 32'hc062c8c6, 32'hc275ff99};
test_output[1863] = '{32'h42b3375b};
test_index[1863] = '{4};
test_input[14912:14919] = '{32'hc24710eb, 32'h42702730, 32'h41de2b44, 32'h41ad91d4, 32'hc26bff23, 32'h42bc6f71, 32'h42c0d8a3, 32'hc16cb366};
test_output[1864] = '{32'h42c0d8a3};
test_index[1864] = '{6};
test_input[14920:14927] = '{32'h42a8e634, 32'hc2c6b51f, 32'hc22e5c22, 32'hc2be7025, 32'h419cbe95, 32'hc202e90d, 32'h4222268f, 32'h4194fdb2};
test_output[1865] = '{32'h42a8e634};
test_index[1865] = '{0};
test_input[14928:14935] = '{32'hc15d44ae, 32'h42878213, 32'hc2b97f29, 32'hc266911a, 32'h41c445be, 32'hc20d03a1, 32'h40c17416, 32'h429060f5};
test_output[1866] = '{32'h429060f5};
test_index[1866] = '{7};
test_input[14936:14943] = '{32'h41c234f3, 32'hc1cf8dd1, 32'hc2933283, 32'hc2ad14be, 32'h409a32b1, 32'hc2bb087d, 32'h42b78134, 32'hc2442e68};
test_output[1867] = '{32'h42b78134};
test_index[1867] = '{6};
test_input[14944:14951] = '{32'hc1c2aa3d, 32'h422e2ac3, 32'hc2033f85, 32'hc1d0de9d, 32'h425b3e8f, 32'h428ecfe9, 32'h423aa03b, 32'h42844654};
test_output[1868] = '{32'h428ecfe9};
test_index[1868] = '{5};
test_input[14952:14959] = '{32'h42849933, 32'h42bc9127, 32'hc161d5fc, 32'hc2be22e8, 32'h426b8e23, 32'h42081531, 32'hc12b8be0, 32'hc1e21424};
test_output[1869] = '{32'h42bc9127};
test_index[1869] = '{1};
test_input[14960:14967] = '{32'hc240f002, 32'hc2c4c66c, 32'h42b5747d, 32'hc2a19580, 32'hc2bfb2c8, 32'hc2408d06, 32'hc29f574b, 32'hc0e7cb4b};
test_output[1870] = '{32'h42b5747d};
test_index[1870] = '{2};
test_input[14968:14975] = '{32'hc2815963, 32'hc2992360, 32'h411c8a6e, 32'h42bc0761, 32'h3fdfead4, 32'hc2a051aa, 32'hc2ad0067, 32'hc20ffc31};
test_output[1871] = '{32'h42bc0761};
test_index[1871] = '{3};
test_input[14976:14983] = '{32'h41f18d17, 32'h421034f1, 32'hc1b02e25, 32'hc262131e, 32'hc2b6a11a, 32'h41535123, 32'h4031e757, 32'hc2bb3454};
test_output[1872] = '{32'h421034f1};
test_index[1872] = '{1};
test_input[14984:14991] = '{32'h417f138c, 32'hbfb56feb, 32'hc083fe80, 32'hc1bac33e, 32'h42661aff, 32'hc1a43bba, 32'h4276a0a0, 32'h42538741};
test_output[1873] = '{32'h4276a0a0};
test_index[1873] = '{6};
test_input[14992:14999] = '{32'hc229ef4f, 32'h41beabe2, 32'hc2b9783c, 32'h41bf89ef, 32'h420e2f5a, 32'hc209c6c1, 32'hc253e9da, 32'h412c2c5d};
test_output[1874] = '{32'h420e2f5a};
test_index[1874] = '{4};
test_input[15000:15007] = '{32'h41ec8b83, 32'h42b359c2, 32'h42187c25, 32'hc2976c25, 32'h3f227e7a, 32'h42437a26, 32'h42c46b58, 32'h42741ec6};
test_output[1875] = '{32'h42c46b58};
test_index[1875] = '{6};
test_input[15008:15015] = '{32'hc299b9e3, 32'hc224e1e4, 32'h42310529, 32'h42032dc9, 32'h4298252a, 32'hc277235a, 32'h4171d7e3, 32'hc173fc62};
test_output[1876] = '{32'h4298252a};
test_index[1876] = '{4};
test_input[15016:15023] = '{32'h4297cb34, 32'hc28d44bd, 32'h42a13fee, 32'hc28b0bd1, 32'h4270d7b2, 32'h41a3487b, 32'hc2bb0ae2, 32'hc1d00983};
test_output[1877] = '{32'h42a13fee};
test_index[1877] = '{2};
test_input[15024:15031] = '{32'h4283edd1, 32'h42b7262d, 32'hc21e8592, 32'h42bef118, 32'hc273e056, 32'hc1c07c91, 32'h409c757a, 32'h418afcbc};
test_output[1878] = '{32'h42bef118};
test_index[1878] = '{3};
test_input[15032:15039] = '{32'hc24abff4, 32'hc2c0df26, 32'hc1b10172, 32'h408b2426, 32'hc1d81cc6, 32'h42673e5a, 32'hc2853948, 32'hc1b5eb7e};
test_output[1879] = '{32'h42673e5a};
test_index[1879] = '{5};
test_input[15040:15047] = '{32'hc11358db, 32'h428b12d9, 32'hc2074196, 32'h4278ae9c, 32'hc0d73825, 32'h424d4528, 32'h42047429, 32'h42a09d1f};
test_output[1880] = '{32'h42a09d1f};
test_index[1880] = '{7};
test_input[15048:15055] = '{32'hc2190196, 32'h42b5dff6, 32'hc19c4190, 32'hc2b1e5bf, 32'hc1a11bcb, 32'h42bc12a8, 32'h421f2490, 32'hc10a3dfe};
test_output[1881] = '{32'h42bc12a8};
test_index[1881] = '{5};
test_input[15056:15063] = '{32'h41f94d54, 32'h4204d4c5, 32'hc2630b9a, 32'h40904b5d, 32'hc2c24d09, 32'hc1bfb000, 32'hc2066abf, 32'h42947121};
test_output[1882] = '{32'h42947121};
test_index[1882] = '{7};
test_input[15064:15071] = '{32'hc23efec1, 32'hc2474958, 32'hbb1f4ea4, 32'hc29675c4, 32'hc2b5df2a, 32'hc2810186, 32'hc066b231, 32'h428014ba};
test_output[1883] = '{32'h428014ba};
test_index[1883] = '{7};
test_input[15072:15079] = '{32'h42122054, 32'hc271665b, 32'hc1ae7a88, 32'hc233d013, 32'hc2274d37, 32'hc1eb3b40, 32'h42bb7c9e, 32'h4292e746};
test_output[1884] = '{32'h42bb7c9e};
test_index[1884] = '{6};
test_input[15080:15087] = '{32'h40b4c534, 32'h4190f3b4, 32'h429829f5, 32'h4284e44d, 32'h42aab13d, 32'h42334746, 32'hc086a7c4, 32'h41fc90b7};
test_output[1885] = '{32'h42aab13d};
test_index[1885] = '{4};
test_input[15088:15095] = '{32'h4144f4ee, 32'h42af4089, 32'h42095717, 32'h42944fd0, 32'hc29ad469, 32'hc29a6730, 32'h41de57b4, 32'h42c05bf7};
test_output[1886] = '{32'h42c05bf7};
test_index[1886] = '{7};
test_input[15096:15103] = '{32'hc292242e, 32'h4284bd7c, 32'hc292ddf2, 32'hc25ec250, 32'h42953d69, 32'h40958b28, 32'h4291f3e1, 32'hc2130cc1};
test_output[1887] = '{32'h42953d69};
test_index[1887] = '{4};
test_input[15104:15111] = '{32'h42b87fde, 32'hc2994788, 32'hc28a55ad, 32'hbff1807e, 32'h3ff25a2f, 32'h422c84c3, 32'hc2bd960c, 32'h42874e22};
test_output[1888] = '{32'h42b87fde};
test_index[1888] = '{0};
test_input[15112:15119] = '{32'h419e60ef, 32'hc2af2864, 32'h41c3cd3a, 32'h426b4c79, 32'hc2146a74, 32'hc2c125a0, 32'h425d4296, 32'h426b1416};
test_output[1889] = '{32'h426b4c79};
test_index[1889] = '{3};
test_input[15120:15127] = '{32'hc2a9f1d8, 32'h42b7ea2a, 32'h42b70161, 32'h41c2430c, 32'hc260c6c0, 32'hc2bbcb1d, 32'hc20a6ef6, 32'hc2c0ef11};
test_output[1890] = '{32'h42b7ea2a};
test_index[1890] = '{1};
test_input[15128:15135] = '{32'h4253b9cf, 32'h40d4f837, 32'h42b3f1bb, 32'h423f96c9, 32'hc2b95293, 32'h42206232, 32'h42a02c81, 32'h42a7c4ff};
test_output[1891] = '{32'h42b3f1bb};
test_index[1891] = '{2};
test_input[15136:15143] = '{32'hc237f2b8, 32'h42b65222, 32'h4286f052, 32'h42bc7e64, 32'h421bb5ee, 32'h42a67849, 32'h42b09ac7, 32'hc255c4c1};
test_output[1892] = '{32'h42bc7e64};
test_index[1892] = '{3};
test_input[15144:15151] = '{32'h429e0c88, 32'h42c60438, 32'hc18bb15c, 32'h42545311, 32'h41aa7221, 32'hc2c4a5df, 32'h41bb767d, 32'h42b10437};
test_output[1893] = '{32'h42c60438};
test_index[1893] = '{1};
test_input[15152:15159] = '{32'h41cd4d35, 32'hc2a0ed82, 32'hc1e50b05, 32'hc261f3b2, 32'hc2890578, 32'h42677b44, 32'h418a3d12, 32'hc20f098a};
test_output[1894] = '{32'h42677b44};
test_index[1894] = '{5};
test_input[15160:15167] = '{32'hc28ba163, 32'h406d9c03, 32'h4253c149, 32'h42b4c45f, 32'h41254a6e, 32'hc2bc7947, 32'hc230164f, 32'h41e4adb0};
test_output[1895] = '{32'h42b4c45f};
test_index[1895] = '{3};
test_input[15168:15175] = '{32'h42159b24, 32'hc1b7e343, 32'h425207ed, 32'h42a74637, 32'hc2b42b18, 32'hc2c547b8, 32'h42034570, 32'hc1a9befd};
test_output[1896] = '{32'h42a74637};
test_index[1896] = '{3};
test_input[15176:15183] = '{32'h4234fe4e, 32'hc2a06731, 32'h4258bdd3, 32'h41bad5df, 32'h42804d75, 32'hc2314aab, 32'h40acb15e, 32'hc1cca015};
test_output[1897] = '{32'h42804d75};
test_index[1897] = '{4};
test_input[15184:15191] = '{32'hc1ec8917, 32'hc22bd88f, 32'hc28dc585, 32'hc18e5b47, 32'h42b429a4, 32'hc272dd91, 32'hc27367db, 32'hc13f5034};
test_output[1898] = '{32'h42b429a4};
test_index[1898] = '{4};
test_input[15192:15199] = '{32'h429a82b0, 32'hc1afbe31, 32'h4287bea3, 32'h42839de6, 32'hc2b8c530, 32'h41953e3b, 32'h41f21aa3, 32'hc1092ab1};
test_output[1899] = '{32'h429a82b0};
test_index[1899] = '{0};
test_input[15200:15207] = '{32'h41ba20cb, 32'hc2586bdf, 32'hc09f5cf9, 32'hc07aa81b, 32'hc197ff4e, 32'h41ffc824, 32'h4231b898, 32'hc2ae1e8f};
test_output[1900] = '{32'h4231b898};
test_index[1900] = '{6};
test_input[15208:15215] = '{32'hc2c70c0c, 32'h42c7c7b7, 32'h4046abf5, 32'h41f7cf79, 32'h42c0b496, 32'hc2aa8d6e, 32'hc276aeef, 32'h409f5e65};
test_output[1901] = '{32'h42c7c7b7};
test_index[1901] = '{1};
test_input[15216:15223] = '{32'h425769c2, 32'h42a44553, 32'h40f9c966, 32'h42b2542e, 32'hc27721be, 32'hc2a68f9a, 32'h4233d1b1, 32'hc28a2382};
test_output[1902] = '{32'h42b2542e};
test_index[1902] = '{3};
test_input[15224:15231] = '{32'h4267d1d7, 32'h41382472, 32'hc2690c0d, 32'h425d01f6, 32'hc2c44033, 32'hc2234085, 32'hc285d1d8, 32'h4279a281};
test_output[1903] = '{32'h4279a281};
test_index[1903] = '{7};
test_input[15232:15239] = '{32'hbe8e3808, 32'hc2af86d7, 32'h419d419e, 32'h428f0f0d, 32'h41e09add, 32'h428a8abd, 32'h421eca24, 32'hc06a27c5};
test_output[1904] = '{32'h428f0f0d};
test_index[1904] = '{3};
test_input[15240:15247] = '{32'hc19a5835, 32'h428c482f, 32'hc20efbc3, 32'h42b1aca2, 32'hc22fa80a, 32'h427b64be, 32'h3d69d5bb, 32'hc1b3bb61};
test_output[1905] = '{32'h42b1aca2};
test_index[1905] = '{3};
test_input[15248:15255] = '{32'h422e9e1f, 32'hc293bd77, 32'h420187ce, 32'hc234274e, 32'h429dce70, 32'h422467ed, 32'h423d584d, 32'h42357d9b};
test_output[1906] = '{32'h429dce70};
test_index[1906] = '{4};
test_input[15256:15263] = '{32'hc16b5205, 32'h41f9d85d, 32'h42a9c376, 32'h42b1f6ea, 32'hc2963e31, 32'hc217f3db, 32'hc20d4b22, 32'hc1d0792f};
test_output[1907] = '{32'h42b1f6ea};
test_index[1907] = '{3};
test_input[15264:15271] = '{32'hc25d3ecb, 32'h429c3a6a, 32'hc2613038, 32'h422f2a02, 32'hc206868a, 32'h4288b425, 32'hc20c9453, 32'h42c504ed};
test_output[1908] = '{32'h42c504ed};
test_index[1908] = '{7};
test_input[15272:15279] = '{32'hc2b94a12, 32'h428506b1, 32'h4236df9b, 32'hc1cacd0d, 32'h41486848, 32'h42aef847, 32'hc27fc792, 32'h425a7ca2};
test_output[1909] = '{32'h42aef847};
test_index[1909] = '{5};
test_input[15280:15287] = '{32'h42c13c3b, 32'h427b29e6, 32'h4251e186, 32'h427c66c2, 32'hc22cffb7, 32'h4293d0e9, 32'hc23b103d, 32'h41eb95d4};
test_output[1910] = '{32'h42c13c3b};
test_index[1910] = '{0};
test_input[15288:15295] = '{32'h42371102, 32'hc1d1de7a, 32'hc1dcf06c, 32'hc1c93535, 32'h42700b52, 32'h4209e4cc, 32'hc1878925, 32'h41dd8228};
test_output[1911] = '{32'h42700b52};
test_index[1911] = '{4};
test_input[15296:15303] = '{32'hc0cecb69, 32'h428266ae, 32'hc23ee62b, 32'hc22164f2, 32'h4297efc5, 32'hc252aaff, 32'h426bb0e2, 32'hc2c3978c};
test_output[1912] = '{32'h4297efc5};
test_index[1912] = '{4};
test_input[15304:15311] = '{32'hc1a5cafb, 32'hc2a52829, 32'h427f5ccd, 32'h42a4a44f, 32'h4119ad23, 32'h428d70ca, 32'h4262a4cd, 32'hc1b8e4a1};
test_output[1913] = '{32'h42a4a44f};
test_index[1913] = '{3};
test_input[15312:15319] = '{32'h42b17529, 32'h42032cf9, 32'hc29d1c23, 32'hc288359c, 32'h423ecd2d, 32'h42a2229d, 32'hc2946092, 32'h40a76383};
test_output[1914] = '{32'h42b17529};
test_index[1914] = '{0};
test_input[15320:15327] = '{32'h42b08702, 32'hc228b39a, 32'h42a9a88f, 32'h426d2eb5, 32'hc2101ad1, 32'h42b0db63, 32'h42bc7b4b, 32'hc28c05c6};
test_output[1915] = '{32'h42bc7b4b};
test_index[1915] = '{6};
test_input[15328:15335] = '{32'h4259d0c2, 32'h4249771b, 32'hc1d14f5a, 32'hc28a5490, 32'h42bc3c65, 32'h4259648e, 32'hc298e731, 32'h425e042c};
test_output[1916] = '{32'h42bc3c65};
test_index[1916] = '{4};
test_input[15336:15343] = '{32'h42921f43, 32'hc1b345ca, 32'h4240b355, 32'h425dec0a, 32'hc2b2a453, 32'h429ddd31, 32'hc29d71d2, 32'hc1373e1f};
test_output[1917] = '{32'h429ddd31};
test_index[1917] = '{5};
test_input[15344:15351] = '{32'hc23641cd, 32'h414f6102, 32'hc2b3872e, 32'h42aace2d, 32'h42be35d0, 32'hc1de976d, 32'h427b7e26, 32'h42141e24};
test_output[1918] = '{32'h42be35d0};
test_index[1918] = '{4};
test_input[15352:15359] = '{32'h421b572f, 32'h42c02569, 32'hc22e3fd4, 32'h4231ece1, 32'h40792061, 32'hc2bf5825, 32'hc20f4f9b, 32'h428de0a2};
test_output[1919] = '{32'h42c02569};
test_index[1919] = '{1};
test_input[15360:15367] = '{32'hc28a6470, 32'h41efe42d, 32'h428a20d7, 32'hc2bedb65, 32'h42b14efd, 32'h4257cf8a, 32'hc1f7dcff, 32'h41e207e5};
test_output[1920] = '{32'h42b14efd};
test_index[1920] = '{4};
test_input[15368:15375] = '{32'h40e40c3d, 32'hc2912427, 32'h42b677c4, 32'h428ff2ce, 32'hc2c28c16, 32'h42944783, 32'h4288302e, 32'hc2c492ab};
test_output[1921] = '{32'h42b677c4};
test_index[1921] = '{2};
test_input[15376:15383] = '{32'h42745566, 32'hc26f2b2c, 32'hc2274289, 32'hc19be64a, 32'hc1ff56a9, 32'hc006404a, 32'hc293d637, 32'h42a4feac};
test_output[1922] = '{32'h42a4feac};
test_index[1922] = '{7};
test_input[15384:15391] = '{32'hc2c5db07, 32'hc249d159, 32'hc000adab, 32'hc17a087a, 32'h42c041a9, 32'h42a41b9d, 32'hc1d3637f, 32'h3ec3030a};
test_output[1923] = '{32'h42c041a9};
test_index[1923] = '{4};
test_input[15392:15399] = '{32'hc205d870, 32'hc146fba6, 32'hc1f190de, 32'h429fa6cc, 32'hc2506d37, 32'h42a05053, 32'hc28439b4, 32'hc1d3d944};
test_output[1924] = '{32'h42a05053};
test_index[1924] = '{5};
test_input[15400:15407] = '{32'h41aaf0e4, 32'hc120317a, 32'hc280fe24, 32'hc1c19aef, 32'h40e3ce49, 32'h42711137, 32'hc29c19ac, 32'hc20d47d7};
test_output[1925] = '{32'h42711137};
test_index[1925] = '{5};
test_input[15408:15415] = '{32'hc1fedda4, 32'hc2a604d1, 32'h41f63ef4, 32'h42b57dde, 32'hc101be01, 32'h42873030, 32'h42800b65, 32'hc1a9e3dc};
test_output[1926] = '{32'h42b57dde};
test_index[1926] = '{3};
test_input[15416:15423] = '{32'hc2815244, 32'h41a99e0d, 32'hc2a2bc2b, 32'hc23f6347, 32'hc1c1a182, 32'h3fd80973, 32'h42204e50, 32'hc208d6ed};
test_output[1927] = '{32'h42204e50};
test_index[1927] = '{6};
test_input[15424:15431] = '{32'h4274b32f, 32'hc2ba43f9, 32'h4119025e, 32'h42ab6b03, 32'h422b4d76, 32'hc2b52edc, 32'h42643bc5, 32'h41883247};
test_output[1928] = '{32'h42ab6b03};
test_index[1928] = '{3};
test_input[15432:15439] = '{32'h40a6b941, 32'hc1a7d357, 32'hc20a095e, 32'h42a7255c, 32'hc2a522c4, 32'h42930a94, 32'h3d9a8db7, 32'hc1420e0e};
test_output[1929] = '{32'h42a7255c};
test_index[1929] = '{3};
test_input[15440:15447] = '{32'h4240837d, 32'h422183e1, 32'h40ba68e1, 32'h4206129a, 32'hc2024174, 32'h41e7f581, 32'hc2b6bffb, 32'h4269d2ed};
test_output[1930] = '{32'h4269d2ed};
test_index[1930] = '{7};
test_input[15448:15455] = '{32'hc2193d26, 32'hc275a8fc, 32'h42c6b70e, 32'h41997889, 32'hc28e2a06, 32'hc20e28d9, 32'h41cc84d2, 32'h42c50e20};
test_output[1931] = '{32'h42c6b70e};
test_index[1931] = '{2};
test_input[15456:15463] = '{32'hc2b56931, 32'hc274d723, 32'h42394d38, 32'h42a3dac5, 32'hc1e90b8e, 32'h415c983e, 32'h42a88718, 32'h4289b807};
test_output[1932] = '{32'h42a88718};
test_index[1932] = '{6};
test_input[15464:15471] = '{32'h42822f5e, 32'hc2bdf191, 32'hc28b5d80, 32'h422b3d56, 32'hc2625816, 32'hc28a6719, 32'h42ac0f3d, 32'hc2a3211a};
test_output[1933] = '{32'h42ac0f3d};
test_index[1933] = '{6};
test_input[15472:15479] = '{32'hc0fb7d55, 32'h41ddff98, 32'hc20b19cc, 32'h41f5ebfa, 32'hc28592d8, 32'hc2bb1fdc, 32'hc18a9cc6, 32'hc23fd420};
test_output[1934] = '{32'h41f5ebfa};
test_index[1934] = '{3};
test_input[15480:15487] = '{32'hc2aa48d9, 32'hc292a159, 32'h429a8b04, 32'h422ec050, 32'h42b3f85a, 32'h4176ca17, 32'h427f83e8, 32'h3fbb8627};
test_output[1935] = '{32'h42b3f85a};
test_index[1935] = '{4};
test_input[15488:15495] = '{32'hc28ff96d, 32'h3f107d31, 32'hc233e0de, 32'h417b2e05, 32'hc26832d3, 32'hc179859f, 32'hc208eab4, 32'h42735a4b};
test_output[1936] = '{32'h42735a4b};
test_index[1936] = '{7};
test_input[15496:15503] = '{32'hc282b4e6, 32'h422b13aa, 32'h42bb283b, 32'hc29d43c5, 32'hc2b8bedf, 32'hc2bc2beb, 32'h426ae8b3, 32'h4256ed7e};
test_output[1937] = '{32'h42bb283b};
test_index[1937] = '{2};
test_input[15504:15511] = '{32'hc1e62764, 32'hc1070630, 32'hc22ae083, 32'h42bdf46d, 32'hc29501d2, 32'h42aafd0d, 32'hc19fa795, 32'h42a9c9a6};
test_output[1938] = '{32'h42bdf46d};
test_index[1938] = '{3};
test_input[15512:15519] = '{32'hc2b64606, 32'hc2afe443, 32'h42bea06b, 32'h414e845d, 32'h428755b2, 32'h4198f648, 32'hc2c14d6e, 32'h428c6fd9};
test_output[1939] = '{32'h42bea06b};
test_index[1939] = '{2};
test_input[15520:15527] = '{32'hc1f4ac5b, 32'hc1e0ec90, 32'h40fead89, 32'h42c02acd, 32'hc27696af, 32'h424a809e, 32'h426f8d66, 32'h4204d83d};
test_output[1940] = '{32'h42c02acd};
test_index[1940] = '{3};
test_input[15528:15535] = '{32'hc2509477, 32'h41ad688d, 32'h42385021, 32'h421be0bb, 32'hc29e66b9, 32'h427027ae, 32'hc28203bb, 32'h427b06e7};
test_output[1941] = '{32'h427b06e7};
test_index[1941] = '{7};
test_input[15536:15543] = '{32'hc262ae03, 32'h41867b6a, 32'h42a9e3b1, 32'hc29d42f7, 32'h422f0092, 32'hc28d3d6f, 32'hbf473ba0, 32'h41c636fd};
test_output[1942] = '{32'h42a9e3b1};
test_index[1942] = '{2};
test_input[15544:15551] = '{32'h42c23eb5, 32'hc2778411, 32'h41e656b8, 32'h423ea091, 32'hc28a85ab, 32'hc2405da9, 32'h429eea1f, 32'h426e6b88};
test_output[1943] = '{32'h42c23eb5};
test_index[1943] = '{0};
test_input[15552:15559] = '{32'h4233de2b, 32'h42bb890f, 32'h42412062, 32'h413748a5, 32'hc2c515f4, 32'hc2a98c48, 32'hc2350afb, 32'h4284df9b};
test_output[1944] = '{32'h42bb890f};
test_index[1944] = '{1};
test_input[15560:15567] = '{32'h421c3964, 32'hc1aa4c1f, 32'h428a70c3, 32'hc28a9071, 32'hc29ec055, 32'h412b1b9c, 32'h40f56860, 32'hc0a92709};
test_output[1945] = '{32'h428a70c3};
test_index[1945] = '{2};
test_input[15568:15575] = '{32'h42334dcd, 32'h4005a0ad, 32'hc2450b7c, 32'hc115ae68, 32'h426e69f0, 32'hc2acba09, 32'h418c1e48, 32'hc29bbe36};
test_output[1946] = '{32'h426e69f0};
test_index[1946] = '{4};
test_input[15576:15583] = '{32'hc2a30778, 32'h4139557c, 32'h41a9aaf6, 32'h3ff93e25, 32'hc1857f1c, 32'h4209968b, 32'h429ba3e0, 32'h428309ad};
test_output[1947] = '{32'h429ba3e0};
test_index[1947] = '{6};
test_input[15584:15591] = '{32'h4297d429, 32'hc2b367b0, 32'hc0b700c5, 32'hbf8bcbfe, 32'hc1d4a3b7, 32'hc2851b87, 32'h42b1f7d5, 32'h429dd253};
test_output[1948] = '{32'h42b1f7d5};
test_index[1948] = '{6};
test_input[15592:15599] = '{32'h40ef694e, 32'hc2b80e20, 32'h4191e844, 32'h4290a39a, 32'h42184148, 32'h41ba6771, 32'h42a93ae3, 32'hc1f57380};
test_output[1949] = '{32'h42a93ae3};
test_index[1949] = '{6};
test_input[15600:15607] = '{32'hc219ad87, 32'hc285876f, 32'hc2b28b57, 32'hc29ec70d, 32'h414365f5, 32'hc2970390, 32'hc1cb3a2f, 32'h40f571a1};
test_output[1950] = '{32'h414365f5};
test_index[1950] = '{4};
test_input[15608:15615] = '{32'h428d132c, 32'hc26d3925, 32'h41b79cc7, 32'h42a322b5, 32'hc2809b59, 32'hc07170c0, 32'h4178d9bc, 32'hc28adfca};
test_output[1951] = '{32'h42a322b5};
test_index[1951] = '{3};
test_input[15616:15623] = '{32'h41a90d2a, 32'hc2c1067c, 32'h4272b5ed, 32'h41b3f605, 32'h41fec6db, 32'h41c2d9ab, 32'hc21b8667, 32'hc12edd2f};
test_output[1952] = '{32'h4272b5ed};
test_index[1952] = '{2};
test_input[15624:15631] = '{32'h4244767e, 32'h425d38cd, 32'hc11c1740, 32'hc2aa6e2b, 32'h42bc1b96, 32'h42bb8c15, 32'hc283ee4d, 32'hc2870553};
test_output[1953] = '{32'h42bc1b96};
test_index[1953] = '{4};
test_input[15632:15639] = '{32'hc2c1c651, 32'hc2bee9a8, 32'hc2448f38, 32'hc282e1a4, 32'hc24bf801, 32'h4245f103, 32'hc1c112e9, 32'hc2c0f4d1};
test_output[1954] = '{32'h4245f103};
test_index[1954] = '{5};
test_input[15640:15647] = '{32'hc23f8f5a, 32'h42afc885, 32'h4216e075, 32'hc226eef4, 32'hc11e8fee, 32'hc1bde6e5, 32'hc22876b5, 32'h42b3906c};
test_output[1955] = '{32'h42b3906c};
test_index[1955] = '{7};
test_input[15648:15655] = '{32'h422f2408, 32'hc105b314, 32'h42b0cf15, 32'hc2bd606f, 32'hc2983b98, 32'hc1c4c887, 32'h410324d6, 32'hc2873ab8};
test_output[1956] = '{32'h42b0cf15};
test_index[1956] = '{2};
test_input[15656:15663] = '{32'h41a68e8a, 32'hc2ab087f, 32'h42be5801, 32'h4251805b, 32'hc2c5d465, 32'hc1ea7196, 32'h42776b6e, 32'h42b73741};
test_output[1957] = '{32'h42be5801};
test_index[1957] = '{2};
test_input[15664:15671] = '{32'h427eb8fb, 32'hbe44412b, 32'h42915d83, 32'h408800cf, 32'h42b76dbd, 32'hc1bb763e, 32'h4279fddc, 32'hc140c248};
test_output[1958] = '{32'h42b76dbd};
test_index[1958] = '{4};
test_input[15672:15679] = '{32'h41f1bd20, 32'hc2bcfbb4, 32'h42bdd5d5, 32'hc1d78cdb, 32'hc2185052, 32'hc1ac79ce, 32'hc2b352b1, 32'hc2795618};
test_output[1959] = '{32'h42bdd5d5};
test_index[1959] = '{2};
test_input[15680:15687] = '{32'hc240c242, 32'h41d09cd2, 32'hc2720008, 32'hc150d2bb, 32'hc274a15e, 32'h42ab4dab, 32'h3e108b8f, 32'h4266d631};
test_output[1960] = '{32'h42ab4dab};
test_index[1960] = '{5};
test_input[15688:15695] = '{32'hc2b9f6b3, 32'hc0cb7a52, 32'h42053d02, 32'h427567b9, 32'h42b87f99, 32'hc0f7de47, 32'h4295cbce, 32'hc2a55fed};
test_output[1961] = '{32'h42b87f99};
test_index[1961] = '{4};
test_input[15696:15703] = '{32'hc1de4abe, 32'h4119ce45, 32'h4281773a, 32'h41a0677a, 32'h420a84e7, 32'h428f5962, 32'h422e2406, 32'hc25efd8e};
test_output[1962] = '{32'h428f5962};
test_index[1962] = '{5};
test_input[15704:15711] = '{32'h41de1498, 32'hc2bf6be7, 32'h42191333, 32'h424ea15c, 32'h42269f27, 32'h41927cb6, 32'hc1d5119c, 32'hc1899259};
test_output[1963] = '{32'h424ea15c};
test_index[1963] = '{3};
test_input[15712:15719] = '{32'hc296fa3d, 32'hc27cfcad, 32'h41e294d9, 32'h4227f0ba, 32'hc2a28e28, 32'h42959b8e, 32'hc2250072, 32'hc0e9c176};
test_output[1964] = '{32'h42959b8e};
test_index[1964] = '{5};
test_input[15720:15727] = '{32'h426ec199, 32'hc2994558, 32'hc28d73d0, 32'hc296dfa9, 32'hc29d5a2e, 32'hc1890d70, 32'hc29b1ed2, 32'h42c694ec};
test_output[1965] = '{32'h42c694ec};
test_index[1965] = '{7};
test_input[15728:15735] = '{32'h42ba1239, 32'h416447e2, 32'hc032a27a, 32'hc233b29b, 32'h428fed42, 32'hc2340ca6, 32'h4247700c, 32'h420c2258};
test_output[1966] = '{32'h42ba1239};
test_index[1966] = '{0};
test_input[15736:15743] = '{32'hc285c623, 32'h42bdb26c, 32'h426e4d2d, 32'hc1bf23ae, 32'hc14c5751, 32'hc26e0aec, 32'h4211ffdc, 32'hc17afc68};
test_output[1967] = '{32'h42bdb26c};
test_index[1967] = '{1};
test_input[15744:15751] = '{32'h42687862, 32'hc1c74b00, 32'h4229e6ae, 32'h4208e26d, 32'hc114af5f, 32'hc2b606f0, 32'h40e9fdb9, 32'hc2436831};
test_output[1968] = '{32'h42687862};
test_index[1968] = '{0};
test_input[15752:15759] = '{32'hc20f5128, 32'hc263f04e, 32'hc28f22a1, 32'h42674798, 32'h4283f64a, 32'h4231cefe, 32'hc1f5dbc8, 32'h42b7de18};
test_output[1969] = '{32'h42b7de18};
test_index[1969] = '{7};
test_input[15760:15767] = '{32'hc2b4055d, 32'hc202e65d, 32'h426719f8, 32'hc1d17edc, 32'h42a35459, 32'h422f2287, 32'hc156f715, 32'hc2a12ac2};
test_output[1970] = '{32'h42a35459};
test_index[1970] = '{4};
test_input[15768:15775] = '{32'hc294c1bc, 32'hc2c34d0a, 32'h42c30fa6, 32'h4289ab8c, 32'hc24cb329, 32'h420df5d0, 32'hc23a2b08, 32'hc1aea23c};
test_output[1971] = '{32'h42c30fa6};
test_index[1971] = '{2};
test_input[15776:15783] = '{32'hc26aeac4, 32'h42813f37, 32'hc1de3adc, 32'h41a263ee, 32'h42bb8a86, 32'hc1dceec8, 32'hc2428bb0, 32'hc0e003f9};
test_output[1972] = '{32'h42bb8a86};
test_index[1972] = '{4};
test_input[15784:15791] = '{32'h4058f65c, 32'hc1ccaab0, 32'hc27d67fc, 32'h42bcb162, 32'h422294dc, 32'hc2c1ba20, 32'hc1c992dd, 32'hc29db6ed};
test_output[1973] = '{32'h42bcb162};
test_index[1973] = '{3};
test_input[15792:15799] = '{32'h42ae802f, 32'h42c3ae43, 32'h3fab0558, 32'hc135a491, 32'hc2a34128, 32'h4241a685, 32'hc1a90173, 32'h4222e536};
test_output[1974] = '{32'h42c3ae43};
test_index[1974] = '{1};
test_input[15800:15807] = '{32'h4287bd1f, 32'h42138e17, 32'hc28d2994, 32'hc27b45b4, 32'hc1336cfc, 32'h41eee828, 32'h421bafed, 32'hc2af57d5};
test_output[1975] = '{32'h4287bd1f};
test_index[1975] = '{0};
test_input[15808:15815] = '{32'h42a0b216, 32'h40f94663, 32'hbf66ceca, 32'hc09b3700, 32'h42699175, 32'h42b98eb2, 32'hc214de50, 32'hc26bf836};
test_output[1976] = '{32'h42b98eb2};
test_index[1976] = '{5};
test_input[15816:15823] = '{32'h415d0df7, 32'h3f30c296, 32'hc27f146f, 32'h420c92ff, 32'hc27a7350, 32'h4157ae7d, 32'h41800c25, 32'hc23cbd3b};
test_output[1977] = '{32'h420c92ff};
test_index[1977] = '{3};
test_input[15824:15831] = '{32'h4114ab5b, 32'h420b590e, 32'hc2b1e375, 32'h42b3d6c6, 32'hc1c8f3fa, 32'h41cbd117, 32'h422d6ac9, 32'h420f87c4};
test_output[1978] = '{32'h42b3d6c6};
test_index[1978] = '{3};
test_input[15832:15839] = '{32'hc20172b9, 32'h4243400b, 32'h404dab0c, 32'hc2c1e1a3, 32'hc15dad29, 32'h4291d05b, 32'hc21db5a5, 32'hc1956f69};
test_output[1979] = '{32'h4291d05b};
test_index[1979] = '{5};
test_input[15840:15847] = '{32'h41c82871, 32'h42205027, 32'h425e0174, 32'h42b96d86, 32'h4209439b, 32'hc1b83a39, 32'h42203dbe, 32'hc12142a5};
test_output[1980] = '{32'h42b96d86};
test_index[1980] = '{3};
test_input[15848:15855] = '{32'hc16844b2, 32'hc24061d5, 32'h42aec899, 32'h419cab52, 32'h42802171, 32'hc02d4243, 32'hc21c6108, 32'h4164ab90};
test_output[1981] = '{32'h42aec899};
test_index[1981] = '{2};
test_input[15856:15863] = '{32'hc2447f5d, 32'h4200b7d1, 32'hc1bd8cb6, 32'h42c72a9c, 32'h41721432, 32'h42338705, 32'hc2bad24b, 32'h427446b3};
test_output[1982] = '{32'h42c72a9c};
test_index[1982] = '{3};
test_input[15864:15871] = '{32'hc1e93061, 32'h4168b57d, 32'h40c0c452, 32'h42ba7683, 32'h42b03d3a, 32'h42785d16, 32'h429dcdfe, 32'h41207f10};
test_output[1983] = '{32'h42ba7683};
test_index[1983] = '{3};
test_input[15872:15879] = '{32'hc2ad2e92, 32'h41cc5242, 32'h4286a177, 32'hc289a052, 32'hc2b3371c, 32'h42a89f50, 32'h42c7d218, 32'hc1897981};
test_output[1984] = '{32'h42c7d218};
test_index[1984] = '{6};
test_input[15880:15887] = '{32'h42aa90fb, 32'hc26e6e52, 32'hc1b09251, 32'h420307bb, 32'hc2b380de, 32'h4134ac8f, 32'hc2a4cdd0, 32'h423f1f6e};
test_output[1985] = '{32'h42aa90fb};
test_index[1985] = '{0};
test_input[15888:15895] = '{32'hc252d052, 32'h42211487, 32'hc2b0a9ef, 32'h426458f1, 32'h42aa6510, 32'hc2250dea, 32'hc20c8106, 32'hc2a071af};
test_output[1986] = '{32'h42aa6510};
test_index[1986] = '{4};
test_input[15896:15903] = '{32'h42255bf4, 32'hc20160d4, 32'h42804826, 32'hbf64bf01, 32'hc2c73f97, 32'hc10d09b2, 32'hc2b65b09, 32'hc284e5d5};
test_output[1987] = '{32'h42804826};
test_index[1987] = '{2};
test_input[15904:15911] = '{32'hc25e70d8, 32'h42bcdd5e, 32'hc290cc6b, 32'h4274edfe, 32'h42772d9d, 32'hc24b2cbe, 32'hc2401117, 32'h423591e4};
test_output[1988] = '{32'h42bcdd5e};
test_index[1988] = '{1};
test_input[15912:15919] = '{32'hc18625dd, 32'h425eb2f1, 32'hc2c24f81, 32'h4216f8b3, 32'hc19f58bc, 32'h408d720d, 32'h422306d4, 32'hc29c4817};
test_output[1989] = '{32'h425eb2f1};
test_index[1989] = '{1};
test_input[15920:15927] = '{32'hc2b0ad65, 32'hc270e95b, 32'h42886989, 32'h41fcf9ad, 32'hc0d9dc1f, 32'h41bd4726, 32'h422ca31a, 32'h4271e340};
test_output[1990] = '{32'h42886989};
test_index[1990] = '{2};
test_input[15928:15935] = '{32'h42458724, 32'h4125dbeb, 32'h41190ba2, 32'h41dc8484, 32'hc047d3a4, 32'hc2957e0d, 32'hc2493d53, 32'hc2a46420};
test_output[1991] = '{32'h42458724};
test_index[1991] = '{0};
test_input[15936:15943] = '{32'hc290e7b3, 32'h42ae0878, 32'h421eec29, 32'h42a3f430, 32'h428a44b7, 32'h422f75ea, 32'hc268f30e, 32'h42bc76ee};
test_output[1992] = '{32'h42bc76ee};
test_index[1992] = '{7};
test_input[15944:15951] = '{32'hc288b8e1, 32'hc1dd9ce5, 32'hc23a91e5, 32'h42055670, 32'h41c19385, 32'h4056d5d0, 32'hc20dda5c, 32'hc290259e};
test_output[1993] = '{32'h42055670};
test_index[1993] = '{3};
test_input[15952:15959] = '{32'hc0b07ca8, 32'h4151e9ef, 32'h42835921, 32'h42977003, 32'h429466b4, 32'hc209a0d2, 32'hc223e694, 32'hc21bfdd5};
test_output[1994] = '{32'h42977003};
test_index[1994] = '{3};
test_input[15960:15967] = '{32'h41799c08, 32'hc09eb5c7, 32'hc2a5bda6, 32'h42165ae9, 32'h3f7bdefd, 32'hc2b507f3, 32'h3eb94548, 32'h41e4a996};
test_output[1995] = '{32'h42165ae9};
test_index[1995] = '{3};
test_input[15968:15975] = '{32'h42b246e3, 32'hc28fae0f, 32'hc1a7cac1, 32'hc1f8d1fe, 32'hc2b53ccb, 32'h42b216a3, 32'h4295c78f, 32'h422cc5e8};
test_output[1996] = '{32'h42b246e3};
test_index[1996] = '{0};
test_input[15976:15983] = '{32'hc18f1c11, 32'h410c0e9c, 32'hc29a5848, 32'h428b98fb, 32'h427841ca, 32'h41de226f, 32'hc07f4311, 32'hc218d9de};
test_output[1997] = '{32'h428b98fb};
test_index[1997] = '{3};
test_input[15984:15991] = '{32'hc2511634, 32'h420221fb, 32'h42bdbf49, 32'hc157f406, 32'hc26f3cbf, 32'h41308f37, 32'h427186e4, 32'hc284c121};
test_output[1998] = '{32'h42bdbf49};
test_index[1998] = '{2};
test_input[15992:15999] = '{32'hc1cb74eb, 32'h411ef711, 32'h42b47c38, 32'hc1827eff, 32'h423c7df0, 32'hc240d601, 32'hc2b66f3b, 32'h42293064};
test_output[1999] = '{32'h42b47c38};
test_index[1999] = '{2};
test_input[16000:16007] = '{32'hc1a22ebf, 32'h418cf2b7, 32'h42a384d9, 32'hc298ab83, 32'hc292a286, 32'hc0ade0b7, 32'hc1c77804, 32'h421b6776};
test_output[2000] = '{32'h42a384d9};
test_index[2000] = '{2};
test_input[16008:16015] = '{32'h4275edbc, 32'hc2a858d6, 32'hc2c5269c, 32'h41a24681, 32'hc2a396ca, 32'hc1e3e8a4, 32'hc2836fd2, 32'hc07a855d};
test_output[2001] = '{32'h4275edbc};
test_index[2001] = '{0};
test_input[16016:16023] = '{32'h42abf26d, 32'hc2511887, 32'hc289e563, 32'hc1d7c922, 32'hc270b69b, 32'h42b60df1, 32'h4290005c, 32'hc2c2e9e0};
test_output[2002] = '{32'h42b60df1};
test_index[2002] = '{5};
test_input[16024:16031] = '{32'hc215cbd8, 32'hc170c95c, 32'hc252ce6e, 32'hc26629fd, 32'hc295cc5b, 32'h425e513e, 32'hc27ba28a, 32'h4251288d};
test_output[2003] = '{32'h425e513e};
test_index[2003] = '{5};
test_input[16032:16039] = '{32'h42bf381a, 32'hc2a6997d, 32'hc2c150b9, 32'hc2c4caa9, 32'hc2384584, 32'hc2a0c965, 32'hc23af1a0, 32'hc2975a89};
test_output[2004] = '{32'h42bf381a};
test_index[2004] = '{0};
test_input[16040:16047] = '{32'hc1f40a26, 32'h42ae09ad, 32'h4194ec23, 32'hc2073ac3, 32'hc2b5a6bf, 32'hc0fe89bf, 32'h41b02fb3, 32'hc2bffc93};
test_output[2005] = '{32'h42ae09ad};
test_index[2005] = '{1};
test_input[16048:16055] = '{32'hc2167cb5, 32'h42932122, 32'h42c6006a, 32'hc1f0350e, 32'h4223c2d7, 32'h4256bd5a, 32'h428c7500, 32'h418b4541};
test_output[2006] = '{32'h42c6006a};
test_index[2006] = '{2};
test_input[16056:16063] = '{32'hc1ac68f2, 32'hc1d9eefb, 32'h4288365e, 32'h41a35c13, 32'h4219e897, 32'h4248c4de, 32'hc18186c3, 32'h4290710a};
test_output[2007] = '{32'h4290710a};
test_index[2007] = '{7};
test_input[16064:16071] = '{32'hc16d0b3d, 32'h42822f4b, 32'h4212f6d1, 32'hc1b9d816, 32'h4116ad59, 32'h428e5b4d, 32'h4172c467, 32'h426ce2fd};
test_output[2008] = '{32'h428e5b4d};
test_index[2008] = '{5};
test_input[16072:16079] = '{32'hc2a3dfac, 32'h42630cef, 32'hbe8b1f3e, 32'h4112c5b4, 32'hc229e7eb, 32'hc258fe01, 32'hc2539cca, 32'hc19cdb62};
test_output[2009] = '{32'h42630cef};
test_index[2009] = '{1};
test_input[16080:16087] = '{32'hc2c52eb7, 32'hc28fa425, 32'hc22584e9, 32'h42368ad8, 32'h4260bbf9, 32'h425eec06, 32'hc2654137, 32'hc22db3e1};
test_output[2010] = '{32'h4260bbf9};
test_index[2010] = '{4};
test_input[16088:16095] = '{32'h42a8e613, 32'hc236ab51, 32'h41eaa27b, 32'h421e3023, 32'hc254a086, 32'hc1feaff8, 32'h4253f7d4, 32'hc2c3668f};
test_output[2011] = '{32'h42a8e613};
test_index[2011] = '{0};
test_input[16096:16103] = '{32'hc29d28b7, 32'hc263d2ce, 32'hc1886099, 32'hc1848af8, 32'hc0547b3f, 32'h4111b94f, 32'h40d425db, 32'hc11e6d6c};
test_output[2012] = '{32'h4111b94f};
test_index[2012] = '{5};
test_input[16104:16111] = '{32'hc28c23d3, 32'h42a49554, 32'h4238c039, 32'h42a22ec9, 32'hc1a1f743, 32'h4284feb9, 32'hc2009456, 32'h425db550};
test_output[2013] = '{32'h42a49554};
test_index[2013] = '{1};
test_input[16112:16119] = '{32'hc2720c21, 32'h425d2764, 32'h41c3715d, 32'hc2acfcd4, 32'h4161fb3a, 32'h4295176d, 32'hc2063b05, 32'hc2c40260};
test_output[2014] = '{32'h4295176d};
test_index[2014] = '{5};
test_input[16120:16127] = '{32'hc1553170, 32'h423f8f0a, 32'h4275ef6b, 32'hc29b5910, 32'h429c9595, 32'h41d9273f, 32'hc094184b, 32'hc21ef036};
test_output[2015] = '{32'h429c9595};
test_index[2015] = '{4};
test_input[16128:16135] = '{32'h40a34b19, 32'h41ac42b4, 32'hc27e417c, 32'hc1b62531, 32'hc28b23ce, 32'hc28d29d7, 32'hc267f2c6, 32'h42ab99b1};
test_output[2016] = '{32'h42ab99b1};
test_index[2016] = '{7};
test_input[16136:16143] = '{32'hc2395e75, 32'hc2bce37c, 32'h4211a5a3, 32'hc23ea53e, 32'hc2563015, 32'hc27c00a3, 32'h3fbc1ced, 32'h425e4e51};
test_output[2017] = '{32'h425e4e51};
test_index[2017] = '{7};
test_input[16144:16151] = '{32'h403709bc, 32'h428b607b, 32'hc23d1656, 32'h3ea0ae13, 32'h429cea72, 32'hc18c07a8, 32'h42913426, 32'h42253b34};
test_output[2018] = '{32'h429cea72};
test_index[2018] = '{4};
test_input[16152:16159] = '{32'h40539e11, 32'h42a03b3d, 32'h42ac35b8, 32'hc2137ec3, 32'hc255a2af, 32'hc117de7b, 32'h42b58181, 32'h42b99fb0};
test_output[2019] = '{32'h42b99fb0};
test_index[2019] = '{7};
test_input[16160:16167] = '{32'h420e9d63, 32'hc2932aff, 32'h40057852, 32'h429eee95, 32'h4236c835, 32'h421b3820, 32'h42c2bd28, 32'h424cacaf};
test_output[2020] = '{32'h42c2bd28};
test_index[2020] = '{6};
test_input[16168:16175] = '{32'hc2aef3cf, 32'hc26c9e8e, 32'hc226c92b, 32'h428ae927, 32'h41e552b6, 32'h42a27b31, 32'hc21e1510, 32'hc2abef6e};
test_output[2021] = '{32'h42a27b31};
test_index[2021] = '{5};
test_input[16176:16183] = '{32'hc2ae0cd3, 32'h41e8511b, 32'hc2ac8c80, 32'h40a01908, 32'h42486ce7, 32'hc1ac30e8, 32'h429becc0, 32'h42855c15};
test_output[2022] = '{32'h429becc0};
test_index[2022] = '{6};
test_input[16184:16191] = '{32'h4296aa2a, 32'hc1bae7cf, 32'hc2ade575, 32'h42b01770, 32'h42c7d94d, 32'hc1a311c8, 32'hc2ad0595, 32'h3fd1cac2};
test_output[2023] = '{32'h42c7d94d};
test_index[2023] = '{4};
test_input[16192:16199] = '{32'h42a76f28, 32'h421dbffa, 32'h42a91cdb, 32'h40edf38a, 32'hc09a54a6, 32'hbfd99e01, 32'h425677c1, 32'hc2b50d0c};
test_output[2024] = '{32'h42a91cdb};
test_index[2024] = '{2};
test_input[16200:16207] = '{32'h422f7ffa, 32'h42c2a9a4, 32'hc0cd8d24, 32'h414abb05, 32'h423297d2, 32'hc29786c3, 32'h409ca785, 32'h42814010};
test_output[2025] = '{32'h42c2a9a4};
test_index[2025] = '{1};
test_input[16208:16215] = '{32'hc26540c2, 32'hc0a07858, 32'h42098c13, 32'hc15ad55b, 32'hc28ee0b9, 32'h42ade246, 32'h421aa67d, 32'h42807a30};
test_output[2026] = '{32'h42ade246};
test_index[2026] = '{5};
test_input[16216:16223] = '{32'h42a1cf55, 32'hc271ef9c, 32'hc18eb806, 32'h4250d674, 32'hc1eabb0a, 32'hc252c875, 32'h42625fdb, 32'h41e790fd};
test_output[2027] = '{32'h42a1cf55};
test_index[2027] = '{0};
test_input[16224:16231] = '{32'h429c9059, 32'h428f12ae, 32'h4205f507, 32'h428e2c3e, 32'hc25d26ea, 32'hc20abbaa, 32'hc1d999f1, 32'h41f4e2fa};
test_output[2028] = '{32'h429c9059};
test_index[2028] = '{0};
test_input[16232:16239] = '{32'hc2b28752, 32'hc20ea6de, 32'hc236b9cd, 32'hc26bab0e, 32'h423c6121, 32'h429d9984, 32'hc2855b52, 32'h42afd473};
test_output[2029] = '{32'h42afd473};
test_index[2029] = '{7};
test_input[16240:16247] = '{32'hc2c48cdb, 32'hc232449a, 32'h421f26d3, 32'h42ba26e7, 32'hc22be909, 32'h426820a8, 32'hc2b9a739, 32'h421ca78d};
test_output[2030] = '{32'h42ba26e7};
test_index[2030] = '{3};
test_input[16248:16255] = '{32'h42b86c8d, 32'h41506ecd, 32'hc1759e6a, 32'h42996ae5, 32'h42950d05, 32'hc296a119, 32'h42549f75, 32'h422babce};
test_output[2031] = '{32'h42b86c8d};
test_index[2031] = '{0};
test_input[16256:16263] = '{32'h429537a2, 32'h42119743, 32'hc1bd6466, 32'h41b51eb7, 32'h42bb9313, 32'h421f98dd, 32'h40911242, 32'h414347a8};
test_output[2032] = '{32'h42bb9313};
test_index[2032] = '{4};
test_input[16264:16271] = '{32'hc2bee0fd, 32'hc2360b46, 32'h42af52ba, 32'h423bf5df, 32'h42a8de0a, 32'h42073716, 32'h4200e0f8, 32'hc0f736ee};
test_output[2033] = '{32'h42af52ba};
test_index[2033] = '{2};
test_input[16272:16279] = '{32'hc2af74d0, 32'h42b664a9, 32'hc2620ef4, 32'hc2a1c1bb, 32'h41fdbe3e, 32'h40ed7d14, 32'h42b05d2b, 32'h429968aa};
test_output[2034] = '{32'h42b664a9};
test_index[2034] = '{1};
test_input[16280:16287] = '{32'hc1354d01, 32'h426f54f6, 32'hc2767b4f, 32'h42901147, 32'h42b050d0, 32'h416f9325, 32'h42a77bfb, 32'hc1d94cb4};
test_output[2035] = '{32'h42b050d0};
test_index[2035] = '{4};
test_input[16288:16295] = '{32'h418f10dc, 32'hc1e8c42b, 32'h42a3d3c7, 32'h4290e695, 32'hc186b68e, 32'hc229deca, 32'hc18f6632, 32'h4215727b};
test_output[2036] = '{32'h42a3d3c7};
test_index[2036] = '{2};
test_input[16296:16303] = '{32'hc299c61f, 32'hc08c3a79, 32'hc2a01b9b, 32'h4237a49c, 32'hc20a1763, 32'h42be45a6, 32'hc270c309, 32'hc2abb550};
test_output[2037] = '{32'h42be45a6};
test_index[2037] = '{5};
test_input[16304:16311] = '{32'h428e250b, 32'hc2192817, 32'hc2a267e8, 32'h421e7111, 32'hc28738c3, 32'hbf9367ac, 32'h421ca067, 32'h41126ca4};
test_output[2038] = '{32'h428e250b};
test_index[2038] = '{0};
test_input[16312:16319] = '{32'h42b389bc, 32'h42b9a6f1, 32'h422ab358, 32'hc0a1ead4, 32'hc2884972, 32'h4257c683, 32'h4261003c, 32'hc24f2399};
test_output[2039] = '{32'h42b9a6f1};
test_index[2039] = '{1};
test_input[16320:16327] = '{32'h40f9ce1f, 32'h42178dce, 32'hc26b9692, 32'hc2c6a0bb, 32'hc208c231, 32'h4272e2e7, 32'hc2838994, 32'h4274e29b};
test_output[2040] = '{32'h4274e29b};
test_index[2040] = '{7};
test_input[16328:16335] = '{32'h42c643e5, 32'h41a39ca8, 32'h4133f61f, 32'h429decc7, 32'hc27c79c7, 32'h4177a093, 32'h4185921d, 32'hc2849473};
test_output[2041] = '{32'h42c643e5};
test_index[2041] = '{0};
test_input[16336:16343] = '{32'hc29ed846, 32'hc1d41b0c, 32'h41edb80f, 32'hc2c1809d, 32'h40a619d9, 32'h42aea9cc, 32'h42a7c67a, 32'h428bb381};
test_output[2042] = '{32'h42aea9cc};
test_index[2042] = '{5};
test_input[16344:16351] = '{32'h4287126a, 32'h41df390e, 32'hc1eb3aff, 32'hc2afcb5e, 32'h426e3e5f, 32'hc28de718, 32'hc252c38c, 32'hc1d64afb};
test_output[2043] = '{32'h4287126a};
test_index[2043] = '{0};
test_input[16352:16359] = '{32'h4211df10, 32'hc1be06cd, 32'hc0bb65d5, 32'hc09709d2, 32'hbf92337a, 32'h41d63155, 32'hc12d1026, 32'h41dd23c1};
test_output[2044] = '{32'h4211df10};
test_index[2044] = '{0};
test_input[16360:16367] = '{32'hc2ad86b2, 32'h4167be8e, 32'hc18c670f, 32'h42bb6b24, 32'hc291acce, 32'h42b2154e, 32'h42b83ce7, 32'hc1b1f0eb};
test_output[2045] = '{32'h42bb6b24};
test_index[2045] = '{3};
test_input[16368:16375] = '{32'hc0ae1860, 32'hc1c0fed8, 32'hc28c1b7f, 32'h42a21b4e, 32'h42000173, 32'hc1782293, 32'hbf361cc8, 32'h4289b19d};
test_output[2046] = '{32'h42a21b4e};
test_index[2046] = '{3};
test_input[16376:16383] = '{32'hc2a2f1b3, 32'h41d2384f, 32'h42aceef2, 32'h41e6f734, 32'hc2b9db72, 32'hc209010d, 32'hc28c7ae3, 32'hc22329d9};
test_output[2047] = '{32'h42aceef2};
test_index[2047] = '{2};
test_input[16384:16391] = '{32'hc2bc4c45, 32'h416dfa10, 32'hc2af339b, 32'h4296ca9c, 32'h42535c67, 32'h42bd8c97, 32'h4223e75f, 32'hc2b24fea};
test_output[2048] = '{32'h42bd8c97};
test_index[2048] = '{5};
test_input[16392:16399] = '{32'h41a97aee, 32'h42b54b90, 32'hc187206b, 32'hc287e062, 32'hc2a484d0, 32'h400e32a1, 32'h425df419, 32'h418f4d2e};
test_output[2049] = '{32'h42b54b90};
test_index[2049] = '{1};
test_input[16400:16407] = '{32'hc12c6022, 32'h4298b008, 32'hc2316529, 32'h4237de11, 32'h423e75d8, 32'h42c4c44e, 32'h42b6541f, 32'hc2a0a1b3};
test_output[2050] = '{32'h42c4c44e};
test_index[2050] = '{5};
test_input[16408:16415] = '{32'hc15589c4, 32'h42a2c07d, 32'hc2b8023e, 32'hc1a99079, 32'hc1d500a7, 32'hc2674d9b, 32'h42305004, 32'hc2936f47};
test_output[2051] = '{32'h42a2c07d};
test_index[2051] = '{1};
test_input[16416:16423] = '{32'hc227824e, 32'hc2728de5, 32'h4243f95a, 32'h42ba42b6, 32'h428ad292, 32'h41ed7565, 32'h4049b863, 32'hc2a8abe1};
test_output[2052] = '{32'h42ba42b6};
test_index[2052] = '{3};
test_input[16424:16431] = '{32'h418b9f86, 32'h426f1bf9, 32'h42a87ba8, 32'h426d4f46, 32'h41d6c62e, 32'hc11f662a, 32'hc2b376b4, 32'hc231f3cd};
test_output[2053] = '{32'h42a87ba8};
test_index[2053] = '{2};
test_input[16432:16439] = '{32'hc01fc1f0, 32'h41f7a542, 32'hc1f9780d, 32'hc22d14e5, 32'hc173ab17, 32'h422a9ac0, 32'h420d91fb, 32'h42692c61};
test_output[2054] = '{32'h42692c61};
test_index[2054] = '{7};
test_input[16440:16447] = '{32'hc23632e7, 32'h4180f004, 32'hc2b0d27c, 32'h4229190b, 32'h42a99710, 32'h420471f7, 32'h42bae58a, 32'h41ccee17};
test_output[2055] = '{32'h42bae58a};
test_index[2055] = '{6};
test_input[16448:16455] = '{32'hc24138e0, 32'hc18bed29, 32'hc1152c68, 32'hc272b695, 32'hc1b2684b, 32'hc240a0b5, 32'hc2baa2b0, 32'hc112d330};
test_output[2056] = '{32'hc112d330};
test_index[2056] = '{7};
test_input[16456:16463] = '{32'h4266b887, 32'h42559ab6, 32'hc2c5f8fa, 32'hc2b88187, 32'hc2c49248, 32'hc1d73a23, 32'hc1ff6022, 32'hc1b69967};
test_output[2057] = '{32'h4266b887};
test_index[2057] = '{0};
test_input[16464:16471] = '{32'hc2b2298a, 32'h42b8f08b, 32'h41ad06f8, 32'h3fbf7991, 32'hc2b96d09, 32'h42c032d9, 32'h421a378e, 32'h41d5e6ef};
test_output[2058] = '{32'h42c032d9};
test_index[2058] = '{5};
test_input[16472:16479] = '{32'hc2c64238, 32'h420a9bc5, 32'hc1841a5f, 32'hc230df7b, 32'hc295187d, 32'h426cb211, 32'h402febd3, 32'hc185fe48};
test_output[2059] = '{32'h426cb211};
test_index[2059] = '{5};
test_input[16480:16487] = '{32'hc2239c4a, 32'hc2abe903, 32'hc29fe084, 32'hbf1fdd57, 32'hc2a3c4f0, 32'h42251d0a, 32'h42bb3346, 32'h4294b40a};
test_output[2060] = '{32'h42bb3346};
test_index[2060] = '{6};
test_input[16488:16495] = '{32'h426e4a6c, 32'h426333e5, 32'hc255e384, 32'h428dee08, 32'h4283f966, 32'hc24f6e72, 32'h42130c1d, 32'hc294ed8f};
test_output[2061] = '{32'h428dee08};
test_index[2061] = '{3};
test_input[16496:16503] = '{32'h415c69c2, 32'hc20afff2, 32'hc162e648, 32'hc19e37ce, 32'hc2c05efa, 32'h42ac2333, 32'h42a80d16, 32'h426da945};
test_output[2062] = '{32'h42ac2333};
test_index[2062] = '{5};
test_input[16504:16511] = '{32'hc253a321, 32'hc22d9da8, 32'h42931e66, 32'hc1c2c9c2, 32'h425b2ef1, 32'h423f4929, 32'hc293e082, 32'h421688c4};
test_output[2063] = '{32'h42931e66};
test_index[2063] = '{2};
test_input[16512:16519] = '{32'h426f25e8, 32'hbea9dbb6, 32'hc1a30d44, 32'hc288dbbf, 32'hc2393f53, 32'h4218ec81, 32'h428b04e5, 32'h422dcc74};
test_output[2064] = '{32'h428b04e5};
test_index[2064] = '{6};
test_input[16520:16527] = '{32'hc2ad5263, 32'hc2c33510, 32'h4280ac34, 32'hc2c7ca25, 32'h41ccbca8, 32'h41bbbf5d, 32'h42a79366, 32'hc2bb7d09};
test_output[2065] = '{32'h42a79366};
test_index[2065] = '{6};
test_input[16528:16535] = '{32'h4288bd3e, 32'h4207ccba, 32'hc2060d7f, 32'hc25ea9b6, 32'hc20ab5dd, 32'h4297e1f4, 32'h42a982a1, 32'hc235caaf};
test_output[2066] = '{32'h42a982a1};
test_index[2066] = '{6};
test_input[16536:16543] = '{32'h4223e4e9, 32'hc101c088, 32'hc283cb6f, 32'hbfacc4cf, 32'hc29dc619, 32'h424d991c, 32'h41d79c25, 32'h42838df6};
test_output[2067] = '{32'h42838df6};
test_index[2067] = '{7};
test_input[16544:16551] = '{32'h42bf7d63, 32'h429b74be, 32'hc26ed94a, 32'h421c13bc, 32'hc255181a, 32'h4285682b, 32'hc23bba66, 32'hc2c11c55};
test_output[2068] = '{32'h42bf7d63};
test_index[2068] = '{0};
test_input[16552:16559] = '{32'h42b89c9c, 32'hc11f1543, 32'hc2804c83, 32'h427c13df, 32'hc215e72e, 32'h41f18463, 32'hc2b9d9f8, 32'hc29f4a64};
test_output[2069] = '{32'h42b89c9c};
test_index[2069] = '{0};
test_input[16560:16567] = '{32'h42aab803, 32'hc2c604d3, 32'hc1aed890, 32'h42a87faf, 32'h41989603, 32'hc2957a18, 32'hc1b170ba, 32'h428b765a};
test_output[2070] = '{32'h42aab803};
test_index[2070] = '{0};
test_input[16568:16575] = '{32'hc2957ea1, 32'hbfac2d10, 32'h429364b3, 32'hc25beb64, 32'h428fc0e6, 32'hc2ba5fbc, 32'hc25ef98a, 32'h41b66954};
test_output[2071] = '{32'h429364b3};
test_index[2071] = '{2};
test_input[16576:16583] = '{32'h42a5f980, 32'hc27c984a, 32'hc23cda56, 32'hc282fadd, 32'h4229e8c7, 32'hc2336036, 32'hc289ff9f, 32'hc294a9d0};
test_output[2072] = '{32'h42a5f980};
test_index[2072] = '{0};
test_input[16584:16591] = '{32'h420eb7d8, 32'hc24bf736, 32'hc09f2ba4, 32'h42a4a9fb, 32'hc2952f9a, 32'hc23acbaa, 32'h42a9b146, 32'hc1234242};
test_output[2073] = '{32'h42a9b146};
test_index[2073] = '{6};
test_input[16592:16599] = '{32'hc290d532, 32'h4270554b, 32'h40e3c792, 32'h42c7d118, 32'hc2988d95, 32'h423de70e, 32'hc128812f, 32'h41b31087};
test_output[2074] = '{32'h42c7d118};
test_index[2074] = '{3};
test_input[16600:16607] = '{32'hc2c07a55, 32'hc2b45c09, 32'hc23f9da9, 32'hc18ab2c3, 32'hc10b6ce0, 32'hc2088ffe, 32'h428c7855, 32'hc289a616};
test_output[2075] = '{32'h428c7855};
test_index[2075] = '{6};
test_input[16608:16615] = '{32'hc256adad, 32'h424b327f, 32'hc27d33b8, 32'h4099fb06, 32'hc291394e, 32'h428b2ed6, 32'hc1c5c017, 32'h42c1b47e};
test_output[2076] = '{32'h42c1b47e};
test_index[2076] = '{7};
test_input[16616:16623] = '{32'hc1ac204f, 32'hc113b567, 32'h4250c4b9, 32'hc1848955, 32'h42c40f6c, 32'hc2bb6957, 32'h423bbe5f, 32'h41175bcd};
test_output[2077] = '{32'h42c40f6c};
test_index[2077] = '{4};
test_input[16624:16631] = '{32'h4189260c, 32'hc18aec49, 32'h41e1e2e0, 32'h41c9999f, 32'h425e4fcd, 32'h4213ec11, 32'hc2c6800c, 32'h409cc420};
test_output[2078] = '{32'h425e4fcd};
test_index[2078] = '{4};
test_input[16632:16639] = '{32'hc20a00f6, 32'hc27fce17, 32'h41b69562, 32'h4258cae7, 32'h41376e8f, 32'h407788e5, 32'hc28c062c, 32'h4230d530};
test_output[2079] = '{32'h4258cae7};
test_index[2079] = '{3};
test_input[16640:16647] = '{32'hc2b48f41, 32'hc16c74a9, 32'hc2c3b12d, 32'hc2371580, 32'hc2842dce, 32'h413fddf9, 32'hc225860a, 32'h4201f036};
test_output[2080] = '{32'h4201f036};
test_index[2080] = '{7};
test_input[16648:16655] = '{32'h42c72838, 32'hc2be7671, 32'h418d6759, 32'h42286c3b, 32'hc2212220, 32'hc2bc2e3e, 32'h412b6564, 32'hc11245f4};
test_output[2081] = '{32'h42c72838};
test_index[2081] = '{0};
test_input[16656:16663] = '{32'hc11f9d6c, 32'hc286f4e5, 32'h42293b44, 32'h42424ba2, 32'h42475d2c, 32'hc2be8ae8, 32'hc2243803, 32'hc2010bfd};
test_output[2082] = '{32'h42475d2c};
test_index[2082] = '{4};
test_input[16664:16671] = '{32'h42a004c1, 32'h4287bc31, 32'h4024c8ca, 32'h41f2d1dc, 32'h4224ba20, 32'h42b873be, 32'hc26a16bf, 32'hc2498d55};
test_output[2083] = '{32'h42b873be};
test_index[2083] = '{5};
test_input[16672:16679] = '{32'hc2c7de8f, 32'hc22483b1, 32'hc1a6ea78, 32'h425d7449, 32'hc2620adc, 32'h42123056, 32'h42bd25af, 32'h417daffb};
test_output[2084] = '{32'h42bd25af};
test_index[2084] = '{6};
test_input[16680:16687] = '{32'hc1039499, 32'h42694f81, 32'hbf8100b2, 32'h42ab534a, 32'h4282a067, 32'hc2c7ad69, 32'h42997c04, 32'h41ee6455};
test_output[2085] = '{32'h42ab534a};
test_index[2085] = '{3};
test_input[16688:16695] = '{32'hc22d79e3, 32'h410a11b8, 32'h428d4e92, 32'h42848084, 32'h420eae31, 32'hc1a39f98, 32'h4275423c, 32'hc29a3205};
test_output[2086] = '{32'h428d4e92};
test_index[2086] = '{2};
test_input[16696:16703] = '{32'hc20f7e08, 32'h420f9e81, 32'h4298b8e5, 32'hc2c1d3e6, 32'h42a550fa, 32'h4235bab1, 32'hc135fb46, 32'hc2a04f10};
test_output[2087] = '{32'h42a550fa};
test_index[2087] = '{4};
test_input[16704:16711] = '{32'hc292599f, 32'hc28b34df, 32'hc251039c, 32'h42ad7496, 32'h42bc55f7, 32'hc1adf346, 32'hc2ac6f4d, 32'h41bdabe2};
test_output[2088] = '{32'h42bc55f7};
test_index[2088] = '{4};
test_input[16712:16719] = '{32'h428ea0ce, 32'hc2483ab6, 32'hc2812020, 32'hc25fd70e, 32'h40a6f051, 32'h42b17fda, 32'h425ff61d, 32'h413570f7};
test_output[2089] = '{32'h42b17fda};
test_index[2089] = '{5};
test_input[16720:16727] = '{32'hc19ab74a, 32'h413492b8, 32'h3ee7d23a, 32'h42449242, 32'hc1c61788, 32'hc2babfbf, 32'h429fe8cd, 32'h4158ba04};
test_output[2090] = '{32'h429fe8cd};
test_index[2090] = '{6};
test_input[16728:16735] = '{32'h42c181ac, 32'h425690f2, 32'hc164b828, 32'h42c49eb7, 32'hc18680b5, 32'h41e5af2e, 32'h42912853, 32'h4089314e};
test_output[2091] = '{32'h42c49eb7};
test_index[2091] = '{3};
test_input[16736:16743] = '{32'hc226e938, 32'hc295aa08, 32'hc29a921f, 32'hc2098fe8, 32'h422a16ae, 32'h4271a8ce, 32'hc2aa6789, 32'hc2ba5ab4};
test_output[2092] = '{32'h4271a8ce};
test_index[2092] = '{5};
test_input[16744:16751] = '{32'hc25e8cfb, 32'hc037dddf, 32'hc209245c, 32'hc07077cf, 32'hc21462a2, 32'hc0d67b13, 32'hc2b613f4, 32'hc1145a2f};
test_output[2093] = '{32'hc037dddf};
test_index[2093] = '{1};
test_input[16752:16759] = '{32'h42a07cd7, 32'h410eb6bc, 32'hc02b6f8d, 32'h42aa65e1, 32'h4229ca6c, 32'hc178d902, 32'h42931a44, 32'h41c21c5c};
test_output[2094] = '{32'h42aa65e1};
test_index[2094] = '{3};
test_input[16760:16767] = '{32'hc2324aeb, 32'h41f5154b, 32'h42046e3a, 32'hc2b64626, 32'h414640e7, 32'hc2c79f41, 32'hc28dd380, 32'h4297e392};
test_output[2095] = '{32'h4297e392};
test_index[2095] = '{7};
test_input[16768:16775] = '{32'h3fe6728b, 32'h42b6b9d2, 32'h42858543, 32'h425f81be, 32'h4217c055, 32'h428da85c, 32'h4185f715, 32'hc1f61297};
test_output[2096] = '{32'h42b6b9d2};
test_index[2096] = '{1};
test_input[16776:16783] = '{32'h4095f1ce, 32'h42a37ec8, 32'h42652616, 32'h4298a9f0, 32'h408c9804, 32'h413ce51a, 32'h4295de25, 32'hc22ee40b};
test_output[2097] = '{32'h42a37ec8};
test_index[2097] = '{1};
test_input[16784:16791] = '{32'h42a6047b, 32'hc2668e49, 32'h42a09410, 32'hc2433c42, 32'hc2405ef4, 32'h42b7b58c, 32'h42937406, 32'h42a0776a};
test_output[2098] = '{32'h42b7b58c};
test_index[2098] = '{5};
test_input[16792:16799] = '{32'hc0aa1329, 32'hc2c071be, 32'hc2a70c19, 32'h42901761, 32'hc2853c76, 32'hc202507e, 32'h40a4cd93, 32'h41d84eef};
test_output[2099] = '{32'h42901761};
test_index[2099] = '{3};
test_input[16800:16807] = '{32'h42394fc9, 32'hc0b506a1, 32'h429e5860, 32'h42c0292c, 32'hc2671ba1, 32'hc1aee07f, 32'hc2bd8136, 32'hc29ae995};
test_output[2100] = '{32'h42c0292c};
test_index[2100] = '{3};
test_input[16808:16815] = '{32'hc2615bf4, 32'h41ef11ce, 32'h426664f9, 32'hc2b6e3d0, 32'hc2b3a944, 32'hc1e99765, 32'h42abc0e1, 32'hc2601fc7};
test_output[2101] = '{32'h42abc0e1};
test_index[2101] = '{6};
test_input[16816:16823] = '{32'h42685450, 32'hc1438827, 32'h4293bf6a, 32'h42916137, 32'hc20e73a9, 32'h424bf68a, 32'h41d9c857, 32'hc2c386a1};
test_output[2102] = '{32'h4293bf6a};
test_index[2102] = '{2};
test_input[16824:16831] = '{32'h421cb056, 32'hc20284f4, 32'h421e1c25, 32'hc2b92c73, 32'hc21ea4f6, 32'hc2a56b7d, 32'hc236243b, 32'hc1252c96};
test_output[2103] = '{32'h421e1c25};
test_index[2103] = '{2};
test_input[16832:16839] = '{32'hc0ba4290, 32'hc1e8dc77, 32'h41b3b76d, 32'hc1bff52d, 32'h42416f81, 32'h4204ff64, 32'h42a8f003, 32'hc2b65b3c};
test_output[2104] = '{32'h42a8f003};
test_index[2104] = '{6};
test_input[16840:16847] = '{32'hc117a3ad, 32'hc1c6491c, 32'hc2b98ce5, 32'hc1abe086, 32'hc2422466, 32'h42292968, 32'hc16f491c, 32'h4202e66b};
test_output[2105] = '{32'h42292968};
test_index[2105] = '{5};
test_input[16848:16855] = '{32'hc26b53ad, 32'h42c1d0fc, 32'hc28a3087, 32'hc19a85d3, 32'hc24e1f27, 32'h427d275c, 32'h424a2e85, 32'h420452d8};
test_output[2106] = '{32'h42c1d0fc};
test_index[2106] = '{1};
test_input[16856:16863] = '{32'hc19096fa, 32'h428c7339, 32'h420ccb09, 32'hc20bb4e2, 32'hc2658b51, 32'hc2bcb611, 32'hc18d8332, 32'hc24d603c};
test_output[2107] = '{32'h428c7339};
test_index[2107] = '{1};
test_input[16864:16871] = '{32'hc284cd7a, 32'h4184be63, 32'h42c0a6b5, 32'hc29a1e23, 32'h420063d0, 32'h42628df7, 32'h420227f6, 32'h42a6be97};
test_output[2108] = '{32'h42c0a6b5};
test_index[2108] = '{2};
test_input[16872:16879] = '{32'hc2179b47, 32'hc29f1138, 32'h4298e874, 32'h42bca85e, 32'h42be4f43, 32'h42931966, 32'h42341947, 32'hc1ae8487};
test_output[2109] = '{32'h42be4f43};
test_index[2109] = '{4};
test_input[16880:16887] = '{32'h415b2fa7, 32'hc2b2a632, 32'h4296a107, 32'hc1ee829d, 32'hc27bb030, 32'h4190036e, 32'hc23fe0cd, 32'hc0279c1c};
test_output[2110] = '{32'h4296a107};
test_index[2110] = '{2};
test_input[16888:16895] = '{32'h4099c10b, 32'h428ce3e5, 32'hc23e3a44, 32'hc2b87e6e, 32'hc26bdeb2, 32'hc23d2db5, 32'hc1631a46, 32'h42705313};
test_output[2111] = '{32'h428ce3e5};
test_index[2111] = '{1};
test_input[16896:16903] = '{32'hc218ffea, 32'h4221cfb6, 32'hc1e7adf1, 32'h423844af, 32'h42aa0c50, 32'hc295acbc, 32'h42714ef7, 32'hc282a109};
test_output[2112] = '{32'h42aa0c50};
test_index[2112] = '{4};
test_input[16904:16911] = '{32'hc2b07e1e, 32'h428b9637, 32'h42314861, 32'h42453984, 32'h428d7835, 32'h4064df7c, 32'hc28687aa, 32'h41f36501};
test_output[2113] = '{32'h428d7835};
test_index[2113] = '{4};
test_input[16912:16919] = '{32'hc1a82d83, 32'hc26a42f9, 32'hc28c5a0c, 32'hc2310680, 32'hc2a4482e, 32'hc06f6f9d, 32'hc2437ef1, 32'h42925a7c};
test_output[2114] = '{32'h42925a7c};
test_index[2114] = '{7};
test_input[16920:16927] = '{32'hc289db1d, 32'h423d071a, 32'hc21a3b9a, 32'h42a23a36, 32'h40072bc6, 32'h42671b0e, 32'hc2b24b48, 32'hc27e92b0};
test_output[2115] = '{32'h42a23a36};
test_index[2115] = '{3};
test_input[16928:16935] = '{32'hc1cea62a, 32'h41efd487, 32'h4192eb6b, 32'hc245a481, 32'hc1fc9c23, 32'h424bdeb8, 32'hc26eaeb7, 32'h42abd830};
test_output[2116] = '{32'h42abd830};
test_index[2116] = '{7};
test_input[16936:16943] = '{32'hc25e352d, 32'h42a053d4, 32'hc1964d49, 32'h42641e09, 32'h422cf1a1, 32'h427b9475, 32'h424af32d, 32'h42846d62};
test_output[2117] = '{32'h42a053d4};
test_index[2117] = '{1};
test_input[16944:16951] = '{32'h42b4ae10, 32'hc24f53f3, 32'h4197d235, 32'h428c506f, 32'h41f80220, 32'h422fbdae, 32'h42108ba4, 32'h42a8f252};
test_output[2118] = '{32'h42b4ae10};
test_index[2118] = '{0};
test_input[16952:16959] = '{32'h4240d07b, 32'hc0531212, 32'hc2aa4ea2, 32'hc1ce3da5, 32'hc2a29986, 32'h428ccf25, 32'h4191f1ef, 32'h42c4011d};
test_output[2119] = '{32'h42c4011d};
test_index[2119] = '{7};
test_input[16960:16967] = '{32'hc1cc8aad, 32'hbfda278e, 32'h42925533, 32'h4184f97e, 32'h42790de0, 32'hc25466a5, 32'hc2840191, 32'h41aee9c7};
test_output[2120] = '{32'h42925533};
test_index[2120] = '{2};
test_input[16968:16975] = '{32'h42ace795, 32'hc276f298, 32'hc20f9af7, 32'h42bbb70a, 32'hbf0e43ad, 32'hc28c2b0c, 32'h41ade3fd, 32'hc2bee2d2};
test_output[2121] = '{32'h42bbb70a};
test_index[2121] = '{3};
test_input[16976:16983] = '{32'h423ff1f0, 32'hc23f10f8, 32'hc173ae5e, 32'hc0af6fd2, 32'hc2b992c0, 32'hc2b333b5, 32'h424595c6, 32'h42ace1fe};
test_output[2122] = '{32'h42ace1fe};
test_index[2122] = '{7};
test_input[16984:16991] = '{32'h41fe9d3d, 32'hc274683b, 32'hc219b2da, 32'h42c4da89, 32'hc2a62c5f, 32'h3fa3adeb, 32'h42ab5c3a, 32'hc20b9ecb};
test_output[2123] = '{32'h42c4da89};
test_index[2123] = '{3};
test_input[16992:16999] = '{32'h420c1706, 32'hc26f6839, 32'h423969fb, 32'hc00979db, 32'hc09a28b1, 32'h427ffe5f, 32'hc2a78034, 32'h4205dd80};
test_output[2124] = '{32'h427ffe5f};
test_index[2124] = '{5};
test_input[17000:17007] = '{32'h42b9bfa7, 32'hc2c653d0, 32'hc1d0b1e7, 32'hc2962db2, 32'hc24d0fe6, 32'h42c35181, 32'hc22189fe, 32'h41c88287};
test_output[2125] = '{32'h42c35181};
test_index[2125] = '{5};
test_input[17008:17015] = '{32'hc2a75edd, 32'hc2491c43, 32'hc28ec010, 32'h42b3d7c2, 32'hc09cd08c, 32'hc29136a8, 32'h421e5602, 32'h42a3e86e};
test_output[2126] = '{32'h42b3d7c2};
test_index[2126] = '{3};
test_input[17016:17023] = '{32'hc28fe44b, 32'h42636378, 32'hc1010026, 32'h42a6bf89, 32'hc0b70960, 32'hc180c7d7, 32'h4297a520, 32'hc17c97e5};
test_output[2127] = '{32'h42a6bf89};
test_index[2127] = '{3};
test_input[17024:17031] = '{32'hc284569d, 32'h41a9e3cd, 32'h429a2656, 32'hc0c4e118, 32'hc15cb62c, 32'h4201f959, 32'h419489f4, 32'hc1913d18};
test_output[2128] = '{32'h429a2656};
test_index[2128] = '{2};
test_input[17032:17039] = '{32'h4197aa89, 32'hc24db497, 32'h4187d3da, 32'hc22ec5f6, 32'h423ae524, 32'hc235c685, 32'h42c20a77, 32'h41a5f937};
test_output[2129] = '{32'h42c20a77};
test_index[2129] = '{6};
test_input[17040:17047] = '{32'h42a1566a, 32'h425c5fca, 32'h42660ee2, 32'hc2a0280f, 32'hc2279f8b, 32'h42226b42, 32'hc2b75696, 32'hc29f7414};
test_output[2130] = '{32'h42a1566a};
test_index[2130] = '{0};
test_input[17048:17055] = '{32'hc285cf1a, 32'hc1a09f4f, 32'hc29bd27f, 32'hc2bc8b81, 32'hc1725047, 32'hc1ca25f8, 32'h41ffedde, 32'h4190366b};
test_output[2131] = '{32'h41ffedde};
test_index[2131] = '{6};
test_input[17056:17063] = '{32'h425dc0f3, 32'h41a85a4f, 32'hc28feb29, 32'h42b8a13c, 32'h42a04ba8, 32'h41f7a954, 32'hc2c0e2e1, 32'h41e4950f};
test_output[2132] = '{32'h42b8a13c};
test_index[2132] = '{3};
test_input[17064:17071] = '{32'h415c42d2, 32'h429fd83d, 32'hc2bbdeb6, 32'hc297c89d, 32'h42ba0baf, 32'h420de077, 32'hc2b5781b, 32'hc201c199};
test_output[2133] = '{32'h42ba0baf};
test_index[2133] = '{4};
test_input[17072:17079] = '{32'h4294a845, 32'hc1f2c586, 32'h41df83e5, 32'hc1978f79, 32'hc156020d, 32'h41c0d2ff, 32'hc2bd4425, 32'hc1b659d5};
test_output[2134] = '{32'h4294a845};
test_index[2134] = '{0};
test_input[17080:17087] = '{32'h402a124a, 32'hc1e32f51, 32'hc2797398, 32'hc1ba834d, 32'h412c0003, 32'hc2a4b964, 32'hc10b7947, 32'h41c31f53};
test_output[2135] = '{32'h41c31f53};
test_index[2135] = '{7};
test_input[17088:17095] = '{32'hc1c40d3f, 32'hc2a68a83, 32'hc27e9240, 32'hc23ffd67, 32'h4265447a, 32'h422ea851, 32'hc2c4b2fb, 32'h4096ebf1};
test_output[2136] = '{32'h4265447a};
test_index[2136] = '{4};
test_input[17096:17103] = '{32'hc2aa5552, 32'hc2a681ae, 32'hc11ef9cf, 32'h41b18566, 32'h42a65121, 32'h42337cbf, 32'hc2bd125e, 32'h41bc9b52};
test_output[2137] = '{32'h42a65121};
test_index[2137] = '{4};
test_input[17104:17111] = '{32'hc1a06c59, 32'h42534462, 32'hc1e09a4f, 32'h42058cb5, 32'h422bfce3, 32'hc29873a2, 32'h42bb57eb, 32'h42b0c6e5};
test_output[2138] = '{32'h42bb57eb};
test_index[2138] = '{6};
test_input[17112:17119] = '{32'h418d6d56, 32'hc1812111, 32'h4216bddb, 32'h423897c1, 32'h40fc88a7, 32'h42a38bd4, 32'h426e26cc, 32'hc19b5ff3};
test_output[2139] = '{32'h42a38bd4};
test_index[2139] = '{5};
test_input[17120:17127] = '{32'h429e509c, 32'hc2170c30, 32'h4196b969, 32'hc09e4d4d, 32'h42877c1c, 32'hc261fe26, 32'h41428828, 32'h420e6074};
test_output[2140] = '{32'h429e509c};
test_index[2140] = '{0};
test_input[17128:17135] = '{32'h41bf9347, 32'h425ebae1, 32'hc1d4db09, 32'h42ab565f, 32'h4204f615, 32'h4209a3ec, 32'h42c63e84, 32'hc2c55492};
test_output[2141] = '{32'h42c63e84};
test_index[2141] = '{6};
test_input[17136:17143] = '{32'h42b7756a, 32'h42451348, 32'h42777cf1, 32'hc1294ec8, 32'hc28d1c61, 32'hc2224633, 32'hc2000e50, 32'h41b586aa};
test_output[2142] = '{32'h42b7756a};
test_index[2142] = '{0};
test_input[17144:17151] = '{32'hc2a4944d, 32'hc2b6e9ae, 32'h411cdc9b, 32'hc11fcb0c, 32'hc2622741, 32'h42652989, 32'hc26317c7, 32'hc270c4bd};
test_output[2143] = '{32'h42652989};
test_index[2143] = '{5};
test_input[17152:17159] = '{32'hc27e1a55, 32'hc29bf53d, 32'h42ac616f, 32'h40a591aa, 32'hc27ad2c0, 32'hc246ed6a, 32'hc07697b5, 32'h403c604e};
test_output[2144] = '{32'h42ac616f};
test_index[2144] = '{2};
test_input[17160:17167] = '{32'hc29e69bc, 32'h4049e6be, 32'hc2a3de4c, 32'hc2a2f23e, 32'hc29383e9, 32'h40f87e69, 32'h420d5bf9, 32'h428cfc26};
test_output[2145] = '{32'h428cfc26};
test_index[2145] = '{7};
test_input[17168:17175] = '{32'hc1ce14fe, 32'h429d488b, 32'hc279ae3d, 32'h42a76c94, 32'hc0031caa, 32'h422f1547, 32'h42c6197d, 32'h42886f65};
test_output[2146] = '{32'h42c6197d};
test_index[2146] = '{6};
test_input[17176:17183] = '{32'h41b24d5d, 32'h40d2ff0b, 32'h42a02518, 32'hc2a91db7, 32'h40973f5a, 32'h422a5af4, 32'hc11f723b, 32'h42c2be42};
test_output[2147] = '{32'h42c2be42};
test_index[2147] = '{7};
test_input[17184:17191] = '{32'h40843576, 32'hc2090def, 32'hc24e3757, 32'h423e483b, 32'hc1d10c5a, 32'h426c53d6, 32'h423dcec1, 32'h429a6f74};
test_output[2148] = '{32'h429a6f74};
test_index[2148] = '{7};
test_input[17192:17199] = '{32'hc28fb56c, 32'hc28af33b, 32'h42c2a032, 32'h426f2b7b, 32'hc25d4e77, 32'h4253a306, 32'h42a4a734, 32'h42a5939b};
test_output[2149] = '{32'h42c2a032};
test_index[2149] = '{2};
test_input[17200:17207] = '{32'hc1912a4d, 32'h42062f99, 32'h429fcbde, 32'h42b0cd0b, 32'hc167184e, 32'h41a585c6, 32'h40be8a07, 32'hc2a10e8e};
test_output[2150] = '{32'h42b0cd0b};
test_index[2150] = '{3};
test_input[17208:17215] = '{32'hc287c8d0, 32'h42ac7a34, 32'h42815807, 32'hc289373b, 32'hc20cdd63, 32'hc22b68f3, 32'h42a6a710, 32'hc288aa2e};
test_output[2151] = '{32'h42ac7a34};
test_index[2151] = '{1};
test_input[17216:17223] = '{32'hc1f957aa, 32'h42bb6acc, 32'hc228dd45, 32'hc2914dcd, 32'hc2a799fe, 32'h426e0a63, 32'h423a84dd, 32'hc25c7027};
test_output[2152] = '{32'h42bb6acc};
test_index[2152] = '{1};
test_input[17224:17231] = '{32'h40a32577, 32'h420c83bf, 32'hc2b50db4, 32'hc0def08b, 32'h4220bf29, 32'hc20e17cb, 32'hc2371c1f, 32'h42b0fca4};
test_output[2153] = '{32'h42b0fca4};
test_index[2153] = '{7};
test_input[17232:17239] = '{32'hc2827619, 32'h42c474f1, 32'hc23a692d, 32'hc0895548, 32'hc2c428f4, 32'hc2c3fc34, 32'hc197827b, 32'hc28884cc};
test_output[2154] = '{32'h42c474f1};
test_index[2154] = '{1};
test_input[17240:17247] = '{32'hc21a13a7, 32'hc1393fcb, 32'hc1141e33, 32'hc1bc630a, 32'h4245d272, 32'h3e90b33b, 32'hc25d1ebd, 32'h42978428};
test_output[2155] = '{32'h42978428};
test_index[2155] = '{7};
test_input[17248:17255] = '{32'h4188e1d2, 32'h42a7cd17, 32'h42bebb47, 32'h408f8088, 32'hc2a36638, 32'hc1d0138d, 32'hc25a1068, 32'hc22d8178};
test_output[2156] = '{32'h42bebb47};
test_index[2156] = '{2};
test_input[17256:17263] = '{32'hc0ae1205, 32'h41e4f810, 32'hc2a57509, 32'h42ba7884, 32'hc1d52873, 32'h40ac67f1, 32'hc16728c7, 32'h42c3bed8};
test_output[2157] = '{32'h42c3bed8};
test_index[2157] = '{7};
test_input[17264:17271] = '{32'h400b39d9, 32'h417e8bba, 32'h42c4b288, 32'h425e8d24, 32'hc194b1ae, 32'hc1d02e06, 32'hc2788f13, 32'hc1ae38a9};
test_output[2158] = '{32'h42c4b288};
test_index[2158] = '{2};
test_input[17272:17279] = '{32'h42b4c4f0, 32'hc256aa26, 32'h42beadce, 32'hc18cc68b, 32'hc2a9e753, 32'hc2adb058, 32'h4205dc80, 32'hc2c07206};
test_output[2159] = '{32'h42beadce};
test_index[2159] = '{2};
test_input[17280:17287] = '{32'h41c6df68, 32'h42567122, 32'h4196b259, 32'h42aae2ca, 32'h3dad30e1, 32'h421d09bf, 32'hc102dee6, 32'hc257553b};
test_output[2160] = '{32'h42aae2ca};
test_index[2160] = '{3};
test_input[17288:17295] = '{32'hc28feb28, 32'h421800a6, 32'hc0aceed9, 32'hc2ab6425, 32'h40ee28f2, 32'h42b0b5e9, 32'hc08c769c, 32'hc24c35e6};
test_output[2161] = '{32'h42b0b5e9};
test_index[2161] = '{5};
test_input[17296:17303] = '{32'hc24d0b58, 32'hc21ede1c, 32'h42ba47fb, 32'h41ba9708, 32'hc246b988, 32'hc09263be, 32'h41d9624f, 32'hc1b9bdfd};
test_output[2162] = '{32'h42ba47fb};
test_index[2162] = '{2};
test_input[17304:17311] = '{32'hc22a1b99, 32'h4136acd7, 32'h427f2f25, 32'h426f6108, 32'hc0a13b64, 32'hc2749cd0, 32'hc2a5d314, 32'h424c873e};
test_output[2163] = '{32'h427f2f25};
test_index[2163] = '{2};
test_input[17312:17319] = '{32'hc2207bf6, 32'h423f8a9f, 32'h3fa38807, 32'h42461702, 32'h40c8b8c1, 32'h424318ba, 32'h42b5968c, 32'hc22cbb18};
test_output[2164] = '{32'h42b5968c};
test_index[2164] = '{6};
test_input[17320:17327] = '{32'h42a70ff3, 32'h42327e4e, 32'h419192a8, 32'h42c2a406, 32'hc06aa7ad, 32'h42a9c3da, 32'hc2ab7e64, 32'hc24d0464};
test_output[2165] = '{32'h42c2a406};
test_index[2165] = '{3};
test_input[17328:17335] = '{32'hc2939504, 32'h41f62f1d, 32'h429275a9, 32'h429f6016, 32'h42b1f68f, 32'h413b3420, 32'hc2c1bee8, 32'hc2969aae};
test_output[2166] = '{32'h42b1f68f};
test_index[2166] = '{4};
test_input[17336:17343] = '{32'hc228253e, 32'hc2b84e9c, 32'h42bae534, 32'h41e05d8e, 32'hc238c9d9, 32'h4291c7dc, 32'hc280ecaa, 32'hc22131e4};
test_output[2167] = '{32'h42bae534};
test_index[2167] = '{2};
test_input[17344:17351] = '{32'h42207dc4, 32'h428aa9c2, 32'hc2bdeafe, 32'hc2a470f6, 32'hc2177996, 32'hc1fd48e1, 32'hc297e95e, 32'hc293d507};
test_output[2168] = '{32'h428aa9c2};
test_index[2168] = '{1};
test_input[17352:17359] = '{32'hc2885cc5, 32'hc243610a, 32'hc242bc6a, 32'h421ea564, 32'hc1f76dc9, 32'h42605486, 32'hc09900e5, 32'hc22b5dc6};
test_output[2169] = '{32'h42605486};
test_index[2169] = '{5};
test_input[17360:17367] = '{32'h428955c6, 32'hc235bed8, 32'h422fdd0a, 32'hc23d7cff, 32'h42b61694, 32'h420f4bf3, 32'h421c2ae9, 32'hc266cf66};
test_output[2170] = '{32'h42b61694};
test_index[2170] = '{4};
test_input[17368:17375] = '{32'hc2a1518d, 32'hc2980aa9, 32'hc24c0a53, 32'h41d8a79f, 32'h427f9d09, 32'h4278f5dd, 32'h4198ddd6, 32'h429189c5};
test_output[2171] = '{32'h429189c5};
test_index[2171] = '{7};
test_input[17376:17383] = '{32'h4208945f, 32'h416fc13f, 32'hc2051bf5, 32'hc2c1aa91, 32'h4274bbe6, 32'h4298937f, 32'h41b4d78b, 32'hc29274d9};
test_output[2172] = '{32'h4298937f};
test_index[2172] = '{5};
test_input[17384:17391] = '{32'hc2722d1e, 32'h428e3bf7, 32'h42c59b67, 32'h42186543, 32'hc0bf0c0d, 32'h42995f88, 32'hc2b3b01b, 32'hc2ac51dc};
test_output[2173] = '{32'h42c59b67};
test_index[2173] = '{2};
test_input[17392:17399] = '{32'hc2a3eeaf, 32'h425cbd19, 32'h415afb74, 32'h4273361a, 32'h41f404db, 32'hc2c10f12, 32'hc1cb1f76, 32'hc297a9ef};
test_output[2174] = '{32'h4273361a};
test_index[2174] = '{3};
test_input[17400:17407] = '{32'hc27b3313, 32'h42aa04bb, 32'h414816b0, 32'h42afb073, 32'h4274e7d2, 32'h4293e7a4, 32'hc14b658f, 32'hc27f4657};
test_output[2175] = '{32'h42afb073};
test_index[2175] = '{3};
test_input[17408:17415] = '{32'hc15eb372, 32'hc28c6d33, 32'h4271db51, 32'h41aea1c6, 32'h417de8f0, 32'h421b0ea7, 32'h41877ce8, 32'h42a36323};
test_output[2176] = '{32'h42a36323};
test_index[2176] = '{7};
test_input[17416:17423] = '{32'hc2be02ad, 32'h424da9fb, 32'hc2a86f42, 32'h42103170, 32'hc05e743c, 32'hc289150d, 32'h42c798ca, 32'h428313fc};
test_output[2177] = '{32'h42c798ca};
test_index[2177] = '{6};
test_input[17424:17431] = '{32'h426b8083, 32'hc0d0fe87, 32'hc238ee9a, 32'h420394b9, 32'h41dff8a1, 32'hc229a17c, 32'h428c2373, 32'h42976c50};
test_output[2178] = '{32'h42976c50};
test_index[2178] = '{7};
test_input[17432:17439] = '{32'hc29d976e, 32'h4034369c, 32'h42aed6bb, 32'hc14eacb3, 32'hc2a34ab6, 32'h422527a2, 32'hc05d7de9, 32'h41fb4cc5};
test_output[2179] = '{32'h42aed6bb};
test_index[2179] = '{2};
test_input[17440:17447] = '{32'hc2b19a22, 32'hc29d8a6e, 32'hc21846a9, 32'h42a06b9e, 32'h41622f86, 32'h4141e9ba, 32'h411a5394, 32'h429d1b57};
test_output[2180] = '{32'h42a06b9e};
test_index[2180] = '{3};
test_input[17448:17455] = '{32'hc29814bb, 32'h42a654d7, 32'h4258e50b, 32'hc22a6284, 32'h429a1e01, 32'hbf9fa53d, 32'hc2bca1b9, 32'hc2c176f1};
test_output[2181] = '{32'h42a654d7};
test_index[2181] = '{1};
test_input[17456:17463] = '{32'h41d7c291, 32'h427f9205, 32'h415dce94, 32'hc221619a, 32'hc13d6667, 32'h42c31cb8, 32'h41ca384f, 32'h425b290e};
test_output[2182] = '{32'h42c31cb8};
test_index[2182] = '{5};
test_input[17464:17471] = '{32'h42c08a78, 32'h42b2fb45, 32'h42a2de54, 32'hc23590b3, 32'h42a1e7cc, 32'h424b670a, 32'h42adc737, 32'hc206f706};
test_output[2183] = '{32'h42c08a78};
test_index[2183] = '{0};
test_input[17472:17479] = '{32'h412fc9ab, 32'h3f88fca9, 32'h422e9cd0, 32'h42bea7dd, 32'h416b5b17, 32'h428569f3, 32'h42b238b8, 32'hc26af50b};
test_output[2184] = '{32'h42bea7dd};
test_index[2184] = '{3};
test_input[17480:17487] = '{32'h418fd94d, 32'h3f56c3af, 32'h42ae0372, 32'h429b7a1a, 32'hc1982458, 32'hc121dfb6, 32'h42686ad9, 32'hc1caacba};
test_output[2185] = '{32'h42ae0372};
test_index[2185] = '{2};
test_input[17488:17495] = '{32'hc2a0c42a, 32'hc2892572, 32'h41adc565, 32'h427e83fc, 32'h4046972f, 32'h411a18bc, 32'h42057a0e, 32'hc2654a88};
test_output[2186] = '{32'h427e83fc};
test_index[2186] = '{3};
test_input[17496:17503] = '{32'hc2301008, 32'hc291da85, 32'h41837835, 32'h42872d46, 32'h429ebafa, 32'hc217f703, 32'hc2b17fa1, 32'h429d7d2f};
test_output[2187] = '{32'h429ebafa};
test_index[2187] = '{4};
test_input[17504:17511] = '{32'hc1e0a6a7, 32'h42884cef, 32'hc28075d0, 32'h42bc2204, 32'h41356aaf, 32'hc10d942a, 32'hc1b0005f, 32'hc0cf320a};
test_output[2188] = '{32'h42bc2204};
test_index[2188] = '{3};
test_input[17512:17519] = '{32'hc27a8e67, 32'h42c4ad38, 32'h42c3d761, 32'hc234949d, 32'h4105af0d, 32'h42349877, 32'hc1284f32, 32'hc250f2dc};
test_output[2189] = '{32'h42c4ad38};
test_index[2189] = '{1};
test_input[17520:17527] = '{32'hc2a75e64, 32'hc207501c, 32'hc29b2bb4, 32'h4291814b, 32'h428c89fd, 32'h416d4799, 32'h421f464c, 32'h423fa9ce};
test_output[2190] = '{32'h4291814b};
test_index[2190] = '{3};
test_input[17528:17535] = '{32'hc155d434, 32'hc28e100f, 32'hc287a825, 32'hc24d787b, 32'hc260b3c2, 32'hc2508abe, 32'h42087216, 32'h42aa0525};
test_output[2191] = '{32'h42aa0525};
test_index[2191] = '{7};
test_input[17536:17543] = '{32'hc1fc4377, 32'h41c0c96a, 32'hc289e8f1, 32'hc221a6e9, 32'h42ab713c, 32'h42162766, 32'hc2b5630d, 32'hc2aef26b};
test_output[2192] = '{32'h42ab713c};
test_index[2192] = '{4};
test_input[17544:17551] = '{32'hc2c5c94d, 32'hc1e62072, 32'hc2743255, 32'hc1ac3703, 32'hc28f79f0, 32'h418dadd7, 32'h42af2f12, 32'hc2b925d4};
test_output[2193] = '{32'h42af2f12};
test_index[2193] = '{6};
test_input[17552:17559] = '{32'h42af993a, 32'hc2b2d848, 32'hc2b4007c, 32'h41828f8c, 32'h42b9396b, 32'hc22a2e49, 32'h42a99ad4, 32'hc124234d};
test_output[2194] = '{32'h42b9396b};
test_index[2194] = '{4};
test_input[17560:17567] = '{32'hc2a874f4, 32'hc2155ac5, 32'h429e0307, 32'h42c42de1, 32'h42486031, 32'h426f8c99, 32'h42791ae2, 32'h40daaa5a};
test_output[2195] = '{32'h42c42de1};
test_index[2195] = '{3};
test_input[17568:17575] = '{32'hc25d35d0, 32'hc15fa544, 32'hc243bb26, 32'hc1dca40d, 32'h42ba4cd8, 32'hc1dfb91a, 32'hc2ac5931, 32'h427d9d05};
test_output[2196] = '{32'h42ba4cd8};
test_index[2196] = '{4};
test_input[17576:17583] = '{32'hc084751c, 32'hc2bc28d6, 32'hc22758ce, 32'h42becc10, 32'hc1efd621, 32'h4225a6fb, 32'h414534c2, 32'hc25fcc87};
test_output[2197] = '{32'h42becc10};
test_index[2197] = '{3};
test_input[17584:17591] = '{32'hc25b22a5, 32'h41a8e7be, 32'hc25cabf2, 32'hc27e6541, 32'h427ce63e, 32'hc26caf32, 32'h4226b753, 32'h42a11307};
test_output[2198] = '{32'h42a11307};
test_index[2198] = '{7};
test_input[17592:17599] = '{32'h42a9581d, 32'h4199f23d, 32'hc2b0df9f, 32'hc2b5ba57, 32'hc2681829, 32'h428730b9, 32'hc1186a9e, 32'hc2578439};
test_output[2199] = '{32'h42a9581d};
test_index[2199] = '{0};
test_input[17600:17607] = '{32'h41c93644, 32'h4221a153, 32'hc1cf1cab, 32'hc2407ec3, 32'hc241ac9d, 32'hc1216abf, 32'hc1ddc3e9, 32'hc0f0de7b};
test_output[2200] = '{32'h4221a153};
test_index[2200] = '{1};
test_input[17608:17615] = '{32'h423dfdaf, 32'h42068f0b, 32'hc2858868, 32'h42b15955, 32'hc01bdad2, 32'hc21ecb14, 32'h42920dd2, 32'hc2a6762a};
test_output[2201] = '{32'h42b15955};
test_index[2201] = '{3};
test_input[17616:17623] = '{32'hc2aa88cc, 32'hc2ac28a8, 32'hc1b048c2, 32'hc1306410, 32'hc04263be, 32'h429a8e9e, 32'hbd8041a0, 32'h421037c1};
test_output[2202] = '{32'h429a8e9e};
test_index[2202] = '{5};
test_input[17624:17631] = '{32'hc2c1fbf2, 32'hc1dc2950, 32'hc1b56553, 32'h40e15a83, 32'h42703188, 32'hc2973f88, 32'hc277e11a, 32'h424659fd};
test_output[2203] = '{32'h42703188};
test_index[2203] = '{4};
test_input[17632:17639] = '{32'h42a91ce8, 32'h424c2ad5, 32'h40b66160, 32'hc29d0ddb, 32'h424bcd4f, 32'h42ae69b6, 32'h42996c2d, 32'hc28d59da};
test_output[2204] = '{32'h42ae69b6};
test_index[2204] = '{5};
test_input[17640:17647] = '{32'h42c6767a, 32'h41ede90f, 32'hc2694a36, 32'hc1f85e8b, 32'h42abe634, 32'hc156d785, 32'hc244cb73, 32'h402556f5};
test_output[2205] = '{32'h42c6767a};
test_index[2205] = '{0};
test_input[17648:17655] = '{32'h41179bd5, 32'hc197c8fe, 32'h418ef663, 32'h42087587, 32'h41d783ff, 32'h427dc65b, 32'hc26ffb52, 32'hc2944702};
test_output[2206] = '{32'h427dc65b};
test_index[2206] = '{5};
test_input[17656:17663] = '{32'h4203b335, 32'h41385d67, 32'h420206ba, 32'hc289a3fc, 32'hc26644a1, 32'hc131b4f9, 32'hc148438f, 32'h42b9fb74};
test_output[2207] = '{32'h42b9fb74};
test_index[2207] = '{7};
test_input[17664:17671] = '{32'h41dfd992, 32'hc2824671, 32'hc2686689, 32'h41a33dd5, 32'hc282e090, 32'hc28b8be1, 32'h422bf51b, 32'h41810b64};
test_output[2208] = '{32'h422bf51b};
test_index[2208] = '{6};
test_input[17672:17679] = '{32'hc19f1940, 32'hc2a1c5bd, 32'h425a0a27, 32'h4149c1da, 32'h428dfab3, 32'h41f04055, 32'hc2bdf181, 32'hc279832e};
test_output[2209] = '{32'h428dfab3};
test_index[2209] = '{4};
test_input[17680:17687] = '{32'hc1356cd9, 32'hc20b1207, 32'h42a9c74d, 32'h40143847, 32'hc2257495, 32'hc2b3d9c4, 32'hc1e71f12, 32'h42ba4f52};
test_output[2210] = '{32'h42ba4f52};
test_index[2210] = '{7};
test_input[17688:17695] = '{32'hc1d8159b, 32'h420e4bed, 32'h420338e1, 32'hc2c1cbc8, 32'hc290c86d, 32'h42c1ac87, 32'h3fd9075c, 32'hc252789d};
test_output[2211] = '{32'h42c1ac87};
test_index[2211] = '{5};
test_input[17696:17703] = '{32'h4208caa8, 32'hc29d2312, 32'h42b731b4, 32'h4209af5d, 32'h429d8c63, 32'hc2714719, 32'hc24392e0, 32'h4290f605};
test_output[2212] = '{32'h42b731b4};
test_index[2212] = '{2};
test_input[17704:17711] = '{32'hc285ccf0, 32'hc13402f4, 32'hc26f6594, 32'h4213285a, 32'hc182ddbd, 32'hc204352f, 32'hc0848bbb, 32'h407dd53f};
test_output[2213] = '{32'h4213285a};
test_index[2213] = '{3};
test_input[17712:17719] = '{32'hc2504f78, 32'h42b39706, 32'h423f4fcb, 32'hc2896465, 32'hc240b634, 32'h40460dd5, 32'h4229c0c7, 32'h42991623};
test_output[2214] = '{32'h42b39706};
test_index[2214] = '{1};
test_input[17720:17727] = '{32'h42a9a702, 32'h428f3612, 32'h42678cad, 32'hc288dc56, 32'hc235c1cc, 32'hc28060b1, 32'hc2396fd8, 32'hc1867539};
test_output[2215] = '{32'h42a9a702};
test_index[2215] = '{0};
test_input[17728:17735] = '{32'h41ff5ef8, 32'hc28dda33, 32'hc2bda6a0, 32'hc0e01719, 32'h429d04d9, 32'h4260c554, 32'h42477013, 32'h3f2e38f0};
test_output[2216] = '{32'h429d04d9};
test_index[2216] = '{4};
test_input[17736:17743] = '{32'h4204912d, 32'h42254aa5, 32'hc2831517, 32'h41288041, 32'hc23f6a6e, 32'hc29e7658, 32'h423d4a9b, 32'hc21bad78};
test_output[2217] = '{32'h423d4a9b};
test_index[2217] = '{6};
test_input[17744:17751] = '{32'hc19ca0cd, 32'hc1f19932, 32'hc267f215, 32'hc2942f35, 32'h41eb8a6b, 32'hc2949639, 32'h42b442c5, 32'h42ac7230};
test_output[2218] = '{32'h42b442c5};
test_index[2218] = '{6};
test_input[17752:17759] = '{32'h4249dd2c, 32'h42c5ddf7, 32'hc28ea0d5, 32'hc1d17252, 32'h41ff1c46, 32'hc2a2d0f1, 32'hc1f28768, 32'hc2be834d};
test_output[2219] = '{32'h42c5ddf7};
test_index[2219] = '{1};
test_input[17760:17767] = '{32'hc2929b67, 32'hc27c9c73, 32'hbf29ddb0, 32'h426f24f5, 32'hc211371b, 32'hc21772b3, 32'hc1d083fb, 32'h4296ce55};
test_output[2220] = '{32'h4296ce55};
test_index[2220] = '{7};
test_input[17768:17775] = '{32'hc29860e9, 32'hc18a355e, 32'h424d0d29, 32'hc2a205ff, 32'h4255360c, 32'h427bbaab, 32'h41ca9c0a, 32'hc28e479e};
test_output[2221] = '{32'h427bbaab};
test_index[2221] = '{5};
test_input[17776:17783] = '{32'h41e91eae, 32'h41a65a49, 32'hc2617ab4, 32'h4013893f, 32'hc28baf1a, 32'hc016faea, 32'hc254a347, 32'hc23a9b25};
test_output[2222] = '{32'h41e91eae};
test_index[2222] = '{0};
test_input[17784:17791] = '{32'hc21cfd47, 32'hc1945e68, 32'h428cb565, 32'h429998f2, 32'h41e4d75b, 32'h41525672, 32'h42a9fcaf, 32'h42a042f1};
test_output[2223] = '{32'h42a9fcaf};
test_index[2223] = '{6};
test_input[17792:17799] = '{32'h419e8c11, 32'h41d50452, 32'hc07e982e, 32'h42347ad5, 32'h426016d2, 32'hc2baf154, 32'hc250fce2, 32'hc2ad1b86};
test_output[2224] = '{32'h426016d2};
test_index[2224] = '{4};
test_input[17800:17807] = '{32'hc2c5360b, 32'hc2bbdde3, 32'h42c40b92, 32'hc262e040, 32'h42a186be, 32'h41a2c125, 32'hc2a382c3, 32'h422aa1a1};
test_output[2225] = '{32'h42c40b92};
test_index[2225] = '{2};
test_input[17808:17815] = '{32'h41e2bef6, 32'h41b6cc57, 32'hc12b9077, 32'h419e32bb, 32'hc1863d19, 32'h429bae1e, 32'hc1baefad, 32'hc2ba71aa};
test_output[2226] = '{32'h429bae1e};
test_index[2226] = '{5};
test_input[17816:17823] = '{32'h4293bbd5, 32'h426997c2, 32'h421bb92b, 32'h42019496, 32'hc19de08b, 32'h3f6682a3, 32'hc0e7d273, 32'h422c6b90};
test_output[2227] = '{32'h4293bbd5};
test_index[2227] = '{0};
test_input[17824:17831] = '{32'h421bb58c, 32'h42820074, 32'hc266b520, 32'h42a8f1e2, 32'h425655d0, 32'h42458feb, 32'h40906eb6, 32'h428bb541};
test_output[2228] = '{32'h42a8f1e2};
test_index[2228] = '{3};
test_input[17832:17839] = '{32'hc2bf5c9b, 32'h42731408, 32'h42a2a712, 32'h42aa2c29, 32'hc2258371, 32'h42a374fd, 32'h41c5f76e, 32'hc2ae6fe3};
test_output[2229] = '{32'h42aa2c29};
test_index[2229] = '{3};
test_input[17840:17847] = '{32'hc2a42cad, 32'h4297cbcf, 32'hc2b67372, 32'hc21652ea, 32'h429c946e, 32'h422e96fd, 32'hc0352a9e, 32'hc2948bf6};
test_output[2230] = '{32'h429c946e};
test_index[2230] = '{4};
test_input[17848:17855] = '{32'h425d0b98, 32'h4176d6c3, 32'hc2bc3cc9, 32'h42be558b, 32'hc21228db, 32'hc259129d, 32'h42a6ca48, 32'hc24d05c1};
test_output[2231] = '{32'h42be558b};
test_index[2231] = '{3};
test_input[17856:17863] = '{32'h3f243d95, 32'hc21797eb, 32'hc29a0c70, 32'h427ecb04, 32'h428522f9, 32'h401ac9ef, 32'hc2583a08, 32'h42590017};
test_output[2232] = '{32'h428522f9};
test_index[2232] = '{4};
test_input[17864:17871] = '{32'hc2961aa3, 32'h42b07562, 32'h40e7eb9d, 32'hc1cbf687, 32'h42554404, 32'hc2abce48, 32'h41a0a43f, 32'h42c5b37d};
test_output[2233] = '{32'h42c5b37d};
test_index[2233] = '{7};
test_input[17872:17879] = '{32'hc2b634aa, 32'h429eb9d7, 32'hc249bcd7, 32'h3f56ed5c, 32'h42842171, 32'h41cf18cd, 32'h428c0be3, 32'h428f25f8};
test_output[2234] = '{32'h429eb9d7};
test_index[2234] = '{1};
test_input[17880:17887] = '{32'hc184180f, 32'hc2305424, 32'h42538539, 32'hc2a66a11, 32'hc2a65305, 32'hc256b6e8, 32'h415db741, 32'hc0d4c804};
test_output[2235] = '{32'h42538539};
test_index[2235] = '{2};
test_input[17888:17895] = '{32'h42563775, 32'hc28f9660, 32'hc1a6f4a2, 32'h4199ce5a, 32'hc2a9ae33, 32'hc2aaf10e, 32'h4287ad6d, 32'h40e87c9d};
test_output[2236] = '{32'h4287ad6d};
test_index[2236] = '{6};
test_input[17896:17903] = '{32'h402f949f, 32'h42aa203d, 32'hc2558ab3, 32'hc2ab405c, 32'h422560b2, 32'h4101cf01, 32'h429fc5a4, 32'h40512f45};
test_output[2237] = '{32'h42aa203d};
test_index[2237] = '{1};
test_input[17904:17911] = '{32'h42a0da5c, 32'h425e0943, 32'h42533ddb, 32'h4059c5ca, 32'h4290afa4, 32'h4200d91e, 32'hbff21f21, 32'hbffc2608};
test_output[2238] = '{32'h42a0da5c};
test_index[2238] = '{0};
test_input[17912:17919] = '{32'h427ad2e0, 32'h4278c693, 32'h425ab47a, 32'h424ce722, 32'hc1dfb735, 32'h41ae691b, 32'h428ee99e, 32'h41a0ace6};
test_output[2239] = '{32'h428ee99e};
test_index[2239] = '{6};
test_input[17920:17927] = '{32'hc2372ce8, 32'h4281d6bc, 32'hc02059a4, 32'hc2a35206, 32'h41f3d0f6, 32'h4246bbe3, 32'hc216897e, 32'hc2bd4d5c};
test_output[2240] = '{32'h4281d6bc};
test_index[2240] = '{1};
test_input[17928:17935] = '{32'h4198d760, 32'h420f3de1, 32'h4290f11c, 32'hc17d043b, 32'h42989101, 32'h40ea07fd, 32'h42a7f435, 32'hc2a26f4a};
test_output[2241] = '{32'h42a7f435};
test_index[2241] = '{6};
test_input[17936:17943] = '{32'hc1f288a7, 32'hc23c2c7b, 32'hc20b5bbc, 32'hc2536a06, 32'hc2645960, 32'h428423e4, 32'hc254e856, 32'h42c0b444};
test_output[2242] = '{32'h42c0b444};
test_index[2242] = '{7};
test_input[17944:17951] = '{32'h42828c7e, 32'hc22c14b8, 32'h426b116b, 32'h411b0a3b, 32'hc1a88432, 32'h424cb2a0, 32'h42b19fd6, 32'h42692305};
test_output[2243] = '{32'h42b19fd6};
test_index[2243] = '{6};
test_input[17952:17959] = '{32'h42a9f897, 32'hc1599ddb, 32'h414c748f, 32'h42a38dc5, 32'hc27fdbc0, 32'hc282caf4, 32'h410ad9f8, 32'h4135d035};
test_output[2244] = '{32'h42a9f897};
test_index[2244] = '{0};
test_input[17960:17967] = '{32'h41dde0e7, 32'hc29e5476, 32'hc19741f3, 32'h428c4543, 32'h42a8e2e9, 32'hc2c6d595, 32'h422df9a6, 32'h41ffef10};
test_output[2245] = '{32'h42a8e2e9};
test_index[2245] = '{4};
test_input[17968:17975] = '{32'hc260b7a4, 32'hc28df59e, 32'hc1a44c51, 32'hc2bced9f, 32'hc01f53ef, 32'hc2bff2cc, 32'h4282361f, 32'h42ab2ef1};
test_output[2246] = '{32'h42ab2ef1};
test_index[2246] = '{7};
test_input[17976:17983] = '{32'hc2849e73, 32'h4194d711, 32'hc29e00f4, 32'hc0d2770f, 32'hc1f3a120, 32'hc15fd370, 32'hc1f8b880, 32'hc2b54290};
test_output[2247] = '{32'h4194d711};
test_index[2247] = '{1};
test_input[17984:17991] = '{32'hc28d970c, 32'h426db0b3, 32'hc1c4fe7c, 32'hc0dc3862, 32'h421b7dbc, 32'h42613cee, 32'hc1b789b5, 32'hc2516065};
test_output[2248] = '{32'h426db0b3};
test_index[2248] = '{1};
test_input[17992:17999] = '{32'h41ecb23a, 32'h429e4b82, 32'h42030705, 32'hc28fbd60, 32'hc28b1112, 32'hc141ecc7, 32'hc247b937, 32'h427adc1f};
test_output[2249] = '{32'h429e4b82};
test_index[2249] = '{1};
test_input[18000:18007] = '{32'hc232cdf5, 32'h42c7542f, 32'hc15dc678, 32'hbf978d6e, 32'hc27a5873, 32'hc1940c5b, 32'h41cab97f, 32'h41b5c167};
test_output[2250] = '{32'h42c7542f};
test_index[2250] = '{1};
test_input[18008:18015] = '{32'h421d8beb, 32'h42968ba7, 32'hc2b6c669, 32'hc17dd80e, 32'h41c71fc2, 32'h4210f66b, 32'hbeda2a23, 32'h4287d899};
test_output[2251] = '{32'h42968ba7};
test_index[2251] = '{1};
test_input[18016:18023] = '{32'h42a3883c, 32'hc1817a08, 32'hc29d0679, 32'hc1fe319c, 32'h42c13c98, 32'hc1d38e6d, 32'hc140a27e, 32'h429d0a0f};
test_output[2252] = '{32'h42c13c98};
test_index[2252] = '{4};
test_input[18024:18031] = '{32'hc2295a19, 32'hc2c0179a, 32'h42b0d284, 32'hc22176d2, 32'hc1c0b7b9, 32'h42522143, 32'hc2924a90, 32'h42c26e0e};
test_output[2253] = '{32'h42c26e0e};
test_index[2253] = '{7};
test_input[18032:18039] = '{32'h42ad9efd, 32'h42935579, 32'h42ba818c, 32'hc108d1d6, 32'h42c5b725, 32'hc0938a39, 32'h4217fa52, 32'h41fa5e5b};
test_output[2254] = '{32'h42c5b725};
test_index[2254] = '{4};
test_input[18040:18047] = '{32'h429ed493, 32'h4274b4d7, 32'hc22b9951, 32'hc2a29ba1, 32'h4288d350, 32'hc2a9d4d0, 32'h429c15d8, 32'hc1e7b4e3};
test_output[2255] = '{32'h429ed493};
test_index[2255] = '{0};
test_input[18048:18055] = '{32'hc0608a1e, 32'h418c3c9c, 32'h41c8781d, 32'h42c7c020, 32'h3fdf6114, 32'h42a66696, 32'hc23c00bc, 32'hc2c2d131};
test_output[2256] = '{32'h42c7c020};
test_index[2256] = '{3};
test_input[18056:18063] = '{32'hc1d334bd, 32'h427afc86, 32'hc12856e9, 32'h42ac63d9, 32'h417458c0, 32'hc19b88d1, 32'hc1c82bfd, 32'h409eb07e};
test_output[2257] = '{32'h42ac63d9};
test_index[2257] = '{3};
test_input[18064:18071] = '{32'hc298357b, 32'h418f63f3, 32'h41bdd069, 32'h41de1da8, 32'hc252a387, 32'hc282ea5b, 32'hc254e6a6, 32'hc2881663};
test_output[2258] = '{32'h41de1da8};
test_index[2258] = '{3};
test_input[18072:18079] = '{32'h412898d9, 32'h4271ce82, 32'hc2b2e852, 32'h420646ce, 32'hc2268828, 32'hbff03290, 32'h41d49a3b, 32'hc2ab0487};
test_output[2259] = '{32'h4271ce82};
test_index[2259] = '{1};
test_input[18080:18087] = '{32'h421c25ac, 32'hc1dc5b9f, 32'h428d69b6, 32'h42917c19, 32'h401b9648, 32'hc20d55d7, 32'hc2abdaaa, 32'hc2c34ad4};
test_output[2260] = '{32'h42917c19};
test_index[2260] = '{3};
test_input[18088:18095] = '{32'hc176ea5b, 32'h42adbe25, 32'h42b401e0, 32'h42a9a712, 32'h400bd9b0, 32'hc22b450f, 32'h412379b1, 32'hc23d81e5};
test_output[2261] = '{32'h42b401e0};
test_index[2261] = '{2};
test_input[18096:18103] = '{32'hc2281f2d, 32'hc01b2c83, 32'hc22abdbf, 32'h40c0370a, 32'h40f3e86e, 32'h41ed63a2, 32'h427a0b14, 32'h42a35da1};
test_output[2262] = '{32'h42a35da1};
test_index[2262] = '{7};
test_input[18104:18111] = '{32'h4186780e, 32'hc2a3f9a2, 32'h3fc6b22a, 32'h428a8c61, 32'h4184daab, 32'h42c7c040, 32'h4214772e, 32'h4281b6c2};
test_output[2263] = '{32'h42c7c040};
test_index[2263] = '{5};
test_input[18112:18119] = '{32'hc2b199a3, 32'h4228a437, 32'h42bbb27f, 32'hc1017622, 32'h426ec5a4, 32'h3ff6c77b, 32'h40a17e31, 32'h42043a54};
test_output[2264] = '{32'h42bbb27f};
test_index[2264] = '{2};
test_input[18120:18127] = '{32'hc2ab1704, 32'hc2a57834, 32'hc135f521, 32'hc10390ca, 32'hc232ff4a, 32'hc280ab66, 32'hc2b1d74d, 32'hc28508e7};
test_output[2265] = '{32'hc10390ca};
test_index[2265] = '{3};
test_input[18128:18135] = '{32'h4237c1ed, 32'hc2887792, 32'h42b7b531, 32'h42618862, 32'h428a21b3, 32'h42860961, 32'hc2678f6c, 32'h4232a806};
test_output[2266] = '{32'h42b7b531};
test_index[2266] = '{2};
test_input[18136:18143] = '{32'hc2b371af, 32'hc194424a, 32'hc1f59935, 32'hc003c0e0, 32'h422cfceb, 32'h41e692e7, 32'hc1a18fa7, 32'h42964afb};
test_output[2267] = '{32'h42964afb};
test_index[2267] = '{7};
test_input[18144:18151] = '{32'h4128dd0f, 32'hc2c37f9a, 32'h426146ba, 32'h40809fa7, 32'h426d82a6, 32'h418a7907, 32'h4102c5dc, 32'h42592a88};
test_output[2268] = '{32'h426d82a6};
test_index[2268] = '{4};
test_input[18152:18159] = '{32'h41b54a16, 32'hc23095bc, 32'hc156698c, 32'hc2878a4e, 32'h423d2e79, 32'h42a90c68, 32'hc26d5938, 32'h42703045};
test_output[2269] = '{32'h42a90c68};
test_index[2269] = '{5};
test_input[18160:18167] = '{32'h424bb152, 32'h42c3c13f, 32'h420738c4, 32'hc1b7b829, 32'hc290f180, 32'h42952c55, 32'h42a0f426, 32'h42069a6d};
test_output[2270] = '{32'h42c3c13f};
test_index[2270] = '{1};
test_input[18168:18175] = '{32'hc2b5c163, 32'h4229df52, 32'hc1c2aa48, 32'hc16a5f71, 32'hc2002d8d, 32'h41107cf3, 32'hc25db590, 32'hc1ddbb7a};
test_output[2271] = '{32'h4229df52};
test_index[2271] = '{1};
test_input[18176:18183] = '{32'h3f51feec, 32'hc2096c24, 32'hc191735c, 32'h429ecae4, 32'hc28c8ea0, 32'h423278d6, 32'h4274cd67, 32'hc295a7fb};
test_output[2272] = '{32'h429ecae4};
test_index[2272] = '{3};
test_input[18184:18191] = '{32'h42810930, 32'hc20f1292, 32'hc28c006b, 32'hc237278d, 32'h4204736d, 32'h41b12734, 32'h420ab775, 32'hc2c44eb1};
test_output[2273] = '{32'h42810930};
test_index[2273] = '{0};
test_input[18192:18199] = '{32'h41ab0317, 32'hc291aae0, 32'h42be87a2, 32'hc214806a, 32'hc1d72112, 32'h42b8eb48, 32'h42687f7e, 32'h42559d1e};
test_output[2274] = '{32'h42be87a2};
test_index[2274] = '{2};
test_input[18200:18207] = '{32'h42308027, 32'hc1961a7a, 32'hc174841d, 32'h429c4392, 32'h411b9ff7, 32'hc203c33e, 32'hc2ac7394, 32'hc1c02244};
test_output[2275] = '{32'h429c4392};
test_index[2275] = '{3};
test_input[18208:18215] = '{32'hc2917499, 32'hc195a1a1, 32'hc2246f6e, 32'hc204a73d, 32'h419c2fec, 32'hc2a4f916, 32'h42c05016, 32'hc2295e22};
test_output[2276] = '{32'h42c05016};
test_index[2276] = '{6};
test_input[18216:18223] = '{32'hc28f1ec3, 32'h417c4194, 32'hc221c49e, 32'h429d125d, 32'hc1d48bf4, 32'h41b2c84f, 32'h401b4d54, 32'hc2c4d4c5};
test_output[2277] = '{32'h429d125d};
test_index[2277] = '{3};
test_input[18224:18231] = '{32'h41c7a042, 32'hc26d2d14, 32'hc2a52946, 32'h41a3e89d, 32'hc2ab2b3b, 32'h42b5f2cc, 32'hc24d4602, 32'h41b1d3c9};
test_output[2278] = '{32'h42b5f2cc};
test_index[2278] = '{5};
test_input[18232:18239] = '{32'hc20e7d8e, 32'hc224c9df, 32'hbe7a63cc, 32'hc2c79fb9, 32'h426829f2, 32'h41995e81, 32'h42b202da, 32'hc2174710};
test_output[2279] = '{32'h42b202da};
test_index[2279] = '{6};
test_input[18240:18247] = '{32'h42a9f4c1, 32'hc194db59, 32'hc1d19f77, 32'h42701313, 32'h41cb83d8, 32'h42b3e984, 32'hc2c08d7c, 32'h428a7d28};
test_output[2280] = '{32'h42b3e984};
test_index[2280] = '{5};
test_input[18248:18255] = '{32'h42a3eae6, 32'hc14ec5bf, 32'h41bdd323, 32'h42c5f2ef, 32'h42292c2a, 32'hc252ce24, 32'h4281cf49, 32'hc208041e};
test_output[2281] = '{32'h42c5f2ef};
test_index[2281] = '{3};
test_input[18256:18263] = '{32'h427e9f2e, 32'h41fbc5fe, 32'h428594da, 32'hc2c5fa78, 32'hc2b94049, 32'hc29a24b8, 32'hc28a27a5, 32'hc1318323};
test_output[2282] = '{32'h428594da};
test_index[2282] = '{2};
test_input[18264:18271] = '{32'hc2b2394f, 32'hc1a5db3a, 32'hc1219ee0, 32'hc263192b, 32'hc2a62f5d, 32'h426be789, 32'hc1d9fee9, 32'h4228abef};
test_output[2283] = '{32'h426be789};
test_index[2283] = '{5};
test_input[18272:18279] = '{32'h4171973e, 32'hc2b52187, 32'hc28348a0, 32'hc22e000c, 32'hc1a10f8f, 32'hc2622610, 32'hc2a483a2, 32'h42a2ab5b};
test_output[2284] = '{32'h42a2ab5b};
test_index[2284] = '{7};
test_input[18280:18287] = '{32'hc2c5d2d8, 32'h40ac2dea, 32'h4297a129, 32'h424b0f3e, 32'hc1f498f5, 32'hc1e5a1df, 32'h42ac13c4, 32'hc299b493};
test_output[2285] = '{32'h42ac13c4};
test_index[2285] = '{6};
test_input[18288:18295] = '{32'h4291debb, 32'h424c2592, 32'hc209a9f2, 32'h40be4147, 32'hc1b5336c, 32'hc2a9c801, 32'hc104305c, 32'hc14567d3};
test_output[2286] = '{32'h4291debb};
test_index[2286] = '{0};
test_input[18296:18303] = '{32'h426cacd7, 32'hc2927aa2, 32'hc2171913, 32'hc1916f02, 32'hc19233bf, 32'hc181dd86, 32'hc28fc97a, 32'hc2a93227};
test_output[2287] = '{32'h426cacd7};
test_index[2287] = '{0};
test_input[18304:18311] = '{32'hc284aad8, 32'hc2924dfb, 32'h428a0003, 32'hc280d63f, 32'hc28e5033, 32'h42abb8f4, 32'hc2129e0e, 32'h42c7d95c};
test_output[2288] = '{32'h42c7d95c};
test_index[2288] = '{7};
test_input[18312:18319] = '{32'h4268ed31, 32'h3f256d3f, 32'hc22ae532, 32'hc2826d08, 32'h428a9026, 32'hc2b3deab, 32'h42bcf673, 32'h42213152};
test_output[2289] = '{32'h42bcf673};
test_index[2289] = '{6};
test_input[18320:18327] = '{32'hc2b9d27d, 32'hc1b31a6d, 32'hc24e5a77, 32'hc21cdda1, 32'hc1a49d48, 32'hc01dcc09, 32'hc2935678, 32'h422a61f9};
test_output[2290] = '{32'h422a61f9};
test_index[2290] = '{7};
test_input[18328:18335] = '{32'hc298a1c2, 32'h409ada17, 32'h42126979, 32'h41d46fd6, 32'h4279dc56, 32'hc237054f, 32'hc19c53b5, 32'h42bd5493};
test_output[2291] = '{32'h42bd5493};
test_index[2291] = '{7};
test_input[18336:18343] = '{32'h41656dad, 32'h428c9c21, 32'h4233c1bc, 32'hc28b2d72, 32'hc26319c8, 32'h418b27e0, 32'hc1d1ea8d, 32'h42c0e03f};
test_output[2292] = '{32'h42c0e03f};
test_index[2292] = '{7};
test_input[18344:18351] = '{32'h3f8365f0, 32'h42bea4b2, 32'h42121de8, 32'h40834f4b, 32'hc202bb04, 32'hc0cef451, 32'h42ad640c, 32'h42837d61};
test_output[2293] = '{32'h42bea4b2};
test_index[2293] = '{1};
test_input[18352:18359] = '{32'hc288cd41, 32'h42b9ac87, 32'hc24fcc99, 32'hc26cf759, 32'h4294dd0b, 32'h427c6c85, 32'hc28b4629, 32'h4161a8f9};
test_output[2294] = '{32'h42b9ac87};
test_index[2294] = '{1};
test_input[18360:18367] = '{32'hc1ef060d, 32'h41a84c1c, 32'hc2845489, 32'h42021818, 32'h3e898d18, 32'hc21e0c44, 32'hc1a4bcd1, 32'h40e70222};
test_output[2295] = '{32'h42021818};
test_index[2295] = '{3};
test_input[18368:18375] = '{32'hc175ffa0, 32'h4119585c, 32'h4283f397, 32'hc24ce029, 32'h42b33f95, 32'h4117fdcc, 32'hc117d66a, 32'h428bad57};
test_output[2296] = '{32'h42b33f95};
test_index[2296] = '{4};
test_input[18376:18383] = '{32'hc24dce82, 32'hc266e415, 32'hc2bd554e, 32'hc2989820, 32'h42bbf088, 32'h425178a5, 32'h4286160c, 32'h423fc73c};
test_output[2297] = '{32'h42bbf088};
test_index[2297] = '{4};
test_input[18384:18391] = '{32'h4287278d, 32'h402c19b1, 32'h4292d2dc, 32'h429ed405, 32'h424e9b3b, 32'h42617f98, 32'h42ab3c26, 32'h40de9079};
test_output[2298] = '{32'h42ab3c26};
test_index[2298] = '{6};
test_input[18392:18399] = '{32'h41d6a9e9, 32'h40cce86d, 32'h421a697f, 32'h4291e6f2, 32'h421f5f7c, 32'h42414dfd, 32'hc287cb56, 32'hc2c69616};
test_output[2299] = '{32'h4291e6f2};
test_index[2299] = '{3};
test_input[18400:18407] = '{32'hc1d69411, 32'hc03024c5, 32'h41dbf7ce, 32'h426ec37e, 32'hc28e3965, 32'hc1d3aa18, 32'hc268469b, 32'hc19a54b0};
test_output[2300] = '{32'h426ec37e};
test_index[2300] = '{3};
test_input[18408:18415] = '{32'h417695aa, 32'hc26c2d19, 32'hc24579de, 32'hc2a09865, 32'hc1903989, 32'h41b3dcc7, 32'h4264925b, 32'hc2a4dede};
test_output[2301] = '{32'h4264925b};
test_index[2301] = '{6};
test_input[18416:18423] = '{32'h424f9f8c, 32'h4296ac33, 32'hc2c0e57f, 32'hc0a6fd37, 32'h41a55fa1, 32'h422e089c, 32'h41fd2e47, 32'hc11593fc};
test_output[2302] = '{32'h4296ac33};
test_index[2302] = '{1};
test_input[18424:18431] = '{32'hc2975250, 32'h4177a4d7, 32'h41a56f3d, 32'hc28f2b2c, 32'hc1ffa679, 32'hbfbefd8e, 32'hc22dcf68, 32'hc25d06f0};
test_output[2303] = '{32'h41a56f3d};
test_index[2303] = '{2};
test_input[18432:18439] = '{32'h4238037e, 32'h42c13220, 32'h41c02c9b, 32'hc1fad7c3, 32'h42ad946e, 32'h41a63e2a, 32'hc24cca56, 32'hc2a78aab};
test_output[2304] = '{32'h42c13220};
test_index[2304] = '{1};
test_input[18440:18447] = '{32'h4215cfac, 32'hc23375f0, 32'h42aa1c2a, 32'hc22da92d, 32'h42abd546, 32'h42984ac2, 32'h42816506, 32'hc23f7c8b};
test_output[2305] = '{32'h42abd546};
test_index[2305] = '{4};
test_input[18448:18455] = '{32'hc22e9c68, 32'hc23b71d8, 32'hc2ba7062, 32'h41dc913a, 32'hc2a69422, 32'h424d2e52, 32'hc29ea293, 32'hc1cacf1a};
test_output[2306] = '{32'h424d2e52};
test_index[2306] = '{5};
test_input[18456:18463] = '{32'hc052cfec, 32'hc1c1ada3, 32'h4284cefa, 32'h41d48521, 32'hc28bce08, 32'hc27f0724, 32'hc2804498, 32'hc1a1cebc};
test_output[2307] = '{32'h4284cefa};
test_index[2307] = '{2};
test_input[18464:18471] = '{32'h42b419f8, 32'hc2a253f6, 32'hc2470c1a, 32'hc0ddbcd7, 32'h4282aa57, 32'hc2ba17bb, 32'h4222d27c, 32'hc1f8d1be};
test_output[2308] = '{32'h42b419f8};
test_index[2308] = '{0};
test_input[18472:18479] = '{32'h429839a6, 32'h42c217ed, 32'h4203956b, 32'h4079d859, 32'hc05981a1, 32'h42afb60a, 32'h42c05c4c, 32'h41729245};
test_output[2309] = '{32'h42c217ed};
test_index[2309] = '{1};
test_input[18480:18487] = '{32'hc21e66ac, 32'hc0283531, 32'hc1327c1a, 32'h4208c17b, 32'hc2355c25, 32'hc19753a9, 32'h4110e5b6, 32'h42c5cc35};
test_output[2310] = '{32'h42c5cc35};
test_index[2310] = '{7};
test_input[18488:18495] = '{32'h42c041ce, 32'h41fbb534, 32'hc22d1983, 32'h4268362c, 32'hc29b0053, 32'hc1d53103, 32'hc249f881, 32'h4265e857};
test_output[2311] = '{32'h42c041ce};
test_index[2311] = '{0};
test_input[18496:18503] = '{32'h41bca3f8, 32'h423d2753, 32'h42c209a2, 32'hc1cbd90c, 32'hc2a73390, 32'h42c49c21, 32'h42ad04a9, 32'h41014cab};
test_output[2312] = '{32'h42c49c21};
test_index[2312] = '{5};
test_input[18504:18511] = '{32'h426c506a, 32'hc2b71eba, 32'h422d3cc6, 32'hc20440bc, 32'hc2a2c5df, 32'hc29833dc, 32'hc25d97ed, 32'h40a055b4};
test_output[2313] = '{32'h426c506a};
test_index[2313] = '{0};
test_input[18512:18519] = '{32'hc1478661, 32'h42672f91, 32'hc2ab7d70, 32'hc1d87d34, 32'h41a5bb48, 32'hc11ffc40, 32'h42c1d8ac, 32'hc00b5fbc};
test_output[2314] = '{32'h42c1d8ac};
test_index[2314] = '{6};
test_input[18520:18527] = '{32'hc262706c, 32'h42ae6f87, 32'h426fdd8d, 32'h429ec82c, 32'hc161670a, 32'h41010c7d, 32'hc1b08fa0, 32'h42c582d6};
test_output[2315] = '{32'h42c582d6};
test_index[2315] = '{7};
test_input[18528:18535] = '{32'hc1d6ff5a, 32'h402033c4, 32'hc101e3b2, 32'hc2293124, 32'h40b9ba95, 32'hc2ae7c4d, 32'h42acd582, 32'hc27e6498};
test_output[2316] = '{32'h42acd582};
test_index[2316] = '{6};
test_input[18536:18543] = '{32'hc2c610aa, 32'hc285f593, 32'hc29dcf18, 32'hc2a7fe2b, 32'h421e23d7, 32'hc290235b, 32'h428edb6e, 32'h424c23da};
test_output[2317] = '{32'h428edb6e};
test_index[2317] = '{6};
test_input[18544:18551] = '{32'h41f5019e, 32'h42634213, 32'hc28042ea, 32'h424ce674, 32'h42b73b11, 32'h41d0f086, 32'h41fe0ade, 32'hc25b4078};
test_output[2318] = '{32'h42b73b11};
test_index[2318] = '{4};
test_input[18552:18559] = '{32'hc1406e13, 32'hc279392b, 32'h413bc531, 32'hc2682d1f, 32'hc0b1b3ce, 32'hc10ec903, 32'h42074820, 32'hc253cd9c};
test_output[2319] = '{32'h42074820};
test_index[2319] = '{6};
test_input[18560:18567] = '{32'hc1539aa3, 32'hbe2824d5, 32'hc24bea6e, 32'h42738e01, 32'hc2910feb, 32'h401c5c9f, 32'hbff51403, 32'hc25b0be9};
test_output[2320] = '{32'h42738e01};
test_index[2320] = '{3};
test_input[18568:18575] = '{32'h40dd75fc, 32'hc19504cc, 32'hc23be2b6, 32'h42c4fb73, 32'h425f428b, 32'h41f23cbb, 32'h4273b69f, 32'hc2a9c843};
test_output[2321] = '{32'h42c4fb73};
test_index[2321] = '{3};
test_input[18576:18583] = '{32'h428bf2f1, 32'hc2a94a61, 32'h42a14c89, 32'h42c110bf, 32'h41dbd275, 32'h422520e7, 32'h42c1855f, 32'h42be8b71};
test_output[2322] = '{32'h42c1855f};
test_index[2322] = '{6};
test_input[18584:18591] = '{32'h42a9ea13, 32'h4126d18b, 32'h419a4ec8, 32'hc0e2a1b0, 32'h42111974, 32'h42b13e27, 32'h417a6813, 32'h414d31ae};
test_output[2323] = '{32'h42b13e27};
test_index[2323] = '{5};
test_input[18592:18599] = '{32'h41e9b8dd, 32'h42a832e6, 32'h428f5312, 32'hc2c172d4, 32'h41cc88f4, 32'h4299097a, 32'hc1962c1f, 32'hc241b0fb};
test_output[2324] = '{32'h42a832e6};
test_index[2324] = '{1};
test_input[18600:18607] = '{32'hc229e0a5, 32'hc2469e77, 32'h429ea4e4, 32'hc16089f9, 32'h42847436, 32'hc11e8353, 32'hc1393238, 32'h41e68a38};
test_output[2325] = '{32'h429ea4e4};
test_index[2325] = '{2};
test_input[18608:18615] = '{32'h412ccd99, 32'hc2a5562c, 32'h42a413e9, 32'hc1318a78, 32'h425be74c, 32'hc26f1295, 32'h42098048, 32'hc2a035f7};
test_output[2326] = '{32'h42a413e9};
test_index[2326] = '{2};
test_input[18616:18623] = '{32'h4227b3a3, 32'hc101d35e, 32'h41f9823a, 32'hc2956466, 32'hc2aab9e3, 32'h42c6a031, 32'hc29e4eae, 32'h40db58de};
test_output[2327] = '{32'h42c6a031};
test_index[2327] = '{5};
test_input[18624:18631] = '{32'h429a3ff5, 32'h42080087, 32'h42442bf0, 32'hc2c287c7, 32'hc2a7fa3d, 32'hc1d4bf23, 32'h42b27b37, 32'hc24468d8};
test_output[2328] = '{32'h42b27b37};
test_index[2328] = '{6};
test_input[18632:18639] = '{32'h42983887, 32'hc26bbf13, 32'h42035c11, 32'hc1b4974e, 32'hc254d92b, 32'h410b3ac7, 32'hc0d3b525, 32'hc2a0ff29};
test_output[2329] = '{32'h42983887};
test_index[2329] = '{0};
test_input[18640:18647] = '{32'hc262c60a, 32'hc23da44d, 32'hc000e428, 32'h42844ec9, 32'hc2a4622f, 32'hc2769a7a, 32'hc24183bd, 32'hbf02b2ad};
test_output[2330] = '{32'h42844ec9};
test_index[2330] = '{3};
test_input[18648:18655] = '{32'h42547bf3, 32'hc1defdc8, 32'hc2274663, 32'h4182a2d6, 32'hc2c6bbf8, 32'hc28a5b56, 32'hc2b06478, 32'hc28f1bd1};
test_output[2331] = '{32'h42547bf3};
test_index[2331] = '{0};
test_input[18656:18663] = '{32'h42ad6124, 32'h4292405f, 32'hc2aa1040, 32'hc26efcc0, 32'hc29b55e1, 32'h4295cf72, 32'hc115a074, 32'h415735c0};
test_output[2332] = '{32'h42ad6124};
test_index[2332] = '{0};
test_input[18664:18671] = '{32'hc1268f0c, 32'h41ae141e, 32'h42bf27b4, 32'h41f95643, 32'hc1b26d13, 32'h42808110, 32'hc2adb917, 32'hc2a5854c};
test_output[2333] = '{32'h42bf27b4};
test_index[2333] = '{2};
test_input[18672:18679] = '{32'hc28ca2c9, 32'hc24213a7, 32'hc246c4a4, 32'h41413a33, 32'h40a8474a, 32'h40bd125f, 32'h42c55dc2, 32'hc2326af3};
test_output[2334] = '{32'h42c55dc2};
test_index[2334] = '{6};
test_input[18680:18687] = '{32'hc199c8e3, 32'h3e87ad35, 32'hc2045599, 32'h429a9f3e, 32'hc0de05ff, 32'h42a6cf54, 32'hc21d72f2, 32'hc281f41b};
test_output[2335] = '{32'h42a6cf54};
test_index[2335] = '{5};
test_input[18688:18695] = '{32'h41056bf7, 32'h42418c8c, 32'h40ca4774, 32'h4161d8c9, 32'h40c824c0, 32'hc28776dd, 32'hc270cd6c, 32'hc249420d};
test_output[2336] = '{32'h42418c8c};
test_index[2336] = '{1};
test_input[18696:18703] = '{32'hc285284b, 32'h42a8f2cd, 32'hc1831ca1, 32'h41e75b9a, 32'h424627a9, 32'h413275be, 32'h429a7a51, 32'h42a49b30};
test_output[2337] = '{32'h42a8f2cd};
test_index[2337] = '{1};
test_input[18704:18711] = '{32'h4244a8a4, 32'hc240180c, 32'h4236c088, 32'hc0abd388, 32'hc284eca7, 32'h42be1749, 32'h42ba1917, 32'h41464b97};
test_output[2338] = '{32'h42be1749};
test_index[2338] = '{5};
test_input[18712:18719] = '{32'hc201c13c, 32'hc28b21e5, 32'hc270507c, 32'h428af302, 32'h429d2510, 32'h4215e7a9, 32'h4277d084, 32'hc26f8061};
test_output[2339] = '{32'h429d2510};
test_index[2339] = '{4};
test_input[18720:18727] = '{32'hc1237f09, 32'h422563f0, 32'h4023e0ae, 32'h412a6959, 32'hc1d3bb0b, 32'hc2557b49, 32'h42be5d27, 32'hc2066b76};
test_output[2340] = '{32'h42be5d27};
test_index[2340] = '{6};
test_input[18728:18735] = '{32'h4220b75a, 32'h42095faf, 32'hc2a8dc81, 32'h42133bd9, 32'hc01e16f5, 32'h42b65575, 32'h429462a6, 32'h4287ed75};
test_output[2341] = '{32'h42b65575};
test_index[2341] = '{5};
test_input[18736:18743] = '{32'h405a3854, 32'h426f9859, 32'hc28f8f87, 32'h428868c6, 32'h4101ad9b, 32'h42b07af9, 32'hc1d6bea6, 32'h426cc99f};
test_output[2342] = '{32'h42b07af9};
test_index[2342] = '{5};
test_input[18744:18751] = '{32'hc2c5b92f, 32'hc2952906, 32'hc2c7dd90, 32'h42a09bce, 32'hc296ae1a, 32'h417ad46b, 32'hc2bd3deb, 32'hc2573b27};
test_output[2343] = '{32'h42a09bce};
test_index[2343] = '{3};
test_input[18752:18759] = '{32'h42a3b53a, 32'hc243c0e4, 32'hc273cee9, 32'h42892a17, 32'h4265ca11, 32'h4031b152, 32'hc2bcb5e5, 32'h40c5a5f7};
test_output[2344] = '{32'h42a3b53a};
test_index[2344] = '{0};
test_input[18760:18767] = '{32'h42a16aa5, 32'hc1cb3449, 32'hc276946c, 32'h4294028e, 32'hc11f1ddf, 32'h42ab9947, 32'h42a59381, 32'hc08bb450};
test_output[2345] = '{32'h42ab9947};
test_index[2345] = '{5};
test_input[18768:18775] = '{32'hc2285c8a, 32'hc1f473c9, 32'h429ca2a3, 32'h423297c6, 32'hc1a2f59b, 32'h41acad4f, 32'hc205547b, 32'hc1a1953d};
test_output[2346] = '{32'h429ca2a3};
test_index[2346] = '{2};
test_input[18776:18783] = '{32'h42bc68a6, 32'hc2574214, 32'h425cb389, 32'h42172f5f, 32'hc2b4b2d3, 32'hc237128c, 32'hbfdfe845, 32'h42a61109};
test_output[2347] = '{32'h42bc68a6};
test_index[2347] = '{0};
test_input[18784:18791] = '{32'h418f35f5, 32'h4231a1c9, 32'hc2a04385, 32'h41c3ad46, 32'h425e2228, 32'hc0d16a5b, 32'h419f9f91, 32'hc29e4966};
test_output[2348] = '{32'h425e2228};
test_index[2348] = '{4};
test_input[18792:18799] = '{32'hc25e27a6, 32'hc262d41a, 32'h4224ea5b, 32'hc206bfec, 32'h42ad4a8a, 32'hc22660a3, 32'hc29c40a8, 32'hc23106f6};
test_output[2349] = '{32'h42ad4a8a};
test_index[2349] = '{4};
test_input[18800:18807] = '{32'h426c8e9e, 32'h42a1ac34, 32'h41d0fafd, 32'hc24ca1a7, 32'h42b7bd9d, 32'hc118385d, 32'h42398acd, 32'hc1b1e5ce};
test_output[2350] = '{32'h42b7bd9d};
test_index[2350] = '{4};
test_input[18808:18815] = '{32'h42583a43, 32'hc19d58e0, 32'hc24fe2ad, 32'hc29028d7, 32'h41a55999, 32'h4281aa8a, 32'h415d0655, 32'hc29b92e1};
test_output[2351] = '{32'h4281aa8a};
test_index[2351] = '{5};
test_input[18816:18823] = '{32'hc18184cd, 32'h4287ac09, 32'hc2269112, 32'h41c8ce8e, 32'h42917062, 32'hc24ade65, 32'h428a85b9, 32'hc20facf0};
test_output[2352] = '{32'h42917062};
test_index[2352] = '{4};
test_input[18824:18831] = '{32'hc23a320a, 32'h428e891f, 32'hc2bbc305, 32'hc2b7c901, 32'hc2a9f7d1, 32'h42b39357, 32'h42872a78, 32'h42468668};
test_output[2353] = '{32'h42b39357};
test_index[2353] = '{5};
test_input[18832:18839] = '{32'h423cff01, 32'h42c253ae, 32'hc07b681c, 32'h41e44ee8, 32'h4016c99a, 32'hc2c11344, 32'h42314571, 32'h41d87eeb};
test_output[2354] = '{32'h42c253ae};
test_index[2354] = '{1};
test_input[18840:18847] = '{32'h4103d01e, 32'hc240b975, 32'h4228fc46, 32'h4270392c, 32'hc28c6ec6, 32'h42b6adf6, 32'hc2ac965d, 32'hc25079ec};
test_output[2355] = '{32'h42b6adf6};
test_index[2355] = '{5};
test_input[18848:18855] = '{32'h4231dfa0, 32'hc0a8016c, 32'hc1a1f625, 32'hc29c5d34, 32'h42097161, 32'hc07bcf6f, 32'hc2697270, 32'h42a8f44e};
test_output[2356] = '{32'h42a8f44e};
test_index[2356] = '{7};
test_input[18856:18863] = '{32'hc2a77ee0, 32'hc10daaf0, 32'hc2b28e01, 32'h42a814e1, 32'h429b7df5, 32'h42406428, 32'h42655276, 32'hc289d31e};
test_output[2357] = '{32'h42a814e1};
test_index[2357] = '{3};
test_input[18864:18871] = '{32'hc18ca09f, 32'hc21260f0, 32'hc2478a27, 32'hc2c489eb, 32'h4166460a, 32'hc20eb19b, 32'hc19c3223, 32'hc1952d14};
test_output[2358] = '{32'h4166460a};
test_index[2358] = '{4};
test_input[18872:18879] = '{32'h4138250c, 32'hc23672b4, 32'hc2bb74e6, 32'h42b6d771, 32'h428f8e7d, 32'hc2b5851c, 32'hc2a9a670, 32'hc225bce6};
test_output[2359] = '{32'h42b6d771};
test_index[2359] = '{3};
test_input[18880:18887] = '{32'h42c17726, 32'hc1827a4f, 32'h4221028b, 32'h42065cb2, 32'hc29a5197, 32'hc2aea94f, 32'hc27d6e02, 32'hc117462d};
test_output[2360] = '{32'h42c17726};
test_index[2360] = '{0};
test_input[18888:18895] = '{32'hc1253015, 32'h428019c9, 32'hc1bf3725, 32'hc2a0956c, 32'h42a7560c, 32'h42929f5a, 32'hc2a79db0, 32'h41166cbd};
test_output[2361] = '{32'h42a7560c};
test_index[2361] = '{4};
test_input[18896:18903] = '{32'h3f28149c, 32'hc2bf54e4, 32'hc23d8dd3, 32'h42a0cadf, 32'h42b1b80b, 32'h4288c1ad, 32'hc25a94af, 32'hc25716dc};
test_output[2362] = '{32'h42b1b80b};
test_index[2362] = '{4};
test_input[18904:18911] = '{32'hc24a3f0e, 32'h42087dbc, 32'hc1fd9d4c, 32'hbea0ad8f, 32'hc0710962, 32'hc1af5930, 32'hc26685fc, 32'h4202935e};
test_output[2363] = '{32'h42087dbc};
test_index[2363] = '{1};
test_input[18912:18919] = '{32'hc1f090c8, 32'hc24e708a, 32'h3fe4d10b, 32'hc21405ab, 32'h4008d273, 32'hc20b1071, 32'h42713a13, 32'h42c3b76e};
test_output[2364] = '{32'h42c3b76e};
test_index[2364] = '{7};
test_input[18920:18927] = '{32'hc2b421b8, 32'hc298ad39, 32'h420fcbdd, 32'hc2c3af42, 32'hc1da34c3, 32'hc2ae9473, 32'h4238948e, 32'hc2ba2daa};
test_output[2365] = '{32'h4238948e};
test_index[2365] = '{6};
test_input[18928:18935] = '{32'hc1b7619e, 32'hc26366df, 32'h426c80a7, 32'h41a86ec3, 32'hc25b0bd9, 32'hc2a3d204, 32'hc2152545, 32'hc2864d6b};
test_output[2366] = '{32'h426c80a7};
test_index[2366] = '{2};
test_input[18936:18943] = '{32'hc2a08164, 32'h42a2c7ee, 32'hc2af5810, 32'hc1f78e32, 32'hc0d7aff0, 32'h4246c979, 32'h42a6229b, 32'hc2c22f93};
test_output[2367] = '{32'h42a6229b};
test_index[2367] = '{6};
test_input[18944:18951] = '{32'h42a48621, 32'h42c634a4, 32'h420ac154, 32'hc2966394, 32'h42962ef0, 32'hc28d0e38, 32'hc0c28592, 32'hc252a374};
test_output[2368] = '{32'h42c634a4};
test_index[2368] = '{1};
test_input[18952:18959] = '{32'h424c1ae6, 32'hc17e8987, 32'hc1c2670c, 32'hc1927a1c, 32'h419f5eb9, 32'h42115b2a, 32'hc13a64f3, 32'hc20192a9};
test_output[2369] = '{32'h424c1ae6};
test_index[2369] = '{0};
test_input[18960:18967] = '{32'h4210302a, 32'hc1d8e56a, 32'h41f58eed, 32'hc1bb652d, 32'hc27efb40, 32'hc1cd1db1, 32'h429ec9e6, 32'h42a7eb36};
test_output[2370] = '{32'h42a7eb36};
test_index[2370] = '{7};
test_input[18968:18975] = '{32'h42b1054e, 32'hc1bcf57e, 32'hc180943c, 32'h423fe926, 32'hbfb95e25, 32'hc294c970, 32'hc203e5b1, 32'h42b082f2};
test_output[2371] = '{32'h42b1054e};
test_index[2371] = '{0};
test_input[18976:18983] = '{32'hc2a6e644, 32'h3ee4154f, 32'hbf38132b, 32'h42c3f22b, 32'hc16d4ac2, 32'hc1e29841, 32'hc23d0411, 32'hc2abeb32};
test_output[2372] = '{32'h42c3f22b};
test_index[2372] = '{3};
test_input[18984:18991] = '{32'h41ab9a13, 32'h424a708c, 32'h40d897e6, 32'hc28858e4, 32'h42b48adf, 32'hc2ac0b6e, 32'h42b13436, 32'h418dfca3};
test_output[2373] = '{32'h42b48adf};
test_index[2373] = '{4};
test_input[18992:18999] = '{32'hc2bd32de, 32'hc2b13644, 32'h429ceed1, 32'h42315b8e, 32'hc2a3ac4e, 32'h42a4c001, 32'hc2b91203, 32'hc29bcfa1};
test_output[2374] = '{32'h42a4c001};
test_index[2374] = '{5};
test_input[19000:19007] = '{32'h426f62fb, 32'h422d598b, 32'hc23971a9, 32'hc0b77e67, 32'h4069731b, 32'hc100caf6, 32'hc29aac2c, 32'hc18f1c29};
test_output[2375] = '{32'h426f62fb};
test_index[2375] = '{0};
test_input[19008:19015] = '{32'h420c955f, 32'hc2c7df39, 32'h417bd85f, 32'hc136afde, 32'hc28030b3, 32'h3e09d48b, 32'h42af4e81, 32'h42c2aa69};
test_output[2376] = '{32'h42c2aa69};
test_index[2376] = '{7};
test_input[19016:19023] = '{32'h410e4e9e, 32'h425ae5f6, 32'h4274d5b8, 32'hc21669a3, 32'h423f1057, 32'h4277509c, 32'h3f2fff77, 32'hc2c68373};
test_output[2377] = '{32'h4277509c};
test_index[2377] = '{5};
test_input[19024:19031] = '{32'hc1c02ca1, 32'h41b1b132, 32'h41a03be2, 32'hc26942d8, 32'hc2836f79, 32'hc0f548d8, 32'h42c2ae55, 32'h426173ec};
test_output[2378] = '{32'h42c2ae55};
test_index[2378] = '{6};
test_input[19032:19039] = '{32'h426d17e0, 32'h40ec25f0, 32'h42032083, 32'h4228727b, 32'hc2aa26cd, 32'h42923b8f, 32'h412a8a4a, 32'h425869fd};
test_output[2379] = '{32'h42923b8f};
test_index[2379] = '{5};
test_input[19040:19047] = '{32'h41958657, 32'h428bcd5f, 32'hc0d01a9d, 32'hc10a0948, 32'hc2a0d424, 32'hc28bd8a8, 32'h41b7f3e8, 32'hc20c2544};
test_output[2380] = '{32'h428bcd5f};
test_index[2380] = '{1};
test_input[19048:19055] = '{32'hc185190d, 32'hc274b7b2, 32'hc1a36ee4, 32'h41ea927a, 32'hc2c57614, 32'hc25154c7, 32'h417db627, 32'h417bac23};
test_output[2381] = '{32'h41ea927a};
test_index[2381] = '{3};
test_input[19056:19063] = '{32'h42c520af, 32'hc1269b0f, 32'hc2a34b71, 32'h4278ed5e, 32'h428f2366, 32'hc24dc890, 32'h42a5b99b, 32'h4280d715};
test_output[2382] = '{32'h42c520af};
test_index[2382] = '{0};
test_input[19064:19071] = '{32'h401c749c, 32'hc221354e, 32'h4282b69a, 32'h42bb2f93, 32'h41ac8df3, 32'h420d17d4, 32'h4272ca1a, 32'hc2ae3ec4};
test_output[2383] = '{32'h42bb2f93};
test_index[2383] = '{3};
test_input[19072:19079] = '{32'h42530c5b, 32'hc26148e4, 32'h4123ea40, 32'hc2443064, 32'hc2c1feba, 32'h4254b44e, 32'hc2099ad3, 32'hc27aabc5};
test_output[2384] = '{32'h4254b44e};
test_index[2384] = '{5};
test_input[19080:19087] = '{32'hc2897615, 32'hc2a5bfa3, 32'h41ed89ff, 32'hc1a382b3, 32'h4293a8e2, 32'hbf4549db, 32'hc2bfd34d, 32'hc13555a4};
test_output[2385] = '{32'h4293a8e2};
test_index[2385] = '{4};
test_input[19088:19095] = '{32'hc1949850, 32'hc17acc1c, 32'h42a0d8ed, 32'hc1f7b34e, 32'h422c6ebc, 32'hc2b68ce1, 32'h4264ab7a, 32'h42a1745b};
test_output[2386] = '{32'h42a1745b};
test_index[2386] = '{7};
test_input[19096:19103] = '{32'h421ab940, 32'h42b26b25, 32'hc15127f3, 32'h420cc1d1, 32'h4281958d, 32'hc29ea20b, 32'hc16741d4, 32'hc1034514};
test_output[2387] = '{32'h42b26b25};
test_index[2387] = '{1};
test_input[19104:19111] = '{32'h42a4abf7, 32'hc274b1c0, 32'hc1a1e9a5, 32'h42c1ef6e, 32'hc28d4e26, 32'h41bce573, 32'h3fae9733, 32'h41ab4aa5};
test_output[2388] = '{32'h42c1ef6e};
test_index[2388] = '{3};
test_input[19112:19119] = '{32'h429900fc, 32'hc20815a4, 32'h41011c1c, 32'h41dc910f, 32'hc28c710a, 32'hc2c58174, 32'hc22c666e, 32'h40e67bb8};
test_output[2389] = '{32'h429900fc};
test_index[2389] = '{0};
test_input[19120:19127] = '{32'h4239fd23, 32'h42300ca9, 32'h42afb770, 32'hc2c09e2d, 32'hc25c3888, 32'hc19a7843, 32'h42c68ec8, 32'hc21e165e};
test_output[2390] = '{32'h42c68ec8};
test_index[2390] = '{6};
test_input[19128:19135] = '{32'hc1bf235e, 32'hc2145435, 32'hc1c603b7, 32'h426b4607, 32'hc287e57a, 32'h41c4fc4e, 32'h42bebb49, 32'h42451e77};
test_output[2391] = '{32'h42bebb49};
test_index[2391] = '{6};
test_input[19136:19143] = '{32'h41da909e, 32'h4196d423, 32'hc26df430, 32'hc1fd4dcd, 32'hc1bbcaba, 32'hc1aceda8, 32'h424b0ecd, 32'h42aa701d};
test_output[2392] = '{32'h42aa701d};
test_index[2392] = '{7};
test_input[19144:19151] = '{32'hc286cac3, 32'h4283d851, 32'h41a56672, 32'hc2171b77, 32'h41cedec9, 32'h42651aca, 32'hc1ad9065, 32'h41b5c1ca};
test_output[2393] = '{32'h4283d851};
test_index[2393] = '{1};
test_input[19152:19159] = '{32'hc25a0c4f, 32'hc2bfa860, 32'h42a59bbc, 32'hc22ba52f, 32'h42816b41, 32'h4295ba89, 32'hc2a76bc6, 32'h42c45715};
test_output[2394] = '{32'h42c45715};
test_index[2394] = '{7};
test_input[19160:19167] = '{32'hc27cf60c, 32'h42844865, 32'hc2984b22, 32'hc24a62fb, 32'h41fbfc71, 32'hc08282e8, 32'h421da633, 32'h41508492};
test_output[2395] = '{32'h42844865};
test_index[2395] = '{1};
test_input[19168:19175] = '{32'h42031a0f, 32'h4085ffcd, 32'hc263d36b, 32'h3fb31298, 32'hc19bb4f9, 32'h428bfd02, 32'h41d98ca8, 32'hc29ac6ae};
test_output[2396] = '{32'h428bfd02};
test_index[2396] = '{5};
test_input[19176:19183] = '{32'hc23587bd, 32'hc0b597b6, 32'hc1b0cef2, 32'hc075f4c1, 32'hc1bf1096, 32'hc26183ee, 32'h4191ce63, 32'h42a8ca58};
test_output[2397] = '{32'h42a8ca58};
test_index[2397] = '{7};
test_input[19184:19191] = '{32'h42ba070f, 32'hc2c2b89d, 32'h427ce635, 32'h42c78fcd, 32'hc174d1fa, 32'hc2add690, 32'hc2b6c5ee, 32'hc1b7e0d8};
test_output[2398] = '{32'h42c78fcd};
test_index[2398] = '{3};
test_input[19192:19199] = '{32'h42aeb501, 32'hc2500c90, 32'hc22468f1, 32'h416c380c, 32'h419e27e4, 32'h4294e974, 32'h4194eb0a, 32'h3ef8db03};
test_output[2399] = '{32'h42aeb501};
test_index[2399] = '{0};
test_input[19200:19207] = '{32'hc050a47d, 32'h429c980e, 32'h42bd3d6e, 32'hc2a17082, 32'h428b9aa8, 32'h412be65d, 32'h419d95aa, 32'hc2baf57f};
test_output[2400] = '{32'h42bd3d6e};
test_index[2400] = '{2};
test_input[19208:19215] = '{32'h424abc25, 32'h413b43b0, 32'h41ac616d, 32'hc1905877, 32'h4252ec7a, 32'hc18df0ee, 32'hc2bd67b2, 32'hc28a273a};
test_output[2401] = '{32'h4252ec7a};
test_index[2401] = '{4};
test_input[19216:19223] = '{32'hc1a745ba, 32'h42ab115f, 32'h425b1dfe, 32'hc1c08d5f, 32'hc29df85a, 32'hc2922c0d, 32'hc2034bda, 32'hc28dd389};
test_output[2402] = '{32'h42ab115f};
test_index[2402] = '{1};
test_input[19224:19231] = '{32'hc2841c8e, 32'h4212bfaf, 32'hc269f5f5, 32'h42c2223e, 32'h42b9c115, 32'h42a7398e, 32'hc21f72d3, 32'hc288ec85};
test_output[2403] = '{32'h42c2223e};
test_index[2403] = '{3};
test_input[19232:19239] = '{32'hc20df553, 32'h42936ede, 32'hc0276a9a, 32'hc25d92b5, 32'h40440ebb, 32'hc28e42c3, 32'h422f9b72, 32'hc2bc2317};
test_output[2404] = '{32'h42936ede};
test_index[2404] = '{1};
test_input[19240:19247] = '{32'h4097e8bf, 32'hc123e285, 32'hc2a80097, 32'h42704f53, 32'hc27882fb, 32'hc26fc114, 32'h424ae25a, 32'h4156607d};
test_output[2405] = '{32'h42704f53};
test_index[2405] = '{3};
test_input[19248:19255] = '{32'h40840839, 32'h41e655e6, 32'hc2bd7712, 32'h4221c0e5, 32'hc266e2b0, 32'hc0c52fd4, 32'h42a645e8, 32'hc2a3f908};
test_output[2406] = '{32'h42a645e8};
test_index[2406] = '{6};
test_input[19256:19263] = '{32'hc21079fa, 32'hc2c54e6c, 32'h42b9c626, 32'h429e5e65, 32'h41f23a99, 32'hc1708597, 32'hc20dc195, 32'h41430f7f};
test_output[2407] = '{32'h42b9c626};
test_index[2407] = '{2};
test_input[19264:19271] = '{32'h42aee809, 32'h4270366d, 32'h4239e4d4, 32'hc1ab0dd6, 32'h42a26998, 32'h42c5c3ef, 32'hc29ce956, 32'h42a5ffc4};
test_output[2408] = '{32'h42c5c3ef};
test_index[2408] = '{5};
test_input[19272:19279] = '{32'hc14561f9, 32'hc2508ba1, 32'hc2a1faf3, 32'h423e90f5, 32'h428d57dd, 32'h42b4408d, 32'hc2824419, 32'hc2950300};
test_output[2409] = '{32'h42b4408d};
test_index[2409] = '{5};
test_input[19280:19287] = '{32'hc25c2913, 32'hc20bb236, 32'hc2b9ad46, 32'hc2258003, 32'h425c0c85, 32'h42bc3d26, 32'hc1315501, 32'h42073926};
test_output[2410] = '{32'h42bc3d26};
test_index[2410] = '{5};
test_input[19288:19295] = '{32'hc1131b68, 32'h424698e0, 32'h42b510c0, 32'h42c36749, 32'hc22bd1a8, 32'h429fda4d, 32'h42bff076, 32'h41c77d0c};
test_output[2411] = '{32'h42c36749};
test_index[2411] = '{3};
test_input[19296:19303] = '{32'h42171a53, 32'hc256a4d5, 32'hc2bcae63, 32'h42137ea8, 32'hc1eda285, 32'h42c5bb1d, 32'h4158ae0a, 32'h3e69c6e8};
test_output[2412] = '{32'h42c5bb1d};
test_index[2412] = '{5};
test_input[19304:19311] = '{32'h414df1eb, 32'h41941f4f, 32'h40514e77, 32'h419f4b8a, 32'hc2b827ba, 32'h41333c46, 32'hc2ad3472, 32'h42473dab};
test_output[2413] = '{32'h42473dab};
test_index[2413] = '{7};
test_input[19312:19319] = '{32'h4236c03c, 32'hc20ec50f, 32'h429190b0, 32'h4184478a, 32'hc215e498, 32'h42b23631, 32'hc2689ab4, 32'h4229d93e};
test_output[2414] = '{32'h42b23631};
test_index[2414] = '{5};
test_input[19320:19327] = '{32'hc24d7b19, 32'hc0b89916, 32'hc2802513, 32'h428b170f, 32'hc1935fd4, 32'h41b99087, 32'h4233af92, 32'hc2aae74a};
test_output[2415] = '{32'h428b170f};
test_index[2415] = '{3};
test_input[19328:19335] = '{32'hc25becd7, 32'h426189e9, 32'hc286d9c1, 32'hc2baf4cd, 32'h429fcbc8, 32'hc242d75b, 32'h42a10030, 32'h40a84249};
test_output[2416] = '{32'h42a10030};
test_index[2416] = '{6};
test_input[19336:19343] = '{32'hc29dfea3, 32'h4256fe20, 32'hc1184cd2, 32'h4117b6c2, 32'hc2be3008, 32'h42809a0b, 32'h4287df91, 32'h4266cf88};
test_output[2417] = '{32'h4287df91};
test_index[2417] = '{6};
test_input[19344:19351] = '{32'hc202d8aa, 32'h4212d840, 32'h41ce4f51, 32'h42b3112f, 32'hc2622c02, 32'h40f39771, 32'hc26c1810, 32'hc13ae4b1};
test_output[2418] = '{32'h42b3112f};
test_index[2418] = '{3};
test_input[19352:19359] = '{32'h4103d55b, 32'hc29077b6, 32'hc1b2a6a8, 32'h42ab8b0a, 32'h422dc043, 32'h42aecf7d, 32'hc21f3389, 32'h429ad980};
test_output[2419] = '{32'h42aecf7d};
test_index[2419] = '{5};
test_input[19360:19367] = '{32'h41c5b725, 32'hc22f8f7a, 32'hc2132df8, 32'h4256af71, 32'h429a946e, 32'hc1a3abe7, 32'hc13d9948, 32'hc0bb25db};
test_output[2420] = '{32'h429a946e};
test_index[2420] = '{4};
test_input[19368:19375] = '{32'hc2af97b2, 32'h41c69682, 32'h41e4c603, 32'h42476b84, 32'hc16636d5, 32'hc2bc0a9b, 32'hc23dcf36, 32'h42c37e28};
test_output[2421] = '{32'h42c37e28};
test_index[2421] = '{7};
test_input[19376:19383] = '{32'hc29959c8, 32'h4287985c, 32'hc0dfd45e, 32'h42b92c89, 32'h425cf9ba, 32'hc10db7e2, 32'h40e3dd2b, 32'hc28b960b};
test_output[2422] = '{32'h42b92c89};
test_index[2422] = '{3};
test_input[19384:19391] = '{32'h4296067a, 32'hc27dee57, 32'hc18623db, 32'h41fc0bfb, 32'hc236d4f1, 32'hc2391bc6, 32'h42191515, 32'hc28fde0d};
test_output[2423] = '{32'h4296067a};
test_index[2423] = '{0};
test_input[19392:19399] = '{32'h4105235d, 32'hc2058873, 32'h4013bde7, 32'h4284cd5e, 32'h41aa9265, 32'h4289c22b, 32'hc2b8bd75, 32'h4214cc21};
test_output[2424] = '{32'h4289c22b};
test_index[2424] = '{5};
test_input[19400:19407] = '{32'h425dde1f, 32'h426d0cd8, 32'hc1eee9af, 32'h4198e8fe, 32'h422c6171, 32'h41c02faa, 32'h41de63c1, 32'h426ef5e4};
test_output[2425] = '{32'h426ef5e4};
test_index[2425] = '{7};
test_input[19408:19415] = '{32'hc1adf989, 32'hc28428cb, 32'hc29b0d8e, 32'h424b36e6, 32'hc25c97b6, 32'hbf7ad98c, 32'hc253d16b, 32'h42873f47};
test_output[2426] = '{32'h42873f47};
test_index[2426] = '{7};
test_input[19416:19423] = '{32'hc2c2d39d, 32'hc28c23be, 32'hc2994fe0, 32'h42bceb01, 32'hc2189c8b, 32'h428b8600, 32'h422add0d, 32'hc28ab60f};
test_output[2427] = '{32'h42bceb01};
test_index[2427] = '{3};
test_input[19424:19431] = '{32'h424c176d, 32'hc29a1bf7, 32'hc29bec4a, 32'hc2aa844f, 32'h424f8caf, 32'hc2501dd5, 32'h41c64297, 32'hc21a04e1};
test_output[2428] = '{32'h424f8caf};
test_index[2428] = '{4};
test_input[19432:19439] = '{32'hc23edf84, 32'h420ad6ec, 32'h4291fefc, 32'h4142c8d8, 32'h426e188d, 32'h41e783d8, 32'h4297bc93, 32'h429f95bd};
test_output[2429] = '{32'h429f95bd};
test_index[2429] = '{7};
test_input[19440:19447] = '{32'hc291babb, 32'h42b79d82, 32'hc2992856, 32'hc22904fa, 32'hc2704b44, 32'h3fcfb515, 32'hc28cb31c, 32'h423ecc2f};
test_output[2430] = '{32'h42b79d82};
test_index[2430] = '{1};
test_input[19448:19455] = '{32'hc2317fda, 32'hc2af1c48, 32'hc21a9383, 32'hc1ae2008, 32'hc20045ab, 32'hc2745e8a, 32'hc28bef90, 32'hc10b9666};
test_output[2431] = '{32'hc10b9666};
test_index[2431] = '{7};
test_input[19456:19463] = '{32'hc25de93e, 32'hc2244b56, 32'hc1a4e6f7, 32'hbf10b565, 32'hc1ebf069, 32'h4018f65b, 32'h41492b57, 32'hc277fe87};
test_output[2432] = '{32'h41492b57};
test_index[2432] = '{6};
test_input[19464:19471] = '{32'h42055ca6, 32'hc21d55d6, 32'hc08fb7e7, 32'h42273c73, 32'hc22595f4, 32'h42c38e6a, 32'h4273a0d6, 32'hc29107c8};
test_output[2433] = '{32'h42c38e6a};
test_index[2433] = '{5};
test_input[19472:19479] = '{32'h420d16e5, 32'hc29ad3fa, 32'hc2a4f845, 32'h423ff971, 32'hc2b2fe89, 32'hc254f6b3, 32'hc085e4bc, 32'hc29dbc21};
test_output[2434] = '{32'h423ff971};
test_index[2434] = '{3};
test_input[19480:19487] = '{32'h428ce0a4, 32'h42059995, 32'hc2bd1519, 32'hc2c23403, 32'hc13802c6, 32'h4251758e, 32'h400647d7, 32'hc2769ac8};
test_output[2435] = '{32'h428ce0a4};
test_index[2435] = '{0};
test_input[19488:19495] = '{32'hc2485959, 32'hc27d8e38, 32'h42bc6e5e, 32'h3fe34bdb, 32'h40c1c035, 32'h423ea2d6, 32'h3f901a45, 32'hc026e001};
test_output[2436] = '{32'h42bc6e5e};
test_index[2436] = '{2};
test_input[19496:19503] = '{32'h4151f0a7, 32'h42111fe8, 32'h413897c8, 32'h42b53c71, 32'h417998a9, 32'hc2bd074f, 32'hc08db31b, 32'h41625d48};
test_output[2437] = '{32'h42b53c71};
test_index[2437] = '{3};
test_input[19504:19511] = '{32'h41dae554, 32'h42518606, 32'hc299806e, 32'h416bc4b5, 32'hc29f053e, 32'h42465753, 32'hc2678eca, 32'h4237aeb1};
test_output[2438] = '{32'h42518606};
test_index[2438] = '{1};
test_input[19512:19519] = '{32'hc2850f00, 32'h42c115a6, 32'h417071c8, 32'hc231f8fc, 32'hc2b9514b, 32'h426ea4f5, 32'h4163629f, 32'hc28de36f};
test_output[2439] = '{32'h42c115a6};
test_index[2439] = '{1};
test_input[19520:19527] = '{32'h426c4aa4, 32'h42a87eb2, 32'hc2b010bd, 32'h428572f4, 32'h422a5a99, 32'h426bc4e2, 32'hc27c57dc, 32'hc2924aa0};
test_output[2440] = '{32'h42a87eb2};
test_index[2440] = '{1};
test_input[19528:19535] = '{32'h424bec6d, 32'hc290fb7a, 32'hc231665f, 32'hc2735404, 32'h41d4043e, 32'hc19ad592, 32'hc2a14030, 32'h41af4a44};
test_output[2441] = '{32'h424bec6d};
test_index[2441] = '{0};
test_input[19536:19543] = '{32'h42897d96, 32'hc2a63242, 32'hc2a54b3f, 32'hc246b905, 32'hc2ba7bee, 32'hc05177a1, 32'hc28520ad, 32'h4210dc53};
test_output[2442] = '{32'h42897d96};
test_index[2442] = '{0};
test_input[19544:19551] = '{32'hc2a4c0e8, 32'hc2a821ef, 32'h428393d9, 32'h42b84365, 32'hc28539d6, 32'h420a0f05, 32'hc1f92cf2, 32'h41a55b9e};
test_output[2443] = '{32'h42b84365};
test_index[2443] = '{3};
test_input[19552:19559] = '{32'hc2221341, 32'hc20200d0, 32'h427e9a73, 32'h4171afc5, 32'hc1b86cf0, 32'h42bf2b25, 32'h4293ea8f, 32'h429a3176};
test_output[2444] = '{32'h42bf2b25};
test_index[2444] = '{5};
test_input[19560:19567] = '{32'h422586ac, 32'hc282b930, 32'hc2afb6a9, 32'h41b05843, 32'h42098676, 32'h41aafcf4, 32'hc0666af4, 32'h4293a85d};
test_output[2445] = '{32'h4293a85d};
test_index[2445] = '{7};
test_input[19568:19575] = '{32'h42b1e0c5, 32'h4246014d, 32'hc051016a, 32'h428e6fec, 32'hc28be49a, 32'hc2a70a4e, 32'h42878ffc, 32'h4225dc77};
test_output[2446] = '{32'h42b1e0c5};
test_index[2446] = '{0};
test_input[19576:19583] = '{32'h42aae911, 32'hc20d4cc8, 32'h420109c8, 32'hc10b97d3, 32'h42147f6b, 32'hc245bdaa, 32'hc20a4b8f, 32'h42af1720};
test_output[2447] = '{32'h42af1720};
test_index[2447] = '{7};
test_input[19584:19591] = '{32'hc015dcce, 32'h42980a70, 32'hc1e37141, 32'hc18fc69b, 32'hc1ee1d5f, 32'h420470bf, 32'hc1e452fc, 32'h4240540d};
test_output[2448] = '{32'h42980a70};
test_index[2448] = '{1};
test_input[19592:19599] = '{32'h428b2c59, 32'h423582ea, 32'hc20bb3ca, 32'hc196258c, 32'hc190c25c, 32'hc2c7169c, 32'hc2909829, 32'hc2c20fbf};
test_output[2449] = '{32'h428b2c59};
test_index[2449] = '{0};
test_input[19600:19607] = '{32'h4187429a, 32'hc2a1d146, 32'h42829fb1, 32'hc2b4757e, 32'h412e8abc, 32'h42879e5c, 32'h4272d360, 32'h42aeaaab};
test_output[2450] = '{32'h42aeaaab};
test_index[2450] = '{7};
test_input[19608:19615] = '{32'h3f1d3bc7, 32'hc2b68155, 32'hc28b8ae2, 32'h428ea321, 32'hc2827f13, 32'h41a6dfc8, 32'h417936a0, 32'h42a4b004};
test_output[2451] = '{32'h42a4b004};
test_index[2451] = '{7};
test_input[19616:19623] = '{32'hc1333c58, 32'hc055e6fd, 32'h42bfe412, 32'h42bcb7c3, 32'hc28b50b6, 32'h42a873c8, 32'h42b276ec, 32'hc2c3355a};
test_output[2452] = '{32'h42bfe412};
test_index[2452] = '{2};
test_input[19624:19631] = '{32'hc0e90619, 32'h42c74062, 32'h42c5afcf, 32'h41fa4121, 32'h42c1c50a, 32'h42935305, 32'h4203009a, 32'hc287dedf};
test_output[2453] = '{32'h42c74062};
test_index[2453] = '{1};
test_input[19632:19639] = '{32'hc2b4bc73, 32'hc0451bcc, 32'hc126556e, 32'hc29b762c, 32'h42355e39, 32'hc23c8af4, 32'h41783e5c, 32'hc208e140};
test_output[2454] = '{32'h42355e39};
test_index[2454] = '{4};
test_input[19640:19647] = '{32'hc26992ae, 32'hc2c6383b, 32'hc2a098c5, 32'hc292ea8e, 32'h419fe8e4, 32'h4271cd60, 32'hc2bb8ace, 32'h415fe7e3};
test_output[2455] = '{32'h4271cd60};
test_index[2455] = '{5};
test_input[19648:19655] = '{32'h428e0705, 32'hc1ce9ef5, 32'hc110fe58, 32'h42617fb6, 32'hc2afb7b5, 32'h4160e865, 32'h41a29844, 32'h42100817};
test_output[2456] = '{32'h428e0705};
test_index[2456] = '{0};
test_input[19656:19663] = '{32'hc1892502, 32'hc2290cd0, 32'hc2bb4b3e, 32'hc2a6b8f9, 32'hc0eec7f2, 32'hc0ebac67, 32'h42c0c2fe, 32'h415f7b95};
test_output[2457] = '{32'h42c0c2fe};
test_index[2457] = '{6};
test_input[19664:19671] = '{32'hc147b265, 32'hc2816011, 32'hc2b04d76, 32'hc28db27e, 32'h429e1ff3, 32'hc2895098, 32'h427d0a31, 32'hc107dc38};
test_output[2458] = '{32'h429e1ff3};
test_index[2458] = '{4};
test_input[19672:19679] = '{32'h4239d4d7, 32'hc2ba046f, 32'h42c66487, 32'hc2a5d949, 32'h4223b6d1, 32'hc19b7bee, 32'hc1602731, 32'hc2011b0b};
test_output[2459] = '{32'h42c66487};
test_index[2459] = '{2};
test_input[19680:19687] = '{32'hc05f63dd, 32'hc25a51bb, 32'hc282fd46, 32'h3f4f3c91, 32'hc260c20c, 32'hc25a74be, 32'hc281d7b7, 32'hc1b8073d};
test_output[2460] = '{32'h3f4f3c91};
test_index[2460] = '{3};
test_input[19688:19695] = '{32'h429bf266, 32'hc2b6308f, 32'hc2004666, 32'hc140dea4, 32'h42a49970, 32'hc2695940, 32'hc2822666, 32'h42616a5a};
test_output[2461] = '{32'h42a49970};
test_index[2461] = '{4};
test_input[19696:19703] = '{32'h42aa4cab, 32'hc1e46f03, 32'h42714449, 32'h3fde8af8, 32'h425b7cf3, 32'h42856aa0, 32'hc056ac3e, 32'h426d9af8};
test_output[2462] = '{32'h42aa4cab};
test_index[2462] = '{0};
test_input[19704:19711] = '{32'h42aebc34, 32'h42a7ba20, 32'hc2958682, 32'h428c21c6, 32'hc2384438, 32'hc26f2a12, 32'h42a1c451, 32'h42129d67};
test_output[2463] = '{32'h42aebc34};
test_index[2463] = '{0};
test_input[19712:19719] = '{32'hc1d20d97, 32'h423a6e2c, 32'hc255e778, 32'h412d36b7, 32'hc296d9cb, 32'h424f7b51, 32'h4288d5b4, 32'hc2a41371};
test_output[2464] = '{32'h4288d5b4};
test_index[2464] = '{6};
test_input[19720:19727] = '{32'h4264781f, 32'h4281c3d5, 32'h4122521f, 32'hc2a8b004, 32'hc2bafe47, 32'hc1287b7d, 32'hc292a406, 32'h42c14f98};
test_output[2465] = '{32'h42c14f98};
test_index[2465] = '{7};
test_input[19728:19735] = '{32'h42182f9c, 32'h42182d2c, 32'h42b0675d, 32'h4202f0a1, 32'h42180355, 32'hc1de9aa6, 32'hc26c6242, 32'hc1c9562e};
test_output[2466] = '{32'h42b0675d};
test_index[2466] = '{2};
test_input[19736:19743] = '{32'hc0818778, 32'hc1aef2c7, 32'hc2bfc3ec, 32'h41f81604, 32'hc2a9e4fe, 32'h425aa556, 32'h42996605, 32'h41c315a2};
test_output[2467] = '{32'h42996605};
test_index[2467] = '{6};
test_input[19744:19751] = '{32'hc214ea00, 32'h42c0916d, 32'h41055bb1, 32'hc24c47e3, 32'h425c8c30, 32'h4109c092, 32'h4234c359, 32'h41b33add};
test_output[2468] = '{32'h42c0916d};
test_index[2468] = '{1};
test_input[19752:19759] = '{32'h42a33f75, 32'hc16c6fae, 32'h41dd168c, 32'h428e1086, 32'h4287dc79, 32'h41a577ff, 32'h41cbad0f, 32'h4277cde5};
test_output[2469] = '{32'h42a33f75};
test_index[2469] = '{0};
test_input[19760:19767] = '{32'hc257d5cc, 32'hc200bc0a, 32'h427250fd, 32'hc1eaaae5, 32'h421bba26, 32'hc2b6f1c1, 32'hc2207077, 32'hc19b7171};
test_output[2470] = '{32'h427250fd};
test_index[2470] = '{2};
test_input[19768:19775] = '{32'hc28bb897, 32'h417314f0, 32'h42af18d0, 32'hc28d6a54, 32'hc2c5a17d, 32'hc25a78f7, 32'h42b6df4c, 32'hc24b08de};
test_output[2471] = '{32'h42b6df4c};
test_index[2471] = '{6};
test_input[19776:19783] = '{32'h4223e1e5, 32'h42106ed7, 32'h41cb582e, 32'h42c1cff8, 32'h428d2e12, 32'hc2538992, 32'hc198c7f4, 32'hc291d932};
test_output[2472] = '{32'h42c1cff8};
test_index[2472] = '{3};
test_input[19784:19791] = '{32'hc26cff62, 32'hc205fd02, 32'hc1a76d36, 32'h4193c066, 32'h426eb724, 32'h420a2c40, 32'hc2b8fd93, 32'h413696a1};
test_output[2473] = '{32'h426eb724};
test_index[2473] = '{4};
test_input[19792:19799] = '{32'hc118c103, 32'hc193d3cd, 32'h422e1eb9, 32'hc1a54134, 32'h40914f24, 32'h41a10a5a, 32'h42a2c70b, 32'hc14903a4};
test_output[2474] = '{32'h42a2c70b};
test_index[2474] = '{6};
test_input[19800:19807] = '{32'h4297d048, 32'h4291216e, 32'hc209077a, 32'hc0d94f7d, 32'hc2b91dc7, 32'hc263cfa9, 32'h428c9499, 32'hc24ba445};
test_output[2475] = '{32'h4297d048};
test_index[2475] = '{0};
test_input[19808:19815] = '{32'h425c4888, 32'hbf0dcf44, 32'hc221a343, 32'h420a85e4, 32'h42ba8619, 32'h4288862f, 32'h428431f6, 32'hc20d024d};
test_output[2476] = '{32'h42ba8619};
test_index[2476] = '{4};
test_input[19816:19823] = '{32'h41ca7eea, 32'hc1e924fb, 32'hc2b97619, 32'hc1ff2fa7, 32'hc23c429d, 32'hc2c4d19c, 32'h42034b44, 32'hc141c948};
test_output[2477] = '{32'h42034b44};
test_index[2477] = '{6};
test_input[19824:19831] = '{32'h42c112ea, 32'h418c37d8, 32'h42a7df3f, 32'hc29c4a13, 32'h41da690e, 32'hc2b5959f, 32'hc2bc8e78, 32'h41b352ce};
test_output[2478] = '{32'h42c112ea};
test_index[2478] = '{0};
test_input[19832:19839] = '{32'h424cb556, 32'hc2798fea, 32'hc22e3f4e, 32'h40eca9b8, 32'hc2a8fa26, 32'hc2085bd6, 32'hc21885b2, 32'hc2637fd7};
test_output[2479] = '{32'h424cb556};
test_index[2479] = '{0};
test_input[19840:19847] = '{32'h412bff82, 32'h41c6f5c3, 32'h42518c83, 32'hc2b55180, 32'hc25f522f, 32'hc149725d, 32'h412cd866, 32'hc23a5105};
test_output[2480] = '{32'h42518c83};
test_index[2480] = '{2};
test_input[19848:19855] = '{32'h4280b943, 32'h42b7de0c, 32'hc0a723c7, 32'hc2b43f69, 32'h413acc4d, 32'h421a22a2, 32'h42921015, 32'h42ade487};
test_output[2481] = '{32'h42b7de0c};
test_index[2481] = '{1};
test_input[19856:19863] = '{32'h4228b455, 32'h4293f817, 32'h422c016c, 32'h42c5d524, 32'hc2236e52, 32'h4206a54d, 32'h424a8c1c, 32'hc1d5c20a};
test_output[2482] = '{32'h42c5d524};
test_index[2482] = '{3};
test_input[19864:19871] = '{32'hc13ecbcf, 32'hc11508c6, 32'h4247bee3, 32'h42184e99, 32'h414ad826, 32'hc27143ef, 32'h4298b00f, 32'hc2385ffa};
test_output[2483] = '{32'h4298b00f};
test_index[2483] = '{6};
test_input[19872:19879] = '{32'hc2078841, 32'hc0a48b10, 32'hc186f877, 32'h428aa802, 32'hc1a85770, 32'hc2a321f8, 32'h42a329bf, 32'hc136ea57};
test_output[2484] = '{32'h42a329bf};
test_index[2484] = '{6};
test_input[19880:19887] = '{32'h40b7c5cc, 32'hc2b9fa1b, 32'h42156286, 32'h416c64b2, 32'h428150d2, 32'hc2afc029, 32'h41ece329, 32'hc10f89eb};
test_output[2485] = '{32'h428150d2};
test_index[2485] = '{4};
test_input[19888:19895] = '{32'hc2380d51, 32'hc29dbc80, 32'h4230fd95, 32'h427b0bc0, 32'hc2941cc2, 32'hc25c2834, 32'h42a77b41, 32'h42b5b0a8};
test_output[2486] = '{32'h42b5b0a8};
test_index[2486] = '{7};
test_input[19896:19903] = '{32'hc2a57aea, 32'hc2781648, 32'hc2877788, 32'h429c756c, 32'hc288a31c, 32'hc2bb7f9b, 32'hc2974123, 32'h429a10fe};
test_output[2487] = '{32'h429c756c};
test_index[2487] = '{3};
test_input[19904:19911] = '{32'hc284854e, 32'hc2b5e4df, 32'h41e2adcd, 32'h40452dff, 32'hc2805e69, 32'h428ee92e, 32'h41b892b1, 32'h419c60c6};
test_output[2488] = '{32'h428ee92e};
test_index[2488] = '{5};
test_input[19912:19919] = '{32'hc252dbab, 32'hc14026cb, 32'h4214e7f5, 32'h42b5a570, 32'h4298ef21, 32'h428c2a0b, 32'h40f14008, 32'hc2630b5e};
test_output[2489] = '{32'h42b5a570};
test_index[2489] = '{3};
test_input[19920:19927] = '{32'hc1c34005, 32'hc293cf33, 32'h41b6c928, 32'h42c5d126, 32'h419e0ad1, 32'hc20f9fac, 32'h427c4ee6, 32'h42b7b8d1};
test_output[2490] = '{32'h42c5d126};
test_index[2490] = '{3};
test_input[19928:19935] = '{32'h42867250, 32'h3f8b51af, 32'h40c839a2, 32'h429abf5d, 32'hc2221d98, 32'h410db19f, 32'h419670cf, 32'hc233d9da};
test_output[2491] = '{32'h429abf5d};
test_index[2491] = '{3};
test_input[19936:19943] = '{32'h427cb75f, 32'h429499b2, 32'h42625a8b, 32'h40fd61bd, 32'hc27e60ad, 32'hc287cb49, 32'h42a9fffd, 32'hc27b1845};
test_output[2492] = '{32'h42a9fffd};
test_index[2492] = '{6};
test_input[19944:19951] = '{32'h4284f359, 32'h41d6f250, 32'h42862af3, 32'h42a66997, 32'hc298ccf5, 32'hc2b72f23, 32'h423bbde9, 32'h41452203};
test_output[2493] = '{32'h42a66997};
test_index[2493] = '{3};
test_input[19952:19959] = '{32'h41b03ee2, 32'hc1cbe0ec, 32'hc2c50b67, 32'hc23b531d, 32'h42675059, 32'hc141fd1a, 32'hc28dd27a, 32'hc190bb0c};
test_output[2494] = '{32'h42675059};
test_index[2494] = '{4};
test_input[19960:19967] = '{32'h4211dff3, 32'hc233f629, 32'hc274b75f, 32'h4278493c, 32'hc07bf2e3, 32'hc147cb9f, 32'h4099101f, 32'hc14cd8ef};
test_output[2495] = '{32'h4278493c};
test_index[2495] = '{3};
test_input[19968:19975] = '{32'h420c16e0, 32'h429d6068, 32'hc2c6a50c, 32'hc2a4a01f, 32'h41b81430, 32'hc25c146b, 32'hc2ae057e, 32'h42564ff4};
test_output[2496] = '{32'h429d6068};
test_index[2496] = '{1};
test_input[19976:19983] = '{32'h42a307c6, 32'h4281376a, 32'h4244d42e, 32'h42b14e34, 32'h42a0215e, 32'h42937861, 32'h42a9e6c0, 32'hc0a12507};
test_output[2497] = '{32'h42b14e34};
test_index[2497] = '{3};
test_input[19984:19991] = '{32'hc20e8b6f, 32'h425600a5, 32'h42bb0b7c, 32'hc28cee1f, 32'h4196f005, 32'h42064e29, 32'h4225d4b2, 32'hc15baaf8};
test_output[2498] = '{32'h42bb0b7c};
test_index[2498] = '{2};
test_input[19992:19999] = '{32'hc28ff2d2, 32'hc2a878ea, 32'h41098c31, 32'hc19249ac, 32'hc18e0330, 32'hc2b484a4, 32'h40a2875d, 32'h4253c638};
test_output[2499] = '{32'h4253c638};
test_index[2499] = '{7};
test_input[20000:20007] = '{32'h4203230e, 32'hc2c5f1c1, 32'h42b4dcfb, 32'h421a8fce, 32'hc2409c0f, 32'h425c553b, 32'h419bf32c, 32'hc205a918};
test_output[2500] = '{32'h42b4dcfb};
test_index[2500] = '{2};
test_input[20008:20015] = '{32'h424800d1, 32'hc29386ce, 32'hc2b3a558, 32'h428638b7, 32'hc28e1303, 32'hc25a86ba, 32'h41fe4324, 32'h42663f6d};
test_output[2501] = '{32'h428638b7};
test_index[2501] = '{3};
test_input[20016:20023] = '{32'h4272d595, 32'h42c02330, 32'h42c4cb3b, 32'hc199c95f, 32'h427f9e5e, 32'h42a446f3, 32'h4204359f, 32'hc11ed965};
test_output[2502] = '{32'h42c4cb3b};
test_index[2502] = '{2};
test_input[20024:20031] = '{32'h428bad65, 32'hc26e5c20, 32'h41854bef, 32'hc2a57416, 32'hc28e7aa5, 32'h42b21d14, 32'hc23a37de, 32'hc1f02b79};
test_output[2503] = '{32'h42b21d14};
test_index[2503] = '{5};
test_input[20032:20039] = '{32'hc2a3970a, 32'h42247d0b, 32'h42a8dab1, 32'h42b6b45f, 32'hc290a9df, 32'h42a1cbd3, 32'h41d72bf5, 32'h412d0ed7};
test_output[2504] = '{32'h42b6b45f};
test_index[2504] = '{3};
test_input[20040:20047] = '{32'h425608bb, 32'hc2394d81, 32'h41d4f506, 32'h428fb4ea, 32'hc2c5a72e, 32'hc2c159e0, 32'hc21fbdf8, 32'h41385dfc};
test_output[2505] = '{32'h428fb4ea};
test_index[2505] = '{3};
test_input[20048:20055] = '{32'h415f9151, 32'h428cd9a1, 32'h426a6b33, 32'h424805f9, 32'h41f295c7, 32'h413fef6f, 32'h42a4ffe9, 32'h42c67f2c};
test_output[2506] = '{32'h42c67f2c};
test_index[2506] = '{7};
test_input[20056:20063] = '{32'h426f082e, 32'h420f6d28, 32'hc10dcfc5, 32'h42c0bacc, 32'h427fc5ae, 32'h4186d52f, 32'h42aabc03, 32'h41be74bb};
test_output[2507] = '{32'h42c0bacc};
test_index[2507] = '{3};
test_input[20064:20071] = '{32'h42a1baa4, 32'hc20a9397, 32'h426aca69, 32'h3f041200, 32'h41828067, 32'h4230a473, 32'hc2b37b92, 32'h423c625d};
test_output[2508] = '{32'h42a1baa4};
test_index[2508] = '{0};
test_input[20072:20079] = '{32'h429acbda, 32'hc181145b, 32'h41a83996, 32'hc20974e5, 32'hc29f2206, 32'h42994552, 32'hc2a1ff2a, 32'hc263863e};
test_output[2509] = '{32'h429acbda};
test_index[2509] = '{0};
test_input[20080:20087] = '{32'hc20cb56f, 32'hc2c3c21b, 32'h420bbba3, 32'hc2616ac2, 32'h4236baf4, 32'hc1e52861, 32'hc1cb9cd9, 32'h424dab0c};
test_output[2510] = '{32'h424dab0c};
test_index[2510] = '{7};
test_input[20088:20095] = '{32'hc28e2a0f, 32'h411da713, 32'h42605e3d, 32'hc297470f, 32'hc2ac9d1c, 32'h41575180, 32'hc17c0c87, 32'h420c24af};
test_output[2511] = '{32'h42605e3d};
test_index[2511] = '{2};
test_input[20096:20103] = '{32'hc218219e, 32'h42968f0b, 32'h410caca9, 32'hc23a8b40, 32'h428ec196, 32'hc1f3d315, 32'h42728b8f, 32'h424c9ff1};
test_output[2512] = '{32'h42968f0b};
test_index[2512] = '{1};
test_input[20104:20111] = '{32'hc1ab14fc, 32'hc2afbdeb, 32'h4177ad49, 32'hc0c58b2e, 32'hc25d9207, 32'h423d2197, 32'h41de5c22, 32'h4277ca74};
test_output[2513] = '{32'h4277ca74};
test_index[2513] = '{7};
test_input[20112:20119] = '{32'h42973d3b, 32'h41abfde8, 32'hc20e901d, 32'h405e229b, 32'h42058f3d, 32'hc26f1c32, 32'h4240db64, 32'h4266eb0b};
test_output[2514] = '{32'h42973d3b};
test_index[2514] = '{0};
test_input[20120:20127] = '{32'hc2b7156c, 32'hc2b28ee5, 32'h40a52cda, 32'h4265cd97, 32'h41c1f7df, 32'h4123a95d, 32'hc2abfef7, 32'h414d463d};
test_output[2515] = '{32'h4265cd97};
test_index[2515] = '{3};
test_input[20128:20135] = '{32'h429ba403, 32'h42c4a4ae, 32'h41547ab1, 32'hc242b5ba, 32'h42c06f56, 32'hc21dcd60, 32'h42ae275e, 32'hc1b71892};
test_output[2516] = '{32'h42c4a4ae};
test_index[2516] = '{1};
test_input[20136:20143] = '{32'hc2017547, 32'h41bb1ae9, 32'h41821d5d, 32'h4285e8eb, 32'h42426659, 32'hc0880f48, 32'h4019d92b, 32'h42c2d78b};
test_output[2517] = '{32'h42c2d78b};
test_index[2517] = '{7};
test_input[20144:20151] = '{32'h42b56c35, 32'hc2a83935, 32'hc2c4f7d3, 32'hc2bfe303, 32'hc28060fa, 32'h412da4a3, 32'h428c75a2, 32'h411b0407};
test_output[2518] = '{32'h42b56c35};
test_index[2518] = '{0};
test_input[20152:20159] = '{32'hc26a74c0, 32'hc18ee279, 32'h42943500, 32'h42aea34a, 32'h41f160cb, 32'h4247637b, 32'hc1dd1f55, 32'hc220b707};
test_output[2519] = '{32'h42aea34a};
test_index[2519] = '{3};
test_input[20160:20167] = '{32'h42c5fa46, 32'hc080a403, 32'h4210964f, 32'h42c109ae, 32'h4275db66, 32'hc11d1a7b, 32'h429e03bb, 32'h420589c0};
test_output[2520] = '{32'h42c5fa46};
test_index[2520] = '{0};
test_input[20168:20175] = '{32'h4288ceb1, 32'hc2ac4fae, 32'hc2b2b86a, 32'h4197500d, 32'h428812f4, 32'h429d5c97, 32'hc24e2edd, 32'hc200736a};
test_output[2521] = '{32'h429d5c97};
test_index[2521] = '{5};
test_input[20176:20183] = '{32'hc202396f, 32'hc198cc35, 32'h42bf1bb2, 32'h4264f218, 32'h420bd4f8, 32'hc1ba5550, 32'h429ccc34, 32'hc264db18};
test_output[2522] = '{32'h42bf1bb2};
test_index[2522] = '{2};
test_input[20184:20191] = '{32'h423e6f8f, 32'h4299a5de, 32'hc2a5c743, 32'h41cc2d84, 32'hc2a9ab58, 32'h419a96ef, 32'h42a334ec, 32'hc28ed04f};
test_output[2523] = '{32'h42a334ec};
test_index[2523] = '{6};
test_input[20192:20199] = '{32'hc16cebe1, 32'hc25a1e09, 32'hc22c0395, 32'h420ebae5, 32'hc2ac5087, 32'hc22bc1b8, 32'hc25f4d55, 32'h4274ade7};
test_output[2524] = '{32'h4274ade7};
test_index[2524] = '{7};
test_input[20200:20207] = '{32'hc27542ca, 32'hc0e8bf61, 32'hc265fc79, 32'hc210eda9, 32'h3f2a8835, 32'h4175c9e4, 32'hc12bab91, 32'hc289a5c0};
test_output[2525] = '{32'h4175c9e4};
test_index[2525] = '{5};
test_input[20208:20215] = '{32'h427999b0, 32'h422be2af, 32'hc0b2cc80, 32'hc2bb5ddb, 32'hc119061b, 32'hc17c62d2, 32'hc1120666, 32'hbe7c2f4f};
test_output[2526] = '{32'h427999b0};
test_index[2526] = '{0};
test_input[20216:20223] = '{32'h40d5af17, 32'h4208e46a, 32'h408d8b44, 32'h427f9350, 32'h4118b902, 32'h40fcd1ce, 32'h40e980e5, 32'h41003c82};
test_output[2527] = '{32'h427f9350};
test_index[2527] = '{3};
test_input[20224:20231] = '{32'hc2bc4605, 32'hc29d424f, 32'hc240d1a5, 32'hc2b1d326, 32'h42bdb9fc, 32'h424c79c7, 32'h42940a6f, 32'hc1ed7554};
test_output[2528] = '{32'h42bdb9fc};
test_index[2528] = '{4};
test_input[20232:20239] = '{32'h41b370b9, 32'hc2a5850b, 32'hc1bbc25f, 32'h425b5e03, 32'hc1db4b3d, 32'hc2b7bfe8, 32'h4215c4d7, 32'h4246ca5a};
test_output[2529] = '{32'h425b5e03};
test_index[2529] = '{3};
test_input[20240:20247] = '{32'hc202e573, 32'h41e10e8e, 32'h411f221e, 32'h4216a8dd, 32'hc27ea5f8, 32'hc2a6a005, 32'hc21186f6, 32'hc2a7aaa1};
test_output[2530] = '{32'h4216a8dd};
test_index[2530] = '{3};
test_input[20248:20255] = '{32'h42b7d397, 32'h40a9737b, 32'h42991f85, 32'h42300729, 32'hc2b34572, 32'hc1c6eb66, 32'h41a56038, 32'h42ac4b7d};
test_output[2531] = '{32'h42b7d397};
test_index[2531] = '{0};
test_input[20256:20263] = '{32'hc2ab71e8, 32'hc250dbc1, 32'hc20401ce, 32'hbfe09524, 32'hc23bc10e, 32'hc2a87966, 32'h42161fa8, 32'hc1c2d010};
test_output[2532] = '{32'h42161fa8};
test_index[2532] = '{6};
test_input[20264:20271] = '{32'hc2319f54, 32'hc2ac38b6, 32'h42565179, 32'hc213a926, 32'h41b869b3, 32'h400ca6b7, 32'hc25aca2d, 32'h42740a72};
test_output[2533] = '{32'h42740a72};
test_index[2533] = '{7};
test_input[20272:20279] = '{32'h4262e326, 32'h419a97f0, 32'hc2b1a082, 32'h425ebf20, 32'hc2b91326, 32'hc2a413bb, 32'h41a5c0c8, 32'h42acd794};
test_output[2534] = '{32'h42acd794};
test_index[2534] = '{7};
test_input[20280:20287] = '{32'h428ac6fb, 32'hc2bdc8c0, 32'hc280ae8c, 32'h4276191d, 32'h42acf5c6, 32'h419affc6, 32'h428a0654, 32'hc2333105};
test_output[2535] = '{32'h42acf5c6};
test_index[2535] = '{4};
test_input[20288:20295] = '{32'hc2582965, 32'hc2c7d2d0, 32'h42c48b44, 32'hc259deba, 32'hc272612c, 32'hc23e00d5, 32'h42729d0a, 32'h42b3450c};
test_output[2536] = '{32'h42c48b44};
test_index[2536] = '{2};
test_input[20296:20303] = '{32'hc27fdb37, 32'hc228c8a7, 32'hc28978dc, 32'h42a9de02, 32'hc2c29cba, 32'hc1e2b7d9, 32'h42bd96e0, 32'hc2419247};
test_output[2537] = '{32'h42bd96e0};
test_index[2537] = '{6};
test_input[20304:20311] = '{32'h426b7521, 32'hc0eaae9e, 32'hc1d5426a, 32'hc24a5ee5, 32'h42878f94, 32'hc2787125, 32'h41360a6f, 32'h4267a412};
test_output[2538] = '{32'h42878f94};
test_index[2538] = '{4};
test_input[20312:20319] = '{32'h42044f6f, 32'hc2a13d59, 32'hc1c91666, 32'hc2849198, 32'hc29d5cc0, 32'hc12ae5be, 32'h42009559, 32'hc1885ead};
test_output[2539] = '{32'h42044f6f};
test_index[2539] = '{0};
test_input[20320:20327] = '{32'hc24ef297, 32'h429d3fff, 32'h415af171, 32'hc28808b7, 32'h4270b2a5, 32'hc1e75bdc, 32'hc2c2b2fc, 32'h42789cda};
test_output[2540] = '{32'h429d3fff};
test_index[2540] = '{1};
test_input[20328:20335] = '{32'hc2c742a0, 32'h42a7dc16, 32'hc17942da, 32'hc2a2e315, 32'hc108d2d7, 32'h421e3d9d, 32'hc1d90385, 32'hc2a0beee};
test_output[2541] = '{32'h42a7dc16};
test_index[2541] = '{1};
test_input[20336:20343] = '{32'hc1190016, 32'h408afbb8, 32'h42b08527, 32'h4215ee06, 32'hc2611f10, 32'hc1e6997c, 32'hc2b55a23, 32'hc2a8aba2};
test_output[2542] = '{32'h42b08527};
test_index[2542] = '{2};
test_input[20344:20351] = '{32'hc2259305, 32'hc180736b, 32'hc14234ba, 32'hc05ce337, 32'hc25d02aa, 32'hc205f038, 32'hc25da2f8, 32'hc2157e23};
test_output[2543] = '{32'hc05ce337};
test_index[2543] = '{3};
test_input[20352:20359] = '{32'h41814e2b, 32'h42c521ef, 32'h4187c434, 32'hc22c6845, 32'h42c7273e, 32'hc1c8344e, 32'h4271f773, 32'hc119067c};
test_output[2544] = '{32'h42c7273e};
test_index[2544] = '{4};
test_input[20360:20367] = '{32'hc28bf7a4, 32'h42c406fa, 32'hc224f0e5, 32'hc263762f, 32'hc2355704, 32'h4264793f, 32'h40e1eb0d, 32'hc263ee1b};
test_output[2545] = '{32'h42c406fa};
test_index[2545] = '{1};
test_input[20368:20375] = '{32'h42adcfda, 32'hc17cca5e, 32'h41ffa182, 32'h428a4c06, 32'h4246d492, 32'h417f3c08, 32'h41988ce3, 32'h42456d31};
test_output[2546] = '{32'h42adcfda};
test_index[2546] = '{0};
test_input[20376:20383] = '{32'hbecd8bea, 32'hc2139bbd, 32'h413ab62f, 32'hc249ea1c, 32'hc266ef72, 32'hc271998b, 32'hc179d319, 32'h4235f916};
test_output[2547] = '{32'h4235f916};
test_index[2547] = '{7};
test_input[20384:20391] = '{32'hc1a8c479, 32'hc296d621, 32'h41b9b1ed, 32'hc28d6d59, 32'hc1414ab3, 32'h42a647cd, 32'hc22bf088, 32'h40e64126};
test_output[2548] = '{32'h42a647cd};
test_index[2548] = '{5};
test_input[20392:20399] = '{32'h41dd6f5a, 32'h4258bf2b, 32'hc161eaab, 32'hc2ad6a3a, 32'h4184d684, 32'h42b6fb4a, 32'hc079304f, 32'hc1947b6b};
test_output[2549] = '{32'h42b6fb4a};
test_index[2549] = '{5};
test_input[20400:20407] = '{32'hc2719a1e, 32'h42407d42, 32'hc2c3b56e, 32'hc08c648b, 32'h426089ae, 32'hc216907b, 32'h3fb16711, 32'hc17e6921};
test_output[2550] = '{32'h426089ae};
test_index[2550] = '{4};
test_input[20408:20415] = '{32'hc1c244da, 32'hc23e950b, 32'h428fb9ab, 32'h4207e6dd, 32'h42001da0, 32'hc222974a, 32'h429bddac, 32'h428cda0f};
test_output[2551] = '{32'h429bddac};
test_index[2551] = '{6};
test_input[20416:20423] = '{32'hc293f25b, 32'hc2afe28a, 32'h42af1841, 32'hc29eeee1, 32'h410a69c4, 32'h40c3f642, 32'hc24ac056, 32'h421a0c1b};
test_output[2552] = '{32'h42af1841};
test_index[2552] = '{2};
test_input[20424:20431] = '{32'hc20d1c57, 32'hc0c6e310, 32'h42683bb2, 32'hc1e2cb4e, 32'h42970741, 32'hc21b9eac, 32'hc2baba49, 32'h42ab2966};
test_output[2553] = '{32'h42ab2966};
test_index[2553] = '{7};
test_input[20432:20439] = '{32'h428e6de5, 32'hc1ec3324, 32'h419e1cec, 32'h424903af, 32'h4173feaf, 32'h426863a8, 32'hc2b8a718, 32'hc183c13d};
test_output[2554] = '{32'h428e6de5};
test_index[2554] = '{0};
test_input[20440:20447] = '{32'hc21ef82b, 32'hc1ad9c86, 32'hc2b31745, 32'hc2644a01, 32'h3f10b978, 32'hbf871b15, 32'hc2957dea, 32'hc01a5d62};
test_output[2555] = '{32'h3f10b978};
test_index[2555] = '{4};
test_input[20448:20455] = '{32'h42c39b13, 32'hc2c236cb, 32'h42c7ab74, 32'hc279ae63, 32'hc2af7caf, 32'h4282548b, 32'h41af6dcf, 32'hc25afb54};
test_output[2556] = '{32'h42c7ab74};
test_index[2556] = '{2};
test_input[20456:20463] = '{32'h41b232ea, 32'h41b5d1b3, 32'hc2aff129, 32'hc2a9eae8, 32'hc1f36cf5, 32'h42c76dfd, 32'h42748396, 32'hc2a32342};
test_output[2557] = '{32'h42c76dfd};
test_index[2557] = '{5};
test_input[20464:20471] = '{32'hc2a1e313, 32'hc2b46d86, 32'hc1d34526, 32'h415362f6, 32'hc2b8e2a4, 32'hc1c1843b, 32'hc2b52d12, 32'hc0e4d11b};
test_output[2558] = '{32'h415362f6};
test_index[2558] = '{3};
test_input[20472:20479] = '{32'hc27fec57, 32'h421a98c4, 32'h42a1d53c, 32'h40237ff2, 32'h408e320b, 32'h41457fe7, 32'hc1e938b3, 32'h4102ca34};
test_output[2559] = '{32'h42a1d53c};
test_index[2559] = '{2};
test_input[20480:20487] = '{32'hc296ae22, 32'h423d2fc5, 32'h426d50e4, 32'h419b59be, 32'h42a8efe5, 32'h42351b20, 32'hc2b9b3d7, 32'h41cc5133};
test_output[2560] = '{32'h42a8efe5};
test_index[2560] = '{4};
test_input[20488:20495] = '{32'hc294e3db, 32'h3fd39884, 32'h42892dcc, 32'hbf3227aa, 32'h4103902c, 32'h4297f968, 32'hc2b5d027, 32'h42c10f8d};
test_output[2561] = '{32'h42c10f8d};
test_index[2561] = '{7};
test_input[20496:20503] = '{32'hc22d3463, 32'h42c3eb71, 32'hc10415f4, 32'h429dbd89, 32'hbfe54940, 32'hc2c62334, 32'hc26ff76f, 32'hc2bc84b7};
test_output[2562] = '{32'h42c3eb71};
test_index[2562] = '{1};
test_input[20504:20511] = '{32'hc07e8fbb, 32'h4004a32c, 32'hc25ba19d, 32'h420e2166, 32'hc21d176c, 32'hc1ccfd39, 32'h428509fb, 32'hc2bbdf10};
test_output[2563] = '{32'h428509fb};
test_index[2563] = '{6};
test_input[20512:20519] = '{32'hc1e88a26, 32'h42af80c5, 32'h41ff491c, 32'h4020ea2a, 32'h41441d0a, 32'h42a7b2ec, 32'hc2181339, 32'hc2416adb};
test_output[2564] = '{32'h42af80c5};
test_index[2564] = '{1};
test_input[20520:20527] = '{32'hc1487e9e, 32'hc2a90bb1, 32'hc18b3f84, 32'hc25ad02a, 32'hc28b3c9d, 32'hc242fa99, 32'hc1378578, 32'hc22a55f0};
test_output[2565] = '{32'hc1378578};
test_index[2565] = '{6};
test_input[20528:20535] = '{32'hc29333dd, 32'h42a69f71, 32'h42242032, 32'h429fe6fd, 32'hc2ac2acd, 32'h41a38a48, 32'hc253da1b, 32'hc21724a2};
test_output[2566] = '{32'h42a69f71};
test_index[2566] = '{1};
test_input[20536:20543] = '{32'hc2466eef, 32'h428f9d97, 32'hc03c2cb4, 32'hc27962c4, 32'h4215b341, 32'hc2970a72, 32'hc28a9a3a, 32'h429fc65e};
test_output[2567] = '{32'h429fc65e};
test_index[2567] = '{7};
test_input[20544:20551] = '{32'h42aa9d6c, 32'hc222bb26, 32'h4197f705, 32'hc25ee8c9, 32'h41dc93da, 32'hc0d0babe, 32'h42022f7f, 32'h42af2225};
test_output[2568] = '{32'h42af2225};
test_index[2568] = '{7};
test_input[20552:20559] = '{32'hc01e9bbc, 32'hc24b2fa5, 32'hc1e44976, 32'hc1005f69, 32'h41b02338, 32'h3d7acda2, 32'hc27bb7f9, 32'hc2c34526};
test_output[2569] = '{32'h41b02338};
test_index[2569] = '{4};
test_input[20560:20567] = '{32'hc29d6e26, 32'h41c5e361, 32'h42210043, 32'hc261ed6e, 32'h42848ebd, 32'hc244b020, 32'hc261c87a, 32'hc2183a71};
test_output[2570] = '{32'h42848ebd};
test_index[2570] = '{4};
test_input[20568:20575] = '{32'h4224550a, 32'hc15883d3, 32'hc2484f6a, 32'hc27b21fb, 32'hc286d7aa, 32'hc239d2b6, 32'h41cdb1a7, 32'hc25159bb};
test_output[2571] = '{32'h4224550a};
test_index[2571] = '{0};
test_input[20576:20583] = '{32'h42ad695b, 32'h42ae5528, 32'hc0a8fd11, 32'h41ebc8fa, 32'h41a4a78f, 32'h42ba272f, 32'h419294cd, 32'h41b3cf7d};
test_output[2572] = '{32'h42ba272f};
test_index[2572] = '{5};
test_input[20584:20591] = '{32'h427bb472, 32'hc2b42ab7, 32'hc0442615, 32'hc22a2595, 32'hc20f7cf0, 32'h428fbda2, 32'h4214c70e, 32'hc220ba3c};
test_output[2573] = '{32'h428fbda2};
test_index[2573] = '{5};
test_input[20592:20599] = '{32'hc02c95b4, 32'h4292e239, 32'hc2c1228a, 32'h42863d3c, 32'hc24e476c, 32'h42b536ed, 32'h424a489a, 32'h4115bbec};
test_output[2574] = '{32'h42b536ed};
test_index[2574] = '{5};
test_input[20600:20607] = '{32'hc1e45091, 32'h42210419, 32'h412bd083, 32'h41708bc1, 32'h42bf5e7b, 32'h424beef6, 32'hc2b61bcb, 32'h4225ee2a};
test_output[2575] = '{32'h42bf5e7b};
test_index[2575] = '{4};
test_input[20608:20615] = '{32'hc2924e73, 32'h41975c0c, 32'h42a2bdaf, 32'hc0eb1278, 32'h41e00939, 32'hc298b41c, 32'hc266b8c5, 32'h4248c29c};
test_output[2576] = '{32'h42a2bdaf};
test_index[2576] = '{2};
test_input[20616:20623] = '{32'h42a3b9fe, 32'hc2a8abb0, 32'h42a64b20, 32'h42295cb8, 32'h41f8ed33, 32'h410b1119, 32'hc281f515, 32'hc19fc3dc};
test_output[2577] = '{32'h42a64b20};
test_index[2577] = '{2};
test_input[20624:20631] = '{32'hc1825d96, 32'h4222fd73, 32'hc2a32c20, 32'hc2bcd5df, 32'h4024c4eb, 32'h42964c34, 32'h42a61a2b, 32'h42c19de0};
test_output[2578] = '{32'h42c19de0};
test_index[2578] = '{7};
test_input[20632:20639] = '{32'hc1498929, 32'hc23f554d, 32'hc249f147, 32'hc294ba37, 32'hc0527f43, 32'h41ebab4e, 32'hc2953664, 32'hc2472897};
test_output[2579] = '{32'h41ebab4e};
test_index[2579] = '{5};
test_input[20640:20647] = '{32'hc28daa90, 32'hc26e73b0, 32'hc1f2540f, 32'h41e988b6, 32'h42a228c0, 32'h4245c484, 32'h424d44f6, 32'hc0a3692d};
test_output[2580] = '{32'h42a228c0};
test_index[2580] = '{4};
test_input[20648:20655] = '{32'h4269dc4e, 32'hc2b82ffe, 32'h42c46f34, 32'h4204cf58, 32'h42784ea8, 32'hc1013704, 32'hc2480404, 32'h4134e478};
test_output[2581] = '{32'h42c46f34};
test_index[2581] = '{2};
test_input[20656:20663] = '{32'h3f26f109, 32'h42688f21, 32'hc2735a1b, 32'hc2aa385c, 32'h42bf3fd1, 32'hc25e6c14, 32'hc28300b8, 32'hc1663526};
test_output[2582] = '{32'h42bf3fd1};
test_index[2582] = '{4};
test_input[20664:20671] = '{32'hc208b19f, 32'h4160b3de, 32'h425fa24a, 32'hc2c76b1b, 32'hc1f542a5, 32'h3f3fc443, 32'h41f818dd, 32'h420ac2d7};
test_output[2583] = '{32'h425fa24a};
test_index[2583] = '{2};
test_input[20672:20679] = '{32'hc261cbcf, 32'h41fb90c6, 32'hc2bae410, 32'hc293e12a, 32'hc1cd64d9, 32'hc16d8340, 32'hc0f59cc5, 32'hc18c05ba};
test_output[2584] = '{32'h41fb90c6};
test_index[2584] = '{1};
test_input[20680:20687] = '{32'h426432d3, 32'hc29250df, 32'h42114aaa, 32'hc1e24f94, 32'h418db0ea, 32'h4258dcc6, 32'hc28ee414, 32'h426d5d29};
test_output[2585] = '{32'h426d5d29};
test_index[2585] = '{7};
test_input[20688:20695] = '{32'h4235c4a2, 32'hc2482e5b, 32'h42196244, 32'h42b181de, 32'hc202719f, 32'h4295b93e, 32'h41c6d0b0, 32'hc23c40d7};
test_output[2586] = '{32'h42b181de};
test_index[2586] = '{3};
test_input[20696:20703] = '{32'hc25ca860, 32'hc24d4986, 32'h42c67a1a, 32'h4267df67, 32'hc2726978, 32'hc276a9f9, 32'h40c94c68, 32'h41b94aa8};
test_output[2587] = '{32'h42c67a1a};
test_index[2587] = '{2};
test_input[20704:20711] = '{32'hc28170f0, 32'h42bc6e89, 32'h4207a4a1, 32'h42aee172, 32'hc2ae1748, 32'h42825b4c, 32'hc2b06a5c, 32'hc2c353f0};
test_output[2588] = '{32'h42bc6e89};
test_index[2588] = '{1};
test_input[20712:20719] = '{32'h41811edc, 32'hc2bcbc43, 32'h414c1ef0, 32'h424b5fa7, 32'hc2170cfd, 32'hc28b16a2, 32'h41739f8e, 32'hc2539638};
test_output[2589] = '{32'h424b5fa7};
test_index[2589] = '{3};
test_input[20720:20727] = '{32'hbfdd80b9, 32'hc1f50d01, 32'h42ac4663, 32'h427a95d8, 32'hc1be31bd, 32'hc1aa485d, 32'hc2a1196a, 32'h42a1838d};
test_output[2590] = '{32'h42ac4663};
test_index[2590] = '{2};
test_input[20728:20735] = '{32'h42b5a28f, 32'hc2362c3d, 32'h42b54384, 32'hc2bafbd9, 32'hc0e1ad2f, 32'h42a3e77f, 32'hc2798724, 32'h42bed7b3};
test_output[2591] = '{32'h42bed7b3};
test_index[2591] = '{7};
test_input[20736:20743] = '{32'h41d01f80, 32'h41ad4e03, 32'h42b3b00a, 32'hc1806fc5, 32'h427aedff, 32'hc2148c70, 32'hc234a0f6, 32'hc22ec4f6};
test_output[2592] = '{32'h42b3b00a};
test_index[2592] = '{2};
test_input[20744:20751] = '{32'h408167d2, 32'hc2216f34, 32'hc25f47ab, 32'h42c625f1, 32'hc26d1541, 32'h42402131, 32'hc2901252, 32'h42b33890};
test_output[2593] = '{32'h42c625f1};
test_index[2593] = '{3};
test_input[20752:20759] = '{32'hc2537ee0, 32'hc2040afe, 32'h42a78306, 32'hc21bc176, 32'hc2bb95e5, 32'h4273732a, 32'h41b75437, 32'h42712dfc};
test_output[2594] = '{32'h42a78306};
test_index[2594] = '{2};
test_input[20760:20767] = '{32'hc219e168, 32'h42748282, 32'h415a46e8, 32'h42c16c4f, 32'h42b54643, 32'h423539f3, 32'hc252a122, 32'h42168f81};
test_output[2595] = '{32'h42c16c4f};
test_index[2595] = '{3};
test_input[20768:20775] = '{32'h41ca7dab, 32'hc2932fbe, 32'h40e60eab, 32'hc11c5731, 32'hc28af15d, 32'h4153a35f, 32'hc1ca126a, 32'h41cfac67};
test_output[2596] = '{32'h41cfac67};
test_index[2596] = '{7};
test_input[20776:20783] = '{32'h427d1346, 32'h4200f7c8, 32'hc23b0a73, 32'hc1b57339, 32'h3fa0673f, 32'h423021d9, 32'hc206e505, 32'h424c5c3c};
test_output[2597] = '{32'h427d1346};
test_index[2597] = '{0};
test_input[20784:20791] = '{32'hc09718b3, 32'hc1acd835, 32'h426e62df, 32'hc1c6f9cb, 32'hc26d6db4, 32'h425e400a, 32'hc2771766, 32'h429c5a91};
test_output[2598] = '{32'h429c5a91};
test_index[2598] = '{7};
test_input[20792:20799] = '{32'hc2840951, 32'hc0d8d6f2, 32'hc16e985b, 32'h40c89d9e, 32'hc299f772, 32'h42b04366, 32'h42a3b24a, 32'h42293168};
test_output[2599] = '{32'h42b04366};
test_index[2599] = '{5};
test_input[20800:20807] = '{32'h4275d0cb, 32'h4263ecf6, 32'hc284855b, 32'hc23948b6, 32'h42237ebf, 32'h425d5090, 32'h425ead86, 32'h41ba51d1};
test_output[2600] = '{32'h4275d0cb};
test_index[2600] = '{0};
test_input[20808:20815] = '{32'h427ea264, 32'hc1d13496, 32'h42b5d9b5, 32'h42982895, 32'h425f920c, 32'hc22f6e03, 32'hc15f8af1, 32'hc144cf4c};
test_output[2601] = '{32'h42b5d9b5};
test_index[2601] = '{2};
test_input[20816:20823] = '{32'hc2a79ca5, 32'hbffc0cd6, 32'h41afca2a, 32'hc0079c47, 32'h4103a54f, 32'h425328dc, 32'h41c57d4c, 32'h42369d2f};
test_output[2602] = '{32'h425328dc};
test_index[2602] = '{5};
test_input[20824:20831] = '{32'hc27a2c92, 32'hc23068e2, 32'h4110ad8f, 32'h42339116, 32'hc2580cb5, 32'h41ff9973, 32'hbfce0073, 32'h4217b616};
test_output[2603] = '{32'h42339116};
test_index[2603] = '{3};
test_input[20832:20839] = '{32'h423c12e1, 32'h4201bdc9, 32'h425a5274, 32'h422411ba, 32'h420098c4, 32'hc2844d71, 32'hc22615c4, 32'hc281d0e2};
test_output[2604] = '{32'h425a5274};
test_index[2604] = '{2};
test_input[20840:20847] = '{32'hc246410e, 32'hc028e328, 32'hc21fa3e5, 32'hc293e4f1, 32'hc1b2cdb1, 32'h418f9662, 32'hc2897484, 32'hc225738c};
test_output[2605] = '{32'h418f9662};
test_index[2605] = '{5};
test_input[20848:20855] = '{32'hc2a8d3c2, 32'hc2bc6d58, 32'hc26ac56a, 32'h40da10ec, 32'hc23c3313, 32'hc2a6a382, 32'h429aece2, 32'hc28280e3};
test_output[2606] = '{32'h429aece2};
test_index[2606] = '{6};
test_input[20856:20863] = '{32'h41c112cd, 32'hc0966e4e, 32'h408b9c68, 32'h42738d78, 32'hc2b70913, 32'h42b8a9c5, 32'hc2626908, 32'hc082e33a};
test_output[2607] = '{32'h42b8a9c5};
test_index[2607] = '{5};
test_input[20864:20871] = '{32'hc1ee9b97, 32'h421ebdfb, 32'h41a9e7c7, 32'hc1ecf6b3, 32'hc2b58bb4, 32'h428fec93, 32'hc21c9dbe, 32'h41817729};
test_output[2608] = '{32'h428fec93};
test_index[2608] = '{5};
test_input[20872:20879] = '{32'hc1f74cd5, 32'h42a11f44, 32'h428be63a, 32'h420da457, 32'h42270615, 32'h428feb9a, 32'h42c45a5f, 32'hc26739e0};
test_output[2609] = '{32'h42c45a5f};
test_index[2609] = '{6};
test_input[20880:20887] = '{32'hc26ed0e9, 32'h4253594b, 32'hc1d0579b, 32'h41943a61, 32'hc2b603aa, 32'h4277b814, 32'hc2687a5b, 32'h4293f184};
test_output[2610] = '{32'h4293f184};
test_index[2610] = '{7};
test_input[20888:20895] = '{32'hc1e0421b, 32'hc2aa680f, 32'hc0965a22, 32'h42a9e689, 32'h41d6d5d1, 32'hc29a64da, 32'hc234a652, 32'hc299ad01};
test_output[2611] = '{32'h42a9e689};
test_index[2611] = '{3};
test_input[20896:20903] = '{32'hc2750964, 32'h419b923d, 32'h40cfc462, 32'h4242fc28, 32'hc1782cd4, 32'h424430fd, 32'hc1c3cd94, 32'hc28d6ca7};
test_output[2612] = '{32'h424430fd};
test_index[2612] = '{5};
test_input[20904:20911] = '{32'h422fff67, 32'hc2a1451d, 32'hc284ada3, 32'hc2aa4252, 32'hc2240480, 32'hc2b7d2e2, 32'hc26f1508, 32'h41b19a81};
test_output[2613] = '{32'h422fff67};
test_index[2613] = '{0};
test_input[20912:20919] = '{32'hc1dd55f8, 32'hc2b281db, 32'h429cf4fe, 32'hc20afdda, 32'hc1f0cd02, 32'h426435ff, 32'hc2288543, 32'hc29eb96c};
test_output[2614] = '{32'h429cf4fe};
test_index[2614] = '{2};
test_input[20920:20927] = '{32'hc0c64e04, 32'hc299276f, 32'hc2141453, 32'hc26556a7, 32'h428eccaf, 32'h4209d82a, 32'h422b7ed7, 32'h41e9d39c};
test_output[2615] = '{32'h428eccaf};
test_index[2615] = '{4};
test_input[20928:20935] = '{32'hc1c18e1d, 32'hc2b637f6, 32'h40f9c525, 32'h423ec640, 32'h4207324e, 32'h41eae792, 32'h42b2aaf2, 32'hc2af6ff0};
test_output[2616] = '{32'h42b2aaf2};
test_index[2616] = '{6};
test_input[20936:20943] = '{32'hc2a16069, 32'hc2885fff, 32'h4204a898, 32'h4211efc6, 32'hc170bb51, 32'h41eb460f, 32'h42942e14, 32'h429ed0e3};
test_output[2617] = '{32'h429ed0e3};
test_index[2617] = '{7};
test_input[20944:20951] = '{32'hc208ad3d, 32'hc249769b, 32'h42bed003, 32'h41e63956, 32'hc2977de2, 32'hc1c6d149, 32'hc15c7740, 32'hc29e599d};
test_output[2618] = '{32'h42bed003};
test_index[2618] = '{2};
test_input[20952:20959] = '{32'h420c3c01, 32'hc2853aca, 32'h42b40fd5, 32'hc20b5e85, 32'hc2634e3b, 32'h41d7cf36, 32'h42071f2c, 32'h4222495f};
test_output[2619] = '{32'h42b40fd5};
test_index[2619] = '{2};
test_input[20960:20967] = '{32'hc280d373, 32'hc255de19, 32'h41f56287, 32'hc1d2d638, 32'hc1a92866, 32'h4105f42c, 32'hc22166ce, 32'hc2c626e9};
test_output[2620] = '{32'h41f56287};
test_index[2620] = '{2};
test_input[20968:20975] = '{32'h41949383, 32'hc158353c, 32'h4287b9d2, 32'h42a5e180, 32'hc2639767, 32'h41f61a6c, 32'hc1cdb627, 32'hbf66aa29};
test_output[2621] = '{32'h42a5e180};
test_index[2621] = '{3};
test_input[20976:20983] = '{32'hc2ba1484, 32'hc2a65e5f, 32'h4266ea4d, 32'h412f308b, 32'h420ea582, 32'h423585d2, 32'h42adc0ea, 32'hc2118817};
test_output[2622] = '{32'h42adc0ea};
test_index[2622] = '{6};
test_input[20984:20991] = '{32'h3f4aaa29, 32'hc0e38805, 32'hc2797bbc, 32'hc2823c4f, 32'hc0b2efcd, 32'hc1d12688, 32'h4283b0f2, 32'h41575c96};
test_output[2623] = '{32'h4283b0f2};
test_index[2623] = '{6};
test_input[20992:20999] = '{32'h4296b0c4, 32'hc2bfd10b, 32'h42211826, 32'hc27748eb, 32'h41a61596, 32'hc2c476b3, 32'h42873a5f, 32'h41a60cf6};
test_output[2624] = '{32'h4296b0c4};
test_index[2624] = '{0};
test_input[21000:21007] = '{32'h428f484b, 32'hc2552247, 32'hc28d5e5e, 32'hc2c2e770, 32'hc2901428, 32'hc09b80eb, 32'hc1f2f92a, 32'hc08a72bb};
test_output[2625] = '{32'h428f484b};
test_index[2625] = '{0};
test_input[21008:21015] = '{32'h4112d542, 32'h3f09c2f2, 32'h4065d791, 32'hc2093414, 32'h42c1264e, 32'h41704760, 32'hc2a65e19, 32'h42239e21};
test_output[2626] = '{32'h42c1264e};
test_index[2626] = '{4};
test_input[21016:21023] = '{32'hc2686dbd, 32'hc1b7c316, 32'hc213b2ed, 32'h41a7049c, 32'hc2c0e5bc, 32'hc27a05fb, 32'hc284d927, 32'h428a1b30};
test_output[2627] = '{32'h428a1b30};
test_index[2627] = '{7};
test_input[21024:21031] = '{32'hc2a279c5, 32'h42839f76, 32'h4244f568, 32'h42099ef7, 32'hc12ddb6f, 32'hc1abf6c1, 32'h4253e30e, 32'hc23785e6};
test_output[2628] = '{32'h42839f76};
test_index[2628] = '{1};
test_input[21032:21039] = '{32'hc1651f02, 32'h4209de72, 32'h420f49b6, 32'hc19e758a, 32'hc2adab4f, 32'h42940da3, 32'h41770eb2, 32'hc2bc4c87};
test_output[2629] = '{32'h42940da3};
test_index[2629] = '{5};
test_input[21040:21047] = '{32'hc118385b, 32'h4298ec11, 32'hc2ae2001, 32'hc10e4b9b, 32'hc219e83a, 32'hc2779755, 32'h42a7bc2b, 32'h421ff7b0};
test_output[2630] = '{32'h42a7bc2b};
test_index[2630] = '{6};
test_input[21048:21055] = '{32'h42c66235, 32'hc2a50298, 32'h42a7773b, 32'hc2a2b58a, 32'h42369ef7, 32'hc2a160c9, 32'hc2093b69, 32'h41ce6eb3};
test_output[2631] = '{32'h42c66235};
test_index[2631] = '{0};
test_input[21056:21063] = '{32'hc2b9b9dd, 32'hc25a68a7, 32'h424b4eb3, 32'h42c460ab, 32'h423f0ed0, 32'h428efd74, 32'h41e49ee9, 32'hc22787fe};
test_output[2632] = '{32'h42c460ab};
test_index[2632] = '{3};
test_input[21064:21071] = '{32'h427e8c36, 32'hc1b3ad0a, 32'hc29f969d, 32'h42353404, 32'h3f0eb66f, 32'h3fc0d954, 32'hc2838065, 32'hc20dd40e};
test_output[2633] = '{32'h427e8c36};
test_index[2633] = '{0};
test_input[21072:21079] = '{32'h41469b62, 32'h41cc0f28, 32'hc2c33bde, 32'hc09deefc, 32'h41c99166, 32'h4176901e, 32'hc2a1b405, 32'h42b9f2e4};
test_output[2634] = '{32'h42b9f2e4};
test_index[2634] = '{7};
test_input[21080:21087] = '{32'hc0aea3b8, 32'hc2bfefb2, 32'h42b5eead, 32'h41f9aa38, 32'h421bc4f3, 32'hc1f51587, 32'hc2b595c1, 32'h42a854a8};
test_output[2635] = '{32'h42b5eead};
test_index[2635] = '{2};
test_input[21088:21095] = '{32'hc29e0f63, 32'hc0937161, 32'h428b207b, 32'hc28889fd, 32'h41cbb4be, 32'h42c421e9, 32'hc2789ba0, 32'hc2568497};
test_output[2636] = '{32'h42c421e9};
test_index[2636] = '{5};
test_input[21096:21103] = '{32'hc038e588, 32'hc2b99ba5, 32'hc18235c9, 32'h42ab298c, 32'h423e4f67, 32'h425efe1e, 32'hc2975f27, 32'h40c8ac3e};
test_output[2637] = '{32'h42ab298c};
test_index[2637] = '{3};
test_input[21104:21111] = '{32'h42296eb4, 32'hc1c03e5f, 32'hc234b386, 32'h41c70aa4, 32'h42533873, 32'h40d294c3, 32'h42641513, 32'h429dd139};
test_output[2638] = '{32'h429dd139};
test_index[2638] = '{7};
test_input[21112:21119] = '{32'h41ab2864, 32'h41ddab73, 32'h427f3085, 32'hc2384826, 32'h42b4e413, 32'hc265fc39, 32'h42c2f0b6, 32'hc242b213};
test_output[2639] = '{32'h42c2f0b6};
test_index[2639] = '{6};
test_input[21120:21127] = '{32'h42b5ce0a, 32'h42b90aef, 32'hc197386f, 32'hbff099f4, 32'h3ec4017c, 32'hc181262a, 32'h428e161b, 32'hc2908423};
test_output[2640] = '{32'h42b90aef};
test_index[2640] = '{1};
test_input[21128:21135] = '{32'h425f56e1, 32'hc2ace41c, 32'h42822711, 32'hc08ae175, 32'hc11641cc, 32'hc29d3a93, 32'h424aeb68, 32'h42be1631};
test_output[2641] = '{32'h42be1631};
test_index[2641] = '{7};
test_input[21136:21143] = '{32'hc16b4f20, 32'hc18b5e62, 32'hc28bb289, 32'hc05b492f, 32'hc1b3512c, 32'h42373a60, 32'hc2338c8f, 32'h42bb8728};
test_output[2642] = '{32'h42bb8728};
test_index[2642] = '{7};
test_input[21144:21151] = '{32'hc1a2b7a0, 32'h41d45b4a, 32'hc1ba6d43, 32'hc2b0b889, 32'h423839c8, 32'hc2bb6048, 32'hc28973b4, 32'h421d13ea};
test_output[2643] = '{32'h423839c8};
test_index[2643] = '{4};
test_input[21152:21159] = '{32'h42c6d697, 32'hc2868389, 32'hc2c48e11, 32'h412690dd, 32'h42a01e50, 32'hc2061a4a, 32'hc295b46e, 32'h428ef92d};
test_output[2644] = '{32'h42c6d697};
test_index[2644] = '{0};
test_input[21160:21167] = '{32'hc1276be7, 32'hc20e1052, 32'hc19453ab, 32'h4298bab3, 32'h42b99b1e, 32'hc2a842e9, 32'hc227f500, 32'hc1e0a5df};
test_output[2645] = '{32'h42b99b1e};
test_index[2645] = '{4};
test_input[21168:21175] = '{32'hc27d36de, 32'h4203df6f, 32'h420cbb02, 32'h42534d72, 32'hc2982e89, 32'hc2a8a027, 32'h42a65e58, 32'h420e62dc};
test_output[2646] = '{32'h42a65e58};
test_index[2646] = '{6};
test_input[21176:21183] = '{32'h42301878, 32'h40bc7916, 32'h41c330a9, 32'h4228a2c1, 32'h40e00ca1, 32'h42c590f6, 32'hc2b6a010, 32'h42a40292};
test_output[2647] = '{32'h42c590f6};
test_index[2647] = '{5};
test_input[21184:21191] = '{32'hc09cffd1, 32'h42c0c6c7, 32'h42b40487, 32'h41992983, 32'hc203517d, 32'h423cac0d, 32'h42bb3ef9, 32'h418d4d56};
test_output[2648] = '{32'h42c0c6c7};
test_index[2648] = '{1};
test_input[21192:21199] = '{32'hc2014fcd, 32'hc2022bec, 32'hc27ab08e, 32'h40ee3b23, 32'hc2ad65c0, 32'h422d87b0, 32'hc2a9d591, 32'hc254022e};
test_output[2649] = '{32'h422d87b0};
test_index[2649] = '{5};
test_input[21200:21207] = '{32'hc169d1b2, 32'hc2577482, 32'h4197aa8b, 32'h42b665c1, 32'hc25a8fb3, 32'hc173b22c, 32'h41b5588c, 32'h41e97bd4};
test_output[2650] = '{32'h42b665c1};
test_index[2650] = '{3};
test_input[21208:21215] = '{32'h427020f9, 32'h40fb4472, 32'h42249b1a, 32'h3fc877d1, 32'h421f26c3, 32'hc2304a7a, 32'h403a0e8d, 32'hc1d2d8dc};
test_output[2651] = '{32'h427020f9};
test_index[2651] = '{0};
test_input[21216:21223] = '{32'hc16eb03c, 32'h414baf29, 32'hc2423420, 32'h421fe4de, 32'hc28f89ef, 32'h42914079, 32'hc2008958, 32'hc19a97a2};
test_output[2652] = '{32'h42914079};
test_index[2652] = '{5};
test_input[21224:21231] = '{32'hc257dc38, 32'hc15e04dd, 32'hc2459da6, 32'hc1bc5e54, 32'h41dc20b1, 32'hc21536d2, 32'h42b4716d, 32'hc298b4ae};
test_output[2653] = '{32'h42b4716d};
test_index[2653] = '{6};
test_input[21232:21239] = '{32'h4209a3ba, 32'h410cf053, 32'h428998a9, 32'h4230fef3, 32'h423699a7, 32'hc2b4b138, 32'hc1efa0a2, 32'hc1a9e955};
test_output[2654] = '{32'h428998a9};
test_index[2654] = '{2};
test_input[21240:21247] = '{32'h4292b22f, 32'hc2ac8621, 32'h42175bfd, 32'h41a5874a, 32'hc28ed46a, 32'hbfd8413e, 32'hc2290b0b, 32'h4187b039};
test_output[2655] = '{32'h4292b22f};
test_index[2655] = '{0};
test_input[21248:21255] = '{32'h429f52f9, 32'h429360ba, 32'hc2bc58f4, 32'hc2807c8b, 32'h42a68c31, 32'h4251c50e, 32'h426eebfc, 32'hc00b5614};
test_output[2656] = '{32'h42a68c31};
test_index[2656] = '{4};
test_input[21256:21263] = '{32'hc2807d0f, 32'h41dc1a3a, 32'hc21b6f94, 32'h4282f4f7, 32'hc19a17d4, 32'hc265d91e, 32'hc24f2fe3, 32'hc21667d3};
test_output[2657] = '{32'h4282f4f7};
test_index[2657] = '{3};
test_input[21264:21271] = '{32'h42bd6acb, 32'h42b86c0a, 32'hc1e09982, 32'h42c3d142, 32'hc24585ac, 32'h41258d44, 32'hc2ad915b, 32'h42af087a};
test_output[2658] = '{32'h42c3d142};
test_index[2658] = '{3};
test_input[21272:21279] = '{32'hc2679c43, 32'h4281d330, 32'h4214c697, 32'h42b3f835, 32'h419af959, 32'hc1b5f20c, 32'hc1dccff9, 32'hc29ecc3d};
test_output[2659] = '{32'h42b3f835};
test_index[2659] = '{3};
test_input[21280:21287] = '{32'h418bf3c3, 32'hc2b1f42c, 32'h42c3153e, 32'hc29e6627, 32'h42c2ccc9, 32'h429f7a67, 32'hc2b70359, 32'h4228acfd};
test_output[2660] = '{32'h42c3153e};
test_index[2660] = '{2};
test_input[21288:21295] = '{32'h41f75d20, 32'h42a01ba1, 32'h422e77d5, 32'h420231ed, 32'hc1b065f8, 32'h40ea83c6, 32'hc2966249, 32'h42a30ea2};
test_output[2661] = '{32'h42a30ea2};
test_index[2661] = '{7};
test_input[21296:21303] = '{32'h40771bee, 32'h4252fbe3, 32'h42b00008, 32'h42932af6, 32'hc26b3776, 32'h4275e515, 32'hc275a14a, 32'hc263a600};
test_output[2662] = '{32'h42b00008};
test_index[2662] = '{2};
test_input[21304:21311] = '{32'hc1fc17d0, 32'h428955bb, 32'h422fa6c9, 32'hc265cfc4, 32'h4273b9ea, 32'hc183f4e8, 32'h42b7f29c, 32'h41bb501a};
test_output[2663] = '{32'h42b7f29c};
test_index[2663] = '{6};
test_input[21312:21319] = '{32'h414b80a8, 32'h4246baea, 32'hc2579362, 32'hc1726ba9, 32'h4228f135, 32'hc1c42001, 32'h41cce8fd, 32'hc2817fe1};
test_output[2664] = '{32'h4246baea};
test_index[2664] = '{1};
test_input[21320:21327] = '{32'hc19fd2ec, 32'h42988e81, 32'hc2a00d7c, 32'hc2989d4f, 32'h42953e42, 32'hc214f22f, 32'hc2c3545f, 32'hc2525139};
test_output[2665] = '{32'h42988e81};
test_index[2665] = '{1};
test_input[21328:21335] = '{32'hc25ec55f, 32'hc2316fb1, 32'h4283b890, 32'hc0c6ef3a, 32'hc213b433, 32'h4276777f, 32'hc1a94af3, 32'hc22f8ffa};
test_output[2666] = '{32'h4283b890};
test_index[2666] = '{2};
test_input[21336:21343] = '{32'hc23825de, 32'hc26e3c81, 32'hc18fc4ba, 32'h414d93de, 32'hc24c6278, 32'hc2266ec6, 32'hc2a47629, 32'hc22bdba2};
test_output[2667] = '{32'h414d93de};
test_index[2667] = '{3};
test_input[21344:21351] = '{32'hc1fc1a1e, 32'h4184f979, 32'hc12f86ed, 32'h42680796, 32'h4188b0fa, 32'hc2125729, 32'h40cf31a6, 32'hc11c043e};
test_output[2668] = '{32'h42680796};
test_index[2668] = '{3};
test_input[21352:21359] = '{32'h4280ce16, 32'h4161ada0, 32'h428c9c0b, 32'hc20ffcd6, 32'hc217512b, 32'h41964714, 32'h429507fb, 32'h423d64d1};
test_output[2669] = '{32'h429507fb};
test_index[2669] = '{6};
test_input[21360:21367] = '{32'hc27b983b, 32'h4277d442, 32'h40f8e6c6, 32'h42c227c0, 32'h40a2e816, 32'h419c8aa4, 32'hc29cecd4, 32'hc1d032b5};
test_output[2670] = '{32'h42c227c0};
test_index[2670] = '{3};
test_input[21368:21375] = '{32'h4260265c, 32'h41929b95, 32'h4103262e, 32'hc212de0f, 32'hc1b996c1, 32'hc1793c17, 32'hc165e56e, 32'hc2b9b83e};
test_output[2671] = '{32'h4260265c};
test_index[2671] = '{0};
test_input[21376:21383] = '{32'h4195715d, 32'h42853eeb, 32'hc2c4d0e6, 32'h41d140d9, 32'hc211c5eb, 32'hc2c2f5d3, 32'hc0e5d03b, 32'hc218471b};
test_output[2672] = '{32'h42853eeb};
test_index[2672] = '{1};
test_input[21384:21391] = '{32'h429009b9, 32'h42116509, 32'hc2ac0421, 32'h41cfe910, 32'hc2a2396c, 32'h4280c342, 32'h4257aa4a, 32'hc04cb6a2};
test_output[2673] = '{32'h429009b9};
test_index[2673] = '{0};
test_input[21392:21399] = '{32'h41dbd663, 32'hc12f0ee0, 32'hc2673494, 32'hc1d4f4d6, 32'hc216e60e, 32'h42a90a7e, 32'h4130501e, 32'hc204413a};
test_output[2674] = '{32'h42a90a7e};
test_index[2674] = '{5};
test_input[21400:21407] = '{32'hc1a3f0e0, 32'h428b06f0, 32'h42a5d427, 32'h42a1b93e, 32'hc20f7f36, 32'h427ebb78, 32'h4181af91, 32'hc2c5e733};
test_output[2675] = '{32'h42a5d427};
test_index[2675] = '{2};
test_input[21408:21415] = '{32'h41907551, 32'h428dc9a7, 32'h41daaacc, 32'hc29bc4b6, 32'hc2123f33, 32'hc24cba3a, 32'hc2c0b8e5, 32'h424febb4};
test_output[2676] = '{32'h428dc9a7};
test_index[2676] = '{1};
test_input[21416:21423] = '{32'hc28e61f1, 32'h42b0c32e, 32'hc2221a26, 32'h4257e4bf, 32'hc2bf87b9, 32'h42458b15, 32'hc2be2be9, 32'hc2a22d09};
test_output[2677] = '{32'h42b0c32e};
test_index[2677] = '{1};
test_input[21424:21431] = '{32'h3fb125fd, 32'hc255edd4, 32'h429376d2, 32'h41f41113, 32'hc2bcf53c, 32'h4262aa07, 32'hc2bc6095, 32'hc1ebe5ee};
test_output[2678] = '{32'h429376d2};
test_index[2678] = '{2};
test_input[21432:21439] = '{32'hc28bec71, 32'h418d8405, 32'h42b00b53, 32'h40d6de1d, 32'hc2ae3888, 32'hc1cfcb1f, 32'hc0e1fd84, 32'h4178e327};
test_output[2679] = '{32'h42b00b53};
test_index[2679] = '{2};
test_input[21440:21447] = '{32'h42658d95, 32'h42916730, 32'hc08ae1bd, 32'h41e9fca6, 32'hc28cc37f, 32'hc2361f2a, 32'hc19d237b, 32'h4207a22e};
test_output[2680] = '{32'h42916730};
test_index[2680] = '{1};
test_input[21448:21455] = '{32'h41f32b7c, 32'h41eb2610, 32'hc1d10880, 32'h4211ef95, 32'hc2a14ae4, 32'hc2008f2d, 32'h4292109b, 32'h42a030f0};
test_output[2681] = '{32'h42a030f0};
test_index[2681] = '{7};
test_input[21456:21463] = '{32'hc29317e3, 32'h4298bb71, 32'hc1645787, 32'hc23dbb52, 32'h428d2920, 32'hc219b6f7, 32'h42c33e62, 32'hc28c501e};
test_output[2682] = '{32'h42c33e62};
test_index[2682] = '{6};
test_input[21464:21471] = '{32'hc12de6df, 32'hc2a1d1b6, 32'hc2b71a1a, 32'hc24f98ef, 32'hc28a5f32, 32'hc21b0d29, 32'hc0b6c695, 32'h42c0738f};
test_output[2683] = '{32'h42c0738f};
test_index[2683] = '{7};
test_input[21472:21479] = '{32'hc1d6ee4f, 32'hc28ee3f6, 32'h41bf81fc, 32'hc2ae7bfa, 32'h422352f4, 32'hc200bcfd, 32'h428c5acc, 32'hc2b6e54e};
test_output[2684] = '{32'h428c5acc};
test_index[2684] = '{6};
test_input[21480:21487] = '{32'h42a51728, 32'hc0b8994f, 32'hc2c1476d, 32'hc285baf3, 32'h4283a7da, 32'hc2ac741a, 32'hc2b318d8, 32'h3f5e768c};
test_output[2685] = '{32'h42a51728};
test_index[2685] = '{0};
test_input[21488:21495] = '{32'h429d6c45, 32'hc2bb9a48, 32'h429f3787, 32'hc26ee1ac, 32'hc281e8ae, 32'hc2af673b, 32'hc18cfac3, 32'hc2b1050d};
test_output[2686] = '{32'h429f3787};
test_index[2686] = '{2};
test_input[21496:21503] = '{32'h42b0dd71, 32'h3fa48071, 32'h414c5b26, 32'h42631f6f, 32'hc1e7b4bd, 32'h4283d46a, 32'hc216c2da, 32'h428357b8};
test_output[2687] = '{32'h42b0dd71};
test_index[2687] = '{0};
test_input[21504:21511] = '{32'h4291dc66, 32'h42469ab1, 32'hc20e1d2b, 32'h42c24947, 32'h41b82f1c, 32'hc26e664b, 32'h42822cbf, 32'hc2a0b764};
test_output[2688] = '{32'h42c24947};
test_index[2688] = '{3};
test_input[21512:21519] = '{32'h4294565e, 32'h4058da9c, 32'h42c34c3b, 32'h427d4c2d, 32'h42016848, 32'hc257f4e9, 32'hc297e95d, 32'h4287846e};
test_output[2689] = '{32'h42c34c3b};
test_index[2689] = '{2};
test_input[21520:21527] = '{32'h405f3943, 32'hc2a7c998, 32'hc2156008, 32'h42821faa, 32'hc2b82aae, 32'hc1667cd9, 32'hc28763f9, 32'hc265f44e};
test_output[2690] = '{32'h42821faa};
test_index[2690] = '{3};
test_input[21528:21535] = '{32'h426e556f, 32'hc29ef97c, 32'hc1c1800a, 32'h4220fce3, 32'h421ec2a6, 32'hc2a6087e, 32'h419bad3a, 32'h3f6937e1};
test_output[2691] = '{32'h426e556f};
test_index[2691] = '{0};
test_input[21536:21543] = '{32'hc2687838, 32'hc1b14791, 32'hc2bb24f0, 32'h4292d89b, 32'h410f90b8, 32'hc2b6cc9d, 32'hc28f86f3, 32'hc2663633};
test_output[2692] = '{32'h4292d89b};
test_index[2692] = '{3};
test_input[21544:21551] = '{32'h42b53bbf, 32'h428a15a5, 32'hc27c4188, 32'hc2c5944d, 32'h423f34f7, 32'h426ffb1f, 32'h40aaf102, 32'hc233273a};
test_output[2693] = '{32'h42b53bbf};
test_index[2693] = '{0};
test_input[21552:21559] = '{32'h42027c90, 32'hc28d7eeb, 32'h418a3076, 32'h42b97e94, 32'hc210da98, 32'hc27f1392, 32'h4146af38, 32'h41fa32ea};
test_output[2694] = '{32'h42b97e94};
test_index[2694] = '{3};
test_input[21560:21567] = '{32'h422956db, 32'h4186d97e, 32'h41d6150e, 32'h41cb50ab, 32'hc1ea4fcc, 32'hc2a694bb, 32'hc2c5919f, 32'hc215d68d};
test_output[2695] = '{32'h422956db};
test_index[2695] = '{0};
test_input[21568:21575] = '{32'h42a3bb82, 32'hc129aba8, 32'h42044f99, 32'h42a62698, 32'h428d8029, 32'hc20338aa, 32'hc19dc5f4, 32'hc1fb3b0a};
test_output[2696] = '{32'h42a62698};
test_index[2696] = '{3};
test_input[21576:21583] = '{32'hc28f0bb2, 32'hc2b00663, 32'hc2791774, 32'hc27cb7b7, 32'h4143f027, 32'hc2acb966, 32'hc182439f, 32'h420c5c87};
test_output[2697] = '{32'h420c5c87};
test_index[2697] = '{7};
test_input[21584:21591] = '{32'hc1c41603, 32'hc2382f88, 32'hc1df9831, 32'hc2a24486, 32'hc279b101, 32'h4175b360, 32'h3d8506d9, 32'h42c639cd};
test_output[2698] = '{32'h42c639cd};
test_index[2698] = '{7};
test_input[21592:21599] = '{32'hc2a5eda8, 32'h4269ed81, 32'h42585039, 32'h428cc828, 32'hc1ec3e95, 32'h4042c3f6, 32'hc1d1f856, 32'h428c0040};
test_output[2699] = '{32'h428cc828};
test_index[2699] = '{3};
test_input[21600:21607] = '{32'hc2b7e3df, 32'hc15976ed, 32'hc2997ae2, 32'h42ab2e72, 32'h42803f21, 32'hc19bc0ed, 32'h42aabcbc, 32'h3e8f2a24};
test_output[2700] = '{32'h42ab2e72};
test_index[2700] = '{3};
test_input[21608:21615] = '{32'hc1a6d484, 32'hc1818442, 32'h40176fb5, 32'h40d969f2, 32'hc192981f, 32'h41802702, 32'h4290b1c7, 32'hc1b9d29c};
test_output[2701] = '{32'h4290b1c7};
test_index[2701] = '{6};
test_input[21616:21623] = '{32'h4227c0af, 32'hc21e2fd7, 32'h41efe0c0, 32'h42156b6b, 32'h42a80db7, 32'h42408bf2, 32'h42a7cd66, 32'hc262e09f};
test_output[2702] = '{32'h42a80db7};
test_index[2702] = '{4};
test_input[21624:21631] = '{32'hc1901d92, 32'hc1b48a5b, 32'h42b7055a, 32'hc29a6edd, 32'hc290c04a, 32'hc2afc500, 32'hbef1fb98, 32'h413a03ba};
test_output[2703] = '{32'h42b7055a};
test_index[2703] = '{2};
test_input[21632:21639] = '{32'hc24518ad, 32'hc15927c7, 32'h42c73cec, 32'hc27ce60f, 32'h421d70b9, 32'hc2109c9c, 32'h41976f00, 32'hc2c4a825};
test_output[2704] = '{32'h42c73cec};
test_index[2704] = '{2};
test_input[21640:21647] = '{32'h4168a486, 32'h42c1e0be, 32'hc20f4343, 32'hc27c7f50, 32'h40ab4c31, 32'hc10ad0eb, 32'h4252c1e2, 32'h41e2aa3e};
test_output[2705] = '{32'h42c1e0be};
test_index[2705] = '{1};
test_input[21648:21655] = '{32'h4206532e, 32'hc2afbf35, 32'hc25aaee0, 32'h418474d5, 32'h428d30a5, 32'hc28a1c74, 32'hc2b3f602, 32'hc260517d};
test_output[2706] = '{32'h428d30a5};
test_index[2706] = '{4};
test_input[21656:21663] = '{32'hc25e4a5c, 32'hc055ab6a, 32'hc24eb22a, 32'h427aa690, 32'hc1b1529d, 32'h4283ec3a, 32'h41df83ca, 32'hc27e593c};
test_output[2707] = '{32'h4283ec3a};
test_index[2707] = '{5};
test_input[21664:21671] = '{32'hc1c0df41, 32'h4229e808, 32'hc283bf87, 32'h42119762, 32'h423d5404, 32'h41dfef25, 32'h422dee76, 32'h429b1193};
test_output[2708] = '{32'h429b1193};
test_index[2708] = '{7};
test_input[21672:21679] = '{32'h42b08bd4, 32'h420bcde1, 32'h42c73dc0, 32'hc1d9a033, 32'hc112e0af, 32'h3d95ac26, 32'hc2b6bd5b, 32'hc26687bc};
test_output[2709] = '{32'h42c73dc0};
test_index[2709] = '{2};
test_input[21680:21687] = '{32'hc2372e3b, 32'hc280ea3c, 32'hc2b370c9, 32'hc0c2a8ec, 32'hc1e97721, 32'h402dab4f, 32'hc1b29947, 32'hc17f76da};
test_output[2710] = '{32'h402dab4f};
test_index[2710] = '{5};
test_input[21688:21695] = '{32'h4253180d, 32'h42c62cc0, 32'h42b3ef61, 32'hc27c93c5, 32'h42490d11, 32'h42c0cab9, 32'h42b9c4e4, 32'h429e94a7};
test_output[2711] = '{32'h42c62cc0};
test_index[2711] = '{1};
test_input[21696:21703] = '{32'h42b037c7, 32'h429cde34, 32'h42b9ced8, 32'hc2a4eba1, 32'hc2ac6b12, 32'hc29a3af4, 32'h4241b664, 32'h42738767};
test_output[2712] = '{32'h42b9ced8};
test_index[2712] = '{2};
test_input[21704:21711] = '{32'h4266058d, 32'h42c4f8bc, 32'hc24b07b3, 32'h42816261, 32'hc289a20f, 32'h420e6a08, 32'hc2c21225, 32'hc2659637};
test_output[2713] = '{32'h42c4f8bc};
test_index[2713] = '{1};
test_input[21712:21719] = '{32'hc2276af0, 32'hc2086766, 32'hc19a9f1f, 32'hc226579b, 32'h3f23bcf1, 32'hc2c2f26f, 32'hbfacc59b, 32'h4153f70c};
test_output[2714] = '{32'h4153f70c};
test_index[2714] = '{7};
test_input[21720:21727] = '{32'h421018b7, 32'h427d5b48, 32'hc29034b2, 32'hc02a9b30, 32'hc28cf17f, 32'h423b9d93, 32'hc1f5f108, 32'hc294c720};
test_output[2715] = '{32'h427d5b48};
test_index[2715] = '{1};
test_input[21728:21735] = '{32'h42279e41, 32'h41832347, 32'hc28f56fe, 32'hc1d645ae, 32'hc22258b9, 32'hc28e5cf5, 32'h4237c602, 32'hc1e2ae32};
test_output[2716] = '{32'h4237c602};
test_index[2716] = '{6};
test_input[21736:21743] = '{32'hc215240c, 32'h40cd6006, 32'hc2b1a358, 32'hc23775c4, 32'h4274d531, 32'h42ba8281, 32'hc2b9936d, 32'h42b7057d};
test_output[2717] = '{32'h42ba8281};
test_index[2717] = '{5};
test_input[21744:21751] = '{32'h422865ee, 32'hc147e6cc, 32'hc294fa91, 32'h42023566, 32'hc1835c2e, 32'h4283959f, 32'hc22dc06e, 32'hc2c19c2c};
test_output[2718] = '{32'h4283959f};
test_index[2718] = '{5};
test_input[21752:21759] = '{32'hc275188b, 32'hc29c7748, 32'h42017d30, 32'hc288919f, 32'hc222e2cb, 32'hc2684857, 32'h42304c75, 32'h42496e8b};
test_output[2719] = '{32'h42496e8b};
test_index[2719] = '{7};
test_input[21760:21767] = '{32'hc2ba30da, 32'h428412eb, 32'hc045c442, 32'h40e03d50, 32'hc2839dda, 32'h41c90e4c, 32'hc0c8188e, 32'hc1d45d40};
test_output[2720] = '{32'h428412eb};
test_index[2720] = '{1};
test_input[21768:21775] = '{32'h4292d0f2, 32'h4208061f, 32'hc0458964, 32'h41fb787c, 32'h421270a8, 32'hc291daf4, 32'h42918796, 32'hc1b81a74};
test_output[2721] = '{32'h4292d0f2};
test_index[2721] = '{0};
test_input[21776:21783] = '{32'h42c5fcbb, 32'h42a7fd76, 32'h426dcdf3, 32'h42a20132, 32'hc27816b3, 32'hc2620d51, 32'h4249ea29, 32'h428b1d2c};
test_output[2722] = '{32'h42c5fcbb};
test_index[2722] = '{0};
test_input[21784:21791] = '{32'h4192a7d7, 32'h4270d7e4, 32'hc273f5cc, 32'hc2848049, 32'h428c492c, 32'h42509eae, 32'h429c720f, 32'hc2b5e304};
test_output[2723] = '{32'h429c720f};
test_index[2723] = '{6};
test_input[21792:21799] = '{32'hc1bb1503, 32'hc197166c, 32'h40573279, 32'h404d879d, 32'h41f99b25, 32'h42c382e4, 32'hc1aff4a3, 32'h4282186a};
test_output[2724] = '{32'h42c382e4};
test_index[2724] = '{5};
test_input[21800:21807] = '{32'hc29f6e96, 32'hc26bd333, 32'h4298abab, 32'h423994c0, 32'hc22c969a, 32'hc20515f9, 32'hc282e8d9, 32'hc1d24926};
test_output[2725] = '{32'h4298abab};
test_index[2725] = '{2};
test_input[21808:21815] = '{32'hc2a33401, 32'hc264dbc8, 32'h42b4f586, 32'h4275fbd8, 32'h420dee0b, 32'hc2bfa677, 32'h429cc98a, 32'hc16a2b8c};
test_output[2726] = '{32'h42b4f586};
test_index[2726] = '{2};
test_input[21816:21823] = '{32'h413e411e, 32'h420d4323, 32'hc2b226a5, 32'h42afae58, 32'h42467d2d, 32'hc251b0fb, 32'h42198007, 32'hc033fc75};
test_output[2727] = '{32'h42afae58};
test_index[2727] = '{3};
test_input[21824:21831] = '{32'hc1a134d2, 32'hc2bfa0b9, 32'hc27b0149, 32'h42bef46a, 32'hc246f3b1, 32'h4213c456, 32'hc1ce626f, 32'h4283087b};
test_output[2728] = '{32'h42bef46a};
test_index[2728] = '{3};
test_input[21832:21839] = '{32'hc29291e5, 32'h42426279, 32'hc2c5e525, 32'hc23d8ceb, 32'h41ed28a4, 32'hc11ee5e1, 32'hc1f197d8, 32'h41ce5f89};
test_output[2729] = '{32'h42426279};
test_index[2729] = '{1};
test_input[21840:21847] = '{32'hc28e81cb, 32'hc26fc628, 32'h420b3962, 32'hc008cc0b, 32'hc2b6ecc0, 32'hc188e9b5, 32'hc202e4b8, 32'hc21e3f06};
test_output[2730] = '{32'h420b3962};
test_index[2730] = '{2};
test_input[21848:21855] = '{32'h42618aee, 32'h42bcf637, 32'h42c0a28e, 32'h42af225c, 32'hc229ddcd, 32'h416cb955, 32'h42b1bb13, 32'hc26d7c53};
test_output[2731] = '{32'h42c0a28e};
test_index[2731] = '{2};
test_input[21856:21863] = '{32'hc1dcf159, 32'hc28ae220, 32'hc2af47d0, 32'hc29981c1, 32'h40b1b6e0, 32'h42acea33, 32'h42b8b1f8, 32'h40f8f1ee};
test_output[2732] = '{32'h42b8b1f8};
test_index[2732] = '{6};
test_input[21864:21871] = '{32'h423e5a64, 32'hc12aa057, 32'h42c02e8f, 32'hc23b688d, 32'h42a0ef2f, 32'hc2a3439d, 32'h4293c772, 32'h410915b2};
test_output[2733] = '{32'h42c02e8f};
test_index[2733] = '{2};
test_input[21872:21879] = '{32'hc2b0a7bd, 32'hc2a7fb7f, 32'hc2744c21, 32'h428db1ab, 32'h411cae12, 32'hc18497c6, 32'hc233f8f1, 32'h42b8b15b};
test_output[2734] = '{32'h42b8b15b};
test_index[2734] = '{7};
test_input[21880:21887] = '{32'h410413c6, 32'hc1f234a6, 32'h410c1097, 32'h41d91acc, 32'h4282fbbe, 32'hc2a07e78, 32'h429c3e40, 32'hbfe9408a};
test_output[2735] = '{32'h429c3e40};
test_index[2735] = '{6};
test_input[21888:21895] = '{32'h40d8e01e, 32'h4260684b, 32'hc23e4191, 32'hc0af7b3d, 32'h42a57e82, 32'h426cba2e, 32'hc2944a37, 32'h429d6185};
test_output[2736] = '{32'h42a57e82};
test_index[2736] = '{4};
test_input[21896:21903] = '{32'h42c39375, 32'hc1656292, 32'hc257abab, 32'h41bcab6a, 32'hc1a6c3b1, 32'hc299b358, 32'hc24fbfc5, 32'hc103959f};
test_output[2737] = '{32'h42c39375};
test_index[2737] = '{0};
test_input[21904:21911] = '{32'hc2098d2e, 32'hc16e330c, 32'hc2774475, 32'h429cf0d3, 32'hc1e01ab5, 32'h417e2374, 32'hc299b333, 32'h42708169};
test_output[2738] = '{32'h429cf0d3};
test_index[2738] = '{3};
test_input[21912:21919] = '{32'h42a1c852, 32'h423e086e, 32'h4260df45, 32'hc1b733b5, 32'h42b61ddd, 32'h41e0963a, 32'h426528a2, 32'h41d85924};
test_output[2739] = '{32'h42b61ddd};
test_index[2739] = '{4};
test_input[21920:21927] = '{32'h42496f1f, 32'hc285fa0e, 32'h42a14e0f, 32'hc150c16f, 32'h42bc6dfc, 32'h42259332, 32'hc09728b8, 32'h4299c2ab};
test_output[2740] = '{32'h42bc6dfc};
test_index[2740] = '{4};
test_input[21928:21935] = '{32'hc2244c1c, 32'h428f9694, 32'h41a6d91a, 32'h428055e2, 32'hc115a92e, 32'h41e1f3fd, 32'hc29d5048, 32'hc29fa051};
test_output[2741] = '{32'h428f9694};
test_index[2741] = '{1};
test_input[21936:21943] = '{32'hc2085bc5, 32'hc299cfdc, 32'hc2ac5c16, 32'h42c66a0d, 32'hc2b16686, 32'h426f277a, 32'hc2c1ea66, 32'h42846ef2};
test_output[2742] = '{32'h42c66a0d};
test_index[2742] = '{3};
test_input[21944:21951] = '{32'h42535ea1, 32'h41c36b8b, 32'hc22703e9, 32'h429c4d84, 32'hc298ba0b, 32'hc26f8c12, 32'h42858835, 32'hc2a9924a};
test_output[2743] = '{32'h429c4d84};
test_index[2743] = '{3};
test_input[21952:21959] = '{32'hc25e7fc6, 32'h425e30aa, 32'h41e4d1a3, 32'hc2895fa5, 32'hc1ac2e87, 32'hc12a775e, 32'hc2b5e641, 32'hbee7a49b};
test_output[2744] = '{32'h425e30aa};
test_index[2744] = '{1};
test_input[21960:21967] = '{32'hc15ba9bd, 32'h424a6f61, 32'hc1d72ca7, 32'h415a6d60, 32'hc29795bd, 32'h421dbe56, 32'hc2b63cc4, 32'h4185e02c};
test_output[2745] = '{32'h424a6f61};
test_index[2745] = '{1};
test_input[21968:21975] = '{32'hc1211a91, 32'h42c3b6c5, 32'h429badf5, 32'h4181b0a1, 32'hc2b96ae6, 32'h425485dc, 32'h42bff699, 32'hc23a92a0};
test_output[2746] = '{32'h42c3b6c5};
test_index[2746] = '{1};
test_input[21976:21983] = '{32'h41356a3f, 32'hc2be1e30, 32'h40c18de5, 32'hc1efd58e, 32'hc21feac8, 32'hc20755f8, 32'hc28f6417, 32'h426abba8};
test_output[2747] = '{32'h426abba8};
test_index[2747] = '{7};
test_input[21984:21991] = '{32'h42523dff, 32'h427f6c9b, 32'hc29f702a, 32'h41dd59ad, 32'h41956ebf, 32'h4295d716, 32'hc19a8599, 32'h40288368};
test_output[2748] = '{32'h4295d716};
test_index[2748] = '{5};
test_input[21992:21999] = '{32'hc27c683b, 32'h4286e4d7, 32'h41277f3c, 32'h4267b081, 32'h4138085b, 32'hc271c6d0, 32'h42198738, 32'hc2b4886f};
test_output[2749] = '{32'h4286e4d7};
test_index[2749] = '{1};
test_input[22000:22007] = '{32'h42b126cc, 32'hc1a05c82, 32'h41b62c50, 32'hc2c7051c, 32'h426c1c0a, 32'hc1ef028c, 32'h41cc39ca, 32'h42944494};
test_output[2750] = '{32'h42b126cc};
test_index[2750] = '{0};
test_input[22008:22015] = '{32'h42b5cd0d, 32'hc297ed32, 32'h413c49d3, 32'h41bd1b0f, 32'h4009b003, 32'h42531f54, 32'h4180015a, 32'h4295937a};
test_output[2751] = '{32'h42b5cd0d};
test_index[2751] = '{0};
test_input[22016:22023] = '{32'h4293dfa6, 32'h4234436f, 32'hc227358e, 32'h3ff5028b, 32'hc184ffd4, 32'hc27865a6, 32'hc2521db1, 32'hc2b5f0d3};
test_output[2752] = '{32'h4293dfa6};
test_index[2752] = '{0};
test_input[22024:22031] = '{32'hbf59437f, 32'hc2308e55, 32'hc25bd86e, 32'h4299f34f, 32'h425d9740, 32'hc271f228, 32'h40025bc5, 32'h428da019};
test_output[2753] = '{32'h4299f34f};
test_index[2753] = '{3};
test_input[22032:22039] = '{32'h41d24888, 32'hc29cc55f, 32'h420ee698, 32'h42a9a7f1, 32'h3d9a0fbc, 32'hc2a13cfd, 32'h41f4deaf, 32'hc23327d5};
test_output[2754] = '{32'h42a9a7f1};
test_index[2754] = '{3};
test_input[22040:22047] = '{32'hc0b60438, 32'hc2801b90, 32'h4020faf3, 32'hc2bd9367, 32'h428d737c, 32'h41ce59b6, 32'hc1c16dab, 32'h40955072};
test_output[2755] = '{32'h428d737c};
test_index[2755] = '{4};
test_input[22048:22055] = '{32'hc215fcf7, 32'hc1ddc632, 32'h42a718cd, 32'hc2b8f28a, 32'hc2be4cef, 32'h4219820b, 32'hc27ebb5c, 32'hc2372c66};
test_output[2756] = '{32'h42a718cd};
test_index[2756] = '{2};
test_input[22056:22063] = '{32'hc2429651, 32'hc2a98ae2, 32'h42adac8a, 32'hc2bb6e00, 32'hc1c26644, 32'hc2798d43, 32'hc26319e9, 32'hc272450a};
test_output[2757] = '{32'h42adac8a};
test_index[2757] = '{2};
test_input[22064:22071] = '{32'hc1882d2a, 32'h40f7da6d, 32'h4254b55d, 32'hc29ebf2a, 32'hc2275d38, 32'hc199ab8c, 32'hc24ad634, 32'hc21ab79f};
test_output[2758] = '{32'h4254b55d};
test_index[2758] = '{2};
test_input[22072:22079] = '{32'h41ba1130, 32'hc295e041, 32'h4235bd60, 32'h42a08635, 32'h42c294c8, 32'h42b27039, 32'h42b77e02, 32'h4115b493};
test_output[2759] = '{32'h42c294c8};
test_index[2759] = '{4};
test_input[22080:22087] = '{32'h424d9fb1, 32'h42b61d2c, 32'hc2254a52, 32'hc26a7d7c, 32'hc265b8ea, 32'h4273865e, 32'hc0ff4d16, 32'hc16ddec4};
test_output[2760] = '{32'h42b61d2c};
test_index[2760] = '{1};
test_input[22088:22095] = '{32'hc1210b1f, 32'hc2367029, 32'h428e313f, 32'hc258f91d, 32'h42aff264, 32'hc2a44dc6, 32'hc2c4ba66, 32'hc11e7460};
test_output[2761] = '{32'h42aff264};
test_index[2761] = '{4};
test_input[22096:22103] = '{32'h424678b6, 32'h42ad36ec, 32'h422a5a95, 32'h428d11cb, 32'h419379cf, 32'h427abce8, 32'h4271d2aa, 32'hc2c1181a};
test_output[2762] = '{32'h42ad36ec};
test_index[2762] = '{1};
test_input[22104:22111] = '{32'h429b558e, 32'hc2805c9f, 32'h4211b2d5, 32'hc206a8a7, 32'h42445fcf, 32'h42c21c82, 32'h409e69cb, 32'hc23201af};
test_output[2763] = '{32'h42c21c82};
test_index[2763] = '{5};
test_input[22112:22119] = '{32'h41f53ded, 32'h41c0a7ec, 32'hc2bb56b3, 32'hc126965e, 32'h41170d88, 32'hc1fea203, 32'h42b1f2f8, 32'h424cc9bb};
test_output[2764] = '{32'h42b1f2f8};
test_index[2764] = '{6};
test_input[22120:22127] = '{32'h419c85aa, 32'h4158cfb5, 32'h4148f673, 32'hc1c75e8e, 32'h42751141, 32'hc1a6d2d7, 32'h409e5120, 32'h42a6cdb8};
test_output[2765] = '{32'h42a6cdb8};
test_index[2765] = '{7};
test_input[22128:22135] = '{32'h41c66c82, 32'h428ae714, 32'hc25cdf93, 32'hc28d9a3c, 32'h428cad61, 32'hc15a4cb5, 32'hc224cccc, 32'h3f6055b6};
test_output[2766] = '{32'h428cad61};
test_index[2766] = '{4};
test_input[22136:22143] = '{32'hc2bc1a0f, 32'h41a23be5, 32'hc13fd71a, 32'h40d4fc94, 32'hc20dc908, 32'h42977b23, 32'hc2bf6a35, 32'hc29fdc43};
test_output[2767] = '{32'h42977b23};
test_index[2767] = '{5};
test_input[22144:22151] = '{32'h4231b671, 32'hc2720114, 32'hc0979d4e, 32'hc20298ce, 32'h421fdf1d, 32'hc1922855, 32'h4287c70e, 32'h429675ba};
test_output[2768] = '{32'h429675ba};
test_index[2768] = '{7};
test_input[22152:22159] = '{32'hc1b49c24, 32'hc28a84ac, 32'h42af4ef2, 32'h4248242f, 32'hc2919491, 32'h4227fa45, 32'h41307e9a, 32'h414af59d};
test_output[2769] = '{32'h42af4ef2};
test_index[2769] = '{2};
test_input[22160:22167] = '{32'h423b30fa, 32'hc09d55f0, 32'h42bb0081, 32'h4280a641, 32'h423b9a28, 32'h4280bbfa, 32'h42596a4b, 32'hc16859f9};
test_output[2770] = '{32'h42bb0081};
test_index[2770] = '{2};
test_input[22168:22175] = '{32'h425e4163, 32'hc2682875, 32'h41c71be4, 32'hc2bd8343, 32'hc180c504, 32'h429352d3, 32'h416f39f8, 32'h426afe74};
test_output[2771] = '{32'h429352d3};
test_index[2771] = '{5};
test_input[22176:22183] = '{32'hc28605b5, 32'h426507c4, 32'hc2bb1c30, 32'h42010dd1, 32'hc266cb12, 32'h42ade129, 32'hc21ef831, 32'h420ed369};
test_output[2772] = '{32'h42ade129};
test_index[2772] = '{5};
test_input[22184:22191] = '{32'h420680b5, 32'hc2be48b0, 32'hc23c23f1, 32'h40e26be5, 32'hc193f568, 32'hc2aaaaa6, 32'hc2b5c143, 32'h405966c0};
test_output[2773] = '{32'h420680b5};
test_index[2773] = '{0};
test_input[22192:22199] = '{32'h42886294, 32'h42a2723d, 32'hc1002740, 32'h4002bd2a, 32'h41d83aff, 32'h4286e9de, 32'h42a7c320, 32'h426cc8c7};
test_output[2774] = '{32'h42a7c320};
test_index[2774] = '{6};
test_input[22200:22207] = '{32'h429aec97, 32'h429ec8e6, 32'h42c29f72, 32'h418d4f74, 32'hbfc1deba, 32'hc2956278, 32'h4281f096, 32'h417b5716};
test_output[2775] = '{32'h42c29f72};
test_index[2775] = '{2};
test_input[22208:22215] = '{32'hc2566e24, 32'hc2b91b8b, 32'hc1cfe920, 32'h4291231e, 32'h41905d4a, 32'hc2666241, 32'hc2a1484c, 32'h421cd4bc};
test_output[2776] = '{32'h4291231e};
test_index[2776] = '{3};
test_input[22216:22223] = '{32'h42a57c93, 32'hc1e816e2, 32'h421ff9dc, 32'hc0c60ad7, 32'h41458062, 32'h42c4edab, 32'hc1ab689d, 32'h425e741e};
test_output[2777] = '{32'h42c4edab};
test_index[2777] = '{5};
test_input[22224:22231] = '{32'h422190fb, 32'h42a3cdd9, 32'h428aec38, 32'h42c11fca, 32'h40dab88a, 32'hc1a0a67c, 32'hc2576894, 32'hc10c7d80};
test_output[2778] = '{32'h42c11fca};
test_index[2778] = '{3};
test_input[22232:22239] = '{32'hc27eca8b, 32'hc2946a45, 32'h429781db, 32'hc203ff0e, 32'hc2a924a3, 32'h423c7d82, 32'h414bd099, 32'h429aa878};
test_output[2779] = '{32'h429aa878};
test_index[2779] = '{7};
test_input[22240:22247] = '{32'hc256f026, 32'h40e41588, 32'h42a38df3, 32'hc15c7177, 32'h42281e3c, 32'hc1ec69ae, 32'h4225084b, 32'h42570d85};
test_output[2780] = '{32'h42a38df3};
test_index[2780] = '{2};
test_input[22248:22255] = '{32'hc2323292, 32'h422f6244, 32'hc27ca74a, 32'hc1d5aa35, 32'h4287f2bd, 32'h420460c6, 32'h42a8b38a, 32'h4227c19c};
test_output[2781] = '{32'h42a8b38a};
test_index[2781] = '{6};
test_input[22256:22263] = '{32'hc2a65110, 32'hc1f0f529, 32'hc18d90aa, 32'h42b6ef50, 32'h423ae496, 32'h42a1c11f, 32'h42986af0, 32'hc2611b70};
test_output[2782] = '{32'h42b6ef50};
test_index[2782] = '{3};
test_input[22264:22271] = '{32'hc22ae143, 32'hc25ff179, 32'hc1f756b0, 32'hc2bec6dc, 32'h423fbf22, 32'h42862998, 32'h429423f6, 32'hc2859cf2};
test_output[2783] = '{32'h429423f6};
test_index[2783] = '{6};
test_input[22272:22279] = '{32'h42c52f83, 32'h4141c0f0, 32'hc1870240, 32'h42337f62, 32'hc2837697, 32'hc248f4ef, 32'hc2641b48, 32'hc26f4904};
test_output[2784] = '{32'h42c52f83};
test_index[2784] = '{0};
test_input[22280:22287] = '{32'h42a069ca, 32'h420e32ee, 32'h4237d387, 32'hc0109ce1, 32'hc12fb320, 32'h3f8abf0a, 32'h42c602a8, 32'h42b1dca0};
test_output[2785] = '{32'h42c602a8};
test_index[2785] = '{6};
test_input[22288:22295] = '{32'hc2b46339, 32'h429d0b00, 32'hc1ae2924, 32'h421aab1c, 32'h42a84817, 32'hc2517dc6, 32'h4087118a, 32'h420c450c};
test_output[2786] = '{32'h42a84817};
test_index[2786] = '{4};
test_input[22296:22303] = '{32'h428261b2, 32'hc1a67b39, 32'h4193081a, 32'hc1d65f6a, 32'hc23ad789, 32'h42b2b123, 32'h417ec4d8, 32'h426eb262};
test_output[2787] = '{32'h42b2b123};
test_index[2787] = '{5};
test_input[22304:22311] = '{32'h42b64722, 32'h42895bbe, 32'h417c6b55, 32'hc26b6aec, 32'hc1415f5d, 32'h4140d436, 32'hc2822c18, 32'h42597d22};
test_output[2788] = '{32'h42b64722};
test_index[2788] = '{0};
test_input[22312:22319] = '{32'hc246afad, 32'hc172251e, 32'h422a2335, 32'hc22449c2, 32'hc2a07134, 32'h42b41473, 32'h4196dc65, 32'hc23c963d};
test_output[2789] = '{32'h42b41473};
test_index[2789] = '{5};
test_input[22320:22327] = '{32'h42160038, 32'h41fb88ac, 32'hc23ebb03, 32'h42b4fc69, 32'hc18737e2, 32'h426ae1f3, 32'h40ea7d29, 32'hc271fd8f};
test_output[2790] = '{32'h42b4fc69};
test_index[2790] = '{3};
test_input[22328:22335] = '{32'hc1880e5d, 32'hc1d4ca2d, 32'hc249a93a, 32'hc26eafc2, 32'h42868818, 32'h41f4a402, 32'h4217e8e0, 32'h4267e231};
test_output[2791] = '{32'h42868818};
test_index[2791] = '{4};
test_input[22336:22343] = '{32'hc2266a91, 32'hc213202e, 32'hc287664b, 32'hc1070127, 32'hc2bb9b59, 32'hc2735e39, 32'hbffb9f6a, 32'h41caee7d};
test_output[2792] = '{32'h41caee7d};
test_index[2792] = '{7};
test_input[22344:22351] = '{32'h42b16202, 32'h4186fbd2, 32'h42297d97, 32'hc1484c79, 32'hc1d72e16, 32'hc2030204, 32'h428ef791, 32'hc08d033c};
test_output[2793] = '{32'h42b16202};
test_index[2793] = '{0};
test_input[22352:22359] = '{32'hc2499fb2, 32'hc1c3d13e, 32'h421166ea, 32'hc2ae9645, 32'h42899c85, 32'hc2c61e74, 32'hc2417d93, 32'hc2b12181};
test_output[2794] = '{32'h42899c85};
test_index[2794] = '{4};
test_input[22360:22367] = '{32'hc226c1eb, 32'hc2997611, 32'hc21a4443, 32'hbfd2e6d7, 32'h421f9bee, 32'hc2956865, 32'hc21525d9, 32'h4045cee6};
test_output[2795] = '{32'h421f9bee};
test_index[2795] = '{4};
test_input[22368:22375] = '{32'hc28aff6b, 32'h41c8fb3b, 32'h42b6c81f, 32'h42aa895c, 32'hc0bc6868, 32'hc262f687, 32'h4214e6de, 32'hc20028b6};
test_output[2796] = '{32'h42b6c81f};
test_index[2796] = '{2};
test_input[22376:22383] = '{32'hc2973995, 32'hc2a023aa, 32'h422bd37b, 32'h427ab40e, 32'hc1d27377, 32'h3e007d54, 32'h42af9bee, 32'hc0f4c472};
test_output[2797] = '{32'h42af9bee};
test_index[2797] = '{6};
test_input[22384:22391] = '{32'hc2bc4367, 32'hc228938d, 32'hc2b23a59, 32'h42946663, 32'h424573ab, 32'h41e6681a, 32'h409902ed, 32'hc1e0e157};
test_output[2798] = '{32'h42946663};
test_index[2798] = '{3};
test_input[22392:22399] = '{32'h42984c01, 32'hc0efa1df, 32'h40ed1d57, 32'hc29fa49d, 32'hc1a0d97e, 32'hc1f238b7, 32'hc157cfbd, 32'hc2c78d76};
test_output[2799] = '{32'h42984c01};
test_index[2799] = '{0};
test_input[22400:22407] = '{32'h40fc68f4, 32'hc25a209c, 32'hc26d4baa, 32'hc1f907e6, 32'h42955fef, 32'h4235363e, 32'h424bda3d, 32'h3ffdf164};
test_output[2800] = '{32'h42955fef};
test_index[2800] = '{4};
test_input[22408:22415] = '{32'hc294177f, 32'h42c1ddae, 32'hc18d39dd, 32'h42375ae6, 32'hc16e6200, 32'h42a9facf, 32'h40ad7b16, 32'hc1d434c4};
test_output[2801] = '{32'h42c1ddae};
test_index[2801] = '{1};
test_input[22416:22423] = '{32'hc2271f1c, 32'hc0cb290a, 32'hc2ac26c7, 32'hc2a07dd0, 32'hbf82fe1b, 32'hc2a92373, 32'hc22cf7bc, 32'hc25faa59};
test_output[2802] = '{32'hbf82fe1b};
test_index[2802] = '{4};
test_input[22424:22431] = '{32'hc228757e, 32'hc2b0170c, 32'h41edbc72, 32'hc2ab698e, 32'hc29d894c, 32'hc1e137de, 32'h425d7bde, 32'h42c363dd};
test_output[2803] = '{32'h42c363dd};
test_index[2803] = '{7};
test_input[22432:22439] = '{32'hc21cda2e, 32'hc28f055e, 32'hc2c0d9ef, 32'h42b57323, 32'h4224b784, 32'hc2a61b73, 32'hc28ec2e3, 32'hc2a0b298};
test_output[2804] = '{32'h42b57323};
test_index[2804] = '{3};
test_input[22440:22447] = '{32'hc17e9b72, 32'hc1823b02, 32'hc21ef299, 32'hc28e89eb, 32'hc28ab166, 32'h418b5262, 32'h42a514c3, 32'h42aadfb2};
test_output[2805] = '{32'h42aadfb2};
test_index[2805] = '{7};
test_input[22448:22455] = '{32'h41b4a74f, 32'h41f317d8, 32'h3f0e2093, 32'hc29cf9cc, 32'h428b7568, 32'hc283c73c, 32'h424710e3, 32'hc207f039};
test_output[2806] = '{32'h428b7568};
test_index[2806] = '{4};
test_input[22456:22463] = '{32'hc244f49a, 32'h4237e6dd, 32'hc2b6710f, 32'h42034701, 32'hc28b450f, 32'hc2c3fa30, 32'h42c6ded1, 32'h42a53900};
test_output[2807] = '{32'h42c6ded1};
test_index[2807] = '{6};
test_input[22464:22471] = '{32'h42bbc519, 32'hc1a6820b, 32'hc29d73d4, 32'h424deae5, 32'hc2c30439, 32'hc1cfa81a, 32'hc26cf0ed, 32'hc2044954};
test_output[2808] = '{32'h42bbc519};
test_index[2808] = '{0};
test_input[22472:22479] = '{32'h429c48ef, 32'h42bde78b, 32'h41c86001, 32'h41e94a25, 32'h41c0d88b, 32'hc18e594f, 32'h4267a7bc, 32'hc20640e0};
test_output[2809] = '{32'h42bde78b};
test_index[2809] = '{1};
test_input[22480:22487] = '{32'h3fd0ef9b, 32'h4270298c, 32'h42949de0, 32'hc2c46d1a, 32'hc203c7d1, 32'hc12119b3, 32'hc21cdb10, 32'h42a101c8};
test_output[2810] = '{32'h42a101c8};
test_index[2810] = '{7};
test_input[22488:22495] = '{32'hc1c382fb, 32'hc27b1967, 32'h42788504, 32'h4264ec9e, 32'h418ce710, 32'h42944874, 32'hc2bbaa5c, 32'h41cc1bf4};
test_output[2811] = '{32'h42944874};
test_index[2811] = '{5};
test_input[22496:22503] = '{32'h42b624ad, 32'hc1a88b3c, 32'h423e808a, 32'hc2b3526b, 32'hc258d2d5, 32'hc191c422, 32'h415eb47f, 32'hc20f8edf};
test_output[2812] = '{32'h42b624ad};
test_index[2812] = '{0};
test_input[22504:22511] = '{32'hc0da367a, 32'h42a19228, 32'hc1e582cf, 32'h422d7644, 32'h41ac1a0e, 32'h42adb7af, 32'hc2aece77, 32'hc263642f};
test_output[2813] = '{32'h42adb7af};
test_index[2813] = '{5};
test_input[22512:22519] = '{32'hc1873a67, 32'hc1c9a003, 32'h4214ae22, 32'h4262e7de, 32'hc1c838df, 32'hc2c3fc69, 32'h41a0b918, 32'h429d93a1};
test_output[2814] = '{32'h429d93a1};
test_index[2814] = '{7};
test_input[22520:22527] = '{32'h41a5e0a7, 32'hc2322025, 32'h423d91c2, 32'h42097966, 32'hc0b1c13b, 32'hc2382916, 32'h42393e59, 32'hc27050cb};
test_output[2815] = '{32'h423d91c2};
test_index[2815] = '{2};
test_input[22528:22535] = '{32'hc240137b, 32'hc238e51b, 32'hc2a1ec06, 32'hc28cf0f4, 32'h42c05fff, 32'hc1515652, 32'h422ad08b, 32'hc297bcf1};
test_output[2816] = '{32'h42c05fff};
test_index[2816] = '{4};
test_input[22536:22543] = '{32'h42321d9b, 32'h41f49acf, 32'h409436df, 32'h4222137d, 32'h4194b7b9, 32'h42871436, 32'h423d6ecf, 32'hc2afadf7};
test_output[2817] = '{32'h42871436};
test_index[2817] = '{5};
test_input[22544:22551] = '{32'hc2abe902, 32'h41258a88, 32'hc2a90a9a, 32'hc2b2716f, 32'hc12773be, 32'hc1ac75cd, 32'hc19540af, 32'h4207ee1f};
test_output[2818] = '{32'h4207ee1f};
test_index[2818] = '{7};
test_input[22552:22559] = '{32'h4251feb7, 32'hc28ba8fa, 32'h42264e85, 32'hc1685b67, 32'hc29133ac, 32'hc29d3e2f, 32'h42430d1c, 32'hc14a8ace};
test_output[2819] = '{32'h4251feb7};
test_index[2819] = '{0};
test_input[22560:22567] = '{32'hc2249a0d, 32'hc13d9d61, 32'hc2b1a8b8, 32'h42a6f47f, 32'hc24f2c75, 32'hc2c2489b, 32'h421a82bf, 32'hc19da023};
test_output[2820] = '{32'h42a6f47f};
test_index[2820] = '{3};
test_input[22568:22575] = '{32'h3f6fd1bb, 32'hc278b397, 32'h4292c751, 32'h42112109, 32'h428f2276, 32'h426e6c43, 32'h428186c3, 32'hc2b0803a};
test_output[2821] = '{32'h4292c751};
test_index[2821] = '{2};
test_input[22576:22583] = '{32'hc201141d, 32'hc183e6c8, 32'h4277d49f, 32'hc2957bc5, 32'hc262935b, 32'hc273691f, 32'h422d3f4c, 32'hc2c454fa};
test_output[2822] = '{32'h4277d49f};
test_index[2822] = '{2};
test_input[22584:22591] = '{32'hc2a0ba80, 32'hc1cdf762, 32'h40be4b45, 32'h426de593, 32'hc2a0d257, 32'h41efcd8e, 32'hc2aedffa, 32'hc2b5eeab};
test_output[2823] = '{32'h426de593};
test_index[2823] = '{3};
test_input[22592:22599] = '{32'hc13d649c, 32'hc29d8780, 32'hc127b6f0, 32'h42befe81, 32'hc2ba39a1, 32'h420e8e86, 32'h42a37cdf, 32'h41b4e8ca};
test_output[2824] = '{32'h42befe81};
test_index[2824] = '{3};
test_input[22600:22607] = '{32'hc22ca458, 32'hc23ea7b2, 32'hc153fa3c, 32'h429083c5, 32'hc2055e08, 32'hc2af37f1, 32'h429dce26, 32'h4280212d};
test_output[2825] = '{32'h429dce26};
test_index[2825] = '{6};
test_input[22608:22615] = '{32'h42853980, 32'hc094039f, 32'hc26c8ef1, 32'hc26eff83, 32'h4293156f, 32'h42bbcb51, 32'h42ac6c34, 32'h4256a415};
test_output[2826] = '{32'h42bbcb51};
test_index[2826] = '{5};
test_input[22616:22623] = '{32'h422f8ade, 32'hc27e9a53, 32'h41daad92, 32'h42bb0e9e, 32'hc1a0840a, 32'h42be7275, 32'hc1d6f8c1, 32'hc2bb8719};
test_output[2827] = '{32'h42be7275};
test_index[2827] = '{5};
test_input[22624:22631] = '{32'h42a44548, 32'h40a69d4f, 32'h41f4b40b, 32'h4232bda7, 32'hc29ecd76, 32'hc12ba528, 32'h418bac4d, 32'hc2730c9d};
test_output[2828] = '{32'h42a44548};
test_index[2828] = '{0};
test_input[22632:22639] = '{32'h4200d1cd, 32'hc2a2b2f4, 32'hc2b84304, 32'hc1dcef14, 32'h42a00972, 32'hc255e4a1, 32'h427ab943, 32'hc2ba4c0c};
test_output[2829] = '{32'h42a00972};
test_index[2829] = '{4};
test_input[22640:22647] = '{32'h42ad6e67, 32'hc1a5b558, 32'h42430cc2, 32'h4198c2d6, 32'h4185d043, 32'hc270827e, 32'h42c4e1f7, 32'h424e2170};
test_output[2830] = '{32'h42c4e1f7};
test_index[2830] = '{6};
test_input[22648:22655] = '{32'hc20d65e3, 32'hc25f8311, 32'h42152cc2, 32'hc2180f78, 32'hc1fb2ce5, 32'hc21f72b7, 32'hc25a786f, 32'hc0ff9bee};
test_output[2831] = '{32'h42152cc2};
test_index[2831] = '{2};
test_input[22656:22663] = '{32'hc27b2f54, 32'h415b1c7a, 32'hc21876e0, 32'h4296eeff, 32'hc15a6af9, 32'h422a7310, 32'hc21b9f25, 32'h42a6c8f7};
test_output[2832] = '{32'h42a6c8f7};
test_index[2832] = '{7};
test_input[22664:22671] = '{32'hc29b4f54, 32'hc2b8465b, 32'h41437f35, 32'h42bbbdb8, 32'h420e7480, 32'h42af9c9d, 32'hc08419d9, 32'hc11072ca};
test_output[2833] = '{32'h42bbbdb8};
test_index[2833] = '{3};
test_input[22672:22679] = '{32'h42b358ad, 32'hc2a9e600, 32'h4227a727, 32'h42937eb2, 32'h4207901c, 32'h42c69f24, 32'h424e10db, 32'hc2a5e6a8};
test_output[2834] = '{32'h42c69f24};
test_index[2834] = '{5};
test_input[22680:22687] = '{32'hc1f095b2, 32'hc2450717, 32'h42b2412e, 32'hc250b512, 32'h418a33ba, 32'h42953f81, 32'h4286c77e, 32'h41ab9649};
test_output[2835] = '{32'h42b2412e};
test_index[2835] = '{2};
test_input[22688:22695] = '{32'hc02cbb92, 32'hc1c5fba9, 32'h4009d5e2, 32'h4296e743, 32'hc28adaa4, 32'h4033968d, 32'hc2a363f9, 32'h424eef04};
test_output[2836] = '{32'h4296e743};
test_index[2836] = '{3};
test_input[22696:22703] = '{32'h41c25c83, 32'hc298232e, 32'hc1453c7d, 32'h3ec19608, 32'h420e72e8, 32'hc285b62c, 32'hc2a60765, 32'h416bfd2b};
test_output[2837] = '{32'h420e72e8};
test_index[2837] = '{4};
test_input[22704:22711] = '{32'h42b240c8, 32'hc2c4eebb, 32'h42848f66, 32'h429e04a7, 32'h421a7c67, 32'hc22399eb, 32'h41f5d8d2, 32'hc293cc07};
test_output[2838] = '{32'h42b240c8};
test_index[2838] = '{0};
test_input[22712:22719] = '{32'hc256b22c, 32'hc29fe58f, 32'h419eab48, 32'hc1abaddb, 32'hc25cfa9a, 32'h418bb721, 32'hc24cd8bf, 32'h4196f7d1};
test_output[2839] = '{32'h419eab48};
test_index[2839] = '{2};
test_input[22720:22727] = '{32'hc2ad05b4, 32'hc208817f, 32'hc29e3eef, 32'h42aa2f05, 32'hbfd83e86, 32'hc1884e9c, 32'hc1e04659, 32'hc1bd1246};
test_output[2840] = '{32'h42aa2f05};
test_index[2840] = '{3};
test_input[22728:22735] = '{32'h422c5403, 32'hc074bea8, 32'hc1c2766d, 32'hc2a6a7b5, 32'hc24040a6, 32'hc1a4ecbd, 32'hc201f488, 32'h421aceba};
test_output[2841] = '{32'h422c5403};
test_index[2841] = '{0};
test_input[22736:22743] = '{32'hc22a42a9, 32'hc253fa7a, 32'hc221e750, 32'h427805e5, 32'hc288c376, 32'hc2a9bc3b, 32'h40fbfce0, 32'h42b3be13};
test_output[2842] = '{32'h42b3be13};
test_index[2842] = '{7};
test_input[22744:22751] = '{32'h42781bea, 32'h428e55ab, 32'h42a16908, 32'h410bd4c7, 32'hc203ea47, 32'hc1467994, 32'hc23b919d, 32'hc2bedcca};
test_output[2843] = '{32'h42a16908};
test_index[2843] = '{2};
test_input[22752:22759] = '{32'hc2856162, 32'h42963840, 32'hc21cc5de, 32'hc20dc9a3, 32'hc292a4be, 32'hc1f4cde6, 32'h41edcb4a, 32'h4297053d};
test_output[2844] = '{32'h4297053d};
test_index[2844] = '{7};
test_input[22760:22767] = '{32'h412c268b, 32'hc282d9ff, 32'h42968a2c, 32'hc105a26a, 32'h42a4e018, 32'hc2413cd2, 32'h40e25806, 32'h42799d4b};
test_output[2845] = '{32'h42a4e018};
test_index[2845] = '{4};
test_input[22768:22775] = '{32'hc249a14c, 32'h40b6eb6c, 32'h41f9871e, 32'h42101a4e, 32'hc2043566, 32'h42a0d8bb, 32'h41b37885, 32'h42332662};
test_output[2846] = '{32'h42a0d8bb};
test_index[2846] = '{5};
test_input[22776:22783] = '{32'hc0c4b99a, 32'h42232bfa, 32'h4134e9f2, 32'hc1b4febd, 32'h4211e8b5, 32'h41a90c41, 32'h42928ff5, 32'h42b45e74};
test_output[2847] = '{32'h42b45e74};
test_index[2847] = '{7};
test_input[22784:22791] = '{32'h424b0e4c, 32'hc294f943, 32'h42a79c17, 32'hc29025ee, 32'hc2c3ca42, 32'hc1f2cffa, 32'hc25c2897, 32'hc11d20e5};
test_output[2848] = '{32'h42a79c17};
test_index[2848] = '{2};
test_input[22792:22799] = '{32'h42874fef, 32'hc2897564, 32'h4196c1d1, 32'h4295298e, 32'h41be7cf5, 32'hc22e004d, 32'h423c25bc, 32'hc29d62bf};
test_output[2849] = '{32'h4295298e};
test_index[2849] = '{3};
test_input[22800:22807] = '{32'hc1184921, 32'hc0e66996, 32'h417bd719, 32'h415d0d04, 32'hc29d0c2c, 32'hc2891637, 32'hc1a3cef4, 32'h42befaac};
test_output[2850] = '{32'h42befaac};
test_index[2850] = '{7};
test_input[22808:22815] = '{32'hc235ce5e, 32'hc1d2c612, 32'hc14f7b4d, 32'hc264e491, 32'h429d5e56, 32'hc2369749, 32'h418d5eb4, 32'h427d9a05};
test_output[2851] = '{32'h429d5e56};
test_index[2851] = '{4};
test_input[22816:22823] = '{32'h42b254d1, 32'h42888b25, 32'h40fce95f, 32'h3f819177, 32'hc1d8f98d, 32'h42a06c0c, 32'h41ee5b97, 32'h41f8389e};
test_output[2852] = '{32'h42b254d1};
test_index[2852] = '{0};
test_input[22824:22831] = '{32'h4291015d, 32'h428b6e24, 32'h4297651e, 32'hc1030dcf, 32'h40d72f83, 32'hc2bdb86f, 32'hc1585c36, 32'h4139e4c9};
test_output[2853] = '{32'h4297651e};
test_index[2853] = '{2};
test_input[22832:22839] = '{32'h42bc12c0, 32'h42951e13, 32'h427077ac, 32'h41f0d5c5, 32'h4291f16b, 32'hc1cfe4ed, 32'h42601072, 32'hbf343430};
test_output[2854] = '{32'h42bc12c0};
test_index[2854] = '{0};
test_input[22840:22847] = '{32'hc0dc58dd, 32'hc1637a18, 32'hc24c9546, 32'h428ac141, 32'hc287a413, 32'hc2a02ac2, 32'hc23f8197, 32'hc1af7b91};
test_output[2855] = '{32'h428ac141};
test_index[2855] = '{3};
test_input[22848:22855] = '{32'h421799f2, 32'hc2b769dc, 32'h4208b508, 32'h427d7b42, 32'hc219c6b8, 32'h42badd6e, 32'h414406cf, 32'h4278336f};
test_output[2856] = '{32'h42badd6e};
test_index[2856] = '{5};
test_input[22856:22863] = '{32'hc28a5dcf, 32'hc12a1fab, 32'h4280d8aa, 32'h42822177, 32'h42a9d499, 32'hc2859c1d, 32'hc20120e8, 32'h42c12f77};
test_output[2857] = '{32'h42c12f77};
test_index[2857] = '{7};
test_input[22864:22871] = '{32'h419fbd2d, 32'h40b604e1, 32'hc221560d, 32'h4284c998, 32'hc227eca2, 32'hc1cb83b1, 32'h4233a93e, 32'h42b58981};
test_output[2858] = '{32'h42b58981};
test_index[2858] = '{7};
test_input[22872:22879] = '{32'hc19a014d, 32'hc27b9491, 32'hc2aa2fe5, 32'h4260cc37, 32'h42171edf, 32'hc23df1a5, 32'hc2b40ebe, 32'hc0120f56};
test_output[2859] = '{32'h4260cc37};
test_index[2859] = '{3};
test_input[22880:22887] = '{32'hc2b96f14, 32'hc10e6387, 32'h4257ff4e, 32'hc0a52618, 32'hc2a0a567, 32'hc186fc1b, 32'h428444c1, 32'hc29157d6};
test_output[2860] = '{32'h428444c1};
test_index[2860] = '{6};
test_input[22888:22895] = '{32'h41c41d3d, 32'h425ba120, 32'h41173000, 32'hc2916016, 32'hc2aee8a6, 32'h407d46de, 32'h42c6fe24, 32'h420dcc17};
test_output[2861] = '{32'h42c6fe24};
test_index[2861] = '{6};
test_input[22896:22903] = '{32'hc15e97d7, 32'hbfaafe4e, 32'h4296d73e, 32'hc2257396, 32'h411c81a9, 32'hc2ad88bc, 32'hc2a9df0c, 32'h42b57525};
test_output[2862] = '{32'h42b57525};
test_index[2862] = '{7};
test_input[22904:22911] = '{32'h429a475e, 32'hc1b67e93, 32'hc2c3cdd9, 32'hc2aad442, 32'hc0593174, 32'h4273b401, 32'hc29d6472, 32'h427327b5};
test_output[2863] = '{32'h429a475e};
test_index[2863] = '{0};
test_input[22912:22919] = '{32'hc1f73a1f, 32'hc2b9e80a, 32'h422e1ac0, 32'h41f88534, 32'h4269dd33, 32'hc03838d7, 32'h428a9f5d, 32'hc2ae53aa};
test_output[2864] = '{32'h428a9f5d};
test_index[2864] = '{6};
test_input[22920:22927] = '{32'hc28c264a, 32'h40845c75, 32'hc19d6985, 32'h42c5c862, 32'hc231a4a4, 32'hc21c106b, 32'h42a20e32, 32'h40d89f61};
test_output[2865] = '{32'h42c5c862};
test_index[2865] = '{3};
test_input[22928:22935] = '{32'hc28f1035, 32'h42102f1c, 32'hc1722ea8, 32'hc28ef7be, 32'h423cd087, 32'h42989254, 32'hc139b2c2, 32'h4239e5f2};
test_output[2866] = '{32'h42989254};
test_index[2866] = '{5};
test_input[22936:22943] = '{32'h421f07f1, 32'hc1aa2ac5, 32'h42ae987a, 32'h429d6227, 32'h42c30dcc, 32'h42b6caed, 32'hc2697a76, 32'hc1289799};
test_output[2867] = '{32'h42c30dcc};
test_index[2867] = '{4};
test_input[22944:22951] = '{32'h418dacd2, 32'hc178a8e6, 32'h4292fdc8, 32'h42a21989, 32'h41f813c5, 32'hc22f6156, 32'hc2c68eb5, 32'hc2b4a1d2};
test_output[2868] = '{32'h42a21989};
test_index[2868] = '{3};
test_input[22952:22959] = '{32'hc2b7fd73, 32'hc1c86fe8, 32'hc1b53f8d, 32'h42966d50, 32'h424dd375, 32'h42b24db0, 32'hc21a9910, 32'hc270aa79};
test_output[2869] = '{32'h42b24db0};
test_index[2869] = '{5};
test_input[22960:22967] = '{32'hc2bb3ed1, 32'h42b9af6b, 32'hc29975a5, 32'hc2a1e984, 32'hc2be3880, 32'hc1528356, 32'h42252944, 32'hc2b21fa7};
test_output[2870] = '{32'h42b9af6b};
test_index[2870] = '{1};
test_input[22968:22975] = '{32'hc244a19f, 32'h4289b8f7, 32'hc2415c8f, 32'hc25019a5, 32'hc1e03c3b, 32'hc2192005, 32'h42b5e0cc, 32'h429a9837};
test_output[2871] = '{32'h42b5e0cc};
test_index[2871] = '{6};
test_input[22976:22983] = '{32'hc250a416, 32'h41518ae7, 32'h42b7c1ef, 32'h412c18fc, 32'h411581ee, 32'hc2b072d1, 32'hc18dbccd, 32'h4280fb47};
test_output[2872] = '{32'h42b7c1ef};
test_index[2872] = '{2};
test_input[22984:22991] = '{32'h41074ee9, 32'h429ea9ba, 32'h41da652f, 32'h429e0700, 32'h42c5f856, 32'h4028793a, 32'hc253d197, 32'h42982806};
test_output[2873] = '{32'h42c5f856};
test_index[2873] = '{4};
test_input[22992:22999] = '{32'hc2a7dd35, 32'hc29337c4, 32'hc2273f2e, 32'hc1a81d51, 32'hc2bac301, 32'hc1afddb8, 32'hc1f6405a, 32'h42c0a033};
test_output[2874] = '{32'h42c0a033};
test_index[2874] = '{7};
test_input[23000:23007] = '{32'h41943152, 32'h424f6b34, 32'h42992cf2, 32'hc1c6bb51, 32'h418ba60e, 32'hc1e2511d, 32'h429c9641, 32'h429926f0};
test_output[2875] = '{32'h429c9641};
test_index[2875] = '{6};
test_input[23008:23015] = '{32'hc2b593e3, 32'h42a0256f, 32'h41a9f2f8, 32'hc2594c4a, 32'hc2117e78, 32'hbee44dcf, 32'h42a54db7, 32'h41df0384};
test_output[2876] = '{32'h42a54db7};
test_index[2876] = '{6};
test_input[23016:23023] = '{32'h41600f8a, 32'hc21eec3d, 32'h3fca09fe, 32'hc281f044, 32'hc28a92c6, 32'hc1262ce1, 32'h412bcdbf, 32'h429e08c8};
test_output[2877] = '{32'h429e08c8};
test_index[2877] = '{7};
test_input[23024:23031] = '{32'hc0200980, 32'h425347ee, 32'h41f165c6, 32'h421f4605, 32'hc22a2f93, 32'h422c4a5d, 32'hc1fdc166, 32'hc2c739fb};
test_output[2878] = '{32'h425347ee};
test_index[2878] = '{1};
test_input[23032:23039] = '{32'h40c327ae, 32'hc27b6a0f, 32'h4286b9fc, 32'h42563312, 32'h42abd00a, 32'h42a6a7a9, 32'h42c59b53, 32'hc2833839};
test_output[2879] = '{32'h42c59b53};
test_index[2879] = '{6};
test_input[23040:23047] = '{32'hc24d94be, 32'hc29726c0, 32'hc22b9761, 32'h429d979e, 32'h41f3f84a, 32'hc2a587f7, 32'hc2506f4e, 32'h41935ab4};
test_output[2880] = '{32'h429d979e};
test_index[2880] = '{3};
test_input[23048:23055] = '{32'h42c3a66f, 32'h41caca67, 32'hc2b0b26c, 32'hc26e060a, 32'h429f05d3, 32'h42ab3278, 32'h42bbf60f, 32'h429d3fb0};
test_output[2881] = '{32'h42c3a66f};
test_index[2881] = '{0};
test_input[23056:23063] = '{32'h422d2ea0, 32'h42721d6e, 32'h41816e0b, 32'h42ac27e2, 32'hc21d6204, 32'hc1fbb99a, 32'hc2640825, 32'hc2bdce8d};
test_output[2882] = '{32'h42ac27e2};
test_index[2882] = '{3};
test_input[23064:23071] = '{32'hc1ef8b26, 32'hc24c4763, 32'h40c06d79, 32'h4262aa69, 32'h41d6b5f1, 32'h40fbbc15, 32'hc230c979, 32'h426d79c5};
test_output[2883] = '{32'h426d79c5};
test_index[2883] = '{7};
test_input[23072:23079] = '{32'h4284e9d4, 32'hc296872c, 32'h427c7054, 32'hc281b6bc, 32'hc200fb31, 32'h40cb6b85, 32'hc2b504bb, 32'h42448647};
test_output[2884] = '{32'h4284e9d4};
test_index[2884] = '{0};
test_input[23080:23087] = '{32'hc199add9, 32'hc2903054, 32'h41302727, 32'hc29bbcb7, 32'h426400a2, 32'h42add1a8, 32'h40892a7e, 32'hc2c0c7a4};
test_output[2885] = '{32'h42add1a8};
test_index[2885] = '{5};
test_input[23088:23095] = '{32'hc22a8552, 32'h408df2ef, 32'hc2c1cf66, 32'h425ced76, 32'hc27eb90a, 32'h428745d5, 32'hc29ebb01, 32'h4156a16c};
test_output[2886] = '{32'h428745d5};
test_index[2886] = '{5};
test_input[23096:23103] = '{32'hc2c5b829, 32'h4188a9f9, 32'h41bdedbf, 32'h4206e4b6, 32'hc282d687, 32'hc207b5cf, 32'h42b109f8, 32'h42049da2};
test_output[2887] = '{32'h42b109f8};
test_index[2887] = '{6};
test_input[23104:23111] = '{32'hc1d14962, 32'h40520227, 32'h41c83f60, 32'hc290df38, 32'hc112c3dc, 32'hc2b0be63, 32'hc2a91148, 32'hc29d8288};
test_output[2888] = '{32'h41c83f60};
test_index[2888] = '{2};
test_input[23112:23119] = '{32'h4263f926, 32'h40249da8, 32'h42526e65, 32'h408604c3, 32'hc2aa404e, 32'h42c6ee21, 32'hc2408ac4, 32'hc269373d};
test_output[2889] = '{32'h42c6ee21};
test_index[2889] = '{5};
test_input[23120:23127] = '{32'hc0a088c4, 32'hc23ebd38, 32'hc2c614d7, 32'hc0fe5fe7, 32'h424c4fb7, 32'hc2b8695c, 32'h4158c48d, 32'h42ac5ffc};
test_output[2890] = '{32'h42ac5ffc};
test_index[2890] = '{7};
test_input[23128:23135] = '{32'hc22801fc, 32'hc1519438, 32'h42bea3b1, 32'h428e06b4, 32'hc0ab582f, 32'hc2abab37, 32'hc2c49168, 32'hc29b535c};
test_output[2891] = '{32'h42bea3b1};
test_index[2891] = '{2};
test_input[23136:23143] = '{32'hc26985e0, 32'hc2b4862c, 32'hc286598c, 32'hc27ada57, 32'hc2bcc010, 32'h42b277c5, 32'h423c0650, 32'hc204b55c};
test_output[2892] = '{32'h42b277c5};
test_index[2892] = '{5};
test_input[23144:23151] = '{32'hc29502f8, 32'h3fb7d39d, 32'hc11e0bd7, 32'h427dc711, 32'hc229f67e, 32'h41cffa85, 32'hc2af61dd, 32'h4204ad03};
test_output[2893] = '{32'h427dc711};
test_index[2893] = '{3};
test_input[23152:23159] = '{32'hc191d066, 32'h42a4a7a9, 32'hc2aa416e, 32'h3ffdf39e, 32'h42b6120c, 32'h4165f398, 32'hc2125141, 32'h420ffa47};
test_output[2894] = '{32'h42b6120c};
test_index[2894] = '{4};
test_input[23160:23167] = '{32'h41589e60, 32'hc296d267, 32'hc264362d, 32'hc1828056, 32'hc1cf28f9, 32'h410fed6b, 32'hc2b4d781, 32'h41de097c};
test_output[2895] = '{32'h41de097c};
test_index[2895] = '{7};
test_input[23168:23175] = '{32'hc05f670f, 32'h40cd2717, 32'h4283a7c5, 32'h42ab23b4, 32'hc2207df7, 32'h4263cce2, 32'h427d8b06, 32'h42b02894};
test_output[2896] = '{32'h42b02894};
test_index[2896] = '{7};
test_input[23176:23183] = '{32'h42717a73, 32'h421426be, 32'hc28096de, 32'hc1f867de, 32'hc29c8d2a, 32'h42b26dd3, 32'h411ff328, 32'hc2aa9aea};
test_output[2897] = '{32'h42b26dd3};
test_index[2897] = '{5};
test_input[23184:23191] = '{32'h40d47a9b, 32'h42ba2003, 32'h4296d46d, 32'hc184455c, 32'hc237c95a, 32'hc2510f29, 32'hc15f83d6, 32'h40f5de5e};
test_output[2898] = '{32'h42ba2003};
test_index[2898] = '{1};
test_input[23192:23199] = '{32'hc23fba41, 32'h421968f8, 32'h42aec2f3, 32'h4295e40a, 32'h42309277, 32'hc2b59ea0, 32'h402c0b1b, 32'hc2bb6261};
test_output[2899] = '{32'h42aec2f3};
test_index[2899] = '{2};
test_input[23200:23207] = '{32'h411c435d, 32'hc1d57b14, 32'hc17f71b4, 32'hc28a5a30, 32'h421e2959, 32'h42057cdd, 32'hc26d3594, 32'h42ae9350};
test_output[2900] = '{32'h42ae9350};
test_index[2900] = '{7};
test_input[23208:23215] = '{32'hc2b57c66, 32'h4280cef3, 32'hc205e54e, 32'hc2046a69, 32'hc24e2f1a, 32'hc289184f, 32'hc19e76c5, 32'h42881cea};
test_output[2901] = '{32'h42881cea};
test_index[2901] = '{7};
test_input[23216:23223] = '{32'hc25a99dc, 32'hc293b6b6, 32'hc0852f02, 32'hc17c7cda, 32'hc19ee2ae, 32'hc196288a, 32'h4280179e, 32'hbf169826};
test_output[2902] = '{32'h4280179e};
test_index[2902] = '{6};
test_input[23224:23231] = '{32'hc20e420b, 32'h42897f61, 32'hc25c46d3, 32'h423944f0, 32'hc2a80b15, 32'h40e1cbf1, 32'h428cad2c, 32'hc259efd0};
test_output[2903] = '{32'h428cad2c};
test_index[2903] = '{6};
test_input[23232:23239] = '{32'hc2aa79b9, 32'h42873c24, 32'h42c647bf, 32'h4265027e, 32'h41a010f9, 32'hc2232f8d, 32'h4299fb42, 32'h41e81d16};
test_output[2904] = '{32'h42c647bf};
test_index[2904] = '{2};
test_input[23240:23247] = '{32'h4147e8f5, 32'hc29f72cf, 32'hc1e8b562, 32'h42bee986, 32'hc2bff2c8, 32'hc1b69b1d, 32'hc292cf6d, 32'hc1aaf73c};
test_output[2905] = '{32'h42bee986};
test_index[2905] = '{3};
test_input[23248:23255] = '{32'h41f1eee3, 32'hc0a27c6b, 32'hc1ce0554, 32'h4242b3fa, 32'h429db275, 32'h4212eae0, 32'h428e8582, 32'hc2986979};
test_output[2906] = '{32'h429db275};
test_index[2906] = '{4};
test_input[23256:23263] = '{32'h42b4e832, 32'h4258f38a, 32'hc22ff5ee, 32'h41fac95a, 32'h42569277, 32'h41e628d6, 32'hc11d6e96, 32'h42c7a0ff};
test_output[2907] = '{32'h42c7a0ff};
test_index[2907] = '{7};
test_input[23264:23271] = '{32'hc2c14946, 32'hc180d9ca, 32'h40bd3066, 32'hc2332eca, 32'h42752334, 32'h42a671d5, 32'hc26a7437, 32'hc290b785};
test_output[2908] = '{32'h42a671d5};
test_index[2908] = '{5};
test_input[23272:23279] = '{32'h40a7811b, 32'hc2b7aa37, 32'hc268217e, 32'h42ab4038, 32'h42796291, 32'h4202740c, 32'hc21e38df, 32'h42940fd2};
test_output[2909] = '{32'h42ab4038};
test_index[2909] = '{3};
test_input[23280:23287] = '{32'hc1bc23f8, 32'hc1bac208, 32'hc27d82cd, 32'hc29db862, 32'hc189fa0b, 32'h42a3238d, 32'h4198eeb6, 32'hc2b1e64d};
test_output[2910] = '{32'h42a3238d};
test_index[2910] = '{5};
test_input[23288:23295] = '{32'h425d563c, 32'hc1aa4485, 32'hc267081b, 32'h429c13e1, 32'hc1fc3c07, 32'hc21e9f6d, 32'h4068c46f, 32'h40967f10};
test_output[2911] = '{32'h429c13e1};
test_index[2911] = '{3};
test_input[23296:23303] = '{32'h42ad8fec, 32'h428a5855, 32'h42778ca5, 32'h40d63bed, 32'hc2a1fec6, 32'h40e901f9, 32'h42af9786, 32'hc2476258};
test_output[2912] = '{32'h42af9786};
test_index[2912] = '{6};
test_input[23304:23311] = '{32'h428e68bf, 32'hc29cbb88, 32'hc2c18a0e, 32'h42b6b45d, 32'h42533292, 32'hc2a7572c, 32'hc2274ef5, 32'hc2984c53};
test_output[2913] = '{32'h42b6b45d};
test_index[2913] = '{3};
test_input[23312:23319] = '{32'h424fbf46, 32'h419c55ac, 32'h41412201, 32'hc230021a, 32'h422f55f3, 32'hc0b9f18f, 32'h42a2c200, 32'hc2433493};
test_output[2914] = '{32'h42a2c200};
test_index[2914] = '{6};
test_input[23320:23327] = '{32'h41908194, 32'h42006f31, 32'hc1e7a197, 32'hc28db56b, 32'h41dc66b7, 32'hc283febb, 32'hc1f11b1a, 32'h41b8ee77};
test_output[2915] = '{32'h42006f31};
test_index[2915] = '{1};
test_input[23328:23335] = '{32'h420b2211, 32'hc2a0fb4d, 32'h429d44f6, 32'h421617e4, 32'h42790476, 32'h4284c7cf, 32'hc25caa9c, 32'hc28743f3};
test_output[2916] = '{32'h429d44f6};
test_index[2916] = '{2};
test_input[23336:23343] = '{32'h42a4b4f6, 32'h42378edd, 32'hc297b3e0, 32'h42afef91, 32'hc24e5371, 32'hc2720ccb, 32'h42c12b05, 32'hc260a534};
test_output[2917] = '{32'h42c12b05};
test_index[2917] = '{6};
test_input[23344:23351] = '{32'h41b2a4a8, 32'hc270ee65, 32'hc2c0875a, 32'hc2730415, 32'hc1320f51, 32'hc15a05aa, 32'h419f099b, 32'h40ebb694};
test_output[2918] = '{32'h41b2a4a8};
test_index[2918] = '{0};
test_input[23352:23359] = '{32'h40e232ef, 32'hc1d4bd19, 32'hc012309b, 32'hc286f62f, 32'hc2207aed, 32'hc1e02d31, 32'hc2c2b4e7, 32'h4266a2ff};
test_output[2919] = '{32'h4266a2ff};
test_index[2919] = '{7};
test_input[23360:23367] = '{32'hc29ba1d0, 32'h426242b0, 32'h42bf96ff, 32'h42399c8a, 32'h41cf3b5d, 32'h4136d3e6, 32'h4299a1ba, 32'h429a3c81};
test_output[2920] = '{32'h42bf96ff};
test_index[2920] = '{2};
test_input[23368:23375] = '{32'hc2b9efe9, 32'hc21d1459, 32'hc27e742b, 32'hc1c312e2, 32'h41d9611d, 32'h41bea352, 32'hc28f0d17, 32'hc2be1e31};
test_output[2921] = '{32'h41d9611d};
test_index[2921] = '{4};
test_input[23376:23383] = '{32'h42b6bd2d, 32'hc2b795f1, 32'hc2c255e6, 32'hc271b9db, 32'hc2c4e102, 32'h428f2ab3, 32'hc1adbb50, 32'hc25cd686};
test_output[2922] = '{32'h42b6bd2d};
test_index[2922] = '{0};
test_input[23384:23391] = '{32'h41d12a98, 32'h42bee78b, 32'h426013cd, 32'h41e69353, 32'hc2b867fa, 32'h4229e196, 32'hc2a22b47, 32'hc2861b4c};
test_output[2923] = '{32'h42bee78b};
test_index[2923] = '{1};
test_input[23392:23399] = '{32'h426b8d6a, 32'h4231a075, 32'hc2959e5b, 32'h41a3953c, 32'h4198958a, 32'hc1927258, 32'hc2be2f81, 32'h420cfd8a};
test_output[2924] = '{32'h426b8d6a};
test_index[2924] = '{0};
test_input[23400:23407] = '{32'h418f2086, 32'h42917c0c, 32'h42263023, 32'hc25a1b53, 32'h42b11a12, 32'hc1725ab0, 32'hc222f271, 32'h420abdd0};
test_output[2925] = '{32'h42b11a12};
test_index[2925] = '{4};
test_input[23408:23415] = '{32'h429c15fb, 32'h4299ee06, 32'hc1ff1c8a, 32'hc2125adf, 32'h4276387d, 32'hc2999ef7, 32'h4195fd30, 32'hc0986814};
test_output[2926] = '{32'h429c15fb};
test_index[2926] = '{0};
test_input[23416:23423] = '{32'hc1db7baf, 32'h429fa398, 32'hc1eabe04, 32'h41a3dcd8, 32'hc2763a42, 32'h42964c0b, 32'h40e1053f, 32'hc29d17b6};
test_output[2927] = '{32'h429fa398};
test_index[2927] = '{1};
test_input[23424:23431] = '{32'hc29cd9d4, 32'hc2404a72, 32'hc287304d, 32'hc0954dd6, 32'hc13579b4, 32'hc2c74bdb, 32'h42acd072, 32'hc251fa04};
test_output[2928] = '{32'h42acd072};
test_index[2928] = '{6};
test_input[23432:23439] = '{32'hc2b226ed, 32'h4241a4e0, 32'h42642eb1, 32'hc296e91e, 32'h423c9d97, 32'hc256e717, 32'hc19a9b59, 32'h428b6ebf};
test_output[2929] = '{32'h428b6ebf};
test_index[2929] = '{7};
test_input[23440:23447] = '{32'h42329d77, 32'h42a468af, 32'h41911e78, 32'hc256650c, 32'hc17a2bee, 32'h42aef78a, 32'h413ca757, 32'hc27eaddf};
test_output[2930] = '{32'h42aef78a};
test_index[2930] = '{5};
test_input[23448:23455] = '{32'h42877dd7, 32'hc2358bf0, 32'h42c0a5bd, 32'hc0f135c8, 32'hc28f0fe7, 32'hc2824e27, 32'hc1aa9207, 32'h42988f18};
test_output[2931] = '{32'h42c0a5bd};
test_index[2931] = '{2};
test_input[23456:23463] = '{32'h42411303, 32'h42a1d7f0, 32'hc2a684f9, 32'hc21186a4, 32'h4280cdf5, 32'h41d68e83, 32'h41e613b0, 32'hc1d8e480};
test_output[2932] = '{32'h42a1d7f0};
test_index[2932] = '{1};
test_input[23464:23471] = '{32'h41eb70c8, 32'h405952b0, 32'hc29403a6, 32'h41354d24, 32'h41fea24a, 32'h42a14dd4, 32'hc083bd18, 32'hc2af2e21};
test_output[2933] = '{32'h42a14dd4};
test_index[2933] = '{5};
test_input[23472:23479] = '{32'h41fa794c, 32'h429c7062, 32'h4224ec64, 32'h42bfdfbd, 32'h42bb5305, 32'h41dc37e3, 32'h42bad844, 32'h411ff747};
test_output[2934] = '{32'h42bfdfbd};
test_index[2934] = '{3};
test_input[23480:23487] = '{32'h429d52be, 32'h423c975d, 32'hc1d27e3f, 32'hc1e6497b, 32'h42afef4b, 32'h413bc226, 32'hc20ef493, 32'h429c1d6b};
test_output[2935] = '{32'h42afef4b};
test_index[2935] = '{4};
test_input[23488:23495] = '{32'hc29845dc, 32'h425e6494, 32'hc260e414, 32'h42abdbef, 32'h42bcc09c, 32'hc2802cd3, 32'hc23d81e6, 32'h422c802f};
test_output[2936] = '{32'h42bcc09c};
test_index[2936] = '{4};
test_input[23496:23503] = '{32'hc1e431fb, 32'h4284fd7f, 32'h41477b96, 32'hc2b5891f, 32'h414182a0, 32'h415a3fcc, 32'h41ab5e33, 32'h42991f91};
test_output[2937] = '{32'h42991f91};
test_index[2937] = '{7};
test_input[23504:23511] = '{32'h413ed59c, 32'hc1bf0f86, 32'hc231b6db, 32'h42a461a9, 32'h42c72105, 32'h4267c55f, 32'hc26e3799, 32'h40c17888};
test_output[2938] = '{32'h42c72105};
test_index[2938] = '{4};
test_input[23512:23519] = '{32'h422c1afd, 32'h4268bedb, 32'hc16c5717, 32'hc1fa5fe4, 32'hc2a3c9cf, 32'hc2256cf5, 32'h424c812b, 32'hc29ccaaf};
test_output[2939] = '{32'h4268bedb};
test_index[2939] = '{1};
test_input[23520:23527] = '{32'h42578f92, 32'hc1a41733, 32'h42537349, 32'h428cfd3d, 32'hc2ba0a29, 32'h4268a8bb, 32'h4213d973, 32'h4169f2ce};
test_output[2940] = '{32'h428cfd3d};
test_index[2940] = '{3};
test_input[23528:23535] = '{32'h427bd310, 32'h404a6b17, 32'h416a2935, 32'h4259481c, 32'hc2a8daaa, 32'h42697074, 32'h42b5b0aa, 32'h428fcac5};
test_output[2941] = '{32'h42b5b0aa};
test_index[2941] = '{6};
test_input[23536:23543] = '{32'hc12203ab, 32'h42967fd8, 32'h422cbb11, 32'h4148cfe6, 32'hbdf7229e, 32'hc29f6ed3, 32'h42661296, 32'h4298a923};
test_output[2942] = '{32'h4298a923};
test_index[2942] = '{7};
test_input[23544:23551] = '{32'hc19105a0, 32'h42ad9f16, 32'h42c35f5b, 32'h41dccb2c, 32'hc09ca67d, 32'hc12c9380, 32'hc25baf19, 32'h3f88f1b8};
test_output[2943] = '{32'h42c35f5b};
test_index[2943] = '{2};
test_input[23552:23559] = '{32'hc2830e5b, 32'hc29db607, 32'h40fe0210, 32'hc2753c1e, 32'h429124ed, 32'hc21cdf3d, 32'hc2a2e5fc, 32'h42bd0036};
test_output[2944] = '{32'h42bd0036};
test_index[2944] = '{7};
test_input[23560:23567] = '{32'h4294cd41, 32'hc2adefcf, 32'h40b05a13, 32'h424ff877, 32'hc186f59f, 32'h40dd1bbf, 32'hc2c6c014, 32'hc23ef0e3};
test_output[2945] = '{32'h4294cd41};
test_index[2945] = '{0};
test_input[23568:23575] = '{32'hc16a4ef6, 32'h4276323d, 32'h42864eb3, 32'h42498377, 32'hc0e06e55, 32'hc280386a, 32'hc2b07f42, 32'hc13e15f4};
test_output[2946] = '{32'h42864eb3};
test_index[2946] = '{2};
test_input[23576:23583] = '{32'h40aaffa8, 32'h42867a7b, 32'h42174a9a, 32'hc1ddd216, 32'hc1cde946, 32'hc2aca4d4, 32'hc23c0324, 32'h429b1130};
test_output[2947] = '{32'h429b1130};
test_index[2947] = '{7};
test_input[23584:23591] = '{32'h42a09935, 32'h42b42c0d, 32'h42bb685e, 32'h40bd4475, 32'hc27a6897, 32'h40dbe8d7, 32'hc0d1c0bb, 32'hc1dd5a41};
test_output[2948] = '{32'h42bb685e};
test_index[2948] = '{2};
test_input[23592:23599] = '{32'h412d82f3, 32'hc2b3d1e7, 32'h408fc783, 32'hc2977a71, 32'hc11b78ca, 32'hc2ad18c6, 32'hc2adb8be, 32'h41f37b84};
test_output[2949] = '{32'h41f37b84};
test_index[2949] = '{7};
test_input[23600:23607] = '{32'h42b6ec44, 32'h42b81310, 32'h42712040, 32'hc2858804, 32'hc27372c7, 32'h42990e3c, 32'h428673d3, 32'hc2532e34};
test_output[2950] = '{32'h42b81310};
test_index[2950] = '{1};
test_input[23608:23615] = '{32'h4299619b, 32'hbf7a49ab, 32'h41bd72f4, 32'h42b6e3de, 32'h42aed7a8, 32'h41ff28d5, 32'h41abe4c8, 32'hc2b4e5ce};
test_output[2951] = '{32'h42b6e3de};
test_index[2951] = '{3};
test_input[23616:23623] = '{32'hc22cbd4e, 32'hbf6a01d5, 32'h41868105, 32'hc29b762a, 32'h41b9fce3, 32'hc1e3e8d8, 32'hc28affca, 32'hc2110d79};
test_output[2952] = '{32'h41b9fce3};
test_index[2952] = '{4};
test_input[23624:23631] = '{32'h428a9f9c, 32'h4297b9e2, 32'h42258581, 32'hc1c573f1, 32'h41b76a63, 32'hc29f86b8, 32'hc2bc7b3c, 32'hc29186d7};
test_output[2953] = '{32'h4297b9e2};
test_index[2953] = '{1};
test_input[23632:23639] = '{32'h422dbd48, 32'hc2b51c97, 32'hc1da0e66, 32'h42aad161, 32'hc20943b8, 32'h41db3bac, 32'h41558715, 32'hc177e9fd};
test_output[2954] = '{32'h42aad161};
test_index[2954] = '{3};
test_input[23640:23647] = '{32'hc2244f63, 32'hc24bb978, 32'h424de247, 32'h4221cedb, 32'hc1f76bee, 32'hc157f068, 32'h425e9981, 32'hc229aeac};
test_output[2955] = '{32'h425e9981};
test_index[2955] = '{6};
test_input[23648:23655] = '{32'h428e0a50, 32'hc1774441, 32'h4176a170, 32'hc1a26ecd, 32'h40b23788, 32'hc231b842, 32'h421545ef, 32'h42c6540d};
test_output[2956] = '{32'h42c6540d};
test_index[2956] = '{7};
test_input[23656:23663] = '{32'h42603d31, 32'hc2366301, 32'h42bce0ee, 32'hc29cf15b, 32'h42197be4, 32'h41e6ac52, 32'h42b0d3b0, 32'hc21e0473};
test_output[2957] = '{32'h42bce0ee};
test_index[2957] = '{2};
test_input[23664:23671] = '{32'h42b03576, 32'h42333696, 32'hc1e30282, 32'hc108e260, 32'hc2831f55, 32'h424fdfd7, 32'h42c4b789, 32'hc26f304a};
test_output[2958] = '{32'h42c4b789};
test_index[2958] = '{6};
test_input[23672:23679] = '{32'hc2041f7e, 32'h426cf8db, 32'h423b0941, 32'h4270e718, 32'hc249c2ae, 32'h41b43ad8, 32'hc29fa9f6, 32'h4215104b};
test_output[2959] = '{32'h4270e718};
test_index[2959] = '{3};
test_input[23680:23687] = '{32'h42645ef8, 32'hc2a14d0b, 32'h4263e8c3, 32'hc16bc643, 32'hc236344f, 32'hc2ae4644, 32'hc0bc1b16, 32'h428678b3};
test_output[2960] = '{32'h428678b3};
test_index[2960] = '{7};
test_input[23688:23695] = '{32'hc1f6381c, 32'hc2bf585b, 32'hc25cf64a, 32'h4119b03c, 32'hc286afe1, 32'hc0e8d6bc, 32'hc20bdc22, 32'hc23f9c06};
test_output[2961] = '{32'h4119b03c};
test_index[2961] = '{3};
test_input[23696:23703] = '{32'h4277c2d7, 32'hc2088dba, 32'hc1ac72d2, 32'h428d848c, 32'hc191df59, 32'h4049eefe, 32'h420c2f4a, 32'hc24f0723};
test_output[2962] = '{32'h428d848c};
test_index[2962] = '{3};
test_input[23704:23711] = '{32'hc2843a42, 32'h426e5d55, 32'hc2ba3ef2, 32'hc2a15c72, 32'hc2b9ef9f, 32'h413e9fea, 32'h40ab3bea, 32'hc2be4a9c};
test_output[2963] = '{32'h426e5d55};
test_index[2963] = '{1};
test_input[23712:23719] = '{32'hc2b4ff6a, 32'hc2b0a2ae, 32'h42a3c63b, 32'hc2c50c13, 32'h411c0d98, 32'hc1971792, 32'h425377f7, 32'hc2a01ebd};
test_output[2964] = '{32'h42a3c63b};
test_index[2964] = '{2};
test_input[23720:23727] = '{32'hc28ad1f7, 32'h41d768e5, 32'h41208d42, 32'hc2b6c663, 32'h42c4bc45, 32'h4284c700, 32'hc22538ce, 32'hc087ed3c};
test_output[2965] = '{32'h42c4bc45};
test_index[2965] = '{4};
test_input[23728:23735] = '{32'h429135d3, 32'h4227c46c, 32'hc26c24bf, 32'h422619f4, 32'h429f6ee8, 32'h4187601b, 32'hc25b423a, 32'hc129a908};
test_output[2966] = '{32'h429f6ee8};
test_index[2966] = '{4};
test_input[23736:23743] = '{32'hc2acaf2c, 32'h429b7b0c, 32'hc1bde707, 32'h40a4fc56, 32'h423c538c, 32'h42bb6079, 32'hc1dcaefc, 32'h4284f3b3};
test_output[2967] = '{32'h42bb6079};
test_index[2967] = '{5};
test_input[23744:23751] = '{32'hc2bbdbf4, 32'h42394694, 32'h420ee096, 32'hc23166a5, 32'h421789a3, 32'h428a6d34, 32'h40dae813, 32'hc19979ca};
test_output[2968] = '{32'h428a6d34};
test_index[2968] = '{5};
test_input[23752:23759] = '{32'h420b2b79, 32'h42a6f645, 32'hc290664d, 32'h428afecf, 32'h42924905, 32'h429a7728, 32'h42a6290b, 32'h42c06945};
test_output[2969] = '{32'h42c06945};
test_index[2969] = '{7};
test_input[23760:23767] = '{32'h40aa1cae, 32'h41b70d0d, 32'h4201ff6c, 32'h423da624, 32'h42abc91e, 32'hc1858354, 32'h42ae4a74, 32'h41a8def1};
test_output[2970] = '{32'h42ae4a74};
test_index[2970] = '{6};
test_input[23768:23775] = '{32'h424d2191, 32'hc1fbe077, 32'hc265585e, 32'hc253890d, 32'hc25c4953, 32'hc25801c9, 32'hc2a21f30, 32'h41c95a00};
test_output[2971] = '{32'h424d2191};
test_index[2971] = '{0};
test_input[23776:23783] = '{32'h42471839, 32'h41c416c0, 32'h424747b7, 32'h41fd5df6, 32'h429f004a, 32'h428944e0, 32'hc1ffd170, 32'hc222c237};
test_output[2972] = '{32'h429f004a};
test_index[2972] = '{4};
test_input[23784:23791] = '{32'h423944ad, 32'h42a786a1, 32'h42b7bd37, 32'h421b2d36, 32'h424718b2, 32'hc25a83ad, 32'hc0dbaff8, 32'h427bafe3};
test_output[2973] = '{32'h42b7bd37};
test_index[2973] = '{2};
test_input[23792:23799] = '{32'hc2bb565b, 32'h42543f6d, 32'hc125a527, 32'h42c2d035, 32'hc2b56f20, 32'h4267b7ff, 32'hc2173b39, 32'h423d4548};
test_output[2974] = '{32'h42c2d035};
test_index[2974] = '{3};
test_input[23800:23807] = '{32'h413259bc, 32'h41a26fbc, 32'h42c701af, 32'hc27f1000, 32'h429f620b, 32'h422d3d11, 32'h426c61a5, 32'hc21aea3f};
test_output[2975] = '{32'h42c701af};
test_index[2975] = '{2};
test_input[23808:23815] = '{32'hc29f4790, 32'h419aa5bb, 32'h4252952b, 32'h427d87b4, 32'hc1941de9, 32'hc15fa867, 32'h42002e00, 32'hc2791da5};
test_output[2976] = '{32'h427d87b4};
test_index[2976] = '{3};
test_input[23816:23823] = '{32'hc07a4fc2, 32'hc29994a5, 32'hbffd41fc, 32'hc04f1c00, 32'hc1ce3db4, 32'hc1e7470f, 32'h429c0199, 32'h429bf43f};
test_output[2977] = '{32'h429c0199};
test_index[2977] = '{6};
test_input[23824:23831] = '{32'h42932915, 32'hc2720594, 32'hc29265e0, 32'h42927a6e, 32'hc276a71c, 32'hc2850d8c, 32'h40681713, 32'h4230326e};
test_output[2978] = '{32'h42932915};
test_index[2978] = '{0};
test_input[23832:23839] = '{32'h4250295a, 32'h42bc1216, 32'hc2928453, 32'hc219559d, 32'h42787fea, 32'h42378264, 32'h41ef2681, 32'h41d01c0c};
test_output[2979] = '{32'h42bc1216};
test_index[2979] = '{1};
test_input[23840:23847] = '{32'hc2c22886, 32'hc2a4fc7f, 32'h42822f65, 32'h415a2dea, 32'hc26321cc, 32'hc2850689, 32'hc170bc5d, 32'hc2a6a696};
test_output[2980] = '{32'h42822f65};
test_index[2980] = '{2};
test_input[23848:23855] = '{32'hc233084a, 32'hc2ad20c7, 32'hc1908aaf, 32'h4224faf6, 32'h4002ec81, 32'hc2b509cd, 32'hc1fe1139, 32'h420d600f};
test_output[2981] = '{32'h4224faf6};
test_index[2981] = '{3};
test_input[23856:23863] = '{32'hc22e17a8, 32'h426c3b32, 32'h4252cc16, 32'hc21a804f, 32'h40f2f728, 32'h40ebe663, 32'h422aaac1, 32'hc2142cab};
test_output[2982] = '{32'h426c3b32};
test_index[2982] = '{1};
test_input[23864:23871] = '{32'hc299a895, 32'hc169ea29, 32'h3f974f08, 32'h42c1d7dd, 32'hc2808f74, 32'hc0f80922, 32'h427e38a9, 32'hc294cb95};
test_output[2983] = '{32'h42c1d7dd};
test_index[2983] = '{3};
test_input[23872:23879] = '{32'hc2bb0fd9, 32'hc25463e4, 32'h42bf9e13, 32'hc2a3ce3a, 32'h427aa440, 32'hc101e2b4, 32'h422d8135, 32'h4259e3cb};
test_output[2984] = '{32'h42bf9e13};
test_index[2984] = '{2};
test_input[23880:23887] = '{32'hc11c2c03, 32'hc1e315f0, 32'h4258dfb9, 32'hc257c29e, 32'h423b1f2b, 32'h429331fb, 32'h421c68f4, 32'h42c3c158};
test_output[2985] = '{32'h42c3c158};
test_index[2985] = '{7};
test_input[23888:23895] = '{32'h429f56b7, 32'h41d94928, 32'hbfa99284, 32'h42c53f89, 32'h4229dcc7, 32'h421dd9cd, 32'hc2a53e06, 32'h42846eec};
test_output[2986] = '{32'h42c53f89};
test_index[2986] = '{3};
test_input[23896:23903] = '{32'hc074d5dd, 32'hc1ad1e99, 32'h4214098a, 32'h42387bda, 32'hc289fa14, 32'h4239c6ee, 32'h4297d3d8, 32'hc20261a7};
test_output[2987] = '{32'h4297d3d8};
test_index[2987] = '{6};
test_input[23904:23911] = '{32'h424d04f7, 32'h41620a8c, 32'hc105d1ae, 32'hc244276b, 32'h3f7b7cd7, 32'hc17ca467, 32'hc2975450, 32'hc23b8ed9};
test_output[2988] = '{32'h424d04f7};
test_index[2988] = '{0};
test_input[23912:23919] = '{32'hc20578cb, 32'hc26c0489, 32'hc06c602c, 32'hc2be06d7, 32'hc2aa4e2d, 32'h428ece00, 32'hc2585a3f, 32'h42adcc41};
test_output[2989] = '{32'h42adcc41};
test_index[2989] = '{7};
test_input[23920:23927] = '{32'hc201f1bc, 32'h4204dd7b, 32'hc1e4584b, 32'h41c60715, 32'hc1868125, 32'hc2ac8685, 32'hc2be0168, 32'h42c1ca1c};
test_output[2990] = '{32'h42c1ca1c};
test_index[2990] = '{7};
test_input[23928:23935] = '{32'h42561359, 32'hc08e24a9, 32'hc0ea277c, 32'hc230e5d9, 32'hc208643d, 32'h428988b0, 32'hc291cd54, 32'hc26fda16};
test_output[2991] = '{32'h428988b0};
test_index[2991] = '{5};
test_input[23936:23943] = '{32'hc112817f, 32'h4201e1c9, 32'h4241c362, 32'h428a9b52, 32'h4278892f, 32'hc1b2208e, 32'hc1b0535c, 32'h413f9d2e};
test_output[2992] = '{32'h428a9b52};
test_index[2992] = '{3};
test_input[23944:23951] = '{32'h4297d12d, 32'h4205dd9c, 32'h42b13cc7, 32'h429c6bb1, 32'hc26e3484, 32'hc21a5808, 32'h4274ae27, 32'h41dbdcf4};
test_output[2993] = '{32'h42b13cc7};
test_index[2993] = '{2};
test_input[23952:23959] = '{32'hc101f2d4, 32'h42817f19, 32'h4148db28, 32'hc27e9339, 32'hc1ce8cb8, 32'hc28bda32, 32'h3f5fa495, 32'hc27f6b6d};
test_output[2994] = '{32'h42817f19};
test_index[2994] = '{1};
test_input[23960:23967] = '{32'h41dfeafd, 32'h425490d4, 32'hc2b5fcf7, 32'h42a819db, 32'hc11c5477, 32'h41dfabc1, 32'h4145e27a, 32'hc2c6ba0f};
test_output[2995] = '{32'h42a819db};
test_index[2995] = '{3};
test_input[23968:23975] = '{32'hc2c1ca03, 32'h421825d7, 32'h42020259, 32'h41c980a2, 32'hc1d9fde4, 32'h42a60238, 32'h42bd5912, 32'hc28dde93};
test_output[2996] = '{32'h42bd5912};
test_index[2996] = '{6};
test_input[23976:23983] = '{32'h422541d4, 32'hc212af70, 32'hc28693c5, 32'hc202889f, 32'h42acf33f, 32'h418ddb63, 32'hc1ee9ffa, 32'h40ccf037};
test_output[2997] = '{32'h42acf33f};
test_index[2997] = '{4};
test_input[23984:23991] = '{32'h427f662f, 32'h420bee9b, 32'h403593a9, 32'hc26d8b64, 32'h42848ba5, 32'hc2947496, 32'h42823a70, 32'hc291d8dd};
test_output[2998] = '{32'h42848ba5};
test_index[2998] = '{4};
test_input[23992:23999] = '{32'hc28d69db, 32'h42963530, 32'h4294d09e, 32'h41101689, 32'h41fd5958, 32'h41a19196, 32'hc2bb6a1e, 32'hc291b183};
test_output[2999] = '{32'h42963530};
test_index[2999] = '{1};
test_input[24000:24007] = '{32'h429a4bc6, 32'hc16f5bf7, 32'h42c7e7ab, 32'h42ab7af7, 32'hc2044cf4, 32'h42aefe0c, 32'h4061a35d, 32'h41f0903e};
test_output[3000] = '{32'h42c7e7ab};
test_index[3000] = '{2};
test_input[24008:24015] = '{32'h4286d980, 32'hc236da40, 32'h41bc0bfe, 32'h41b003d4, 32'hc2b4cfa5, 32'h41a04b10, 32'hc28a2cfe, 32'h42161666};
test_output[3001] = '{32'h4286d980};
test_index[3001] = '{0};
test_input[24016:24023] = '{32'hc266a90b, 32'hc2c1bb16, 32'hc2a03148, 32'h428e1aca, 32'h427e9304, 32'hc28b44bc, 32'hc28bd60f, 32'h418ee4a3};
test_output[3002] = '{32'h428e1aca};
test_index[3002] = '{3};
test_input[24024:24031] = '{32'h41d776bf, 32'hc27e9a40, 32'hc20c4f5c, 32'hc2b2c8c6, 32'hc1198ae1, 32'h42ab0bc1, 32'hc23da636, 32'hc2a4e550};
test_output[3003] = '{32'h42ab0bc1};
test_index[3003] = '{5};
test_input[24032:24039] = '{32'h42ac80bc, 32'hc221f308, 32'h4220bfe6, 32'h423c5ac9, 32'hc22888fa, 32'h42be36a4, 32'h42336711, 32'h41964d98};
test_output[3004] = '{32'h42be36a4};
test_index[3004] = '{5};
test_input[24040:24047] = '{32'hc25b0342, 32'hc2539fd0, 32'hc2c18024, 32'hc16d480d, 32'h404028a4, 32'h4031e551, 32'h4281ba3e, 32'hc240afb8};
test_output[3005] = '{32'h4281ba3e};
test_index[3005] = '{6};
test_input[24048:24055] = '{32'h42c0c375, 32'hc178c98d, 32'h426d28c1, 32'h4280ebfb, 32'h4285de47, 32'h429069dd, 32'hc25735e8, 32'hc021150c};
test_output[3006] = '{32'h42c0c375};
test_index[3006] = '{0};
test_input[24056:24063] = '{32'h42881edc, 32'h40f27e4b, 32'hc299e581, 32'hc2992d0b, 32'h41ae8a0a, 32'h420b6f78, 32'hc29df97e, 32'hbe5f93f4};
test_output[3007] = '{32'h42881edc};
test_index[3007] = '{0};
test_input[24064:24071] = '{32'h42800ecd, 32'hc272cfb1, 32'hc271114f, 32'h41565d0f, 32'hc197aa50, 32'hc12df00a, 32'hc022d327, 32'h4231dc44};
test_output[3008] = '{32'h42800ecd};
test_index[3008] = '{0};
test_input[24072:24079] = '{32'hc2714688, 32'h4114c58f, 32'h41a886ba, 32'h4290458c, 32'hc2c6fa3f, 32'h428a491c, 32'h4273d827, 32'hc23da9ab};
test_output[3009] = '{32'h4290458c};
test_index[3009] = '{3};
test_input[24080:24087] = '{32'h41fda1ce, 32'h4297507d, 32'h41f70d7f, 32'hc18afb69, 32'hc2c295c0, 32'h42c20f96, 32'hc054666c, 32'h4243e244};
test_output[3010] = '{32'h42c20f96};
test_index[3010] = '{5};
test_input[24088:24095] = '{32'h41adc0a9, 32'h42b2be4a, 32'hc207312e, 32'hc27c111b, 32'hc19992ce, 32'h41c8b651, 32'h4271083e, 32'hc24634fc};
test_output[3011] = '{32'h42b2be4a};
test_index[3011] = '{1};
test_input[24096:24103] = '{32'hc2575919, 32'h41ad1d07, 32'h425b67a5, 32'h42af37d0, 32'hc1e827ee, 32'hc2bcff80, 32'h40039f1b, 32'h423c99cf};
test_output[3012] = '{32'h42af37d0};
test_index[3012] = '{3};
test_input[24104:24111] = '{32'h4276c9a8, 32'h4292a8f4, 32'h42a74649, 32'h41a9b4ee, 32'h41fc770b, 32'h429c1ce5, 32'h3fe9be6b, 32'h42957860};
test_output[3013] = '{32'h42a74649};
test_index[3013] = '{2};
test_input[24112:24119] = '{32'h41e433bc, 32'hc24e8ee1, 32'h42140169, 32'h41998641, 32'hc19edc9e, 32'hc2829216, 32'hc2a90065, 32'h41ed2346};
test_output[3014] = '{32'h42140169};
test_index[3014] = '{2};
test_input[24120:24127] = '{32'hc26e2338, 32'h4280abf9, 32'h42be23f2, 32'hc259967b, 32'hc1bd86fb, 32'hc23eea26, 32'h429f101e, 32'h41fc6ed4};
test_output[3015] = '{32'h42be23f2};
test_index[3015] = '{2};
test_input[24128:24135] = '{32'hc2867faa, 32'h4262ed1e, 32'hc296c750, 32'h429f6b30, 32'h42449c8d, 32'h42a6e1ea, 32'hc279aa89, 32'hc1b15e75};
test_output[3016] = '{32'h42a6e1ea};
test_index[3016] = '{5};
test_input[24136:24143] = '{32'hc2463544, 32'hc2241b7d, 32'h42c6de0f, 32'hc2c58fae, 32'h429bdb42, 32'h419a11c8, 32'hc28eeb1c, 32'h40c33ccc};
test_output[3017] = '{32'h42c6de0f};
test_index[3017] = '{2};
test_input[24144:24151] = '{32'hc1a713ca, 32'hc23a1a8f, 32'h428bfe9a, 32'h42a811fa, 32'h421cff6b, 32'hc19ec860, 32'h4235017a, 32'hc2ae676d};
test_output[3018] = '{32'h42a811fa};
test_index[3018] = '{3};
test_input[24152:24159] = '{32'hc1d67f2f, 32'h428418a2, 32'hc133f313, 32'h429111cb, 32'hc11c0ed5, 32'hc29e8203, 32'h42144774, 32'hc276665e};
test_output[3019] = '{32'h429111cb};
test_index[3019] = '{3};
test_input[24160:24167] = '{32'hc1a880fa, 32'hc1f0880a, 32'h4253a168, 32'h42be8435, 32'h411af509, 32'h427c45cf, 32'hc29dbf77, 32'h41f1bd4d};
test_output[3020] = '{32'h42be8435};
test_index[3020] = '{3};
test_input[24168:24175] = '{32'h4153525b, 32'hc28ea24d, 32'h41bbdbed, 32'h42285b48, 32'h41374f29, 32'hc25d0ac1, 32'h42546cac, 32'hc236fcf8};
test_output[3021] = '{32'h42546cac};
test_index[3021] = '{6};
test_input[24176:24183] = '{32'hc2920792, 32'hc2bb7eb1, 32'h42b95252, 32'h422fe5f8, 32'hc2926d27, 32'h429f5f1d, 32'hc26ea7b6, 32'hc274129a};
test_output[3022] = '{32'h42b95252};
test_index[3022] = '{2};
test_input[24184:24191] = '{32'h41570600, 32'h42128d99, 32'hc2c583c0, 32'hc2930189, 32'hc2338e38, 32'hc293ba66, 32'h42b2f912, 32'h42c4d2ff};
test_output[3023] = '{32'h42c4d2ff};
test_index[3023] = '{7};
test_input[24192:24199] = '{32'h42c66d06, 32'hc29af7a4, 32'hc242b3dd, 32'hc22690d5, 32'hc1fd757c, 32'hc21f276a, 32'h42af02e7, 32'hc2b28650};
test_output[3024] = '{32'h42c66d06};
test_index[3024] = '{0};
test_input[24200:24207] = '{32'h424f9138, 32'h42bc6ceb, 32'h4274f153, 32'h417a9b13, 32'hc199e17e, 32'hc2396975, 32'h4131ebf5, 32'hc2b75958};
test_output[3025] = '{32'h42bc6ceb};
test_index[3025] = '{1};
test_input[24208:24215] = '{32'h42a008fb, 32'hc14ad4d4, 32'h417463bc, 32'h416f3ab4, 32'h4295af2a, 32'h42961b51, 32'hc289f762, 32'hc2aceb10};
test_output[3026] = '{32'h42a008fb};
test_index[3026] = '{0};
test_input[24216:24223] = '{32'h42a35afd, 32'h4195f3be, 32'hc1772431, 32'hc2ba0418, 32'h42bd6fff, 32'h40ac8a50, 32'hc28215e1, 32'hc22eb804};
test_output[3027] = '{32'h42bd6fff};
test_index[3027] = '{4};
test_input[24224:24231] = '{32'h4186180b, 32'h42159cc3, 32'h424f3e78, 32'hc2a7f20a, 32'hc2047b68, 32'h429eced9, 32'h42965d25, 32'hc2912b87};
test_output[3028] = '{32'h429eced9};
test_index[3028] = '{5};
test_input[24232:24239] = '{32'h42baa04b, 32'h42aa4ba4, 32'h421604e9, 32'hc2b3e1bd, 32'hc2589186, 32'h40da3d11, 32'h411b47c1, 32'h42962c50};
test_output[3029] = '{32'h42baa04b};
test_index[3029] = '{0};
test_input[24240:24247] = '{32'hc2a53af4, 32'h42055951, 32'hc28cf89d, 32'h3fa082c7, 32'hc27c6922, 32'h42a63b00, 32'hc28d02ca, 32'h4176497f};
test_output[3030] = '{32'h42a63b00};
test_index[3030] = '{5};
test_input[24248:24255] = '{32'h427480bf, 32'hc236e0f1, 32'hc1d612ea, 32'h4201692b, 32'h429c0b75, 32'h42995170, 32'hc224d4af, 32'h42033a2e};
test_output[3031] = '{32'h429c0b75};
test_index[3031] = '{4};
test_input[24256:24263] = '{32'hc1843bfe, 32'hc268b5cc, 32'h429d0fbe, 32'h4176b46b, 32'h42bcf9ea, 32'h40c8134c, 32'hc2b54ae5, 32'hc196a768};
test_output[3032] = '{32'h42bcf9ea};
test_index[3032] = '{4};
test_input[24264:24271] = '{32'h3f3cd7c0, 32'h413601b9, 32'hc244b5cf, 32'h42880d1e, 32'hc0f941de, 32'hc2838563, 32'hc29ba01f, 32'h41c4408c};
test_output[3033] = '{32'h42880d1e};
test_index[3033] = '{3};
test_input[24272:24279] = '{32'hc1fe4b45, 32'h41445fa9, 32'h41207e7c, 32'hc28d3207, 32'h42b4ebe9, 32'hc2ad9efd, 32'hc1c055da, 32'h42487af8};
test_output[3034] = '{32'h42b4ebe9};
test_index[3034] = '{4};
test_input[24280:24287] = '{32'h42b9a7e1, 32'h42b57b33, 32'h41f37ac2, 32'h42c1aac4, 32'h429a1347, 32'hc2904532, 32'hc2333680, 32'hc29802b5};
test_output[3035] = '{32'h42c1aac4};
test_index[3035] = '{3};
test_input[24288:24295] = '{32'h427de1e4, 32'hc23f2220, 32'h429b6ee1, 32'hc14ea210, 32'h423c7a04, 32'hc2459afc, 32'hc28d0854, 32'hc0f148ab};
test_output[3036] = '{32'h429b6ee1};
test_index[3036] = '{2};
test_input[24296:24303] = '{32'hc109ace5, 32'hc247c2d5, 32'h4207f243, 32'hc1dea016, 32'h4213bd49, 32'hc2ba550d, 32'h4281ff96, 32'hc181cbc4};
test_output[3037] = '{32'h4281ff96};
test_index[3037] = '{6};
test_input[24304:24311] = '{32'h4296efc4, 32'hc2a89c54, 32'hc24cafe0, 32'h426cb24c, 32'hc21c8bae, 32'hc24b6c5f, 32'h425b6ce6, 32'hbfc619ad};
test_output[3038] = '{32'h4296efc4};
test_index[3038] = '{0};
test_input[24312:24319] = '{32'h42b0cec6, 32'h41d56942, 32'hc0ea7270, 32'h4137e6d3, 32'h40aaef7b, 32'hc13a5a50, 32'h4253c0ab, 32'h42c3ff52};
test_output[3039] = '{32'h42c3ff52};
test_index[3039] = '{7};
test_input[24320:24327] = '{32'hc16846ad, 32'h428a07e5, 32'hc2410317, 32'hc231c3e4, 32'hc2c14fac, 32'h42955826, 32'hc1abea50, 32'h42906a29};
test_output[3040] = '{32'h42955826};
test_index[3040] = '{5};
test_input[24328:24335] = '{32'hc1712d25, 32'hc29734e0, 32'hc1b76500, 32'hc28252f1, 32'h41506291, 32'h4226365d, 32'hc27ca3db, 32'h425d566e};
test_output[3041] = '{32'h425d566e};
test_index[3041] = '{7};
test_input[24336:24343] = '{32'hc2aa477a, 32'hc2a0a445, 32'hc292f7f4, 32'h42afcd33, 32'h4216da63, 32'h42b38823, 32'hc19d84fa, 32'h41a400ef};
test_output[3042] = '{32'h42b38823};
test_index[3042] = '{5};
test_input[24344:24351] = '{32'h426856cd, 32'hc2996f9d, 32'h429bfe3d, 32'h41e89bc6, 32'h4160b238, 32'hc2986fff, 32'h42954a80, 32'h419985be};
test_output[3043] = '{32'h429bfe3d};
test_index[3043] = '{2};
test_input[24352:24359] = '{32'hc2bb9040, 32'hc24a5791, 32'h42b644e6, 32'h401f4fa8, 32'h419f5348, 32'h420ed99b, 32'h427dce2b, 32'hc0024d2a};
test_output[3044] = '{32'h42b644e6};
test_index[3044] = '{2};
test_input[24360:24367] = '{32'hc27e0731, 32'hc27fa7f6, 32'h420b1595, 32'h42948a4b, 32'h427a5a2d, 32'hc28be5c4, 32'h402a6c74, 32'hc23cd9a6};
test_output[3045] = '{32'h42948a4b};
test_index[3045] = '{3};
test_input[24368:24375] = '{32'hc134ad54, 32'h42368de9, 32'h416c26d3, 32'hc1eb9f7c, 32'h429cc0db, 32'h4174084f, 32'hc2842bd9, 32'hc28eb2aa};
test_output[3046] = '{32'h429cc0db};
test_index[3046] = '{4};
test_input[24376:24383] = '{32'h41ccc58c, 32'h4285a507, 32'hc27677bc, 32'hc0ab1a8c, 32'hc2a864af, 32'hc19225f2, 32'h42bab2af, 32'hc19fcfbb};
test_output[3047] = '{32'h42bab2af};
test_index[3047] = '{6};
test_input[24384:24391] = '{32'hc2547a24, 32'hc229dd39, 32'h41c77363, 32'h425fa5a7, 32'h42b8fb5f, 32'h42a2560c, 32'h421cecca, 32'hc25db22b};
test_output[3048] = '{32'h42b8fb5f};
test_index[3048] = '{4};
test_input[24392:24399] = '{32'h42b724fc, 32'hc219b044, 32'h428360a1, 32'hc260d615, 32'h41aadfd8, 32'h3f906fb3, 32'hc298f52d, 32'hc2001d36};
test_output[3049] = '{32'h42b724fc};
test_index[3049] = '{0};
test_input[24400:24407] = '{32'h4228450a, 32'h41b295b6, 32'hc1fa9c9f, 32'h42a0de7a, 32'h42a7167c, 32'hc2954912, 32'h426de884, 32'hc01fe4d6};
test_output[3050] = '{32'h42a7167c};
test_index[3050] = '{4};
test_input[24408:24415] = '{32'h424dfe3b, 32'h41656e69, 32'h42a11a6d, 32'hc2853bff, 32'hc288f45e, 32'h426922e3, 32'h429ea4d8, 32'h42c726ed};
test_output[3051] = '{32'h42c726ed};
test_index[3051] = '{7};
test_input[24416:24423] = '{32'h41e01f7f, 32'h42492051, 32'hc1d7646c, 32'h42ba393f, 32'hc28b639e, 32'h4287b7de, 32'hc1451985, 32'h42b140a7};
test_output[3052] = '{32'h42ba393f};
test_index[3052] = '{3};
test_input[24424:24431] = '{32'hc0dccb49, 32'h42803ea7, 32'hc18555cf, 32'h41808e86, 32'hc1a5ad47, 32'hc289eeea, 32'h429605da, 32'h42a19553};
test_output[3053] = '{32'h42a19553};
test_index[3053] = '{7};
test_input[24432:24439] = '{32'h3f05e5fb, 32'hc252f913, 32'h42600c09, 32'h427763d0, 32'h424193dd, 32'h410cd059, 32'h42a2103b, 32'hc2759f27};
test_output[3054] = '{32'h42a2103b};
test_index[3054] = '{6};
test_input[24440:24447] = '{32'h42b0e44a, 32'h4294c91d, 32'h42786ad1, 32'h426090c0, 32'hc157130d, 32'h428f6cb4, 32'h4114a4e2, 32'h42481eb0};
test_output[3055] = '{32'h42b0e44a};
test_index[3055] = '{0};
test_input[24448:24455] = '{32'h4124191b, 32'h40cca7f1, 32'h42646385, 32'hc272da4e, 32'hc2992647, 32'h4117a204, 32'hc1cea9c5, 32'hc2a8f8c4};
test_output[3056] = '{32'h42646385};
test_index[3056] = '{2};
test_input[24456:24463] = '{32'hc284ebcb, 32'hc2b47ce8, 32'h42c0cf8f, 32'h42af4f17, 32'hc2947a72, 32'h42972857, 32'h42574d7c, 32'hc19235c6};
test_output[3057] = '{32'h42c0cf8f};
test_index[3057] = '{2};
test_input[24464:24471] = '{32'hc20ed643, 32'h42a76219, 32'hc2aeceeb, 32'hc2704b33, 32'hc1e06950, 32'h425c4873, 32'h42a679ac, 32'hc2222330};
test_output[3058] = '{32'h42a76219};
test_index[3058] = '{1};
test_input[24472:24479] = '{32'hbe1bb4e2, 32'h410fe3bb, 32'hc20832f9, 32'hc29272d4, 32'h428abda5, 32'hc278b197, 32'hc2c7c2c2, 32'hc2aa36a0};
test_output[3059] = '{32'h428abda5};
test_index[3059] = '{4};
test_input[24480:24487] = '{32'hc21ae5e4, 32'h412630ba, 32'hc2958fe2, 32'h42570097, 32'h4270194d, 32'h41ba3f4a, 32'h4252259c, 32'hc2907f45};
test_output[3060] = '{32'h4270194d};
test_index[3060] = '{4};
test_input[24488:24495] = '{32'h428df71b, 32'hc28ac61a, 32'hc1491447, 32'h4249a136, 32'h42528c69, 32'hc2bb5f9c, 32'h4153b6cf, 32'hc1ed9151};
test_output[3061] = '{32'h428df71b};
test_index[3061] = '{0};
test_input[24496:24503] = '{32'hc18fa62c, 32'h429d3d3c, 32'h41490595, 32'hc28dd44e, 32'hc2c3c8c1, 32'h41e7cce2, 32'h427f2bb5, 32'hc2a34d22};
test_output[3062] = '{32'h429d3d3c};
test_index[3062] = '{1};
test_input[24504:24511] = '{32'h4264d8ec, 32'hc15b91b0, 32'h4287b4eb, 32'hc1804142, 32'hc1c16b43, 32'hc267e87c, 32'h41071323, 32'hc28e2fde};
test_output[3063] = '{32'h4287b4eb};
test_index[3063] = '{2};
test_input[24512:24519] = '{32'hc1bd3b36, 32'h42b52ffa, 32'hc1e88a95, 32'h419a95cd, 32'hc29678fc, 32'h40e1a53e, 32'h4227a7fd, 32'h42a01ba8};
test_output[3064] = '{32'h42b52ffa};
test_index[3064] = '{1};
test_input[24520:24527] = '{32'h41a6a891, 32'h41ba944a, 32'h42aca4e4, 32'h428c88ec, 32'hc1ea9d07, 32'h3fe66d4c, 32'h42ac531b, 32'h426eb970};
test_output[3065] = '{32'h42aca4e4};
test_index[3065] = '{2};
test_input[24528:24535] = '{32'h4213dbfb, 32'h4242e594, 32'h42866304, 32'hc2baa5af, 32'h41ea842e, 32'h42ab5797, 32'hc2b557a9, 32'hc106e02b};
test_output[3066] = '{32'h42ab5797};
test_index[3066] = '{5};
test_input[24536:24543] = '{32'h427b347b, 32'h4223ccbc, 32'hc2a83a5a, 32'h426bc004, 32'hc1f25d68, 32'hc08cb6b3, 32'h3f254da8, 32'hc2502470};
test_output[3067] = '{32'h427b347b};
test_index[3067] = '{0};
test_input[24544:24551] = '{32'hc2302851, 32'h429aeff4, 32'hc1c40dfd, 32'h3f4cd9f6, 32'h424730e0, 32'h422720bc, 32'h42ab0609, 32'h421316d6};
test_output[3068] = '{32'h42ab0609};
test_index[3068] = '{6};
test_input[24552:24559] = '{32'hc25dcfef, 32'h42c21bac, 32'hc23d906b, 32'h4267e55b, 32'h4209cbe3, 32'h42c3b5db, 32'h4292baf5, 32'hc225831c};
test_output[3069] = '{32'h42c3b5db};
test_index[3069] = '{5};
test_input[24560:24567] = '{32'h41225a02, 32'hc266bf1d, 32'h42944b82, 32'h42a03df2, 32'hc1dab2f6, 32'h408cb782, 32'h41320b74, 32'hc2793b7f};
test_output[3070] = '{32'h42a03df2};
test_index[3070] = '{3};
test_input[24568:24575] = '{32'hc27eaa51, 32'h428ed547, 32'hc2ba76c0, 32'hc0c8eb4f, 32'h42485434, 32'h42afb6bf, 32'hc21e6325, 32'h421994fb};
test_output[3071] = '{32'h42afb6bf};
test_index[3071] = '{5};
test_input[24576:24583] = '{32'hc2159631, 32'hc221f17f, 32'h42188b0c, 32'h42c190d2, 32'hc1583f07, 32'h4036b221, 32'hc2a0a9f6, 32'hc222c01f};
test_output[3072] = '{32'h42c190d2};
test_index[3072] = '{3};
test_input[24584:24591] = '{32'hc2b523aa, 32'hc2b1a3ac, 32'hc2c7bd61, 32'hc252777a, 32'hbf734708, 32'hc28f0e97, 32'hc2a75e75, 32'h42adb69f};
test_output[3073] = '{32'h42adb69f};
test_index[3073] = '{7};
test_input[24592:24599] = '{32'hc2923b82, 32'h41e0c96b, 32'hc1012fcd, 32'h425d923d, 32'hc29da0a1, 32'hc1d10260, 32'hc2a3d918, 32'h42bb2525};
test_output[3074] = '{32'h42bb2525};
test_index[3074] = '{7};
test_input[24600:24607] = '{32'h42a91886, 32'hc1027b73, 32'h41abd21d, 32'hc23420f9, 32'h42c04976, 32'h42ba8d12, 32'hc20738e3, 32'h429ca304};
test_output[3075] = '{32'h42c04976};
test_index[3075] = '{4};
test_input[24608:24615] = '{32'h421dc1b3, 32'h405a7d1e, 32'h42af19ac, 32'h41eec821, 32'hc2a8dbde, 32'h42a51665, 32'hc0d73f37, 32'hc2b8ea49};
test_output[3076] = '{32'h42af19ac};
test_index[3076] = '{2};
test_input[24616:24623] = '{32'hc29f4f80, 32'hc2b46b0a, 32'hc2656b3d, 32'h428a32dc, 32'hc18744d6, 32'h41f2967a, 32'h4195793f, 32'h403b3097};
test_output[3077] = '{32'h428a32dc};
test_index[3077] = '{3};
test_input[24624:24631] = '{32'h41bdc66a, 32'h4281d02c, 32'h41db582d, 32'hc1a91c6f, 32'h42667b0b, 32'h4194a75d, 32'h4274be38, 32'hc26eae6e};
test_output[3078] = '{32'h4281d02c};
test_index[3078] = '{1};
test_input[24632:24639] = '{32'h428d6b28, 32'h41370b4f, 32'h42bb3cf6, 32'hc27787fb, 32'hc268db60, 32'hc27b539c, 32'h41846c08, 32'h420c67ae};
test_output[3079] = '{32'h42bb3cf6};
test_index[3079] = '{2};
test_input[24640:24647] = '{32'h42050ac0, 32'hc1f0e8f3, 32'h40d93869, 32'h42ac8b04, 32'h4129ae5c, 32'hc28c5f74, 32'hc2672675, 32'hc2abc526};
test_output[3080] = '{32'h42ac8b04};
test_index[3080] = '{3};
test_input[24648:24655] = '{32'hc23f633a, 32'h428f2e80, 32'h428d0aef, 32'hc29dff14, 32'h40ffcb45, 32'hc1d5fc06, 32'h42a95f55, 32'h422baabc};
test_output[3081] = '{32'h42a95f55};
test_index[3081] = '{6};
test_input[24656:24663] = '{32'hc2c16b91, 32'h4225338b, 32'hc0393a25, 32'h40359bd3, 32'h41eef3e8, 32'h425626d2, 32'hc22bbfe7, 32'h4277d4ee};
test_output[3082] = '{32'h4277d4ee};
test_index[3082] = '{7};
test_input[24664:24671] = '{32'hc2b075a8, 32'hc21045a5, 32'h40bd1ce7, 32'hc2b436ed, 32'h42791baf, 32'h3ffc6b46, 32'hc1cde017, 32'h42c2ad0e};
test_output[3083] = '{32'h42c2ad0e};
test_index[3083] = '{7};
test_input[24672:24679] = '{32'hc0802206, 32'h42c10f06, 32'h42a0d4dd, 32'h42a924d6, 32'hc16814ce, 32'hc13c2b9a, 32'hc249e9d5, 32'hc1d01644};
test_output[3084] = '{32'h42c10f06};
test_index[3084] = '{1};
test_input[24680:24687] = '{32'hc1e7c628, 32'h429cc944, 32'hbf3eeeb2, 32'hc2c36280, 32'hc0baac7e, 32'hc27a391f, 32'h423a39bc, 32'h42c03ca5};
test_output[3085] = '{32'h42c03ca5};
test_index[3085] = '{7};
test_input[24688:24695] = '{32'hc28b992b, 32'h4189ec9c, 32'hc18bf10f, 32'h42748dc0, 32'hc2b15f49, 32'h4280ec79, 32'h41331d5b, 32'hc2b9e924};
test_output[3086] = '{32'h4280ec79};
test_index[3086] = '{5};
test_input[24696:24703] = '{32'hc2c15def, 32'hc2b638c6, 32'h42472575, 32'hc1c45a7d, 32'h4081dee1, 32'hc1d89ec3, 32'hc21f1cdf, 32'hc25426bc};
test_output[3087] = '{32'h42472575};
test_index[3087] = '{2};
test_input[24704:24711] = '{32'hc220e041, 32'hc21766bc, 32'h41cff7bf, 32'hc29b6283, 32'hc1bdc9ca, 32'h41ff8996, 32'h42094a7a, 32'h42aa4144};
test_output[3088] = '{32'h42aa4144};
test_index[3088] = '{7};
test_input[24712:24719] = '{32'h428faadb, 32'hc28209b0, 32'hc22e3124, 32'hc2456dfd, 32'hc13a859e, 32'h42bde24e, 32'h426e3048, 32'hc28276dd};
test_output[3089] = '{32'h42bde24e};
test_index[3089] = '{5};
test_input[24720:24727] = '{32'h427fee91, 32'hc1e5f9fc, 32'hc1b1a937, 32'h4234f199, 32'h42bbddb3, 32'hc2a84111, 32'h40e3d1df, 32'hc08907aa};
test_output[3090] = '{32'h42bbddb3};
test_index[3090] = '{4};
test_input[24728:24735] = '{32'h41f2d57e, 32'h41936a1c, 32'h41f0650f, 32'hc15098ae, 32'h42946632, 32'h421baab6, 32'h425e08d4, 32'h4222565d};
test_output[3091] = '{32'h42946632};
test_index[3091] = '{4};
test_input[24736:24743] = '{32'h41f9f8d2, 32'h42095d6e, 32'hc224f279, 32'hc00498ff, 32'hc1a4d63b, 32'hc2a925a2, 32'h4251a4c3, 32'h41ef0a49};
test_output[3092] = '{32'h4251a4c3};
test_index[3092] = '{6};
test_input[24744:24751] = '{32'h42be7c0a, 32'h41ed73ee, 32'h40bcb9d3, 32'h41484147, 32'h42434c6d, 32'hc169d29f, 32'h4293de75, 32'hc260885b};
test_output[3093] = '{32'h42be7c0a};
test_index[3093] = '{0};
test_input[24752:24759] = '{32'hc2a98162, 32'h4092cb7a, 32'hc1b1509b, 32'h424d6ce9, 32'h42858962, 32'h40d18470, 32'h4147c134, 32'hbfc95c37};
test_output[3094] = '{32'h42858962};
test_index[3094] = '{4};
test_input[24760:24767] = '{32'h4220c1d2, 32'h41cb1684, 32'h40b1a0dd, 32'h401a3795, 32'h41a27ea1, 32'hc23f00df, 32'hc1c831e4, 32'hc2be12fa};
test_output[3095] = '{32'h4220c1d2};
test_index[3095] = '{0};
test_input[24768:24775] = '{32'h4189c743, 32'h41809aec, 32'hc225b65c, 32'hc137676e, 32'h428c1f6f, 32'hc1a04776, 32'hc2a39577, 32'hc2854bae};
test_output[3096] = '{32'h428c1f6f};
test_index[3096] = '{4};
test_input[24776:24783] = '{32'hc1cb8543, 32'h42636cea, 32'hc1813eb5, 32'hc0905554, 32'hc1b4fc8d, 32'hc28ccf54, 32'hc20ea6f8, 32'hc1422b74};
test_output[3097] = '{32'h42636cea};
test_index[3097] = '{1};
test_input[24784:24791] = '{32'h4297ed17, 32'h4179978f, 32'h424824ca, 32'h42c63760, 32'hc11ec81a, 32'hc2b07984, 32'hc2861e5f, 32'h422405f4};
test_output[3098] = '{32'h42c63760};
test_index[3098] = '{3};
test_input[24792:24799] = '{32'hc276e696, 32'h42057157, 32'h42b32e8f, 32'h42941875, 32'h4281b093, 32'h42b53774, 32'h426f33f7, 32'hc29b55cc};
test_output[3099] = '{32'h42b53774};
test_index[3099] = '{5};
test_input[24800:24807] = '{32'h41f928be, 32'h42a0d972, 32'hc1fbba56, 32'hc2c6b415, 32'hc270d9af, 32'h42a6c81c, 32'hc2b813bb, 32'hc0b2b2de};
test_output[3100] = '{32'h42a6c81c};
test_index[3100] = '{5};
test_input[24808:24815] = '{32'h42ba21c0, 32'h40073fdc, 32'h423afbf4, 32'hc208a9a1, 32'h42157ca9, 32'h4291317f, 32'h3fbf595b, 32'h41afc662};
test_output[3101] = '{32'h42ba21c0};
test_index[3101] = '{0};
test_input[24816:24823] = '{32'hc237b3cc, 32'h4269e595, 32'hc2387ec2, 32'h42aa4380, 32'h429579cb, 32'h42ab5d53, 32'hc2bba496, 32'h42684842};
test_output[3102] = '{32'h42ab5d53};
test_index[3102] = '{5};
test_input[24824:24831] = '{32'hc21265ed, 32'hc28df16a, 32'h42c1b1a8, 32'hc20c6886, 32'h41ba6eb9, 32'hc2827e3b, 32'h428eff51, 32'h4214e6c9};
test_output[3103] = '{32'h42c1b1a8};
test_index[3103] = '{2};
test_input[24832:24839] = '{32'hc2aed12b, 32'h42606d92, 32'h41c76151, 32'hc2a014b1, 32'h41db890f, 32'hc1b5c6d9, 32'hc20c4275, 32'hc2a4aba4};
test_output[3104] = '{32'h42606d92};
test_index[3104] = '{1};
test_input[24840:24847] = '{32'h4201b1fb, 32'hc1c67216, 32'hc2b4f7da, 32'hc1d34bb3, 32'hc234a4ca, 32'hc2acc9a8, 32'h423fc747, 32'hc23dc7bf};
test_output[3105] = '{32'h423fc747};
test_index[3105] = '{6};
test_input[24848:24855] = '{32'hc21ca539, 32'hc2573e0b, 32'hc2491280, 32'h421e362c, 32'h42b0a6ce, 32'h428e7f43, 32'h42c1ba93, 32'h4172d3aa};
test_output[3106] = '{32'h42c1ba93};
test_index[3106] = '{6};
test_input[24856:24863] = '{32'h42c16cce, 32'h4116b11c, 32'h42ac5b8a, 32'h40cfede5, 32'hc07e404c, 32'hc15befc6, 32'h42680850, 32'hc1ffc09e};
test_output[3107] = '{32'h42c16cce};
test_index[3107] = '{0};
test_input[24864:24871] = '{32'h42bd4859, 32'h4126913f, 32'hc26b4d11, 32'h42277d02, 32'hc265d48a, 32'hc22f19c0, 32'hc2525c9d, 32'h411756f3};
test_output[3108] = '{32'h42bd4859};
test_index[3108] = '{0};
test_input[24872:24879] = '{32'h41bb2aa9, 32'hc25832a6, 32'hc0ddd605, 32'h41db3fc2, 32'hc295693f, 32'hc10984f1, 32'h424773f1, 32'h416cf35c};
test_output[3109] = '{32'h424773f1};
test_index[3109] = '{6};
test_input[24880:24887] = '{32'h4290aad3, 32'h42a46921, 32'h4281e411, 32'h424cb32a, 32'h42bf7d71, 32'h3f742a0b, 32'hc2642a71, 32'h4209f98e};
test_output[3110] = '{32'h42bf7d71};
test_index[3110] = '{4};
test_input[24888:24895] = '{32'hc1aad353, 32'hc20e5bec, 32'h42af308c, 32'hc2731464, 32'h4296ff01, 32'h4186158e, 32'hc2aa614d, 32'h42b719d2};
test_output[3111] = '{32'h42b719d2};
test_index[3111] = '{7};
test_input[24896:24903] = '{32'h42bd5b06, 32'hc20eba77, 32'h42b40f14, 32'h424c9cc1, 32'hc2601669, 32'h42b0df7c, 32'hc2b40804, 32'h41d337e0};
test_output[3112] = '{32'h42bd5b06};
test_index[3112] = '{0};
test_input[24904:24911] = '{32'hc1ef48fe, 32'h428bc752, 32'h42956f5d, 32'hc29d7edd, 32'hc24068db, 32'hc1f2a558, 32'h429e1d28, 32'hc2bb3c1c};
test_output[3113] = '{32'h429e1d28};
test_index[3113] = '{6};
test_input[24912:24919] = '{32'h42a909d5, 32'hc23ff5a4, 32'hc26a4004, 32'h419ae8fb, 32'hc1a838e8, 32'hc206787c, 32'h42b45734, 32'hc277b5f9};
test_output[3114] = '{32'h42b45734};
test_index[3114] = '{6};
test_input[24920:24927] = '{32'hc23c858b, 32'hc1f0546d, 32'h423d14cb, 32'h420b6d5b, 32'hc24dd7da, 32'hc1a6f758, 32'h42b451c9, 32'h423d7245};
test_output[3115] = '{32'h42b451c9};
test_index[3115] = '{6};
test_input[24928:24935] = '{32'h4055db61, 32'h42116cf0, 32'h429985d5, 32'hc2a204bb, 32'hc16f43ae, 32'hc17140c1, 32'hc19f3ac9, 32'h413d53d1};
test_output[3116] = '{32'h429985d5};
test_index[3116] = '{2};
test_input[24936:24943] = '{32'hc20ede8f, 32'hc1643f87, 32'h429d0d30, 32'h42a3cb82, 32'h41a4c1d7, 32'hc25bd2c7, 32'hc2a2ac06, 32'h425f2b77};
test_output[3117] = '{32'h42a3cb82};
test_index[3117] = '{3};
test_input[24944:24951] = '{32'h41dbf378, 32'h4180f270, 32'hc088f824, 32'hc24acfdd, 32'hc0beee66, 32'h41b8ec28, 32'hc15887fa, 32'h4244a3e4};
test_output[3118] = '{32'h4244a3e4};
test_index[3118] = '{7};
test_input[24952:24959] = '{32'h41459cd9, 32'h4298b6fb, 32'h41a71ad4, 32'h429455da, 32'hc284a8aa, 32'hc1c24157, 32'h426e6711, 32'hc2c65d3a};
test_output[3119] = '{32'h4298b6fb};
test_index[3119] = '{1};
test_input[24960:24967] = '{32'hc1feb14c, 32'h41b70af4, 32'h419b59c7, 32'hc2641030, 32'hc26771dd, 32'h42455f56, 32'h4177028e, 32'h429ed210};
test_output[3120] = '{32'h429ed210};
test_index[3120] = '{7};
test_input[24968:24975] = '{32'h407257cc, 32'hc1a8702c, 32'hc29e49c9, 32'h41b2ea03, 32'hc28936ee, 32'h424ac124, 32'h42ae8736, 32'hc2af9f33};
test_output[3121] = '{32'h42ae8736};
test_index[3121] = '{6};
test_input[24976:24983] = '{32'hc2921137, 32'h42679fdd, 32'hc2c4e2bc, 32'h4244dd91, 32'hc27398c4, 32'hc1ef5e09, 32'hc23e7db9, 32'h42306ff0};
test_output[3122] = '{32'h42679fdd};
test_index[3122] = '{1};
test_input[24984:24991] = '{32'h40b59f71, 32'h3ec1618f, 32'hc1b5a5fa, 32'hc2bf3e4d, 32'h42a331a4, 32'h412f8e23, 32'hbf3f80e1, 32'h423ddc5d};
test_output[3123] = '{32'h42a331a4};
test_index[3123] = '{4};
test_input[24992:24999] = '{32'hc2bc7d4c, 32'hc1b9ce98, 32'h3fd24775, 32'h4287b0a2, 32'hc2858d30, 32'h42aaf2c3, 32'hbf1a30bd, 32'hc2825e2c};
test_output[3124] = '{32'h42aaf2c3};
test_index[3124] = '{5};
test_input[25000:25007] = '{32'hc18d0afd, 32'hc284cc8a, 32'hc1ba3d4e, 32'h42be1a62, 32'h4230c31c, 32'h40b19c65, 32'hc1f5b4f0, 32'hc2b884cf};
test_output[3125] = '{32'h42be1a62};
test_index[3125] = '{3};
test_input[25008:25015] = '{32'hc2c70128, 32'h41cabd60, 32'hc1ea3951, 32'hc20cf540, 32'h42ad91fc, 32'h421491f0, 32'hc2704466, 32'h401fe245};
test_output[3126] = '{32'h42ad91fc};
test_index[3126] = '{4};
test_input[25016:25023] = '{32'hc170825d, 32'h4255aab4, 32'h408710ef, 32'h411ae21b, 32'h422b7f45, 32'h421b8e75, 32'hc2a830b0, 32'h418a36ac};
test_output[3127] = '{32'h4255aab4};
test_index[3127] = '{1};
test_input[25024:25031] = '{32'h424304cf, 32'hc0860620, 32'h429ec280, 32'h41ec1530, 32'h4209cbda, 32'h42b9537e, 32'hc21bfb74, 32'hc211e945};
test_output[3128] = '{32'h42b9537e};
test_index[3128] = '{5};
test_input[25032:25039] = '{32'hc17f73d5, 32'hc09f13b3, 32'h42935699, 32'hc14b61cf, 32'h41c5b013, 32'h42be5490, 32'h42b56bb6, 32'h421093a0};
test_output[3129] = '{32'h42be5490};
test_index[3129] = '{5};
test_input[25040:25047] = '{32'hc27ab151, 32'hc0310a29, 32'h41bb9c3d, 32'h422bef80, 32'hc2ab169e, 32'h429e70a6, 32'h42b2d5e9, 32'hc25b9324};
test_output[3130] = '{32'h42b2d5e9};
test_index[3130] = '{6};
test_input[25048:25055] = '{32'hc29e626b, 32'hc2beae1e, 32'hc2125259, 32'h41d74445, 32'h42375f77, 32'h422a436e, 32'hc006597c, 32'hc2846d48};
test_output[3131] = '{32'h42375f77};
test_index[3131] = '{4};
test_input[25056:25063] = '{32'hc1b0a8f5, 32'hc13b9046, 32'h3f9e0730, 32'h42594720, 32'hc156019f, 32'hc215e70c, 32'hc2af7495, 32'hc183bea3};
test_output[3132] = '{32'h42594720};
test_index[3132] = '{3};
test_input[25064:25071] = '{32'h42bbdd17, 32'h42c2ff33, 32'h41d2a835, 32'hc28dc2dc, 32'hc23a722f, 32'h42b1df51, 32'hc29a5bbd, 32'hc195e54f};
test_output[3133] = '{32'h42c2ff33};
test_index[3133] = '{1};
test_input[25072:25079] = '{32'h4209b9b2, 32'h42a33f8e, 32'h42a9fd1d, 32'h420aedae, 32'h4254a3c9, 32'h42688823, 32'hc235e5ee, 32'h410a109e};
test_output[3134] = '{32'h42a9fd1d};
test_index[3134] = '{2};
test_input[25080:25087] = '{32'h422758f0, 32'h428a4bf1, 32'hbfac0ac3, 32'h42379754, 32'hc18e7b26, 32'hc19798c0, 32'hc2c13786, 32'h41dcc820};
test_output[3135] = '{32'h428a4bf1};
test_index[3135] = '{1};
test_input[25088:25095] = '{32'h424b3ad8, 32'hc1f7a4e2, 32'hc1d5a2fc, 32'hc0b43478, 32'hc2a0fe54, 32'h41dba295, 32'hc2ac7986, 32'hc093c422};
test_output[3136] = '{32'h424b3ad8};
test_index[3136] = '{0};
test_input[25096:25103] = '{32'h42782071, 32'hc28a5a36, 32'h4260cf27, 32'hc1c02a06, 32'hc22217c7, 32'hc1488d8a, 32'hc1f2f4d9, 32'h4197f9da};
test_output[3137] = '{32'h42782071};
test_index[3137] = '{0};
test_input[25104:25111] = '{32'h425ee79d, 32'h423a71bf, 32'h421a439d, 32'h3f9a78ce, 32'h4214be12, 32'hc22be295, 32'h41c374e4, 32'hc2ad7e38};
test_output[3138] = '{32'h425ee79d};
test_index[3138] = '{0};
test_input[25112:25119] = '{32'h42486b6b, 32'h4259c1d4, 32'hc250174d, 32'h42805c4e, 32'h4130d07f, 32'h41c6cf1b, 32'hc21e71e7, 32'hc1d5c805};
test_output[3139] = '{32'h42805c4e};
test_index[3139] = '{3};
test_input[25120:25127] = '{32'h42095d35, 32'hc27a9c2a, 32'hc0b0abfc, 32'h42740fac, 32'hc1b6ab6a, 32'h41b0bcac, 32'h42048294, 32'hc24a4c67};
test_output[3140] = '{32'h42740fac};
test_index[3140] = '{3};
test_input[25128:25135] = '{32'h4232cf21, 32'hc1eca2cb, 32'h414e2224, 32'hc1afe680, 32'hc243b74e, 32'hc2449a37, 32'h429bc7c7, 32'hc20c5422};
test_output[3141] = '{32'h429bc7c7};
test_index[3141] = '{6};
test_input[25136:25143] = '{32'h428a934a, 32'hc2b53750, 32'h428ed329, 32'hc277c7d3, 32'hc2836b9c, 32'h42617247, 32'hc29a2071, 32'h4195e3cf};
test_output[3142] = '{32'h428ed329};
test_index[3142] = '{2};
test_input[25144:25151] = '{32'hc2b3cc8a, 32'hc256bd79, 32'hc2849b22, 32'h4190bcc8, 32'h42437e50, 32'hc22672cb, 32'h42b7cf17, 32'hc1660e7a};
test_output[3143] = '{32'h42b7cf17};
test_index[3143] = '{6};
test_input[25152:25159] = '{32'hc2b3d9f7, 32'hc154f572, 32'h413fc644, 32'hc23617fd, 32'h426fb547, 32'hc23a3012, 32'hc2894f14, 32'h42a48e5d};
test_output[3144] = '{32'h42a48e5d};
test_index[3144] = '{7};
test_input[25160:25167] = '{32'h41a4da41, 32'h429fc587, 32'h424b1873, 32'hc18e3dac, 32'hc28337df, 32'h41f1c8a8, 32'h423bad78, 32'h41eb64c5};
test_output[3145] = '{32'h429fc587};
test_index[3145] = '{1};
test_input[25168:25175] = '{32'h42451eba, 32'h42b655e9, 32'hc1eab814, 32'hc11789f3, 32'h42b8badb, 32'h425d358e, 32'hc256b700, 32'h42bb373d};
test_output[3146] = '{32'h42bb373d};
test_index[3146] = '{7};
test_input[25176:25183] = '{32'hc2b01755, 32'h4195172f, 32'hc2b84cb6, 32'h4248715b, 32'h41b03d31, 32'h422dd909, 32'h42297d72, 32'hc137fbfe};
test_output[3147] = '{32'h4248715b};
test_index[3147] = '{3};
test_input[25184:25191] = '{32'hc2148b30, 32'h407785a0, 32'h41a517f2, 32'hc2af1c04, 32'h4241ea44, 32'h42b06df2, 32'h41819957, 32'h3f491255};
test_output[3148] = '{32'h42b06df2};
test_index[3148] = '{5};
test_input[25192:25199] = '{32'hc22211e3, 32'h429bab61, 32'h42b56a9a, 32'h4296bdcb, 32'hc272c484, 32'hc0614f7b, 32'hc2bf61c1, 32'h4283c558};
test_output[3149] = '{32'h42b56a9a};
test_index[3149] = '{2};
test_input[25200:25207] = '{32'hc1fd0a3c, 32'hc2c6dae5, 32'h42a604e1, 32'h41f2b0f9, 32'hc0bf2ceb, 32'h41a0f7a4, 32'hc0d3bd7a, 32'hc1b78023};
test_output[3150] = '{32'h42a604e1};
test_index[3150] = '{2};
test_input[25208:25215] = '{32'hc2bf33ce, 32'h42c3b124, 32'hc11e6a4b, 32'h42beae07, 32'hc27f8dbe, 32'hc004b952, 32'hc2be312d, 32'hc1ae7b24};
test_output[3151] = '{32'h42c3b124};
test_index[3151] = '{1};
test_input[25216:25223] = '{32'h415f96c3, 32'h424adc33, 32'h42b0be77, 32'hc06adfd5, 32'h41ac7c79, 32'h41d9bb55, 32'hc25a0959, 32'hc2849fdf};
test_output[3152] = '{32'h42b0be77};
test_index[3152] = '{2};
test_input[25224:25231] = '{32'hc17a616d, 32'hc29741da, 32'h421860f0, 32'h42b4b3e9, 32'hc2ba01f0, 32'hc26e5154, 32'hc255babb, 32'hc236fa88};
test_output[3153] = '{32'h42b4b3e9};
test_index[3153] = '{3};
test_input[25232:25239] = '{32'hc2b7e4b3, 32'h40c662cf, 32'hc27d3c00, 32'hc1851957, 32'hc2c086dc, 32'h42720cab, 32'hc205ca0c, 32'hc24475dc};
test_output[3154] = '{32'h42720cab};
test_index[3154] = '{5};
test_input[25240:25247] = '{32'h4222df82, 32'hc293d8c2, 32'hc0c88a8d, 32'h42bdc452, 32'h3f8eae28, 32'h41a93592, 32'hc19f7b0e, 32'hc1bd7f4f};
test_output[3155] = '{32'h42bdc452};
test_index[3155] = '{3};
test_input[25248:25255] = '{32'hc2a69941, 32'hc2a19d2d, 32'hc1ee9608, 32'h42232a50, 32'hc16568fa, 32'hc1f38bba, 32'hc2932834, 32'hc2b95df6};
test_output[3156] = '{32'h42232a50};
test_index[3156] = '{3};
test_input[25256:25263] = '{32'hbfb6469c, 32'hc2ac16d5, 32'h4228993e, 32'hc2329daf, 32'hc2b2561f, 32'h42c28fa7, 32'hc1f440ff, 32'hc16ca3e5};
test_output[3157] = '{32'h42c28fa7};
test_index[3157] = '{5};
test_input[25264:25271] = '{32'hc1c2a0b0, 32'hc1d20fe9, 32'hc2799bd2, 32'hc21f5764, 32'h42c2fe58, 32'h42914778, 32'h42648081, 32'hc209e09e};
test_output[3158] = '{32'h42c2fe58};
test_index[3158] = '{4};
test_input[25272:25279] = '{32'h429a2e28, 32'h42c22c8d, 32'hc2a9d6d8, 32'h408226a9, 32'h4298acd2, 32'h4262b43a, 32'h41c0f47c, 32'hc2a83334};
test_output[3159] = '{32'h42c22c8d};
test_index[3159] = '{1};
test_input[25280:25287] = '{32'h4247e485, 32'hc1e94826, 32'h41bab625, 32'h42759d9c, 32'hc2abf4c4, 32'hc25b61c7, 32'h427d8b6f, 32'hc2317739};
test_output[3160] = '{32'h427d8b6f};
test_index[3160] = '{6};
test_input[25288:25295] = '{32'h42900dbd, 32'h41812abf, 32'hc1d83f57, 32'hc2b66fd7, 32'h42aeced4, 32'hc277cddf, 32'h429377ab, 32'h42802965};
test_output[3161] = '{32'h42aeced4};
test_index[3161] = '{4};
test_input[25296:25303] = '{32'hc1bc37e5, 32'hc1344bb6, 32'hc220933f, 32'h41b966dd, 32'hc2b5276c, 32'hc2c5c469, 32'hc2c37752, 32'h4289dd8e};
test_output[3162] = '{32'h4289dd8e};
test_index[3162] = '{7};
test_input[25304:25311] = '{32'h41d3039c, 32'hc1f3be14, 32'hc2b1da94, 32'h42a27b03, 32'hc2157174, 32'h41be5d97, 32'h4279c59e, 32'h42b3aa8f};
test_output[3163] = '{32'h42b3aa8f};
test_index[3163] = '{7};
test_input[25312:25319] = '{32'h41545d0c, 32'h42372918, 32'h4006f6f3, 32'h423393f5, 32'h42ba3b97, 32'h41a3de51, 32'h42c5ba6e, 32'h411451fb};
test_output[3164] = '{32'h42c5ba6e};
test_index[3164] = '{6};
test_input[25320:25327] = '{32'h4238336b, 32'hc19da147, 32'hc2343acc, 32'h42bb0e27, 32'h41c5bd43, 32'h426eb00a, 32'hc1ceb4f4, 32'hc28c1cf5};
test_output[3165] = '{32'h42bb0e27};
test_index[3165] = '{3};
test_input[25328:25335] = '{32'hc185ae41, 32'hc2543d38, 32'h428a36f6, 32'h4156a068, 32'hc2a02ca0, 32'hc1335de1, 32'hc1f2c356, 32'h420bbeae};
test_output[3166] = '{32'h428a36f6};
test_index[3166] = '{2};
test_input[25336:25343] = '{32'hc250033f, 32'hc253f350, 32'hc14f0af3, 32'h419867b1, 32'h4239302b, 32'h4284267c, 32'hc2706dfc, 32'hbfa25833};
test_output[3167] = '{32'h4284267c};
test_index[3167] = '{5};
test_input[25344:25351] = '{32'hc2c7459d, 32'h41c0cff8, 32'h427f39d5, 32'h4266fecf, 32'h42341a24, 32'hc26751b2, 32'h42519392, 32'hc28cdd24};
test_output[3168] = '{32'h427f39d5};
test_index[3168] = '{2};
test_input[25352:25359] = '{32'hc29e21f9, 32'h40ac9c8f, 32'hc2986ca6, 32'hc1cf24f8, 32'hc19471d9, 32'hc155b89b, 32'hc1dd6cb5, 32'hc28b68fb};
test_output[3169] = '{32'h40ac9c8f};
test_index[3169] = '{1};
test_input[25360:25367] = '{32'hc2a3968b, 32'h41cc5fd5, 32'hc14769e7, 32'h416e7271, 32'h42776022, 32'h411b38c7, 32'hc1ce56b0, 32'hc28fe21f};
test_output[3170] = '{32'h42776022};
test_index[3170] = '{4};
test_input[25368:25375] = '{32'hc2210ddc, 32'hc19f0c96, 32'h42c610e5, 32'h413fd14a, 32'h4288fbff, 32'hc29e9176, 32'h4200373c, 32'hc1e0e2d3};
test_output[3171] = '{32'h42c610e5};
test_index[3171] = '{2};
test_input[25376:25383] = '{32'hc1edae94, 32'hc02e07c1, 32'h42935d16, 32'hc2c61beb, 32'h42ae2aac, 32'h42c271ac, 32'hc11eef1e, 32'hc267b8e7};
test_output[3172] = '{32'h42c271ac};
test_index[3172] = '{5};
test_input[25384:25391] = '{32'hc1682e5b, 32'hc1b8028a, 32'hc1af74f2, 32'h42b5681c, 32'hc030bd58, 32'h401f9623, 32'hc0d76dba, 32'h42a1d681};
test_output[3173] = '{32'h42b5681c};
test_index[3173] = '{3};
test_input[25392:25399] = '{32'h428ad5d9, 32'hc22ce0fe, 32'hc284956b, 32'h42677bc4, 32'hc2582567, 32'hc2052468, 32'hc2b49647, 32'hc23798cc};
test_output[3174] = '{32'h428ad5d9};
test_index[3174] = '{0};
test_input[25400:25407] = '{32'hc28314bf, 32'h42063823, 32'hc2860171, 32'hc2a1c0f3, 32'h420c2258, 32'h4263e035, 32'hc1f088dc, 32'h42768ad6};
test_output[3175] = '{32'h42768ad6};
test_index[3175] = '{7};
test_input[25408:25415] = '{32'hc29e15eb, 32'hc2a80388, 32'hc21a9259, 32'hc24e0c2e, 32'hc2c23810, 32'hc2a8af94, 32'h40a9dffc, 32'hc1d4e1b3};
test_output[3176] = '{32'h40a9dffc};
test_index[3176] = '{6};
test_input[25416:25423] = '{32'h41bb1169, 32'hc1872bb0, 32'hc12e6926, 32'hc2a57596, 32'hc20162dc, 32'hc2b98a42, 32'h4204e6ca, 32'hc2c21edf};
test_output[3177] = '{32'h4204e6ca};
test_index[3177] = '{6};
test_input[25424:25431] = '{32'hc1f8dce7, 32'h41f26c1b, 32'h426de733, 32'h420d1fdb, 32'h42301d59, 32'hc2b68df0, 32'hc2bbe114, 32'hc2492512};
test_output[3178] = '{32'h426de733};
test_index[3178] = '{2};
test_input[25432:25439] = '{32'hc22f2aaa, 32'h42b529e5, 32'hc144a500, 32'hc2a5e2ac, 32'hc1cbf0ee, 32'hc2a933e1, 32'hc23bad76, 32'h428d5aef};
test_output[3179] = '{32'h42b529e5};
test_index[3179] = '{1};
test_input[25440:25447] = '{32'hc00b1873, 32'h41d62b40, 32'hc240d125, 32'h405cb915, 32'h424af831, 32'hc098c308, 32'h42379ec7, 32'h42b06253};
test_output[3180] = '{32'h42b06253};
test_index[3180] = '{7};
test_input[25448:25455] = '{32'h42be5893, 32'h3fe94323, 32'hc2c04e2b, 32'h424e66a6, 32'h428c1c5a, 32'h42c31a53, 32'hc28b84cf, 32'h42aad810};
test_output[3181] = '{32'h42c31a53};
test_index[3181] = '{5};
test_input[25456:25463] = '{32'h408eaba2, 32'hc2b970cc, 32'h428c1c03, 32'hc1c251ea, 32'h41af2d0e, 32'h42043e33, 32'h42339608, 32'h4274a3be};
test_output[3182] = '{32'h428c1c03};
test_index[3182] = '{2};
test_input[25464:25471] = '{32'hc143d7bd, 32'hc226ee8e, 32'hc2a5f53f, 32'hc1b26a84, 32'h4184f87b, 32'hc2051a84, 32'h41d7bf02, 32'hc275307b};
test_output[3183] = '{32'h41d7bf02};
test_index[3183] = '{6};
test_input[25472:25479] = '{32'h4280b109, 32'h42b2b745, 32'h423749ac, 32'h4160c0df, 32'h4145bda2, 32'h42717196, 32'h420084e3, 32'h429145b6};
test_output[3184] = '{32'h42b2b745};
test_index[3184] = '{1};
test_input[25480:25487] = '{32'h425ab813, 32'hc2320903, 32'h429cd7a0, 32'hc22acb6a, 32'hc29fd771, 32'h42c551b1, 32'hc17b30d4, 32'hc174b6c8};
test_output[3185] = '{32'h42c551b1};
test_index[3185] = '{5};
test_input[25488:25495] = '{32'h42ab61a8, 32'h4285d5ad, 32'h412d963d, 32'h4262cf31, 32'hc1f77af5, 32'hc1eadff6, 32'h42c5e9e4, 32'h4275cd6a};
test_output[3186] = '{32'h42c5e9e4};
test_index[3186] = '{6};
test_input[25496:25503] = '{32'hc1231378, 32'h420a76dc, 32'hc22f8ed5, 32'hc1d136d8, 32'h427161c3, 32'hc2968716, 32'hc24a4d43, 32'h41785b91};
test_output[3187] = '{32'h427161c3};
test_index[3187] = '{4};
test_input[25504:25511] = '{32'hc294c48f, 32'hc17ee150, 32'hc1e5a1a9, 32'h42beacf6, 32'h420ff086, 32'hc25333fa, 32'h42a1e738, 32'h4210d13e};
test_output[3188] = '{32'h42beacf6};
test_index[3188] = '{3};
test_input[25512:25519] = '{32'h423367ed, 32'hc10b9880, 32'hc218871b, 32'h4261c8df, 32'h4232caca, 32'h40b17317, 32'hc101b4ee, 32'hc2ba5554};
test_output[3189] = '{32'h4261c8df};
test_index[3189] = '{3};
test_input[25520:25527] = '{32'hc2c0705a, 32'h4200c0bc, 32'h4282bf05, 32'h42165712, 32'hc2b99a40, 32'h410f9036, 32'hc269111d, 32'hc1ca0dd8};
test_output[3190] = '{32'h4282bf05};
test_index[3190] = '{2};
test_input[25528:25535] = '{32'h41209af1, 32'hc184f35f, 32'hc1f0fa78, 32'hc20f455e, 32'hc287e948, 32'hc268075d, 32'h42b7f5e2, 32'h420ad13e};
test_output[3191] = '{32'h42b7f5e2};
test_index[3191] = '{6};
test_input[25536:25543] = '{32'h42aa4438, 32'hc229395a, 32'hc27c3134, 32'hc2952d8e, 32'h4244b8fa, 32'hc25621fc, 32'h42c35098, 32'h42361e5b};
test_output[3192] = '{32'h42c35098};
test_index[3192] = '{6};
test_input[25544:25551] = '{32'h4093daf2, 32'h4175dbb6, 32'h42abf18e, 32'hc2b74db1, 32'h42183a55, 32'h41a6f52e, 32'hc2549a36, 32'hc1a35e01};
test_output[3193] = '{32'h42abf18e};
test_index[3193] = '{2};
test_input[25552:25559] = '{32'h42c3a02e, 32'h42bd7317, 32'h427b1bed, 32'hc2b4f8c5, 32'hc29a0f72, 32'h42519fe1, 32'hc23c94da, 32'hc28220d5};
test_output[3194] = '{32'h42c3a02e};
test_index[3194] = '{0};
test_input[25560:25567] = '{32'h41fc8195, 32'hc1ccfcb6, 32'h426fd8b4, 32'hc1993264, 32'h41f0dddb, 32'hc2aca9f6, 32'hc28d3e3a, 32'hc1c2f117};
test_output[3195] = '{32'h426fd8b4};
test_index[3195] = '{2};
test_input[25568:25575] = '{32'hc2c2cd85, 32'h42c6c264, 32'h420c8b77, 32'hc27d338e, 32'hc2b2558d, 32'h41fad979, 32'hc269856f, 32'hc1f21b51};
test_output[3196] = '{32'h42c6c264};
test_index[3196] = '{1};
test_input[25576:25583] = '{32'h4286a21f, 32'h41b327aa, 32'hc2ac52d8, 32'h4280293f, 32'h42bd80fa, 32'hc16b2638, 32'h424477c2, 32'h41e53ee2};
test_output[3197] = '{32'h42bd80fa};
test_index[3197] = '{4};
test_input[25584:25591] = '{32'hc24161bc, 32'hc2568b71, 32'hc28be33c, 32'h42c0d561, 32'hc286c6bd, 32'h42a8e22b, 32'hc2542162, 32'h4128eaa8};
test_output[3198] = '{32'h42c0d561};
test_index[3198] = '{3};
test_input[25592:25599] = '{32'h4190a181, 32'h420504be, 32'h42425f76, 32'h42277226, 32'hc2102068, 32'h40aa11eb, 32'hc21b24dc, 32'hc2467064};
test_output[3199] = '{32'h42425f76};
test_index[3199] = '{2};
test_input[25600:25607] = '{32'hc1e019fc, 32'hc2a80b23, 32'h429040a6, 32'h420b99bb, 32'h42ae7aff, 32'h420e73f4, 32'h41a4a92f, 32'hc28f8319};
test_output[3200] = '{32'h42ae7aff};
test_index[3200] = '{4};
test_input[25608:25615] = '{32'h41cbed0e, 32'hc254b6c9, 32'h4296b0fa, 32'hc2b4589b, 32'h4269e59d, 32'hc285f511, 32'hc28b08e3, 32'hc199ab6b};
test_output[3201] = '{32'h4296b0fa};
test_index[3201] = '{2};
test_input[25616:25623] = '{32'h4294c921, 32'h4284e8e5, 32'hc1893e80, 32'h41081555, 32'hc2588a0f, 32'hc0cb16c6, 32'hc21aebc3, 32'h42c138fc};
test_output[3202] = '{32'h42c138fc};
test_index[3202] = '{7};
test_input[25624:25631] = '{32'hc29c3c26, 32'hc1744ff0, 32'hc2802f6d, 32'hc1dc1ca5, 32'hc29e3d67, 32'h41d328cb, 32'hc282e113, 32'h42958756};
test_output[3203] = '{32'h42958756};
test_index[3203] = '{7};
test_input[25632:25639] = '{32'hc204c9d0, 32'hc2474333, 32'h408b3741, 32'h42a8f97c, 32'h419759e2, 32'hc283bb15, 32'hc192410f, 32'hc00afc42};
test_output[3204] = '{32'h42a8f97c};
test_index[3204] = '{3};
test_input[25640:25647] = '{32'hc20b43a2, 32'hc1f3ec4c, 32'h429a5def, 32'hc20ee873, 32'hc28bdcb8, 32'h41d616f1, 32'h41fe2ede, 32'hc01687cb};
test_output[3205] = '{32'h429a5def};
test_index[3205] = '{2};
test_input[25648:25655] = '{32'hc25a7f50, 32'hbf035277, 32'h428abdc0, 32'h41a09218, 32'hc2b77f9d, 32'h4243b9fc, 32'hc1a41a15, 32'hc2208a87};
test_output[3206] = '{32'h428abdc0};
test_index[3206] = '{2};
test_input[25656:25663] = '{32'hc211ebfc, 32'h42c6f55e, 32'h3f352adb, 32'h4294adfa, 32'h429ea2ca, 32'h42beb62b, 32'hc243ff26, 32'hc2ad5116};
test_output[3207] = '{32'h42c6f55e};
test_index[3207] = '{1};
test_input[25664:25671] = '{32'hc228818a, 32'hc1a4fea1, 32'hc2a17d7b, 32'h42089c22, 32'h422dc5e3, 32'hc03aa107, 32'hc2877699, 32'hc26558bb};
test_output[3208] = '{32'h422dc5e3};
test_index[3208] = '{4};
test_input[25672:25679] = '{32'hc171fd57, 32'h42072ace, 32'h418a41d7, 32'h4265d6b1, 32'hc2b2eae1, 32'hc2835c4f, 32'hc2a1e2a6, 32'hc2bc9980};
test_output[3209] = '{32'h4265d6b1};
test_index[3209] = '{3};
test_input[25680:25687] = '{32'h425d6287, 32'h426af077, 32'h42b5498f, 32'hc1d02268, 32'hc21c582f, 32'hc2bf467c, 32'hc212ab68, 32'h42a2a265};
test_output[3210] = '{32'h42b5498f};
test_index[3210] = '{2};
test_input[25688:25695] = '{32'h41c4e7eb, 32'h41afe761, 32'hc192fb11, 32'hc130dc89, 32'hc2be1f71, 32'hc090deff, 32'h4200543b, 32'hc296242d};
test_output[3211] = '{32'h4200543b};
test_index[3211] = '{6};
test_input[25696:25703] = '{32'h428398f3, 32'hc294e726, 32'h3fc77a6a, 32'hc1591e20, 32'h42a430f7, 32'hc1b8619c, 32'hc192811a, 32'h42b30eed};
test_output[3212] = '{32'h42b30eed};
test_index[3212] = '{7};
test_input[25704:25711] = '{32'hc299a914, 32'hc1c19b7e, 32'h42a76b6d, 32'h417a672b, 32'h42c3c28c, 32'h416afa75, 32'hc1f9ece1, 32'h40cd80c1};
test_output[3213] = '{32'h42c3c28c};
test_index[3213] = '{4};
test_input[25712:25719] = '{32'h429b9502, 32'hc23c6ee9, 32'h40a6e06a, 32'h42896aa4, 32'hc29fe25d, 32'hc22f7e6e, 32'hc2b0e72c, 32'h42b15220};
test_output[3214] = '{32'h42b15220};
test_index[3214] = '{7};
test_input[25720:25727] = '{32'hc266cc49, 32'h42462413, 32'hc2a26344, 32'hc21d53e3, 32'hc15383b3, 32'hc2ae6a93, 32'h3fc57888, 32'hc2574eca};
test_output[3215] = '{32'h42462413};
test_index[3215] = '{1};
test_input[25728:25735] = '{32'h42843f2d, 32'hc2b4585d, 32'hc13757b2, 32'h4201d164, 32'hc13e510b, 32'hc2aac9e4, 32'h424e9d91, 32'h4290bf35};
test_output[3216] = '{32'h4290bf35};
test_index[3216] = '{7};
test_input[25736:25743] = '{32'h423d8457, 32'hc2594a57, 32'hc209792d, 32'h42b1b72d, 32'hc26ba57d, 32'h42a7f6fe, 32'hc1d68195, 32'h4119bcdd};
test_output[3217] = '{32'h42b1b72d};
test_index[3217] = '{3};
test_input[25744:25751] = '{32'h428ebd8b, 32'h42872a6e, 32'hc265f9ae, 32'h42051778, 32'hc1461dc5, 32'hc24e31e3, 32'h41e844d3, 32'h41fc9b3f};
test_output[3218] = '{32'h428ebd8b};
test_index[3218] = '{0};
test_input[25752:25759] = '{32'hc25c724f, 32'hc2a68160, 32'hc199c706, 32'h422cb415, 32'hc209134d, 32'h42a8c6e3, 32'hc23a52a8, 32'h4231c540};
test_output[3219] = '{32'h42a8c6e3};
test_index[3219] = '{5};
test_input[25760:25767] = '{32'h41a09b19, 32'h424e3513, 32'h422475be, 32'h3f6fc3fd, 32'h4255dd19, 32'hc10bb1b7, 32'h42b50f4d, 32'h42420d4a};
test_output[3220] = '{32'h42b50f4d};
test_index[3220] = '{6};
test_input[25768:25775] = '{32'h3fabe865, 32'h411d4b0a, 32'hc29dffa5, 32'h4213c1c4, 32'h42bac815, 32'h4262cbd2, 32'hc291dc34, 32'hc2553713};
test_output[3221] = '{32'h42bac815};
test_index[3221] = '{4};
test_input[25776:25783] = '{32'h4242efe1, 32'hc2b37f3e, 32'hc0c354e4, 32'h423aa531, 32'h41e8fb13, 32'hc246a2e2, 32'h425da7f6, 32'hbeb05fbf};
test_output[3222] = '{32'h425da7f6};
test_index[3222] = '{6};
test_input[25784:25791] = '{32'hc2be87e0, 32'hc2b90ee1, 32'hc2906108, 32'hc2b5ab45, 32'hc2a93a6b, 32'h42b19500, 32'hc1075d7f, 32'hc237b7f4};
test_output[3223] = '{32'h42b19500};
test_index[3223] = '{5};
test_input[25792:25799] = '{32'h427f3f61, 32'h42c7e1ba, 32'hc207fcdc, 32'h4290b72b, 32'h4244b4f7, 32'hc2a181d3, 32'h423e48c1, 32'h408465c1};
test_output[3224] = '{32'h42c7e1ba};
test_index[3224] = '{1};
test_input[25800:25807] = '{32'hc19af949, 32'hc2395a24, 32'h42b78f5d, 32'h426e3e42, 32'hc1a7cced, 32'h42c2b44f, 32'h42315b90, 32'h42a80d83};
test_output[3225] = '{32'h42c2b44f};
test_index[3225] = '{5};
test_input[25808:25815] = '{32'h425b8a91, 32'h40f91d3b, 32'h4241ab83, 32'h41e83490, 32'h40edbb2d, 32'h41b0ada2, 32'h413f39bd, 32'hc25f9442};
test_output[3226] = '{32'h425b8a91};
test_index[3226] = '{0};
test_input[25816:25823] = '{32'h42304436, 32'hc1556fe1, 32'h41f72141, 32'h40526b2e, 32'hc25d13d3, 32'hc29c8962, 32'hc22d6d59, 32'h4198123c};
test_output[3227] = '{32'h42304436};
test_index[3227] = '{0};
test_input[25824:25831] = '{32'h429d09e9, 32'hc1f83204, 32'h4270fa65, 32'h42942ac6, 32'hc09aeca6, 32'hc057e99d, 32'h42b8d566, 32'hc26ff3f6};
test_output[3228] = '{32'h42b8d566};
test_index[3228] = '{6};
test_input[25832:25839] = '{32'h42ade58e, 32'hc28591a9, 32'h3fdc44e9, 32'hc292c6cd, 32'h42582b4e, 32'hc2adac65, 32'hc28ed14e, 32'h418747db};
test_output[3229] = '{32'h42ade58e};
test_index[3229] = '{0};
test_input[25840:25847] = '{32'hc29874ef, 32'hc2a212d2, 32'hc08216e6, 32'h420e685f, 32'h425f5481, 32'h41f40b88, 32'hc1079263, 32'hc06c477c};
test_output[3230] = '{32'h425f5481};
test_index[3230] = '{4};
test_input[25848:25855] = '{32'hc2a4d5da, 32'hc0fc6e39, 32'h42bd040d, 32'h3e896a1f, 32'h42a0a5f6, 32'h4264f629, 32'hc2aca8da, 32'h4251ee19};
test_output[3231] = '{32'h42bd040d};
test_index[3231] = '{2};
test_input[25856:25863] = '{32'h426524f5, 32'hc256d574, 32'hc2944380, 32'h4207e227, 32'hc237ab64, 32'hc1149dc2, 32'h41db4149, 32'h42b464d4};
test_output[3232] = '{32'h42b464d4};
test_index[3232] = '{7};
test_input[25864:25871] = '{32'hc223f215, 32'hc25bbc7a, 32'h42b72d13, 32'hc189dcf3, 32'hc2bc37de, 32'hc2bfdede, 32'h422b7919, 32'h40800f9f};
test_output[3233] = '{32'h42b72d13};
test_index[3233] = '{2};
test_input[25872:25879] = '{32'h42363afe, 32'hc20b785d, 32'hc18ba9a3, 32'h42c29857, 32'h429fc54a, 32'hc259986e, 32'h429e02c0, 32'hc285a652};
test_output[3234] = '{32'h42c29857};
test_index[3234] = '{3};
test_input[25880:25887] = '{32'h428425c2, 32'h41b3807c, 32'h42883ff5, 32'hc10658f0, 32'hc2a38722, 32'h4285a2d2, 32'h42c65b12, 32'h42acb416};
test_output[3235] = '{32'h42c65b12};
test_index[3235] = '{6};
test_input[25888:25895] = '{32'hc1c4e7d6, 32'hc2c77a34, 32'h42888292, 32'h42bcc295, 32'h4282327e, 32'hc28d3b68, 32'h41f0124f, 32'hc196c1e9};
test_output[3236] = '{32'h42bcc295};
test_index[3236] = '{3};
test_input[25896:25903] = '{32'hc2b3f6ce, 32'h4240bed4, 32'hc08c39be, 32'hc13e8d24, 32'h42bfd777, 32'h42623cae, 32'hc2af4ba6, 32'h4194ef4c};
test_output[3237] = '{32'h42bfd777};
test_index[3237] = '{4};
test_input[25904:25911] = '{32'h425e3450, 32'hc0094a96, 32'h422acab2, 32'h4278de12, 32'h419198fc, 32'hc21be1c2, 32'hc10599a2, 32'h426b0cc2};
test_output[3238] = '{32'h4278de12};
test_index[3238] = '{3};
test_input[25912:25919] = '{32'h42b8880c, 32'hc0795ebc, 32'hc2c3df43, 32'hc12d21a9, 32'hc2b584fd, 32'h42389f91, 32'h40ae83c3, 32'hc2157cc6};
test_output[3239] = '{32'h42b8880c};
test_index[3239] = '{0};
test_input[25920:25927] = '{32'h42b1bafb, 32'hc2a3017c, 32'h4214f167, 32'hc28d36db, 32'h4166d1ff, 32'h42a0da3c, 32'hc11cf478, 32'hc2a28cfb};
test_output[3240] = '{32'h42b1bafb};
test_index[3240] = '{0};
test_input[25928:25935] = '{32'h425fab91, 32'hc2ac5238, 32'hc212592b, 32'h4229d0b2, 32'hc1949220, 32'hc26376a8, 32'h429b0cdf, 32'h3fdaf806};
test_output[3241] = '{32'h429b0cdf};
test_index[3241] = '{6};
test_input[25936:25943] = '{32'hc26565c3, 32'h42b1e36b, 32'h41ebd57e, 32'hc288334c, 32'h429e8f9e, 32'hc28a2cfe, 32'hc290c8cc, 32'h4280e9ac};
test_output[3242] = '{32'h42b1e36b};
test_index[3242] = '{1};
test_input[25944:25951] = '{32'hc25bf37e, 32'h424afe11, 32'h42728a8f, 32'hc1477955, 32'h402bea05, 32'h42bb5bcf, 32'h4253e543, 32'hc2bce259};
test_output[3243] = '{32'h42bb5bcf};
test_index[3243] = '{5};
test_input[25952:25959] = '{32'h424df3bf, 32'h4040736a, 32'hc293c38e, 32'h41d480ae, 32'h42a9614f, 32'hc195e10c, 32'h42875a7b, 32'hc2b0b284};
test_output[3244] = '{32'h42a9614f};
test_index[3244] = '{4};
test_input[25960:25967] = '{32'hc28a1089, 32'h42564001, 32'h415146c6, 32'h42b4eeca, 32'hc2834bc6, 32'h41997fc5, 32'h41b29148, 32'h42a0bcbd};
test_output[3245] = '{32'h42b4eeca};
test_index[3245] = '{3};
test_input[25968:25975] = '{32'hc1c576ea, 32'hc170575b, 32'hc0e52e75, 32'h41996473, 32'hc2bc52be, 32'h417d383e, 32'h426a7e28, 32'hc25dad61};
test_output[3246] = '{32'h426a7e28};
test_index[3246] = '{6};
test_input[25976:25983] = '{32'hc25d6baa, 32'h426f630b, 32'hc22b0891, 32'h414f409c, 32'h42403ef0, 32'h42b26198, 32'hc218b768, 32'h429cad09};
test_output[3247] = '{32'h42b26198};
test_index[3247] = '{5};
test_input[25984:25991] = '{32'hc2bb59b1, 32'hc2898fc9, 32'hc1995e19, 32'h429c49b2, 32'h42c77d7f, 32'h4194ad8a, 32'hc1aeae6b, 32'hc21bff1d};
test_output[3248] = '{32'h42c77d7f};
test_index[3248] = '{4};
test_input[25992:25999] = '{32'hc270ff3b, 32'hc18ba34f, 32'h427602ca, 32'hc263e177, 32'h42a22640, 32'hc178bd0d, 32'hc2b5c166, 32'hc211f0d3};
test_output[3249] = '{32'h42a22640};
test_index[3249] = '{4};
test_input[26000:26007] = '{32'hc1705ba1, 32'hc292a936, 32'h41456e31, 32'hc126f97f, 32'h41e96a19, 32'h42a1594a, 32'h41a8f63c, 32'h42a3e27d};
test_output[3250] = '{32'h42a3e27d};
test_index[3250] = '{7};
test_input[26008:26015] = '{32'hc26816b8, 32'h42877649, 32'hc25fd813, 32'h428e0512, 32'hc21eb739, 32'hc23528ac, 32'hc2b75755, 32'hc23d2bdd};
test_output[3251] = '{32'h428e0512};
test_index[3251] = '{3};
test_input[26016:26023] = '{32'h42b9c284, 32'hc1605aaf, 32'h426022b5, 32'h42195a53, 32'hc2016866, 32'h42694d68, 32'h4299bac7, 32'h42872360};
test_output[3252] = '{32'h42b9c284};
test_index[3252] = '{0};
test_input[26024:26031] = '{32'h429d45dc, 32'h42815e8e, 32'h42b5b2fd, 32'hc26275b6, 32'h41e74f20, 32'hc249d7ef, 32'h4093e957, 32'h423f6679};
test_output[3253] = '{32'h42b5b2fd};
test_index[3253] = '{2};
test_input[26032:26039] = '{32'h4293a661, 32'h42a3af18, 32'h42479a4d, 32'hc13336ff, 32'h42940388, 32'h40804d0a, 32'h42516dbc, 32'h41dddbe5};
test_output[3254] = '{32'h42a3af18};
test_index[3254] = '{1};
test_input[26040:26047] = '{32'h4193d9bf, 32'hc223c22e, 32'hc2ab44ef, 32'h42bd259d, 32'hc2848e49, 32'h41f07535, 32'hc21a9648, 32'h426cc264};
test_output[3255] = '{32'h42bd259d};
test_index[3255] = '{3};
test_input[26048:26055] = '{32'h4293e49f, 32'hc2115067, 32'hc2a83599, 32'hc2be134c, 32'hc2a646f2, 32'h4205f396, 32'hc28e6941, 32'h42a0bcac};
test_output[3256] = '{32'h42a0bcac};
test_index[3256] = '{7};
test_input[26056:26063] = '{32'h42358d5c, 32'h418d4de4, 32'hc1f5161d, 32'hc29787d2, 32'hc1a73e65, 32'hc0a8ac98, 32'h42b27505, 32'hc114b6e0};
test_output[3257] = '{32'h42b27505};
test_index[3257] = '{6};
test_input[26064:26071] = '{32'hc19f4b5f, 32'h42969010, 32'h42627c00, 32'h425f564e, 32'hc27d4b66, 32'h42138849, 32'hc2b08875, 32'h412eb709};
test_output[3258] = '{32'h42969010};
test_index[3258] = '{1};
test_input[26072:26079] = '{32'hc12814f5, 32'h410106fc, 32'hc1efc931, 32'hc18e55ac, 32'hc2b303e2, 32'hc23c5df7, 32'hc2958a53, 32'h42201cc9};
test_output[3259] = '{32'h42201cc9};
test_index[3259] = '{7};
test_input[26080:26087] = '{32'h4213d8d1, 32'h42b1e1c5, 32'hc00e01c9, 32'hc26b6cf5, 32'h42211d37, 32'h42bc0d51, 32'h41810a11, 32'h42210503};
test_output[3260] = '{32'h42bc0d51};
test_index[3260] = '{5};
test_input[26088:26095] = '{32'h4231e63f, 32'hc1d1f262, 32'h4113d965, 32'h420995af, 32'hc21e7e3d, 32'h42b57fa6, 32'h414f6d49, 32'h420d00e1};
test_output[3261] = '{32'h42b57fa6};
test_index[3261] = '{5};
test_input[26096:26103] = '{32'hc0caa633, 32'h424b3510, 32'hc1cbafae, 32'h4254f288, 32'h411fd6a6, 32'hc278ab8a, 32'h42382516, 32'hc17a3f0d};
test_output[3262] = '{32'h4254f288};
test_index[3262] = '{3};
test_input[26104:26111] = '{32'h3fcbca13, 32'hc24dae6f, 32'h41ece921, 32'hc2c4bf21, 32'hc0c88646, 32'hc19da633, 32'hc210f8fc, 32'hc1827c1d};
test_output[3263] = '{32'h41ece921};
test_index[3263] = '{2};
test_input[26112:26119] = '{32'hc2ad2f6c, 32'hc2c759b6, 32'hc2c3baa0, 32'h4226b0d1, 32'h4149509a, 32'h41b85747, 32'h429d57ee, 32'h423a913c};
test_output[3264] = '{32'h429d57ee};
test_index[3264] = '{6};
test_input[26120:26127] = '{32'hc10aac07, 32'h408166d6, 32'h42b033cc, 32'h42c20c34, 32'hc12640aa, 32'h4231f641, 32'h42c63502, 32'hc0b9b7a4};
test_output[3265] = '{32'h42c63502};
test_index[3265] = '{6};
test_input[26128:26135] = '{32'h41ff3ce9, 32'hc28081ef, 32'h41f59342, 32'hc17de5d2, 32'h3f1ccf47, 32'hc2382bf8, 32'h414ffe38, 32'h40c6afb6};
test_output[3266] = '{32'h41ff3ce9};
test_index[3266] = '{0};
test_input[26136:26143] = '{32'h42b74e5a, 32'hc293d175, 32'h4248e5f3, 32'hbff10784, 32'h42b788e3, 32'h42bbf414, 32'hc27b9dc4, 32'h41dd5cf3};
test_output[3267] = '{32'h42bbf414};
test_index[3267] = '{5};
test_input[26144:26151] = '{32'h41da94e8, 32'h42b0531b, 32'hc23fcfdb, 32'h4214f3f5, 32'h40375f93, 32'hc1b36302, 32'h41ebadfb, 32'h42928348};
test_output[3268] = '{32'h42b0531b};
test_index[3268] = '{1};
test_input[26152:26159] = '{32'hc120c266, 32'h428f5c30, 32'hc2b5fe40, 32'hc2902292, 32'hc2280e20, 32'h4285ba61, 32'h425cc729, 32'h4239b697};
test_output[3269] = '{32'h428f5c30};
test_index[3269] = '{1};
test_input[26160:26167] = '{32'h40eb8006, 32'h429216cf, 32'hc2933fb3, 32'hc257c0f7, 32'hc14ec821, 32'hc1e2bf76, 32'hc22dc603, 32'h412f5965};
test_output[3270] = '{32'h429216cf};
test_index[3270] = '{1};
test_input[26168:26175] = '{32'hc1390b53, 32'hc2c0b8f9, 32'h41edbe65, 32'hc13bb611, 32'h4294b7e0, 32'hc2a92f1a, 32'hc2acaca2, 32'hc10f1f5d};
test_output[3271] = '{32'h4294b7e0};
test_index[3271] = '{4};
test_input[26176:26183] = '{32'h425f6492, 32'h40c5ce06, 32'hc29ec079, 32'hc2942c60, 32'h414fc75a, 32'h422031e8, 32'hc15916df, 32'hc2af9820};
test_output[3272] = '{32'h425f6492};
test_index[3272] = '{0};
test_input[26184:26191] = '{32'h417012c9, 32'hc13617c3, 32'hc28096ea, 32'h4153e011, 32'hc288c66b, 32'h426a32b8, 32'hc275c9fb, 32'hc2385fbe};
test_output[3273] = '{32'h426a32b8};
test_index[3273] = '{5};
test_input[26192:26199] = '{32'hc00c76b2, 32'hbfa07009, 32'h429c41ae, 32'h425ff9b7, 32'hc2b16cd0, 32'hc29bb357, 32'h42aa895c, 32'h4256646d};
test_output[3274] = '{32'h42aa895c};
test_index[3274] = '{6};
test_input[26200:26207] = '{32'hc274136b, 32'hc20d8d9e, 32'hc2932cef, 32'hc21ab26c, 32'h42830cf9, 32'hc215dd5b, 32'hc2c11e8f, 32'hc0b09722};
test_output[3275] = '{32'h42830cf9};
test_index[3275] = '{4};
test_input[26208:26215] = '{32'hc2350dde, 32'hc23c1847, 32'h42ab50a3, 32'hc2971466, 32'h400a1436, 32'hc1877ee5, 32'hc28eb31a, 32'hc105082f};
test_output[3276] = '{32'h42ab50a3};
test_index[3276] = '{2};
test_input[26216:26223] = '{32'hc28d807e, 32'h4252ced4, 32'hc21f42c3, 32'h4292fa6d, 32'h424189d0, 32'h412e8fe9, 32'hc23484a2, 32'h40751021};
test_output[3277] = '{32'h4292fa6d};
test_index[3277] = '{3};
test_input[26224:26231] = '{32'h427867ab, 32'h429d32fa, 32'h42bb3abf, 32'hc1e08bdf, 32'h420e9773, 32'h4238dc95, 32'h41c7817f, 32'hc1ba5c96};
test_output[3278] = '{32'h42bb3abf};
test_index[3278] = '{2};
test_input[26232:26239] = '{32'hc2c2ecaa, 32'h42b31d83, 32'hc2b68a2f, 32'h41cbb815, 32'h40118fea, 32'hc2937ce7, 32'hc287bf8a, 32'hc2ab365f};
test_output[3279] = '{32'h42b31d83};
test_index[3279] = '{1};
test_input[26240:26247] = '{32'hc2471303, 32'h4283e870, 32'h418bbd70, 32'h41a90622, 32'h422b9e6e, 32'hc1886700, 32'h421eb5fd, 32'h4219d4b9};
test_output[3280] = '{32'h4283e870};
test_index[3280] = '{1};
test_input[26248:26255] = '{32'h410c895d, 32'hc17b6bb4, 32'h42b1723d, 32'h42039815, 32'hc29ba14e, 32'h428be859, 32'hc287cd98, 32'hc12bc829};
test_output[3281] = '{32'h42b1723d};
test_index[3281] = '{2};
test_input[26256:26263] = '{32'hc2b3a013, 32'h42ae5b74, 32'h40007472, 32'hc0ff705f, 32'hc2bbdccd, 32'h418d0fc2, 32'h417686db, 32'h42b195c9};
test_output[3282] = '{32'h42b195c9};
test_index[3282] = '{7};
test_input[26264:26271] = '{32'hc1c0e816, 32'hc21c96b0, 32'h4246e696, 32'h42b4317d, 32'hc2bc4d83, 32'hc2380664, 32'h4242db2c, 32'h4213df7d};
test_output[3283] = '{32'h42b4317d};
test_index[3283] = '{3};
test_input[26272:26279] = '{32'h3e773cfe, 32'hbf92fc1d, 32'hc1294273, 32'hc0f74205, 32'h42bc69b4, 32'h41b4e7c3, 32'hc2bd837a, 32'hc21244a3};
test_output[3284] = '{32'h42bc69b4};
test_index[3284] = '{4};
test_input[26280:26287] = '{32'h416a3bcd, 32'hc2bfaa97, 32'h41f108d7, 32'h42aea815, 32'hc1e22600, 32'hc2a42864, 32'h425ee95e, 32'hc2c5e1b4};
test_output[3285] = '{32'h42aea815};
test_index[3285] = '{3};
test_input[26288:26295] = '{32'hc2b64a8a, 32'h429a3a66, 32'h4285abc8, 32'h428c3c55, 32'h423ab7b4, 32'hc2b9e1d4, 32'h428e537d, 32'hc1c5371b};
test_output[3286] = '{32'h429a3a66};
test_index[3286] = '{1};
test_input[26296:26303] = '{32'hc16596d5, 32'hc2654ed0, 32'h4264d142, 32'h42784c30, 32'hc1db2c0f, 32'hc14b0b5f, 32'hc258ebc8, 32'hc24aa38f};
test_output[3287] = '{32'h42784c30};
test_index[3287] = '{3};
test_input[26304:26311] = '{32'hc1440c65, 32'h42b3fedc, 32'h42aafada, 32'hc19ca110, 32'h4019293f, 32'h42890b26, 32'hc1b661d5, 32'hc28bc085};
test_output[3288] = '{32'h42b3fedc};
test_index[3288] = '{1};
test_input[26312:26319] = '{32'hc2c08965, 32'hc2c1419c, 32'h42820b85, 32'hc29c8cba, 32'hc2a697c3, 32'hc294dfce, 32'hc280a682, 32'hc27f556c};
test_output[3289] = '{32'h42820b85};
test_index[3289] = '{2};
test_input[26320:26327] = '{32'hc2aa60f0, 32'h3f88999a, 32'hc1e7f153, 32'hc298106b, 32'h4138edff, 32'hbf1c0613, 32'hc2bc20fc, 32'h42985517};
test_output[3290] = '{32'h42985517};
test_index[3290] = '{7};
test_input[26328:26335] = '{32'hc179adfd, 32'hc1747d3b, 32'hc28798f7, 32'h41817286, 32'h41a4f81d, 32'h428a7179, 32'h423b3428, 32'h420a2167};
test_output[3291] = '{32'h428a7179};
test_index[3291] = '{5};
test_input[26336:26343] = '{32'hc2b806ed, 32'h429b605c, 32'hc29959b6, 32'hc1b9a21a, 32'hc2b009f6, 32'h402e9630, 32'hc2363b1f, 32'h413e9683};
test_output[3292] = '{32'h429b605c};
test_index[3292] = '{1};
test_input[26344:26351] = '{32'hc2887018, 32'h41de7448, 32'h412d1749, 32'h42c617e8, 32'hc28ad162, 32'hc2480afb, 32'hc2953bc6, 32'h424f02a8};
test_output[3293] = '{32'h42c617e8};
test_index[3293] = '{3};
test_input[26352:26359] = '{32'h42883afa, 32'hc2361360, 32'hc2502209, 32'hc1a1b80c, 32'h411f733e, 32'h42932f46, 32'hc2620a89, 32'h401bf0b5};
test_output[3294] = '{32'h42932f46};
test_index[3294] = '{5};
test_input[26360:26367] = '{32'hc23e2514, 32'hc1c57a9d, 32'h42b96f04, 32'h422b3ca6, 32'h42baa10d, 32'hc1eb4100, 32'h41d4079a, 32'hc136d5f8};
test_output[3295] = '{32'h42baa10d};
test_index[3295] = '{4};
test_input[26368:26375] = '{32'h4203b802, 32'hc2810a4a, 32'hc26c1c29, 32'h426b79f0, 32'h42ba626e, 32'hc2963d70, 32'hc260cd3a, 32'hbebddfca};
test_output[3296] = '{32'h42ba626e};
test_index[3296] = '{4};
test_input[26376:26383] = '{32'h42a7f440, 32'h424bf218, 32'hc2aa4fc0, 32'h42280a9c, 32'hc2a6899f, 32'h4289c26e, 32'hc19ed766, 32'h42945834};
test_output[3297] = '{32'h42a7f440};
test_index[3297] = '{0};
test_input[26384:26391] = '{32'h41bb027a, 32'h42b2d164, 32'hc1fef1ab, 32'hc2b14f59, 32'hc2136a2e, 32'h42a4821e, 32'hc0987b8d, 32'h422a7792};
test_output[3298] = '{32'h42b2d164};
test_index[3298] = '{1};
test_input[26392:26399] = '{32'h426413e0, 32'h42aa25cf, 32'h42340cde, 32'h4120d95a, 32'h42b3c54b, 32'hc2c2bfd8, 32'hc29b4a17, 32'hc2529e03};
test_output[3299] = '{32'h42b3c54b};
test_index[3299] = '{4};
test_input[26400:26407] = '{32'hc15887a9, 32'hc1a279e5, 32'hc2c06865, 32'hc1f4a6b4, 32'hc1fa77b6, 32'hc248419f, 32'hc1a78d28, 32'hc1a67cb5};
test_output[3300] = '{32'hc15887a9};
test_index[3300] = '{0};
test_input[26408:26415] = '{32'hc05008d8, 32'hc22228a5, 32'h42c2ea34, 32'h42aeb1ef, 32'hc0bb6f97, 32'hc135fd6f, 32'hc2a0e71d, 32'h42bfc2ae};
test_output[3301] = '{32'h42c2ea34};
test_index[3301] = '{2};
test_input[26416:26423] = '{32'hbfc6b7f6, 32'h425c39ea, 32'hc21b3c99, 32'hc2a7da92, 32'hc28fc652, 32'h41823b9e, 32'h4217f465, 32'h42ba6fd9};
test_output[3302] = '{32'h42ba6fd9};
test_index[3302] = '{7};
test_input[26424:26431] = '{32'h42351480, 32'h41c48219, 32'h42868e4f, 32'h42706cba, 32'h42c05523, 32'hc285640b, 32'h41f86f78, 32'hc25e7a5f};
test_output[3303] = '{32'h42c05523};
test_index[3303] = '{4};
test_input[26432:26439] = '{32'hc2c574f9, 32'h422f261c, 32'hc148af2a, 32'hc2aac008, 32'h4204b8d2, 32'h420c4229, 32'h3fd9d48c, 32'h429ec87f};
test_output[3304] = '{32'h429ec87f};
test_index[3304] = '{7};
test_input[26440:26447] = '{32'hc283d42f, 32'hc2b49b82, 32'hc237b59c, 32'h41ef66de, 32'h42990ae5, 32'h42196d61, 32'h429b2237, 32'h41048d3d};
test_output[3305] = '{32'h429b2237};
test_index[3305] = '{6};
test_input[26448:26455] = '{32'h413aba2c, 32'h4291b8ef, 32'hc29c19e3, 32'h410cb1ae, 32'hc2907e7e, 32'hc2c725a0, 32'hc2a5aae2, 32'h40ac4be2};
test_output[3306] = '{32'h4291b8ef};
test_index[3306] = '{1};
test_input[26456:26463] = '{32'h42c690f6, 32'hc2a0120d, 32'h4236f298, 32'h42b62fe8, 32'h41cb7ea8, 32'hc2065a52, 32'h428145da, 32'hc20208a4};
test_output[3307] = '{32'h42c690f6};
test_index[3307] = '{0};
test_input[26464:26471] = '{32'h41d1dd07, 32'hc2a35823, 32'hc292628d, 32'h42943b23, 32'h42a02312, 32'h42a8264a, 32'hc0614595, 32'h42bbcb25};
test_output[3308] = '{32'h42bbcb25};
test_index[3308] = '{7};
test_input[26472:26479] = '{32'h425a7c43, 32'h420178ba, 32'h42a3e0f1, 32'h42a5e72d, 32'hc1c29416, 32'h42b46cd0, 32'hc2958665, 32'h422024e6};
test_output[3309] = '{32'h42b46cd0};
test_index[3309] = '{5};
test_input[26480:26487] = '{32'h4222faea, 32'hc2a83426, 32'hc2b41004, 32'hc25c3c65, 32'h40f6e597, 32'h40dcdaa6, 32'h42b7536b, 32'hc2850ea6};
test_output[3310] = '{32'h42b7536b};
test_index[3310] = '{6};
test_input[26488:26495] = '{32'h41f61ad7, 32'hc25ffd09, 32'h41b65b8c, 32'h42be5625, 32'hc28bb3b4, 32'hc2af704f, 32'h41a34a1a, 32'h424ae03d};
test_output[3311] = '{32'h42be5625};
test_index[3311] = '{3};
test_input[26496:26503] = '{32'hc231dd69, 32'hc23b1c50, 32'hc2c6af16, 32'hc2b9bb15, 32'hc2651e85, 32'hc0cab34c, 32'hc2a97ae8, 32'h420b551c};
test_output[3312] = '{32'h420b551c};
test_index[3312] = '{7};
test_input[26504:26511] = '{32'h42c72eda, 32'hc148f023, 32'hc174337c, 32'h4285c1bb, 32'hc2b40313, 32'h428a75f2, 32'h428474b8, 32'h40d1db07};
test_output[3313] = '{32'h42c72eda};
test_index[3313] = '{0};
test_input[26512:26519] = '{32'hc2a116f7, 32'hc2b0b473, 32'h424790d2, 32'h41743c1a, 32'hc2bc7054, 32'hc267044b, 32'h429d1cdc, 32'h42ba9418};
test_output[3314] = '{32'h42ba9418};
test_index[3314] = '{7};
test_input[26520:26527] = '{32'h420c9c3c, 32'hc2af5c81, 32'hc2166e51, 32'hc29a1cae, 32'hc296f4be, 32'h40c53f06, 32'hc2aa1c1d, 32'hc26a7cab};
test_output[3315] = '{32'h420c9c3c};
test_index[3315] = '{0};
test_input[26528:26535] = '{32'h42bd5d5d, 32'h42a7dda6, 32'hc20297f4, 32'hbf3ffd39, 32'hc29659bf, 32'h4214d31a, 32'hc05881e1, 32'hc1a72a42};
test_output[3316] = '{32'h42bd5d5d};
test_index[3316] = '{0};
test_input[26536:26543] = '{32'hc2c46fde, 32'hc0c13fba, 32'hc20d2e08, 32'h422df39b, 32'h427bb746, 32'h42a2f5a9, 32'h41dcc4cd, 32'hc11b36d1};
test_output[3317] = '{32'h42a2f5a9};
test_index[3317] = '{5};
test_input[26544:26551] = '{32'hc29aa0e0, 32'hc28b3ac5, 32'hc2be240f, 32'hc1cd68ed, 32'hc233a286, 32'h42ae5c4a, 32'hc290fa1a, 32'hc26619b7};
test_output[3318] = '{32'h42ae5c4a};
test_index[3318] = '{5};
test_input[26552:26559] = '{32'hc2bd930a, 32'hc2ade597, 32'hc218e91d, 32'hc239c4a2, 32'h42bae1bb, 32'h42c6d99a, 32'hc28eff98, 32'h42a719e5};
test_output[3319] = '{32'h42c6d99a};
test_index[3319] = '{5};
test_input[26560:26567] = '{32'h42c7af89, 32'hc2959a32, 32'hc2a69f9a, 32'h42335982, 32'hc2876a69, 32'h4237ac52, 32'hc189c541, 32'h41a06061};
test_output[3320] = '{32'h42c7af89};
test_index[3320] = '{0};
test_input[26568:26575] = '{32'h411e5e94, 32'h4271c26a, 32'hc25785bf, 32'h41aa7838, 32'hc268b0ed, 32'hc2b073de, 32'hc2af8d70, 32'hc18836a8};
test_output[3321] = '{32'h4271c26a};
test_index[3321] = '{1};
test_input[26576:26583] = '{32'h419ff640, 32'h42a1bceb, 32'hc08a4fcc, 32'hc29a1667, 32'h42b32ff9, 32'h4288d828, 32'h40546e93, 32'hc1d710f6};
test_output[3322] = '{32'h42b32ff9};
test_index[3322] = '{4};
test_input[26584:26591] = '{32'h41b03a0d, 32'hc1adfac1, 32'h42318c07, 32'h42b6866b, 32'h424d972a, 32'h4273ab66, 32'hc00d3248, 32'h4249ac96};
test_output[3323] = '{32'h42b6866b};
test_index[3323] = '{3};
test_input[26592:26599] = '{32'h428f5fe8, 32'hc16e9241, 32'hc2800b76, 32'hc1b610eb, 32'hc05a1235, 32'h41c4e9db, 32'h42ad10ab, 32'h422f19b2};
test_output[3324] = '{32'h42ad10ab};
test_index[3324] = '{6};
test_input[26600:26607] = '{32'h420bc74b, 32'h420f57f8, 32'h420d7750, 32'hc2bad8cc, 32'h42731b5f, 32'hc0a36ed3, 32'hc1cf0674, 32'hc249b31b};
test_output[3325] = '{32'h42731b5f};
test_index[3325] = '{4};
test_input[26608:26615] = '{32'h42517db0, 32'hc26dbd6a, 32'hc2b39dca, 32'h4263aea9, 32'hc219c87e, 32'h42c44047, 32'h4225f85f, 32'hc2af7417};
test_output[3326] = '{32'h42c44047};
test_index[3326] = '{5};
test_input[26616:26623] = '{32'hc2c30c86, 32'hc23b4da3, 32'hc1928084, 32'hc2178751, 32'hc22a016a, 32'hc2c083ce, 32'h4226793c, 32'h4242f496};
test_output[3327] = '{32'h4242f496};
test_index[3327] = '{7};
test_input[26624:26631] = '{32'h42ac9f63, 32'hc2451b8a, 32'h429164cd, 32'h421379b9, 32'h4284cb69, 32'hc2232595, 32'hc25647b3, 32'h428b4507};
test_output[3328] = '{32'h42ac9f63};
test_index[3328] = '{0};
test_input[26632:26639] = '{32'hc2bd1375, 32'h42267a4b, 32'hc1cc91c9, 32'hc1bdaa7b, 32'h426afa37, 32'hc2b2c9aa, 32'h428f94b2, 32'h4273f596};
test_output[3329] = '{32'h428f94b2};
test_index[3329] = '{6};
test_input[26640:26647] = '{32'h4157d51c, 32'hc29488bb, 32'hc1f2d363, 32'h4200a366, 32'h419b0091, 32'h41ac4340, 32'h422b042e, 32'hc29cae6e};
test_output[3330] = '{32'h422b042e};
test_index[3330] = '{6};
test_input[26648:26655] = '{32'hc24dc931, 32'hc14c4fe2, 32'hc2910ff3, 32'h428a1c0a, 32'h42592095, 32'hc2559576, 32'hc20ee2a4, 32'h42127672};
test_output[3331] = '{32'h428a1c0a};
test_index[3331] = '{3};
test_input[26656:26663] = '{32'hc2828057, 32'hc253c4fe, 32'h405ce688, 32'hc22de69b, 32'h42b2dace, 32'hc23530bf, 32'h424c1545, 32'hc27e6bb1};
test_output[3332] = '{32'h42b2dace};
test_index[3332] = '{4};
test_input[26664:26671] = '{32'hc2c0f945, 32'hc29e7454, 32'hc2bc35eb, 32'hc294c734, 32'hc29a1aa8, 32'hc0ee0fa2, 32'hc2860b93, 32'h42a7d2ea};
test_output[3333] = '{32'h42a7d2ea};
test_index[3333] = '{7};
test_input[26672:26679] = '{32'h42636806, 32'h42249c6f, 32'hc1838633, 32'h42c30ab0, 32'h418bf08c, 32'hc23df5b6, 32'h42b67ab9, 32'h425b2108};
test_output[3334] = '{32'h42c30ab0};
test_index[3334] = '{3};
test_input[26680:26687] = '{32'h41ce5fe8, 32'h4271ed96, 32'h41d4003b, 32'hc0668b5a, 32'h42622878, 32'hc203fbd3, 32'hc20f9548, 32'h41c76cd1};
test_output[3335] = '{32'h4271ed96};
test_index[3335] = '{1};
test_input[26688:26695] = '{32'hc18d4569, 32'h41bb0ace, 32'hc1884b71, 32'h42561ffa, 32'hc279fbf1, 32'h40fb3881, 32'hc2ad335d, 32'hc1e38eae};
test_output[3336] = '{32'h42561ffa};
test_index[3336] = '{3};
test_input[26696:26703] = '{32'hc250af9d, 32'hc2045d9c, 32'hc1b6ed8f, 32'h423f3892, 32'h3eb5893f, 32'h420a9f34, 32'h40108a3f, 32'hc1a89c6d};
test_output[3337] = '{32'h423f3892};
test_index[3337] = '{3};
test_input[26704:26711] = '{32'h40ff7e83, 32'h42656ff4, 32'hc1a59cd1, 32'hc29b2d87, 32'h416a8a7e, 32'h4025b584, 32'hc1ffe118, 32'h40251868};
test_output[3338] = '{32'h42656ff4};
test_index[3338] = '{1};
test_input[26712:26719] = '{32'h41d28576, 32'hc0f78256, 32'hc28f90af, 32'hc17891b3, 32'h40896276, 32'h4114ce61, 32'hc1a84409, 32'h42960692};
test_output[3339] = '{32'h42960692};
test_index[3339] = '{7};
test_input[26720:26727] = '{32'h428155d2, 32'hc28647de, 32'h4268631f, 32'hc212f37b, 32'hc00be21a, 32'h419a8e0e, 32'hc19c1b13, 32'h4080282c};
test_output[3340] = '{32'h428155d2};
test_index[3340] = '{0};
test_input[26728:26735] = '{32'h42c1ca55, 32'hc1d74ebe, 32'hc20daf30, 32'h42596c3d, 32'h41de3e01, 32'hc24ac30c, 32'h427b945e, 32'h41fd3edc};
test_output[3341] = '{32'h42c1ca55};
test_index[3341] = '{0};
test_input[26736:26743] = '{32'hc2939af5, 32'hc2973037, 32'hc2765ee5, 32'hc22dc7d4, 32'hc26d1ec4, 32'h42b7b418, 32'h421f3092, 32'h428916eb};
test_output[3342] = '{32'h42b7b418};
test_index[3342] = '{5};
test_input[26744:26751] = '{32'h421bbc66, 32'h41e23311, 32'hc2c4f36d, 32'hc261233e, 32'h41808110, 32'h424db374, 32'h3fb95748, 32'h424e41df};
test_output[3343] = '{32'h424e41df};
test_index[3343] = '{7};
test_input[26752:26759] = '{32'hc2b504d0, 32'h4195c45b, 32'hc29212d5, 32'hc29e0d9e, 32'hc240a87d, 32'h4243c25e, 32'hc2b499b2, 32'hc1db2279};
test_output[3344] = '{32'h4243c25e};
test_index[3344] = '{5};
test_input[26760:26767] = '{32'h424b798c, 32'hc2277e8c, 32'h4293c017, 32'h42492986, 32'h42a7b55d, 32'hc244d90f, 32'h42942383, 32'h419f8dec};
test_output[3345] = '{32'h42a7b55d};
test_index[3345] = '{4};
test_input[26768:26775] = '{32'h4290b8ff, 32'h423da2e3, 32'h427ff503, 32'h42435863, 32'hc1b4a60e, 32'h42136609, 32'hc29126cc, 32'hc28e14c0};
test_output[3346] = '{32'h4290b8ff};
test_index[3346] = '{0};
test_input[26776:26783] = '{32'hc250bb8f, 32'h41bd6365, 32'h41696bf9, 32'hc18d9352, 32'h42231881, 32'h42266d22, 32'h422d0ae1, 32'hc2c3b930};
test_output[3347] = '{32'h422d0ae1};
test_index[3347] = '{6};
test_input[26784:26791] = '{32'hc28af12d, 32'hc265988f, 32'h3fe09e91, 32'hc26476f7, 32'hc2a361f6, 32'h4158eb81, 32'hc2b668a6, 32'hc25b6e96};
test_output[3348] = '{32'h4158eb81};
test_index[3348] = '{5};
test_input[26792:26799] = '{32'h428d7df8, 32'hc214fd31, 32'h41dde956, 32'hc292b692, 32'hc2b25d05, 32'h428ac0c0, 32'hc2a5c155, 32'hc2b6dc82};
test_output[3349] = '{32'h428d7df8};
test_index[3349] = '{0};
test_input[26800:26807] = '{32'h41805436, 32'hc0662f56, 32'hc1e88d09, 32'h429a920e, 32'hc2886ff8, 32'h4094b5b1, 32'h428d16e9, 32'hc2b1f85c};
test_output[3350] = '{32'h429a920e};
test_index[3350] = '{3};
test_input[26808:26815] = '{32'h41984161, 32'h4123af77, 32'h42ac910e, 32'h421345bf, 32'hc253bc02, 32'h42c005e2, 32'h4242b383, 32'hc1936049};
test_output[3351] = '{32'h42c005e2};
test_index[3351] = '{5};
test_input[26816:26823] = '{32'hc28f0859, 32'hc24acc06, 32'hbed33107, 32'h429663ea, 32'h42816933, 32'hc15e057b, 32'hc22707d7, 32'h427c144c};
test_output[3352] = '{32'h429663ea};
test_index[3352] = '{3};
test_input[26824:26831] = '{32'hc2596365, 32'h42969e99, 32'h41eac51a, 32'h4248eaf8, 32'hc24ac3c3, 32'hc28bef41, 32'hc167be31, 32'h42040911};
test_output[3353] = '{32'h42969e99};
test_index[3353] = '{1};
test_input[26832:26839] = '{32'h4271c133, 32'h423d0ba8, 32'hc23aea6e, 32'h42a6c497, 32'h42a26f7b, 32'hc245e08a, 32'h4155ead6, 32'hc2b15ab5};
test_output[3354] = '{32'h42a6c497};
test_index[3354] = '{3};
test_input[26840:26847] = '{32'h423517a5, 32'h425b22a3, 32'h414650b1, 32'h429b605f, 32'h42ab1af7, 32'hc236830b, 32'hc29dca31, 32'h42af4929};
test_output[3355] = '{32'h42af4929};
test_index[3355] = '{7};
test_input[26848:26855] = '{32'h41c9f774, 32'h42c3509a, 32'hc28a19f3, 32'hc22e8eaf, 32'hc145334d, 32'h42a8076f, 32'hc17b16ff, 32'h4266e0a1};
test_output[3356] = '{32'h42c3509a};
test_index[3356] = '{1};
test_input[26856:26863] = '{32'h41e54263, 32'h41a757e4, 32'h42b525aa, 32'h42c3b909, 32'h42b0de79, 32'h42b89649, 32'h42ab763f, 32'h41982d48};
test_output[3357] = '{32'h42c3b909};
test_index[3357] = '{3};
test_input[26864:26871] = '{32'h425b92ca, 32'hc25be72b, 32'hc280583e, 32'hc2a8a305, 32'hc246b896, 32'hc253c264, 32'hbf965906, 32'h42b6fed7};
test_output[3358] = '{32'h42b6fed7};
test_index[3358] = '{7};
test_input[26872:26879] = '{32'h42ad0891, 32'h4293c708, 32'hc291ed3b, 32'hc28a52a0, 32'h42877b9a, 32'h425f406f, 32'h4208b7d8, 32'hc1c8b78e};
test_output[3359] = '{32'h42ad0891};
test_index[3359] = '{0};
test_input[26880:26887] = '{32'h428e550e, 32'h4196785e, 32'h41e727cf, 32'h4239793f, 32'hc258691c, 32'hc2234e01, 32'h4253a178, 32'hc25b4e00};
test_output[3360] = '{32'h428e550e};
test_index[3360] = '{0};
test_input[26888:26895] = '{32'hc2180fb0, 32'h4280b23c, 32'hc2a01acb, 32'hc2303a26, 32'h4237686a, 32'hc235cd7b, 32'h426c6fce, 32'h4170b1c6};
test_output[3361] = '{32'h4280b23c};
test_index[3361] = '{1};
test_input[26896:26903] = '{32'h42091b5d, 32'h42937ad9, 32'h4123c018, 32'hc129e041, 32'h415b1216, 32'hc2a4f6ca, 32'h42113716, 32'h3ca2764d};
test_output[3362] = '{32'h42937ad9};
test_index[3362] = '{1};
test_input[26904:26911] = '{32'hc1ed787a, 32'hbff66cb9, 32'h429960b7, 32'h4209d97b, 32'h42768a8c, 32'h41a347c6, 32'h41911aad, 32'h40e2bd27};
test_output[3363] = '{32'h429960b7};
test_index[3363] = '{2};
test_input[26912:26919] = '{32'hc24f59e3, 32'h424824b4, 32'hc13d6d3c, 32'hc1834040, 32'h41dcc4b4, 32'hc26a429b, 32'hc229676f, 32'hbfaee636};
test_output[3364] = '{32'h424824b4};
test_index[3364] = '{1};
test_input[26920:26927] = '{32'hc2af7b2e, 32'h4258d17b, 32'h42af113f, 32'hc156b820, 32'h424aaf92, 32'hc2a095cb, 32'h41bc74d5, 32'h424b3940};
test_output[3365] = '{32'h42af113f};
test_index[3365] = '{2};
test_input[26928:26935] = '{32'h41a8d0ff, 32'h4296514d, 32'hc1c472b6, 32'h42860710, 32'h42a0456b, 32'h40f4ccf6, 32'h413167b1, 32'hc22cbd3b};
test_output[3366] = '{32'h42a0456b};
test_index[3366] = '{4};
test_input[26936:26943] = '{32'hc21bbb7a, 32'h41367a67, 32'h4104290f, 32'h42b096d6, 32'h42aeb7a1, 32'hc29d5260, 32'hc298a344, 32'hc1dffa3b};
test_output[3367] = '{32'h42b096d6};
test_index[3367] = '{3};
test_input[26944:26951] = '{32'hc224a767, 32'h42c0cf6c, 32'hc28c29b5, 32'h417bf123, 32'h428352e2, 32'hc277f7d7, 32'hc2b9654e, 32'hc2c6e7b5};
test_output[3368] = '{32'h42c0cf6c};
test_index[3368] = '{1};
test_input[26952:26959] = '{32'h42981213, 32'h42a20d25, 32'hc29cd73e, 32'hc2b08b7c, 32'hc1bbe015, 32'hc2b7f4ed, 32'hc264e70e, 32'hc26e97ce};
test_output[3369] = '{32'h42a20d25};
test_index[3369] = '{1};
test_input[26960:26967] = '{32'h42c32d1d, 32'h42b09d94, 32'h4299f399, 32'hc15b029a, 32'hc280ff2f, 32'h4215f937, 32'h420e997f, 32'hc05b852b};
test_output[3370] = '{32'h42c32d1d};
test_index[3370] = '{0};
test_input[26968:26975] = '{32'hc21457df, 32'hbfb635f5, 32'hc25f2f60, 32'h42037ff5, 32'hbeaef511, 32'hc22158da, 32'hc0d53e3f, 32'h40f5618a};
test_output[3371] = '{32'h42037ff5};
test_index[3371] = '{3};
test_input[26976:26983] = '{32'hc18c7b0e, 32'hc23b0c8f, 32'h426880da, 32'hc27059a1, 32'hc2a8c2cc, 32'h425f4490, 32'hc2b1959a, 32'h424e88ae};
test_output[3372] = '{32'h426880da};
test_index[3372] = '{2};
test_input[26984:26991] = '{32'hc1c17855, 32'hc2877129, 32'hc297bf3b, 32'h42ab6724, 32'hc2c0062b, 32'h429794c7, 32'h42c1ae14, 32'h428b8112};
test_output[3373] = '{32'h42c1ae14};
test_index[3373] = '{6};
test_input[26992:26999] = '{32'h420f231e, 32'hc28c3478, 32'hc2218aeb, 32'h4284f224, 32'hc16cca67, 32'hc2896d56, 32'h429a4cae, 32'h422a676a};
test_output[3374] = '{32'h429a4cae};
test_index[3374] = '{6};
test_input[27000:27007] = '{32'h42954b81, 32'hc28bbc85, 32'hc2234e1f, 32'h4215e226, 32'hc29e62c9, 32'h41d20341, 32'hc240c960, 32'h42c3fae9};
test_output[3375] = '{32'h42c3fae9};
test_index[3375] = '{7};
test_input[27008:27015] = '{32'h41051c80, 32'hc24f53b0, 32'h4235534d, 32'h422f6d32, 32'h42b34b79, 32'hc16b13e1, 32'hc235639d, 32'hc18efbdb};
test_output[3376] = '{32'h42b34b79};
test_index[3376] = '{4};
test_input[27016:27023] = '{32'hc241bc92, 32'hc1cc46ed, 32'h42b75684, 32'hc28663e3, 32'hc0593955, 32'hc28a939b, 32'hc277f60f, 32'hc23ccce5};
test_output[3377] = '{32'h42b75684};
test_index[3377] = '{2};
test_input[27024:27031] = '{32'hc2020e66, 32'hc1828f23, 32'hc28a755e, 32'h419bfc6c, 32'h420586fc, 32'hc181bfdd, 32'hc2bb754e, 32'hc1b69830};
test_output[3378] = '{32'h420586fc};
test_index[3378] = '{4};
test_input[27032:27039] = '{32'hc15c25d2, 32'hc2537aca, 32'hc22ed4ba, 32'hc1f5eb3c, 32'h4152ebb4, 32'hc29394bd, 32'hc2c3b357, 32'hc2a1af6a};
test_output[3379] = '{32'h4152ebb4};
test_index[3379] = '{4};
test_input[27040:27047] = '{32'h3f5fef08, 32'h4256b1a3, 32'h425ddb44, 32'hc24fdd94, 32'hc29234d9, 32'hc29b0a76, 32'h42006371, 32'h4269277c};
test_output[3380] = '{32'h4269277c};
test_index[3380] = '{7};
test_input[27048:27055] = '{32'hc2a36b4c, 32'h42c0a948, 32'h42313e08, 32'h3f973099, 32'hbec7b75b, 32'h421dd89b, 32'hc1cf967e, 32'hc2298f57};
test_output[3381] = '{32'h42c0a948};
test_index[3381] = '{1};
test_input[27056:27063] = '{32'hc185a23f, 32'h42206fdc, 32'h40ab1220, 32'h4235617d, 32'hc23f0550, 32'h42876d38, 32'hc2957af4, 32'hc20f43b1};
test_output[3382] = '{32'h42876d38};
test_index[3382] = '{5};
test_input[27064:27071] = '{32'h429e3559, 32'h4206126c, 32'hc02e94ea, 32'hc2c3ed81, 32'h427d8571, 32'hc28e3c6e, 32'h425262bb, 32'hc2a35970};
test_output[3383] = '{32'h429e3559};
test_index[3383] = '{0};
test_input[27072:27079] = '{32'h42b1104f, 32'hc09b33ee, 32'hc2b2f112, 32'hc282b191, 32'h4268797b, 32'hc29c2a33, 32'hc249f2f3, 32'hc2bbccdc};
test_output[3384] = '{32'h42b1104f};
test_index[3384] = '{0};
test_input[27080:27087] = '{32'h41adc3e2, 32'hc241f2ef, 32'h425b4c03, 32'h42b4a4de, 32'hc1c8b5fe, 32'hc2853e6b, 32'h41e58997, 32'hc28d1e73};
test_output[3385] = '{32'h42b4a4de};
test_index[3385] = '{3};
test_input[27088:27095] = '{32'hc206fa35, 32'h42b4605d, 32'h40910f5d, 32'h423f6b4b, 32'h42a87695, 32'h41b1a039, 32'hc2837708, 32'h427e0eaf};
test_output[3386] = '{32'h42b4605d};
test_index[3386] = '{1};
test_input[27096:27103] = '{32'h41a4dbce, 32'hc2b10dd1, 32'hc2b0fc4b, 32'h3f0c7899, 32'h423ae14c, 32'hc2afd93c, 32'hc28a3294, 32'hc2936166};
test_output[3387] = '{32'h423ae14c};
test_index[3387] = '{4};
test_input[27104:27111] = '{32'hc23f0c5e, 32'h42c17c8a, 32'h41b907d3, 32'h4139cd07, 32'hc2a4c78d, 32'hbeff09bf, 32'h415dc527, 32'h42c325e5};
test_output[3388] = '{32'h42c325e5};
test_index[3388] = '{7};
test_input[27112:27119] = '{32'hc0db643e, 32'h42a89af1, 32'hc29a74a0, 32'hc1cd6eb7, 32'hc276f6ac, 32'hc117f7bb, 32'hc2a53d64, 32'h425eaf0a};
test_output[3389] = '{32'h42a89af1};
test_index[3389] = '{1};
test_input[27120:27127] = '{32'hc173a8d8, 32'h3d8cc46a, 32'h42c467d6, 32'h428a169b, 32'hc22d3af8, 32'h42c535a6, 32'h42b74e9d, 32'hc282001e};
test_output[3390] = '{32'h42c535a6};
test_index[3390] = '{5};
test_input[27128:27135] = '{32'h428e65e9, 32'h42b2e540, 32'hc2ac9cc7, 32'h42a34e89, 32'h429d8963, 32'hc234752a, 32'hc15d1534, 32'hc2290206};
test_output[3391] = '{32'h42b2e540};
test_index[3391] = '{1};
test_input[27136:27143] = '{32'h42b73946, 32'hc2c5f3b5, 32'hc1dfa66f, 32'h42bed389, 32'hc2c230d2, 32'hc20506a6, 32'hc280e5a9, 32'hc1d96e8d};
test_output[3392] = '{32'h42bed389};
test_index[3392] = '{3};
test_input[27144:27151] = '{32'hc24e6080, 32'hc25a30cd, 32'hc2688bd7, 32'h42bfbae7, 32'hc23a3dcd, 32'h427dfb0b, 32'hc1ab622b, 32'hc232d737};
test_output[3393] = '{32'h42bfbae7};
test_index[3393] = '{3};
test_input[27152:27159] = '{32'hc2bdb033, 32'h4244386a, 32'hc217ce10, 32'h426998d4, 32'hc2c3cf96, 32'h41fa83e6, 32'hc2a60eea, 32'h40edbdac};
test_output[3394] = '{32'h426998d4};
test_index[3394] = '{3};
test_input[27160:27167] = '{32'hc29c1120, 32'hc211ff8b, 32'hc2a0b191, 32'hc2b75c21, 32'hc2b40e5d, 32'h42134f03, 32'hbf8545c3, 32'hc2aa1259};
test_output[3395] = '{32'h42134f03};
test_index[3395] = '{5};
test_input[27168:27175] = '{32'h42836497, 32'h42b7e7a2, 32'h415a37da, 32'hc265cfb4, 32'h420cd4b3, 32'hc2717a6f, 32'h42886efc, 32'hc29bdecc};
test_output[3396] = '{32'h42b7e7a2};
test_index[3396] = '{1};
test_input[27176:27183] = '{32'hc2a9783b, 32'hc107905d, 32'h42297aac, 32'hc264d24e, 32'h412536d2, 32'hc21539cb, 32'hc2a46d2a, 32'hc28ff044};
test_output[3397] = '{32'h42297aac};
test_index[3397] = '{2};
test_input[27184:27191] = '{32'hc26e92b0, 32'hc280ce8d, 32'h42aeb00b, 32'hc1917cd1, 32'hc0880be8, 32'hc0a1188f, 32'hc123acd0, 32'h42a56574};
test_output[3398] = '{32'h42aeb00b};
test_index[3398] = '{2};
test_input[27192:27199] = '{32'hc245eed5, 32'h4241aa3d, 32'hc1919d72, 32'hc2796607, 32'hc20f7aec, 32'hc2936051, 32'h421f36ee, 32'h412fe95e};
test_output[3399] = '{32'h4241aa3d};
test_index[3399] = '{1};
test_input[27200:27207] = '{32'hc2c0fcb4, 32'hc1bdd66d, 32'h41d94562, 32'hc28095a9, 32'h4226262f, 32'h3fabebc4, 32'hc2977b64, 32'h41a9ca15};
test_output[3400] = '{32'h4226262f};
test_index[3400] = '{4};
test_input[27208:27215] = '{32'hc2866a28, 32'hc2ab21de, 32'h42a9a802, 32'hc27a0dbe, 32'h4226e177, 32'hc24cc065, 32'hc2af0235, 32'h4163973b};
test_output[3401] = '{32'h42a9a802};
test_index[3401] = '{2};
test_input[27216:27223] = '{32'hc299d3b9, 32'h41d99c33, 32'hc2786fe0, 32'h418d6bb8, 32'hc242bd2a, 32'h42a2dfeb, 32'h42b5ad28, 32'hc1ca7b01};
test_output[3402] = '{32'h42b5ad28};
test_index[3402] = '{6};
test_input[27224:27231] = '{32'hc090f03e, 32'h3f84c252, 32'hc0ff182e, 32'hc1dddb37, 32'h4270dafd, 32'h428130eb, 32'hc28c219f, 32'h42bea8f7};
test_output[3403] = '{32'h42bea8f7};
test_index[3403] = '{7};
test_input[27232:27239] = '{32'hc2722f50, 32'h42bcd0a8, 32'h427bd354, 32'h42b5358a, 32'h4299893f, 32'hc268abcd, 32'h42918eed, 32'hc2ad8758};
test_output[3404] = '{32'h42bcd0a8};
test_index[3404] = '{1};
test_input[27240:27247] = '{32'h42b89963, 32'hc1c4cfeb, 32'h423a4060, 32'hc25945be, 32'h428b3252, 32'h42ba3310, 32'hc2a51d3b, 32'h42c56823};
test_output[3405] = '{32'h42c56823};
test_index[3405] = '{7};
test_input[27248:27255] = '{32'h4221bd00, 32'hc2a65fc2, 32'hc29bb519, 32'h42aeb8c0, 32'h410a7077, 32'hc1f2cdfc, 32'hc1d174e0, 32'hc247309c};
test_output[3406] = '{32'h42aeb8c0};
test_index[3406] = '{3};
test_input[27256:27263] = '{32'hc19e1de2, 32'h41f3740c, 32'h42104508, 32'hc25e4329, 32'hc0b39639, 32'h4296c1f3, 32'hc11ad61c, 32'h41e1bfea};
test_output[3407] = '{32'h4296c1f3};
test_index[3407] = '{5};
test_input[27264:27271] = '{32'h4267c7e1, 32'h423c463e, 32'hc2a2d217, 32'hc2b62ec4, 32'hc28f09fc, 32'hc217479c, 32'h4156614e, 32'h41efa913};
test_output[3408] = '{32'h4267c7e1};
test_index[3408] = '{0};
test_input[27272:27279] = '{32'h41923497, 32'hc29728d2, 32'hc2b70a66, 32'hc2aa3771, 32'h42aae044, 32'hc1c6f53a, 32'hc1caee64, 32'h42300a0b};
test_output[3409] = '{32'h42aae044};
test_index[3409] = '{4};
test_input[27280:27287] = '{32'hc28b7da8, 32'hc27f4b06, 32'hc26710a2, 32'h41bba262, 32'h42ab6261, 32'hbe438c96, 32'h420c2eeb, 32'hc1e66680};
test_output[3410] = '{32'h42ab6261};
test_index[3410] = '{4};
test_input[27288:27295] = '{32'hc20f3fdc, 32'h4273d5c6, 32'h40fb44f5, 32'h41e21f26, 32'hc2ac9eee, 32'hc19e93bb, 32'hc1a7f1f3, 32'h42222a90};
test_output[3411] = '{32'h4273d5c6};
test_index[3411] = '{1};
test_input[27296:27303] = '{32'h4299667a, 32'hc2828273, 32'h42a817c6, 32'hc1acbefd, 32'hc09c150b, 32'h42c06539, 32'h4215178f, 32'h4145f9f6};
test_output[3412] = '{32'h42c06539};
test_index[3412] = '{5};
test_input[27304:27311] = '{32'hc287b66f, 32'hc2b4b5bd, 32'hc28e30f3, 32'h3ef870c3, 32'h42aec7a0, 32'hc25a82fe, 32'h41a7440d, 32'h41851c56};
test_output[3413] = '{32'h42aec7a0};
test_index[3413] = '{4};
test_input[27312:27319] = '{32'h42c39c6a, 32'h41a267bd, 32'hc289cc14, 32'h41f920aa, 32'hc0d8656b, 32'hc19f554e, 32'hc224ba7f, 32'h415a0521};
test_output[3414] = '{32'h42c39c6a};
test_index[3414] = '{0};
test_input[27320:27327] = '{32'hc27ddffe, 32'h40b44463, 32'h42042448, 32'h402d0d9d, 32'hc2aab005, 32'hc13c61ba, 32'h4191aa68, 32'h4245b835};
test_output[3415] = '{32'h4245b835};
test_index[3415] = '{7};
test_input[27328:27335] = '{32'h4110e24d, 32'hc2b0ab57, 32'h42b13322, 32'hc1752402, 32'h41b90642, 32'hc2587bd2, 32'h42825576, 32'h4293b1ef};
test_output[3416] = '{32'h42b13322};
test_index[3416] = '{2};
test_input[27336:27343] = '{32'hc2af5282, 32'hc27d4b03, 32'hc2210ac8, 32'hc28d6b19, 32'hc1ab5a89, 32'h42bf62ce, 32'h42bd00c7, 32'h424245de};
test_output[3417] = '{32'h42bf62ce};
test_index[3417] = '{5};
test_input[27344:27351] = '{32'hc2bab889, 32'h41379070, 32'hc2bdfca6, 32'hc157a178, 32'h429189a5, 32'hc29f17ad, 32'h42846494, 32'h4197e0f3};
test_output[3418] = '{32'h429189a5};
test_index[3418] = '{4};
test_input[27352:27359] = '{32'h4201ee84, 32'hc25cb062, 32'h42ab2e6c, 32'h42249f0b, 32'hc2370d37, 32'h42019f13, 32'hc2c1ede6, 32'hc282b7cf};
test_output[3419] = '{32'h42ab2e6c};
test_index[3419] = '{2};
test_input[27360:27367] = '{32'h4274d0ae, 32'hc2bd82e9, 32'h42a44489, 32'h42c750a2, 32'hc1a90554, 32'h41e3c3ff, 32'hbf135284, 32'hc283e8e8};
test_output[3420] = '{32'h42c750a2};
test_index[3420] = '{3};
test_input[27368:27375] = '{32'h429878c9, 32'h42003fea, 32'h421da352, 32'hc26cac87, 32'h427e2cba, 32'h41ed4f2e, 32'h4031953d, 32'h411a87b0};
test_output[3421] = '{32'h429878c9};
test_index[3421] = '{0};
test_input[27376:27383] = '{32'h428d2409, 32'h41f0235c, 32'hc2b7748b, 32'h4174c44b, 32'hc258861d, 32'hc2b241b8, 32'h424aa1cc, 32'h429208de};
test_output[3422] = '{32'h429208de};
test_index[3422] = '{7};
test_input[27384:27391] = '{32'hc2bf8a3f, 32'hc0a51cbe, 32'h428c85ba, 32'h429e87c2, 32'h42a56d29, 32'h42a60dce, 32'hc2a7cb5e, 32'h41ea0e69};
test_output[3423] = '{32'h42a60dce};
test_index[3423] = '{5};
test_input[27392:27399] = '{32'h42886026, 32'hc2498355, 32'h4285518a, 32'hc15f70a7, 32'h422ad431, 32'hc28d904b, 32'h41ec3621, 32'h4271d824};
test_output[3424] = '{32'h42886026};
test_index[3424] = '{0};
test_input[27400:27407] = '{32'h422f301d, 32'hc2b68cfa, 32'hc14e3b11, 32'h412c7fe2, 32'h418000ab, 32'h429ae617, 32'hc2be8f0a, 32'h414c519c};
test_output[3425] = '{32'h429ae617};
test_index[3425] = '{5};
test_input[27408:27415] = '{32'hc1ea78f2, 32'hc2083e0b, 32'hc2a9915c, 32'h4222902a, 32'hc2a00508, 32'hc1baf399, 32'h3f6e063b, 32'hc20ac6be};
test_output[3426] = '{32'h4222902a};
test_index[3426] = '{3};
test_input[27416:27423] = '{32'hc2b016c8, 32'h40c16f36, 32'hc25dd3f0, 32'h42263193, 32'hc2b5e79f, 32'hc2a18f09, 32'hc2c161f5, 32'hc29d6984};
test_output[3427] = '{32'h42263193};
test_index[3427] = '{3};
test_input[27424:27431] = '{32'h42c71b38, 32'h4222075b, 32'h42b668e5, 32'hc216f341, 32'hc290e25f, 32'hc21de58f, 32'h40bc805c, 32'hc20b6e44};
test_output[3428] = '{32'h42c71b38};
test_index[3428] = '{0};
test_input[27432:27439] = '{32'hc19e24b1, 32'h4298cec6, 32'hc0d05749, 32'hc2c3892b, 32'h424b2364, 32'h42a1822e, 32'h420ccd40, 32'h42197671};
test_output[3429] = '{32'h42a1822e};
test_index[3429] = '{5};
test_input[27440:27447] = '{32'hc2ade61c, 32'h42a8c842, 32'h42c5d1ac, 32'hc22c3c19, 32'hc2542a26, 32'h427ae833, 32'hc1415655, 32'h41f9b775};
test_output[3430] = '{32'h42c5d1ac};
test_index[3430] = '{2};
test_input[27448:27455] = '{32'hc249d66d, 32'h42b045e9, 32'hc2a694b7, 32'hc1cbc8cb, 32'hc0c6270d, 32'hc2bcc467, 32'hc29999b5, 32'hc1bceb22};
test_output[3431] = '{32'h42b045e9};
test_index[3431] = '{1};
test_input[27456:27463] = '{32'hc2a47a5e, 32'hc28f42f4, 32'h42465aa1, 32'h427d7634, 32'hc2a33cd5, 32'hc1bebc51, 32'hc2176b79, 32'h422af5ed};
test_output[3432] = '{32'h427d7634};
test_index[3432] = '{3};
test_input[27464:27471] = '{32'h42b5502b, 32'h421a29c0, 32'h42a918ca, 32'h42beac20, 32'hc28ba28e, 32'hc29b54da, 32'h42a92987, 32'hc29f183d};
test_output[3433] = '{32'h42beac20};
test_index[3433] = '{3};
test_input[27472:27479] = '{32'h426d23c8, 32'hc2bbdcbf, 32'hc2c7601e, 32'hc2716bf1, 32'hc27ab092, 32'h42c44d83, 32'h41398459, 32'hc2c22ffd};
test_output[3434] = '{32'h42c44d83};
test_index[3434] = '{5};
test_input[27480:27487] = '{32'hc11e181b, 32'hc2c67532, 32'h42b7c9d5, 32'h410436cb, 32'h411dc23b, 32'hc253e80b, 32'h42adb583, 32'hc0491275};
test_output[3435] = '{32'h42b7c9d5};
test_index[3435] = '{2};
test_input[27488:27495] = '{32'hc265fe5a, 32'h42c479b0, 32'h425b6e5e, 32'h429723d9, 32'hc28c72bd, 32'h42399f9c, 32'hc2873336, 32'h41f1c8a3};
test_output[3436] = '{32'h42c479b0};
test_index[3436] = '{1};
test_input[27496:27503] = '{32'hc2c72edf, 32'hc2b9a8eb, 32'hc20e6729, 32'hc2b99b75, 32'hc250928c, 32'hc2423129, 32'h426e95ff, 32'h42a7535a};
test_output[3437] = '{32'h42a7535a};
test_index[3437] = '{7};
test_input[27504:27511] = '{32'h42989950, 32'hc170a182, 32'hc1de88f3, 32'hc2b96d4c, 32'hc1964cd0, 32'hc288cef3, 32'h41384d18, 32'hc27ee7b7};
test_output[3438] = '{32'h42989950};
test_index[3438] = '{0};
test_input[27512:27519] = '{32'hc2bb0ef1, 32'h429f01f7, 32'hc2aa63dd, 32'hc203642e, 32'h419f85e7, 32'h42887224, 32'h41ccfef9, 32'hc2368ce8};
test_output[3439] = '{32'h429f01f7};
test_index[3439] = '{1};
test_input[27520:27527] = '{32'hc2ab0b2c, 32'h4269e443, 32'hc0f1fea6, 32'hc1933457, 32'h428cf7c1, 32'h425b8506, 32'hc250d4b9, 32'h425b1ac3};
test_output[3440] = '{32'h428cf7c1};
test_index[3440] = '{4};
test_input[27528:27535] = '{32'hc2af4985, 32'h410cdfca, 32'hc2a1ad6d, 32'hc2806e49, 32'h429ab9c0, 32'h42a14e4c, 32'h427fb725, 32'hc0e56d8b};
test_output[3441] = '{32'h42a14e4c};
test_index[3441] = '{5};
test_input[27536:27543] = '{32'hc2722a92, 32'h428edfed, 32'hc26b38b6, 32'h42bddc5c, 32'h425b7734, 32'hc1845f01, 32'h41fd1bb8, 32'h42927dd5};
test_output[3442] = '{32'h42bddc5c};
test_index[3442] = '{3};
test_input[27544:27551] = '{32'h42b3904a, 32'hc25da331, 32'h42262606, 32'hc2924fbb, 32'h41d5d357, 32'h427e9d59, 32'hc2954a5c, 32'hc229efee};
test_output[3443] = '{32'h42b3904a};
test_index[3443] = '{0};
test_input[27552:27559] = '{32'h4186f96a, 32'h42c22456, 32'hc213ce2c, 32'h4284c33d, 32'h4297840e, 32'hc1b8388d, 32'hc242278e, 32'h42672ee0};
test_output[3444] = '{32'h42c22456};
test_index[3444] = '{1};
test_input[27560:27567] = '{32'hc1cce41b, 32'hc27a190d, 32'hc1d973e8, 32'hc21b1aa8, 32'hc1041f33, 32'h424f0c58, 32'h42aa5fa7, 32'hc18c85fd};
test_output[3445] = '{32'h42aa5fa7};
test_index[3445] = '{6};
test_input[27568:27575] = '{32'hc27b2aec, 32'hc23e05d9, 32'hc207f77a, 32'h4180efeb, 32'hc10a6998, 32'hc290b69f, 32'h4220ad9b, 32'hc2447a2b};
test_output[3446] = '{32'h4220ad9b};
test_index[3446] = '{6};
test_input[27576:27583] = '{32'hc2873a3a, 32'hc22bdd76, 32'h427f0872, 32'h42c52006, 32'h42a24221, 32'h4276664b, 32'h3f5eb7ba, 32'h41f90f22};
test_output[3447] = '{32'h42c52006};
test_index[3447] = '{3};
test_input[27584:27591] = '{32'h41ff8760, 32'h42bd1f46, 32'h42148d69, 32'h42507fe9, 32'hc1c85da6, 32'hc287603b, 32'h3f969e1e, 32'hc29aaae0};
test_output[3448] = '{32'h42bd1f46};
test_index[3448] = '{1};
test_input[27592:27599] = '{32'h428795fe, 32'h4204539f, 32'hc29dc72f, 32'hc25acab8, 32'h4228f7eb, 32'hc29ceb6a, 32'h3fc0460c, 32'hc29465ec};
test_output[3449] = '{32'h428795fe};
test_index[3449] = '{0};
test_input[27600:27607] = '{32'h42578a53, 32'h4093b536, 32'hc20291a9, 32'h4276cbbf, 32'hc25ecf71, 32'hc28e55ca, 32'hc2845f91, 32'h421fb9d3};
test_output[3450] = '{32'h4276cbbf};
test_index[3450] = '{3};
test_input[27608:27615] = '{32'h427b5677, 32'hc1bb1402, 32'hc2b5f464, 32'h4256ee2d, 32'h42a562ec, 32'h422306ac, 32'h42acaabe, 32'h42c0083a};
test_output[3451] = '{32'h42c0083a};
test_index[3451] = '{7};
test_input[27616:27623] = '{32'hc1aeeb93, 32'h42109295, 32'hc2a7ca01, 32'h42311c43, 32'hc25ba9d9, 32'h42573ee8, 32'hc132e23f, 32'hc141150a};
test_output[3452] = '{32'h42573ee8};
test_index[3452] = '{5};
test_input[27624:27631] = '{32'h423701e2, 32'hc2b96091, 32'hc22df316, 32'h42b0b1f5, 32'h41b1378f, 32'hc24af3fa, 32'h420c769e, 32'hc1f8d544};
test_output[3453] = '{32'h42b0b1f5};
test_index[3453] = '{3};
test_input[27632:27639] = '{32'hc1cbe5eb, 32'h4274507e, 32'h42949530, 32'h42b02837, 32'hc1fbd513, 32'h4285bf23, 32'hc2832ad2, 32'h41884c37};
test_output[3454] = '{32'h42b02837};
test_index[3454] = '{3};
test_input[27640:27647] = '{32'h4184abb7, 32'hc210c0b2, 32'hc24fd9ca, 32'hc28aa75c, 32'hc1b2c368, 32'hc2ac0ebe, 32'hc27e189c, 32'h42abcba4};
test_output[3455] = '{32'h42abcba4};
test_index[3455] = '{7};
test_input[27648:27655] = '{32'hc22ce9d6, 32'h42a18dcd, 32'hc29b0bc3, 32'h42bf24cf, 32'h41f3ee2e, 32'hc1dddc6e, 32'h42b2431d, 32'hc2b62da9};
test_output[3456] = '{32'h42bf24cf};
test_index[3456] = '{3};
test_input[27656:27663] = '{32'h4200412c, 32'h4227570e, 32'h41faab41, 32'hc284ea17, 32'h42944dc1, 32'h42c62bf7, 32'h42350570, 32'hc29cb75d};
test_output[3457] = '{32'h42c62bf7};
test_index[3457] = '{5};
test_input[27664:27671] = '{32'hc1107dca, 32'h424a2856, 32'h422c45d1, 32'h40304bde, 32'h4160d283, 32'h42272dac, 32'hc1af2f6c, 32'hc29db50d};
test_output[3458] = '{32'h424a2856};
test_index[3458] = '{1};
test_input[27672:27679] = '{32'h424bbf43, 32'h4285bab9, 32'hc17b6407, 32'h4281c724, 32'hc28b6a18, 32'hc249b518, 32'h41a10ed0, 32'hc0ae8c5e};
test_output[3459] = '{32'h4285bab9};
test_index[3459] = '{1};
test_input[27680:27687] = '{32'h421be09a, 32'hc228cb50, 32'h41088292, 32'h41e5a2b9, 32'h42a54614, 32'hc29b451e, 32'h4237356b, 32'hc22393a9};
test_output[3460] = '{32'h42a54614};
test_index[3460] = '{4};
test_input[27688:27695] = '{32'hc2665a6d, 32'hc27edc04, 32'hc0db8f9c, 32'h41f32717, 32'h42a15597, 32'hc29f3426, 32'hc1275ba6, 32'hc2893e86};
test_output[3461] = '{32'h42a15597};
test_index[3461] = '{4};
test_input[27696:27703] = '{32'hc2bed44d, 32'hc280e0a6, 32'hc2b7aed4, 32'hc2bc2513, 32'h429677bb, 32'h41c2bb75, 32'h42489919, 32'hc24d671c};
test_output[3462] = '{32'h429677bb};
test_index[3462] = '{4};
test_input[27704:27711] = '{32'h42343f59, 32'hc2adc992, 32'h428a32b0, 32'h4190f7ee, 32'hc2389548, 32'h42c27044, 32'h42aeda51, 32'h421b828b};
test_output[3463] = '{32'h42c27044};
test_index[3463] = '{5};
test_input[27712:27719] = '{32'h4253eccc, 32'hc29005bd, 32'hc0fe7697, 32'hc21a7ed1, 32'hc20ce0c7, 32'hc24ae6a1, 32'h413d653b, 32'hc2b50996};
test_output[3464] = '{32'h4253eccc};
test_index[3464] = '{0};
test_input[27720:27727] = '{32'h415b8f0c, 32'h4248f948, 32'h419684e8, 32'h422018d9, 32'h41211b5f, 32'hc1cac5d9, 32'h429541af, 32'h428d4551};
test_output[3465] = '{32'h429541af};
test_index[3465] = '{6};
test_input[27728:27735] = '{32'h42139f01, 32'h401e05fa, 32'hc288bd52, 32'hc1186611, 32'hc1f83278, 32'h4238cd39, 32'h414d9119, 32'h424a64cc};
test_output[3466] = '{32'h424a64cc};
test_index[3466] = '{7};
test_input[27736:27743] = '{32'hc1f5cf6a, 32'hc1302712, 32'hc24e11f6, 32'h4289dde5, 32'h41bb0756, 32'hc19386b6, 32'hc24fa09f, 32'hc26f0fc9};
test_output[3467] = '{32'h4289dde5};
test_index[3467] = '{3};
test_input[27744:27751] = '{32'hc2c329f1, 32'hc2aee47a, 32'hc2142b8b, 32'hc29c1f8e, 32'h41c14b12, 32'hc23192b8, 32'hc1965f89, 32'h42bdc6e8};
test_output[3468] = '{32'h42bdc6e8};
test_index[3468] = '{7};
test_input[27752:27759] = '{32'hc24471f3, 32'h42980e1c, 32'hc172366f, 32'hc1c148b0, 32'hc2558a49, 32'h424b4e07, 32'h410d48ac, 32'hc29e8efe};
test_output[3469] = '{32'h42980e1c};
test_index[3469] = '{1};
test_input[27760:27767] = '{32'h42972163, 32'hc182ee1b, 32'hc2632c2d, 32'h41c9e5a0, 32'hc12a2630, 32'hc212daba, 32'h427b89b2, 32'h42193efb};
test_output[3470] = '{32'h42972163};
test_index[3470] = '{0};
test_input[27768:27775] = '{32'h428658ac, 32'hc10b7f3e, 32'hc2ad9a21, 32'h420adeab, 32'hc1b81a53, 32'hc2b7857a, 32'h41f1d231, 32'hc24c7e57};
test_output[3471] = '{32'h428658ac};
test_index[3471] = '{0};
test_input[27776:27783] = '{32'h42a6f84e, 32'h429f170c, 32'h41919d18, 32'hc26f9d7b, 32'hc19f4696, 32'hc2b7c266, 32'h4298dae0, 32'hc28c13c1};
test_output[3472] = '{32'h42a6f84e};
test_index[3472] = '{0};
test_input[27784:27791] = '{32'hc2ab39a0, 32'hc1961192, 32'h429989dd, 32'h4232d133, 32'hc2695eb8, 32'h41786330, 32'h426402e2, 32'hc28cc2dc};
test_output[3473] = '{32'h429989dd};
test_index[3473] = '{2};
test_input[27792:27799] = '{32'hc2a01cad, 32'hc2c77e78, 32'h4268b5ff, 32'hc1474297, 32'h419225b4, 32'h41a8e9b4, 32'h41af9ca6, 32'h42b00d76};
test_output[3474] = '{32'h42b00d76};
test_index[3474] = '{7};
test_input[27800:27807] = '{32'h42877eb1, 32'h42744309, 32'h42b34631, 32'hc224ebba, 32'h413bbcf0, 32'h42b506c1, 32'h429ac484, 32'h421338df};
test_output[3475] = '{32'h42b506c1};
test_index[3475] = '{5};
test_input[27808:27815] = '{32'h428e952d, 32'h4265a020, 32'h41e3bae1, 32'hc2c1b96c, 32'hc259fa99, 32'hc28a10fa, 32'h42bdffad, 32'hc2af99e6};
test_output[3476] = '{32'h42bdffad};
test_index[3476] = '{6};
test_input[27816:27823] = '{32'hc29accb7, 32'h41ec7423, 32'h429f69a1, 32'h429a5b79, 32'h42b6ce8f, 32'h42627ded, 32'hc1ec4784, 32'h4280a61d};
test_output[3477] = '{32'h42b6ce8f};
test_index[3477] = '{4};
test_input[27824:27831] = '{32'hc2830111, 32'h424d06a4, 32'hc2899628, 32'h42b26175, 32'h4162c96a, 32'h4243dc61, 32'h4240148d, 32'hc2547a35};
test_output[3478] = '{32'h42b26175};
test_index[3478] = '{3};
test_input[27832:27839] = '{32'h41d49aa3, 32'h42a37619, 32'hc2b7ab35, 32'hc285eb93, 32'hc043b476, 32'h41ce3574, 32'h41b5c51b, 32'hc1c7224a};
test_output[3479] = '{32'h42a37619};
test_index[3479] = '{1};
test_input[27840:27847] = '{32'h42a4a68a, 32'hc0efcdeb, 32'h40c71837, 32'h425e0ff6, 32'h41bdae9f, 32'hc29b4906, 32'h42c7e630, 32'hc15c1dd4};
test_output[3480] = '{32'h42c7e630};
test_index[3480] = '{6};
test_input[27848:27855] = '{32'hc0d63829, 32'hc1e91292, 32'hc222a791, 32'h42265197, 32'hc24fec6b, 32'hc2c3896e, 32'hc2c56bec, 32'h418c6849};
test_output[3481] = '{32'h42265197};
test_index[3481] = '{3};
test_input[27856:27863] = '{32'h41e6cbe5, 32'hc2a0a292, 32'h4212d99b, 32'h42aa6e5c, 32'h4230c926, 32'h41fcc777, 32'hc2820024, 32'hc1bdcb45};
test_output[3482] = '{32'h42aa6e5c};
test_index[3482] = '{3};
test_input[27864:27871] = '{32'hc258d055, 32'h42b8d416, 32'hc2acf17b, 32'h429a0495, 32'hc29fb35b, 32'hc283eea9, 32'hc299dd9a, 32'h42a51837};
test_output[3483] = '{32'h42b8d416};
test_index[3483] = '{1};
test_input[27872:27879] = '{32'h411549cf, 32'h429f1298, 32'h41d4f7f4, 32'hc18d29a1, 32'h420dc6e3, 32'hc2c71de1, 32'h4229a6f1, 32'hc23fd34c};
test_output[3484] = '{32'h429f1298};
test_index[3484] = '{1};
test_input[27880:27887] = '{32'h41444518, 32'hc16a8fff, 32'hc2aca5c0, 32'hc2760725, 32'hc22f2f50, 32'h4291cb31, 32'h40ea2e62, 32'h42092b02};
test_output[3485] = '{32'h4291cb31};
test_index[3485] = '{5};
test_input[27888:27895] = '{32'hc1bfa16f, 32'h427441df, 32'h4210cd4c, 32'h42a33410, 32'h42993a13, 32'h42873e1d, 32'hc255e668, 32'h425e87b8};
test_output[3486] = '{32'h42a33410};
test_index[3486] = '{3};
test_input[27896:27903] = '{32'hc2b01ffe, 32'h41dcdc43, 32'hc09417ab, 32'h422ae5f4, 32'h420ecc63, 32'h42c26ae5, 32'h42a8c653, 32'h40d4c5b8};
test_output[3487] = '{32'h42c26ae5};
test_index[3487] = '{5};
test_input[27904:27911] = '{32'h42bfad2e, 32'h42a46687, 32'hc2a4b00c, 32'hc2635a97, 32'h429e6025, 32'h405b6487, 32'hc2909940, 32'hc2c18fdc};
test_output[3488] = '{32'h42bfad2e};
test_index[3488] = '{0};
test_input[27912:27919] = '{32'h42bee165, 32'h419f7488, 32'hc29e0928, 32'hc131e986, 32'hc2311717, 32'hc282814f, 32'hc2bc60d7, 32'h424c89ec};
test_output[3489] = '{32'h42bee165};
test_index[3489] = '{0};
test_input[27920:27927] = '{32'hc27c3325, 32'hc14991ad, 32'hc2b7fc28, 32'hc2a7ec70, 32'hc25ea842, 32'h41d1434d, 32'hc1a39f87, 32'h42996f0d};
test_output[3490] = '{32'h42996f0d};
test_index[3490] = '{7};
test_input[27928:27935] = '{32'h41865ac3, 32'h427e0a44, 32'h42028885, 32'hc2b42394, 32'hc1af48be, 32'h429cbca0, 32'h42403b8b, 32'h429f5877};
test_output[3491] = '{32'h429f5877};
test_index[3491] = '{7};
test_input[27936:27943] = '{32'h428fbc21, 32'hc26479c2, 32'hc1cbb6aa, 32'hc0dd0ea4, 32'h401def2d, 32'h42769a73, 32'hc220131f, 32'hc2a5e14e};
test_output[3492] = '{32'h428fbc21};
test_index[3492] = '{0};
test_input[27944:27951] = '{32'hc2c7f6a1, 32'h422e46df, 32'h421c156c, 32'h410067a4, 32'hc08edc20, 32'hc2c318f0, 32'hc2b19a3b, 32'hc1d1d4fe};
test_output[3493] = '{32'h422e46df};
test_index[3493] = '{1};
test_input[27952:27959] = '{32'hc2579506, 32'hc209c700, 32'hc2c7fcd4, 32'h42c432df, 32'hc1dcffde, 32'hc196774a, 32'hc267ef97, 32'hbf8414b0};
test_output[3494] = '{32'h42c432df};
test_index[3494] = '{3};
test_input[27960:27967] = '{32'h42895dde, 32'hc2409e7a, 32'h41e8c0f0, 32'h42a5c80e, 32'hc225388c, 32'h4291e3b9, 32'hc23a0f3e, 32'hc1cfb57f};
test_output[3495] = '{32'h42a5c80e};
test_index[3495] = '{3};
test_input[27968:27975] = '{32'h4281a3c9, 32'hc12de624, 32'h42848a1a, 32'h3fcebe03, 32'h421c38c7, 32'hc1ebc1c9, 32'h42446a1d, 32'h422eae12};
test_output[3496] = '{32'h42848a1a};
test_index[3496] = '{2};
test_input[27976:27983] = '{32'h429cf74c, 32'hc29c4962, 32'h41996480, 32'hc2340dca, 32'hc1723de0, 32'h416f8383, 32'hc2a97eef, 32'h428e3c0c};
test_output[3497] = '{32'h429cf74c};
test_index[3497] = '{0};
test_input[27984:27991] = '{32'hc1aecc5f, 32'hc134a804, 32'h429ceb3f, 32'h4233f68a, 32'hc16af5e3, 32'hc2a5529c, 32'h41ada588, 32'h424e8cac};
test_output[3498] = '{32'h429ceb3f};
test_index[3498] = '{2};
test_input[27992:27999] = '{32'hc265c0aa, 32'h42b231a7, 32'h42868735, 32'hc2968aed, 32'hc18cc9b2, 32'h42b7ab78, 32'h41bccd20, 32'hc299843d};
test_output[3499] = '{32'h42b7ab78};
test_index[3499] = '{5};
test_input[28000:28007] = '{32'h41bf2908, 32'h3d9e55a8, 32'h41dc2ea0, 32'hc2b083f5, 32'hc29e2028, 32'hc0a97b02, 32'hc22dcecb, 32'hc21808b8};
test_output[3500] = '{32'h41dc2ea0};
test_index[3500] = '{2};
test_input[28008:28015] = '{32'h428c2591, 32'hc236362c, 32'h409c86c1, 32'hc245011a, 32'hc28a6ae5, 32'hc2312bf2, 32'h4245606e, 32'h4249eae2};
test_output[3501] = '{32'h428c2591};
test_index[3501] = '{0};
test_input[28016:28023] = '{32'h42012a2b, 32'h42a663d0, 32'h424036eb, 32'hc2764c75, 32'h41094c46, 32'h42902cf3, 32'h424f7059, 32'h42b49f65};
test_output[3502] = '{32'h42b49f65};
test_index[3502] = '{7};
test_input[28024:28031] = '{32'hc2a66872, 32'hc29c90e9, 32'hc2b12ad1, 32'hc15bda24, 32'h4269cf14, 32'hc2111b55, 32'hc2805a9f, 32'hc1e48eb8};
test_output[3503] = '{32'h4269cf14};
test_index[3503] = '{4};
test_input[28032:28039] = '{32'h42b24ea2, 32'hc259b723, 32'hc222612f, 32'hc235c69f, 32'hc22150cb, 32'h42045aa9, 32'hc236ac38, 32'h4108c3f4};
test_output[3504] = '{32'h42b24ea2};
test_index[3504] = '{0};
test_input[28040:28047] = '{32'h42b5d65d, 32'h42500d00, 32'hc22977e1, 32'h400020a4, 32'h4174e50f, 32'h40ed63f3, 32'hc29ae807, 32'h4210cbd3};
test_output[3505] = '{32'h42b5d65d};
test_index[3505] = '{0};
test_input[28048:28055] = '{32'h41a9b04c, 32'hc132630d, 32'hc2b0144b, 32'hbffdce46, 32'hc274b928, 32'hc2395361, 32'h42ae1fe1, 32'h4108b51c};
test_output[3506] = '{32'h42ae1fe1};
test_index[3506] = '{6};
test_input[28056:28063] = '{32'hc1b4ee89, 32'hc27c2dd1, 32'hc2592e24, 32'hc108cf0a, 32'h4202f8bb, 32'hc2a27856, 32'hbf9a4de1, 32'h42bfe82a};
test_output[3507] = '{32'h42bfe82a};
test_index[3507] = '{7};
test_input[28064:28071] = '{32'h419ce2f0, 32'hc2803963, 32'hc17ec5a8, 32'h425c5a31, 32'hc2aaaa6c, 32'h41396e5c, 32'hc1ac1d0b, 32'hc2b3a4e7};
test_output[3508] = '{32'h425c5a31};
test_index[3508] = '{3};
test_input[28072:28079] = '{32'hc24966c7, 32'h4259806a, 32'hc25d7133, 32'hc2a61197, 32'h41dcb3ac, 32'h42b41a3b, 32'hc1c6dfcc, 32'h41042fde};
test_output[3509] = '{32'h42b41a3b};
test_index[3509] = '{5};
test_input[28080:28087] = '{32'hc12d4829, 32'h422d46cd, 32'hc282746a, 32'h413c9e18, 32'hc2b765ed, 32'h41aa0bf1, 32'h42324ae9, 32'hc25a948d};
test_output[3510] = '{32'h42324ae9};
test_index[3510] = '{6};
test_input[28088:28095] = '{32'hc274ee93, 32'hc2414166, 32'hc2128bd8, 32'h42a411e0, 32'hc24d7bf4, 32'h42a33925, 32'hc2b945fa, 32'h4273e3f9};
test_output[3511] = '{32'h42a411e0};
test_index[3511] = '{3};
test_input[28096:28103] = '{32'hc2b31d81, 32'hc0c4c885, 32'hc24324ce, 32'h42a7fe19, 32'hc27435c8, 32'hc0ddf6ef, 32'h42ae12fb, 32'hc24f573e};
test_output[3512] = '{32'h42ae12fb};
test_index[3512] = '{6};
test_input[28104:28111] = '{32'h41beef94, 32'h42ae4b34, 32'hc13ab3b6, 32'hc0b69b6d, 32'hc2bee6ed, 32'hc2c74627, 32'hbef227cd, 32'h42c63909};
test_output[3513] = '{32'h42c63909};
test_index[3513] = '{7};
test_input[28112:28119] = '{32'hc0a30ea6, 32'hc2a504e7, 32'hc2a7804b, 32'h41bf1ef3, 32'h41723106, 32'hc20c57a4, 32'hc2732386, 32'h429e52fc};
test_output[3514] = '{32'h429e52fc};
test_index[3514] = '{7};
test_input[28120:28127] = '{32'h4211234e, 32'hc2bf0c29, 32'hc195c2aa, 32'h4297077a, 32'hc28c1ae4, 32'h4165c0d8, 32'h416ffe60, 32'h41f79066};
test_output[3515] = '{32'h4297077a};
test_index[3515] = '{3};
test_input[28128:28135] = '{32'hc1a4a127, 32'hc14c4848, 32'h42343a12, 32'hc18e3f64, 32'h42b9b3b0, 32'h42807a86, 32'hc2a81ae6, 32'h426eb0d1};
test_output[3516] = '{32'h42b9b3b0};
test_index[3516] = '{4};
test_input[28136:28143] = '{32'hc2aeb478, 32'hbf2e6bc9, 32'h4238eac3, 32'hc1bf6e90, 32'hc1c36cc3, 32'hc21ff75a, 32'hc23dba06, 32'h428f0e36};
test_output[3517] = '{32'h428f0e36};
test_index[3517] = '{7};
test_input[28144:28151] = '{32'hc2a007ea, 32'h412e524a, 32'h41489790, 32'h4260e93c, 32'hc29da47c, 32'h425ca455, 32'h4279266c, 32'h4200cc7f};
test_output[3518] = '{32'h4279266c};
test_index[3518] = '{6};
test_input[28152:28159] = '{32'hc1961bc3, 32'h4228a150, 32'hc21cc9e5, 32'h42407c33, 32'hc1a20ac2, 32'hc275d5f1, 32'hc2835fd2, 32'hc225c1ad};
test_output[3519] = '{32'h42407c33};
test_index[3519] = '{3};
test_input[28160:28167] = '{32'hc2a15762, 32'h42a43a31, 32'h42c50926, 32'h41b35550, 32'hc1bc897a, 32'hc22bfea7, 32'h4220f7ce, 32'h419368c1};
test_output[3520] = '{32'h42c50926};
test_index[3520] = '{2};
test_input[28168:28175] = '{32'hc20bc0fb, 32'hc146023a, 32'h427290e3, 32'hc0f1455a, 32'hc174095e, 32'h415077b0, 32'hbeeec61d, 32'hc18574b5};
test_output[3521] = '{32'h427290e3};
test_index[3521] = '{2};
test_input[28176:28183] = '{32'hc2b46cb0, 32'hc120b610, 32'hc2c5ad9d, 32'hc2741735, 32'hc21049e9, 32'hc2a306d9, 32'hc17c3fda, 32'hc2325145};
test_output[3522] = '{32'hc120b610};
test_index[3522] = '{1};
test_input[28184:28191] = '{32'hc299b2b4, 32'hc2a0679b, 32'h4299d104, 32'hc297c0d0, 32'h42163d3d, 32'h415f7dd5, 32'hc27eaa66, 32'h42ab3d7a};
test_output[3523] = '{32'h42ab3d7a};
test_index[3523] = '{7};
test_input[28192:28199] = '{32'h41ef3e18, 32'h4285f7c7, 32'hc28d486b, 32'hc25430e3, 32'h41e0636b, 32'h42c02f37, 32'hc1f2e30c, 32'h42493ff0};
test_output[3524] = '{32'h42c02f37};
test_index[3524] = '{5};
test_input[28200:28207] = '{32'h41c51185, 32'hc293cda9, 32'h41e0b7a3, 32'hc2a780f1, 32'h42b284e5, 32'h42975674, 32'h42aa8ddf, 32'hc2905f89};
test_output[3525] = '{32'h42b284e5};
test_index[3525] = '{4};
test_input[28208:28215] = '{32'hc2540c87, 32'hc2957d08, 32'hc23b8399, 32'hc2ad6d3e, 32'h428f663e, 32'h420a2875, 32'hc0d0f0c2, 32'h40ec9dfe};
test_output[3526] = '{32'h428f663e};
test_index[3526] = '{4};
test_input[28216:28223] = '{32'hc2815346, 32'hc2a443d2, 32'h42487280, 32'h424e4217, 32'h4129a21e, 32'hc1510398, 32'hc01e3f51, 32'hc2b96d08};
test_output[3527] = '{32'h424e4217};
test_index[3527] = '{3};
test_input[28224:28231] = '{32'hc19f37a2, 32'h41e9aa7b, 32'h42a632aa, 32'hc1fa1741, 32'hc27a8332, 32'hc2adff2a, 32'h423522c6, 32'h42c5869f};
test_output[3528] = '{32'h42c5869f};
test_index[3528] = '{7};
test_input[28232:28239] = '{32'h4244e313, 32'hc278d7e1, 32'hc061e80d, 32'h41ed57ef, 32'hc0bcf787, 32'hc1efaa96, 32'h42be60f3, 32'h423de7e6};
test_output[3529] = '{32'h42be60f3};
test_index[3529] = '{6};
test_input[28240:28247] = '{32'h413d15c5, 32'h41d9e764, 32'h4216087b, 32'hc1e2893d, 32'hc2952667, 32'h4284d998, 32'hc29bd7fa, 32'h422b57c8};
test_output[3530] = '{32'h4284d998};
test_index[3530] = '{5};
test_input[28248:28255] = '{32'h42c5bcc9, 32'h42859ef1, 32'h429e486e, 32'hc2aabd9b, 32'h42ba5d68, 32'hc2535184, 32'hc164fab0, 32'h40b56c92};
test_output[3531] = '{32'h42c5bcc9};
test_index[3531] = '{0};
test_input[28256:28263] = '{32'h4289724d, 32'h428e88f5, 32'h42c6896e, 32'h4278e987, 32'h4182c61d, 32'hc2588799, 32'h42a3efee, 32'hc2c2ba55};
test_output[3532] = '{32'h42c6896e};
test_index[3532] = '{2};
test_input[28264:28271] = '{32'hc23fae5e, 32'hc1f78699, 32'h40286a9e, 32'h41389e8f, 32'hc2ac1cb8, 32'h4264bdf9, 32'h41b6b3b3, 32'hc2670290};
test_output[3533] = '{32'h4264bdf9};
test_index[3533] = '{5};
test_input[28272:28279] = '{32'h42883b1b, 32'hc2ac05ed, 32'hc2877a8c, 32'hc1ce573b, 32'h411f9dc8, 32'hc203fa2f, 32'h42012d8d, 32'h41d17b2a};
test_output[3534] = '{32'h42883b1b};
test_index[3534] = '{0};
test_input[28280:28287] = '{32'h4289fdad, 32'hc138de1a, 32'hc24c0123, 32'hbf6c7dc6, 32'h42c6f689, 32'hc2a8ee72, 32'hc116e2d3, 32'h417dafd0};
test_output[3535] = '{32'h42c6f689};
test_index[3535] = '{4};
test_input[28288:28295] = '{32'hc23abac0, 32'hc2b4a92d, 32'hc2c2e91a, 32'h42353932, 32'h42b099bd, 32'hc232332b, 32'h424387b6, 32'hc29fc9cd};
test_output[3536] = '{32'h42b099bd};
test_index[3536] = '{4};
test_input[28296:28303] = '{32'hc1157826, 32'hc164bbdb, 32'h426b949a, 32'h400fe749, 32'hc2822c7f, 32'hc22aa7ff, 32'h4087d2a7, 32'h41d03ea0};
test_output[3537] = '{32'h426b949a};
test_index[3537] = '{2};
test_input[28304:28311] = '{32'hc27a78d2, 32'h41bceb38, 32'hc27a98a7, 32'hc06b8f0b, 32'hc1fd4345, 32'h42563799, 32'hc2870565, 32'hc25a1a0b};
test_output[3538] = '{32'h42563799};
test_index[3538] = '{5};
test_input[28312:28319] = '{32'hc28306cb, 32'h4108cb09, 32'h427a740d, 32'h427598c3, 32'h41f03107, 32'hc1f4b534, 32'hc27bf801, 32'hc15fd8b3};
test_output[3539] = '{32'h427a740d};
test_index[3539] = '{2};
test_input[28320:28327] = '{32'h4078a7d5, 32'h41577ff4, 32'h41aaa98e, 32'h424297fc, 32'h428e338f, 32'h41aea913, 32'h426f01cd, 32'hc225b932};
test_output[3540] = '{32'h428e338f};
test_index[3540] = '{4};
test_input[28328:28335] = '{32'h4263e260, 32'h421eefd1, 32'hc28f8e9c, 32'h41f6bc5f, 32'hc14d28e5, 32'hc0099cc1, 32'hc27a4e8e, 32'h4260d776};
test_output[3541] = '{32'h4263e260};
test_index[3541] = '{0};
test_input[28336:28343] = '{32'h42581ab1, 32'h42ad57bc, 32'h428fa8ef, 32'hc1948a86, 32'h41ec762d, 32'hc28b66d2, 32'h42018343, 32'h4284e2ff};
test_output[3542] = '{32'h42ad57bc};
test_index[3542] = '{1};
test_input[28344:28351] = '{32'h4285fb8f, 32'hc2768f7a, 32'hc206ff82, 32'h3c50f0d4, 32'h4174cb8d, 32'hc2b3a73b, 32'hc2b96061, 32'h40940e6a};
test_output[3543] = '{32'h4285fb8f};
test_index[3543] = '{0};
test_input[28352:28359] = '{32'h408a105d, 32'hc23341ce, 32'hc291a0fc, 32'hc139e9e9, 32'hc2946d04, 32'h413f63dd, 32'hc239cf0b, 32'h421ae9fd};
test_output[3544] = '{32'h421ae9fd};
test_index[3544] = '{7};
test_input[28360:28367] = '{32'hc1e8609f, 32'hc2865def, 32'h422e1832, 32'hc265b1f2, 32'hc2044096, 32'hc29de495, 32'hc2615245, 32'hc22a9f04};
test_output[3545] = '{32'h422e1832};
test_index[3545] = '{2};
test_input[28368:28375] = '{32'h42bcb576, 32'h420f4251, 32'h40c75e8d, 32'hc2a376c4, 32'h425b4f1e, 32'hc2716817, 32'h428bc9cb, 32'h4248cc81};
test_output[3546] = '{32'h42bcb576};
test_index[3546] = '{0};
test_input[28376:28383] = '{32'h4198c0ed, 32'hc2a4848b, 32'hc1d5ec0c, 32'h4246aeda, 32'hc226c2f4, 32'h421790b2, 32'h4285aeb1, 32'hc2bc7470};
test_output[3547] = '{32'h4285aeb1};
test_index[3547] = '{6};
test_input[28384:28391] = '{32'h422f56e8, 32'hc2a400e1, 32'h42a63976, 32'h428d9ddd, 32'hc157a951, 32'h420bd563, 32'hc25516ef, 32'hc2c2bb8b};
test_output[3548] = '{32'h42a63976};
test_index[3548] = '{2};
test_input[28392:28399] = '{32'h40b13525, 32'hc1272f4c, 32'h42ae36cc, 32'h4217062c, 32'h42b8fc70, 32'hc2a24b24, 32'h42c6f77e, 32'hc265c702};
test_output[3549] = '{32'h42c6f77e};
test_index[3549] = '{6};
test_input[28400:28407] = '{32'h4161ec9e, 32'h4191d6db, 32'h4265836b, 32'hc285ab91, 32'hc15c9dde, 32'hc1a961e6, 32'hc2356f42, 32'hc25345ec};
test_output[3550] = '{32'h4265836b};
test_index[3550] = '{2};
test_input[28408:28415] = '{32'h42b349be, 32'h42849a02, 32'hbf5344c9, 32'hc2bd029f, 32'h42c24fdf, 32'hc2a92fab, 32'hc2aeff44, 32'h42aaee59};
test_output[3551] = '{32'h42c24fdf};
test_index[3551] = '{4};
test_input[28416:28423] = '{32'h425f81c2, 32'h42b3ce9e, 32'hbfb8566d, 32'h42c3ae89, 32'hc2aeb2f5, 32'h4267a8d6, 32'hc02d6daf, 32'hc22bfa3e};
test_output[3552] = '{32'h42c3ae89};
test_index[3552] = '{3};
test_input[28424:28431] = '{32'hc20bb05d, 32'h4255c8b1, 32'h42b6e02c, 32'hc27dcb23, 32'hc2c70d99, 32'hc1b2c997, 32'hc1c775a7, 32'h4230109f};
test_output[3553] = '{32'h42b6e02c};
test_index[3553] = '{2};
test_input[28432:28439] = '{32'hc2c1cbcb, 32'h411727a1, 32'hc2a872cb, 32'h421d22d4, 32'h4192fa86, 32'hc2be25b5, 32'hc299865f, 32'hc21b0391};
test_output[3554] = '{32'h421d22d4};
test_index[3554] = '{3};
test_input[28440:28447] = '{32'h42b04efd, 32'h42a0731d, 32'hbf9ffbcf, 32'hc01a485a, 32'h41d1e306, 32'h42a22b0a, 32'h418ca819, 32'hc196ed91};
test_output[3555] = '{32'h42b04efd};
test_index[3555] = '{0};
test_input[28448:28455] = '{32'h424ddbdf, 32'h425b8471, 32'h426f9451, 32'h42923222, 32'h426a7f9c, 32'hc21c3ace, 32'h402f0e32, 32'h425019e9};
test_output[3556] = '{32'h42923222};
test_index[3556] = '{3};
test_input[28456:28463] = '{32'hc2496e47, 32'h4017ab37, 32'h41930f60, 32'hc1a6cdb4, 32'h42477fd1, 32'hc22d3518, 32'hc20e0a8a, 32'hc2af1ced};
test_output[3557] = '{32'h42477fd1};
test_index[3557] = '{4};
test_input[28464:28471] = '{32'hc1e5f602, 32'h41dc8a65, 32'hc25f692f, 32'hc2694ef9, 32'hc2bc52b8, 32'hc1a1e9ca, 32'h422a16a7, 32'hc298e948};
test_output[3558] = '{32'h422a16a7};
test_index[3558] = '{6};
test_input[28472:28479] = '{32'hc263fc03, 32'h4224698f, 32'h41d65bb4, 32'h429212d9, 32'h42b82ebf, 32'hc1cf3eec, 32'h41ba4298, 32'hc2880e23};
test_output[3559] = '{32'h42b82ebf};
test_index[3559] = '{4};
test_input[28480:28487] = '{32'h42a7d22d, 32'h4210db09, 32'h42a9398d, 32'hc1740047, 32'h420c5ded, 32'hc285ef01, 32'h42ab046f, 32'h4249ea1e};
test_output[3560] = '{32'h42ab046f};
test_index[3560] = '{6};
test_input[28488:28495] = '{32'hc2b600b6, 32'h41cd149e, 32'h4226f9b5, 32'h42c17b20, 32'h425098bd, 32'h4245d813, 32'h42b41d63, 32'hc202fe7a};
test_output[3561] = '{32'h42c17b20};
test_index[3561] = '{3};
test_input[28496:28503] = '{32'h42448658, 32'hc2ada823, 32'hc29273a4, 32'hc281f6b6, 32'hc2241a27, 32'h420c8e6f, 32'h4295623e, 32'hc2732552};
test_output[3562] = '{32'h4295623e};
test_index[3562] = '{6};
test_input[28504:28511] = '{32'h4201166d, 32'h422689ee, 32'hc263e990, 32'hbf4e4cb0, 32'h42c1621c, 32'h42846c80, 32'h41ae656d, 32'h4254c95f};
test_output[3563] = '{32'h42c1621c};
test_index[3563] = '{4};
test_input[28512:28519] = '{32'hc08d0a72, 32'hc28bf013, 32'h41892c43, 32'hc2452732, 32'hc033916c, 32'hc28f9abc, 32'hc2556583, 32'h419e3d7a};
test_output[3564] = '{32'h419e3d7a};
test_index[3564] = '{7};
test_input[28520:28527] = '{32'h4290b1ad, 32'h422bceae, 32'h416b769d, 32'h4270bfa9, 32'hc1adbef0, 32'hc29c80f4, 32'h42419a7a, 32'h417b1be6};
test_output[3565] = '{32'h4290b1ad};
test_index[3565] = '{0};
test_input[28528:28535] = '{32'h41d626fc, 32'h3f7c71b9, 32'hc2a68ac3, 32'hc29ccd4a, 32'h403678de, 32'hc07a5e9e, 32'h4169b9d8, 32'hc28357ec};
test_output[3566] = '{32'h41d626fc};
test_index[3566] = '{0};
test_input[28536:28543] = '{32'h42c66615, 32'h424bf98b, 32'hc0b4e007, 32'hc2b5f356, 32'h42b75d27, 32'h42bc05f2, 32'hc2bb560c, 32'h42c264dd};
test_output[3567] = '{32'h42c66615};
test_index[3567] = '{0};
test_input[28544:28551] = '{32'hc127d9ec, 32'h418aa225, 32'h429f9689, 32'h42c792e5, 32'h42c7c53e, 32'hc2127adc, 32'h4286d94a, 32'h426a8bf1};
test_output[3568] = '{32'h42c7c53e};
test_index[3568] = '{4};
test_input[28552:28559] = '{32'h41d30b72, 32'h42278664, 32'h4245e52a, 32'h419b6da6, 32'hc1534066, 32'hc23148b9, 32'h41c25ae2, 32'h4246bd81};
test_output[3569] = '{32'h4246bd81};
test_index[3569] = '{7};
test_input[28560:28567] = '{32'h42455648, 32'hc138e0a2, 32'h42c724a1, 32'h406d8c5c, 32'hc2c790da, 32'hc2236f6e, 32'hc2a74d43, 32'hc247bf52};
test_output[3570] = '{32'h42c724a1};
test_index[3570] = '{2};
test_input[28568:28575] = '{32'h42366e0f, 32'h41ebae0b, 32'h40e73bde, 32'h40507cdc, 32'h422b767d, 32'hc25f99f7, 32'h42c7046e, 32'h411098c3};
test_output[3571] = '{32'h42c7046e};
test_index[3571] = '{6};
test_input[28576:28583] = '{32'hc103e7a2, 32'hc277156c, 32'hc2af5542, 32'h41ef3025, 32'h41fd4dcc, 32'h42b0258e, 32'hc1588cf2, 32'hc1aeb284};
test_output[3572] = '{32'h42b0258e};
test_index[3572] = '{5};
test_input[28584:28591] = '{32'hc27c8ad6, 32'hc2c70dd8, 32'hc151cfed, 32'hc2299c05, 32'hc29c99fb, 32'hc2ad85a3, 32'hbfe8f51b, 32'hc2c5f520};
test_output[3573] = '{32'hbfe8f51b};
test_index[3573] = '{6};
test_input[28592:28599] = '{32'hc2994aa5, 32'h421406d8, 32'h42b79366, 32'h41a6ccfc, 32'hc12b6fdc, 32'hc292ada5, 32'hc284fbc3, 32'hc2acbd1c};
test_output[3574] = '{32'h42b79366};
test_index[3574] = '{2};
test_input[28600:28607] = '{32'hbf0f1f00, 32'hc25e07ff, 32'h42609da8, 32'hc21ef56c, 32'h41dd012f, 32'hc2723d4a, 32'h42709a77, 32'h42780085};
test_output[3575] = '{32'h42780085};
test_index[3575] = '{7};
test_input[28608:28615] = '{32'hc21b765a, 32'hc1749c8d, 32'h4231bd93, 32'hc2256ee0, 32'h41a6629c, 32'h3fb57368, 32'h41be2980, 32'hc2abbe33};
test_output[3576] = '{32'h4231bd93};
test_index[3576] = '{2};
test_input[28616:28623] = '{32'h4234f0d2, 32'hc127bacf, 32'hc2a3e1d4, 32'hc221d846, 32'hc2004aca, 32'hc244cc69, 32'hc2acb8fa, 32'h424f7d23};
test_output[3577] = '{32'h424f7d23};
test_index[3577] = '{7};
test_input[28624:28631] = '{32'hc219e1b1, 32'h424e218a, 32'hc0ceb4df, 32'h42991260, 32'h427dfcd1, 32'h4274dbdd, 32'hc240f2cb, 32'h4178be58};
test_output[3578] = '{32'h42991260};
test_index[3578] = '{3};
test_input[28632:28639] = '{32'h42090f69, 32'hc2b4c540, 32'h428969f8, 32'h42b80ac2, 32'h4299e38f, 32'h41c95bee, 32'hc2861025, 32'hc1dd9f16};
test_output[3579] = '{32'h42b80ac2};
test_index[3579] = '{3};
test_input[28640:28647] = '{32'hc20da80b, 32'hc2b8f22a, 32'h4287612f, 32'h42b5b1be, 32'hc2b2516d, 32'hc269363f, 32'h3d8eacbb, 32'h4180bcc1};
test_output[3580] = '{32'h42b5b1be};
test_index[3580] = '{3};
test_input[28648:28655] = '{32'h424c2604, 32'h418d41a2, 32'h41bc8145, 32'h41e1e6d6, 32'h4239ec67, 32'h41a5c144, 32'h41104772, 32'hc26c33ec};
test_output[3581] = '{32'h424c2604};
test_index[3581] = '{0};
test_input[28656:28663] = '{32'hc22f8db5, 32'hc2375c79, 32'hc188d626, 32'h4248a1cf, 32'h42675735, 32'h41819c21, 32'h41cdd0af, 32'hc28a5e36};
test_output[3582] = '{32'h42675735};
test_index[3582] = '{4};
test_input[28664:28671] = '{32'hc1921ec0, 32'hc294d280, 32'hc28da60b, 32'hc270518c, 32'hc266ed04, 32'hc2b98327, 32'h42a78aa8, 32'hc25f4ef5};
test_output[3583] = '{32'h42a78aa8};
test_index[3583] = '{6};
test_input[28672:28679] = '{32'h42abf7cf, 32'h424d287a, 32'h42c7c967, 32'hc2af1887, 32'h4203508b, 32'h4205930e, 32'h42bb2252, 32'hc2615960};
test_output[3584] = '{32'h42c7c967};
test_index[3584] = '{2};
test_input[28680:28687] = '{32'hc2ab9511, 32'h428cd9b2, 32'hc2b0c453, 32'h42748493, 32'hc2293671, 32'hc1c67bc9, 32'hc18ed76d, 32'hc0aa3533};
test_output[3585] = '{32'h428cd9b2};
test_index[3585] = '{1};
test_input[28688:28695] = '{32'h428680f4, 32'h41265f8f, 32'h424bc6c0, 32'h3ea6a13a, 32'hc29595f9, 32'h42be0361, 32'hc2271623, 32'h41649e60};
test_output[3586] = '{32'h42be0361};
test_index[3586] = '{5};
test_input[28696:28703] = '{32'hc2b1e889, 32'h42aff3a1, 32'h4243d3c2, 32'h42a11614, 32'hc2236839, 32'h42205e3e, 32'h429e4c6c, 32'hc2bd8b42};
test_output[3587] = '{32'h42aff3a1};
test_index[3587] = '{1};
test_input[28704:28711] = '{32'hc2330243, 32'h42ad0556, 32'h421976a2, 32'h422ef3a5, 32'h42c41768, 32'h4253146a, 32'h42af31ac, 32'hc291a8c4};
test_output[3588] = '{32'h42c41768};
test_index[3588] = '{4};
test_input[28712:28719] = '{32'h42ba7eba, 32'hc180fad3, 32'hc201413c, 32'h42ac30db, 32'h421a7807, 32'hc2a037c0, 32'hc27282e8, 32'h4273a435};
test_output[3589] = '{32'h42ba7eba};
test_index[3589] = '{0};
test_input[28720:28727] = '{32'h4181c324, 32'h429fd6b1, 32'h427a26fd, 32'h423fc829, 32'hc2bccb1e, 32'h42483278, 32'hc2c76ddb, 32'h424b8e8a};
test_output[3590] = '{32'h429fd6b1};
test_index[3590] = '{1};
test_input[28728:28735] = '{32'h4292e1eb, 32'h42be51f0, 32'h41bcf29f, 32'hc26bf6da, 32'h42c11466, 32'hc26dde9a, 32'h42382450, 32'h42599864};
test_output[3591] = '{32'h42c11466};
test_index[3591] = '{4};
test_input[28736:28743] = '{32'h4230e5f8, 32'h413ebbfb, 32'h42b11aff, 32'hc2a8e9df, 32'hc2bf13e8, 32'hc2990217, 32'hc21d6951, 32'hc29021d9};
test_output[3592] = '{32'h42b11aff};
test_index[3592] = '{2};
test_input[28744:28751] = '{32'hbf84a8e0, 32'h4285bfe4, 32'h4293895f, 32'hc215cdb7, 32'h42388b7f, 32'hc241c687, 32'h41d33913, 32'hc24da97d};
test_output[3593] = '{32'h4293895f};
test_index[3593] = '{2};
test_input[28752:28759] = '{32'hc2aafbfe, 32'hc13bf69c, 32'hc2c7c2c8, 32'hc2862551, 32'h4296a4d9, 32'hc0bbfe8d, 32'hc20dd74b, 32'hc20388bd};
test_output[3594] = '{32'h4296a4d9};
test_index[3594] = '{4};
test_input[28760:28767] = '{32'hc18947ee, 32'h429d19f1, 32'h428a8b12, 32'h4281a702, 32'hc249fe27, 32'hc1c14fcf, 32'hc2b78303, 32'hc290a0df};
test_output[3595] = '{32'h429d19f1};
test_index[3595] = '{1};
test_input[28768:28775] = '{32'h4219290d, 32'hc2b935a7, 32'hc128f1d3, 32'hc21f9656, 32'hc1f5939d, 32'hc0a69252, 32'hc24ca0dd, 32'hc1b323f3};
test_output[3596] = '{32'h4219290d};
test_index[3596] = '{0};
test_input[28776:28783] = '{32'hc272b606, 32'h4290148f, 32'h42913e2a, 32'hc12e1f02, 32'h4285d679, 32'h4292225a, 32'h42727433, 32'hc12d6824};
test_output[3597] = '{32'h4292225a};
test_index[3597] = '{5};
test_input[28784:28791] = '{32'hc2656220, 32'h42899603, 32'h42b63bfc, 32'hc2abd73e, 32'hc2b9eb58, 32'hc088b929, 32'hc1597527, 32'hc2ab4303};
test_output[3598] = '{32'h42b63bfc};
test_index[3598] = '{2};
test_input[28792:28799] = '{32'h429c29ba, 32'h420af631, 32'hc19a7b86, 32'hc1033563, 32'hc2aed41d, 32'hc26557d6, 32'hc1819f8a, 32'h42716c72};
test_output[3599] = '{32'h429c29ba};
test_index[3599] = '{0};
test_input[28800:28807] = '{32'h413f4a43, 32'hc0fc35c4, 32'h428e04aa, 32'h42b5f1d9, 32'h42873009, 32'hc1cd0b69, 32'hc26403cb, 32'hc2048ff5};
test_output[3600] = '{32'h42b5f1d9};
test_index[3600] = '{3};
test_input[28808:28815] = '{32'h4211bf71, 32'h422242f4, 32'hc2bff823, 32'hc2bc446e, 32'h42ba76ce, 32'hc278208e, 32'hc23ad298, 32'h429ea80c};
test_output[3601] = '{32'h42ba76ce};
test_index[3601] = '{4};
test_input[28816:28823] = '{32'h42462475, 32'h4075e6f4, 32'hc1fca9a9, 32'hc2280a6f, 32'hc1c052c5, 32'hc0b70981, 32'h42a48dbb, 32'h42715423};
test_output[3602] = '{32'h42a48dbb};
test_index[3602] = '{6};
test_input[28824:28831] = '{32'hc2ae0d68, 32'h41fac0af, 32'hc26cc496, 32'h41c27142, 32'h42b5c423, 32'hc2a4aa98, 32'h42869fd8, 32'hc105f801};
test_output[3603] = '{32'h42b5c423};
test_index[3603] = '{4};
test_input[28832:28839] = '{32'hc2924334, 32'hc2b16680, 32'h42bd65c2, 32'h41a5c745, 32'hc1b142ba, 32'h428a456b, 32'h40fa03bb, 32'hc1b18ce3};
test_output[3604] = '{32'h42bd65c2};
test_index[3604] = '{2};
test_input[28840:28847] = '{32'hc17c6995, 32'h422f7106, 32'h410b7289, 32'h42091f01, 32'hc0a920b3, 32'hc2661041, 32'hc2a72499, 32'h422e676c};
test_output[3605] = '{32'h422f7106};
test_index[3605] = '{1};
test_input[28848:28855] = '{32'h42651189, 32'hc1712c51, 32'hc238372e, 32'h429b2831, 32'hc27f5cca, 32'hc2b74742, 32'hc1a09656, 32'h42272f5d};
test_output[3606] = '{32'h429b2831};
test_index[3606] = '{3};
test_input[28856:28863] = '{32'h4299d8fb, 32'h429b686f, 32'hc22a3f36, 32'h41f2066d, 32'hc2675d59, 32'h41e101db, 32'h420ca782, 32'hc1f5ea7c};
test_output[3607] = '{32'h429b686f};
test_index[3607] = '{1};
test_input[28864:28871] = '{32'h428b3325, 32'h42382d84, 32'h417e6fd3, 32'h4239b609, 32'h41471916, 32'h429701bd, 32'hc10e33a8, 32'hc0bc5357};
test_output[3608] = '{32'h429701bd};
test_index[3608] = '{5};
test_input[28872:28879] = '{32'h427fc930, 32'h4278c603, 32'hc2bd4553, 32'h40a61dfb, 32'h42b4eb6e, 32'hc06a01c5, 32'h41a7d941, 32'h42b738cf};
test_output[3609] = '{32'h42b738cf};
test_index[3609] = '{7};
test_input[28880:28887] = '{32'h42a3bb1f, 32'hc1569db3, 32'hc290a635, 32'h4235c691, 32'h42bdfd1f, 32'h4227ec65, 32'h42b626cc, 32'h41e95418};
test_output[3610] = '{32'h42bdfd1f};
test_index[3610] = '{4};
test_input[28888:28895] = '{32'h42257c1d, 32'hc2a65f59, 32'hc2770f9a, 32'h4215d6ce, 32'h426ab8d9, 32'h429f7f36, 32'h42c17d4a, 32'hc26e64c3};
test_output[3611] = '{32'h42c17d4a};
test_index[3611] = '{6};
test_input[28896:28903] = '{32'hc1d43b1d, 32'hc09efe3e, 32'h428ca685, 32'h42bf19e4, 32'h429de157, 32'h4260da09, 32'hbfc26970, 32'h4297dc2c};
test_output[3612] = '{32'h42bf19e4};
test_index[3612] = '{3};
test_input[28904:28911] = '{32'hc276fb86, 32'hc2b04a6a, 32'h40b501f9, 32'h3f3eb1b1, 32'hc22f7a5a, 32'h42c5bba0, 32'h426db24d, 32'hc2c4dd99};
test_output[3613] = '{32'h42c5bba0};
test_index[3613] = '{5};
test_input[28912:28919] = '{32'h42589b16, 32'h41897600, 32'h427b293a, 32'h4262216b, 32'h418c6ad5, 32'hc2b5155f, 32'hc2210f32, 32'h42bd85fe};
test_output[3614] = '{32'h42bd85fe};
test_index[3614] = '{7};
test_input[28920:28927] = '{32'hc2171432, 32'h42c12bb7, 32'h4233f898, 32'hc0385482, 32'hc208db2b, 32'h4251f87c, 32'hc2561701, 32'h42311e79};
test_output[3615] = '{32'h42c12bb7};
test_index[3615] = '{1};
test_input[28928:28935] = '{32'h41bc6c1a, 32'hc2545a4e, 32'h42873f7c, 32'h42b71ec1, 32'hc11d802d, 32'h42287e1e, 32'hc299960f, 32'h408c08ce};
test_output[3616] = '{32'h42b71ec1};
test_index[3616] = '{3};
test_input[28936:28943] = '{32'h424a5a5a, 32'h42832cf6, 32'hc2a533d7, 32'hc2c431f7, 32'hc221146e, 32'h423a6cfc, 32'h40aabad6, 32'hc0b3036c};
test_output[3617] = '{32'h42832cf6};
test_index[3617] = '{1};
test_input[28944:28951] = '{32'h424e57b0, 32'h42abfbed, 32'hc289f411, 32'h429db44c, 32'h421abadc, 32'h4214ae24, 32'hc1506f3d, 32'h4228260d};
test_output[3618] = '{32'h42abfbed};
test_index[3618] = '{1};
test_input[28952:28959] = '{32'hc2a030de, 32'hc278d36e, 32'hc2a4ac53, 32'h427a06ff, 32'hc19a87ff, 32'h42881a6e, 32'h418551a4, 32'hc21f7995};
test_output[3619] = '{32'h42881a6e};
test_index[3619] = '{5};
test_input[28960:28967] = '{32'h4222d605, 32'hc2711bd8, 32'hc213027f, 32'h425c26cc, 32'hc28ef1ba, 32'h4221d692, 32'h42abdedc, 32'h3f903fd1};
test_output[3620] = '{32'h42abdedc};
test_index[3620] = '{6};
test_input[28968:28975] = '{32'hc161d0ec, 32'h42a89381, 32'hc2976903, 32'h4226a435, 32'h429ac957, 32'h419426ec, 32'h42b69680, 32'h4217ec8b};
test_output[3621] = '{32'h42b69680};
test_index[3621] = '{6};
test_input[28976:28983] = '{32'hc2ab85c8, 32'hc2bf9bda, 32'hc2af554f, 32'h428c92a0, 32'h41f52301, 32'hc25c0807, 32'hc1ac69fc, 32'h4277ee2d};
test_output[3622] = '{32'h428c92a0};
test_index[3622] = '{3};
test_input[28984:28991] = '{32'hc2bf6de9, 32'h42659243, 32'h4014bf7a, 32'h42af94b8, 32'hc196a022, 32'h41bd8860, 32'hc18195a7, 32'h42915e57};
test_output[3623] = '{32'h42af94b8};
test_index[3623] = '{3};
test_input[28992:28999] = '{32'hc1000922, 32'h426b314c, 32'hc229bea3, 32'hc272d9bc, 32'hc1f9ec5a, 32'hc2bed60e, 32'h40bd8aaf, 32'hc23e236d};
test_output[3624] = '{32'h426b314c};
test_index[3624] = '{1};
test_input[29000:29007] = '{32'hc21a751b, 32'hc28c82dd, 32'h4113d845, 32'h3fe051c5, 32'hc2b6ed53, 32'h424c6c80, 32'h419a054f, 32'h42a08a98};
test_output[3625] = '{32'h42a08a98};
test_index[3625] = '{7};
test_input[29008:29015] = '{32'hc28f9b65, 32'hc1e26de4, 32'h427782ba, 32'hc2a408a4, 32'h426b210e, 32'h4268eb04, 32'h41bff5e8, 32'h42b3a498};
test_output[3626] = '{32'h42b3a498};
test_index[3626] = '{7};
test_input[29016:29023] = '{32'hc236cf64, 32'h421dc131, 32'hc2b24b9b, 32'h42bc32e4, 32'hc12e5751, 32'h42b9af83, 32'hc26c80a4, 32'hc22ed764};
test_output[3627] = '{32'h42bc32e4};
test_index[3627] = '{3};
test_input[29024:29031] = '{32'h420bf884, 32'hc1ea0371, 32'hc292d994, 32'h41b73b1d, 32'hc2003060, 32'hc2403ebb, 32'hc009fb70, 32'h423f8f42};
test_output[3628] = '{32'h423f8f42};
test_index[3628] = '{7};
test_input[29032:29039] = '{32'hc2a1fbed, 32'h413a5e46, 32'hc1e406c6, 32'h42b4bc4b, 32'h423bbc6d, 32'hc297f899, 32'hc25c84c0, 32'h40e1307e};
test_output[3629] = '{32'h42b4bc4b};
test_index[3629] = '{3};
test_input[29040:29047] = '{32'hc0e3e5a5, 32'hc2b133ca, 32'h4152dc65, 32'hc2a20af1, 32'h4205da0a, 32'hc26849d0, 32'h422d9387, 32'h42b12188};
test_output[3630] = '{32'h42b12188};
test_index[3630] = '{7};
test_input[29048:29055] = '{32'h425dbc39, 32'hc2324179, 32'hc19717a4, 32'hc2496646, 32'h429a4bd4, 32'h429180d8, 32'hc2a38a30, 32'h425ab53c};
test_output[3631] = '{32'h429a4bd4};
test_index[3631] = '{4};
test_input[29056:29063] = '{32'h4265d802, 32'hc29ff804, 32'h42859247, 32'h415f71ea, 32'hc1a79bd2, 32'hc293933f, 32'hc23c1538, 32'hc2a34da9};
test_output[3632] = '{32'h42859247};
test_index[3632] = '{2};
test_input[29064:29071] = '{32'h414d9b7e, 32'hc1319977, 32'h42bd91fa, 32'hc288bc5f, 32'h40e6a521, 32'h408590a4, 32'hc2acc384, 32'hc2a3a73f};
test_output[3633] = '{32'h42bd91fa};
test_index[3633] = '{2};
test_input[29072:29079] = '{32'h4209c6da, 32'hc28928cd, 32'h41566e9d, 32'h41f2f03b, 32'h4115869c, 32'hc285469a, 32'hc1447381, 32'h42742167};
test_output[3634] = '{32'h42742167};
test_index[3634] = '{7};
test_input[29080:29087] = '{32'h4291aee6, 32'h41d2894d, 32'hc2486499, 32'h42ae55d2, 32'hc097e06a, 32'h41af4d03, 32'hc2819790, 32'hbfebf099};
test_output[3635] = '{32'h42ae55d2};
test_index[3635] = '{3};
test_input[29088:29095] = '{32'h42134a8d, 32'hc263af62, 32'h42b67fe0, 32'h42a50416, 32'hc217980d, 32'hbf059045, 32'h4266958b, 32'hc180f459};
test_output[3636] = '{32'h42b67fe0};
test_index[3636] = '{2};
test_input[29096:29103] = '{32'hc11ca14e, 32'hc27df0f5, 32'hc1b69236, 32'h42c69c7b, 32'h4294ce95, 32'hc240563b, 32'hc220ec96, 32'hc21a7f97};
test_output[3637] = '{32'h42c69c7b};
test_index[3637] = '{3};
test_input[29104:29111] = '{32'h421dcf36, 32'hbec472a5, 32'h42a271ce, 32'hc147ddec, 32'h4218b14d, 32'hc2c2373a, 32'h42648ada, 32'h428e5e10};
test_output[3638] = '{32'h42a271ce};
test_index[3638] = '{2};
test_input[29112:29119] = '{32'h42a3fdab, 32'h4206a67b, 32'hc1c65ee6, 32'hc285616f, 32'hc2774fa4, 32'hc284a6d1, 32'h42654581, 32'h4143a660};
test_output[3639] = '{32'h42a3fdab};
test_index[3639] = '{0};
test_input[29120:29127] = '{32'h3fed12eb, 32'h4215b932, 32'hc2afa425, 32'h41eb1db0, 32'hc0f2c7d7, 32'hc2a5b382, 32'h4287f194, 32'hc28c22e7};
test_output[3640] = '{32'h4287f194};
test_index[3640] = '{6};
test_input[29128:29135] = '{32'hc1e42c69, 32'hc2b6db8b, 32'h4136c8ae, 32'hc1e9aeae, 32'h42a521d1, 32'hc23b9e8e, 32'h42b18702, 32'h422287db};
test_output[3641] = '{32'h42b18702};
test_index[3641] = '{6};
test_input[29136:29143] = '{32'h41957b29, 32'h416c0ef6, 32'h421d1207, 32'hc2bef1fe, 32'h424f78e2, 32'hc224316e, 32'hc2accd19, 32'h42098051};
test_output[3642] = '{32'h424f78e2};
test_index[3642] = '{4};
test_input[29144:29151] = '{32'h42669eb4, 32'hc294c95a, 32'hc299a2ea, 32'hc16c4c45, 32'hc14d88dd, 32'hc2b26ef4, 32'hc1e52ad8, 32'hc2c34b48};
test_output[3643] = '{32'h42669eb4};
test_index[3643] = '{0};
test_input[29152:29159] = '{32'h424107a5, 32'h42988da1, 32'h4233c26d, 32'h41cad06a, 32'hc16c3793, 32'hc1957ae5, 32'h42792f8a, 32'h421a99c6};
test_output[3644] = '{32'h42988da1};
test_index[3644] = '{1};
test_input[29160:29167] = '{32'h4162ba22, 32'hc2c48e50, 32'hc1b701d1, 32'h4160e52a, 32'hc1bb3983, 32'hc1eb3f51, 32'h428bda8b, 32'hc219db60};
test_output[3645] = '{32'h428bda8b};
test_index[3645] = '{6};
test_input[29168:29175] = '{32'h41f86962, 32'h41dba03e, 32'hc2b338de, 32'h42b0abc0, 32'h42199301, 32'hc1feb77f, 32'h41b2c0f7, 32'h4294dbcc};
test_output[3646] = '{32'h42b0abc0};
test_index[3646] = '{3};
test_input[29176:29183] = '{32'hc2bfff50, 32'h42a6192e, 32'h42144bce, 32'hc260df47, 32'hc13f715d, 32'h41d2ee11, 32'hc268d7d7, 32'h40033cb0};
test_output[3647] = '{32'h42a6192e};
test_index[3647] = '{1};
test_input[29184:29191] = '{32'hc28d2e53, 32'h4228d6ca, 32'hc2255cc7, 32'h42a6ce79, 32'hc1b6eeb0, 32'hc28dd4a1, 32'hc2c718a5, 32'hc2206ce3};
test_output[3648] = '{32'h42a6ce79};
test_index[3648] = '{3};
test_input[29192:29199] = '{32'hc1b315fc, 32'hc1c7d2ad, 32'h428d6b9f, 32'hc29ab69d, 32'hc1e3a0e0, 32'h4267cade, 32'h429a7cd9, 32'h419821c3};
test_output[3649] = '{32'h429a7cd9};
test_index[3649] = '{6};
test_input[29200:29207] = '{32'h4108f2a6, 32'hc2311e21, 32'hc236c0b8, 32'hc2038443, 32'h42c14cc5, 32'h420dfefa, 32'h422265e0, 32'hc2ad9627};
test_output[3650] = '{32'h42c14cc5};
test_index[3650] = '{4};
test_input[29208:29215] = '{32'hc2640f2d, 32'hc289b9ee, 32'h4290dc06, 32'hc15d1c18, 32'hbf3b03d9, 32'hc28c3018, 32'hc2a6a57a, 32'hc21d7551};
test_output[3651] = '{32'h4290dc06};
test_index[3651] = '{2};
test_input[29216:29223] = '{32'hc280483d, 32'h426aaa91, 32'h424b687a, 32'h415a8869, 32'hc169558c, 32'h406fd151, 32'h424a5c2c, 32'h41a24139};
test_output[3652] = '{32'h426aaa91};
test_index[3652] = '{1};
test_input[29224:29231] = '{32'hc164df4c, 32'hc1cc84d6, 32'hc27a0e9b, 32'hc2aff22d, 32'h40dfe01a, 32'h42a29d06, 32'h41c95fb6, 32'h42618942};
test_output[3653] = '{32'h42a29d06};
test_index[3653] = '{5};
test_input[29232:29239] = '{32'h42723e03, 32'h410ab284, 32'hc288782e, 32'hc2a35b95, 32'h42729e91, 32'hc2929571, 32'hc2b12dbc, 32'hc2ada5d7};
test_output[3654] = '{32'h42729e91};
test_index[3654] = '{4};
test_input[29240:29247] = '{32'h422c0cc1, 32'h42bd32e8, 32'h423f2202, 32'hc1e8e611, 32'hc1425382, 32'h42aee37b, 32'h42b79ca2, 32'h4209b2fa};
test_output[3655] = '{32'h42bd32e8};
test_index[3655] = '{1};
test_input[29248:29255] = '{32'h4213703c, 32'h421f914a, 32'hc2b518f3, 32'h418217b0, 32'h427e35a6, 32'h41d7282d, 32'hc2ba04ec, 32'h42808a56};
test_output[3656] = '{32'h42808a56};
test_index[3656] = '{7};
test_input[29256:29263] = '{32'h413a7713, 32'h41757674, 32'hc285786f, 32'h40b3b3b9, 32'hc1e142c1, 32'h400bd67d, 32'h42b3b3c0, 32'hc29053a6};
test_output[3657] = '{32'h42b3b3c0};
test_index[3657] = '{6};
test_input[29264:29271] = '{32'hc1be8834, 32'h4241cc83, 32'h424de252, 32'h42bcc817, 32'hc24f4ab1, 32'h428d0747, 32'hc286c234, 32'h42936b84};
test_output[3658] = '{32'h42bcc817};
test_index[3658] = '{3};
test_input[29272:29279] = '{32'h4274ddbf, 32'h42b1303e, 32'h42ae8e5c, 32'h42adca70, 32'h42af5f45, 32'hc1119e61, 32'h42ab6abb, 32'hc2282b07};
test_output[3659] = '{32'h42b1303e};
test_index[3659] = '{1};
test_input[29280:29287] = '{32'h42209ed1, 32'h42b9cced, 32'hc262fb86, 32'hc1996a06, 32'hc1813eeb, 32'hc1922493, 32'hc2046cf6, 32'hc20d86f1};
test_output[3660] = '{32'h42b9cced};
test_index[3660] = '{1};
test_input[29288:29295] = '{32'hc1f9177d, 32'hc2926a72, 32'h4230e86f, 32'h426de3e2, 32'h41677c52, 32'h41ecb18c, 32'h42b15653, 32'h41f06970};
test_output[3661] = '{32'h42b15653};
test_index[3661] = '{6};
test_input[29296:29303] = '{32'hc2bee464, 32'h42c0097a, 32'hbfce1f16, 32'hc2455733, 32'hc2b5cf99, 32'hc2b051f5, 32'hc2235f08, 32'h4239841d};
test_output[3662] = '{32'h42c0097a};
test_index[3662] = '{1};
test_input[29304:29311] = '{32'hc28005db, 32'h421b3723, 32'hc2a22eea, 32'hc23a997d, 32'h42afc109, 32'h41a91852, 32'h411999e2, 32'h42447ef0};
test_output[3663] = '{32'h42afc109};
test_index[3663] = '{4};
test_input[29312:29319] = '{32'hc1fe3857, 32'h428efecd, 32'hc11e10d3, 32'hc2859a3f, 32'h41bb146a, 32'hc28325b1, 32'h418dac34, 32'hc2a503e3};
test_output[3664] = '{32'h428efecd};
test_index[3664] = '{1};
test_input[29320:29327] = '{32'hc25dd9e4, 32'h4220b5e8, 32'hc22250f2, 32'h42b1e0a3, 32'h40a11be9, 32'hc276fff5, 32'hc24d2cbb, 32'h42b1cc3b};
test_output[3665] = '{32'h42b1e0a3};
test_index[3665] = '{3};
test_input[29328:29335] = '{32'hc1adda60, 32'hc1b5e665, 32'hc25f7bf7, 32'hc2b4bbaf, 32'h41720143, 32'h4189c264, 32'h425963dd, 32'h41cf0813};
test_output[3666] = '{32'h425963dd};
test_index[3666] = '{6};
test_input[29336:29343] = '{32'hc23f4a48, 32'h42a386b3, 32'h42c7dcf2, 32'h41cb1102, 32'h412fe403, 32'h420be315, 32'hc2347a5e, 32'h41f219ef};
test_output[3667] = '{32'h42c7dcf2};
test_index[3667] = '{2};
test_input[29344:29351] = '{32'h42b43dfa, 32'h428dc730, 32'hc28707a6, 32'hc1f765d8, 32'hc2b0b59f, 32'h4276dbfa, 32'h41a52633, 32'hc1afc70e};
test_output[3668] = '{32'h42b43dfa};
test_index[3668] = '{0};
test_input[29352:29359] = '{32'h41fcc689, 32'h4290a1de, 32'h4261b411, 32'h426f829e, 32'h42c41993, 32'h420f76ce, 32'hc20e8a66, 32'h42586cc5};
test_output[3669] = '{32'h42c41993};
test_index[3669] = '{4};
test_input[29360:29367] = '{32'h424ce917, 32'h4009c4e9, 32'hc23ee69c, 32'h41b8e6da, 32'h4292d04e, 32'hc22ac4cb, 32'hc2862415, 32'h41885455};
test_output[3670] = '{32'h4292d04e};
test_index[3670] = '{4};
test_input[29368:29375] = '{32'hbfd677b1, 32'hc2857024, 32'hc224c870, 32'h41552cb9, 32'h4222fb08, 32'h420c26e5, 32'hc2423c9f, 32'h4192ac07};
test_output[3671] = '{32'h4222fb08};
test_index[3671] = '{4};
test_input[29376:29383] = '{32'hc272803c, 32'h424734d8, 32'hc25f5026, 32'h4211a7f3, 32'hc2388708, 32'hc2368e3c, 32'hc1b663f9, 32'h419885a4};
test_output[3672] = '{32'h424734d8};
test_index[3672] = '{1};
test_input[29384:29391] = '{32'hc2aa55c8, 32'h42a466a7, 32'hc2367f6c, 32'h42c5ab0d, 32'h429a8841, 32'hc17caeb3, 32'hc1254247, 32'hc2a7a1b0};
test_output[3673] = '{32'h42c5ab0d};
test_index[3673] = '{3};
test_input[29392:29399] = '{32'h41b5ae9f, 32'h429564e9, 32'h42b4d636, 32'hc109c34c, 32'hc29455ae, 32'h4249a0f3, 32'hc2b13b45, 32'hc2b8be39};
test_output[3674] = '{32'h42b4d636};
test_index[3674] = '{2};
test_input[29400:29407] = '{32'h42ab29f7, 32'hc11c0c72, 32'hc28ef166, 32'h4279a511, 32'h40d833e4, 32'h42bda16b, 32'h4149dcd2, 32'hc20f0652};
test_output[3675] = '{32'h42bda16b};
test_index[3675] = '{5};
test_input[29408:29415] = '{32'h40e43ce0, 32'hc294f6c7, 32'h42aab685, 32'h41ae0543, 32'hc238ea20, 32'hc2c31ead, 32'h42bc1dd5, 32'hc2aec7e2};
test_output[3676] = '{32'h42bc1dd5};
test_index[3676] = '{6};
test_input[29416:29423] = '{32'hc1b13bda, 32'h42314dc7, 32'h4284d356, 32'h41caeb2a, 32'h428b1e00, 32'hc156383e, 32'hc2825842, 32'h4216e749};
test_output[3677] = '{32'h428b1e00};
test_index[3677] = '{4};
test_input[29424:29431] = '{32'hc263b994, 32'h429e3238, 32'hc273e618, 32'h41cb4b2e, 32'h42b3196d, 32'hc23d82f4, 32'hc25f2237, 32'hc2342c2f};
test_output[3678] = '{32'h42b3196d};
test_index[3678] = '{4};
test_input[29432:29439] = '{32'hc1bc75cd, 32'hc22aa53b, 32'h42b361bc, 32'hc0979e53, 32'h42999bf1, 32'h42c4ad9e, 32'h419c0092, 32'h4178580b};
test_output[3679] = '{32'h42c4ad9e};
test_index[3679] = '{5};
test_input[29440:29447] = '{32'hc29a7e44, 32'hc284f688, 32'hc22acb10, 32'h427e501e, 32'h425583f6, 32'h421f86e9, 32'h419286ed, 32'hc266555c};
test_output[3680] = '{32'h427e501e};
test_index[3680] = '{3};
test_input[29448:29455] = '{32'h42c26061, 32'h42c6718f, 32'hc165f3c0, 32'h418571f4, 32'hc1caf454, 32'h421cd262, 32'h42a9a9d2, 32'h42aee245};
test_output[3681] = '{32'h42c6718f};
test_index[3681] = '{1};
test_input[29456:29463] = '{32'hc29614f9, 32'hc189abbe, 32'hbfa0d5eb, 32'h419cf960, 32'h423277e3, 32'h41f5b661, 32'h429a24c1, 32'hc2070ced};
test_output[3682] = '{32'h429a24c1};
test_index[3682] = '{6};
test_input[29464:29471] = '{32'h4237b091, 32'h40fbfbda, 32'h42593339, 32'h422145fd, 32'hc2aa6728, 32'hc11fc802, 32'h41cb1eab, 32'hc205a7df};
test_output[3683] = '{32'h42593339};
test_index[3683] = '{2};
test_input[29472:29479] = '{32'h42a22838, 32'h42a50469, 32'hc24b5f0a, 32'h42181d9a, 32'h4266533f, 32'hc2878882, 32'h42ae2eed, 32'hbf8a1602};
test_output[3684] = '{32'h42ae2eed};
test_index[3684] = '{6};
test_input[29480:29487] = '{32'h41c60684, 32'hbfb0be04, 32'hc1bd555c, 32'h42c5feac, 32'hc22eea4d, 32'h429718eb, 32'hc2bf801d, 32'hc27022fb};
test_output[3685] = '{32'h42c5feac};
test_index[3685] = '{3};
test_input[29488:29495] = '{32'hc22bd212, 32'h40501412, 32'hc2ae153b, 32'hc1c0b529, 32'hc29c5644, 32'h429ebb05, 32'h42beb8ac, 32'hc223e0be};
test_output[3686] = '{32'h42beb8ac};
test_index[3686] = '{6};
test_input[29496:29503] = '{32'h42a577a7, 32'hc1b7eac3, 32'h4162c90f, 32'h422c8034, 32'hc1a061b8, 32'hc2a4fd90, 32'hc2a2eeda, 32'h4164b634};
test_output[3687] = '{32'h42a577a7};
test_index[3687] = '{0};
test_input[29504:29511] = '{32'h4232df5f, 32'hc1f745d4, 32'hc2a62093, 32'h426f8041, 32'hc0cf0269, 32'h42c66b62, 32'hc240e3e8, 32'h42bc22e5};
test_output[3688] = '{32'h42c66b62};
test_index[3688] = '{5};
test_input[29512:29519] = '{32'h41e473f5, 32'h420a2d2d, 32'hc1c80977, 32'h4254dfa5, 32'hc2b97bd3, 32'hc2258fab, 32'h421e024b, 32'hc23ab10c};
test_output[3689] = '{32'h4254dfa5};
test_index[3689] = '{3};
test_input[29520:29527] = '{32'hc2a8ae91, 32'h42871e31, 32'h4217ba76, 32'hc28cc484, 32'h422f7809, 32'hc1ab7b89, 32'h421ac2ef, 32'h421cbc1b};
test_output[3690] = '{32'h42871e31};
test_index[3690] = '{1};
test_input[29528:29535] = '{32'h420565bd, 32'hc18beecc, 32'h42867677, 32'h4247fd45, 32'h421af408, 32'hc208b034, 32'hc20f308b, 32'h42219205};
test_output[3691] = '{32'h42867677};
test_index[3691] = '{2};
test_input[29536:29543] = '{32'h413f348c, 32'hc2c60f21, 32'hc29c0ae1, 32'hc1ab4b94, 32'hc28c44b3, 32'h4293b840, 32'h42b9864e, 32'hc2abed18};
test_output[3692] = '{32'h42b9864e};
test_index[3692] = '{6};
test_input[29544:29551] = '{32'h40bb1417, 32'hc0a22614, 32'hc07dc85d, 32'h41c94c8c, 32'h421e9806, 32'hc227aa10, 32'h427b34a4, 32'hc07e3c43};
test_output[3693] = '{32'h427b34a4};
test_index[3693] = '{6};
test_input[29552:29559] = '{32'hc283a880, 32'h408381e9, 32'h4275c40e, 32'hc2a7a666, 32'h428c4dd8, 32'hc280eb41, 32'hc1d56376, 32'h41b3e1b2};
test_output[3694] = '{32'h428c4dd8};
test_index[3694] = '{4};
test_input[29560:29567] = '{32'hc2988e31, 32'h42c28e02, 32'hc1b1be30, 32'hc1fc0ca1, 32'h41af9def, 32'hc1b33d1c, 32'h3e791a2f, 32'hc198e4e4};
test_output[3695] = '{32'h42c28e02};
test_index[3695] = '{1};
test_input[29568:29575] = '{32'h42878fba, 32'h42815b35, 32'hc28b600c, 32'hc0d03653, 32'h40092cc6, 32'hc2b4f641, 32'hc239cea6, 32'hc2810bf1};
test_output[3696] = '{32'h42878fba};
test_index[3696] = '{0};
test_input[29576:29583] = '{32'h424e9bdc, 32'hc1f5d934, 32'h41d716da, 32'h3fba83f5, 32'hc1598167, 32'hbfd86739, 32'hc29f1aa0, 32'h41ac91d1};
test_output[3697] = '{32'h424e9bdc};
test_index[3697] = '{0};
test_input[29584:29591] = '{32'hbedcd655, 32'h42aaa29c, 32'h42581fdb, 32'hc2b5777f, 32'hc214dcae, 32'h4296af94, 32'h423c443f, 32'hc2c71257};
test_output[3698] = '{32'h42aaa29c};
test_index[3698] = '{1};
test_input[29592:29599] = '{32'hc15919ea, 32'hc2bdadee, 32'hc1b75ceb, 32'hc2b3da97, 32'hc20c6e8d, 32'hc26529e0, 32'hc20e427a, 32'hc1c8d0f0};
test_output[3699] = '{32'hc15919ea};
test_index[3699] = '{0};
test_input[29600:29607] = '{32'hc2b1c338, 32'h4192d934, 32'hc2393d85, 32'hc1b3d5d4, 32'h4241c3dd, 32'h42aacfb0, 32'hc260aa77, 32'h41a1ca48};
test_output[3700] = '{32'h42aacfb0};
test_index[3700] = '{5};
test_input[29608:29615] = '{32'hc1a5d00c, 32'hc20c5052, 32'hc16604a0, 32'hc2916c55, 32'hc223b926, 32'hc2279b7a, 32'h4191e233, 32'h42a20bf4};
test_output[3701] = '{32'h42a20bf4};
test_index[3701] = '{7};
test_input[29616:29623] = '{32'hc2abe004, 32'h41c64efd, 32'hc26b7f28, 32'hc1a008ac, 32'h428eb0d2, 32'hc1934e29, 32'hc11cccf2, 32'h42726176};
test_output[3702] = '{32'h428eb0d2};
test_index[3702] = '{4};
test_input[29624:29631] = '{32'h42b2aabb, 32'h40bf780b, 32'hc239a5e4, 32'h429b9b06, 32'hc205dee8, 32'hc2846e8f, 32'hc2499951, 32'h41018ce2};
test_output[3703] = '{32'h42b2aabb};
test_index[3703] = '{0};
test_input[29632:29639] = '{32'h4222aa70, 32'h4150176a, 32'h42bbea12, 32'hc2aa220b, 32'h42071531, 32'hc231c3be, 32'hc2a5d8d5, 32'h4265bbb3};
test_output[3704] = '{32'h42bbea12};
test_index[3704] = '{2};
test_input[29640:29647] = '{32'hc28dbd63, 32'hc21b055a, 32'h426762ac, 32'hc28fa1ba, 32'hc236fcb9, 32'hc2c7ac16, 32'h42ae70d6, 32'h41f7b910};
test_output[3705] = '{32'h42ae70d6};
test_index[3705] = '{6};
test_input[29648:29655] = '{32'h428fabcd, 32'h42b92078, 32'h41b5ef6b, 32'h4275ae89, 32'hc2c3e689, 32'h4187721d, 32'hc1993ac5, 32'hc1f8269d};
test_output[3706] = '{32'h42b92078};
test_index[3706] = '{1};
test_input[29656:29663] = '{32'hc2b04dd8, 32'h42523cb1, 32'h4240d10a, 32'h424e0105, 32'h4282a1d9, 32'hc00f65ca, 32'h42bde3ff, 32'hc2a08638};
test_output[3707] = '{32'h42bde3ff};
test_index[3707] = '{6};
test_input[29664:29671] = '{32'h42c36aab, 32'h41d7fde5, 32'hc1acf108, 32'hc2bc29be, 32'h4256a226, 32'h42a29247, 32'hc28a9001, 32'hc19145bd};
test_output[3708] = '{32'h42c36aab};
test_index[3708] = '{0};
test_input[29672:29679] = '{32'h419cc459, 32'hc2ae521d, 32'h41050b0f, 32'hc0d6185b, 32'h4298759a, 32'h420cd780, 32'hc1ebc162, 32'h4284fde7};
test_output[3709] = '{32'h4298759a};
test_index[3709] = '{4};
test_input[29680:29687] = '{32'h42b194eb, 32'h42a78650, 32'h42a27a7f, 32'h42356e3e, 32'hc285fa5a, 32'h42c70661, 32'hc2be5928, 32'h42b6d485};
test_output[3710] = '{32'h42c70661};
test_index[3710] = '{5};
test_input[29688:29695] = '{32'hc28a9373, 32'h4015cd8d, 32'hc1164636, 32'hc223a3e1, 32'hc2a8e102, 32'h42765e8c, 32'h4261e849, 32'hc297f633};
test_output[3711] = '{32'h42765e8c};
test_index[3711] = '{5};
test_input[29696:29703] = '{32'h426997b6, 32'hc0f54f6a, 32'hc2ab6d8a, 32'hc13b70a4, 32'hc0322976, 32'h429308d1, 32'h422ec18e, 32'h429b84e9};
test_output[3712] = '{32'h429b84e9};
test_index[3712] = '{7};
test_input[29704:29711] = '{32'hc2b57629, 32'h42be0ff9, 32'hbf893bcd, 32'h4237e538, 32'h42b2ca4a, 32'h42a85029, 32'h42048dee, 32'h4297110e};
test_output[3713] = '{32'h42be0ff9};
test_index[3713] = '{1};
test_input[29712:29719] = '{32'hc21cb157, 32'h41cfdb00, 32'hc1276440, 32'h429e64d8, 32'hc2b1d95d, 32'h41eac69c, 32'h40ab5056, 32'hc21482b5};
test_output[3714] = '{32'h429e64d8};
test_index[3714] = '{3};
test_input[29720:29727] = '{32'hbece20f1, 32'h42792d7b, 32'hc280c8ba, 32'h42adea65, 32'h404c0590, 32'h42326658, 32'h42afb03a, 32'hc118dbd5};
test_output[3715] = '{32'h42afb03a};
test_index[3715] = '{6};
test_input[29728:29735] = '{32'hc0b5083e, 32'hbf8a7e36, 32'hc24108e0, 32'hc1afce55, 32'hc114b788, 32'hc20e6b67, 32'hc23bef91, 32'hc2ab3da9};
test_output[3716] = '{32'hbf8a7e36};
test_index[3716] = '{1};
test_input[29736:29743] = '{32'hc20d76a2, 32'hc232b2ca, 32'h42c090b3, 32'h4254d350, 32'h421236fe, 32'hc2af04e5, 32'hc2a55364, 32'h422db726};
test_output[3717] = '{32'h42c090b3};
test_index[3717] = '{2};
test_input[29744:29751] = '{32'h4011dec3, 32'h41120adc, 32'h41730b8d, 32'h42bd48ed, 32'h42b1a446, 32'hc0054508, 32'h42c41d9e, 32'h414aac4e};
test_output[3718] = '{32'h42c41d9e};
test_index[3718] = '{6};
test_input[29752:29759] = '{32'h42655d8d, 32'h4299c8ef, 32'hc2a62441, 32'hc2c5430e, 32'h41bf2914, 32'hc293c088, 32'hc184c0fa, 32'hc18a2542};
test_output[3719] = '{32'h4299c8ef};
test_index[3719] = '{1};
test_input[29760:29767] = '{32'hc1bcd630, 32'h42801e33, 32'h40b163a9, 32'hc188a975, 32'h41d376fd, 32'h42b30b8e, 32'hc2c2222e, 32'hc28076c0};
test_output[3720] = '{32'h42b30b8e};
test_index[3720] = '{5};
test_input[29768:29775] = '{32'hc281f428, 32'hc28e0fc1, 32'h42aaabf5, 32'hc2b990e1, 32'hc21c73fd, 32'h421246ec, 32'hc2410a70, 32'h42ab5d2b};
test_output[3721] = '{32'h42ab5d2b};
test_index[3721] = '{7};
test_input[29776:29783] = '{32'hc108104e, 32'hc27c4b58, 32'h42407a20, 32'h42c3cc7c, 32'h41efad6d, 32'h405a4e44, 32'h420326bd, 32'hc25c384c};
test_output[3722] = '{32'h42c3cc7c};
test_index[3722] = '{3};
test_input[29784:29791] = '{32'h41ce62b3, 32'hc25261b1, 32'h42717d48, 32'h3fa1cda8, 32'h429e8ebb, 32'hc1f59431, 32'h42bf2a2e, 32'h428d177e};
test_output[3723] = '{32'h42bf2a2e};
test_index[3723] = '{6};
test_input[29792:29799] = '{32'h42bd303a, 32'h4229425b, 32'hc29eb1c4, 32'h41babe72, 32'h41cb6e65, 32'h429986d3, 32'h424f1216, 32'hc28d6947};
test_output[3724] = '{32'h42bd303a};
test_index[3724] = '{0};
test_input[29800:29807] = '{32'hc089e9dc, 32'hc26a23eb, 32'h42acd2a1, 32'h42084f10, 32'hc294f62e, 32'h426d9d0d, 32'h429f2595, 32'h42745506};
test_output[3725] = '{32'h42acd2a1};
test_index[3725] = '{2};
test_input[29808:29815] = '{32'hc1ed5f0d, 32'h42898706, 32'hc13a5d93, 32'h42b40e92, 32'hc18a3293, 32'h41ef4af4, 32'h428d5190, 32'h42561f53};
test_output[3726] = '{32'h42b40e92};
test_index[3726] = '{3};
test_input[29816:29823] = '{32'h42b6e3a0, 32'h413cd7ea, 32'h42bb9466, 32'hc0db2265, 32'h42c47f85, 32'h42bc1875, 32'hc2bfaee3, 32'h42c271da};
test_output[3727] = '{32'h42c47f85};
test_index[3727] = '{4};
test_input[29824:29831] = '{32'hc2886b52, 32'hc2a748ac, 32'hc01023be, 32'h41ba3837, 32'h42413ed5, 32'hc0ec427b, 32'h423f895b, 32'hc27a8016};
test_output[3728] = '{32'h42413ed5};
test_index[3728] = '{4};
test_input[29832:29839] = '{32'hc257f30a, 32'h4250c7e4, 32'h428ace8f, 32'h41b03f4f, 32'hc16f28f3, 32'hc29c88f6, 32'hc29effd4, 32'hc2c207b7};
test_output[3729] = '{32'h428ace8f};
test_index[3729] = '{2};
test_input[29840:29847] = '{32'h4208397b, 32'hc206861c, 32'h41c1e3fd, 32'h41b41c56, 32'hc298705b, 32'h4238bccb, 32'h42bbd593, 32'h422122d0};
test_output[3730] = '{32'h42bbd593};
test_index[3730] = '{6};
test_input[29848:29855] = '{32'hc297876d, 32'hc2844328, 32'h41bf8806, 32'h411952ff, 32'h424c8c4b, 32'h4142abc2, 32'h428e3a59, 32'hc29d4dd8};
test_output[3731] = '{32'h428e3a59};
test_index[3731] = '{6};
test_input[29856:29863] = '{32'h429b4b46, 32'h427ead18, 32'hc26e7b4a, 32'hc2943209, 32'h40bd7c06, 32'h424f5cc8, 32'hc2a54f5a, 32'h3fb749f5};
test_output[3732] = '{32'h429b4b46};
test_index[3732] = '{0};
test_input[29864:29871] = '{32'hc20e2970, 32'hc1cb694c, 32'hc1ced0be, 32'hc25f0bfa, 32'h4132f093, 32'h4281e372, 32'hc0682c79, 32'hc151b7c1};
test_output[3733] = '{32'h4281e372};
test_index[3733] = '{5};
test_input[29872:29879] = '{32'h4286fcec, 32'hc2bad6f0, 32'h42805a40, 32'hc2c69e11, 32'hc2b9984b, 32'h4218d81d, 32'h41ece5f7, 32'h4283f604};
test_output[3734] = '{32'h4286fcec};
test_index[3734] = '{0};
test_input[29880:29887] = '{32'h42a03bb7, 32'h42b12992, 32'hc28c4721, 32'h42b49d12, 32'h419db06f, 32'h4246eb93, 32'hc13a7ea2, 32'h42326a0f};
test_output[3735] = '{32'h42b49d12};
test_index[3735] = '{3};
test_input[29888:29895] = '{32'hc2482796, 32'hc2a54ab6, 32'hc1bc12bf, 32'h421bc616, 32'h41f58f1e, 32'h42a2da2b, 32'h42348857, 32'h42bff77e};
test_output[3736] = '{32'h42bff77e};
test_index[3736] = '{7};
test_input[29896:29903] = '{32'h411a849a, 32'hc1f1bade, 32'hc20f4859, 32'hc22f64f1, 32'hc138fd32, 32'h42138033, 32'hc295f9af, 32'hc25bf519};
test_output[3737] = '{32'h42138033};
test_index[3737] = '{5};
test_input[29904:29911] = '{32'h42be132f, 32'hc22d80f0, 32'h42c0b530, 32'hc26adb45, 32'hc081b6cc, 32'h4228b202, 32'h41bef982, 32'h429453d2};
test_output[3738] = '{32'h42c0b530};
test_index[3738] = '{2};
test_input[29912:29919] = '{32'h42afae74, 32'h42b3cc6c, 32'h3f6b9b70, 32'h4298fb3a, 32'hc2aa47d4, 32'hc08dfdac, 32'h424781ee, 32'h41444eb5};
test_output[3739] = '{32'h42b3cc6c};
test_index[3739] = '{1};
test_input[29920:29927] = '{32'hc2b887a3, 32'hc28b673e, 32'hc21272dd, 32'h4256a112, 32'hc265b33c, 32'h41e143b4, 32'hc0957d3e, 32'hc29e49ff};
test_output[3740] = '{32'h4256a112};
test_index[3740] = '{3};
test_input[29928:29935] = '{32'h42c4203b, 32'h42aab018, 32'hc181c0a2, 32'hc1e94556, 32'h421a2d02, 32'hc2b058bb, 32'hc2a37b30, 32'h41eb5217};
test_output[3741] = '{32'h42c4203b};
test_index[3741] = '{0};
test_input[29936:29943] = '{32'h41c90036, 32'h3f34c4bc, 32'h4241d718, 32'hc1b68aca, 32'h42559b77, 32'h42a32044, 32'hc2121946, 32'hc2248a81};
test_output[3742] = '{32'h42a32044};
test_index[3742] = '{5};
test_input[29944:29951] = '{32'h429fd6bc, 32'h420c5548, 32'h4298fcb7, 32'h4292fb18, 32'h42807975, 32'hc28942e2, 32'hc12cb174, 32'hc1446f0b};
test_output[3743] = '{32'h429fd6bc};
test_index[3743] = '{0};
test_input[29952:29959] = '{32'hc1970cc3, 32'h420fa276, 32'hc2007fd3, 32'hc2b53406, 32'hc2338011, 32'hc20eff68, 32'h42c52be4, 32'h41688bf3};
test_output[3744] = '{32'h42c52be4};
test_index[3744] = '{6};
test_input[29960:29967] = '{32'hc291bf10, 32'hc28fa852, 32'hc2912943, 32'h421d627e, 32'hc20ba923, 32'hc26c4666, 32'hc292cc6e, 32'hc217b653};
test_output[3745] = '{32'h421d627e};
test_index[3745] = '{3};
test_input[29968:29975] = '{32'h41b5cca2, 32'hc090ee18, 32'hc2971d25, 32'h427e6e22, 32'h427d0f03, 32'hc228b4c5, 32'h42c3e314, 32'h42ac75f4};
test_output[3746] = '{32'h42c3e314};
test_index[3746] = '{6};
test_input[29976:29983] = '{32'hc2927b94, 32'hc229d157, 32'hc013396d, 32'hc270ecb3, 32'h42650d6a, 32'hc2453bed, 32'hc2af9886, 32'hc2082cf0};
test_output[3747] = '{32'h42650d6a};
test_index[3747] = '{4};
test_input[29984:29991] = '{32'hc25d0dd1, 32'hc22a26a2, 32'hc2bf3822, 32'hc2b32a51, 32'h41b19da2, 32'h4281b420, 32'hc1af2cbe, 32'hc2886c11};
test_output[3748] = '{32'h4281b420};
test_index[3748] = '{5};
test_input[29992:29999] = '{32'h42701eff, 32'h413e6cc9, 32'hc20f7279, 32'hc251f865, 32'h427d41e7, 32'hc224f9dd, 32'hc237d6e4, 32'h42a88bfd};
test_output[3749] = '{32'h42a88bfd};
test_index[3749] = '{7};
test_input[30000:30007] = '{32'h429a51da, 32'h42b99f7b, 32'hc2c7ca81, 32'hc29f1caf, 32'hc2712614, 32'hc28d09d1, 32'hc29b6a24, 32'hc2545257};
test_output[3750] = '{32'h42b99f7b};
test_index[3750] = '{1};
test_input[30008:30015] = '{32'h428567ee, 32'hc24ec11c, 32'h41d31452, 32'h42bd4377, 32'hc2011c1c, 32'hc27df55c, 32'h3e3a97aa, 32'hc2839bb2};
test_output[3751] = '{32'h42bd4377};
test_index[3751] = '{3};
test_input[30016:30023] = '{32'hc2a8b3ea, 32'h42ba9fc7, 32'h41bc3d3d, 32'h425b1ed8, 32'h4264d8dd, 32'h4232a594, 32'hc1e196ec, 32'h421baae7};
test_output[3752] = '{32'h42ba9fc7};
test_index[3752] = '{1};
test_input[30024:30031] = '{32'hbfc6923f, 32'hc2b4665a, 32'h413d6093, 32'h41f645b9, 32'hc2064d84, 32'hc23aad45, 32'hc2c4013f, 32'hc28e27e7};
test_output[3753] = '{32'h41f645b9};
test_index[3753] = '{3};
test_input[30032:30039] = '{32'h41e47a90, 32'hc2580970, 32'h411fde4f, 32'hc1b7a4d5, 32'h413aaf5f, 32'hc21caf26, 32'h425f5b68, 32'hc1882ff2};
test_output[3754] = '{32'h425f5b68};
test_index[3754] = '{6};
test_input[30040:30047] = '{32'hc1ba4f71, 32'hc170eabc, 32'hc22584dc, 32'h3fcda795, 32'h41a41106, 32'h4215215d, 32'h41a6d95e, 32'hc09feed5};
test_output[3755] = '{32'h4215215d};
test_index[3755] = '{5};
test_input[30048:30055] = '{32'hc25b968d, 32'hc1fc4ce1, 32'hc2601d38, 32'hc2551962, 32'hc160972b, 32'h42acac68, 32'hc165722b, 32'hc10ec326};
test_output[3756] = '{32'h42acac68};
test_index[3756] = '{5};
test_input[30056:30063] = '{32'hc23d578d, 32'hc2abff54, 32'h423f2e1e, 32'h42a663dd, 32'hc21e7eae, 32'hc2632d87, 32'h42569456, 32'hc239160f};
test_output[3757] = '{32'h42a663dd};
test_index[3757] = '{3};
test_input[30064:30071] = '{32'hc20ad69c, 32'hc1e29fb5, 32'hc2149e92, 32'h429b2c5f, 32'h3fb18392, 32'h42c65100, 32'hc0a1b946, 32'h41bbc175};
test_output[3758] = '{32'h42c65100};
test_index[3758] = '{5};
test_input[30072:30079] = '{32'h42b59dd0, 32'h42b6f7d4, 32'hc1c5b236, 32'hc2a0dc71, 32'hc2bc1b60, 32'h42bc9c53, 32'hc21b24e8, 32'h422396be};
test_output[3759] = '{32'h42bc9c53};
test_index[3759] = '{5};
test_input[30080:30087] = '{32'hc2859302, 32'hc23f3978, 32'h4024cebd, 32'hc1faef13, 32'h42c152ae, 32'h42984e3d, 32'h42b3649b, 32'h420d4d6a};
test_output[3760] = '{32'h42c152ae};
test_index[3760] = '{4};
test_input[30088:30095] = '{32'h4267b033, 32'h3f2c0e2d, 32'h428fe08a, 32'hc298f7a4, 32'hc1cd66e5, 32'hc2a09b3f, 32'hc1953683, 32'h42c5beba};
test_output[3761] = '{32'h42c5beba};
test_index[3761] = '{7};
test_input[30096:30103] = '{32'h41c15562, 32'h41f863c4, 32'hc27f7449, 32'h425e06e5, 32'h42a5f469, 32'hc2ad4ed6, 32'h42aac379, 32'h42ab07ff};
test_output[3762] = '{32'h42ab07ff};
test_index[3762] = '{7};
test_input[30104:30111] = '{32'h41a98ccf, 32'hc2b0f188, 32'hc2385d8a, 32'hc1db1be7, 32'hc261c870, 32'hc1af383b, 32'h42a78523, 32'h428de621};
test_output[3763] = '{32'h42a78523};
test_index[3763] = '{6};
test_input[30112:30119] = '{32'hc2bbca67, 32'h4230faad, 32'h42b8832f, 32'hc1d0246c, 32'hc28b3517, 32'h42900163, 32'h42b1e0ef, 32'h42adeb9a};
test_output[3764] = '{32'h42b8832f};
test_index[3764] = '{2};
test_input[30120:30127] = '{32'hc24b07e9, 32'hc2ba4597, 32'hc140c678, 32'hc2a73f7a, 32'hc2c7207a, 32'h4043b114, 32'hbfdee607, 32'h4193d56d};
test_output[3765] = '{32'h4193d56d};
test_index[3765] = '{7};
test_input[30128:30135] = '{32'h4130026f, 32'h4211a86a, 32'hc2a15f7e, 32'hc246c9b8, 32'hc2bed2aa, 32'hc139ba48, 32'h4154bd8c, 32'hc23650da};
test_output[3766] = '{32'h4211a86a};
test_index[3766] = '{1};
test_input[30136:30143] = '{32'h416dc8cb, 32'hc2b7566e, 32'hc2906c5f, 32'h41b9184b, 32'h41fbc996, 32'h4175320b, 32'h42b19359, 32'h42b1cd61};
test_output[3767] = '{32'h42b1cd61};
test_index[3767] = '{7};
test_input[30144:30151] = '{32'hc2346efe, 32'h40e43382, 32'hc2b088b7, 32'h418b5222, 32'hc2888367, 32'hc2c2ec2b, 32'h426073bb, 32'h41a0de66};
test_output[3768] = '{32'h426073bb};
test_index[3768] = '{6};
test_input[30152:30159] = '{32'hc18aff49, 32'hc1ead2bb, 32'hc165718d, 32'hc253ca6f, 32'h426f5f72, 32'hc1b53ef6, 32'hc2b0da0a, 32'hc19104d2};
test_output[3769] = '{32'h426f5f72};
test_index[3769] = '{4};
test_input[30160:30167] = '{32'h42029db8, 32'h4296bf66, 32'hbfc3ce6f, 32'h4292bbf2, 32'h41ec2663, 32'h42c55ef0, 32'h41c913b0, 32'h416898f3};
test_output[3770] = '{32'h42c55ef0};
test_index[3770] = '{5};
test_input[30168:30175] = '{32'hc2c6378e, 32'hc0d63d42, 32'hc2b1b868, 32'h429ad441, 32'h425a9f14, 32'hc27d9def, 32'hc2922563, 32'h42a8a710};
test_output[3771] = '{32'h42a8a710};
test_index[3771] = '{7};
test_input[30176:30183] = '{32'h4262fc33, 32'hc2314165, 32'hc0b2a873, 32'h422337fb, 32'hc1cdffc9, 32'h42b09f56, 32'h413a6254, 32'hc1dad0ba};
test_output[3772] = '{32'h42b09f56};
test_index[3772] = '{5};
test_input[30184:30191] = '{32'h42ad67c1, 32'hc21bacec, 32'h429479c8, 32'hc298b06f, 32'h42c23341, 32'hc1e4a07b, 32'h4228e15a, 32'h4159d6a5};
test_output[3773] = '{32'h42c23341};
test_index[3773] = '{4};
test_input[30192:30199] = '{32'h42064cb6, 32'h426a15f1, 32'h42123bdc, 32'hc2c66c96, 32'h41e6b0b3, 32'hc24631b3, 32'hc2a01f85, 32'hc2c58794};
test_output[3774] = '{32'h426a15f1};
test_index[3774] = '{1};
test_input[30200:30207] = '{32'hc0f86d3e, 32'h42154756, 32'hc1edd54f, 32'hbf894a2e, 32'hc295965e, 32'hc2bfa645, 32'hc29ea374, 32'hc269ce32};
test_output[3775] = '{32'h42154756};
test_index[3775] = '{1};
test_input[30208:30215] = '{32'hc101b4a0, 32'h424f85c5, 32'hc15c51be, 32'hc22bb11c, 32'h429d4c5e, 32'hc293c9e3, 32'hc296dfc0, 32'hc258e1f7};
test_output[3776] = '{32'h429d4c5e};
test_index[3776] = '{4};
test_input[30216:30223] = '{32'hc02a60a8, 32'hc2c69e50, 32'h40f945a1, 32'h420eee13, 32'hc2185132, 32'h42564b1c, 32'h42462bd3, 32'h42949ab5};
test_output[3777] = '{32'h42949ab5};
test_index[3777] = '{7};
test_input[30224:30231] = '{32'hc2740d44, 32'h428c5e4f, 32'hc1bec90e, 32'hc1f5d927, 32'h41f2e227, 32'hc25e898d, 32'h423c54ad, 32'h4214674f};
test_output[3778] = '{32'h428c5e4f};
test_index[3778] = '{1};
test_input[30232:30239] = '{32'hc2677047, 32'hc2716185, 32'h42abcf01, 32'h41a6ea13, 32'hc25a2865, 32'hc2a31049, 32'h421df8a6, 32'hc2b4ea3d};
test_output[3779] = '{32'h42abcf01};
test_index[3779] = '{2};
test_input[30240:30247] = '{32'h42adffa2, 32'h420139ac, 32'hc2a346cf, 32'h42bd2913, 32'h429b8802, 32'h4095296d, 32'h42a1e163, 32'hbe355685};
test_output[3780] = '{32'h42bd2913};
test_index[3780] = '{3};
test_input[30248:30255] = '{32'h42937812, 32'hc16254cf, 32'hc26ea433, 32'h4273c01d, 32'hc1c6234c, 32'h41bc0906, 32'hc2856b25, 32'h428a2792};
test_output[3781] = '{32'h42937812};
test_index[3781] = '{0};
test_input[30256:30263] = '{32'hc281ef91, 32'h42a9fa18, 32'hc24a181c, 32'hc066555d, 32'hc1b9c12b, 32'hc2c6a48b, 32'h42756be8, 32'hc2955cdf};
test_output[3782] = '{32'h42a9fa18};
test_index[3782] = '{1};
test_input[30264:30271] = '{32'hc24cb90c, 32'h40c460a3, 32'h42ab9291, 32'h42315d74, 32'hc2005843, 32'h4004ea42, 32'hc2554057, 32'h42c73b7d};
test_output[3783] = '{32'h42c73b7d};
test_index[3783] = '{7};
test_input[30272:30279] = '{32'hc1bfa566, 32'hc2c18a4c, 32'h42c023db, 32'hc0cd2dec, 32'h42440c50, 32'hc2934159, 32'h421d41ae, 32'h3fc69182};
test_output[3784] = '{32'h42c023db};
test_index[3784] = '{2};
test_input[30280:30287] = '{32'h42c15e93, 32'h4218befe, 32'hc2382b79, 32'h42187f65, 32'hc26f8055, 32'h41c615bd, 32'h425ec56c, 32'h4215d502};
test_output[3785] = '{32'h42c15e93};
test_index[3785] = '{0};
test_input[30288:30295] = '{32'hc2498688, 32'hc2b0e33d, 32'hc295c442, 32'h416e7afa, 32'h4045af3e, 32'h42869205, 32'hc2838f32, 32'h4194041d};
test_output[3786] = '{32'h42869205};
test_index[3786] = '{5};
test_input[30296:30303] = '{32'hc1a109dc, 32'h421a9080, 32'hc1dc791e, 32'h42af4a26, 32'h429b1ead, 32'hc1879855, 32'hc287a8cb, 32'hc11a88ce};
test_output[3787] = '{32'h42af4a26};
test_index[3787] = '{3};
test_input[30304:30311] = '{32'h4253edca, 32'h426cd0d7, 32'h41ef48a1, 32'hc1c330df, 32'h4270b4a0, 32'h42241e21, 32'h413e22d7, 32'h429d8b21};
test_output[3788] = '{32'h429d8b21};
test_index[3788] = '{7};
test_input[30312:30319] = '{32'hc1d0510b, 32'hc28ac497, 32'h428fe0e6, 32'hc0d7daf6, 32'hc181592d, 32'hc274058a, 32'hc264bbd7, 32'hc0b0df21};
test_output[3789] = '{32'h428fe0e6};
test_index[3789] = '{2};
test_input[30320:30327] = '{32'h428a8fae, 32'h42342e19, 32'hc208b46f, 32'hc2a8b346, 32'h411e09c7, 32'hc2686076, 32'hc12a68db, 32'h41c73246};
test_output[3790] = '{32'h428a8fae};
test_index[3790] = '{0};
test_input[30328:30335] = '{32'h41b5d74c, 32'h429af221, 32'hc19eea91, 32'h418415f7, 32'hc1891298, 32'h429fe1bc, 32'hc2768c8c, 32'hc2b08795};
test_output[3791] = '{32'h429fe1bc};
test_index[3791] = '{5};
test_input[30336:30343] = '{32'hc2c6fb91, 32'hc294d553, 32'hc22782a6, 32'hc0cb391c, 32'h41e12d35, 32'hc0b84fe8, 32'h41b29ed8, 32'hc179c334};
test_output[3792] = '{32'h41e12d35};
test_index[3792] = '{4};
test_input[30344:30351] = '{32'hc2b7c201, 32'h429427f9, 32'h41804c85, 32'h4191d294, 32'h42a06c97, 32'h424394a9, 32'hc2a03093, 32'h42a7d3aa};
test_output[3793] = '{32'h42a7d3aa};
test_index[3793] = '{7};
test_input[30352:30359] = '{32'h42539fb1, 32'h40a8bfdd, 32'h41bf7d85, 32'h42087408, 32'h411769fe, 32'hc256263f, 32'h3e0e39d9, 32'hc1a2d592};
test_output[3794] = '{32'h42539fb1};
test_index[3794] = '{0};
test_input[30360:30367] = '{32'hc263f117, 32'h41e35565, 32'h424c6d85, 32'hc1bbcf01, 32'hc1e97e6d, 32'h429d94ab, 32'hc2862839, 32'h429d280c};
test_output[3795] = '{32'h429d94ab};
test_index[3795] = '{5};
test_input[30368:30375] = '{32'h422655bd, 32'h425b39e1, 32'hc2bb94cd, 32'hc28a54c3, 32'hc20508a7, 32'hc28f51b9, 32'h4264c983, 32'h4257e7c6};
test_output[3796] = '{32'h4264c983};
test_index[3796] = '{6};
test_input[30376:30383] = '{32'h42518b52, 32'hc21faa89, 32'hc2924702, 32'hc199453a, 32'hc2ae618f, 32'hc26fd44b, 32'hc1e24280, 32'hc2176d7f};
test_output[3797] = '{32'h42518b52};
test_index[3797] = '{0};
test_input[30384:30391] = '{32'h4212df18, 32'h423afc91, 32'h40b94ba4, 32'hc2c68d49, 32'h4293c882, 32'h410ba6d9, 32'hc2818569, 32'hc204e983};
test_output[3798] = '{32'h4293c882};
test_index[3798] = '{4};
test_input[30392:30399] = '{32'h41d05662, 32'h40202e7d, 32'hc2047c50, 32'hc27c759e, 32'h41cbb9ae, 32'h4194de56, 32'h428a6201, 32'h4223c958};
test_output[3799] = '{32'h428a6201};
test_index[3799] = '{6};
test_input[30400:30407] = '{32'h42997165, 32'hc28e2223, 32'h4283293b, 32'hc2a301ca, 32'hc22692d4, 32'hc0c497ec, 32'h42c31a15, 32'h4122234c};
test_output[3800] = '{32'h42c31a15};
test_index[3800] = '{6};
test_input[30408:30415] = '{32'h42b14646, 32'hc29f5846, 32'hbfbe3922, 32'h42a81038, 32'hc1f9a336, 32'hc29ed9a4, 32'h42b0e5a1, 32'h417a2ed2};
test_output[3801] = '{32'h42b14646};
test_index[3801] = '{0};
test_input[30416:30423] = '{32'h42a46379, 32'h41fe6ea2, 32'h419ff987, 32'hc189fab8, 32'h415e7227, 32'hc2934bb8, 32'hc1e280b1, 32'h4181966b};
test_output[3802] = '{32'h42a46379};
test_index[3802] = '{0};
test_input[30424:30431] = '{32'hc00c6f5f, 32'h42bf8810, 32'h425a267c, 32'h42863b25, 32'hc2197986, 32'h42881463, 32'hc2507d76, 32'h42325774};
test_output[3803] = '{32'h42bf8810};
test_index[3803] = '{1};
test_input[30432:30439] = '{32'h3fc26086, 32'hc0c0a34e, 32'hc28884af, 32'hc1365102, 32'hc2612542, 32'hc22de581, 32'h423eb2f9, 32'h42abc4f2};
test_output[3804] = '{32'h42abc4f2};
test_index[3804] = '{7};
test_input[30440:30447] = '{32'h40af262d, 32'hc08c52d9, 32'h42a0561c, 32'hc21b6618, 32'hc19641f1, 32'hc2a05aaf, 32'hc270c63d, 32'h42a09eeb};
test_output[3805] = '{32'h42a09eeb};
test_index[3805] = '{7};
test_input[30448:30455] = '{32'h418ed512, 32'hc25ba165, 32'hc1d49d8c, 32'h42aa1f46, 32'hc11c47b4, 32'h4223b60a, 32'h4235e2ed, 32'hc2735091};
test_output[3806] = '{32'h42aa1f46};
test_index[3806] = '{3};
test_input[30456:30463] = '{32'h41fac811, 32'h42729ef7, 32'hc2647104, 32'h413b1dfb, 32'hc1bdba39, 32'h4291a6f7, 32'hc0e3e19e, 32'h42bd792b};
test_output[3807] = '{32'h42bd792b};
test_index[3807] = '{7};
test_input[30464:30471] = '{32'hc23076a8, 32'hc1967e80, 32'hc21ac5f5, 32'hc24f7cf0, 32'h4297e66c, 32'hc23a7346, 32'h4019acf8, 32'hc2af3891};
test_output[3808] = '{32'h4297e66c};
test_index[3808] = '{4};
test_input[30472:30479] = '{32'h42144bc4, 32'h4109a57f, 32'hc28e6cf9, 32'hc2c013c8, 32'hc14956c0, 32'hc2a9db26, 32'hc251b230, 32'hc295d5bb};
test_output[3809] = '{32'h42144bc4};
test_index[3809] = '{0};
test_input[30480:30487] = '{32'h4084204d, 32'h4105905c, 32'h4242e615, 32'hc2300ee8, 32'h42b84af8, 32'hc2728c29, 32'h41ebd57c, 32'hc22160d9};
test_output[3810] = '{32'h42b84af8};
test_index[3810] = '{4};
test_input[30488:30495] = '{32'h41f79508, 32'h41ee0b58, 32'h3fd2c697, 32'h429b1937, 32'h41df2821, 32'hc23918fc, 32'hc235e857, 32'h421e3a60};
test_output[3811] = '{32'h429b1937};
test_index[3811] = '{3};
test_input[30496:30503] = '{32'h42bc7958, 32'h424cf596, 32'hc202f15d, 32'h423f837b, 32'h42212ded, 32'hc0cf81eb, 32'h418e3cb6, 32'hc2c486bf};
test_output[3812] = '{32'h42bc7958};
test_index[3812] = '{0};
test_input[30504:30511] = '{32'hc1bc583e, 32'hc2992733, 32'h4131caaf, 32'hc24679a7, 32'h421e2924, 32'hc2a21da1, 32'hc29deb54, 32'hc2b86da6};
test_output[3813] = '{32'h421e2924};
test_index[3813] = '{4};
test_input[30512:30519] = '{32'h42831425, 32'h423feb9f, 32'h42497593, 32'hc26de3c7, 32'hc2a9731f, 32'hc2c13043, 32'h4121ca63, 32'hc08eed97};
test_output[3814] = '{32'h42831425};
test_index[3814] = '{0};
test_input[30520:30527] = '{32'hc28a0bc1, 32'hc177e540, 32'h42c27adc, 32'hc2b7aee9, 32'hc2c21002, 32'h3f9d13d8, 32'hc295777b, 32'h42af869b};
test_output[3815] = '{32'h42c27adc};
test_index[3815] = '{2};
test_input[30528:30535] = '{32'h4109a3cd, 32'hc2ba6c75, 32'hc28c167c, 32'hc0b32e11, 32'h428f4382, 32'h42b35fa3, 32'hc285a51f, 32'hc1287ce3};
test_output[3816] = '{32'h42b35fa3};
test_index[3816] = '{5};
test_input[30536:30543] = '{32'h42a5da41, 32'h41a22ec6, 32'hc2241cf5, 32'hc1de9217, 32'h4285d2eb, 32'hc2c558ed, 32'hbe91d193, 32'hc1af4e13};
test_output[3817] = '{32'h42a5da41};
test_index[3817] = '{0};
test_input[30544:30551] = '{32'hc13c3cbb, 32'hc2bfe9e5, 32'hc1651682, 32'h4062328b, 32'h3e976e15, 32'h415a244b, 32'h41d63674, 32'h42476bba};
test_output[3818] = '{32'h42476bba};
test_index[3818] = '{7};
test_input[30552:30559] = '{32'hc24b82a5, 32'hc182d56d, 32'hc21d9bd3, 32'h42b65b89, 32'h41fd8df3, 32'hc1a9bc62, 32'hc1132e2e, 32'h42b3d857};
test_output[3819] = '{32'h42b65b89};
test_index[3819] = '{3};
test_input[30560:30567] = '{32'h4298b456, 32'hc23aab9d, 32'h42a75736, 32'h41126ea5, 32'hc2900b3f, 32'hc2864c84, 32'h424b101c, 32'hc1fad7b9};
test_output[3820] = '{32'h42a75736};
test_index[3820] = '{2};
test_input[30568:30575] = '{32'hc2bb53e7, 32'h42b47756, 32'h4169cc9d, 32'hc2bc2069, 32'hc1fd57e6, 32'hc29d29c6, 32'h42013abe, 32'h42a14f07};
test_output[3821] = '{32'h42b47756};
test_index[3821] = '{1};
test_input[30576:30583] = '{32'h4277b3df, 32'h426289bd, 32'hc2b370d2, 32'h422c8c75, 32'hc2515d2e, 32'h42a682fa, 32'hc29cd4e4, 32'hc2b4d630};
test_output[3822] = '{32'h42a682fa};
test_index[3822] = '{5};
test_input[30584:30591] = '{32'h429d5f38, 32'h3e8406c3, 32'hc2860a27, 32'hc0966401, 32'h426ab958, 32'hc10ef2ae, 32'h40ba885e, 32'h4085177e};
test_output[3823] = '{32'h429d5f38};
test_index[3823] = '{0};
test_input[30592:30599] = '{32'hc272e3aa, 32'h42b43705, 32'h42a9bc3e, 32'h410721da, 32'hc2b2fe33, 32'hc2a4f505, 32'hc294feaa, 32'h4287a87c};
test_output[3824] = '{32'h42b43705};
test_index[3824] = '{1};
test_input[30600:30607] = '{32'h41539d05, 32'hc291c701, 32'hc21521ef, 32'hc011a72a, 32'h42bfa104, 32'h41b2dbee, 32'hc1adcb55, 32'h4166ff07};
test_output[3825] = '{32'h42bfa104};
test_index[3825] = '{4};
test_input[30608:30615] = '{32'hc2a02872, 32'hc1e18fb9, 32'hc1897c0e, 32'hc184ea1f, 32'h4219ffc1, 32'hc2b94424, 32'h428cb5eb, 32'hc2a93f4f};
test_output[3826] = '{32'h428cb5eb};
test_index[3826] = '{6};
test_input[30616:30623] = '{32'h4265dc39, 32'hc16a92b2, 32'h42693219, 32'h427e8afb, 32'h40068e6f, 32'hc19a0c2e, 32'hc2b30516, 32'hc2ac5dc5};
test_output[3827] = '{32'h427e8afb};
test_index[3827] = '{3};
test_input[30624:30631] = '{32'hc270f4cb, 32'hc13cb42a, 32'h4279f11b, 32'hc1f7aeec, 32'hc2304d50, 32'hc127a9ed, 32'hc19ad351, 32'hc1f95bd7};
test_output[3828] = '{32'h4279f11b};
test_index[3828] = '{2};
test_input[30632:30639] = '{32'h4291a96c, 32'hc29c9d72, 32'h42915a22, 32'h4260d1ad, 32'hbecc830c, 32'hc2854bdb, 32'hc27d3661, 32'h42bbc270};
test_output[3829] = '{32'h42bbc270};
test_index[3829] = '{7};
test_input[30640:30647] = '{32'hc169c471, 32'h40a48d92, 32'hc2bba364, 32'hc23eff23, 32'h41c79b40, 32'h42af67ce, 32'hbedb608a, 32'h423ecafd};
test_output[3830] = '{32'h42af67ce};
test_index[3830] = '{5};
test_input[30648:30655] = '{32'h418b7e5f, 32'hc29ec839, 32'hc2977161, 32'hc263f89f, 32'h4242c05c, 32'h42204ae9, 32'hc06043a5, 32'h420cfb0d};
test_output[3831] = '{32'h4242c05c};
test_index[3831] = '{4};
test_input[30656:30663] = '{32'h42c40548, 32'hc1ed1c8c, 32'hc21b0711, 32'hc2016474, 32'h41fadb3c, 32'h41e1b9a9, 32'hc2349300, 32'hc22f3932};
test_output[3832] = '{32'h42c40548};
test_index[3832] = '{0};
test_input[30664:30671] = '{32'hc1cb1ef2, 32'h42905dba, 32'h42508aad, 32'hc1a276ec, 32'h418b7162, 32'hc24181c2, 32'h42811b46, 32'hc24f7cb8};
test_output[3833] = '{32'h42905dba};
test_index[3833] = '{1};
test_input[30672:30679] = '{32'h42c5a628, 32'h428ee9ff, 32'h41e4051d, 32'h4299280b, 32'h42348a31, 32'hc12e35d4, 32'hc2b4e122, 32'hc2acdae5};
test_output[3834] = '{32'h42c5a628};
test_index[3834] = '{0};
test_input[30680:30687] = '{32'h42ac64ea, 32'h4296ba8b, 32'hc2b7339e, 32'hc28c42af, 32'h42b58380, 32'hc2b610f1, 32'h42963d6c, 32'hc2b28f87};
test_output[3835] = '{32'h42b58380};
test_index[3835] = '{4};
test_input[30688:30695] = '{32'h429a2f5b, 32'hc1ee7114, 32'hc1eda205, 32'hc2bdca26, 32'h4275b960, 32'h419d3380, 32'hc20136e2, 32'hc28a13ca};
test_output[3836] = '{32'h429a2f5b};
test_index[3836] = '{0};
test_input[30696:30703] = '{32'hc1ec498f, 32'h426f69f6, 32'hc1846801, 32'h42b25aca, 32'hc20531df, 32'h4095fe02, 32'h41677427, 32'hc1eb3ab5};
test_output[3837] = '{32'h42b25aca};
test_index[3837] = '{3};
test_input[30704:30711] = '{32'h429670b0, 32'hc1e4aa74, 32'hc28f9582, 32'hc2a3ad89, 32'h41c7f734, 32'h41bc71de, 32'h429b0d39, 32'h4267a562};
test_output[3838] = '{32'h429b0d39};
test_index[3838] = '{6};
test_input[30712:30719] = '{32'h429b8d79, 32'h3eb71bdf, 32'h41c4bd36, 32'hc21a3009, 32'hc1ebc9a1, 32'hc26ddaee, 32'h41d5f246, 32'hc2c1cba8};
test_output[3839] = '{32'h429b8d79};
test_index[3839] = '{0};
test_input[30720:30727] = '{32'h42b60772, 32'hc28d71d0, 32'h4243a324, 32'h4125c5bc, 32'hc1935274, 32'hc2a658a3, 32'h40fc9584, 32'hc23231f1};
test_output[3840] = '{32'h42b60772};
test_index[3840] = '{0};
test_input[30728:30735] = '{32'hc2c54fbc, 32'hc2c0e591, 32'h41e0e4af, 32'h41631265, 32'hc1d1f7f1, 32'hc2a92c0e, 32'hc2552b8a, 32'h4263708a};
test_output[3841] = '{32'h4263708a};
test_index[3841] = '{7};
test_input[30736:30743] = '{32'hc2198347, 32'h424baa54, 32'hc275947c, 32'hc2b5f65e, 32'hc2520713, 32'h42c3a9b9, 32'hc26d3d90, 32'hc2429e33};
test_output[3842] = '{32'h42c3a9b9};
test_index[3842] = '{5};
test_input[30744:30751] = '{32'h42732726, 32'hc2704964, 32'h42060d79, 32'h42a39ca0, 32'hc25fae1b, 32'h40925f53, 32'hc138501a, 32'hc19d9e8f};
test_output[3843] = '{32'h42a39ca0};
test_index[3843] = '{3};
test_input[30752:30759] = '{32'h42812457, 32'hc2159c40, 32'h42832e4e, 32'hc2c19863, 32'h42b04d13, 32'h420f8c02, 32'h42bd97e9, 32'hc10fa2fb};
test_output[3844] = '{32'h42bd97e9};
test_index[3844] = '{6};
test_input[30760:30767] = '{32'hc22d1446, 32'h42c6e4d9, 32'hc1ad13b9, 32'hc2990598, 32'hc12b9a8c, 32'hc2a24711, 32'hc2499db0, 32'h429fc665};
test_output[3845] = '{32'h42c6e4d9};
test_index[3845] = '{1};
test_input[30768:30775] = '{32'hc26aee46, 32'h429543ec, 32'hc225fb72, 32'h41dd47a9, 32'h42b22029, 32'h4278731c, 32'hc24641c3, 32'hc28e0707};
test_output[3846] = '{32'h42b22029};
test_index[3846] = '{4};
test_input[30776:30783] = '{32'h423b447d, 32'h42489a43, 32'h428ce65f, 32'hc283ef68, 32'h42b4a336, 32'h426fbbbd, 32'hc09a3015, 32'h41ba4dce};
test_output[3847] = '{32'h42b4a336};
test_index[3847] = '{4};
test_input[30784:30791] = '{32'h42986731, 32'h41b1e709, 32'h42adea9b, 32'hc2888e84, 32'hc2993c52, 32'hc2bd57fe, 32'h42b391fa, 32'hc1c61376};
test_output[3848] = '{32'h42b391fa};
test_index[3848] = '{6};
test_input[30792:30799] = '{32'hc2b7da98, 32'h42c0a9d2, 32'hc06181c2, 32'hc2525271, 32'h4236a021, 32'hc2b4e67a, 32'hc2a3058e, 32'hc1ddae12};
test_output[3849] = '{32'h42c0a9d2};
test_index[3849] = '{1};
test_input[30800:30807] = '{32'h403f2bdb, 32'h421af336, 32'h4188055f, 32'h429e923f, 32'hc296814d, 32'hc2c4eedf, 32'h42925fbf, 32'hc29ddb28};
test_output[3850] = '{32'h429e923f};
test_index[3850] = '{3};
test_input[30808:30815] = '{32'h426e8f48, 32'h412f1721, 32'hc22a9d5f, 32'hc1b9a965, 32'h42be6eba, 32'hc0fa1e26, 32'h42518ff4, 32'hc2392ac5};
test_output[3851] = '{32'h42be6eba};
test_index[3851] = '{4};
test_input[30816:30823] = '{32'hc299a55a, 32'h42a7b303, 32'hc21041c3, 32'hc26167a5, 32'hc2c36454, 32'hc29a6e55, 32'h4208e39a, 32'hc148e6c6};
test_output[3852] = '{32'h42a7b303};
test_index[3852] = '{1};
test_input[30824:30831] = '{32'hc20d71d4, 32'h4278adfd, 32'h42ab6892, 32'h42b0ee64, 32'h4195285f, 32'hc1e07815, 32'hc228a299, 32'hc1c9d848};
test_output[3853] = '{32'h42b0ee64};
test_index[3853] = '{3};
test_input[30832:30839] = '{32'hc2902090, 32'hc231f589, 32'h42682071, 32'hc21f4d28, 32'h4295fdfc, 32'h42a0b73c, 32'h4214d665, 32'hc2842d10};
test_output[3854] = '{32'h42a0b73c};
test_index[3854] = '{5};
test_input[30840:30847] = '{32'hc125a16d, 32'hc2afc6aa, 32'hc2608413, 32'h422ca6fe, 32'h4188c411, 32'h40be4815, 32'h422c174b, 32'hc22051e2};
test_output[3855] = '{32'h422ca6fe};
test_index[3855] = '{3};
test_input[30848:30855] = '{32'h42af24fe, 32'hc1a88fec, 32'hc2ba0501, 32'hc2c3f29e, 32'hc1911314, 32'h42c33480, 32'hc1a8cfe8, 32'hc29360a2};
test_output[3856] = '{32'h42c33480};
test_index[3856] = '{5};
test_input[30856:30863] = '{32'h429992df, 32'h42bcd2a5, 32'h42885608, 32'h419eae45, 32'h4150d594, 32'hc2885a25, 32'h42b2e6fc, 32'h412116ad};
test_output[3857] = '{32'h42bcd2a5};
test_index[3857] = '{1};
test_input[30864:30871] = '{32'h42af6235, 32'h40b86203, 32'h40834dc7, 32'h41c8f550, 32'h429ec05f, 32'h4290fca4, 32'h41e19970, 32'h42bae1bb};
test_output[3858] = '{32'h42bae1bb};
test_index[3858] = '{7};
test_input[30872:30879] = '{32'h412d8d2a, 32'hc1e7e6d2, 32'h422f6d69, 32'h41ad4d9d, 32'hc1797fc0, 32'hc217649b, 32'hc1cabba4, 32'hc27a4db3};
test_output[3859] = '{32'h422f6d69};
test_index[3859] = '{2};
test_input[30880:30887] = '{32'hc20415f9, 32'h42523382, 32'hc2806b2a, 32'hbfbaa417, 32'hc276f13c, 32'h41ab36f6, 32'h40a71d8f, 32'h423d679a};
test_output[3860] = '{32'h42523382};
test_index[3860] = '{1};
test_input[30888:30895] = '{32'hc26a8d6b, 32'hc21debdc, 32'hc20ebe9b, 32'hc10d5414, 32'hc2265a34, 32'h418f569e, 32'hc2a92853, 32'hc1087ce1};
test_output[3861] = '{32'h418f569e};
test_index[3861] = '{5};
test_input[30896:30903] = '{32'hc29df3b1, 32'hc1e0357c, 32'hbfea574a, 32'h418d05d7, 32'h41acfa92, 32'h425884a8, 32'h3f7d3ab2, 32'hc1e99a93};
test_output[3862] = '{32'h425884a8};
test_index[3862] = '{5};
test_input[30904:30911] = '{32'h423e10fc, 32'h4275a8cf, 32'hc2bffd0c, 32'hc1a069ac, 32'h42b0c083, 32'hc218f06e, 32'h428353a1, 32'h421b5963};
test_output[3863] = '{32'h42b0c083};
test_index[3863] = '{4};
test_input[30912:30919] = '{32'h41d5870c, 32'hc1906340, 32'h429310a9, 32'hc2c08193, 32'hc2964357, 32'hc2a087ab, 32'h422221a5, 32'h426b788a};
test_output[3864] = '{32'h429310a9};
test_index[3864] = '{2};
test_input[30920:30927] = '{32'hc20a3960, 32'h41a929fd, 32'hc2abb6a8, 32'hc28ed024, 32'h424aae3d, 32'h427952fe, 32'h4235637c, 32'h42809b91};
test_output[3865] = '{32'h42809b91};
test_index[3865] = '{7};
test_input[30928:30935] = '{32'hc29c69d0, 32'h41a77960, 32'h42c22eba, 32'h42069277, 32'h42bac18a, 32'h40713ea4, 32'h41429167, 32'hc1e9b993};
test_output[3866] = '{32'h42c22eba};
test_index[3866] = '{2};
test_input[30936:30943] = '{32'h424154ca, 32'h424ce379, 32'hc277fcb9, 32'hc22bdc41, 32'h427e7cae, 32'hc268f710, 32'hc2983ed8, 32'hc27ef2fc};
test_output[3867] = '{32'h427e7cae};
test_index[3867] = '{4};
test_input[30944:30951] = '{32'hc2abbef6, 32'h42b1d542, 32'h42c3022c, 32'hc21dc155, 32'hc2025c94, 32'hc1fbbabb, 32'hc27b6846, 32'hc287e411};
test_output[3868] = '{32'h42c3022c};
test_index[3868] = '{2};
test_input[30952:30959] = '{32'hc0581833, 32'hc2807fd8, 32'hc228bfa7, 32'h426d55c4, 32'h420f29ac, 32'h425add35, 32'h41e9cb71, 32'hc2047067};
test_output[3869] = '{32'h426d55c4};
test_index[3869] = '{3};
test_input[30960:30967] = '{32'hc06f93ee, 32'hc282fef2, 32'h42a6b8c4, 32'h42b776fb, 32'hc22a2196, 32'h41ea84ee, 32'hc245228e, 32'hc294562e};
test_output[3870] = '{32'h42b776fb};
test_index[3870] = '{3};
test_input[30968:30975] = '{32'h4264d585, 32'hc20f24fc, 32'h42092478, 32'hc1481ee4, 32'hc1482db5, 32'h4231ed35, 32'h4139fd4e, 32'hc08c5d5e};
test_output[3871] = '{32'h4264d585};
test_index[3871] = '{0};
test_input[30976:30983] = '{32'h420c6c46, 32'h41320ff1, 32'hc22dbd5e, 32'hc2083e8d, 32'h423d0274, 32'hc18b7598, 32'hc2c3d583, 32'hc2aa1b16};
test_output[3872] = '{32'h423d0274};
test_index[3872] = '{4};
test_input[30984:30991] = '{32'h3fb0703c, 32'h4123784d, 32'hc20f7cab, 32'h411a9d38, 32'h42bcd598, 32'h425966d1, 32'h419936e7, 32'h42183871};
test_output[3873] = '{32'h42bcd598};
test_index[3873] = '{4};
test_input[30992:30999] = '{32'hc10350e4, 32'h42a7f493, 32'h41c053b9, 32'hbff937ff, 32'hc1b67c30, 32'h424bc5c0, 32'h42a338c9, 32'h4123ecde};
test_output[3874] = '{32'h42a7f493};
test_index[3874] = '{1};
test_input[31000:31007] = '{32'hc2aa5ebe, 32'h41cfaf94, 32'hc2452f31, 32'h409c112c, 32'hc151f0da, 32'hc253a191, 32'h42330fe6, 32'h426e7fcf};
test_output[3875] = '{32'h426e7fcf};
test_index[3875] = '{7};
test_input[31008:31015] = '{32'hc1fcb192, 32'h4236418c, 32'hc28c1375, 32'h42b22537, 32'hc1b5aa0d, 32'h4270e3eb, 32'hc1fd0c5f, 32'hc2afda9d};
test_output[3876] = '{32'h42b22537};
test_index[3876] = '{3};
test_input[31016:31023] = '{32'hc2bcf346, 32'h42a9b546, 32'h4240582b, 32'h42832a06, 32'hc29939d8, 32'hc1851727, 32'h42b08656, 32'h4285f65f};
test_output[3877] = '{32'h42b08656};
test_index[3877] = '{6};
test_input[31024:31031] = '{32'hc2b5bfde, 32'h4295e7ad, 32'hc2ae802c, 32'hc0c94508, 32'h4254a305, 32'hc293f0f8, 32'hc2abb0fe, 32'h42bb21cf};
test_output[3878] = '{32'h42bb21cf};
test_index[3878] = '{7};
test_input[31032:31039] = '{32'hc1ba24ff, 32'hc22b282f, 32'hc25a57e9, 32'h4199db6b, 32'h423f1e3c, 32'hc29836a8, 32'h41078078, 32'hc29555fe};
test_output[3879] = '{32'h423f1e3c};
test_index[3879] = '{4};
test_input[31040:31047] = '{32'h40ff85ac, 32'hc2c23eed, 32'h42942eb1, 32'h42c032a1, 32'hc2b50851, 32'h41b6315b, 32'hc257e107, 32'h411a611e};
test_output[3880] = '{32'h42c032a1};
test_index[3880] = '{3};
test_input[31048:31055] = '{32'hc29a532c, 32'h41c2bed8, 32'h42b1846d, 32'h42c79d82, 32'hc23447de, 32'hc1ced626, 32'h41bf2fc2, 32'hc28554e7};
test_output[3881] = '{32'h42c79d82};
test_index[3881] = '{3};
test_input[31056:31063] = '{32'hc243d757, 32'h425bec9a, 32'h41dcd4f3, 32'h42232ffe, 32'h429ff828, 32'hc26bc779, 32'h3f8ec901, 32'hc1ce81a9};
test_output[3882] = '{32'h429ff828};
test_index[3882] = '{4};
test_input[31064:31071] = '{32'hc022a2b8, 32'hc1aebc3a, 32'hc26745c2, 32'h42c11244, 32'hc2bb08f5, 32'hc104bcc5, 32'h42c75280, 32'h42910a6f};
test_output[3883] = '{32'h42c75280};
test_index[3883] = '{6};
test_input[31072:31079] = '{32'hc2a9e892, 32'hc2aa5238, 32'h42af4b29, 32'h4285dfc1, 32'h42231e22, 32'hc1e18153, 32'hc1bcf365, 32'h418055dc};
test_output[3884] = '{32'h42af4b29};
test_index[3884] = '{2};
test_input[31080:31087] = '{32'h42bfa37a, 32'hc289b08a, 32'hc2615dca, 32'hc28a1b14, 32'h42a40d49, 32'h42409d62, 32'hc29b8e0d, 32'h418d20f1};
test_output[3885] = '{32'h42bfa37a};
test_index[3885] = '{0};
test_input[31088:31095] = '{32'hc2a3bcf5, 32'h4129428b, 32'hc2b09f93, 32'h429cb548, 32'h400c29c7, 32'h42523f57, 32'hc2a8a735, 32'h42422350};
test_output[3886] = '{32'h429cb548};
test_index[3886] = '{3};
test_input[31096:31103] = '{32'hc2591b18, 32'hc129ce63, 32'h42aecff3, 32'h429208b3, 32'h4245aa6d, 32'hc1a568c6, 32'hc1d35684, 32'h42b27c9c};
test_output[3887] = '{32'h42b27c9c};
test_index[3887] = '{7};
test_input[31104:31111] = '{32'h40951f1a, 32'h42ab5e20, 32'h41130c13, 32'h4216ce53, 32'h4248b481, 32'h4148bd4c, 32'hc1a8f685, 32'hc28059a8};
test_output[3888] = '{32'h42ab5e20};
test_index[3888] = '{1};
test_input[31112:31119] = '{32'h42a8a8cd, 32'hc1e47bd0, 32'hc1cec4dc, 32'hc2a2d9b5, 32'h408cae63, 32'hc29cbe8b, 32'hc1d340a1, 32'h424df71e};
test_output[3889] = '{32'h42a8a8cd};
test_index[3889] = '{0};
test_input[31120:31127] = '{32'hc180645f, 32'h424fb0ff, 32'hc09d3eda, 32'hc157ec99, 32'h4126e03f, 32'hc2aea9a2, 32'h42b34713, 32'h427ccc53};
test_output[3890] = '{32'h42b34713};
test_index[3890] = '{6};
test_input[31128:31135] = '{32'h424469a8, 32'hc2771a58, 32'h3f694ad1, 32'hc246932f, 32'hc2247d9d, 32'hc2138f05, 32'h4289f9f3, 32'hc286b708};
test_output[3891] = '{32'h4289f9f3};
test_index[3891] = '{6};
test_input[31136:31143] = '{32'h400a0b92, 32'hc2a6fd6c, 32'hc2707cc1, 32'hc118eba9, 32'h42950bbc, 32'hc29f087e, 32'hc20e4a3e, 32'hbf6ed7e9};
test_output[3892] = '{32'h42950bbc};
test_index[3892] = '{4};
test_input[31144:31151] = '{32'hc28006e5, 32'h41902522, 32'hc2b5b179, 32'h42321eef, 32'hc2013048, 32'h3ed48956, 32'h42ad904e, 32'hc10d56d6};
test_output[3893] = '{32'h42ad904e};
test_index[3893] = '{6};
test_input[31152:31159] = '{32'hc21e77a7, 32'h42824df4, 32'hc24b76c4, 32'hc2c25ea0, 32'h4280fe4c, 32'hc2934186, 32'hc22700f8, 32'h42437125};
test_output[3894] = '{32'h42824df4};
test_index[3894] = '{1};
test_input[31160:31167] = '{32'h42794f10, 32'h42c2d7a5, 32'hc142ace0, 32'hc2b3e4c0, 32'hc18d3c6c, 32'hc28fc3ca, 32'hc228e917, 32'h414addba};
test_output[3895] = '{32'h42c2d7a5};
test_index[3895] = '{1};
test_input[31168:31175] = '{32'hc16828a9, 32'hc2c483a0, 32'h428dd3b5, 32'h421af3ad, 32'hc29dec51, 32'h42575f1c, 32'h4255567c, 32'hc20bf1a8};
test_output[3896] = '{32'h428dd3b5};
test_index[3896] = '{2};
test_input[31176:31183] = '{32'h42719ec7, 32'hc103972a, 32'hc2869cf2, 32'h4219b3c7, 32'h42b1f60f, 32'h425c1293, 32'h429e9119, 32'h42c46b86};
test_output[3897] = '{32'h42c46b86};
test_index[3897] = '{7};
test_input[31184:31191] = '{32'h42bb23b1, 32'h414f87fc, 32'hc110315f, 32'h427b8b7f, 32'h42acfa82, 32'hc21ac319, 32'hc2936306, 32'h41db829b};
test_output[3898] = '{32'h42bb23b1};
test_index[3898] = '{0};
test_input[31192:31199] = '{32'hc08bd9a2, 32'hc2b1d2d3, 32'h4208c11c, 32'hc2759bdc, 32'h422f26b1, 32'hc277e64b, 32'hc1e96387, 32'hc1ba9285};
test_output[3899] = '{32'h422f26b1};
test_index[3899] = '{4};
test_input[31200:31207] = '{32'h3f23c188, 32'h428269ff, 32'hc2856d90, 32'h4211a228, 32'hc2ad1b16, 32'hc2387506, 32'hc1a8a756, 32'hc2ada4cc};
test_output[3900] = '{32'h428269ff};
test_index[3900] = '{1};
test_input[31208:31215] = '{32'hc21e6f82, 32'hc2915159, 32'hc2497cab, 32'hc1c0b3e1, 32'hc1e961cb, 32'hc24984d3, 32'hc1b67490, 32'hc2954657};
test_output[3901] = '{32'hc1b67490};
test_index[3901] = '{6};
test_input[31216:31223] = '{32'hc142ea3c, 32'h411bfdd0, 32'hc2b98aee, 32'h4207f156, 32'h42759f45, 32'hc269cd29, 32'h403ffde1, 32'h429561ff};
test_output[3902] = '{32'h429561ff};
test_index[3902] = '{7};
test_input[31224:31231] = '{32'h4251f464, 32'hc270f7d0, 32'h40b1d9fc, 32'hc256eb2f, 32'hc29a4704, 32'hc1e337bf, 32'h4259134b, 32'hc29247ec};
test_output[3903] = '{32'h4259134b};
test_index[3903] = '{6};
test_input[31232:31239] = '{32'h42b08208, 32'h41b817e3, 32'hc28ac27a, 32'hc2522bc9, 32'hc2919bf0, 32'h4150987f, 32'hc235ff27, 32'h4262ef04};
test_output[3904] = '{32'h42b08208};
test_index[3904] = '{0};
test_input[31240:31247] = '{32'hc11cd33b, 32'hc2943338, 32'hc2939af6, 32'hc21113ca, 32'hc23bf52b, 32'h42a66a18, 32'hc20fc442, 32'hc1740653};
test_output[3905] = '{32'h42a66a18};
test_index[3905] = '{5};
test_input[31248:31255] = '{32'hc1af42df, 32'h4040df6c, 32'h427b6626, 32'hc29dfd71, 32'h4187aac5, 32'h40372e32, 32'h4070ac94, 32'hc2abcfdc};
test_output[3906] = '{32'h427b6626};
test_index[3906] = '{2};
test_input[31256:31263] = '{32'hc207a8c8, 32'hc2072884, 32'h4208a9a9, 32'hc2511567, 32'hc211652d, 32'hc2063ab5, 32'hc2be1445, 32'h42c3140f};
test_output[3907] = '{32'h42c3140f};
test_index[3907] = '{7};
test_input[31264:31271] = '{32'h418b3689, 32'hc21d0817, 32'h423f556b, 32'hc0f59f7c, 32'h40a89eb2, 32'hc221980d, 32'hc0dd2151, 32'hc1af6353};
test_output[3908] = '{32'h423f556b};
test_index[3908] = '{2};
test_input[31272:31279] = '{32'hc17ea49f, 32'hc1dea7fc, 32'hc194285b, 32'h40d1d98b, 32'h42b092d6, 32'hc2bccba7, 32'hc2b69eb7, 32'h426562bb};
test_output[3909] = '{32'h42b092d6};
test_index[3909] = '{4};
test_input[31280:31287] = '{32'hc18c6d96, 32'h422a0c27, 32'h40a27a01, 32'h4124edf8, 32'hc29e30fa, 32'h421d3ba8, 32'hc2269d02, 32'hc21f1746};
test_output[3910] = '{32'h422a0c27};
test_index[3910] = '{1};
test_input[31288:31295] = '{32'h4226d555, 32'hc239216d, 32'hc2a0aae8, 32'hc222f332, 32'h42bd2c38, 32'hc2c142d0, 32'hc2c2384f, 32'h42b9c245};
test_output[3911] = '{32'h42bd2c38};
test_index[3911] = '{4};
test_input[31296:31303] = '{32'h41bb6eb8, 32'hc158d5a2, 32'hc2a7a5d3, 32'hc2041792, 32'h42889987, 32'hc03f2667, 32'h4274db54, 32'hc2a6ba9e};
test_output[3912] = '{32'h42889987};
test_index[3912] = '{4};
test_input[31304:31311] = '{32'h419cc14f, 32'h424b9596, 32'h428e97b9, 32'h42be6ce0, 32'h42b31ff8, 32'hc1c07d4e, 32'h42b6f995, 32'hc2730d86};
test_output[3913] = '{32'h42be6ce0};
test_index[3913] = '{3};
test_input[31312:31319] = '{32'hc18adcf3, 32'hc2b90024, 32'h42b91747, 32'hc24105b0, 32'h423059b2, 32'hc2561f1e, 32'h425bcda3, 32'h42013fb6};
test_output[3914] = '{32'h42b91747};
test_index[3914] = '{2};
test_input[31320:31327] = '{32'h4296cb88, 32'h42ae76e9, 32'h404162a8, 32'hc1d502c3, 32'h4136352f, 32'hc20d2949, 32'h426a5964, 32'h413caf4b};
test_output[3915] = '{32'h42ae76e9};
test_index[3915] = '{1};
test_input[31328:31335] = '{32'h428219e9, 32'h403d0154, 32'hc1ea5f32, 32'h4209ad03, 32'hc2af7eb8, 32'hc2a81ee0, 32'hc2c1b199, 32'h4223b23b};
test_output[3916] = '{32'h428219e9};
test_index[3916] = '{0};
test_input[31336:31343] = '{32'hc2b8f977, 32'h424a4925, 32'hc2084873, 32'h41d24cc3, 32'hc19a1aba, 32'hc23e270f, 32'h419b15e2, 32'hc1afdf14};
test_output[3917] = '{32'h424a4925};
test_index[3917] = '{1};
test_input[31344:31351] = '{32'h42be9bd3, 32'hc2bc8e58, 32'h4282196f, 32'hc2b21c8f, 32'hc0a53327, 32'hc28834ac, 32'hc29abf80, 32'hc157d35f};
test_output[3918] = '{32'h42be9bd3};
test_index[3918] = '{0};
test_input[31352:31359] = '{32'hc246fdc2, 32'h41fb3516, 32'hc2522ed0, 32'hc28285b9, 32'hc1cf5326, 32'h4252c2e2, 32'hc243186c, 32'h40dd3f03};
test_output[3919] = '{32'h4252c2e2};
test_index[3919] = '{5};
test_input[31360:31367] = '{32'h40b5d249, 32'hc23b7c3b, 32'hc19ef9dd, 32'hc2c1372f, 32'h41b9326e, 32'h426e72b7, 32'hc1b8c818, 32'hc1c465cf};
test_output[3920] = '{32'h426e72b7};
test_index[3920] = '{5};
test_input[31368:31375] = '{32'hc01b2eee, 32'h40e978d6, 32'h4289a328, 32'h42820f2e, 32'h41738938, 32'hc03f2a3f, 32'hc1c2dfb0, 32'hc2b6775f};
test_output[3921] = '{32'h4289a328};
test_index[3921] = '{2};
test_input[31376:31383] = '{32'hbeab6fd8, 32'h4105e989, 32'hc2a0e9f5, 32'h41e2da76, 32'hc29feada, 32'hc0967b21, 32'hc1e92ccd, 32'hc21fd00d};
test_output[3922] = '{32'h41e2da76};
test_index[3922] = '{3};
test_input[31384:31391] = '{32'h4259cd1b, 32'h425318ec, 32'h4271d458, 32'hc03d5b31, 32'h428fac5e, 32'hc1072600, 32'h42aff33f, 32'h42c0b40d};
test_output[3923] = '{32'h42c0b40d};
test_index[3923] = '{7};
test_input[31392:31399] = '{32'h429b0aba, 32'hc263f091, 32'h40dc5eb3, 32'hc28bcf75, 32'hbd83de26, 32'h42b36969, 32'h425f80d3, 32'h41984826};
test_output[3924] = '{32'h42b36969};
test_index[3924] = '{5};
test_input[31400:31407] = '{32'h41dde59a, 32'h42a5bb31, 32'h418a9e88, 32'hc29a794f, 32'hc2909941, 32'hc2afc5b1, 32'hc2c698d2, 32'hc29e2270};
test_output[3925] = '{32'h42a5bb31};
test_index[3925] = '{1};
test_input[31408:31415] = '{32'hc1f7a8f7, 32'hc29d7d38, 32'h42a08269, 32'h4282f136, 32'hc280b179, 32'h42bfc878, 32'h42051157, 32'hc26f5db0};
test_output[3926] = '{32'h42bfc878};
test_index[3926] = '{5};
test_input[31416:31423] = '{32'h4225e181, 32'h42436619, 32'hbf3465e8, 32'h424fe119, 32'h417b97c9, 32'hc26f340c, 32'hc2c47665, 32'h4085112d};
test_output[3927] = '{32'h424fe119};
test_index[3927] = '{3};
test_input[31424:31431] = '{32'hc2544fce, 32'h425ddd1e, 32'hc29f8d58, 32'h41ed5187, 32'hc2a731b9, 32'h424df95c, 32'hc22bf8e7, 32'h4240a3cf};
test_output[3928] = '{32'h425ddd1e};
test_index[3928] = '{1};
test_input[31432:31439] = '{32'h42ba09ed, 32'h42a1ea03, 32'h42896066, 32'hc0768021, 32'h4211aa47, 32'h3fe8e97f, 32'hc23e9dc7, 32'hc2af2b2f};
test_output[3929] = '{32'h42ba09ed};
test_index[3929] = '{0};
test_input[31440:31447] = '{32'hc230cf85, 32'h418aa7c5, 32'hc27485cc, 32'h41812322, 32'hc219f531, 32'hc243f3f8, 32'hc2a1eaf2, 32'h42905588};
test_output[3930] = '{32'h42905588};
test_index[3930] = '{7};
test_input[31448:31455] = '{32'h42a098b9, 32'hc1b52d76, 32'h4263c778, 32'hc1b75121, 32'h42615fc5, 32'hc2a5e0be, 32'h42660736, 32'hc17a2c9c};
test_output[3931] = '{32'h42a098b9};
test_index[3931] = '{0};
test_input[31456:31463] = '{32'h42ae4a5a, 32'hc1b647f7, 32'h42325999, 32'h42839e5d, 32'hc2ac8e3b, 32'hc2b54f44, 32'h42afb452, 32'hc1de6d6c};
test_output[3932] = '{32'h42afb452};
test_index[3932] = '{6};
test_input[31464:31471] = '{32'h42899809, 32'hc1f381f8, 32'h4295a26a, 32'h417fa3aa, 32'hc2b42540, 32'h42b29f11, 32'h425d6410, 32'hc0745ab8};
test_output[3933] = '{32'h42b29f11};
test_index[3933] = '{5};
test_input[31472:31479] = '{32'h41a2332e, 32'h422f00b3, 32'hc2afdea9, 32'hc24d893b, 32'hc2911389, 32'h42049fa1, 32'h41e759db, 32'h418522e5};
test_output[3934] = '{32'h422f00b3};
test_index[3934] = '{1};
test_input[31480:31487] = '{32'h41dcdb8c, 32'h4213627b, 32'h422bedaa, 32'hc0bae630, 32'h41d7c01b, 32'hc1ebb168, 32'hc190013c, 32'hbfbcd770};
test_output[3935] = '{32'h422bedaa};
test_index[3935] = '{2};
test_input[31488:31495] = '{32'h40cd15fa, 32'hc28e3af0, 32'h40fe2b58, 32'hc23d2548, 32'hc26b5c10, 32'h41e41638, 32'h4057bc10, 32'hc28a27e6};
test_output[3936] = '{32'h41e41638};
test_index[3936] = '{5};
test_input[31496:31503] = '{32'h41970d4e, 32'h40face84, 32'hc0b0b8fd, 32'hc221086f, 32'h42bf9ba7, 32'hc2336f63, 32'h426aaa4e, 32'h423d56ec};
test_output[3937] = '{32'h42bf9ba7};
test_index[3937] = '{4};
test_input[31504:31511] = '{32'h421ad207, 32'h41826efa, 32'h4253d76c, 32'h4297da93, 32'hbfb422c1, 32'hc2356a34, 32'h42965ea6, 32'hc20f4a41};
test_output[3938] = '{32'h4297da93};
test_index[3938] = '{3};
test_input[31512:31519] = '{32'hc2609202, 32'h429849cf, 32'h428cb008, 32'h417878b3, 32'hc2b09b48, 32'hc1c93792, 32'h4291bd50, 32'hc2a623b9};
test_output[3939] = '{32'h429849cf};
test_index[3939] = '{1};
test_input[31520:31527] = '{32'h42b1564e, 32'hc28a6db7, 32'h426ef617, 32'hc23f6246, 32'h423b48bc, 32'h4299a3e0, 32'hc2387f9a, 32'h4229cd76};
test_output[3940] = '{32'h42b1564e};
test_index[3940] = '{0};
test_input[31528:31535] = '{32'h42836951, 32'hc2b735f5, 32'h425a522f, 32'h41b56522, 32'h429e4a32, 32'h42aa5981, 32'hc291f046, 32'h412151e5};
test_output[3941] = '{32'h42aa5981};
test_index[3941] = '{5};
test_input[31536:31543] = '{32'hc02b6c7f, 32'hc1407b5c, 32'h42c4e32a, 32'hc2a7a31b, 32'h42b06fbd, 32'h425628e1, 32'hc24c1b9b, 32'hc0db0381};
test_output[3942] = '{32'h42c4e32a};
test_index[3942] = '{2};
test_input[31544:31551] = '{32'h42001749, 32'h4274b8c2, 32'hc2991d9c, 32'hc0dd79aa, 32'hc2a14ec3, 32'hc19226de, 32'hc29820e3, 32'h42b9f900};
test_output[3943] = '{32'h42b9f900};
test_index[3943] = '{7};
test_input[31552:31559] = '{32'h41ead598, 32'h40f1690e, 32'hc11532d5, 32'hc1707f04, 32'h4286f84b, 32'h42b0180e, 32'hc2bbfbe3, 32'hc2ac0ec6};
test_output[3944] = '{32'h42b0180e};
test_index[3944] = '{5};
test_input[31560:31567] = '{32'h424cbc4a, 32'hc2a61384, 32'h420516e7, 32'hc2341023, 32'h4299615e, 32'h3caf5957, 32'hc28a5d1c, 32'hc1d5f2fa};
test_output[3945] = '{32'h4299615e};
test_index[3945] = '{4};
test_input[31568:31575] = '{32'h42468ed1, 32'h41d845b0, 32'h4203d21d, 32'h42a2d0d8, 32'hc293c0c3, 32'h42881c8d, 32'hc23e22ac, 32'h425420f4};
test_output[3946] = '{32'h42a2d0d8};
test_index[3946] = '{3};
test_input[31576:31583] = '{32'hc200b2f4, 32'h425e4f5f, 32'h42262b2c, 32'hc0b5e72a, 32'hc1949b08, 32'h428e9afe, 32'hc1e1412e, 32'h42bd4b84};
test_output[3947] = '{32'h42bd4b84};
test_index[3947] = '{7};
test_input[31584:31591] = '{32'hc20c8538, 32'h425ec2ef, 32'h424e18e6, 32'hc206b660, 32'hc27c8f59, 32'h42be0e71, 32'h411f3f0e, 32'hc18b927d};
test_output[3948] = '{32'h42be0e71};
test_index[3948] = '{5};
test_input[31592:31599] = '{32'h421b0a23, 32'h42b692b2, 32'h425ffb3e, 32'h42bdcb4a, 32'h41c98352, 32'h42b42050, 32'hc1978a56, 32'hc24014ef};
test_output[3949] = '{32'h42bdcb4a};
test_index[3949] = '{3};
test_input[31600:31607] = '{32'hc24bceed, 32'hc24c1cad, 32'h4291ddb4, 32'h429d0684, 32'h41992776, 32'hc1bc5214, 32'h42966c4c, 32'h42303cec};
test_output[3950] = '{32'h429d0684};
test_index[3950] = '{3};
test_input[31608:31615] = '{32'h421deaaf, 32'h42a5629e, 32'h41c62542, 32'h4290a782, 32'h4295f1ca, 32'hc277ac4a, 32'hc2491b39, 32'h4262b339};
test_output[3951] = '{32'h42a5629e};
test_index[3951] = '{1};
test_input[31616:31623] = '{32'hc137f7cf, 32'hc20b4088, 32'h42c18f3c, 32'hc1f3dc69, 32'hc294d33e, 32'hc2016911, 32'h420c9c76, 32'h424177e1};
test_output[3952] = '{32'h42c18f3c};
test_index[3952] = '{2};
test_input[31624:31631] = '{32'hc2811fb6, 32'hc266db5f, 32'hc29a5a0b, 32'h42a4b44a, 32'hc2bfd540, 32'h4192919a, 32'h419d2101, 32'hc1d681e4};
test_output[3953] = '{32'h42a4b44a};
test_index[3953] = '{3};
test_input[31632:31639] = '{32'hc23bdbca, 32'h427e2e03, 32'hc2b70c93, 32'hc2232254, 32'hc2b363b6, 32'h424eda3c, 32'h42995931, 32'h41bed8a9};
test_output[3954] = '{32'h42995931};
test_index[3954] = '{6};
test_input[31640:31647] = '{32'hc203ba0b, 32'h40b0a3eb, 32'hc2740f89, 32'hc234ea95, 32'hc18b1dd9, 32'h428848be, 32'hc2a3d8d8, 32'hc10bee36};
test_output[3955] = '{32'h428848be};
test_index[3955] = '{5};
test_input[31648:31655] = '{32'h42191ded, 32'hc2b232c3, 32'h4281b302, 32'h417cfbe6, 32'h41921896, 32'hc2116bb9, 32'hc20ffe58, 32'h42924679};
test_output[3956] = '{32'h42924679};
test_index[3956] = '{7};
test_input[31656:31663] = '{32'h3f7f2b5f, 32'hc2c19755, 32'h42068de8, 32'hc1f7cdec, 32'h41e1de4b, 32'h41d16b01, 32'hc2a85f08, 32'hc216d7ca};
test_output[3957] = '{32'h42068de8};
test_index[3957] = '{2};
test_input[31664:31671] = '{32'hc0b16e66, 32'h4226e7b5, 32'hc2707178, 32'hc213a02e, 32'hc2aa44f6, 32'h42455a2e, 32'h41593728, 32'hc220f235};
test_output[3958] = '{32'h42455a2e};
test_index[3958] = '{5};
test_input[31672:31679] = '{32'hc27e5ec7, 32'h42a24771, 32'h4259291d, 32'hc2aec93f, 32'hc25b3bec, 32'hc1eadb35, 32'h42a11cf7, 32'hc2a401bb};
test_output[3959] = '{32'h42a24771};
test_index[3959] = '{1};
test_input[31680:31687] = '{32'hc2935525, 32'h42485cab, 32'hc0516104, 32'hc116d3dd, 32'hc298938e, 32'hc2c4c7c9, 32'hc286df95, 32'hc2b41e45};
test_output[3960] = '{32'h42485cab};
test_index[3960] = '{1};
test_input[31688:31695] = '{32'h412292a2, 32'h40f922ae, 32'hc28b6f05, 32'hc11828e5, 32'hc2156c33, 32'h42517045, 32'hc0eec8ac, 32'hc0e90384};
test_output[3961] = '{32'h42517045};
test_index[3961] = '{5};
test_input[31696:31703] = '{32'h417b7371, 32'h42c33773, 32'h3e9d0068, 32'h42a3862b, 32'hc21d617b, 32'hc28b89c0, 32'hc21b21cd, 32'h4272a96d};
test_output[3962] = '{32'h42c33773};
test_index[3962] = '{1};
test_input[31704:31711] = '{32'hc2be4614, 32'hc2b6be73, 32'hc25151ca, 32'hc2885e57, 32'h426e1c60, 32'h41239f6e, 32'h4201bed4, 32'hc056fbec};
test_output[3963] = '{32'h426e1c60};
test_index[3963] = '{4};
test_input[31712:31719] = '{32'hc1a6afd8, 32'h4267294a, 32'h42b5ca94, 32'hc28f12c4, 32'hc17e1301, 32'hc0c879e0, 32'hc080ce89, 32'h423b3119};
test_output[3964] = '{32'h42b5ca94};
test_index[3964] = '{2};
test_input[31720:31727] = '{32'hc290a1b9, 32'h42ad63fd, 32'hc2bcf099, 32'hc29dd5b7, 32'h42c34abe, 32'h42b6cfaf, 32'h42b5d3c5, 32'h425606c0};
test_output[3965] = '{32'h42c34abe};
test_index[3965] = '{4};
test_input[31728:31735] = '{32'h41811b1a, 32'h42c7f5bd, 32'h42902499, 32'h4292a2c5, 32'hc1a04bfa, 32'h42329b87, 32'h41d513bf, 32'h424a4a69};
test_output[3966] = '{32'h42c7f5bd};
test_index[3966] = '{1};
test_input[31736:31743] = '{32'h3f86f60c, 32'h42bb8d32, 32'h4214a8d6, 32'h425e862b, 32'h40f1b6ad, 32'hc291ea12, 32'hc2ba6171, 32'hc15bf414};
test_output[3967] = '{32'h42bb8d32};
test_index[3967] = '{1};
test_input[31744:31751] = '{32'h420ac839, 32'hc24a5d9b, 32'h41e19437, 32'hc2b0e91f, 32'hc298f359, 32'hc27c8ba9, 32'hc28ebd3d, 32'hc2c31b08};
test_output[3968] = '{32'h420ac839};
test_index[3968] = '{0};
test_input[31752:31759] = '{32'hc2bac08d, 32'h42380b9b, 32'h423674ab, 32'h40fa7e57, 32'h40e5cde3, 32'hc1ea5251, 32'h401ede14, 32'hc2a9828a};
test_output[3969] = '{32'h42380b9b};
test_index[3969] = '{1};
test_input[31760:31767] = '{32'hc2b78e4a, 32'h40eff15e, 32'hc28fef6f, 32'h42bf2b2c, 32'hc28146fc, 32'h4251aaab, 32'h42b2ba1b, 32'h41458983};
test_output[3970] = '{32'h42bf2b2c};
test_index[3970] = '{3};
test_input[31768:31775] = '{32'hc2575b0a, 32'hc14f5087, 32'hc247d21c, 32'h42bafb9e, 32'h42925e13, 32'hc1b040f9, 32'h423f0aef, 32'h42852133};
test_output[3971] = '{32'h42bafb9e};
test_index[3971] = '{3};
test_input[31776:31783] = '{32'hc189cc3c, 32'h42afd073, 32'h42958750, 32'h42bc5baf, 32'h42a81c88, 32'hc0db95a1, 32'hc27610b8, 32'h414ec225};
test_output[3972] = '{32'h42bc5baf};
test_index[3972] = '{3};
test_input[31784:31791] = '{32'hc2033088, 32'h41ac8175, 32'h42628e44, 32'h42b850e8, 32'hc21a52a0, 32'h414cc90a, 32'hc2921148, 32'hc2755054};
test_output[3973] = '{32'h42b850e8};
test_index[3973] = '{3};
test_input[31792:31799] = '{32'h41effaaf, 32'h4197a548, 32'h4164549b, 32'hc27567d6, 32'h405e6336, 32'h42880ed4, 32'hc29242c5, 32'h422257ca};
test_output[3974] = '{32'h42880ed4};
test_index[3974] = '{5};
test_input[31800:31807] = '{32'h3fcbb7ef, 32'hc285c63e, 32'h40db067c, 32'hc18b46c4, 32'hc25433fe, 32'h41fbcb03, 32'hc27124bd, 32'h428e41a3};
test_output[3975] = '{32'h428e41a3};
test_index[3975] = '{7};
test_input[31808:31815] = '{32'h42507a34, 32'hc2b24741, 32'h4292bcd4, 32'hc2803c25, 32'h42a71b8c, 32'h42b4f3c5, 32'h41e9804a, 32'hc27b2c0d};
test_output[3976] = '{32'h42b4f3c5};
test_index[3976] = '{5};
test_input[31816:31823] = '{32'h41e65a59, 32'hc2c26a9f, 32'hc2bec53f, 32'h42334b49, 32'h429a5ee1, 32'hc1d96886, 32'hc28820b7, 32'hc21fb8a6};
test_output[3977] = '{32'h429a5ee1};
test_index[3977] = '{4};
test_input[31824:31831] = '{32'hc1a0b89f, 32'h42bf3d8b, 32'h42c35330, 32'hc2be179c, 32'h429b0547, 32'h41bbc51c, 32'h42c22e9d, 32'h42a4af23};
test_output[3978] = '{32'h42c35330};
test_index[3978] = '{2};
test_input[31832:31839] = '{32'hc2a87b0a, 32'hc258596a, 32'hc10c2316, 32'h420fa765, 32'hc267cd99, 32'h42a8cae3, 32'h4299d7aa, 32'hc2169d91};
test_output[3979] = '{32'h42a8cae3};
test_index[3979] = '{5};
test_input[31840:31847] = '{32'hc2864e4c, 32'h41358edc, 32'hc14badd2, 32'hc17d2c24, 32'h413de6e8, 32'h41293983, 32'h425c5f57, 32'hc1b38953};
test_output[3980] = '{32'h425c5f57};
test_index[3980] = '{6};
test_input[31848:31855] = '{32'h41c85e92, 32'hc19686c1, 32'hc1aacedc, 32'h41a88baa, 32'h41221fb6, 32'hc1b7598f, 32'hc24badfd, 32'h42bb55cb};
test_output[3981] = '{32'h42bb55cb};
test_index[3981] = '{7};
test_input[31856:31863] = '{32'h427b5ebe, 32'h429fcc92, 32'h423984fa, 32'h4116b59b, 32'h425e8239, 32'h4154bb10, 32'h422ce17d, 32'hc29e6444};
test_output[3982] = '{32'h429fcc92};
test_index[3982] = '{1};
test_input[31864:31871] = '{32'hc24a65b8, 32'hc248a35a, 32'h42bb90f8, 32'hc2a34e0f, 32'h42a72c46, 32'hc1d0cabf, 32'h42595231, 32'h427d119a};
test_output[3983] = '{32'h42bb90f8};
test_index[3983] = '{2};
test_input[31872:31879] = '{32'h4284f44d, 32'h4229265a, 32'h428ccec7, 32'h41d79769, 32'h425a8883, 32'h4231413b, 32'h423dea4e, 32'h42275af0};
test_output[3984] = '{32'h428ccec7};
test_index[3984] = '{2};
test_input[31880:31887] = '{32'h42178057, 32'h41086248, 32'h42602de2, 32'h4224ffff, 32'h429811d7, 32'hc192ca0f, 32'hc2b4fb34, 32'hc2b77042};
test_output[3985] = '{32'h429811d7};
test_index[3985] = '{4};
test_input[31888:31895] = '{32'hc2811bf1, 32'hc151785c, 32'h429e5468, 32'hc101f52a, 32'hc228707e, 32'h427966b3, 32'hc2c4533f, 32'hc2b5f92a};
test_output[3986] = '{32'h429e5468};
test_index[3986] = '{2};
test_input[31896:31903] = '{32'hc19dd6d6, 32'h42b20d6e, 32'h42376871, 32'h4278fb05, 32'h42b4cc35, 32'hc20472dc, 32'h4184faff, 32'hc2bd4ec0};
test_output[3987] = '{32'h42b4cc35};
test_index[3987] = '{4};
test_input[31904:31911] = '{32'h41e389d2, 32'h421dc654, 32'h4136bf32, 32'h4235b081, 32'hc230ea0d, 32'h42201402, 32'h412ff287, 32'hc29448d0};
test_output[3988] = '{32'h4235b081};
test_index[3988] = '{3};
test_input[31912:31919] = '{32'hc29e3ebc, 32'h4276326f, 32'h42c24242, 32'h42358309, 32'h4231b888, 32'h4276aedd, 32'hc2a06441, 32'h41b2889f};
test_output[3989] = '{32'h42c24242};
test_index[3989] = '{2};
test_input[31920:31927] = '{32'hc28b544f, 32'h4253f75d, 32'h424ad378, 32'h428e75e4, 32'hc2b816fc, 32'h415e38b9, 32'hc27bed4e, 32'hc2c2f68e};
test_output[3990] = '{32'h428e75e4};
test_index[3990] = '{3};
test_input[31928:31935] = '{32'hc27aa440, 32'hc05c818c, 32'hc1890f99, 32'hc0ff6590, 32'h41b7fe94, 32'h42baec07, 32'h3fed6cff, 32'hc25a58ed};
test_output[3991] = '{32'h42baec07};
test_index[3991] = '{5};
test_input[31936:31943] = '{32'h4257a72f, 32'h428a34c8, 32'hc1d7f2ea, 32'hc1a09a4e, 32'hc1f932d2, 32'hc2c55589, 32'hc1607ec7, 32'h4149f5a4};
test_output[3992] = '{32'h428a34c8};
test_index[3992] = '{1};
test_input[31944:31951] = '{32'h4281f2ce, 32'h42b90c30, 32'h42c49255, 32'h42b1cc33, 32'hc2bc9c67, 32'h3f45aa6e, 32'hc2a339d1, 32'h428a36e5};
test_output[3993] = '{32'h42c49255};
test_index[3993] = '{2};
test_input[31952:31959] = '{32'hc2996c16, 32'hc286b6de, 32'h42afd7ca, 32'hc23caa0a, 32'h426bbe78, 32'h42a10f8a, 32'h4285c3fa, 32'hc232f680};
test_output[3994] = '{32'h42afd7ca};
test_index[3994] = '{2};
test_input[31960:31967] = '{32'hc16b712c, 32'h41ceb781, 32'h41477a0f, 32'h42554b10, 32'hc2c19c12, 32'h40bbd76b, 32'hc244bbc1, 32'h41fcbd47};
test_output[3995] = '{32'h42554b10};
test_index[3995] = '{3};
test_input[31968:31975] = '{32'hc272fd5e, 32'hc03d511d, 32'hc135ee98, 32'hc2b4bf1d, 32'h4231e1d3, 32'hc2b9b053, 32'h42012a49, 32'hc296384f};
test_output[3996] = '{32'h4231e1d3};
test_index[3996] = '{4};
test_input[31976:31983] = '{32'h41b062c4, 32'h42bf36dc, 32'hc226b742, 32'hc2113278, 32'h42bd4cba, 32'h41b0d7b9, 32'h40de043d, 32'h42057bfd};
test_output[3997] = '{32'h42bf36dc};
test_index[3997] = '{1};
test_input[31984:31991] = '{32'h418f7a1a, 32'h42947f8f, 32'h428ac607, 32'h42b3a997, 32'hc1f1b23b, 32'h429879b3, 32'hc2226775, 32'hc25a7527};
test_output[3998] = '{32'h42b3a997};
test_index[3998] = '{3};
test_input[31992:31999] = '{32'hc221983e, 32'h42c55e7a, 32'hc1e179d6, 32'hc2b2c2a0, 32'h41cdb6b6, 32'h411944bb, 32'hc28b2d7e, 32'hc227ae94};
test_output[3999] = '{32'h42c55e7a};
test_index[3999] = '{1};
test_input[32000:32007] = '{32'hc288cc36, 32'hc276e426, 32'hc2aa44dd, 32'hc2a8df16, 32'h4255a9a3, 32'hc1e1fee6, 32'h41640a31, 32'hc199e2e5};
test_output[4000] = '{32'h4255a9a3};
test_index[4000] = '{4};
test_input[32008:32015] = '{32'h429c5983, 32'h42716679, 32'h42a573ce, 32'h42c3af12, 32'h41d79394, 32'hc230f5b4, 32'h42aaa17c, 32'h421645c9};
test_output[4001] = '{32'h42c3af12};
test_index[4001] = '{3};
test_input[32016:32023] = '{32'hc0a81238, 32'h4251826a, 32'hc0ecf2b6, 32'h429e8d47, 32'hc2bd921b, 32'hc11433e1, 32'hc2ad1f5e, 32'hc14e52b1};
test_output[4002] = '{32'h429e8d47};
test_index[4002] = '{3};
test_input[32024:32031] = '{32'hc0ecd67e, 32'h4274c5b2, 32'hc2b3a03f, 32'h4216bc15, 32'h424a4335, 32'h41cba5ae, 32'hc2acfec4, 32'hc03e3262};
test_output[4003] = '{32'h4274c5b2};
test_index[4003] = '{1};
test_input[32032:32039] = '{32'hc1a1fee0, 32'hc2b66f49, 32'hbfba1dbe, 32'h423b0e05, 32'hc2b95d82, 32'hc10a995e, 32'hc1dbc548, 32'h423e3c1b};
test_output[4004] = '{32'h423e3c1b};
test_index[4004] = '{7};
test_input[32040:32047] = '{32'hc218f649, 32'h42037b4d, 32'hc212bc6e, 32'hc222e221, 32'hc253e299, 32'h42a88d6d, 32'hc1f969cf, 32'hc2bd1648};
test_output[4005] = '{32'h42a88d6d};
test_index[4005] = '{5};
test_input[32048:32055] = '{32'hc1629002, 32'h413888db, 32'hc1a6d9d5, 32'hc29c5854, 32'hc2416031, 32'hc2148a1b, 32'hc25e6a19, 32'h42626737};
test_output[4006] = '{32'h42626737};
test_index[4006] = '{7};
test_input[32056:32063] = '{32'hc21cd3bb, 32'hc299743d, 32'hbe1110ec, 32'h4197a8a2, 32'hc173bce2, 32'hc2917a7d, 32'hc2bdd027, 32'h429ee79a};
test_output[4007] = '{32'h429ee79a};
test_index[4007] = '{7};
test_input[32064:32071] = '{32'h424f553b, 32'h42b7351d, 32'hc2b5cdad, 32'h428300ea, 32'h42931493, 32'h42b933bd, 32'h425e6132, 32'h41cdf605};
test_output[4008] = '{32'h42b933bd};
test_index[4008] = '{5};
test_input[32072:32079] = '{32'hbfcd9199, 32'hc2bfbbc2, 32'h42153c1c, 32'h40c6599e, 32'hc2835436, 32'hc21598c3, 32'h4282c610, 32'h429f528f};
test_output[4009] = '{32'h429f528f};
test_index[4009] = '{7};
test_input[32080:32087] = '{32'hc1d1ec63, 32'hc27191dd, 32'hc1019f67, 32'hc24113bf, 32'hc1b4f46a, 32'h427b1afe, 32'h42ba17f5, 32'hc2a4b726};
test_output[4010] = '{32'h42ba17f5};
test_index[4010] = '{6};
test_input[32088:32095] = '{32'h42395fb8, 32'hc229c020, 32'hc28dd046, 32'h4105c463, 32'h41e399c1, 32'h42c098df, 32'h42187de1, 32'h42955d71};
test_output[4011] = '{32'h42c098df};
test_index[4011] = '{5};
test_input[32096:32103] = '{32'hc29c5991, 32'hc2bf8afc, 32'h42550931, 32'hc178e0dc, 32'hc2558d4a, 32'hc1147204, 32'hc20420e4, 32'hc21fa6f1};
test_output[4012] = '{32'h42550931};
test_index[4012] = '{2};
test_input[32104:32111] = '{32'h42009588, 32'h425c079f, 32'h427d7e87, 32'hc2acc1b3, 32'h41e3f582, 32'hc273a23c, 32'hc287498b, 32'hc1c6ce2b};
test_output[4013] = '{32'h427d7e87};
test_index[4013] = '{2};
test_input[32112:32119] = '{32'h42186084, 32'hc15793be, 32'hc207764d, 32'hc1fe265a, 32'hc2baa4ae, 32'hc2648778, 32'h42a46f8c, 32'hc2c54281};
test_output[4014] = '{32'h42a46f8c};
test_index[4014] = '{6};
test_input[32120:32127] = '{32'h4286bb9b, 32'h4242e4aa, 32'h419b861a, 32'hc26e9b15, 32'h42b78ca7, 32'h42c3817c, 32'h42a39756, 32'hc2c36dd3};
test_output[4015] = '{32'h42c3817c};
test_index[4015] = '{5};
test_input[32128:32135] = '{32'h42270c47, 32'h42a55a61, 32'hc2199c44, 32'h42b0243b, 32'hc29d665c, 32'h413efdf0, 32'h417e7383, 32'h424cfa3a};
test_output[4016] = '{32'h42b0243b};
test_index[4016] = '{3};
test_input[32136:32143] = '{32'h4233865b, 32'h42c33cda, 32'hc2c7d2dc, 32'hc16496af, 32'hc0130db8, 32'h41eb5805, 32'h42679000, 32'h41ab4bab};
test_output[4017] = '{32'h42c33cda};
test_index[4017] = '{1};
test_input[32144:32151] = '{32'hc10254c4, 32'hc14efd57, 32'hc23fc20d, 32'h42a6c226, 32'h41b13f1d, 32'h41e81f1e, 32'hc28dbbf6, 32'hc29486af};
test_output[4018] = '{32'h42a6c226};
test_index[4018] = '{3};
test_input[32152:32159] = '{32'h420c93f0, 32'h4241875e, 32'hc2663e0b, 32'hc2166b39, 32'hc2c1d321, 32'h421b64a9, 32'hc2a1544e, 32'h42043049};
test_output[4019] = '{32'h4241875e};
test_index[4019] = '{1};
test_input[32160:32167] = '{32'h42c4f0c2, 32'h421d116c, 32'h414c2802, 32'hc28f31ea, 32'hc2396ea0, 32'hc2931347, 32'h426ffda2, 32'h422c6b0b};
test_output[4020] = '{32'h42c4f0c2};
test_index[4020] = '{0};
test_input[32168:32175] = '{32'h42a969f0, 32'hc2bcaf2a, 32'hc2208a2b, 32'h421f8973, 32'h41ce2bf8, 32'h4211128f, 32'hc1a3a287, 32'h42a861b9};
test_output[4021] = '{32'h42a969f0};
test_index[4021] = '{0};
test_input[32176:32183] = '{32'h42bf74a5, 32'hc292f037, 32'h428a7bd7, 32'h3f83b148, 32'hc2c4074e, 32'hc210e262, 32'h418aa790, 32'hc21c6a84};
test_output[4022] = '{32'h42bf74a5};
test_index[4022] = '{0};
test_input[32184:32191] = '{32'h428f66db, 32'h42745ed3, 32'hc2b5981b, 32'h4280fdba, 32'hc2540efb, 32'hc2468311, 32'h42bd01b1, 32'h42c5f9a2};
test_output[4023] = '{32'h42c5f9a2};
test_index[4023] = '{7};
test_input[32192:32199] = '{32'hbfb9a5ec, 32'hc1d9c338, 32'h427ab0b4, 32'hc1b07343, 32'h42abd87a, 32'h42539240, 32'h41c414dd, 32'h42a0e109};
test_output[4024] = '{32'h42abd87a};
test_index[4024] = '{4};
test_input[32200:32207] = '{32'h425724d9, 32'hc142023d, 32'h416b7c9c, 32'h41847d41, 32'hc1134878, 32'hc24c8fdf, 32'h42915658, 32'h416b4361};
test_output[4025] = '{32'h42915658};
test_index[4025] = '{6};
test_input[32208:32215] = '{32'h416841ba, 32'hc15912a1, 32'hc267193f, 32'hc06ed322, 32'hc1f23b28, 32'h42a95272, 32'h422be06c, 32'hc201c318};
test_output[4026] = '{32'h42a95272};
test_index[4026] = '{5};
test_input[32216:32223] = '{32'hc057147b, 32'h4286bbfa, 32'h41d78079, 32'h423b6e76, 32'hc1d85152, 32'hc21182f1, 32'h4259b884, 32'h4138c87a};
test_output[4027] = '{32'h4286bbfa};
test_index[4027] = '{1};
test_input[32224:32231] = '{32'h41f97acd, 32'h42a4c5a6, 32'h4298a8df, 32'hc1df8111, 32'hbffd3c9b, 32'hc24dd469, 32'hc17b78f1, 32'h429db605};
test_output[4028] = '{32'h42a4c5a6};
test_index[4028] = '{1};
test_input[32232:32239] = '{32'h424a4150, 32'hc2b4453e, 32'h418e6c9f, 32'hc260d284, 32'h4211032e, 32'hc21732ef, 32'h42b81134, 32'hc2b1f255};
test_output[4029] = '{32'h42b81134};
test_index[4029] = '{6};
test_input[32240:32247] = '{32'h42851fce, 32'h427300ae, 32'h42a12024, 32'hc2a2fd31, 32'h429cdef6, 32'hc1996f84, 32'hc212c107, 32'h428ecd09};
test_output[4030] = '{32'h42a12024};
test_index[4030] = '{2};
test_input[32248:32255] = '{32'h427cf8b1, 32'h4264f141, 32'hc2246e81, 32'hc294c960, 32'hc181ee1e, 32'h4215a90c, 32'h41a914cb, 32'h428c1dc7};
test_output[4031] = '{32'h428c1dc7};
test_index[4031] = '{7};
test_input[32256:32263] = '{32'hc12fc0b4, 32'h41891650, 32'hc2581c85, 32'h41007754, 32'hc28a31ed, 32'h4245298c, 32'h42bd72fd, 32'hc1e060c8};
test_output[4032] = '{32'h42bd72fd};
test_index[4032] = '{6};
test_input[32264:32271] = '{32'hc29235fa, 32'hc0ab0f0e, 32'hc27de41e, 32'h423973fd, 32'hc1222ced, 32'h42c04b09, 32'h42b7d603, 32'h42804321};
test_output[4033] = '{32'h42c04b09};
test_index[4033] = '{5};
test_input[32272:32279] = '{32'h42a7bb40, 32'hc2be9fbd, 32'h4252669b, 32'h4004a3dd, 32'h4246e2f7, 32'h3ea1418a, 32'h41ca8672, 32'hc23291b2};
test_output[4034] = '{32'h42a7bb40};
test_index[4034] = '{0};
test_input[32280:32287] = '{32'h427b1d63, 32'h423cbd3f, 32'hc18db52d, 32'h418932c0, 32'hc25056b1, 32'h424013d7, 32'hc29bfce4, 32'h400b688e};
test_output[4035] = '{32'h427b1d63};
test_index[4035] = '{0};
test_input[32288:32295] = '{32'h41d1d2d7, 32'h428370e0, 32'h4211ba5e, 32'h42417425, 32'hc1870d51, 32'h41d376fd, 32'hc2ac8bee, 32'h416c3226};
test_output[4036] = '{32'h428370e0};
test_index[4036] = '{1};
test_input[32296:32303] = '{32'hc16519ea, 32'hc1eb36fd, 32'hc227c98f, 32'hc16219bd, 32'hc2917e87, 32'hc2248287, 32'h4253544b, 32'h41cc86d8};
test_output[4037] = '{32'h4253544b};
test_index[4037] = '{6};
test_input[32304:32311] = '{32'hc1bb7087, 32'h42c5fc16, 32'h41b5c01e, 32'hc22ce6da, 32'hc21850f2, 32'hc2a11115, 32'h418fbfac, 32'hc22a65c4};
test_output[4038] = '{32'h42c5fc16};
test_index[4038] = '{1};
test_input[32312:32319] = '{32'hc2b05907, 32'hc2376606, 32'h42c0914b, 32'h420a845a, 32'hc289bdaf, 32'h4238f61b, 32'hc268ddd1, 32'h417163eb};
test_output[4039] = '{32'h42c0914b};
test_index[4039] = '{2};
test_input[32320:32327] = '{32'h42a3f7e4, 32'hc20dab85, 32'h41dcbf8f, 32'h42272d2c, 32'hc142618e, 32'hc24a1125, 32'hc1d0065e, 32'h42990efd};
test_output[4040] = '{32'h42a3f7e4};
test_index[4040] = '{0};
test_input[32328:32335] = '{32'hc291bcdc, 32'h42582988, 32'h42ab7726, 32'hc1fd6709, 32'h426d5815, 32'hc2bb2ff4, 32'hc2b10e81, 32'h42a09979};
test_output[4041] = '{32'h42ab7726};
test_index[4041] = '{2};
test_input[32336:32343] = '{32'h42bb6074, 32'h428ee1cf, 32'h4202cffe, 32'hc288828a, 32'hc1430f10, 32'hc284f0d3, 32'h42bc08cc, 32'hc258083f};
test_output[4042] = '{32'h42bc08cc};
test_index[4042] = '{6};
test_input[32344:32351] = '{32'h42b25216, 32'hc289aa14, 32'hc18d9a1e, 32'hc2a33559, 32'h424c3566, 32'h42a22c58, 32'h42bdf8e6, 32'hc1d092b4};
test_output[4043] = '{32'h42bdf8e6};
test_index[4043] = '{6};
test_input[32352:32359] = '{32'hc21edc8d, 32'hc239c393, 32'hc2b5d7e1, 32'hc1c8e993, 32'h417b7e2f, 32'hbfad3b70, 32'h4207312a, 32'hc2bf4df2};
test_output[4044] = '{32'h4207312a};
test_index[4044] = '{6};
test_input[32360:32367] = '{32'h42a94a66, 32'hc1925c70, 32'h42775403, 32'h41223104, 32'hc0bd595c, 32'h4286ef60, 32'hc208d975, 32'hc2accb7d};
test_output[4045] = '{32'h42a94a66};
test_index[4045] = '{0};
test_input[32368:32375] = '{32'h428c78c7, 32'hc20dfdd1, 32'hc0eb6b32, 32'h42a01481, 32'hc245bf27, 32'h42928c36, 32'h424d1cbf, 32'h415093b3};
test_output[4046] = '{32'h42a01481};
test_index[4046] = '{3};
test_input[32376:32383] = '{32'hc274b96f, 32'h42599124, 32'hc2a39134, 32'h4118b230, 32'h424ab628, 32'hc2a31655, 32'h4295668f, 32'hc2642e91};
test_output[4047] = '{32'h4295668f};
test_index[4047] = '{6};
test_input[32384:32391] = '{32'h4199fb4a, 32'hc04143c7, 32'hc280bca2, 32'hc2106d5f, 32'hc27da860, 32'hc1836d0c, 32'hc12fbd3b, 32'h4223edae};
test_output[4048] = '{32'h4223edae};
test_index[4048] = '{7};
test_input[32392:32399] = '{32'h41a23d88, 32'hc2c236bf, 32'h419940cf, 32'hc237a422, 32'hc2b4e14e, 32'hc227a50d, 32'h410c319d, 32'h42c6bfee};
test_output[4049] = '{32'h42c6bfee};
test_index[4049] = '{7};
test_input[32400:32407] = '{32'hc09d9ac1, 32'h41ed690b, 32'h4290e8f8, 32'h415c6040, 32'hc2301d8d, 32'h423d4513, 32'hc2beb123, 32'h42791b0f};
test_output[4050] = '{32'h4290e8f8};
test_index[4050] = '{2};
test_input[32408:32415] = '{32'h41fb4224, 32'hc2876f21, 32'hc1232666, 32'hc25ea790, 32'hc2a78acf, 32'h41238507, 32'hc268e6ae, 32'hc1f16fc1};
test_output[4051] = '{32'h41fb4224};
test_index[4051] = '{0};
test_input[32416:32423] = '{32'hc2ba0ef3, 32'h420cdb6e, 32'hc19048f4, 32'hc0ed8be0, 32'hc11484dc, 32'h429d446e, 32'hbfc604b1, 32'h42900dd7};
test_output[4052] = '{32'h429d446e};
test_index[4052] = '{5};
test_input[32424:32431] = '{32'hc2120a78, 32'h42bb32bb, 32'hc2923c32, 32'hc2186ec2, 32'hc260bb52, 32'hc23bd33f, 32'hc06a9262, 32'h42a88e7e};
test_output[4053] = '{32'h42bb32bb};
test_index[4053] = '{1};
test_input[32432:32439] = '{32'hc2a3bb45, 32'hc1cd612e, 32'hc19266b6, 32'h3ca1ef5c, 32'hc26924d1, 32'hc2bab4f1, 32'hc16a0237, 32'hc19ddb9f};
test_output[4054] = '{32'h3ca1ef5c};
test_index[4054] = '{3};
test_input[32440:32447] = '{32'hc29f3daf, 32'h42aebefd, 32'h42815593, 32'h423f8fcf, 32'h421a8f04, 32'h42c65aab, 32'h42713bae, 32'h41e1e258};
test_output[4055] = '{32'h42c65aab};
test_index[4055] = '{5};
test_input[32448:32455] = '{32'h423e461e, 32'hc1df6316, 32'hc2bd57e6, 32'hc28be621, 32'h42bf55bb, 32'hc2c2e400, 32'h420a5c94, 32'hc28ee9b1};
test_output[4056] = '{32'h42bf55bb};
test_index[4056] = '{4};
test_input[32456:32463] = '{32'hbffe5f3a, 32'h42194e1c, 32'h41c14384, 32'h42ba2230, 32'h421bdca2, 32'h42987c55, 32'h4255999c, 32'hc239ed8f};
test_output[4057] = '{32'h42ba2230};
test_index[4057] = '{3};
test_input[32464:32471] = '{32'h4283af35, 32'h42b3dda0, 32'hc2c0333f, 32'hc2a21585, 32'h42877c39, 32'hc1f11f84, 32'h4214d4d9, 32'h427f0e50};
test_output[4058] = '{32'h42b3dda0};
test_index[4058] = '{1};
test_input[32472:32479] = '{32'h4281302b, 32'h40888a68, 32'hc236f542, 32'hc2449c90, 32'h424b2fe3, 32'hc288027f, 32'h423b4358, 32'h401f5a83};
test_output[4059] = '{32'h4281302b};
test_index[4059] = '{0};
test_input[32480:32487] = '{32'h423730c8, 32'h41808363, 32'h417f81bb, 32'hc24496a5, 32'h40ad3107, 32'hc2a866b5, 32'hc21a347c, 32'h400ce723};
test_output[4060] = '{32'h423730c8};
test_index[4060] = '{0};
test_input[32488:32495] = '{32'hc1d3762b, 32'h42b27fe9, 32'hc1ae2862, 32'h40b748a1, 32'h420980ec, 32'h4246d86c, 32'hc23dc95f, 32'h41e44d9b};
test_output[4061] = '{32'h42b27fe9};
test_index[4061] = '{1};
test_input[32496:32503] = '{32'hc263ddff, 32'hc1d57125, 32'hc2b29608, 32'hc2b897f1, 32'hc1eee869, 32'hc2bf857e, 32'hc0b4c82c, 32'h42c46482};
test_output[4062] = '{32'h42c46482};
test_index[4062] = '{7};
test_input[32504:32511] = '{32'hc2b44d41, 32'h4297d40e, 32'hc2464215, 32'hc2a5fa66, 32'h42b6179a, 32'h4188fd4b, 32'h409b578f, 32'h42423e7e};
test_output[4063] = '{32'h42b6179a};
test_index[4063] = '{4};
test_input[32512:32519] = '{32'hc2aa5699, 32'h428089d3, 32'h42498d07, 32'hc22b560c, 32'h427dd998, 32'h428ca798, 32'h4232aa17, 32'hc2850d58};
test_output[4064] = '{32'h428ca798};
test_index[4064] = '{5};
test_input[32520:32527] = '{32'h42715876, 32'hc207ed99, 32'hc257040d, 32'h41e68e56, 32'h42371b0a, 32'h422a407e, 32'hc212942f, 32'h42115b94};
test_output[4065] = '{32'h42715876};
test_index[4065] = '{0};
test_input[32528:32535] = '{32'hc0c80189, 32'hbfcca695, 32'hc29a2aca, 32'h42b99a82, 32'h420a0dff, 32'h40f9b370, 32'h42ae549c, 32'hc2a10b46};
test_output[4066] = '{32'h42b99a82};
test_index[4066] = '{3};
test_input[32536:32543] = '{32'h42944a5d, 32'h42315188, 32'h42855cd3, 32'h4194c08d, 32'h423d0523, 32'hc221d046, 32'h40f8c121, 32'h422e45c1};
test_output[4067] = '{32'h42944a5d};
test_index[4067] = '{0};
test_input[32544:32551] = '{32'hc28544ce, 32'h416d28cc, 32'hc13b1313, 32'h40482112, 32'h3f002e98, 32'h42c251e2, 32'h42656f36, 32'h421cc6dd};
test_output[4068] = '{32'h42c251e2};
test_index[4068] = '{5};
test_input[32552:32559] = '{32'h424e29a8, 32'hc232360a, 32'hc2aa6a64, 32'hc28b55bd, 32'hc21af4f0, 32'h427d2059, 32'h4292d805, 32'h4290b1bb};
test_output[4069] = '{32'h4292d805};
test_index[4069] = '{6};
test_input[32560:32567] = '{32'hc105e7b7, 32'hc2b6b706, 32'h4254d994, 32'h4278b4b5, 32'hc2aa7621, 32'hc28b88f0, 32'hc26d24c4, 32'hc21f8c36};
test_output[4070] = '{32'h4278b4b5};
test_index[4070] = '{3};
test_input[32568:32575] = '{32'hc2b3b47d, 32'h42399ec4, 32'hc1a1305d, 32'hc19a89f0, 32'hc2b52109, 32'h428eae5a, 32'hc26226b8, 32'hc2840233};
test_output[4071] = '{32'h428eae5a};
test_index[4071] = '{5};
test_input[32576:32583] = '{32'h428106cc, 32'hc25e3de0, 32'h42109d34, 32'hc1961408, 32'hc168b788, 32'h42156db9, 32'h41c57b02, 32'h4210787f};
test_output[4072] = '{32'h428106cc};
test_index[4072] = '{0};
test_input[32584:32591] = '{32'h41ee4902, 32'h40a8a6eb, 32'hc2acaafa, 32'h429b5392, 32'h426a5ff8, 32'hc2c778d6, 32'hc2804a8e, 32'hc298fe03};
test_output[4073] = '{32'h429b5392};
test_index[4073] = '{3};
test_input[32592:32599] = '{32'h4289a556, 32'hc1f41eb7, 32'hc1a53eeb, 32'h4148569d, 32'hc22da4b6, 32'h42afd3b5, 32'hc2205cc6, 32'hc285b4b0};
test_output[4074] = '{32'h42afd3b5};
test_index[4074] = '{5};
test_input[32600:32607] = '{32'hc2c695f5, 32'hc2692f33, 32'hc235f073, 32'hc13b6609, 32'h41edf6cf, 32'h428c3c28, 32'hc2a4161f, 32'hc24ea0ff};
test_output[4075] = '{32'h428c3c28};
test_index[4075] = '{5};
test_input[32608:32615] = '{32'h40987f28, 32'hc23ce1ae, 32'h4279d9eb, 32'hc2a80a12, 32'h42bad0f3, 32'h4271a2f1, 32'h42416809, 32'hc29c166a};
test_output[4076] = '{32'h42bad0f3};
test_index[4076] = '{4};
test_input[32616:32623] = '{32'h4209306a, 32'h429825b6, 32'hc23d1916, 32'h4254cd5c, 32'h422b5cea, 32'hc20121b9, 32'h424e8ad9, 32'h422c34d3};
test_output[4077] = '{32'h429825b6};
test_index[4077] = '{1};
test_input[32624:32631] = '{32'h40ee1d2a, 32'hc0ffc84c, 32'h42bc077e, 32'h4259f808, 32'h42aed769, 32'hc240d374, 32'h429971f9, 32'h420b3af2};
test_output[4078] = '{32'h42bc077e};
test_index[4078] = '{2};
test_input[32632:32639] = '{32'h4236a555, 32'hc1ac945a, 32'hbe22c23c, 32'hc22022c2, 32'h42078111, 32'hc1d1b04f, 32'hc2562ba4, 32'h426c7884};
test_output[4079] = '{32'h426c7884};
test_index[4079] = '{7};
test_input[32640:32647] = '{32'h42c090da, 32'hc291d50e, 32'hc188acdd, 32'hc116b173, 32'h41ed3470, 32'h4288d640, 32'h42c5feb9, 32'h4281b2c7};
test_output[4080] = '{32'h42c5feb9};
test_index[4080] = '{6};
test_input[32648:32655] = '{32'hc1145b35, 32'h41afdf28, 32'hc2b218bd, 32'hc2948b2b, 32'h421bac9f, 32'hc10d997e, 32'h426f8de6, 32'hc0b85e6f};
test_output[4081] = '{32'h426f8de6};
test_index[4081] = '{6};
test_input[32656:32663] = '{32'hc14d04d6, 32'hc29ee14d, 32'hc27b44c3, 32'h3e20171d, 32'hc1fce9f0, 32'h42223c12, 32'h4212811c, 32'h42b0981a};
test_output[4082] = '{32'h42b0981a};
test_index[4082] = '{7};
test_input[32664:32671] = '{32'hc0490437, 32'hc1b278cb, 32'h424d6d99, 32'h42b17da0, 32'h42724e13, 32'hc2447257, 32'hbf0be458, 32'hc2652753};
test_output[4083] = '{32'h42b17da0};
test_index[4083] = '{3};
test_input[32672:32679] = '{32'h4181e8df, 32'hc21e965a, 32'h427de8a0, 32'h429e8175, 32'hc2c2955f, 32'h42a5bf95, 32'hc29adcbc, 32'hc2a847a1};
test_output[4084] = '{32'h42a5bf95};
test_index[4084] = '{5};
test_input[32680:32687] = '{32'hc20e1b59, 32'hc297d505, 32'hc2a43f8d, 32'hc295a14b, 32'h42b56d49, 32'h42237fad, 32'h41ca22b5, 32'h424ba459};
test_output[4085] = '{32'h42b56d49};
test_index[4085] = '{4};
test_input[32688:32695] = '{32'hc2255d85, 32'h422f721b, 32'h42796fba, 32'hc227421a, 32'hc296a6d2, 32'h4275568a, 32'hc191a4a3, 32'h4271a162};
test_output[4086] = '{32'h42796fba};
test_index[4086] = '{2};
test_input[32696:32703] = '{32'h41929361, 32'hc162bcec, 32'hc2be44fa, 32'hc29a4933, 32'hc2bfdc58, 32'h42a01b38, 32'h4100157c, 32'h40ff304c};
test_output[4087] = '{32'h42a01b38};
test_index[4087] = '{5};
test_input[32704:32711] = '{32'h41dc0971, 32'hc1c8352a, 32'h42626be3, 32'h42a35134, 32'h421f0353, 32'hc19a88b9, 32'hc2adebde, 32'hc29c6bcc};
test_output[4088] = '{32'h42a35134};
test_index[4088] = '{3};
test_input[32712:32719] = '{32'hc2a38a98, 32'hc18299f6, 32'h41ac030b, 32'hc2b0ff02, 32'hc21bedd6, 32'hc1b66b07, 32'h4213ceea, 32'hc239a7dd};
test_output[4089] = '{32'h4213ceea};
test_index[4089] = '{6};
test_input[32720:32727] = '{32'h420f64fc, 32'hc1cddb43, 32'hc283f0c6, 32'hc288bc06, 32'h40fb4320, 32'hc272797a, 32'hc28091b5, 32'h41ef6ce6};
test_output[4090] = '{32'h420f64fc};
test_index[4090] = '{0};
test_input[32728:32735] = '{32'h42331ae7, 32'hc0e8263b, 32'h4154f4b9, 32'hc27775a5, 32'h41467c3c, 32'hc16bd91a, 32'h42bb3596, 32'hc28ea6d1};
test_output[4091] = '{32'h42bb3596};
test_index[4091] = '{6};
test_input[32736:32743] = '{32'h410ebf12, 32'hc1e32e76, 32'h423d802e, 32'hc2418b8a, 32'hc1149f85, 32'h4289d2f0, 32'hc2196b98, 32'hc20fdad7};
test_output[4092] = '{32'h4289d2f0};
test_index[4092] = '{5};
test_input[32744:32751] = '{32'hc1ea7f23, 32'h428d40dc, 32'hc29fe2dc, 32'h41950740, 32'h41d915af, 32'hc2a07b91, 32'hc290e745, 32'h425607e9};
test_output[4093] = '{32'h428d40dc};
test_index[4093] = '{1};
test_input[32752:32759] = '{32'hc2543922, 32'hc2379d30, 32'hc212ce6d, 32'h4230583a, 32'hc28c58e9, 32'h42805956, 32'h4282ae9b, 32'hc28ad8b4};
test_output[4094] = '{32'h4282ae9b};
test_index[4094] = '{6};
test_input[32760:32767] = '{32'h41c07b0c, 32'hc2c791b5, 32'h428f8577, 32'h422a6724, 32'hc0f20c8c, 32'hc0830edc, 32'h410f4ec8, 32'hc183bacf};
test_output[4095] = '{32'h428f8577};
test_index[4095] = '{2};
test_input[32768:32775] = '{32'hc26d3583, 32'h4263941b, 32'h42c74f23, 32'h41e8fd54, 32'h41268fa1, 32'h42bbf921, 32'hc2a5d553, 32'h429f8b8b};
test_output[4096] = '{32'h42c74f23};
test_index[4096] = '{2};
test_input[32776:32783] = '{32'h42349e21, 32'h4237cd87, 32'h426f54d5, 32'hc2585e61, 32'h42b542f9, 32'h41923dcc, 32'h4299b875, 32'hc294f1a2};
test_output[4097] = '{32'h42b542f9};
test_index[4097] = '{4};
test_input[32784:32791] = '{32'hc1c8c058, 32'h4244068b, 32'h42b0e2e1, 32'hc1bc1f43, 32'hc29b79af, 32'h4287d8eb, 32'h42712bd4, 32'hc296f69f};
test_output[4098] = '{32'h42b0e2e1};
test_index[4098] = '{2};
test_input[32792:32799] = '{32'hc2b1dd62, 32'hc2a9ba3c, 32'h428019fb, 32'hc059dd87, 32'h40f23d6b, 32'hc24640c1, 32'hc2ab8c0d, 32'hc21e792b};
test_output[4099] = '{32'h428019fb};
test_index[4099] = '{2};
test_input[32800:32807] = '{32'hc281ad7b, 32'h424dfb78, 32'h3e7c6b69, 32'h4133fbd3, 32'h41bc6dec, 32'hc2220fd4, 32'hc10b9c4d, 32'h4209ee18};
test_output[4100] = '{32'h424dfb78};
test_index[4100] = '{1};
test_input[32808:32815] = '{32'h41bf2260, 32'hc2b73aa2, 32'h41966fdd, 32'hc13444fa, 32'h42b47433, 32'h42c31c76, 32'hc28ec966, 32'hc06b81d3};
test_output[4101] = '{32'h42c31c76};
test_index[4101] = '{5};
test_input[32816:32823] = '{32'h4088c9a9, 32'h4125eef5, 32'hc2619329, 32'hc2c2fc3d, 32'h4246aa0f, 32'h422ba310, 32'hc1847097, 32'h422aaff6};
test_output[4102] = '{32'h4246aa0f};
test_index[4102] = '{4};
test_input[32824:32831] = '{32'h42a0af9c, 32'h42c293e7, 32'h4293dd61, 32'h3eb90946, 32'h426a639d, 32'hc2a972ce, 32'hc2766452, 32'hc2b94992};
test_output[4103] = '{32'h42c293e7};
test_index[4103] = '{1};
test_input[32832:32839] = '{32'h41618365, 32'hc26b1058, 32'h427c085d, 32'h424f5b03, 32'h410d0870, 32'hc26f9825, 32'hc29e64c4, 32'hc29032e7};
test_output[4104] = '{32'h427c085d};
test_index[4104] = '{2};
test_input[32840:32847] = '{32'h423f3f3d, 32'hc218637e, 32'h428627bd, 32'h42a152a5, 32'hc252cbe6, 32'h420172a2, 32'h4244ee5f, 32'h421525e7};
test_output[4105] = '{32'h42a152a5};
test_index[4105] = '{3};
test_input[32848:32855] = '{32'h4168167d, 32'h41eabfac, 32'h425b12b0, 32'h426c35fe, 32'hc2567221, 32'h41af468f, 32'h4238ca62, 32'hc161ed34};
test_output[4106] = '{32'h426c35fe};
test_index[4106] = '{3};
test_input[32856:32863] = '{32'h4234c897, 32'h42c6a3a3, 32'hc27da905, 32'h41797ddd, 32'hc1ff35ef, 32'hc295b81a, 32'hc2855547, 32'h41967455};
test_output[4107] = '{32'h42c6a3a3};
test_index[4107] = '{1};
test_input[32864:32871] = '{32'hbf6bba2d, 32'h414cabb9, 32'hc2a448d5, 32'hc22b5b31, 32'hc28c7e42, 32'h3f15af52, 32'h4292b325, 32'hc22b69ed};
test_output[4108] = '{32'h4292b325};
test_index[4108] = '{6};
test_input[32872:32879] = '{32'hc2309adf, 32'hc299c268, 32'h42424ba4, 32'h41e0065f, 32'h408fcc58, 32'h429e1b3f, 32'h41fcd267, 32'h42bb5cd3};
test_output[4109] = '{32'h42bb5cd3};
test_index[4109] = '{7};
test_input[32880:32887] = '{32'hc26fd552, 32'h40ca0e15, 32'hc2682799, 32'hc28b50f1, 32'hc2bb3b50, 32'h410597a7, 32'h41b707a0, 32'hc19898e8};
test_output[4110] = '{32'h41b707a0};
test_index[4110] = '{6};
test_input[32888:32895] = '{32'hc2839a0a, 32'hc2494ec8, 32'hc2a5d4ad, 32'h42074840, 32'hc27b3376, 32'h422c03f8, 32'hc25aabe6, 32'h42be9e35};
test_output[4111] = '{32'h42be9e35};
test_index[4111] = '{7};
test_input[32896:32903] = '{32'h410bef84, 32'h4297f33a, 32'hc2138077, 32'h41dab1ba, 32'h428e48de, 32'hc26c701f, 32'hc2c1fa23, 32'hc10b585a};
test_output[4112] = '{32'h4297f33a};
test_index[4112] = '{1};
test_input[32904:32911] = '{32'h425aa5a1, 32'h42778e5c, 32'hc2a52ce5, 32'hc2147804, 32'hc1654a06, 32'hc245314d, 32'h4186faf5, 32'hc286d437};
test_output[4113] = '{32'h42778e5c};
test_index[4113] = '{1};
test_input[32912:32919] = '{32'h41d855b7, 32'h428d2394, 32'hc26d8c32, 32'h428be663, 32'hc10d92f5, 32'hc2970226, 32'hc22249a9, 32'hc1e0a293};
test_output[4114] = '{32'h428d2394};
test_index[4114] = '{1};
test_input[32920:32927] = '{32'h4213649a, 32'h42af0df2, 32'h423ad292, 32'h42bc673a, 32'hc28d849b, 32'hc14f206a, 32'h42c2a27f, 32'h42aa76ec};
test_output[4115] = '{32'h42c2a27f};
test_index[4115] = '{6};
test_input[32928:32935] = '{32'hc206bffb, 32'hc2bd60d0, 32'hc2b51572, 32'hc1972b38, 32'hc20a433e, 32'h42b8d08d, 32'h41ba007f, 32'hc1c4d202};
test_output[4116] = '{32'h42b8d08d};
test_index[4116] = '{5};
test_input[32936:32943] = '{32'hc238acab, 32'h42ab0311, 32'hc2b0a800, 32'h4279e834, 32'h403226e6, 32'h423fcb1e, 32'hc24600f2, 32'hc2c39986};
test_output[4117] = '{32'h42ab0311};
test_index[4117] = '{1};
test_input[32944:32951] = '{32'hc2bdea25, 32'h40903749, 32'h4280231e, 32'h42afffa6, 32'h3f83781c, 32'h41af414b, 32'h42994c3b, 32'h4215d323};
test_output[4118] = '{32'h42afffa6};
test_index[4118] = '{3};
test_input[32952:32959] = '{32'hc1cc4000, 32'h4277577a, 32'hc215e45e, 32'hc0249f38, 32'hc23a578b, 32'h4285cc68, 32'h42b28b7e, 32'hc235ef12};
test_output[4119] = '{32'h42b28b7e};
test_index[4119] = '{6};
test_input[32960:32967] = '{32'h41feb54c, 32'hc2c24182, 32'h412d44a3, 32'hc1db1ea2, 32'h41fd9077, 32'hc2adc3c7, 32'h42862f46, 32'hc19b1476};
test_output[4120] = '{32'h42862f46};
test_index[4120] = '{6};
test_input[32968:32975] = '{32'hc20cc698, 32'h42953049, 32'h426c72e3, 32'hc1d95a54, 32'h41c649ef, 32'h42075c96, 32'h4208df5d, 32'hc28f64ae};
test_output[4121] = '{32'h42953049};
test_index[4121] = '{1};
test_input[32976:32983] = '{32'h42c367bb, 32'hc2b23401, 32'hc2b49c64, 32'h42186cf4, 32'hc2baf756, 32'h4299a78e, 32'hc19d1092, 32'hc1989c06};
test_output[4122] = '{32'h42c367bb};
test_index[4122] = '{0};
test_input[32984:32991] = '{32'h42b49589, 32'h4295e8e2, 32'h41e8319c, 32'h42c152b5, 32'hc12ef0f4, 32'h42aa4147, 32'h42c3dc89, 32'h427de250};
test_output[4123] = '{32'h42c3dc89};
test_index[4123] = '{6};
test_input[32992:32999] = '{32'h423b1f4f, 32'hc23693ad, 32'h4229404c, 32'hc2b979bf, 32'h41917b94, 32'hc2af2313, 32'h424e4171, 32'hc1929c4d};
test_output[4124] = '{32'h424e4171};
test_index[4124] = '{6};
test_input[33000:33007] = '{32'h411abad2, 32'h41d694ad, 32'h428c73df, 32'hc1b0b675, 32'h424e524f, 32'hc28a3969, 32'h428fed1f, 32'hc1afb972};
test_output[4125] = '{32'h428fed1f};
test_index[4125] = '{6};
test_input[33008:33015] = '{32'h41b40e51, 32'hc1107daa, 32'h42a8e653, 32'hc288f816, 32'h4267600a, 32'hc228189f, 32'h422bbd91, 32'h42b008f3};
test_output[4126] = '{32'h42b008f3};
test_index[4126] = '{7};
test_input[33016:33023] = '{32'hc23ad021, 32'h41b9881a, 32'h422fd61b, 32'h428a8553, 32'hc2c386e1, 32'hc2ab1e3e, 32'h41d6e410, 32'hc273c111};
test_output[4127] = '{32'h428a8553};
test_index[4127] = '{3};
test_input[33024:33031] = '{32'h3fc32c72, 32'hc20e96aa, 32'hc21a8ca6, 32'h40b9f043, 32'hc29d5cb9, 32'h419f7f9b, 32'h4281caca, 32'hc27d46e5};
test_output[4128] = '{32'h4281caca};
test_index[4128] = '{6};
test_input[33032:33039] = '{32'h42966d0e, 32'h42a6b376, 32'h41b3af6f, 32'hc1e8ddad, 32'hc288378a, 32'hc091c1b7, 32'h429acfbd, 32'hc1f9a5da};
test_output[4129] = '{32'h42a6b376};
test_index[4129] = '{1};
test_input[33040:33047] = '{32'h40ebeb1a, 32'h41a245a1, 32'h3fbf7dc2, 32'hc250ff87, 32'h422e9e34, 32'h40af4038, 32'h42142219, 32'hc2544bce};
test_output[4130] = '{32'h422e9e34};
test_index[4130] = '{4};
test_input[33048:33055] = '{32'h42c12d23, 32'h4215f76b, 32'h420304e7, 32'h4081900c, 32'h42a7771f, 32'hc26b89eb, 32'hc17f51ce, 32'hc179f9c0};
test_output[4131] = '{32'h42c12d23};
test_index[4131] = '{0};
test_input[33056:33063] = '{32'hc055e2ac, 32'hc29224b6, 32'h4122cd12, 32'h414a867f, 32'hc298f39e, 32'hc276838b, 32'hc16966e4, 32'h420e59d5};
test_output[4132] = '{32'h420e59d5};
test_index[4132] = '{7};
test_input[33064:33071] = '{32'hc1142658, 32'hc200a85c, 32'h42b60ab9, 32'hc2603196, 32'hc29b070a, 32'hc2845e61, 32'h411138f4, 32'hc172e77d};
test_output[4133] = '{32'h42b60ab9};
test_index[4133] = '{2};
test_input[33072:33079] = '{32'h40d91d46, 32'hc177b6aa, 32'hc1849666, 32'h42bbfd5b, 32'h42671544, 32'hbfcb27a0, 32'h4231098c, 32'hc1f5679a};
test_output[4134] = '{32'h42bbfd5b};
test_index[4134] = '{3};
test_input[33080:33087] = '{32'hc2b5e1f3, 32'h40d5fe4c, 32'hc1e14aaa, 32'h4214ffd3, 32'h429bec90, 32'h425f0eab, 32'h4222c7e0, 32'hc28d211b};
test_output[4135] = '{32'h429bec90};
test_index[4135] = '{4};
test_input[33088:33095] = '{32'hc00e61f3, 32'h422e26c8, 32'h42683e37, 32'hc2befd11, 32'h426100fb, 32'hc1cdcd0f, 32'h420478d2, 32'h42068a97};
test_output[4136] = '{32'h42683e37};
test_index[4136] = '{2};
test_input[33096:33103] = '{32'hc26b47a1, 32'h428364bf, 32'h4032c7a0, 32'h42addc97, 32'hc291ba98, 32'hc29ac149, 32'hc2bdd84f, 32'hc1a289b1};
test_output[4137] = '{32'h42addc97};
test_index[4137] = '{3};
test_input[33104:33111] = '{32'h4251afc6, 32'h42888f4b, 32'h4224850b, 32'h42bba55f, 32'hc234d13a, 32'hc2c673dd, 32'hc2b17acc, 32'hc2c15cfa};
test_output[4138] = '{32'h42bba55f};
test_index[4138] = '{3};
test_input[33112:33119] = '{32'h4297da8e, 32'h42828798, 32'h42b62f16, 32'h42a9ab38, 32'hc24f5532, 32'hc25dc673, 32'h42358a61, 32'hc2b47343};
test_output[4139] = '{32'h42b62f16};
test_index[4139] = '{2};
test_input[33120:33127] = '{32'hc29082b6, 32'hc2b0dd82, 32'h42a4903f, 32'hc25057e0, 32'h41d2b1cb, 32'h426fe28f, 32'hc1a94fdd, 32'h426901eb};
test_output[4140] = '{32'h42a4903f};
test_index[4140] = '{2};
test_input[33128:33135] = '{32'hc1b9061c, 32'hc159fe74, 32'hc287efb2, 32'hc18da13c, 32'h409a0244, 32'hc1a7e4fe, 32'hc23cdecb, 32'hc2540d9c};
test_output[4141] = '{32'h409a0244};
test_index[4141] = '{4};
test_input[33136:33143] = '{32'hc298f02d, 32'h421b5f4f, 32'hc220448b, 32'h40d895bd, 32'h42157e5e, 32'h429bb48a, 32'hc1c32610, 32'h423ca5a1};
test_output[4142] = '{32'h429bb48a};
test_index[4142] = '{5};
test_input[33144:33151] = '{32'hc2808aa6, 32'h42aa022e, 32'hc1ad1204, 32'h4218dfcb, 32'hc20bf19d, 32'h40bdae8d, 32'hc27e2782, 32'h42781f44};
test_output[4143] = '{32'h42aa022e};
test_index[4143] = '{1};
test_input[33152:33159] = '{32'hc242c4a8, 32'h42a8b883, 32'h4289ec05, 32'hc2b7fbe3, 32'hc2b70288, 32'h41aa7a64, 32'h42282ae2, 32'hc06eba27};
test_output[4144] = '{32'h42a8b883};
test_index[4144] = '{1};
test_input[33160:33167] = '{32'h42c6b170, 32'h42a9bd69, 32'h41ea8b18, 32'h42a16e22, 32'hc291439f, 32'h429ca869, 32'hc2b591dd, 32'hbf4a80be};
test_output[4145] = '{32'h42c6b170};
test_index[4145] = '{0};
test_input[33168:33175] = '{32'h4215822b, 32'hc29419b8, 32'h42a4eabe, 32'hc2c74832, 32'h429bf706, 32'hc21e3aa7, 32'h42636884, 32'hc01c19b6};
test_output[4146] = '{32'h42a4eabe};
test_index[4146] = '{2};
test_input[33176:33183] = '{32'h429eed50, 32'hc27043d2, 32'h425e43a9, 32'h4257ad29, 32'h42c57e34, 32'h41b9b988, 32'hc2afa64a, 32'h3ea8d5fb};
test_output[4147] = '{32'h42c57e34};
test_index[4147] = '{4};
test_input[33184:33191] = '{32'hc125643d, 32'hc2bf833e, 32'h41e35f77, 32'hc2c55af5, 32'h4202141f, 32'h42b21382, 32'h4277db13, 32'h4201880c};
test_output[4148] = '{32'h42b21382};
test_index[4148] = '{5};
test_input[33192:33199] = '{32'hc15a023a, 32'h424c1a82, 32'h41ca410b, 32'hc2c10786, 32'hc219edfd, 32'h42627701, 32'h4288db70, 32'h41d486af};
test_output[4149] = '{32'h4288db70};
test_index[4149] = '{6};
test_input[33200:33207] = '{32'hc2b7c532, 32'h40cd3736, 32'h42a3fff2, 32'h41ec1f31, 32'hc0ee0bec, 32'hc2969402, 32'h425fb3bf, 32'hc2ab2c51};
test_output[4150] = '{32'h42a3fff2};
test_index[4150] = '{2};
test_input[33208:33215] = '{32'hc0de7f76, 32'h4281d73f, 32'h42bfbd54, 32'h40d16f62, 32'hc19cb702, 32'h41885bd7, 32'h428d552f, 32'hc1d6e6ef};
test_output[4151] = '{32'h42bfbd54};
test_index[4151] = '{2};
test_input[33216:33223] = '{32'h42b7cc55, 32'hc27ddc82, 32'hc1b25079, 32'h40adb120, 32'hc1040d6e, 32'h42aa0c2e, 32'hc2b1a1ca, 32'h41092641};
test_output[4152] = '{32'h42b7cc55};
test_index[4152] = '{0};
test_input[33224:33231] = '{32'hc1ccb888, 32'hc1d3e593, 32'hc21f606a, 32'h423832fe, 32'h41df6ffd, 32'h428042f4, 32'hc227a274, 32'hc28dc864};
test_output[4153] = '{32'h428042f4};
test_index[4153] = '{5};
test_input[33232:33239] = '{32'h4267384a, 32'h429f9a9b, 32'h408ffca2, 32'h42980654, 32'h42610bc9, 32'h41b25e28, 32'h403058c4, 32'h41a479e2};
test_output[4154] = '{32'h429f9a9b};
test_index[4154] = '{1};
test_input[33240:33247] = '{32'h425776c7, 32'h423c15e8, 32'hc2a3960d, 32'h425628eb, 32'hc1ca2844, 32'hc2036181, 32'h424ed2cd, 32'h42962522};
test_output[4155] = '{32'h42962522};
test_index[4155] = '{7};
test_input[33248:33255] = '{32'hc2a666a1, 32'h41407502, 32'h41182fdd, 32'h429bb4cc, 32'h42aff27d, 32'h425c7ebd, 32'hc1a1664e, 32'hc06f6220};
test_output[4156] = '{32'h42aff27d};
test_index[4156] = '{4};
test_input[33256:33263] = '{32'h42b74cc5, 32'hc227aad2, 32'hc28374d7, 32'hc09b263d, 32'h429bb87a, 32'hc2b9db20, 32'h42ad8d6b, 32'h420b370f};
test_output[4157] = '{32'h42b74cc5};
test_index[4157] = '{0};
test_input[33264:33271] = '{32'hc2b51c5c, 32'h42440105, 32'hc296ae1b, 32'hc21eb34e, 32'h4252a2a2, 32'h40e7aca3, 32'h41e93290, 32'hc0f6f516};
test_output[4158] = '{32'h4252a2a2};
test_index[4158] = '{4};
test_input[33272:33279] = '{32'hc24a043f, 32'hc2c41bdf, 32'h4222dcbd, 32'h410afcc5, 32'h418d3999, 32'hc23eb87a, 32'hc284c6ea, 32'hc261ff0a};
test_output[4159] = '{32'h4222dcbd};
test_index[4159] = '{2};
test_input[33280:33287] = '{32'h42771856, 32'hc1934b1d, 32'hc2997ff8, 32'h4270fa52, 32'h4182bcbd, 32'hc242c783, 32'h42c211e2, 32'h429384cf};
test_output[4160] = '{32'h42c211e2};
test_index[4160] = '{6};
test_input[33288:33295] = '{32'hc2a30109, 32'hc2300a19, 32'hc29ac4fa, 32'hc27ba0e0, 32'hc2a4dee8, 32'h4130b6bc, 32'h422a7031, 32'hc24d05e9};
test_output[4161] = '{32'h422a7031};
test_index[4161] = '{6};
test_input[33296:33303] = '{32'hc2c13f55, 32'hc04445cd, 32'hc2a95e5b, 32'h41a5e971, 32'hc29ae7ba, 32'hc22a2e9a, 32'h4042dcef, 32'hc2ab7165};
test_output[4162] = '{32'h41a5e971};
test_index[4162] = '{3};
test_input[33304:33311] = '{32'h420e1d25, 32'hc29bfa35, 32'hc2ab61bb, 32'h42950cbd, 32'h424de2e1, 32'h418eb74a, 32'h428e30f0, 32'h406305ed};
test_output[4163] = '{32'h42950cbd};
test_index[4163] = '{3};
test_input[33312:33319] = '{32'hc28f5ea0, 32'hc298e532, 32'h42391535, 32'hc2b7f16a, 32'h42789579, 32'h40d2d3d9, 32'hc255b8a4, 32'h421f3eee};
test_output[4164] = '{32'h42789579};
test_index[4164] = '{4};
test_input[33320:33327] = '{32'hc13d1dc0, 32'hc1c031b6, 32'hc0df5846, 32'hc2b24d2a, 32'h4123c6c7, 32'hc240a7b0, 32'h41aa58b0, 32'hc200db01};
test_output[4165] = '{32'h41aa58b0};
test_index[4165] = '{6};
test_input[33328:33335] = '{32'hc20a8e72, 32'h41dc1f27, 32'hc24f97ab, 32'hc1ec4144, 32'h420a663d, 32'h42b6a1b5, 32'hc239c21f, 32'hc1e9d510};
test_output[4166] = '{32'h42b6a1b5};
test_index[4166] = '{5};
test_input[33336:33343] = '{32'h41692b9f, 32'h4284c5d0, 32'h427567d1, 32'h42586ba7, 32'h4296b258, 32'hc2b362d7, 32'hc2a74c2a, 32'hc1924f13};
test_output[4167] = '{32'h4296b258};
test_index[4167] = '{4};
test_input[33344:33351] = '{32'hc279671d, 32'hc1fa55a5, 32'hc28d971e, 32'h4212bc06, 32'h4274002b, 32'h41ed5f93, 32'h428e75a0, 32'h42c7bc20};
test_output[4168] = '{32'h42c7bc20};
test_index[4168] = '{7};
test_input[33352:33359] = '{32'h42288d51, 32'h42a8ee84, 32'hc19002e3, 32'hc290e746, 32'hc1db16bc, 32'hc2aa0709, 32'h4248b4bf, 32'hc28f295d};
test_output[4169] = '{32'h42a8ee84};
test_index[4169] = '{1};
test_input[33360:33367] = '{32'h414d2a7f, 32'h428f66ea, 32'h4224c22a, 32'h423032fb, 32'hc2b27462, 32'hc255cc3a, 32'h42b30c12, 32'hc283196d};
test_output[4170] = '{32'h42b30c12};
test_index[4170] = '{6};
test_input[33368:33375] = '{32'hc225aa69, 32'h4284abd7, 32'hc26aa643, 32'hc1135033, 32'h424234c3, 32'h4249695b, 32'h4222f1d7, 32'hc29bf4c9};
test_output[4171] = '{32'h4284abd7};
test_index[4171] = '{1};
test_input[33376:33383] = '{32'h41556749, 32'hc2868fe6, 32'h429740a9, 32'hc2943ead, 32'hc247945d, 32'h41a6b1f0, 32'h40685a67, 32'hc223c5d3};
test_output[4172] = '{32'h429740a9};
test_index[4172] = '{2};
test_input[33384:33391] = '{32'h422ff141, 32'h42519d80, 32'h401a655f, 32'hc2943d1c, 32'hc1af7733, 32'hc29e3f13, 32'hc2b64035, 32'h41161526};
test_output[4173] = '{32'h42519d80};
test_index[4173] = '{1};
test_input[33392:33399] = '{32'h415817d7, 32'hc23653ff, 32'hc25cae46, 32'h426ab12e, 32'hc291dfad, 32'hc25e78a3, 32'hc1646d20, 32'hc0dc9d9f};
test_output[4174] = '{32'h426ab12e};
test_index[4174] = '{3};
test_input[33400:33407] = '{32'h42527065, 32'hc204fd5d, 32'hc1d72ab5, 32'hc21e3962, 32'hc232987e, 32'h42a25dab, 32'hc27516d8, 32'h4226c4f3};
test_output[4175] = '{32'h42a25dab};
test_index[4175] = '{5};
test_input[33408:33415] = '{32'hc246d500, 32'hc1b22447, 32'h41f2c2a1, 32'h4247d6c5, 32'h422c0d46, 32'hc1a31fcf, 32'h425f5233, 32'hc292296b};
test_output[4176] = '{32'h425f5233};
test_index[4176] = '{6};
test_input[33416:33423] = '{32'hc12932a3, 32'hc23e2329, 32'h424ee29b, 32'h41be1d8b, 32'hc2c6e403, 32'h3ff5de88, 32'h42502177, 32'hc280a1d5};
test_output[4177] = '{32'h42502177};
test_index[4177] = '{6};
test_input[33424:33431] = '{32'h41be957a, 32'h4264322d, 32'hc28c6b01, 32'h41a74d6c, 32'hc2084f8a, 32'hc0b7fc47, 32'h4265781b, 32'h42092912};
test_output[4178] = '{32'h4265781b};
test_index[4178] = '{6};
test_input[33432:33439] = '{32'hc2919338, 32'h42a5d980, 32'hc10c46a7, 32'h412b288e, 32'h4069b34b, 32'hc1037af8, 32'hc2b22d16, 32'hbf32e582};
test_output[4179] = '{32'h42a5d980};
test_index[4179] = '{1};
test_input[33440:33447] = '{32'h41c982a2, 32'hc0d8895c, 32'h42b4881d, 32'h4295e32f, 32'h408d945d, 32'hc2885f5d, 32'hc1ef47ff, 32'h42c773d8};
test_output[4180] = '{32'h42c773d8};
test_index[4180] = '{7};
test_input[33448:33455] = '{32'h4255feac, 32'hc167fd72, 32'h42397620, 32'h425bf5a5, 32'hc1a53d5a, 32'hc2b4fd58, 32'h428ee97d, 32'hc286ef8c};
test_output[4181] = '{32'h428ee97d};
test_index[4181] = '{6};
test_input[33456:33463] = '{32'hc293a58f, 32'h42c17a70, 32'hc1dbd9a9, 32'h42a1fc25, 32'h406ac456, 32'h4207ede8, 32'h4246202a, 32'h4282bfae};
test_output[4182] = '{32'h42c17a70};
test_index[4182] = '{1};
test_input[33464:33471] = '{32'hc2b5fc3a, 32'hc2b23653, 32'hc29e5c9f, 32'hc10f6af3, 32'hc2a49776, 32'h42560c43, 32'hc28bb65b, 32'h42b9aa80};
test_output[4183] = '{32'h42b9aa80};
test_index[4183] = '{7};
test_input[33472:33479] = '{32'hc1489156, 32'h4153732a, 32'hc2783756, 32'hc24c47f1, 32'h41d5024c, 32'h4017c714, 32'h4216bf0b, 32'h42b51a4b};
test_output[4184] = '{32'h42b51a4b};
test_index[4184] = '{7};
test_input[33480:33487] = '{32'h429cc7db, 32'h4265c271, 32'hc2b18bba, 32'h42b9ca62, 32'h42981fe1, 32'h427116aa, 32'h41a35b7b, 32'hc116b2a0};
test_output[4185] = '{32'h42b9ca62};
test_index[4185] = '{3};
test_input[33488:33495] = '{32'h422b0c86, 32'h42c1deb5, 32'hc1f8f931, 32'h412f38ab, 32'h4283558b, 32'hc271a196, 32'hc0a8d3d1, 32'h422a6ab5};
test_output[4186] = '{32'h42c1deb5};
test_index[4186] = '{1};
test_input[33496:33503] = '{32'hc196ec58, 32'h4287244c, 32'hc234bc57, 32'h42a3715f, 32'hc12b1db0, 32'h419d9513, 32'h42c5db88, 32'hc2b2c011};
test_output[4187] = '{32'h42c5db88};
test_index[4187] = '{6};
test_input[33504:33511] = '{32'hc2021ca3, 32'h421d7c6a, 32'h424dd11d, 32'h42421fea, 32'hc2048ea2, 32'h4174c4c4, 32'hc073527c, 32'h42b1db1f};
test_output[4188] = '{32'h42b1db1f};
test_index[4188] = '{7};
test_input[33512:33519] = '{32'h42a26c52, 32'hc15e3d2d, 32'hc2a91a39, 32'h42197f22, 32'h41f52605, 32'h42ab25a0, 32'h42b8deb1, 32'h42207348};
test_output[4189] = '{32'h42b8deb1};
test_index[4189] = '{6};
test_input[33520:33527] = '{32'hc2a66407, 32'hc25f8277, 32'hc067c28e, 32'h413f33f9, 32'hc2b14851, 32'h41b93769, 32'hc2a39305, 32'h42267172};
test_output[4190] = '{32'h42267172};
test_index[4190] = '{7};
test_input[33528:33535] = '{32'hc2b2aa80, 32'hc2b64841, 32'hc2401dc2, 32'hc11e7155, 32'h428ab789, 32'hc2231955, 32'h42c2da58, 32'hc29eb730};
test_output[4191] = '{32'h42c2da58};
test_index[4191] = '{6};
test_input[33536:33543] = '{32'hc29ca17c, 32'h42090728, 32'hc18e7e57, 32'hc2a3a575, 32'hc288dbd3, 32'h3ff051d8, 32'h42761e43, 32'hc17de0d4};
test_output[4192] = '{32'h42761e43};
test_index[4192] = '{6};
test_input[33544:33551] = '{32'h410c5d0a, 32'h423d78a7, 32'hc2107c83, 32'hc2c628c7, 32'h42a9a506, 32'h417becd0, 32'hc2bff715, 32'h42582718};
test_output[4193] = '{32'h42a9a506};
test_index[4193] = '{4};
test_input[33552:33559] = '{32'hc2703de1, 32'h421ae5bb, 32'hc2781b1c, 32'h4293719b, 32'h42345ad8, 32'hc2c5f968, 32'h428c737a, 32'h4241c2d0};
test_output[4194] = '{32'h4293719b};
test_index[4194] = '{3};
test_input[33560:33567] = '{32'h429cc648, 32'hc200cfa1, 32'h42b0fb85, 32'hc260019c, 32'h42b905ca, 32'h429b3830, 32'h428bcc51, 32'hc2968696};
test_output[4195] = '{32'h42b905ca};
test_index[4195] = '{4};
test_input[33568:33575] = '{32'hc1c732ac, 32'h4107504a, 32'hc29e2bbd, 32'h42823c38, 32'hc1d13a20, 32'h41a74263, 32'h405220a2, 32'hc2ac3897};
test_output[4196] = '{32'h42823c38};
test_index[4196] = '{3};
test_input[33576:33583] = '{32'h411e8f8b, 32'hc1b57669, 32'h4101e040, 32'h417594b8, 32'hc090d6d4, 32'h423cc623, 32'hc2181fca, 32'hc12f41b2};
test_output[4197] = '{32'h423cc623};
test_index[4197] = '{5};
test_input[33584:33591] = '{32'hc282e8f6, 32'h429dcc5d, 32'hc10ac3f5, 32'hc2b6f82c, 32'h424105e3, 32'h42b6f058, 32'hc2a06e6a, 32'h4257fcd3};
test_output[4198] = '{32'h42b6f058};
test_index[4198] = '{5};
test_input[33592:33599] = '{32'hc29e0d0a, 32'h4281a1c6, 32'h420272e4, 32'hc1e8122a, 32'h42769723, 32'hc0f825c3, 32'hc2bad081, 32'hc22cc105};
test_output[4199] = '{32'h4281a1c6};
test_index[4199] = '{1};
test_input[33600:33607] = '{32'hc1bfb78a, 32'hc0432afd, 32'h429a79fc, 32'h41914a2f, 32'h422e3e42, 32'h4197e523, 32'h410de4b3, 32'h42bfafc8};
test_output[4200] = '{32'h42bfafc8};
test_index[4200] = '{7};
test_input[33608:33615] = '{32'hc1b60ecd, 32'h4221b362, 32'h42c5e04b, 32'h4281b4f6, 32'hc2bfc30d, 32'hc1f4df4d, 32'h42255364, 32'hc0cc2142};
test_output[4201] = '{32'h42c5e04b};
test_index[4201] = '{2};
test_input[33616:33623] = '{32'hc273fea4, 32'hc24974a5, 32'h4298b51b, 32'h4043b1a3, 32'hc2b7b009, 32'hc2c161ce, 32'hc1b412a4, 32'h42a78ea9};
test_output[4202] = '{32'h42a78ea9};
test_index[4202] = '{7};
test_input[33624:33631] = '{32'hc2a40bb9, 32'hc2a71c43, 32'hc1fe1351, 32'hc1fd8155, 32'hc2ad57cb, 32'hc0838072, 32'hbeb90786, 32'hc2bdb800};
test_output[4203] = '{32'hbeb90786};
test_index[4203] = '{6};
test_input[33632:33639] = '{32'h420c5964, 32'hc2bdbf69, 32'hc1c7a5a6, 32'h4122a05a, 32'h42b8bbe8, 32'h41239a32, 32'h42004179, 32'hc2c6c4bb};
test_output[4204] = '{32'h42b8bbe8};
test_index[4204] = '{4};
test_input[33640:33647] = '{32'h40bf580c, 32'h41e75c42, 32'h421419eb, 32'hc0ba3671, 32'hc279f9fe, 32'hc29ea203, 32'h421b95fd, 32'hc29b5f84};
test_output[4205] = '{32'h421b95fd};
test_index[4205] = '{6};
test_input[33648:33655] = '{32'hc0e505ad, 32'hc25ce970, 32'h420b799f, 32'h42c5cef2, 32'hc21d5c7d, 32'h40f57ed1, 32'hc1ecc38e, 32'h426361f2};
test_output[4206] = '{32'h42c5cef2};
test_index[4206] = '{3};
test_input[33656:33663] = '{32'hc189bd91, 32'hc1559590, 32'hc2b79557, 32'h42c1b5db, 32'hc235a01d, 32'h4240959a, 32'hc19190c7, 32'hc28c5ca8};
test_output[4207] = '{32'h42c1b5db};
test_index[4207] = '{3};
test_input[33664:33671] = '{32'hc270b16b, 32'h40cfd2fa, 32'h42983fd3, 32'hc1a154db, 32'hc0a15217, 32'hc168b556, 32'h4279f58c, 32'hc1a4f2a2};
test_output[4208] = '{32'h42983fd3};
test_index[4208] = '{2};
test_input[33672:33679] = '{32'hc2793cfd, 32'hc2c43082, 32'hc16a2fe6, 32'hc14fd3cf, 32'hc2b72297, 32'hc1cb0bc8, 32'h428b4ff5, 32'hc18640f0};
test_output[4209] = '{32'h428b4ff5};
test_index[4209] = '{6};
test_input[33680:33687] = '{32'h4284b37c, 32'h422abe98, 32'hc2957342, 32'hc28db5ab, 32'h42c52278, 32'hc27b1827, 32'hc1c6ab92, 32'h423d6803};
test_output[4210] = '{32'h42c52278};
test_index[4210] = '{4};
test_input[33688:33695] = '{32'h42ba2872, 32'hc282f4a5, 32'hc1e7a6ce, 32'h4274b9af, 32'hc2b0adab, 32'hc2442094, 32'hc2662463, 32'h4297f6a6};
test_output[4211] = '{32'h42ba2872};
test_index[4211] = '{0};
test_input[33696:33703] = '{32'hc1f584bf, 32'hc0100812, 32'h425e637c, 32'h42892033, 32'hc17c628a, 32'h410d99dc, 32'h427be68b, 32'hc2c4e144};
test_output[4212] = '{32'h42892033};
test_index[4212] = '{3};
test_input[33704:33711] = '{32'hc1dad4c6, 32'h42aa8634, 32'h41408f20, 32'h42bfbf9a, 32'h419880d3, 32'hc250f1c7, 32'h40c7d1a4, 32'hc2b6a9da};
test_output[4213] = '{32'h42bfbf9a};
test_index[4213] = '{3};
test_input[33712:33719] = '{32'h422b94c1, 32'h423b3782, 32'hc23ea7dd, 32'hc29f5a42, 32'h42247eab, 32'h41285db0, 32'h42850778, 32'h41f684f2};
test_output[4214] = '{32'h42850778};
test_index[4214] = '{6};
test_input[33720:33727] = '{32'h42628db3, 32'hc2bcc895, 32'h4200877b, 32'h41f72bc8, 32'h4181af1a, 32'hc2a69778, 32'hc2b464c3, 32'h4192299e};
test_output[4215] = '{32'h42628db3};
test_index[4215] = '{0};
test_input[33728:33735] = '{32'hc2946fdc, 32'hc2b934b8, 32'hc2896725, 32'h427246f0, 32'h4262e074, 32'hc0d54db1, 32'hc20840e2, 32'h41663c29};
test_output[4216] = '{32'h427246f0};
test_index[4216] = '{3};
test_input[33736:33743] = '{32'h429c6e79, 32'hc24ae89c, 32'hc29e10f0, 32'h426ee324, 32'h426a8ed4, 32'h42aa2515, 32'hc18af529, 32'h41e77a8d};
test_output[4217] = '{32'h42aa2515};
test_index[4217] = '{5};
test_input[33744:33751] = '{32'hc09efaff, 32'h4236ac3b, 32'hc2a1c462, 32'h426adda5, 32'hc2158f3b, 32'hc27447da, 32'h42990ffb, 32'hc2a987f2};
test_output[4218] = '{32'h42990ffb};
test_index[4218] = '{6};
test_input[33752:33759] = '{32'hc2011f1e, 32'h4256aac3, 32'hc2a4796a, 32'h424f3b49, 32'hc2c25fee, 32'h42879010, 32'h41876522, 32'hc2667ff9};
test_output[4219] = '{32'h42879010};
test_index[4219] = '{5};
test_input[33760:33767] = '{32'h41c55092, 32'hc295048f, 32'h4254603b, 32'hc1a0e731, 32'h421e1861, 32'hc1e7e24f, 32'h41003ede, 32'hbffd3df2};
test_output[4220] = '{32'h4254603b};
test_index[4220] = '{2};
test_input[33768:33775] = '{32'h4220e8d5, 32'hc11b94ca, 32'h423a6c09, 32'hc2bd63ff, 32'hc203be5f, 32'hc22e77e0, 32'h429046ad, 32'hc2b7a130};
test_output[4221] = '{32'h429046ad};
test_index[4221] = '{6};
test_input[33776:33783] = '{32'h422bbc94, 32'hc291e246, 32'hc227b7d8, 32'hc1992735, 32'h42912539, 32'hc20c7162, 32'hc1b61012, 32'h41bd64e4};
test_output[4222] = '{32'h42912539};
test_index[4222] = '{4};
test_input[33784:33791] = '{32'hc2655d62, 32'hc26b619e, 32'hc1b06997, 32'hc1503870, 32'h4138cb98, 32'h41df9242, 32'h40d4fa60, 32'hc2b40bb6};
test_output[4223] = '{32'h41df9242};
test_index[4223] = '{5};
test_input[33792:33799] = '{32'h41955857, 32'hc2a63dbe, 32'hc1e178df, 32'h40d1b5f5, 32'h425c78a9, 32'h4256ab15, 32'h4211a6bd, 32'h42933b1d};
test_output[4224] = '{32'h42933b1d};
test_index[4224] = '{7};
test_input[33800:33807] = '{32'h41ac9cf0, 32'h429d6a40, 32'hc2b0d452, 32'h429498aa, 32'hc27e47cc, 32'h428ff450, 32'h41cdbde2, 32'hc29cc866};
test_output[4225] = '{32'h429d6a40};
test_index[4225] = '{1};
test_input[33808:33815] = '{32'h41af2d00, 32'hc2c397f7, 32'h421c3e8e, 32'hc285e9d0, 32'hc297d19a, 32'hc28504a4, 32'hc2c11390, 32'hc2bcc8ce};
test_output[4226] = '{32'h421c3e8e};
test_index[4226] = '{2};
test_input[33816:33823] = '{32'h40534740, 32'h42916402, 32'hc08ebf1f, 32'h42a533d8, 32'h42b81eab, 32'hc23c3809, 32'h419ae7f6, 32'h41e0b146};
test_output[4227] = '{32'h42b81eab};
test_index[4227] = '{4};
test_input[33824:33831] = '{32'hc082e9ec, 32'h41bbc652, 32'hc1864e92, 32'h429301ed, 32'h42b8a023, 32'hc14f5a6e, 32'hc109f627, 32'hc14232c3};
test_output[4228] = '{32'h42b8a023};
test_index[4228] = '{4};
test_input[33832:33839] = '{32'hc07e3550, 32'hc1cb84a7, 32'hc25f421a, 32'h41cfdf36, 32'hc2623013, 32'h4189ffae, 32'hc126a7be, 32'h424b0e13};
test_output[4229] = '{32'h424b0e13};
test_index[4229] = '{7};
test_input[33840:33847] = '{32'h42a44841, 32'h41a046b6, 32'hc2b9e311, 32'h42b9b73c, 32'hc2c665f0, 32'hc2c16f18, 32'h41aa3f0a, 32'h417485e9};
test_output[4230] = '{32'h42b9b73c};
test_index[4230] = '{3};
test_input[33848:33855] = '{32'hc282f64f, 32'hc2b62990, 32'h426bf2d7, 32'hc243790b, 32'hc1ef4112, 32'hc19ee3e9, 32'hc1773bdf, 32'hc1191850};
test_output[4231] = '{32'h426bf2d7};
test_index[4231] = '{2};
test_input[33856:33863] = '{32'h428909f2, 32'hc256bf84, 32'hc21079ea, 32'h42381884, 32'h40da2891, 32'h429a8098, 32'h420809c4, 32'h42a5e073};
test_output[4232] = '{32'h42a5e073};
test_index[4232] = '{7};
test_input[33864:33871] = '{32'hc0271f26, 32'h41b1af66, 32'h42785e24, 32'h4290b0a0, 32'h414b7b0f, 32'hc2c6d9a7, 32'h42841402, 32'h4271c57c};
test_output[4233] = '{32'h4290b0a0};
test_index[4233] = '{3};
test_input[33872:33879] = '{32'hc26e3fcb, 32'h40cd2624, 32'hc2a0c733, 32'h42a92133, 32'hc1b3f5ed, 32'hc26e1a3a, 32'hc2221100, 32'hc08412f1};
test_output[4234] = '{32'h42a92133};
test_index[4234] = '{3};
test_input[33880:33887] = '{32'h42c69bbe, 32'h41312d99, 32'hc296de91, 32'hc2644404, 32'h42b8abb9, 32'h4252b37a, 32'h42b52d68, 32'h426af77c};
test_output[4235] = '{32'h42c69bbe};
test_index[4235] = '{0};
test_input[33888:33895] = '{32'h42a8ae64, 32'hc2918199, 32'h420f492f, 32'hc1e0d500, 32'h41f70d83, 32'h426bc109, 32'h42490ad5, 32'hc293d953};
test_output[4236] = '{32'h42a8ae64};
test_index[4236] = '{0};
test_input[33896:33903] = '{32'hc2c363c3, 32'hc27c3201, 32'hc20f0eec, 32'hc1e258eb, 32'h414f6776, 32'h422113f6, 32'h42598ac7, 32'h4278303d};
test_output[4237] = '{32'h4278303d};
test_index[4237] = '{7};
test_input[33904:33911] = '{32'h414e42f1, 32'hc0c6f4d1, 32'h41764001, 32'h426d670a, 32'h42aadbec, 32'hc27d9750, 32'hbfcda94c, 32'hc233dc93};
test_output[4238] = '{32'h42aadbec};
test_index[4238] = '{4};
test_input[33912:33919] = '{32'hc286e5bf, 32'h4150bfba, 32'hc2b9aa1d, 32'hc26a5be0, 32'hc2a00c60, 32'hc1308bef, 32'hc256ee1a, 32'h41a3a846};
test_output[4239] = '{32'h41a3a846};
test_index[4239] = '{7};
test_input[33920:33927] = '{32'h41de4384, 32'h40f45671, 32'hc1146802, 32'hc28cc80e, 32'hc218e720, 32'hc2ad95c4, 32'h42bfe776, 32'h42454179};
test_output[4240] = '{32'h42bfe776};
test_index[4240] = '{6};
test_input[33928:33935] = '{32'h40a3f0c2, 32'hc295d06e, 32'h42a14ab3, 32'hc2b267aa, 32'h427647ad, 32'h42b6bdf4, 32'hc25d921f, 32'hbfd70f1b};
test_output[4241] = '{32'h42b6bdf4};
test_index[4241] = '{5};
test_input[33936:33943] = '{32'hc22cf034, 32'h41fe87e0, 32'hc2307130, 32'hc28f8696, 32'hc291021d, 32'h419b42dc, 32'h40f8703d, 32'hc2a211f9};
test_output[4242] = '{32'h41fe87e0};
test_index[4242] = '{1};
test_input[33944:33951] = '{32'h42491d6d, 32'h4208e410, 32'hc2874fbe, 32'h42c49f3f, 32'h42162e9e, 32'h412ca550, 32'h424a1ee5, 32'h420c3e9c};
test_output[4243] = '{32'h42c49f3f};
test_index[4243] = '{3};
test_input[33952:33959] = '{32'hc25e197a, 32'h42ab02cb, 32'h427475bb, 32'h426df969, 32'hc0c829a3, 32'hc28850d9, 32'hc2b27ca5, 32'h420ff35c};
test_output[4244] = '{32'h42ab02cb};
test_index[4244] = '{1};
test_input[33960:33967] = '{32'hc2c3f65c, 32'hc2274b85, 32'h42125036, 32'h421991f8, 32'h420e83bb, 32'hc11b8693, 32'h4236f194, 32'h42a85ad5};
test_output[4245] = '{32'h42a85ad5};
test_index[4245] = '{7};
test_input[33968:33975] = '{32'hc1e639ce, 32'hc29c4ef7, 32'hc1c43c11, 32'hc26ed2a8, 32'hc2abee06, 32'hc2a21c7d, 32'hc20a2b23, 32'h42915aaf};
test_output[4246] = '{32'h42915aaf};
test_index[4246] = '{7};
test_input[33976:33983] = '{32'hc2c66135, 32'hc297ce56, 32'hc21faf90, 32'h424a2515, 32'hc2b6f375, 32'h41df63f3, 32'h3fc1a2ab, 32'hc2b279bd};
test_output[4247] = '{32'h424a2515};
test_index[4247] = '{3};
test_input[33984:33991] = '{32'h42451f44, 32'h4279a8c9, 32'h421cce85, 32'h4287ca15, 32'h429bd427, 32'h428b012d, 32'hc28711b1, 32'hc2b8b0de};
test_output[4248] = '{32'h429bd427};
test_index[4248] = '{4};
test_input[33992:33999] = '{32'h428ab188, 32'h424666e8, 32'hc2a516f3, 32'h42b0ca06, 32'h41b07051, 32'h404eedec, 32'h4254a985, 32'h42b7f499};
test_output[4249] = '{32'h42b7f499};
test_index[4249] = '{7};
test_input[34000:34007] = '{32'h4073d888, 32'hc1fd22fd, 32'h41c96af4, 32'hc2a2f659, 32'hc24815b4, 32'h425c5655, 32'hc2c74b27, 32'h42792bde};
test_output[4250] = '{32'h42792bde};
test_index[4250] = '{7};
test_input[34008:34015] = '{32'h42a1caa4, 32'h41d1edf9, 32'hc244d99d, 32'h42b2ef3e, 32'hc28252f5, 32'hc2809b9d, 32'h41df7177, 32'hc22ed0fe};
test_output[4251] = '{32'h42b2ef3e};
test_index[4251] = '{3};
test_input[34016:34023] = '{32'h429ab093, 32'h42ad0193, 32'h424bcf2a, 32'hc25c2723, 32'h419b6e6d, 32'h4295f862, 32'hc2a299cc, 32'hc188bd65};
test_output[4252] = '{32'h42ad0193};
test_index[4252] = '{1};
test_input[34024:34031] = '{32'h422263df, 32'h42a758da, 32'hc2bff88b, 32'hc28bd261, 32'h4285d9d8, 32'h42164207, 32'h42bd8251, 32'h41a6b072};
test_output[4253] = '{32'h42bd8251};
test_index[4253] = '{6};
test_input[34032:34039] = '{32'hc14797c5, 32'hc20f69b2, 32'hc2c2182e, 32'h425a17c0, 32'hc22b84d9, 32'hc1c5c8fd, 32'h40966255, 32'h42a6a4fc};
test_output[4254] = '{32'h42a6a4fc};
test_index[4254] = '{7};
test_input[34040:34047] = '{32'hc2b7d3ed, 32'hc17601f7, 32'h41f62a56, 32'hc19a3cd3, 32'h42b377d7, 32'hbef7a50e, 32'h416d4962, 32'hc20f5e12};
test_output[4255] = '{32'h42b377d7};
test_index[4255] = '{4};
test_input[34048:34055] = '{32'h42b074c7, 32'hc2bb1edd, 32'hc15a1756, 32'hc158d9a7, 32'h414d45c4, 32'hc2430a3c, 32'hc270b1ad, 32'hc27e8276};
test_output[4256] = '{32'h42b074c7};
test_index[4256] = '{0};
test_input[34056:34063] = '{32'hc1c34e61, 32'hc2c1eb4a, 32'h4254da92, 32'hc18ee320, 32'h419e3c75, 32'hc2937706, 32'h4152d6e2, 32'h428224c4};
test_output[4257] = '{32'h428224c4};
test_index[4257] = '{7};
test_input[34064:34071] = '{32'h42a40f03, 32'h4261debf, 32'h42040aff, 32'h4046c3ee, 32'hc2bac576, 32'hc2b3dd27, 32'hc2a2d4ff, 32'hc2af420f};
test_output[4258] = '{32'h42a40f03};
test_index[4258] = '{0};
test_input[34072:34079] = '{32'h4182d46e, 32'h4124b313, 32'hc2ba308e, 32'hc281e9a1, 32'hc2bfad40, 32'hc1104781, 32'h4223c10c, 32'hc15a1d62};
test_output[4259] = '{32'h4223c10c};
test_index[4259] = '{6};
test_input[34080:34087] = '{32'hc1e077a3, 32'hc2766448, 32'h42449f3c, 32'h42644f9f, 32'h4281e315, 32'h421ceaff, 32'h4231c6ed, 32'hc1108e9c};
test_output[4260] = '{32'h4281e315};
test_index[4260] = '{4};
test_input[34088:34095] = '{32'h41ec13f1, 32'hc25cedc9, 32'h41c71c70, 32'h4183df58, 32'h42c58827, 32'hc2b1533c, 32'h3fa238fd, 32'h42270f67};
test_output[4261] = '{32'h42c58827};
test_index[4261] = '{4};
test_input[34096:34103] = '{32'hc2c2cf45, 32'hc2a5d6e9, 32'h41d8f891, 32'hc1fc6d7c, 32'h41c0db41, 32'hc22b7307, 32'hc21965b8, 32'hc19aaa47};
test_output[4262] = '{32'h41d8f891};
test_index[4262] = '{2};
test_input[34104:34111] = '{32'hc20b65e2, 32'hc238788c, 32'h41e6f380, 32'h4252d472, 32'h414f7b0b, 32'hc2ba9b4c, 32'h42af0b26, 32'h42005c28};
test_output[4263] = '{32'h42af0b26};
test_index[4263] = '{6};
test_input[34112:34119] = '{32'hc2668c65, 32'hc11acfe9, 32'h422b440c, 32'h423e1ccd, 32'hc13550d6, 32'hc2c19fd0, 32'h41552d99, 32'h4265b267};
test_output[4264] = '{32'h4265b267};
test_index[4264] = '{7};
test_input[34120:34127] = '{32'h42b3c06f, 32'hc039276a, 32'h42a41aa0, 32'hc12384d1, 32'h404d062c, 32'hc2988db8, 32'hc1b09e15, 32'h41ed2c9e};
test_output[4265] = '{32'h42b3c06f};
test_index[4265] = '{0};
test_input[34128:34135] = '{32'hc2b310d0, 32'hc237ad9f, 32'h42432c7b, 32'hc29c8108, 32'hc0ebeedc, 32'hc18e4428, 32'h42bad52f, 32'hc2af60ae};
test_output[4266] = '{32'h42bad52f};
test_index[4266] = '{6};
test_input[34136:34143] = '{32'h428bab1d, 32'h421a4c6f, 32'h425d8a27, 32'h42babd94, 32'hc1d1826e, 32'hc1583717, 32'hc2795404, 32'hc2a156a6};
test_output[4267] = '{32'h42babd94};
test_index[4267] = '{3};
test_input[34144:34151] = '{32'h407fa58e, 32'hbf9f855f, 32'h42c2a0c2, 32'hc276b8b8, 32'h41bed24e, 32'hc1f94a74, 32'h4222011a, 32'h42806229};
test_output[4268] = '{32'h42c2a0c2};
test_index[4268] = '{2};
test_input[34152:34159] = '{32'hc1fe79a4, 32'hc29a2c48, 32'hc291616a, 32'h42ae919d, 32'hc28f0e1d, 32'h4243ab67, 32'h422be8df, 32'hc280b468};
test_output[4269] = '{32'h42ae919d};
test_index[4269] = '{3};
test_input[34160:34167] = '{32'h42879281, 32'h4140a471, 32'hc18cd9fe, 32'h41b66c9c, 32'h4145bbd6, 32'h429fdce2, 32'hc1a14f4a, 32'hc21ce445};
test_output[4270] = '{32'h429fdce2};
test_index[4270] = '{5};
test_input[34168:34175] = '{32'hc1f83a91, 32'hc1c27e4a, 32'h4233cfb3, 32'hc29b46ac, 32'hc2735c3c, 32'h4255a001, 32'hc2a5c344, 32'hc12d9451};
test_output[4271] = '{32'h4255a001};
test_index[4271] = '{5};
test_input[34176:34183] = '{32'h426d15d9, 32'h41d42871, 32'hc26d85c7, 32'h41e50666, 32'hc20832c9, 32'h42b22080, 32'hc1563571, 32'hc2446347};
test_output[4272] = '{32'h42b22080};
test_index[4272] = '{5};
test_input[34184:34191] = '{32'h42881905, 32'hc1209714, 32'hc20a4d43, 32'hc1c282b7, 32'hc28ffe26, 32'h41e43383, 32'h42c0b02b, 32'hc2c00b2e};
test_output[4273] = '{32'h42c0b02b};
test_index[4273] = '{6};
test_input[34192:34199] = '{32'h422de8be, 32'h428a5463, 32'hc28fdc7b, 32'hc204796d, 32'h42a33f41, 32'h4232284b, 32'hc221edf6, 32'h4244319b};
test_output[4274] = '{32'h42a33f41};
test_index[4274] = '{4};
test_input[34200:34207] = '{32'h429fb9de, 32'h41d34237, 32'hc22783c3, 32'hc2b3a829, 32'h40329aed, 32'h42b694a8, 32'h428dd1a2, 32'hc2120937};
test_output[4275] = '{32'h42b694a8};
test_index[4275] = '{5};
test_input[34208:34215] = '{32'hc1aba605, 32'hc2959eb2, 32'h429d5604, 32'hc1abea29, 32'h428b6314, 32'h42802cda, 32'h42c53f5c, 32'hc169ce00};
test_output[4276] = '{32'h42c53f5c};
test_index[4276] = '{6};
test_input[34216:34223] = '{32'hc1c3bb85, 32'hc295c050, 32'h4217c6b5, 32'hc26a6892, 32'hc20e4658, 32'h42b72410, 32'h423aa7f8, 32'h41119ce1};
test_output[4277] = '{32'h42b72410};
test_index[4277] = '{5};
test_input[34224:34231] = '{32'hc294719b, 32'hc2b1774f, 32'hc286858d, 32'h3ec4d054, 32'hc23441b4, 32'hc2b53bf3, 32'hc179034c, 32'hc109eba4};
test_output[4278] = '{32'h3ec4d054};
test_index[4278] = '{3};
test_input[34232:34239] = '{32'hc28ffc24, 32'h41a22f57, 32'hc1f1c172, 32'h410c8a44, 32'h420b15f6, 32'h41d1c711, 32'h424c8c6d, 32'h423a7c40};
test_output[4279] = '{32'h424c8c6d};
test_index[4279] = '{6};
test_input[34240:34247] = '{32'h42297397, 32'hc23f74e3, 32'hc27a57ad, 32'h4220bac1, 32'hc227b7f1, 32'hc2b109fb, 32'hc225c2a3, 32'hc1d672fa};
test_output[4280] = '{32'h42297397};
test_index[4280] = '{0};
test_input[34248:34255] = '{32'h42548b42, 32'hc220525a, 32'hc233a317, 32'h4271143d, 32'h426bf3bb, 32'hc204f634, 32'h425c57a1, 32'h4188a669};
test_output[4281] = '{32'h4271143d};
test_index[4281] = '{3};
test_input[34256:34263] = '{32'h4297b909, 32'hc2814f54, 32'h42b66b2f, 32'hc28e0c2d, 32'hc29c09d0, 32'hbf458b70, 32'hc0fbe881, 32'h42635777};
test_output[4282] = '{32'h42b66b2f};
test_index[4282] = '{2};
test_input[34264:34271] = '{32'h41f62a5b, 32'h42909ca2, 32'hc26dc370, 32'h422a834b, 32'h42434a21, 32'hc2757993, 32'hc26f2c90, 32'h42a190df};
test_output[4283] = '{32'h42a190df};
test_index[4283] = '{7};
test_input[34272:34279] = '{32'h428fa838, 32'hc0d003ea, 32'hc29d7afd, 32'h4297f887, 32'h427ad8d8, 32'hc1e4e3f9, 32'hc209fdfb, 32'hc273c62c};
test_output[4284] = '{32'h4297f887};
test_index[4284] = '{3};
test_input[34280:34287] = '{32'h4263310f, 32'h423a1264, 32'hc14bc9a0, 32'hc251caf7, 32'hc287d97c, 32'hc2742041, 32'h429711b0, 32'h4288a8d3};
test_output[4285] = '{32'h429711b0};
test_index[4285] = '{6};
test_input[34288:34295] = '{32'hc2881a7e, 32'hc24ad5d8, 32'h428455c8, 32'hc23954e6, 32'h417eb068, 32'hc19138f8, 32'h42c4a952, 32'hc2b956ed};
test_output[4286] = '{32'h42c4a952};
test_index[4286] = '{6};
test_input[34296:34303] = '{32'h4250d17c, 32'h42862697, 32'h4125ff87, 32'hc26bc495, 32'h42656ad8, 32'h41af7f90, 32'hc2978526, 32'hc13a1169};
test_output[4287] = '{32'h42862697};
test_index[4287] = '{1};
test_input[34304:34311] = '{32'h42a30b1a, 32'hc1a213d6, 32'h42ac6e7e, 32'h42a7972e, 32'hc20a5435, 32'h41b2d8e4, 32'hc1d0f0bf, 32'h42141b4e};
test_output[4288] = '{32'h42ac6e7e};
test_index[4288] = '{2};
test_input[34312:34319] = '{32'h42677a4c, 32'hc23690e4, 32'h42c27b11, 32'h421e4a3b, 32'hc2950aa5, 32'hc2bb04f1, 32'h4288bff8, 32'h40ee8b73};
test_output[4289] = '{32'h42c27b11};
test_index[4289] = '{2};
test_input[34320:34327] = '{32'h42441365, 32'h4289f8d4, 32'h40fe8223, 32'h426675b7, 32'h417d0500, 32'h4244fb8a, 32'h40d53958, 32'hc1b68898};
test_output[4290] = '{32'h4289f8d4};
test_index[4290] = '{1};
test_input[34328:34335] = '{32'hc28e872f, 32'h42aa2df3, 32'h42af26bd, 32'hc2bb217f, 32'h42af107e, 32'hc2867c3f, 32'h42755dd2, 32'h421875de};
test_output[4291] = '{32'h42af26bd};
test_index[4291] = '{2};
test_input[34336:34343] = '{32'hc12bf117, 32'h42b70695, 32'h4296aacd, 32'hc25a7ddd, 32'hc19eb16d, 32'h42a8afc6, 32'hbfd19af8, 32'hc1de77e7};
test_output[4292] = '{32'h42b70695};
test_index[4292] = '{1};
test_input[34344:34351] = '{32'hc1f2b8a7, 32'hc275152a, 32'hc228d9d3, 32'h417c4828, 32'h42addf10, 32'hc121650e, 32'hc2a723d3, 32'hc042da99};
test_output[4293] = '{32'h42addf10};
test_index[4293] = '{4};
test_input[34352:34359] = '{32'hc29989dd, 32'h42c1eeb3, 32'h3f13d173, 32'hc27f526f, 32'hc24e602f, 32'hc2b449bd, 32'hc2952311, 32'h42038114};
test_output[4294] = '{32'h42c1eeb3};
test_index[4294] = '{1};
test_input[34360:34367] = '{32'h40fa905d, 32'hc13780c0, 32'h41b496fc, 32'hc18f7c42, 32'hc22ae603, 32'h42b1e958, 32'h415dc524, 32'hc2af917f};
test_output[4295] = '{32'h42b1e958};
test_index[4295] = '{5};
test_input[34368:34375] = '{32'hc2a80657, 32'h4283fe8f, 32'h42afdd0d, 32'hc2b0efec, 32'h42709413, 32'h41c998a5, 32'h42bc33a7, 32'hc208d478};
test_output[4296] = '{32'h42bc33a7};
test_index[4296] = '{6};
test_input[34376:34383] = '{32'hc260b5fc, 32'h41f8d900, 32'h4284aa45, 32'hc2a3062f, 32'hc2556ff0, 32'hc2b9baa2, 32'hc26c6d47, 32'h41a73c1d};
test_output[4297] = '{32'h4284aa45};
test_index[4297] = '{2};
test_input[34384:34391] = '{32'h40d60426, 32'h42b19f15, 32'hc165fa06, 32'hc2b784bd, 32'h42840032, 32'h42a7e301, 32'h425b5d87, 32'h423250e2};
test_output[4298] = '{32'h42b19f15};
test_index[4298] = '{1};
test_input[34392:34399] = '{32'hc2bb701f, 32'hc2aa1521, 32'h421ce2ba, 32'hc21a2129, 32'hc209c2bf, 32'h42454614, 32'h4096fd87, 32'hc16e15f2};
test_output[4299] = '{32'h42454614};
test_index[4299] = '{5};
test_input[34400:34407] = '{32'h428aff23, 32'h422e3d57, 32'h428e2dc8, 32'hc28b69ae, 32'hc1e49d91, 32'h42a05c3e, 32'h421eb1ac, 32'h42b5beff};
test_output[4300] = '{32'h42b5beff};
test_index[4300] = '{7};
test_input[34408:34415] = '{32'hc2af4ecd, 32'hc1275e76, 32'hc2867c79, 32'hc219cbcf, 32'h42c4f8dd, 32'h42965ab7, 32'h410c1881, 32'h426c83b1};
test_output[4301] = '{32'h42c4f8dd};
test_index[4301] = '{4};
test_input[34416:34423] = '{32'h420bb2b5, 32'hc1f25b22, 32'hc2800ac7, 32'h41a011d1, 32'hc2c000d1, 32'hc20741e2, 32'h4252d5ce, 32'hc23f4220};
test_output[4302] = '{32'h4252d5ce};
test_index[4302] = '{6};
test_input[34424:34431] = '{32'hbfedb8a6, 32'hc0cf4807, 32'hc20f22e9, 32'h41bda9dd, 32'h42a8ba20, 32'hc29537c5, 32'h428b8b27, 32'hc236f3e7};
test_output[4303] = '{32'h42a8ba20};
test_index[4303] = '{4};
test_input[34432:34439] = '{32'h42bc1d50, 32'hc2baee7e, 32'h42795002, 32'hc2966da4, 32'h416d88dc, 32'hc23993ad, 32'h42657a50, 32'hc0cdb087};
test_output[4304] = '{32'h42bc1d50};
test_index[4304] = '{0};
test_input[34440:34447] = '{32'hc29aef56, 32'h42938488, 32'h42c7be2f, 32'hc277537e, 32'hc29b2319, 32'hc242a3bf, 32'h42c128a6, 32'h42b2bf9d};
test_output[4305] = '{32'h42c7be2f};
test_index[4305] = '{2};
test_input[34448:34455] = '{32'hc14c4fd4, 32'h42142810, 32'hc2003d18, 32'hc1c4bf3b, 32'h42a1beb0, 32'h42acd41d, 32'h41c82308, 32'hc2ab3acc};
test_output[4306] = '{32'h42acd41d};
test_index[4306] = '{5};
test_input[34456:34463] = '{32'hc10d3767, 32'h429910af, 32'hc1e136ed, 32'h4210e481, 32'h42c18511, 32'hc06d4bde, 32'hc2bdbf13, 32'hc21e45da};
test_output[4307] = '{32'h42c18511};
test_index[4307] = '{4};
test_input[34464:34471] = '{32'hc24849a1, 32'h426c5f1f, 32'hc0cd78a4, 32'h3e7c1974, 32'h429fde12, 32'hc20a70c4, 32'hc13e3cd3, 32'hc1ec7ed7};
test_output[4308] = '{32'h429fde12};
test_index[4308] = '{4};
test_input[34472:34479] = '{32'hc2701e1f, 32'h419e55db, 32'h427a8a2d, 32'h408a7cd4, 32'hc2c22b5d, 32'h4239bab0, 32'hc2c7fbba, 32'hc21f9b5f};
test_output[4309] = '{32'h427a8a2d};
test_index[4309] = '{2};
test_input[34480:34487] = '{32'h4280f10d, 32'hc28c2ed6, 32'hc1238e9e, 32'hc2801882, 32'h428990fa, 32'hc15b177e, 32'hc0b88743, 32'hc2a00873};
test_output[4310] = '{32'h428990fa};
test_index[4310] = '{4};
test_input[34488:34495] = '{32'hc2aa9199, 32'h40bee73c, 32'h4217fc87, 32'hc292cd1b, 32'h421c2e72, 32'hc25182d5, 32'hc21bd057, 32'h41668354};
test_output[4311] = '{32'h421c2e72};
test_index[4311] = '{4};
test_input[34496:34503] = '{32'hc1f374a2, 32'h41d06423, 32'h423b8f7b, 32'hc1e35740, 32'h41ef0c7e, 32'h4199bd56, 32'hc282fe12, 32'hc2807b22};
test_output[4312] = '{32'h423b8f7b};
test_index[4312] = '{2};
test_input[34504:34511] = '{32'hc2a48902, 32'hc29dcb85, 32'hc2312f53, 32'hc1a104d0, 32'h42987fb0, 32'h41085ab6, 32'h428a76d1, 32'h4024a2ae};
test_output[4313] = '{32'h42987fb0};
test_index[4313] = '{4};
test_input[34512:34519] = '{32'hc0ee2f2f, 32'hc2233661, 32'h415f5a1c, 32'hc20b0323, 32'h42818228, 32'hc2905dee, 32'hc1fc1a04, 32'hc180751b};
test_output[4314] = '{32'h42818228};
test_index[4314] = '{4};
test_input[34520:34527] = '{32'h424de1c5, 32'h41908dc4, 32'hc293bfd4, 32'h42092e14, 32'hc1fc34de, 32'hc265b94e, 32'h42ac6dc4, 32'hc2a11c33};
test_output[4315] = '{32'h42ac6dc4};
test_index[4315] = '{6};
test_input[34528:34535] = '{32'h421480a5, 32'h42136e59, 32'h4296f032, 32'hc2abb1bf, 32'h42a06365, 32'hc2a3e721, 32'h42b5cd3d, 32'hc2923fcb};
test_output[4316] = '{32'h42b5cd3d};
test_index[4316] = '{6};
test_input[34536:34543] = '{32'hc12b9ef5, 32'h4266cec8, 32'h42685131, 32'h42817ed8, 32'hc1877ad9, 32'h4021c7da, 32'h42012e83, 32'hc2bf304d};
test_output[4317] = '{32'h42817ed8};
test_index[4317] = '{3};
test_input[34544:34551] = '{32'h41d46cfe, 32'hc2b24ba7, 32'hc2a7b7ef, 32'h429fc7ed, 32'hc217cc07, 32'h42958517, 32'hc140d621, 32'h4287540c};
test_output[4318] = '{32'h429fc7ed};
test_index[4318] = '{3};
test_input[34552:34559] = '{32'hc27b9436, 32'h42a49f38, 32'h411272fa, 32'h42262034, 32'hc202b1af, 32'hc279d326, 32'hc138644c, 32'hc22df0c8};
test_output[4319] = '{32'h42a49f38};
test_index[4319] = '{1};
test_input[34560:34567] = '{32'hc200021b, 32'h3feae63b, 32'hc27aa19b, 32'hc170e750, 32'hc25e6005, 32'h423c8b60, 32'hc042a694, 32'h42be1c16};
test_output[4320] = '{32'h42be1c16};
test_index[4320] = '{7};
test_input[34568:34575] = '{32'h428167d7, 32'hc28c2e4e, 32'h42a877bb, 32'hc2abd111, 32'hc25dda12, 32'h40365df7, 32'h3f60491f, 32'hc29abd96};
test_output[4321] = '{32'h42a877bb};
test_index[4321] = '{2};
test_input[34576:34583] = '{32'h42999486, 32'hc20e0034, 32'h4281e85c, 32'h41a4e504, 32'h425fc054, 32'h427fcb1d, 32'h40fc25d5, 32'hc2248501};
test_output[4322] = '{32'h42999486};
test_index[4322] = '{0};
test_input[34584:34591] = '{32'hc29da120, 32'hc267d37c, 32'h4253ff7a, 32'h41b13a07, 32'h42340c89, 32'h4201973e, 32'h428f1215, 32'hc28de1c7};
test_output[4323] = '{32'h428f1215};
test_index[4323] = '{6};
test_input[34592:34599] = '{32'h42964cb8, 32'hc26e316b, 32'h425c7223, 32'hc2674484, 32'h429f1a9d, 32'h429c1a12, 32'hc25cfd9e, 32'h41874e72};
test_output[4324] = '{32'h429f1a9d};
test_index[4324] = '{4};
test_input[34600:34607] = '{32'hc2b32794, 32'hc18da531, 32'hc2a9f0a8, 32'hc24fd72e, 32'h42859a62, 32'hc21a7cee, 32'hc2992416, 32'h4241802d};
test_output[4325] = '{32'h42859a62};
test_index[4325] = '{4};
test_input[34608:34615] = '{32'h42b58b91, 32'h42b036e0, 32'h42525ec2, 32'h41a7b2b9, 32'h424ff103, 32'hc28c3f76, 32'h401b4f6f, 32'hc29fb1e9};
test_output[4326] = '{32'h42b58b91};
test_index[4326] = '{0};
test_input[34616:34623] = '{32'h3feace89, 32'hc1783bc3, 32'hc1ea965c, 32'h42b403e5, 32'hc2c408eb, 32'hc299d5ba, 32'hc24d7e9f, 32'hc1b2c963};
test_output[4327] = '{32'h42b403e5};
test_index[4327] = '{3};
test_input[34624:34631] = '{32'h410689c4, 32'hc295159d, 32'h429d7efa, 32'hc2b5f457, 32'hc1d59d6b, 32'hc1dee1c3, 32'hc08a4537, 32'h4096116a};
test_output[4328] = '{32'h429d7efa};
test_index[4328] = '{2};
test_input[34632:34639] = '{32'hc1d84c86, 32'hc17280ac, 32'h426e3e69, 32'h42bb9d6e, 32'hc1bb3d14, 32'h426cffae, 32'hc17df31d, 32'h42838321};
test_output[4329] = '{32'h42bb9d6e};
test_index[4329] = '{3};
test_input[34640:34647] = '{32'hc264c50d, 32'hc2895f80, 32'hc28eb0ad, 32'h42bac448, 32'h418ce7c1, 32'h42868319, 32'hc1be2893, 32'h42b3e2ff};
test_output[4330] = '{32'h42bac448};
test_index[4330] = '{3};
test_input[34648:34655] = '{32'h42b77092, 32'h41273994, 32'hc23930d6, 32'h42b1bdaf, 32'h42119435, 32'hc2b55068, 32'hc295221a, 32'h428f32d0};
test_output[4331] = '{32'h42b77092};
test_index[4331] = '{0};
test_input[34656:34663] = '{32'hc2a650ed, 32'hc21095e2, 32'hc1150b6b, 32'h428ac100, 32'h41df1d61, 32'hc284ec89, 32'hc2456f8f, 32'h42bd62ef};
test_output[4332] = '{32'h42bd62ef};
test_index[4332] = '{7};
test_input[34664:34671] = '{32'hc29cb01e, 32'h4282bd64, 32'hc2498f8b, 32'h41e98f43, 32'h41980b49, 32'h418e8995, 32'h42b7b2cb, 32'h42abbb73};
test_output[4333] = '{32'h42b7b2cb};
test_index[4333] = '{6};
test_input[34672:34679] = '{32'h416a5c76, 32'h418b751c, 32'hc284ec29, 32'hc2c2be43, 32'h4291cc1d, 32'hc118de96, 32'h42c6ec9c, 32'hc29056d2};
test_output[4334] = '{32'h42c6ec9c};
test_index[4334] = '{6};
test_input[34680:34687] = '{32'hc2542dd9, 32'hc2c24ed2, 32'hc2c71303, 32'hc01ae6c3, 32'hc266b00d, 32'h4116e9ea, 32'h42a061bb, 32'hc039cabb};
test_output[4335] = '{32'h42a061bb};
test_index[4335] = '{6};
test_input[34688:34695] = '{32'hc15b9952, 32'h42642922, 32'hc2001213, 32'hc2badc10, 32'hc1c883f0, 32'hc1d7ff41, 32'h428a58da, 32'hc1bb004e};
test_output[4336] = '{32'h428a58da};
test_index[4336] = '{6};
test_input[34696:34703] = '{32'hc28b854b, 32'hc20b0afc, 32'h408abeff, 32'hc2c24021, 32'h427183cb, 32'hc27493df, 32'hc16232a7, 32'h41b22fe6};
test_output[4337] = '{32'h427183cb};
test_index[4337] = '{4};
test_input[34704:34711] = '{32'h4284b6a1, 32'hc225d3be, 32'hc10d21fd, 32'h4214c8d9, 32'h42887334, 32'h42afee8f, 32'hc1db145a, 32'h422c4610};
test_output[4338] = '{32'h42afee8f};
test_index[4338] = '{5};
test_input[34712:34719] = '{32'hbfdff7a1, 32'hc2530f1d, 32'hc1e05ca3, 32'hc2652850, 32'h42c57552, 32'hc260517e, 32'hc29c28ae, 32'h409be097};
test_output[4339] = '{32'h42c57552};
test_index[4339] = '{4};
test_input[34720:34727] = '{32'h42a3449f, 32'h422b1cec, 32'h41f13de9, 32'hc2ad19f8, 32'hc2b401ce, 32'h42668636, 32'h42c4ad65, 32'hc0a11db1};
test_output[4340] = '{32'h42c4ad65};
test_index[4340] = '{6};
test_input[34728:34735] = '{32'hc194c290, 32'hc2a36a98, 32'h41907910, 32'hc28da13a, 32'h4219e64b, 32'h3e1a58f1, 32'hc22e9f6a, 32'hc1f6463e};
test_output[4341] = '{32'h4219e64b};
test_index[4341] = '{4};
test_input[34736:34743] = '{32'hc26ea14f, 32'hc2b20995, 32'hc23c5ce9, 32'h3fa64bdc, 32'hc14e2bf1, 32'hc2b21832, 32'h422a7c07, 32'h41cb1248};
test_output[4342] = '{32'h422a7c07};
test_index[4342] = '{6};
test_input[34744:34751] = '{32'hc2210547, 32'h40fa5c0c, 32'h424fc38f, 32'h42b35037, 32'hc0a63eb2, 32'hc2344ba0, 32'h421268e9, 32'hc2894ed3};
test_output[4343] = '{32'h42b35037};
test_index[4343] = '{3};
test_input[34752:34759] = '{32'h42404384, 32'hc29292ca, 32'h4196d801, 32'hc29e38cb, 32'h42511d3c, 32'hc2930527, 32'h420820f0, 32'h424805a5};
test_output[4344] = '{32'h42511d3c};
test_index[4344] = '{4};
test_input[34760:34767] = '{32'hc15adfa8, 32'h41c10f95, 32'hc1a104e3, 32'hc2a74aff, 32'h415abf6f, 32'hc2129fc3, 32'h42c33dd4, 32'hc2c432cd};
test_output[4345] = '{32'h42c33dd4};
test_index[4345] = '{6};
test_input[34768:34775] = '{32'h429f629c, 32'h42331813, 32'hc2c5e8d4, 32'h429ba0f4, 32'h3ff9dc19, 32'hc284ef14, 32'hc2a12b1f, 32'hc286e60c};
test_output[4346] = '{32'h429f629c};
test_index[4346] = '{0};
test_input[34776:34783] = '{32'h42b61319, 32'h412b7e01, 32'h3d311a50, 32'h429a9c5a, 32'h427bd52e, 32'h42336810, 32'h41800c4d, 32'h4282bcaf};
test_output[4347] = '{32'h42b61319};
test_index[4347] = '{0};
test_input[34784:34791] = '{32'hc131ce9c, 32'hc28c9233, 32'hc17db1b3, 32'hc2bbe159, 32'hc20a7db8, 32'h4219b4c4, 32'h42a1231f, 32'hbea79768};
test_output[4348] = '{32'h42a1231f};
test_index[4348] = '{6};
test_input[34792:34799] = '{32'h42a8a420, 32'h42b047d3, 32'hc207a35e, 32'hc262e76b, 32'hc2c4cbea, 32'h3fbe1cc8, 32'hc2975c45, 32'h3e3ef905};
test_output[4349] = '{32'h42b047d3};
test_index[4349] = '{1};
test_input[34800:34807] = '{32'hc2a204b4, 32'hc28094fe, 32'hc2b72fe5, 32'hc142ced4, 32'hc09505b3, 32'hc2c01463, 32'hc2b59826, 32'hc28d0a23};
test_output[4350] = '{32'hc09505b3};
test_index[4350] = '{4};
test_input[34808:34815] = '{32'hc2b0c720, 32'hc271aaee, 32'h428dcebe, 32'h419d1f25, 32'hc2627b69, 32'hc2727d75, 32'hc2024982, 32'h42bcf4f1};
test_output[4351] = '{32'h42bcf4f1};
test_index[4351] = '{7};
test_input[34816:34823] = '{32'hc17aa1d8, 32'h4186471b, 32'h41d540d0, 32'h41d02b54, 32'h425dc860, 32'hc287ff64, 32'hc232d29e, 32'h413fbf1c};
test_output[4352] = '{32'h425dc860};
test_index[4352] = '{4};
test_input[34824:34831] = '{32'hc241214f, 32'h4225991f, 32'h4233f918, 32'h42be28bb, 32'h41099718, 32'h4272a711, 32'hc1c1a82f, 32'h41e620ff};
test_output[4353] = '{32'h42be28bb};
test_index[4353] = '{3};
test_input[34832:34839] = '{32'hc2557da1, 32'hc2b49903, 32'hc260bb75, 32'hc1d9cc96, 32'h423d4388, 32'hc061fee6, 32'h40e82148, 32'hc2449415};
test_output[4354] = '{32'h423d4388};
test_index[4354] = '{4};
test_input[34840:34847] = '{32'h424a0af0, 32'hc2afd0b7, 32'hc25f2bae, 32'h4006d013, 32'h41ab9165, 32'h4190ee2c, 32'h4293b913, 32'hc2009b65};
test_output[4355] = '{32'h4293b913};
test_index[4355] = '{6};
test_input[34848:34855] = '{32'hc22e0763, 32'hc28f6369, 32'hc296cc21, 32'hc2718c2f, 32'h41e3c276, 32'hc0b476e6, 32'h42949110, 32'h42c5a890};
test_output[4356] = '{32'h42c5a890};
test_index[4356] = '{7};
test_input[34856:34863] = '{32'hc28ceda2, 32'hc2bacd44, 32'h4251e472, 32'h423c4226, 32'h428585a2, 32'hc2c05faf, 32'h42751150, 32'hc19027d4};
test_output[4357] = '{32'h428585a2};
test_index[4357] = '{4};
test_input[34864:34871] = '{32'hc2a7e9b3, 32'hc2672011, 32'hc2060a6a, 32'hc242d87a, 32'hc29a575b, 32'hc1f4d14d, 32'hc293cb3f, 32'h42bc01dd};
test_output[4358] = '{32'h42bc01dd};
test_index[4358] = '{7};
test_input[34872:34879] = '{32'hc2744c97, 32'hc296e3f1, 32'hc26986b3, 32'h40a015be, 32'hc287b743, 32'h4216a032, 32'hc2044762, 32'hbf768559};
test_output[4359] = '{32'h4216a032};
test_index[4359] = '{5};
test_input[34880:34887] = '{32'hc1849b26, 32'hc1ea2759, 32'hc28324a8, 32'h42a394fd, 32'hc2943cc4, 32'hc23ce1c8, 32'h42803de0, 32'hc281802f};
test_output[4360] = '{32'h42a394fd};
test_index[4360] = '{3};
test_input[34888:34895] = '{32'hc230558f, 32'hc1c1744f, 32'hc1988f4b, 32'hc2804e3d, 32'hc294ea50, 32'hc1c15ef6, 32'hc2832114, 32'h4224e255};
test_output[4361] = '{32'h4224e255};
test_index[4361] = '{7};
test_input[34896:34903] = '{32'hc2a8f43e, 32'h41f1ce73, 32'h41890bdf, 32'hc286816e, 32'hc007360e, 32'hc2c7a298, 32'h424e52aa, 32'h41107fdd};
test_output[4362] = '{32'h424e52aa};
test_index[4362] = '{6};
test_input[34904:34911] = '{32'h42ad3ff5, 32'hc2b550c5, 32'hc2c44268, 32'hc23c52c5, 32'h424cf47e, 32'h4291a0a4, 32'hc1589d2b, 32'hc146c521};
test_output[4363] = '{32'h42ad3ff5};
test_index[4363] = '{0};
test_input[34912:34919] = '{32'h42c002c0, 32'hc2903fdb, 32'hc29fe3fd, 32'hc161f8b5, 32'h427e5b14, 32'h41422207, 32'h4292c36a, 32'h4173aaff};
test_output[4364] = '{32'h42c002c0};
test_index[4364] = '{0};
test_input[34920:34927] = '{32'hc297a119, 32'hc2b240b4, 32'h417887e4, 32'hbeea4b2e, 32'hc0d3be03, 32'hc2b3bf20, 32'hc2456453, 32'hc13e1825};
test_output[4365] = '{32'h417887e4};
test_index[4365] = '{2};
test_input[34928:34935] = '{32'h42809154, 32'hc28fe609, 32'hc26e41dd, 32'hc295549c, 32'h4103fb08, 32'hc2a860ce, 32'hc1a1e88a, 32'h3ff96e81};
test_output[4366] = '{32'h42809154};
test_index[4366] = '{0};
test_input[34936:34943] = '{32'h429d8d1a, 32'hc2c13ed0, 32'hc200230a, 32'h416c8dc3, 32'h42c5052e, 32'hc2113b29, 32'h40b8a2f0, 32'hc2a0859d};
test_output[4367] = '{32'h42c5052e};
test_index[4367] = '{4};
test_input[34944:34951] = '{32'hc2863f82, 32'h40e7cc53, 32'hc2af8259, 32'hc28cccca, 32'h42ad53c4, 32'h42871891, 32'hc2a72f8a, 32'hc2b71a61};
test_output[4368] = '{32'h42ad53c4};
test_index[4368] = '{4};
test_input[34952:34959] = '{32'h4288f1ef, 32'hc1e41988, 32'hc116ad36, 32'hc29aa25f, 32'h41103455, 32'h4171efd1, 32'hc117075e, 32'hc276b158};
test_output[4369] = '{32'h4288f1ef};
test_index[4369] = '{0};
test_input[34960:34967] = '{32'h42058bc1, 32'h424101a4, 32'hc2598e78, 32'h42a0b4f4, 32'hc15c988f, 32'h3f4ae881, 32'h42446f9b, 32'h42862df6};
test_output[4370] = '{32'h42a0b4f4};
test_index[4370] = '{3};
test_input[34968:34975] = '{32'hc1b81022, 32'hc26d126a, 32'hc2849b13, 32'hc2ae7969, 32'h407c64e0, 32'h42b3a031, 32'hc285b78c, 32'hc22e64de};
test_output[4371] = '{32'h42b3a031};
test_index[4371] = '{5};
test_input[34976:34983] = '{32'hc207a1b3, 32'h42bb00dc, 32'h4230a213, 32'hc2904926, 32'h429bfc46, 32'hc0ac2cb1, 32'hc256cb2c, 32'h400b15e5};
test_output[4372] = '{32'h42bb00dc};
test_index[4372] = '{1};
test_input[34984:34991] = '{32'h41b92db9, 32'h41bf9a21, 32'h42bbf442, 32'hc18be296, 32'h42014059, 32'h423eb330, 32'hc10170d2, 32'hc241e71f};
test_output[4373] = '{32'h42bbf442};
test_index[4373] = '{2};
test_input[34992:34999] = '{32'hc1d05995, 32'h41ad07ef, 32'hc2a8b927, 32'hc22622e3, 32'hc1b2197e, 32'h428d2fde, 32'hc2624b81, 32'hc2850b62};
test_output[4374] = '{32'h428d2fde};
test_index[4374] = '{5};
test_input[35000:35007] = '{32'h41f7b368, 32'hc20e03fb, 32'h41b6eff5, 32'hc2c74f20, 32'hc2a3378d, 32'hc1946738, 32'h41ae3b86, 32'h42448d4a};
test_output[4375] = '{32'h42448d4a};
test_index[4375] = '{7};
test_input[35008:35015] = '{32'h42ad38d5, 32'h427d2b10, 32'hc217a670, 32'h428415ef, 32'hc20aca7c, 32'h4264d9e7, 32'h41b72a34, 32'hc2b2edcb};
test_output[4376] = '{32'h42ad38d5};
test_index[4376] = '{0};
test_input[35016:35023] = '{32'hc2a1061d, 32'h42a2e949, 32'h40497f58, 32'h4294507a, 32'h40d74879, 32'h42a8d0b5, 32'h42a4849d, 32'h41b380c5};
test_output[4377] = '{32'h42a8d0b5};
test_index[4377] = '{5};
test_input[35024:35031] = '{32'h420b8971, 32'h415a6d08, 32'h4201fb9e, 32'hc288a38d, 32'h428cb201, 32'hc2320fb3, 32'hc06af2be, 32'h40011d19};
test_output[4378] = '{32'h428cb201};
test_index[4378] = '{4};
test_input[35032:35039] = '{32'hc1f0a1ad, 32'h42900f66, 32'hc0090cb5, 32'h423b22e9, 32'h42c7b025, 32'h42c2fcfe, 32'h41ea1e0a, 32'hc207a40e};
test_output[4379] = '{32'h42c7b025};
test_index[4379] = '{4};
test_input[35040:35047] = '{32'hc2a4c952, 32'h41d370fb, 32'hc28c1872, 32'hc277ebca, 32'hc27965e1, 32'hc1eb1311, 32'hc229f0ba, 32'hc2a4f931};
test_output[4380] = '{32'h41d370fb};
test_index[4380] = '{1};
test_input[35048:35055] = '{32'hc2424b3b, 32'h428378a2, 32'hc2095226, 32'h4298f9aa, 32'h42753a48, 32'h42be3973, 32'h427727e2, 32'h418d711c};
test_output[4381] = '{32'h42be3973};
test_index[4381] = '{5};
test_input[35056:35063] = '{32'hc097b075, 32'h42167f75, 32'hc1f1d539, 32'h42875561, 32'h42c0cd72, 32'hc17a991e, 32'h3f8e73ff, 32'h41e43539};
test_output[4382] = '{32'h42c0cd72};
test_index[4382] = '{4};
test_input[35064:35071] = '{32'h42a7251d, 32'h42632994, 32'h42bf566c, 32'h41cb3a99, 32'h40234cd6, 32'hc135905a, 32'hc288f5ef, 32'h429d96f9};
test_output[4383] = '{32'h42bf566c};
test_index[4383] = '{2};
test_input[35072:35079] = '{32'h422d1dd1, 32'hc27c2706, 32'h4294bb4f, 32'hc0808ea6, 32'hc18b4e3b, 32'h42855d84, 32'h42a89f0c, 32'h3fa885d1};
test_output[4384] = '{32'h42a89f0c};
test_index[4384] = '{6};
test_input[35080:35087] = '{32'h42b25d32, 32'hc257caf1, 32'h42209de8, 32'hc286bae1, 32'h407f6fa0, 32'h423e7de8, 32'hc1fd11ed, 32'h41be8b5b};
test_output[4385] = '{32'h42b25d32};
test_index[4385] = '{0};
test_input[35088:35095] = '{32'hc109143e, 32'h42ab3178, 32'hc2a7f8ab, 32'hc20f26c5, 32'h4281822f, 32'h42851844, 32'h4187656b, 32'h4277b1ce};
test_output[4386] = '{32'h42ab3178};
test_index[4386] = '{1};
test_input[35096:35103] = '{32'h425fefd2, 32'hbfbc3532, 32'hc26c50f1, 32'h4236ed67, 32'h422b2bae, 32'h4197f942, 32'h429a6130, 32'h42341507};
test_output[4387] = '{32'h429a6130};
test_index[4387] = '{6};
test_input[35104:35111] = '{32'h4297d1c4, 32'h4294426a, 32'h41e7571f, 32'h40a25da6, 32'hc2211a9f, 32'hc2918f58, 32'hbe7945ee, 32'h40f6109b};
test_output[4388] = '{32'h4297d1c4};
test_index[4388] = '{0};
test_input[35112:35119] = '{32'h42afcc6b, 32'h41cc456d, 32'h42aea33b, 32'hc123e5ac, 32'hc02844da, 32'hc261c89b, 32'h429031fc, 32'h41a90b41};
test_output[4389] = '{32'h42afcc6b};
test_index[4389] = '{0};
test_input[35120:35127] = '{32'h42afb427, 32'h42921e53, 32'hc22d8dfb, 32'h3fafa2ed, 32'h40e2743a, 32'h42a38d6d, 32'hc175c40e, 32'h41c7887c};
test_output[4390] = '{32'h42afb427};
test_index[4390] = '{0};
test_input[35128:35135] = '{32'h429a6c7b, 32'hc29147c4, 32'h416c1bb5, 32'hc29704b6, 32'h40b8d947, 32'h42b2cb3d, 32'hc0b183e9, 32'h3f8c75ff};
test_output[4391] = '{32'h42b2cb3d};
test_index[4391] = '{5};
test_input[35136:35143] = '{32'h41675aa8, 32'hc2bb3788, 32'h4294dea2, 32'h419e126a, 32'hc21d4d51, 32'hc0192151, 32'hc268a41f, 32'hc1aabd32};
test_output[4392] = '{32'h4294dea2};
test_index[4392] = '{2};
test_input[35144:35151] = '{32'hc1d50f9a, 32'h42287cea, 32'h42ac7339, 32'hc2c23fde, 32'hc1334be1, 32'h41b863db, 32'h4211e2e7, 32'hc1e17c5f};
test_output[4393] = '{32'h42ac7339};
test_index[4393] = '{2};
test_input[35152:35159] = '{32'hc249e7ba, 32'h3fc82baa, 32'h42aef98a, 32'hc22efa1e, 32'hbfe377d9, 32'hc25eeb8d, 32'hc23e43bb, 32'h42a5615e};
test_output[4394] = '{32'h42aef98a};
test_index[4394] = '{2};
test_input[35160:35167] = '{32'hc2322943, 32'h422714f3, 32'h40decb76, 32'hbf8eca2f, 32'hc2c0308d, 32'hc25432a9, 32'h41a7e021, 32'h427069ce};
test_output[4395] = '{32'h427069ce};
test_index[4395] = '{7};
test_input[35168:35175] = '{32'hc29b78e4, 32'hc227fd63, 32'h42082527, 32'hc105ffc6, 32'h4155fe71, 32'hc0e38b69, 32'h428cc0bb, 32'hc21cc07c};
test_output[4396] = '{32'h428cc0bb};
test_index[4396] = '{6};
test_input[35176:35183] = '{32'h42325b2b, 32'hc0065cb2, 32'hc1e87a3a, 32'hc2bc0c9b, 32'h4280c513, 32'h41a47bc8, 32'hc217f22b, 32'h42978e02};
test_output[4397] = '{32'h42978e02};
test_index[4397] = '{7};
test_input[35184:35191] = '{32'hc2b27616, 32'h422c9ea1, 32'h421b513f, 32'hc0d53847, 32'hc26f0fc9, 32'h419c3cc8, 32'hc17ab5ef, 32'h424cc5c9};
test_output[4398] = '{32'h424cc5c9};
test_index[4398] = '{7};
test_input[35192:35199] = '{32'hc2a5a58a, 32'h42bb7c71, 32'h422a4a03, 32'h41c8af4b, 32'hc251d954, 32'h41823755, 32'h42be4133, 32'h42c1c68b};
test_output[4399] = '{32'h42c1c68b};
test_index[4399] = '{7};
test_input[35200:35207] = '{32'hc2bd89c1, 32'h4223e97e, 32'hc1ebf68a, 32'hc229cb39, 32'hc1c8fef9, 32'hc04b664d, 32'h4280f89d, 32'h4215a90d};
test_output[4400] = '{32'h4280f89d};
test_index[4400] = '{6};
test_input[35208:35215] = '{32'hc2003348, 32'h423d7b5c, 32'hbe5deb97, 32'hc213837f, 32'h42a192fd, 32'h428741c9, 32'hc282a281, 32'h4213a827};
test_output[4401] = '{32'h42a192fd};
test_index[4401] = '{4};
test_input[35216:35223] = '{32'h425fa068, 32'hc240864a, 32'h41829ff0, 32'h42c511ea, 32'hc2a3cd2e, 32'hc0b4cb6b, 32'h42c370a7, 32'h426b618a};
test_output[4402] = '{32'h42c511ea};
test_index[4402] = '{3};
test_input[35224:35231] = '{32'h420a5564, 32'hc16a0bb9, 32'hc16d7f5f, 32'hc2c31109, 32'hc12cf25b, 32'hc13f5541, 32'hc290418e, 32'h41939e0d};
test_output[4403] = '{32'h420a5564};
test_index[4403] = '{0};
test_input[35232:35239] = '{32'hc06f2f84, 32'h428d9f0b, 32'hbf9d19be, 32'h41746705, 32'h4238293b, 32'h4248d20b, 32'hc2be3973, 32'hc1d78463};
test_output[4404] = '{32'h428d9f0b};
test_index[4404] = '{1};
test_input[35240:35247] = '{32'hc24d117f, 32'h424e9512, 32'h42386a82, 32'h42c79692, 32'h429884f0, 32'hc28af06d, 32'hc1478e8a, 32'h413e8bbf};
test_output[4405] = '{32'h42c79692};
test_index[4405] = '{3};
test_input[35248:35255] = '{32'hc22d7ac2, 32'hc1fc0f64, 32'h40c32518, 32'hc1cc9c57, 32'h42b37ab4, 32'h40451c2b, 32'hbfb6ee9c, 32'h4194e785};
test_output[4406] = '{32'h42b37ab4};
test_index[4406] = '{4};
test_input[35256:35263] = '{32'h42ab5b23, 32'hc2ac46de, 32'hc284b1bf, 32'hc18c79d0, 32'h417bed2d, 32'h42c0e01d, 32'h42845ce2, 32'h428ceebf};
test_output[4407] = '{32'h42c0e01d};
test_index[4407] = '{5};
test_input[35264:35271] = '{32'h416b2048, 32'h4255af24, 32'h426ca620, 32'h427cd2cf, 32'h4205611e, 32'hc11132dd, 32'h41acb662, 32'hc2c37784};
test_output[4408] = '{32'h427cd2cf};
test_index[4408] = '{3};
test_input[35272:35279] = '{32'hc17b274b, 32'h41ac84c3, 32'h4279c2bd, 32'h41e1d278, 32'hc2acd9bb, 32'h411b603b, 32'hc2bba2d8, 32'hc22b4853};
test_output[4409] = '{32'h4279c2bd};
test_index[4409] = '{2};
test_input[35280:35287] = '{32'hc2a13890, 32'h3f287bc6, 32'h42a7242f, 32'h425acc75, 32'hc200b209, 32'h42ae73b2, 32'hc11bae2c, 32'hc2b56021};
test_output[4410] = '{32'h42ae73b2};
test_index[4410] = '{5};
test_input[35288:35295] = '{32'h422ccbdc, 32'h411fdc64, 32'h41b92a0b, 32'hc1549527, 32'h42338116, 32'hc2997a15, 32'hc2559dbf, 32'hc2863739};
test_output[4411] = '{32'h42338116};
test_index[4411] = '{4};
test_input[35296:35303] = '{32'hc2867ba3, 32'h419d2f20, 32'hc28ce7ee, 32'h4268cf02, 32'hc1cb3c4c, 32'hc19ef4c2, 32'hc28649fc, 32'hc2732439};
test_output[4412] = '{32'h4268cf02};
test_index[4412] = '{3};
test_input[35304:35311] = '{32'hc234808b, 32'h42a9fc90, 32'hc2940e07, 32'hc2bd48ec, 32'h422954d1, 32'h42a34d96, 32'h421d74e6, 32'hc2a7e219};
test_output[4413] = '{32'h42a9fc90};
test_index[4413] = '{1};
test_input[35312:35319] = '{32'hc242d6ce, 32'hc286a9c6, 32'h42854c5f, 32'h42b745a9, 32'h42b7cb28, 32'h4223e45b, 32'h41cf5bda, 32'h42b283ad};
test_output[4414] = '{32'h42b7cb28};
test_index[4414] = '{4};
test_input[35320:35327] = '{32'h429dd0d5, 32'h42aa3e5b, 32'h422aef63, 32'h42692923, 32'hc0ad8fa1, 32'h41bdf139, 32'hc0155527, 32'h42b6d9b2};
test_output[4415] = '{32'h42b6d9b2};
test_index[4415] = '{7};
test_input[35328:35335] = '{32'h4275a46c, 32'h41132c96, 32'hc299860e, 32'hbdf18e0b, 32'hc2aefac0, 32'h428d28e5, 32'hc1079617, 32'hc2331898};
test_output[4416] = '{32'h428d28e5};
test_index[4416] = '{5};
test_input[35336:35343] = '{32'hc28c2a7a, 32'h42b03587, 32'hc2b66725, 32'h428cb03b, 32'h41a4328b, 32'h41cb1d16, 32'h41978f12, 32'hc206c211};
test_output[4417] = '{32'h42b03587};
test_index[4417] = '{1};
test_input[35344:35351] = '{32'h4255baf6, 32'h40561993, 32'hc1e59f48, 32'h42c03f32, 32'hc1b31fbf, 32'hc1c982bb, 32'h410fe50d, 32'h429c8610};
test_output[4418] = '{32'h42c03f32};
test_index[4418] = '{3};
test_input[35352:35359] = '{32'hc0c84d21, 32'hc240c8e8, 32'h41318084, 32'h4176000d, 32'hc2487bd9, 32'hc22dfcae, 32'h40e945e3, 32'hc1800eee};
test_output[4419] = '{32'h4176000d};
test_index[4419] = '{3};
test_input[35360:35367] = '{32'hc237eedd, 32'h41b96a5e, 32'hc25191f3, 32'hc252be2f, 32'hc2b1dcc8, 32'h420a3a25, 32'hc2adfeb2, 32'hc132a294};
test_output[4420] = '{32'h420a3a25};
test_index[4420] = '{5};
test_input[35368:35375] = '{32'hc21af301, 32'h41402ee2, 32'hc2c203b6, 32'h4285d9bf, 32'hc1cbf96f, 32'h42a41cee, 32'hc24af3d8, 32'h4177b654};
test_output[4421] = '{32'h42a41cee};
test_index[4421] = '{5};
test_input[35376:35383] = '{32'hc23daba3, 32'hc256cd87, 32'h42c0000f, 32'hc2134712, 32'hc28f1009, 32'h4292e061, 32'hc1bb9230, 32'hc26692d4};
test_output[4422] = '{32'h42c0000f};
test_index[4422] = '{2};
test_input[35384:35391] = '{32'hc117f971, 32'h4279266b, 32'hc1b387c1, 32'hc25e2ef7, 32'h40e549dc, 32'h40a60e05, 32'hc1c62fb7, 32'hc2420ecc};
test_output[4423] = '{32'h4279266b};
test_index[4423] = '{1};
test_input[35392:35399] = '{32'h41cacad8, 32'h40ca5917, 32'h41282916, 32'hc10118b0, 32'h4102333b, 32'h42b63ae4, 32'hc2373e7b, 32'hc22050ec};
test_output[4424] = '{32'h42b63ae4};
test_index[4424] = '{5};
test_input[35400:35407] = '{32'hc29a2d29, 32'hc2b70f7f, 32'h427ab0f2, 32'hc2b108e9, 32'h40b3e880, 32'h42479fbe, 32'h4102f8b2, 32'h42afc487};
test_output[4425] = '{32'h42afc487};
test_index[4425] = '{7};
test_input[35408:35415] = '{32'h427dd972, 32'h42adcbbd, 32'hc101ccd2, 32'h428d11fb, 32'h429b55d4, 32'hc2ac31fb, 32'hc2090e8d, 32'h4278317b};
test_output[4426] = '{32'h42adcbbd};
test_index[4426] = '{1};
test_input[35416:35423] = '{32'hc276f9cb, 32'hc13ac9f4, 32'hc2282e88, 32'h423763a4, 32'hc24bd4b4, 32'h41dc3c5d, 32'hc1f60da4, 32'hc279d43d};
test_output[4427] = '{32'h423763a4};
test_index[4427] = '{3};
test_input[35424:35431] = '{32'hbfe5d8a0, 32'hc20aafcb, 32'hc2901db9, 32'hc249b85e, 32'hc281deed, 32'hc295b7fb, 32'h42a03557, 32'hc15e1463};
test_output[4428] = '{32'h42a03557};
test_index[4428] = '{6};
test_input[35432:35439] = '{32'hc26a41eb, 32'hc1b20bb9, 32'h425e3c45, 32'hc2a6292a, 32'h419f24cd, 32'hc291180e, 32'h42b60085, 32'h3f55e31d};
test_output[4429] = '{32'h42b60085};
test_index[4429] = '{6};
test_input[35440:35447] = '{32'hc2884abf, 32'hc23fb583, 32'hc2b48925, 32'h42a1cef7, 32'h4281ff0d, 32'hc264ba21, 32'h4297d92e, 32'hc2a1c0a9};
test_output[4430] = '{32'h42a1cef7};
test_index[4430] = '{3};
test_input[35448:35455] = '{32'h414e9f84, 32'hc19ae9b6, 32'hc25a48b7, 32'hc237c81b, 32'h41e0ef01, 32'h420901ce, 32'h424842ec, 32'hc03ad241};
test_output[4431] = '{32'h424842ec};
test_index[4431] = '{6};
test_input[35456:35463] = '{32'h42af1eb4, 32'hc2a73267, 32'h3f5fdf83, 32'h42411e0c, 32'hc2c7f63d, 32'h42317ecb, 32'hc217904b, 32'h41265700};
test_output[4432] = '{32'h42af1eb4};
test_index[4432] = '{0};
test_input[35464:35471] = '{32'h42af98f1, 32'h42317573, 32'hbfc3a4ed, 32'h3d8bf7eb, 32'h4206e09f, 32'hc29ec4c7, 32'hc2955d06, 32'hc285b590};
test_output[4433] = '{32'h42af98f1};
test_index[4433] = '{0};
test_input[35472:35479] = '{32'h41cfe697, 32'h41f40003, 32'hc1a39574, 32'h41fbabc5, 32'h3f2e61bf, 32'hc299f444, 32'hc200b707, 32'hc29594dc};
test_output[4434] = '{32'h41fbabc5};
test_index[4434] = '{3};
test_input[35480:35487] = '{32'h42838e6a, 32'h429e6300, 32'hc2c20bf6, 32'h429b32cb, 32'h429dbcec, 32'h413b2c0b, 32'h428f793e, 32'hc29ea59d};
test_output[4435] = '{32'h429e6300};
test_index[4435] = '{1};
test_input[35488:35495] = '{32'h42b71dae, 32'hc2c1c285, 32'h4276de2c, 32'h4223c1ff, 32'hc108c5f3, 32'h42c06fcd, 32'h42a6dae4, 32'h426b7505};
test_output[4436] = '{32'h42c06fcd};
test_index[4436] = '{5};
test_input[35496:35503] = '{32'h423ef120, 32'h42112bfc, 32'h423e80ea, 32'h41f48d0b, 32'hc1e87def, 32'hc22b0d6b, 32'h4255a7b6, 32'hc18adf9e};
test_output[4437] = '{32'h4255a7b6};
test_index[4437] = '{6};
test_input[35504:35511] = '{32'h42761f40, 32'h41f50743, 32'hc1a1344c, 32'h424c45e2, 32'h41f8e5ce, 32'hc24ecf82, 32'h4207acdb, 32'h4116898e};
test_output[4438] = '{32'h42761f40};
test_index[4438] = '{0};
test_input[35512:35519] = '{32'h422a5b9f, 32'hc2b14d2a, 32'hc281643c, 32'h425dbc27, 32'h420d63b2, 32'hc284df13, 32'hc1dc4aff, 32'hc2b45056};
test_output[4439] = '{32'h425dbc27};
test_index[4439] = '{3};
test_input[35520:35527] = '{32'hc062c00d, 32'hc1b666d6, 32'hc23a597c, 32'hc1c34101, 32'hc20cb380, 32'h42c4f5dd, 32'h41a71354, 32'hc2571905};
test_output[4440] = '{32'h42c4f5dd};
test_index[4440] = '{5};
test_input[35528:35535] = '{32'hc18c66a2, 32'hc28a836c, 32'hc2b56d14, 32'hc1f9e778, 32'h4290947c, 32'hc20f2b79, 32'h4215daf4, 32'hc294ac9b};
test_output[4441] = '{32'h4290947c};
test_index[4441] = '{4};
test_input[35536:35543] = '{32'hc2983938, 32'h42bfc4d2, 32'h41bb00ee, 32'hc29abc84, 32'hc224e563, 32'hc247d40b, 32'hc2785b1d, 32'hc28acdf4};
test_output[4442] = '{32'h42bfc4d2};
test_index[4442] = '{1};
test_input[35544:35551] = '{32'h4231df75, 32'h42b5747b, 32'h418a8b31, 32'hc28cab3f, 32'hc2419894, 32'h42acde3e, 32'hc1eb06ca, 32'hc168c27a};
test_output[4443] = '{32'h42b5747b};
test_index[4443] = '{1};
test_input[35552:35559] = '{32'hc221c225, 32'h40bcea61, 32'h42731060, 32'hc2bf8cae, 32'h4246ffc5, 32'h425e13b1, 32'h42b1f1a0, 32'hc1a4435c};
test_output[4444] = '{32'h42b1f1a0};
test_index[4444] = '{6};
test_input[35560:35567] = '{32'hc1916da4, 32'h42895859, 32'h42270bdb, 32'h429c275b, 32'h42174438, 32'h4249048b, 32'hc2165500, 32'h42014345};
test_output[4445] = '{32'h429c275b};
test_index[4445] = '{3};
test_input[35568:35575] = '{32'h42a4ee79, 32'h3f1df3a5, 32'hc0d271d4, 32'h4287e9b7, 32'hc2c14cb0, 32'h4293dad3, 32'hc193729d, 32'h41af574c};
test_output[4446] = '{32'h42a4ee79};
test_index[4446] = '{0};
test_input[35576:35583] = '{32'h429adb93, 32'hc21e6054, 32'h417103d6, 32'hc2aa9037, 32'h428897c2, 32'h422a4492, 32'h41356e2c, 32'hc0ab1609};
test_output[4447] = '{32'h429adb93};
test_index[4447] = '{0};
test_input[35584:35591] = '{32'h421da153, 32'hc28c1251, 32'h4222a41f, 32'h411385c2, 32'hbfc56ca7, 32'hc0a4b5f6, 32'h41ede4ef, 32'hc2af9750};
test_output[4448] = '{32'h4222a41f};
test_index[4448] = '{2};
test_input[35592:35599] = '{32'hc2bf6ae7, 32'h42220e78, 32'h4143f10e, 32'h42501deb, 32'hc2aa5722, 32'h42666f3a, 32'h41ee6b74, 32'h420f2e2b};
test_output[4449] = '{32'h42666f3a};
test_index[4449] = '{5};
test_input[35600:35607] = '{32'hc196844d, 32'h42bbd383, 32'hc24bed2b, 32'h41241f8e, 32'h4259ac7a, 32'hc2604fc4, 32'h41bf89ea, 32'hc2297231};
test_output[4450] = '{32'h42bbd383};
test_index[4450] = '{1};
test_input[35608:35615] = '{32'hc1e88467, 32'h421201d9, 32'hc1a8737f, 32'hc1f4e248, 32'hc2b311e7, 32'hc28b4d1a, 32'h423f17b5, 32'hc2858d1c};
test_output[4451] = '{32'h423f17b5};
test_index[4451] = '{6};
test_input[35616:35623] = '{32'hc16c318d, 32'hc190ab85, 32'hc26056f7, 32'h4174798d, 32'hc2aadfd8, 32'h42840181, 32'h42b6c2bf, 32'h41813cc9};
test_output[4452] = '{32'h42b6c2bf};
test_index[4452] = '{6};
test_input[35624:35631] = '{32'h41b91ed5, 32'hc0f46f22, 32'h418ca33c, 32'hc20b45e4, 32'h429c90ab, 32'h417636f4, 32'h426c09fb, 32'hc23703fa};
test_output[4453] = '{32'h429c90ab};
test_index[4453] = '{4};
test_input[35632:35639] = '{32'h4295124b, 32'hc23854b5, 32'h41d127b0, 32'h426f9ce3, 32'hc2844413, 32'hc25ef356, 32'hc226b3af, 32'hc23153a0};
test_output[4454] = '{32'h4295124b};
test_index[4454] = '{0};
test_input[35640:35647] = '{32'hc2978e44, 32'hc1b6a19c, 32'h4251fed3, 32'hc1d8f855, 32'h429f2889, 32'hc21a4fed, 32'hc26b28b2, 32'h42952c83};
test_output[4455] = '{32'h429f2889};
test_index[4455] = '{4};
test_input[35648:35655] = '{32'h42483c8a, 32'hc20d3ac7, 32'hc2a275b2, 32'h42160401, 32'hc14f5572, 32'hc2ad7696, 32'hc01d37a1, 32'h421bc10e};
test_output[4456] = '{32'h42483c8a};
test_index[4456] = '{0};
test_input[35656:35663] = '{32'hc13853cb, 32'h41c78393, 32'hc26fdee9, 32'hc1cfabc2, 32'h41f508ed, 32'h427bb04a, 32'h420a9fd1, 32'hc1b82800};
test_output[4457] = '{32'h427bb04a};
test_index[4457] = '{5};
test_input[35664:35671] = '{32'h4180dc17, 32'h42295244, 32'hc2181453, 32'h42c1a84b, 32'hc1aadd2d, 32'hc28f17f1, 32'hc2bcd05e, 32'h4234fab9};
test_output[4458] = '{32'h42c1a84b};
test_index[4458] = '{3};
test_input[35672:35679] = '{32'hc1e2cd3b, 32'h4213a23c, 32'hc2b49c5d, 32'hc1d492bd, 32'h42b5e146, 32'hc259044a, 32'hc29f7f17, 32'h41955891};
test_output[4459] = '{32'h42b5e146};
test_index[4459] = '{4};
test_input[35680:35687] = '{32'h419adcba, 32'hc17f9231, 32'hc2a7cd98, 32'hc28db8e4, 32'h42720a5d, 32'h425223e7, 32'h41a65617, 32'hc28918eb};
test_output[4460] = '{32'h42720a5d};
test_index[4460] = '{4};
test_input[35688:35695] = '{32'hc20be091, 32'hc241d1e4, 32'hc1cb38fb, 32'h42c2df66, 32'h4246b505, 32'h4242d7ba, 32'h4157c5a1, 32'hc2426f58};
test_output[4461] = '{32'h42c2df66};
test_index[4461] = '{3};
test_input[35696:35703] = '{32'h4136a53d, 32'h41d33f38, 32'h42c764af, 32'h425cb12b, 32'hc2952f16, 32'hc287900d, 32'hc20ebec4, 32'hc1141e13};
test_output[4462] = '{32'h42c764af};
test_index[4462] = '{2};
test_input[35704:35711] = '{32'hc28dd3fc, 32'h40a88745, 32'h42a63cba, 32'h423de41a, 32'hc12d51bd, 32'h4295cc11, 32'h41b54af9, 32'hc22873f4};
test_output[4463] = '{32'h42a63cba};
test_index[4463] = '{2};
test_input[35712:35719] = '{32'h40790650, 32'h42764d2c, 32'h422e4779, 32'h41007dd6, 32'h429e90ab, 32'hc25c0b8b, 32'h429bb877, 32'h42013f6d};
test_output[4464] = '{32'h429e90ab};
test_index[4464] = '{4};
test_input[35720:35727] = '{32'h4295be80, 32'h40b67e25, 32'h413bc720, 32'h41818435, 32'h425fe609, 32'hc2915886, 32'hc28a58d0, 32'hc2697528};
test_output[4465] = '{32'h4295be80};
test_index[4465] = '{0};
test_input[35728:35735] = '{32'hc1e89605, 32'hc25a062e, 32'hc21a3c1d, 32'h41b308d5, 32'h3fa4df9f, 32'h413e5e09, 32'hc2b3aac0, 32'h41e9d965};
test_output[4466] = '{32'h41e9d965};
test_index[4466] = '{7};
test_input[35736:35743] = '{32'h4002e98a, 32'hc0df8000, 32'h4288941b, 32'hc1a67a2d, 32'h41f71815, 32'h41c84317, 32'h4266a723, 32'hc1bac055};
test_output[4467] = '{32'h4288941b};
test_index[4467] = '{2};
test_input[35744:35751] = '{32'hc29aedb4, 32'hc2898745, 32'h42b7a715, 32'hc2088a18, 32'hc08d9290, 32'hc1e132cf, 32'hbf2fbb5b, 32'hc147e18b};
test_output[4468] = '{32'h42b7a715};
test_index[4468] = '{2};
test_input[35752:35759] = '{32'h42895d14, 32'hc1e2a0a8, 32'h42c57cbe, 32'hc2b56e0f, 32'hc2b9a0f6, 32'hc2a49304, 32'h41d10231, 32'h4197be69};
test_output[4469] = '{32'h42c57cbe};
test_index[4469] = '{2};
test_input[35760:35767] = '{32'h405b2e28, 32'hc24f931a, 32'h41c519b0, 32'hc245904a, 32'hc263dc67, 32'hc289d001, 32'h41ed5879, 32'h4283e1cd};
test_output[4470] = '{32'h4283e1cd};
test_index[4470] = '{7};
test_input[35768:35775] = '{32'hc106b86c, 32'hc218b7a2, 32'hc056b25b, 32'hc2ae8953, 32'h429cec94, 32'hc142445f, 32'h3e3ce370, 32'h42919975};
test_output[4471] = '{32'h429cec94};
test_index[4471] = '{4};
test_input[35776:35783] = '{32'hc297f0ba, 32'hc29af595, 32'hc288a165, 32'hc1a9bc35, 32'hc2919907, 32'h427e874e, 32'hc104d9c6, 32'hc25e1f95};
test_output[4472] = '{32'h427e874e};
test_index[4472] = '{5};
test_input[35784:35791] = '{32'hc11a01dc, 32'hc2c7362e, 32'hc1a89568, 32'h4149edd5, 32'h41e0f7b5, 32'hbf9f7281, 32'h4263e1c7, 32'hc18be43a};
test_output[4473] = '{32'h4263e1c7};
test_index[4473] = '{6};
test_input[35792:35799] = '{32'h42256ef5, 32'hbfa46d33, 32'h42688201, 32'hc29f1bc5, 32'hc2b628da, 32'hc22a2acc, 32'hc2b46b1e, 32'h41fa49ca};
test_output[4474] = '{32'h42688201};
test_index[4474] = '{2};
test_input[35800:35807] = '{32'h42a4089f, 32'h4285c4ae, 32'h4254b6a3, 32'hc1d3b213, 32'h428ec4d4, 32'hc29859b0, 32'h42af1387, 32'hc225564b};
test_output[4475] = '{32'h42af1387};
test_index[4475] = '{6};
test_input[35808:35815] = '{32'hc28ef124, 32'h4203f6d2, 32'h42817fac, 32'hc2bf24ee, 32'hc23a7293, 32'h41eb0f42, 32'hc2017380, 32'hc0bae2da};
test_output[4476] = '{32'h42817fac};
test_index[4476] = '{2};
test_input[35816:35823] = '{32'hc1ade24d, 32'hc281887a, 32'h42491eed, 32'h4283233d, 32'h41dc41f9, 32'hc18043a2, 32'h426d7264, 32'h3fc1c94b};
test_output[4477] = '{32'h4283233d};
test_index[4477] = '{3};
test_input[35824:35831] = '{32'hc1e498b9, 32'h428536c7, 32'h40943ee3, 32'h421c51b1, 32'hc28a1e5c, 32'hc1aeb0ed, 32'h42831170, 32'h4291dc2b};
test_output[4478] = '{32'h4291dc2b};
test_index[4478] = '{7};
test_input[35832:35839] = '{32'h428a293b, 32'h42c17584, 32'hc2ac51e4, 32'h421575a4, 32'hc0939ba1, 32'hc28a86d9, 32'h42ac181b, 32'hc2aa8f57};
test_output[4479] = '{32'h42c17584};
test_index[4479] = '{1};
test_input[35840:35847] = '{32'hc1b0e4e7, 32'hc1febd05, 32'h42be2b76, 32'hc29b7eb6, 32'hc0401918, 32'hc1b26703, 32'h42b26670, 32'h422a9c10};
test_output[4480] = '{32'h42be2b76};
test_index[4480] = '{2};
test_input[35848:35855] = '{32'hc29594e4, 32'h412d6d6d, 32'hc292a69d, 32'h42547f67, 32'h41cc23a5, 32'hc1a78e4c, 32'h4284df7d, 32'hc240e131};
test_output[4481] = '{32'h4284df7d};
test_index[4481] = '{6};
test_input[35856:35863] = '{32'hc1b0a566, 32'h428b095b, 32'hc22282d6, 32'h427b5714, 32'h4208931c, 32'hbe84e202, 32'h41808a85, 32'hc218946b};
test_output[4482] = '{32'h428b095b};
test_index[4482] = '{1};
test_input[35864:35871] = '{32'h42b08c3e, 32'hc1ca9fa5, 32'hc28b1375, 32'hc28d53c1, 32'hc258c8ed, 32'h423fb7b9, 32'hc2add79a, 32'hc0729e07};
test_output[4483] = '{32'h42b08c3e};
test_index[4483] = '{0};
test_input[35872:35879] = '{32'h41daeed5, 32'h42bbca19, 32'h426fd3f4, 32'hc2970846, 32'h41d3c20d, 32'h42875cc0, 32'h41e05f90, 32'hc115ac04};
test_output[4484] = '{32'h42bbca19};
test_index[4484] = '{1};
test_input[35880:35887] = '{32'h429182c6, 32'hc2b5c89a, 32'hc28e8a8d, 32'h4062938c, 32'h4086aedb, 32'hc27c4924, 32'hc28f315a, 32'hc20946a6};
test_output[4485] = '{32'h429182c6};
test_index[4485] = '{0};
test_input[35888:35895] = '{32'hc0ec735e, 32'h4232626b, 32'hc10c61ca, 32'hc0a060b4, 32'hc1ab5fe2, 32'hc23afd02, 32'h4251db55, 32'h42129945};
test_output[4486] = '{32'h4251db55};
test_index[4486] = '{6};
test_input[35896:35903] = '{32'h421506c0, 32'hc1eb71db, 32'h428b5ecd, 32'h42a40003, 32'h41e6cefc, 32'hc2b91d5e, 32'h42aa7146, 32'h4270f95f};
test_output[4487] = '{32'h42aa7146};
test_index[4487] = '{6};
test_input[35904:35911] = '{32'h428c8635, 32'h428061e4, 32'h42b6e660, 32'h4021456d, 32'hc1305501, 32'h42b89d4d, 32'h4284d403, 32'hc2023d2e};
test_output[4488] = '{32'h42b89d4d};
test_index[4488] = '{5};
test_input[35912:35919] = '{32'h42935abf, 32'h42c125f7, 32'h41d957ad, 32'hc2168e77, 32'hc28a7a46, 32'hc2bf36e2, 32'hc2855fae, 32'hc28947e9};
test_output[4489] = '{32'h42c125f7};
test_index[4489] = '{1};
test_input[35920:35927] = '{32'h427c1e7f, 32'h4277bce9, 32'h418b57d7, 32'hc292c853, 32'h4298e3d5, 32'h42ab5967, 32'h42c08d92, 32'hc131d68b};
test_output[4490] = '{32'h42c08d92};
test_index[4490] = '{6};
test_input[35928:35935] = '{32'h4117c0a5, 32'h42b61628, 32'h4251162a, 32'h418cfee0, 32'hc2aadf65, 32'hc02a4fb9, 32'hc2282a3e, 32'h41db10c2};
test_output[4491] = '{32'h42b61628};
test_index[4491] = '{1};
test_input[35936:35943] = '{32'hc1819ae9, 32'hc2a2b80e, 32'h42c73e3a, 32'hc27bbadf, 32'h428be43f, 32'h4203078f, 32'h428cf45b, 32'hc1549863};
test_output[4492] = '{32'h42c73e3a};
test_index[4492] = '{2};
test_input[35944:35951] = '{32'hc122ea1b, 32'hc20ddfaf, 32'hc28704e5, 32'hc1870cad, 32'hc2486a20, 32'hc2bb208e, 32'hc1db1ec9, 32'hc28a3434};
test_output[4493] = '{32'hc122ea1b};
test_index[4493] = '{0};
test_input[35952:35959] = '{32'h42a0514e, 32'hc196ddc3, 32'h428524e5, 32'hc2bf1c81, 32'hc2a3a474, 32'h41fd0b23, 32'h4280ac4c, 32'h42b0f2d8};
test_output[4494] = '{32'h42b0f2d8};
test_index[4494] = '{7};
test_input[35960:35967] = '{32'h409bd393, 32'h4257fc28, 32'h4183862e, 32'h41b163fc, 32'hc2a553dd, 32'h424b94e8, 32'hc20e9e64, 32'hc227c220};
test_output[4495] = '{32'h4257fc28};
test_index[4495] = '{1};
test_input[35968:35975] = '{32'hc1776b80, 32'h428c0fc8, 32'h413e3bf0, 32'h4224521b, 32'h412104c1, 32'h42294663, 32'hc02cd96c, 32'hc2a6115b};
test_output[4496] = '{32'h428c0fc8};
test_index[4496] = '{1};
test_input[35976:35983] = '{32'h421de76a, 32'hc255be64, 32'hc2b0c865, 32'h428e7769, 32'h42267de5, 32'hc2a9f3af, 32'h41ff4e97, 32'hc2666781};
test_output[4497] = '{32'h428e7769};
test_index[4497] = '{3};
test_input[35984:35991] = '{32'hc24a043c, 32'hc1aba0f2, 32'h4159dc1d, 32'h413b691b, 32'hc2bddc32, 32'hc287850e, 32'h4290888a, 32'hc2b1e2a5};
test_output[4498] = '{32'h4290888a};
test_index[4498] = '{6};
test_input[35992:35999] = '{32'h42a531a2, 32'hc1afec28, 32'h428ff13f, 32'hc2ba4aa8, 32'hc222f6dc, 32'hc2c2569d, 32'hc2aaa8c9, 32'hc2124f35};
test_output[4499] = '{32'h42a531a2};
test_index[4499] = '{0};
test_input[36000:36007] = '{32'h424a5bf5, 32'hc2988f64, 32'hc169f6fd, 32'h41b4462b, 32'hc2a8e656, 32'hc2c5f318, 32'h42abc911, 32'h42b6a261};
test_output[4500] = '{32'h42b6a261};
test_index[4500] = '{7};
test_input[36008:36015] = '{32'h427e1b32, 32'hc259be77, 32'hc27cc456, 32'hc1e43087, 32'hbe9998c6, 32'hc1bc5a0a, 32'h429f03ad, 32'h41f3380d};
test_output[4501] = '{32'h429f03ad};
test_index[4501] = '{6};
test_input[36016:36023] = '{32'h4208002c, 32'hc21569af, 32'h426094dd, 32'hc2859671, 32'h42af4e38, 32'h41e6f500, 32'hc0bae77c, 32'hc2b81f03};
test_output[4502] = '{32'h42af4e38};
test_index[4502] = '{4};
test_input[36024:36031] = '{32'h41314c32, 32'hc1a2908e, 32'h41faecfd, 32'h4297677e, 32'h42a3db71, 32'h4234fe56, 32'h4229f503, 32'hc284096c};
test_output[4503] = '{32'h42a3db71};
test_index[4503] = '{4};
test_input[36032:36039] = '{32'h4279a5d4, 32'h3fdee19e, 32'h406e26a3, 32'h422bb6d7, 32'hc1d72a67, 32'h42a5c026, 32'hc2886591, 32'h42a6baac};
test_output[4504] = '{32'h42a6baac};
test_index[4504] = '{7};
test_input[36040:36047] = '{32'hc20c3894, 32'hc210473c, 32'hc1b6a71d, 32'hc1a1de2c, 32'hc2329b8e, 32'h41fa50e3, 32'h42693805, 32'h42ab7279};
test_output[4505] = '{32'h42ab7279};
test_index[4505] = '{7};
test_input[36048:36055] = '{32'h42358fb4, 32'hc29320c9, 32'hc2a40d72, 32'hc1d7f895, 32'h4066eb89, 32'h42bde795, 32'h42668a27, 32'hc219f06b};
test_output[4506] = '{32'h42bde795};
test_index[4506] = '{5};
test_input[36056:36063] = '{32'h4287805e, 32'h41a2ed69, 32'h411bd1be, 32'h42102959, 32'h4286e76d, 32'h4287a359, 32'h427ff30b, 32'h4196095d};
test_output[4507] = '{32'h4287a359};
test_index[4507] = '{5};
test_input[36064:36071] = '{32'h4141ddf6, 32'hc2579d96, 32'h42bf28fe, 32'hc222cbbb, 32'h41fdb892, 32'h41fb9ca7, 32'h42c1788f, 32'hc1b72430};
test_output[4508] = '{32'h42c1788f};
test_index[4508] = '{6};
test_input[36072:36079] = '{32'h42152687, 32'h42b9d71b, 32'hc21a8703, 32'hc25b5988, 32'hc1d6ce25, 32'h42844c6b, 32'h425e0d54, 32'h421725b6};
test_output[4509] = '{32'h42b9d71b};
test_index[4509] = '{1};
test_input[36080:36087] = '{32'h4146eda2, 32'hc2188558, 32'hc0f6fcec, 32'hc281d774, 32'hc27e2020, 32'hc2bfb43d, 32'hc29c1740, 32'hc133fc34};
test_output[4510] = '{32'h4146eda2};
test_index[4510] = '{0};
test_input[36088:36095] = '{32'hc1fd9d1b, 32'hc24799ae, 32'hc1dcd578, 32'hc293f36d, 32'h411efb5f, 32'hc29e3836, 32'h42336118, 32'h42c0c596};
test_output[4511] = '{32'h42c0c596};
test_index[4511] = '{7};
test_input[36096:36103] = '{32'h4208dcf7, 32'hc213f387, 32'hc2215c54, 32'hc18cf423, 32'h3ee2213a, 32'h42a65fd2, 32'h4270ba99, 32'hc2aa4e2c};
test_output[4512] = '{32'h42a65fd2};
test_index[4512] = '{5};
test_input[36104:36111] = '{32'h418958f2, 32'h4281269f, 32'hc2a7d004, 32'hc1b1cd63, 32'hc1d5da9a, 32'hc1aea57b, 32'hc2af0dc9, 32'h40d831ad};
test_output[4513] = '{32'h4281269f};
test_index[4513] = '{1};
test_input[36112:36119] = '{32'h42abf681, 32'h427b13b5, 32'h4252af94, 32'hc156ff36, 32'h42b31850, 32'hc2a9689d, 32'h42ba2b3d, 32'hc2107e43};
test_output[4514] = '{32'h42ba2b3d};
test_index[4514] = '{6};
test_input[36120:36127] = '{32'h4298eaf7, 32'h428d76cc, 32'h42413d69, 32'h428aa35b, 32'hc27038e3, 32'hc149e8dd, 32'hc25d65d6, 32'hc13503bc};
test_output[4515] = '{32'h4298eaf7};
test_index[4515] = '{0};
test_input[36128:36135] = '{32'hc2aa4df6, 32'hc1b33b5b, 32'hc2574734, 32'hc2a52316, 32'hc206831d, 32'h3ef91441, 32'h41c2b69e, 32'hc2bf11e6};
test_output[4516] = '{32'h41c2b69e};
test_index[4516] = '{6};
test_input[36136:36143] = '{32'hc0acd061, 32'h418624ce, 32'hc24230d8, 32'hc252ab1a, 32'h424e734f, 32'h42bfee46, 32'hc2bc657d, 32'hc28c272c};
test_output[4517] = '{32'h42bfee46};
test_index[4517] = '{5};
test_input[36144:36151] = '{32'h41d62286, 32'h40d28476, 32'hc200b62f, 32'hc204b6f6, 32'hc2c144b0, 32'h42733273, 32'h4290f907, 32'hc2879478};
test_output[4518] = '{32'h4290f907};
test_index[4518] = '{6};
test_input[36152:36159] = '{32'hc23d4fe4, 32'hc175dec1, 32'h42561954, 32'h428e98d9, 32'hc20da0d9, 32'h42380d7b, 32'hc273882a, 32'hc2979043};
test_output[4519] = '{32'h428e98d9};
test_index[4519] = '{3};
test_input[36160:36167] = '{32'h4295ce3f, 32'hc293acf2, 32'h41046739, 32'h428170e2, 32'hc21037ff, 32'h42bf5d33, 32'hc1751a72, 32'hc2bcd97b};
test_output[4520] = '{32'h42bf5d33};
test_index[4520] = '{5};
test_input[36168:36175] = '{32'hc2ada082, 32'h418fdcaa, 32'hc282d8fc, 32'hc277bde7, 32'hc29b4ca3, 32'hc2c754f1, 32'h41ea86dc, 32'h40b8cc30};
test_output[4521] = '{32'h41ea86dc};
test_index[4521] = '{6};
test_input[36176:36183] = '{32'hc2b51fd0, 32'hc29668dd, 32'h42ae8cbb, 32'h40a6ef7e, 32'hc18311bd, 32'hc26dc83c, 32'hc2b15abd, 32'h40015818};
test_output[4522] = '{32'h42ae8cbb};
test_index[4522] = '{2};
test_input[36184:36191] = '{32'hc2bd3736, 32'h42ab6edd, 32'h42007dc5, 32'hc12fe22d, 32'hc253ee67, 32'h41e9cf12, 32'hc26bdad4, 32'h42a0fdb6};
test_output[4523] = '{32'h42ab6edd};
test_index[4523] = '{1};
test_input[36192:36199] = '{32'h41e8543d, 32'hc2936cb2, 32'h42885d36, 32'h42a3d7f1, 32'h424d59b5, 32'h42beb1a1, 32'h42680dbd, 32'hc29676cc};
test_output[4524] = '{32'h42beb1a1};
test_index[4524] = '{5};
test_input[36200:36207] = '{32'h41f66a88, 32'hc24b680e, 32'h42c1384f, 32'hc203e311, 32'h41961b9d, 32'h4128bf7f, 32'h4296dcee, 32'h41e94b9c};
test_output[4525] = '{32'h42c1384f};
test_index[4525] = '{2};
test_input[36208:36215] = '{32'hc2baccbb, 32'h427be04e, 32'hc2ba632e, 32'hc2054de8, 32'hc1ae6e6c, 32'hc2918d73, 32'h4126ce30, 32'h428c70ad};
test_output[4526] = '{32'h428c70ad};
test_index[4526] = '{7};
test_input[36216:36223] = '{32'h42365e80, 32'h42a0ea1f, 32'h41dcc723, 32'h42260c2d, 32'hc26d9f98, 32'h40008b08, 32'hc19d8bd2, 32'hc278dec2};
test_output[4527] = '{32'h42a0ea1f};
test_index[4527] = '{1};
test_input[36224:36231] = '{32'h42a524cc, 32'h42c160b6, 32'h4181d9c6, 32'hc144815a, 32'h41c748b9, 32'hc287148c, 32'hc15864da, 32'h414ef980};
test_output[4528] = '{32'h42c160b6};
test_index[4528] = '{1};
test_input[36232:36239] = '{32'h42436262, 32'h4291fb38, 32'hc18d0082, 32'h42985210, 32'hc0cebbbe, 32'hc27dca4b, 32'hc2a05828, 32'hc23a6ef5};
test_output[4529] = '{32'h42985210};
test_index[4529] = '{3};
test_input[36240:36247] = '{32'h42162569, 32'hc25bd1eb, 32'h4283d93b, 32'hc2aee0e4, 32'hc261f67a, 32'hc2a58f00, 32'hc2829351, 32'h42375d09};
test_output[4530] = '{32'h4283d93b};
test_index[4530] = '{2};
test_input[36248:36255] = '{32'h425617eb, 32'hc242af5e, 32'hc249dbe8, 32'h424fe819, 32'hc2a110c6, 32'hc2993a76, 32'hc0c9b6f7, 32'hc2bd97c0};
test_output[4531] = '{32'h425617eb};
test_index[4531] = '{0};
test_input[36256:36263] = '{32'h423c4ea2, 32'h42115d55, 32'h429d0dca, 32'hc1a25163, 32'hc2beba7f, 32'hc29aeed3, 32'h422a3d65, 32'hc0af5bcc};
test_output[4532] = '{32'h429d0dca};
test_index[4532] = '{2};
test_input[36264:36271] = '{32'hc24e84e4, 32'hc2879762, 32'h42b02e77, 32'h42c25adf, 32'h41f4819a, 32'hc2b36f2f, 32'h427b2740, 32'hc1e4be7c};
test_output[4533] = '{32'h42c25adf};
test_index[4533] = '{3};
test_input[36272:36279] = '{32'h41d2db2a, 32'hc19dd2b2, 32'hc260f4d8, 32'hc0aba73c, 32'h3fcfefaa, 32'h41f08d7f, 32'hc2bd7c13, 32'h423a41d5};
test_output[4534] = '{32'h423a41d5};
test_index[4534] = '{7};
test_input[36280:36287] = '{32'hc0c0ef55, 32'h42be9ffe, 32'h4272163d, 32'h429fd139, 32'hc282c04e, 32'hbfce88fe, 32'h42412c6b, 32'hc226b46f};
test_output[4535] = '{32'h42be9ffe};
test_index[4535] = '{1};
test_input[36288:36295] = '{32'hc2aa8743, 32'h41e69539, 32'hc1cf1c7b, 32'h425df01f, 32'hc2bb663d, 32'hc28c2a17, 32'h429e3f63, 32'hc1e9c990};
test_output[4536] = '{32'h429e3f63};
test_index[4536] = '{6};
test_input[36296:36303] = '{32'hc1c30d13, 32'h42b0c948, 32'hbd7bb85b, 32'h41a5c676, 32'hc2a0f2fc, 32'h426d3b08, 32'h429cf722, 32'h42bfa4c1};
test_output[4537] = '{32'h42bfa4c1};
test_index[4537] = '{7};
test_input[36304:36311] = '{32'h42c6a6ee, 32'hc2914022, 32'hc21f6eb2, 32'h3f847ecf, 32'hc2c1a7a6, 32'h42675b41, 32'hc2a8f0f9, 32'hc1037a77};
test_output[4538] = '{32'h42c6a6ee};
test_index[4538] = '{0};
test_input[36312:36319] = '{32'hc216876a, 32'h4276bfd0, 32'hc22de348, 32'h42ae7bf9, 32'h42501e90, 32'hc2c35bc6, 32'h4249a7e3, 32'h42b6e734};
test_output[4539] = '{32'h42b6e734};
test_index[4539] = '{7};
test_input[36320:36327] = '{32'h41fed935, 32'h420066e1, 32'h4292a94d, 32'hc26041f2, 32'hc1dc18f0, 32'hc2aa10a9, 32'hc229e546, 32'h4126b72d};
test_output[4540] = '{32'h4292a94d};
test_index[4540] = '{2};
test_input[36328:36335] = '{32'hc07ac4ba, 32'hc1564938, 32'h4275c29b, 32'hc1f3c818, 32'h42a02f3b, 32'h3fdadc2a, 32'hc22f4f20, 32'h4285b85f};
test_output[4541] = '{32'h42a02f3b};
test_index[4541] = '{4};
test_input[36336:36343] = '{32'hc20c36a5, 32'hc2a0146a, 32'h419ac8b4, 32'hc2587095, 32'h424d43be, 32'hc2468b1e, 32'hbe4b5652, 32'h41f69306};
test_output[4542] = '{32'h424d43be};
test_index[4542] = '{4};
test_input[36344:36351] = '{32'h41069fa1, 32'hc228111a, 32'h4240759b, 32'h4232ad62, 32'hc0931afa, 32'hc239a289, 32'h40e530a9, 32'hc2bdc501};
test_output[4543] = '{32'h4240759b};
test_index[4543] = '{2};
test_input[36352:36359] = '{32'hc1346f5a, 32'hc21d4a0c, 32'hc1ecc0bf, 32'h3d1b7cb1, 32'h41d4349e, 32'hc26de1d7, 32'hc22711d2, 32'hc255fce9};
test_output[4544] = '{32'h41d4349e};
test_index[4544] = '{4};
test_input[36360:36367] = '{32'hc1bc1b9e, 32'hc21d6182, 32'hc2bf8653, 32'hc1b2e8d1, 32'h42b04493, 32'hc07effec, 32'h42a3c1e2, 32'h416a21bb};
test_output[4545] = '{32'h42b04493};
test_index[4545] = '{4};
test_input[36368:36375] = '{32'h423683e1, 32'h41bdf67c, 32'hc2438550, 32'h428d152b, 32'h427956d8, 32'hc2bb0ff8, 32'h42683213, 32'h421e53e4};
test_output[4546] = '{32'h428d152b};
test_index[4546] = '{3};
test_input[36376:36383] = '{32'h42352eb9, 32'h42bf0217, 32'hc2866be8, 32'hc203f2f7, 32'h42018cb6, 32'hc21aeec2, 32'hbf0b4a83, 32'h411d1a15};
test_output[4547] = '{32'h42bf0217};
test_index[4547] = '{1};
test_input[36384:36391] = '{32'h42949d19, 32'h417dffea, 32'hc29abf08, 32'hc296d102, 32'hc08af714, 32'h42016d63, 32'h42c76f77, 32'h42936d0c};
test_output[4548] = '{32'h42c76f77};
test_index[4548] = '{6};
test_input[36392:36399] = '{32'h42b44fcd, 32'hc2167656, 32'h4297c5c9, 32'h41bbd4a6, 32'h42ae087f, 32'h42a990a3, 32'hbfd328e5, 32'h428d5c2c};
test_output[4549] = '{32'h42b44fcd};
test_index[4549] = '{0};
test_input[36400:36407] = '{32'hc1392b6a, 32'hc1e01379, 32'hc2908a52, 32'hc2c1f9b2, 32'h42a858d6, 32'h418484b8, 32'h4277d7b5, 32'h428f8559};
test_output[4550] = '{32'h42a858d6};
test_index[4550] = '{4};
test_input[36408:36415] = '{32'h41c917c1, 32'hc2496697, 32'h426ce947, 32'hc16fec6f, 32'h42971cae, 32'h4284b3e1, 32'hc121902d, 32'h41ccd34f};
test_output[4551] = '{32'h42971cae};
test_index[4551] = '{4};
test_input[36416:36423] = '{32'hc23cd8e0, 32'h41effe98, 32'hc2abdff5, 32'hc26b74dd, 32'hc2a819eb, 32'hc29e3771, 32'hc229bff3, 32'h42ac001d};
test_output[4552] = '{32'h42ac001d};
test_index[4552] = '{7};
test_input[36424:36431] = '{32'hc0c0a695, 32'hc18488db, 32'h42224384, 32'h4185f0ac, 32'hc1f47391, 32'hc21f294f, 32'hc1d4198f, 32'h4228e7b8};
test_output[4553] = '{32'h4228e7b8};
test_index[4553] = '{7};
test_input[36432:36439] = '{32'hc20867af, 32'hc01ceb22, 32'h42c44d09, 32'h4229a04c, 32'h41e1f7e5, 32'h41774d36, 32'h415b4ff2, 32'h40bc55b9};
test_output[4554] = '{32'h42c44d09};
test_index[4554] = '{2};
test_input[36440:36447] = '{32'hc2c3d1c6, 32'h42a5fbe4, 32'hc2195220, 32'h427f1360, 32'h40e62a52, 32'h41d906cc, 32'hc287fdde, 32'hc1d4223b};
test_output[4555] = '{32'h42a5fbe4};
test_index[4555] = '{1};
test_input[36448:36455] = '{32'h42224ef2, 32'hc28d2f20, 32'h4210c6dc, 32'hc283296f, 32'hc284403c, 32'h42973ac4, 32'hc1dd7674, 32'h4293afb3};
test_output[4556] = '{32'h42973ac4};
test_index[4556] = '{5};
test_input[36456:36463] = '{32'h42440bd6, 32'h428eb33c, 32'h4224b605, 32'hc01d404c, 32'h40b670f1, 32'hc255f593, 32'h42b47266, 32'h42ae8a00};
test_output[4557] = '{32'h42b47266};
test_index[4557] = '{6};
test_input[36464:36471] = '{32'h429a3946, 32'hc2158e30, 32'hc1a35314, 32'hc283ff5f, 32'hc2a0a44b, 32'h427191c6, 32'hc23f610e, 32'h4227515b};
test_output[4558] = '{32'h429a3946};
test_index[4558] = '{0};
test_input[36472:36479] = '{32'h429d83bc, 32'hc1b74d68, 32'h42c7770a, 32'h41f783de, 32'hc0c54178, 32'hc1bf953b, 32'hc2872ef2, 32'h42714d87};
test_output[4559] = '{32'h42c7770a};
test_index[4559] = '{2};
test_input[36480:36487] = '{32'hc150fc3c, 32'hc2045004, 32'hc299b67b, 32'h41fc09fc, 32'h411c1cbc, 32'hc17a147d, 32'h41b50a47, 32'h40c81a8f};
test_output[4560] = '{32'h41fc09fc};
test_index[4560] = '{3};
test_input[36488:36495] = '{32'hc07b700b, 32'hc2a6c28e, 32'h421fc373, 32'h3fcbb4e0, 32'hc085b483, 32'h42a3cbe9, 32'h42a29c15, 32'hc2300899};
test_output[4561] = '{32'h42a3cbe9};
test_index[4561] = '{5};
test_input[36496:36503] = '{32'hc18a4d60, 32'hc180842f, 32'h429b3b4c, 32'h4253bf28, 32'hc26bf65b, 32'h428d6513, 32'hc09376bb, 32'hc16b767b};
test_output[4562] = '{32'h429b3b4c};
test_index[4562] = '{2};
test_input[36504:36511] = '{32'hc002b11c, 32'hc245dc33, 32'h42427918, 32'hc2ae7bd1, 32'hc29aa194, 32'hc29f8b7d, 32'h41e9c69e, 32'h41cbe47f};
test_output[4563] = '{32'h42427918};
test_index[4563] = '{2};
test_input[36512:36519] = '{32'h4295858d, 32'hc23bff13, 32'hc2c24bfa, 32'hc2a84e85, 32'hc1f31c39, 32'hc20ce998, 32'h42b0b8fd, 32'h425dc9b2};
test_output[4564] = '{32'h42b0b8fd};
test_index[4564] = '{6};
test_input[36520:36527] = '{32'hc2979466, 32'h419c2485, 32'hc2c4b896, 32'h419f6716, 32'hc190a632, 32'h426b1524, 32'hc1e241ee, 32'h42afc90c};
test_output[4565] = '{32'h42afc90c};
test_index[4565] = '{7};
test_input[36528:36535] = '{32'hc18883d0, 32'hc274d1e2, 32'h41036fdb, 32'hc104c81a, 32'hc2669c4d, 32'h420f5a7e, 32'h4266ee0a, 32'hc1aa200b};
test_output[4566] = '{32'h4266ee0a};
test_index[4566] = '{6};
test_input[36536:36543] = '{32'h42c3cd56, 32'hc2972000, 32'hc1864f9b, 32'hc2ba6da7, 32'hc2b61020, 32'h42184cdd, 32'hc266d24e, 32'hc29b3a04};
test_output[4567] = '{32'h42c3cd56};
test_index[4567] = '{0};
test_input[36544:36551] = '{32'h4071fa58, 32'h4230e10b, 32'h429b9a8a, 32'hc1079565, 32'h3f10f8e3, 32'hc2a1e815, 32'h42704729, 32'hc1a8e3f5};
test_output[4568] = '{32'h429b9a8a};
test_index[4568] = '{2};
test_input[36552:36559] = '{32'hc04b3fff, 32'hc1da616c, 32'hc2c1adc0, 32'hc1c570fd, 32'hc1f15bd0, 32'h41eadbb4, 32'hc2a6d935, 32'h4241edf1};
test_output[4569] = '{32'h4241edf1};
test_index[4569] = '{7};
test_input[36560:36567] = '{32'h4289f87a, 32'hc1c796bf, 32'h41597708, 32'hc209c081, 32'hc1c6f9ed, 32'hc0643ae4, 32'h41854dd8, 32'hc1908747};
test_output[4570] = '{32'h4289f87a};
test_index[4570] = '{0};
test_input[36568:36575] = '{32'h41f6009a, 32'hc04bc574, 32'h420afcf0, 32'h419bef72, 32'h42bb52df, 32'hc2b32d87, 32'h418849d6, 32'h42af5ea1};
test_output[4571] = '{32'h42bb52df};
test_index[4571] = '{4};
test_input[36576:36583] = '{32'h41d96105, 32'hc28d4a92, 32'h42ae6757, 32'h4292b86f, 32'hc2b98da2, 32'h41cdb1da, 32'hc060b2ae, 32'hc22bca26};
test_output[4572] = '{32'h42ae6757};
test_index[4572] = '{2};
test_input[36584:36591] = '{32'h4257d191, 32'hc0edead0, 32'h40419dcb, 32'h42085288, 32'hc26a0c2e, 32'hc2a6c0c3, 32'hc1b7e26f, 32'hc2c2f0b8};
test_output[4573] = '{32'h4257d191};
test_index[4573] = '{0};
test_input[36592:36599] = '{32'hc2bbc125, 32'hc11afdee, 32'h4123e25b, 32'h4130fbb7, 32'h42c46c3a, 32'h42099246, 32'hc2991e00, 32'h424c4c0d};
test_output[4574] = '{32'h42c46c3a};
test_index[4574] = '{4};
test_input[36600:36607] = '{32'hc21c6e23, 32'hc060dbb1, 32'hc2989374, 32'hc23bb1f7, 32'hc08421e6, 32'h42490370, 32'h425c93fe, 32'hc1c11dc8};
test_output[4575] = '{32'h425c93fe};
test_index[4575] = '{6};
test_input[36608:36615] = '{32'h41c32b38, 32'h4133cb83, 32'hc1b7479e, 32'hc28920cc, 32'h41416e28, 32'h423ca16a, 32'hc2c7c075, 32'h42adaf6e};
test_output[4576] = '{32'h42adaf6e};
test_index[4576] = '{7};
test_input[36616:36623] = '{32'h42a3ab0a, 32'h42900473, 32'h41f64e2e, 32'hc2647beb, 32'hc1f7345b, 32'h40819ae2, 32'h4286f3c2, 32'hc2bb8af2};
test_output[4577] = '{32'h42a3ab0a};
test_index[4577] = '{0};
test_input[36624:36631] = '{32'hbf7670df, 32'h4228e971, 32'h429c4fdb, 32'hc21c0185, 32'hc2bb43fc, 32'h42963a6d, 32'h4264dc6a, 32'hc14a4b78};
test_output[4578] = '{32'h429c4fdb};
test_index[4578] = '{2};
test_input[36632:36639] = '{32'hc263a21a, 32'hc2173b22, 32'h4005d365, 32'h418b0f7b, 32'hc21d180b, 32'hc0d7202c, 32'hc17f3872, 32'hc2575c70};
test_output[4579] = '{32'h418b0f7b};
test_index[4579] = '{3};
test_input[36640:36647] = '{32'hc245762a, 32'hc1ce394d, 32'hc297f2e4, 32'hc298c4b2, 32'h4192a4a9, 32'hc2974bf8, 32'h42961253, 32'h4222965a};
test_output[4580] = '{32'h42961253};
test_index[4580] = '{6};
test_input[36648:36655] = '{32'h426c184e, 32'h42587be8, 32'h41ca1023, 32'hc2b63f02, 32'h423a2806, 32'hc2c58492, 32'h41132de3, 32'h4294d9d2};
test_output[4581] = '{32'h4294d9d2};
test_index[4581] = '{7};
test_input[36656:36663] = '{32'hc0363d7b, 32'hc2a1ec5a, 32'hc283384b, 32'hc19f6188, 32'h428781e2, 32'hc27021c3, 32'hc2094232, 32'hc23caa17};
test_output[4582] = '{32'h428781e2};
test_index[4582] = '{4};
test_input[36664:36671] = '{32'h41b121e0, 32'hc2950c81, 32'hc2bc83bb, 32'hc2b60d17, 32'hbee2d649, 32'hc2a6737c, 32'hc2660a71, 32'h42877ae7};
test_output[4583] = '{32'h42877ae7};
test_index[4583] = '{7};
test_input[36672:36679] = '{32'h3feeff4e, 32'hc280f1b6, 32'hc24d4883, 32'h4288de0c, 32'hc27b1080, 32'h4298c85f, 32'h410208b7, 32'h423852ca};
test_output[4584] = '{32'h4298c85f};
test_index[4584] = '{5};
test_input[36680:36687] = '{32'h42026196, 32'h41d8c14b, 32'h422f4368, 32'hc22ddee8, 32'h427a0bc1, 32'hc1e554d6, 32'h42a1c39b, 32'h41807a95};
test_output[4585] = '{32'h42a1c39b};
test_index[4585] = '{6};
test_input[36688:36695] = '{32'h42b58193, 32'hc2b92d19, 32'hc0c613ad, 32'h42062f94, 32'hc2b4007f, 32'h42c1ba48, 32'hc2963bcd, 32'h42b181d1};
test_output[4586] = '{32'h42c1ba48};
test_index[4586] = '{5};
test_input[36696:36703] = '{32'h42c3445d, 32'h41ce5dc6, 32'h41bc616d, 32'h42555bb4, 32'hc245e652, 32'hc2b30774, 32'h42bc3c6c, 32'hc16f1310};
test_output[4587] = '{32'h42c3445d};
test_index[4587] = '{0};
test_input[36704:36711] = '{32'h42ae4d07, 32'hc2a26896, 32'h4057ffc1, 32'hc229b980, 32'hc25d2307, 32'hc2aa1408, 32'hc28c167f, 32'hc1e2c8af};
test_output[4588] = '{32'h42ae4d07};
test_index[4588] = '{0};
test_input[36712:36719] = '{32'h415fa04b, 32'h421279b9, 32'h426d5fa3, 32'h42c6c83b, 32'hc2626368, 32'hc1e5d7df, 32'h40fa8a39, 32'hc0fff587};
test_output[4589] = '{32'h42c6c83b};
test_index[4589] = '{3};
test_input[36720:36727] = '{32'h42854a5d, 32'h40afa262, 32'h3fc4cbf2, 32'hc1a56d89, 32'h423efcf5, 32'h41db6c69, 32'hc245e9d2, 32'h42190381};
test_output[4590] = '{32'h42854a5d};
test_index[4590] = '{0};
test_input[36728:36735] = '{32'h42b071df, 32'hc25babb1, 32'h4112473e, 32'h42a026da, 32'hc283f40e, 32'h42911158, 32'h42b65439, 32'hc2af6b81};
test_output[4591] = '{32'h42b65439};
test_index[4591] = '{6};
test_input[36736:36743] = '{32'hc25395d5, 32'h4260ad0d, 32'hc1d9511e, 32'h3feb78f0, 32'hc23ec88e, 32'hc1b66bda, 32'h3f03a93a, 32'hc1fad218};
test_output[4592] = '{32'h4260ad0d};
test_index[4592] = '{1};
test_input[36744:36751] = '{32'hc181bfce, 32'hc194cea5, 32'h41ceee1c, 32'hc2c453af, 32'hc27b15c5, 32'h427c7762, 32'h3ed74f78, 32'h424bfc6a};
test_output[4593] = '{32'h427c7762};
test_index[4593] = '{5};
test_input[36752:36759] = '{32'hc1f08a20, 32'hc2977198, 32'h41032118, 32'hc23d2acf, 32'hc2893241, 32'hc1e7c0d0, 32'hc1aaf606, 32'hc0bc9380};
test_output[4594] = '{32'h41032118};
test_index[4594] = '{2};
test_input[36760:36767] = '{32'hc2b34d7f, 32'hc27f0d6e, 32'h422a3427, 32'hc2b354ee, 32'hc1aa4e2b, 32'hc05ab147, 32'hc22749ba, 32'hc2984f91};
test_output[4595] = '{32'h422a3427};
test_index[4595] = '{2};
test_input[36768:36775] = '{32'h40ae4dd8, 32'hc24e0435, 32'hc032c665, 32'hc2681fcd, 32'h41369be8, 32'hc2034a4b, 32'h428e4065, 32'h41e27984};
test_output[4596] = '{32'h428e4065};
test_index[4596] = '{6};
test_input[36776:36783] = '{32'h418cbbab, 32'hc18f85c8, 32'h4298e4a3, 32'h42265f92, 32'hc21f0f2d, 32'hc267a4bd, 32'hc25e5182, 32'h428c818c};
test_output[4597] = '{32'h4298e4a3};
test_index[4597] = '{2};
test_input[36784:36791] = '{32'hc274cd60, 32'hc2c224dd, 32'hc292f224, 32'h41d4fdee, 32'h414bb8d3, 32'hc2975759, 32'hbfbfbbc7, 32'hc2c761ae};
test_output[4598] = '{32'h41d4fdee};
test_index[4598] = '{3};
test_input[36792:36799] = '{32'hc22b6a83, 32'h4221cede, 32'h428e26b5, 32'hc282631d, 32'hc200b3f6, 32'h42405e8b, 32'h427c0ae0, 32'hc2834117};
test_output[4599] = '{32'h428e26b5};
test_index[4599] = '{2};
test_input[36800:36807] = '{32'h42963dbd, 32'hc24611b8, 32'hc2aa83a0, 32'h41a12445, 32'hc2beefb2, 32'h421886f4, 32'hc1c45956, 32'hc2c18d15};
test_output[4600] = '{32'h42963dbd};
test_index[4600] = '{0};
test_input[36808:36815] = '{32'h4214a1ab, 32'hc15502f1, 32'hc1c31439, 32'hc1d1d69c, 32'h42afdb6a, 32'hc2bfc7f7, 32'h429df041, 32'hc28cf7d4};
test_output[4601] = '{32'h42afdb6a};
test_index[4601] = '{4};
test_input[36816:36823] = '{32'h40c4ba7c, 32'h41b64206, 32'h41aea903, 32'hc255978f, 32'hc1d18883, 32'h40ff9467, 32'h4283393e, 32'h41ae9236};
test_output[4602] = '{32'h4283393e};
test_index[4602] = '{6};
test_input[36824:36831] = '{32'h419e9761, 32'h42bc7356, 32'hc25179a5, 32'hc08ad233, 32'hc268d625, 32'hc1f42e22, 32'h42aaa1c0, 32'hc1c62e19};
test_output[4603] = '{32'h42bc7356};
test_index[4603] = '{1};
test_input[36832:36839] = '{32'hc28e029e, 32'hc1b9650e, 32'hc1afd779, 32'h41a1c7e5, 32'h42333007, 32'hc2a97027, 32'h42b29502, 32'h420e5fd7};
test_output[4604] = '{32'h42b29502};
test_index[4604] = '{6};
test_input[36840:36847] = '{32'hc1133901, 32'h420dcf81, 32'hc2549381, 32'h429df147, 32'hc290309f, 32'h419df15b, 32'hc2ba1eeb, 32'h415928e4};
test_output[4605] = '{32'h429df147};
test_index[4605] = '{3};
test_input[36848:36855] = '{32'h4282676f, 32'h41d2bc4e, 32'hc23c8c7c, 32'h404c9a30, 32'h41f15d67, 32'hc2b85f07, 32'hc2bf8c86, 32'hc2568742};
test_output[4606] = '{32'h4282676f};
test_index[4606] = '{0};
test_input[36856:36863] = '{32'hc178b965, 32'h42c2970d, 32'hc1fbea09, 32'h420b3799, 32'hc2820186, 32'hc162beb1, 32'h408f0e67, 32'h4291b8c6};
test_output[4607] = '{32'h42c2970d};
test_index[4607] = '{1};
test_input[36864:36871] = '{32'h41e55976, 32'hc192596d, 32'hc2a0cfb1, 32'hc09e115b, 32'h41556805, 32'h42bc3afe, 32'hc186d542, 32'hc286b0c6};
test_output[4608] = '{32'h42bc3afe};
test_index[4608] = '{5};
test_input[36872:36879] = '{32'h42738a0b, 32'hc2aac80e, 32'hc2193875, 32'h4000ee8d, 32'h41b2c5ab, 32'hc20e8df1, 32'hc2844ee8, 32'hc2763ada};
test_output[4609] = '{32'h42738a0b};
test_index[4609] = '{0};
test_input[36880:36887] = '{32'h42a0c336, 32'h41a18fd9, 32'h421b4505, 32'hc2963294, 32'hc2666f4a, 32'hc269f14b, 32'hc28f56d4, 32'hc2933070};
test_output[4610] = '{32'h42a0c336};
test_index[4610] = '{0};
test_input[36888:36895] = '{32'hc2c3b970, 32'hc2530e94, 32'h424eda9a, 32'h42998310, 32'h428bab4b, 32'hc21643dd, 32'hc2000d23, 32'h421815eb};
test_output[4611] = '{32'h42998310};
test_index[4611] = '{3};
test_input[36896:36903] = '{32'h42b1f807, 32'hc192ba83, 32'hbff361e3, 32'hc292a841, 32'hc22e7d62, 32'h413f5a4f, 32'hc24a12d0, 32'hc27f210a};
test_output[4612] = '{32'h42b1f807};
test_index[4612] = '{0};
test_input[36904:36911] = '{32'hc09c0808, 32'hc27cf98f, 32'h4266260b, 32'hc2a1218b, 32'hc246856f, 32'hc2ba18d6, 32'hc296fa79, 32'h40dd6185};
test_output[4613] = '{32'h4266260b};
test_index[4613] = '{2};
test_input[36912:36919] = '{32'hc050cf1f, 32'h42bac1ea, 32'h42ad8f90, 32'h4299e9c4, 32'h428fd01b, 32'h41c51d87, 32'hc2c56ca4, 32'h42032b53};
test_output[4614] = '{32'h42bac1ea};
test_index[4614] = '{1};
test_input[36920:36927] = '{32'hc1dcc187, 32'h41db5ed7, 32'h41c45045, 32'h421b23eb, 32'h415f97a9, 32'hc1ba5beb, 32'h4148da72, 32'hc2c74b64};
test_output[4615] = '{32'h421b23eb};
test_index[4615] = '{3};
test_input[36928:36935] = '{32'h427e0ace, 32'hc2961848, 32'hc02b9ef9, 32'h42670274, 32'h41acf25b, 32'hc11968e8, 32'hc1f8f6dd, 32'hc181023f};
test_output[4616] = '{32'h427e0ace};
test_index[4616] = '{0};
test_input[36936:36943] = '{32'h424153dc, 32'hc294102b, 32'hc2b58db6, 32'hc0ac44ce, 32'h413164b6, 32'h428216ed, 32'h422070bb, 32'h41749281};
test_output[4617] = '{32'h428216ed};
test_index[4617] = '{5};
test_input[36944:36951] = '{32'hc2ac56cc, 32'h42bd7974, 32'h42602138, 32'hc2b19801, 32'h428b2c2b, 32'h42b0bf52, 32'hbfb074f3, 32'h40b714b3};
test_output[4618] = '{32'h42bd7974};
test_index[4618] = '{1};
test_input[36952:36959] = '{32'hc2c4ff4e, 32'hc1f329e7, 32'hc2b373dd, 32'hc1b34a9c, 32'h42b31e4c, 32'h40fefefc, 32'h4152bde3, 32'hc284324e};
test_output[4619] = '{32'h42b31e4c};
test_index[4619] = '{4};
test_input[36960:36967] = '{32'hc201f9c0, 32'h4012f7c4, 32'hc20437b6, 32'hc16cb829, 32'h42b84491, 32'h427961db, 32'h3fd8fb94, 32'hc2387be9};
test_output[4620] = '{32'h42b84491};
test_index[4620] = '{4};
test_input[36968:36975] = '{32'hc2ba1157, 32'hc280ac49, 32'h41da3d15, 32'hc27fc8e3, 32'h427c20c9, 32'h418e13d4, 32'hc18724b1, 32'hc2451deb};
test_output[4621] = '{32'h427c20c9};
test_index[4621] = '{4};
test_input[36976:36983] = '{32'h425da17c, 32'h4115da36, 32'h42c4fb61, 32'hbe71179f, 32'h4299d0f3, 32'h41049023, 32'h42bafe11, 32'hc26a2171};
test_output[4622] = '{32'h42c4fb61};
test_index[4622] = '{2};
test_input[36984:36991] = '{32'h42a0e0d2, 32'h4216d29e, 32'h41bca538, 32'h4094fb29, 32'hc280ec80, 32'h42a251ed, 32'h4246af27, 32'hc1c5eef7};
test_output[4623] = '{32'h42a251ed};
test_index[4623] = '{5};
test_input[36992:36999] = '{32'h42141628, 32'h4213f35e, 32'hc2b26e76, 32'hc116bd97, 32'h4280c2b4, 32'hc2c38eae, 32'hc20a2e81, 32'hc261d714};
test_output[4624] = '{32'h4280c2b4};
test_index[4624] = '{4};
test_input[37000:37007] = '{32'h41f10242, 32'hc29e9914, 32'hc1dcb493, 32'hc1941a36, 32'h41fd2fe3, 32'h42b67dc8, 32'hc27d1a05, 32'hc2326cbd};
test_output[4625] = '{32'h42b67dc8};
test_index[4625] = '{5};
test_input[37008:37015] = '{32'h41e0eab0, 32'h4280fbee, 32'hc0f1d36c, 32'h41262adb, 32'h42365c1d, 32'hc2166421, 32'hc22781fc, 32'hc13c0e35};
test_output[4626] = '{32'h4280fbee};
test_index[4626] = '{1};
test_input[37016:37023] = '{32'h40e86567, 32'hc25e8cbf, 32'h3ea36b8f, 32'hc297f4f1, 32'hc2af22b8, 32'h4190f5bc, 32'h42c5e65c, 32'hc2979163};
test_output[4627] = '{32'h42c5e65c};
test_index[4627] = '{6};
test_input[37024:37031] = '{32'hc2750495, 32'hc0e85907, 32'h42b9390d, 32'h420d799f, 32'h4284046a, 32'hc18938e8, 32'hc289f6cf, 32'hc104ee02};
test_output[4628] = '{32'h42b9390d};
test_index[4628] = '{2};
test_input[37032:37039] = '{32'h422b0588, 32'hbd9810f4, 32'h41f504c7, 32'hc238b400, 32'hc24776fd, 32'h4275033a, 32'h42c054d8, 32'h4178b2fa};
test_output[4629] = '{32'h42c054d8};
test_index[4629] = '{6};
test_input[37040:37047] = '{32'h427b6702, 32'h4292bac3, 32'h4146b121, 32'hc0d7d0ee, 32'h427e800d, 32'h42089a9a, 32'hc2b8a3bd, 32'h41341680};
test_output[4630] = '{32'h4292bac3};
test_index[4630] = '{1};
test_input[37048:37055] = '{32'hc1cca804, 32'hc2a4701d, 32'hc297880b, 32'hc067bae7, 32'h4270d944, 32'h42b79ede, 32'hc1f9e024, 32'hc2b34a7a};
test_output[4631] = '{32'h42b79ede};
test_index[4631] = '{5};
test_input[37056:37063] = '{32'hc1aa1c13, 32'h420c69cb, 32'hc2b4cfa3, 32'h422420b0, 32'hc2a5d954, 32'h42a16d7a, 32'hc2bb0aa1, 32'hc281ee5b};
test_output[4632] = '{32'h42a16d7a};
test_index[4632] = '{5};
test_input[37064:37071] = '{32'hc29151a7, 32'h422c0131, 32'h42b29d9f, 32'h41650f4b, 32'h41cb714d, 32'hc2ade128, 32'h428b5405, 32'h42b2f237};
test_output[4633] = '{32'h42b2f237};
test_index[4633] = '{7};
test_input[37072:37079] = '{32'hc15528e7, 32'hc1a58be7, 32'hc08a9110, 32'h427205ae, 32'hc190df76, 32'hc2a4d79f, 32'hc28e7266, 32'hc20a7eba};
test_output[4634] = '{32'h427205ae};
test_index[4634] = '{3};
test_input[37080:37087] = '{32'hc2a38b54, 32'h42b02b7f, 32'h41b16cfe, 32'h4222fec5, 32'h42517410, 32'h42ab3cb1, 32'h42b1031e, 32'hc18e3dfd};
test_output[4635] = '{32'h42b1031e};
test_index[4635] = '{6};
test_input[37088:37095] = '{32'h421ea682, 32'h41256127, 32'h4290e294, 32'hc19ed5bf, 32'h423dca73, 32'hc2288639, 32'hc1c71a2b, 32'h41c7a5fd};
test_output[4636] = '{32'h4290e294};
test_index[4636] = '{2};
test_input[37096:37103] = '{32'h42bbb273, 32'h4291490a, 32'h42b42cd6, 32'hc271c0ef, 32'hc1e6888f, 32'hc25783a2, 32'hc23f319d, 32'h42b9afe6};
test_output[4637] = '{32'h42bbb273};
test_index[4637] = '{0};
test_input[37104:37111] = '{32'hc20f3d68, 32'h42ad0391, 32'h4297d48d, 32'hc0c50819, 32'h410a1696, 32'h42459ff0, 32'h3f37457c, 32'hc202f438};
test_output[4638] = '{32'h42ad0391};
test_index[4638] = '{1};
test_input[37112:37119] = '{32'h42150d6a, 32'hc1cfac43, 32'hc0ac8e96, 32'h42ad64af, 32'h428c7da2, 32'hc28f8b6d, 32'h4292f3e4, 32'h41cf414b};
test_output[4639] = '{32'h42ad64af};
test_index[4639] = '{3};
test_input[37120:37127] = '{32'h428cfd22, 32'h421ecf61, 32'h4204005f, 32'hc1f86596, 32'h427b06c1, 32'h427e4742, 32'hc20fe9e3, 32'hc2c215fe};
test_output[4640] = '{32'h428cfd22};
test_index[4640] = '{0};
test_input[37128:37135] = '{32'hc1794752, 32'h42be0daa, 32'hc29f6540, 32'h419e0446, 32'h41bae660, 32'h42627eee, 32'hc284df23, 32'hc20b9ec4};
test_output[4641] = '{32'h42be0daa};
test_index[4641] = '{1};
test_input[37136:37143] = '{32'h421112bc, 32'hc1d70eef, 32'hc1948e68, 32'h42afd4a8, 32'hc03e7e45, 32'h4272b96f, 32'hc28896eb, 32'hc2bb3908};
test_output[4642] = '{32'h42afd4a8};
test_index[4642] = '{3};
test_input[37144:37151] = '{32'hc27296be, 32'hc1ce9b37, 32'h41d01dad, 32'hc21ccc3d, 32'h4296ef3f, 32'hc1abf4e7, 32'hc2285a30, 32'hc257ead8};
test_output[4643] = '{32'h4296ef3f};
test_index[4643] = '{4};
test_input[37152:37159] = '{32'h41420267, 32'hc070f06e, 32'h42a49ccb, 32'h428bb9cf, 32'h4232aee4, 32'hc2586c4a, 32'h4164bddc, 32'h40fc4b06};
test_output[4644] = '{32'h42a49ccb};
test_index[4644] = '{2};
test_input[37160:37167] = '{32'hc26c725d, 32'h418ca25d, 32'h41d4dcb3, 32'hc1ad6c05, 32'hc09d7185, 32'h429ddfe4, 32'hc1c17af0, 32'hc259af32};
test_output[4645] = '{32'h429ddfe4};
test_index[4645] = '{5};
test_input[37168:37175] = '{32'h421a2416, 32'h41d6ed0a, 32'hc2bcd3e2, 32'hc261d5b3, 32'h42ab61a6, 32'h42099dc4, 32'h4221febd, 32'h422e3138};
test_output[4646] = '{32'h42ab61a6};
test_index[4646] = '{4};
test_input[37176:37183] = '{32'h42abe5a3, 32'h41ed94f3, 32'hc201936d, 32'h42959870, 32'hc2a61469, 32'hc27fc76b, 32'hc005542c, 32'h42c4d6f3};
test_output[4647] = '{32'h42c4d6f3};
test_index[4647] = '{7};
test_input[37184:37191] = '{32'h426d3832, 32'h42c61e06, 32'hc0f0f98b, 32'h420efd4d, 32'hc289d23e, 32'h42bc2632, 32'h42b295ba, 32'h4116a227};
test_output[4648] = '{32'h42c61e06};
test_index[4648] = '{1};
test_input[37192:37199] = '{32'hc1982023, 32'h41f2cfff, 32'hc19a4071, 32'h4219354a, 32'hc1c4fd90, 32'h40d9eda8, 32'hc2376a02, 32'hc249ec96};
test_output[4649] = '{32'h4219354a};
test_index[4649] = '{3};
test_input[37200:37207] = '{32'hc2094e11, 32'h42c37f23, 32'h42493ce4, 32'h4270835c, 32'h4241285c, 32'hc2b7890e, 32'h42be5fb6, 32'hc28d72bb};
test_output[4650] = '{32'h42c37f23};
test_index[4650] = '{1};
test_input[37208:37215] = '{32'hc186ca63, 32'hc18a5018, 32'hc16de114, 32'h4282bcbf, 32'h419a6124, 32'h4123c49a, 32'hc21da982, 32'hc2415577};
test_output[4651] = '{32'h4282bcbf};
test_index[4651] = '{3};
test_input[37216:37223] = '{32'hc18866b4, 32'hc242bfeb, 32'hc21c9371, 32'hc2b9a235, 32'h42704ff5, 32'h42b600e4, 32'hc224cda9, 32'h423fc315};
test_output[4652] = '{32'h42b600e4};
test_index[4652] = '{5};
test_input[37224:37231] = '{32'hc2abcb21, 32'hc1da03df, 32'hc28a4b4f, 32'h42489f90, 32'hc2b67353, 32'h42b602c7, 32'h428c640a, 32'hc1cf824c};
test_output[4653] = '{32'h42b602c7};
test_index[4653] = '{5};
test_input[37232:37239] = '{32'hc281501c, 32'h4200166c, 32'h422f6ee2, 32'h4275de32, 32'hc29eec58, 32'hc18a2884, 32'h41cf63c7, 32'hc254d8fd};
test_output[4654] = '{32'h4275de32};
test_index[4654] = '{3};
test_input[37240:37247] = '{32'h426c8e46, 32'h411d79f0, 32'h412a3881, 32'hc2829da0, 32'h42a6e43d, 32'hc1d2618a, 32'hc29c7c03, 32'hbdcb7a40};
test_output[4655] = '{32'h42a6e43d};
test_index[4655] = '{4};
test_input[37248:37255] = '{32'hc284432d, 32'h426d1037, 32'hc0c664e0, 32'h42c6105b, 32'hc2c24e75, 32'hc107aa05, 32'h428aa3c0, 32'hc2a7ada3};
test_output[4656] = '{32'h42c6105b};
test_index[4656] = '{3};
test_input[37256:37263] = '{32'hc1706626, 32'hc1d29724, 32'hc22aeba1, 32'h427b72f1, 32'hc257a8a6, 32'h4256921c, 32'h4240b07e, 32'h415aeef7};
test_output[4657] = '{32'h427b72f1};
test_index[4657] = '{3};
test_input[37264:37271] = '{32'hc1e61b0b, 32'hc2b1cb87, 32'hc2930589, 32'h402730f1, 32'h4288ae4b, 32'hc28a7382, 32'h3f4b4d8a, 32'h42b24341};
test_output[4658] = '{32'h42b24341};
test_index[4658] = '{7};
test_input[37272:37279] = '{32'h42accaf2, 32'hc21ed70f, 32'hc217d5c7, 32'h42b19f25, 32'hc2c4d0f9, 32'hc19b9b4a, 32'h419d7765, 32'h428fc0b3};
test_output[4659] = '{32'h42b19f25};
test_index[4659] = '{3};
test_input[37280:37287] = '{32'hc2797262, 32'h42b86080, 32'h4196acd1, 32'hc277326b, 32'h42bd381a, 32'h420d16a9, 32'h41ad534e, 32'h41de9035};
test_output[4660] = '{32'h42bd381a};
test_index[4660] = '{4};
test_input[37288:37295] = '{32'hc265322e, 32'h421fb7d4, 32'h41f94cd3, 32'hc21cd2dd, 32'hc1f7b0d7, 32'h429bae40, 32'hc29ec584, 32'h429d7096};
test_output[4661] = '{32'h429d7096};
test_index[4661] = '{7};
test_input[37296:37303] = '{32'hc25440d9, 32'h42c31a82, 32'hc2a84639, 32'h4278e04e, 32'hc29c6e0b, 32'hc2779da6, 32'h42c239e1, 32'h425285c7};
test_output[4662] = '{32'h42c31a82};
test_index[4662] = '{1};
test_input[37304:37311] = '{32'h418f86e8, 32'hc24391db, 32'h42828964, 32'h41cec2f8, 32'hc2003312, 32'hc2c1e7dc, 32'h4285093a, 32'hc1e0dace};
test_output[4663] = '{32'h4285093a};
test_index[4663] = '{6};
test_input[37312:37319] = '{32'hc29fc47c, 32'hc12afc95, 32'hc2b75f1e, 32'h429679cd, 32'h420bed97, 32'h42a52495, 32'hc210c076, 32'hc26da049};
test_output[4664] = '{32'h42a52495};
test_index[4664] = '{5};
test_input[37320:37327] = '{32'h42859661, 32'h423205ed, 32'hc16fc61d, 32'hc2a8a06d, 32'hc28d87e4, 32'hc2a018d0, 32'hc2c30387, 32'hc2579966};
test_output[4665] = '{32'h42859661};
test_index[4665] = '{0};
test_input[37328:37335] = '{32'h42bae4fd, 32'hc221f71f, 32'h40c06085, 32'h42b98b38, 32'h42b99692, 32'h40de1f91, 32'hc24cdc26, 32'h42807111};
test_output[4666] = '{32'h42bae4fd};
test_index[4666] = '{0};
test_input[37336:37343] = '{32'h4204ed72, 32'hc2301e75, 32'h427cd9bc, 32'hc29473b3, 32'hc28e03d5, 32'h42b41fcf, 32'hc29a10e7, 32'h4277c1e9};
test_output[4667] = '{32'h42b41fcf};
test_index[4667] = '{5};
test_input[37344:37351] = '{32'h427cdab9, 32'hc2bded83, 32'hc2036dd2, 32'hc293ab00, 32'h4240cba4, 32'h42920ca5, 32'h403bae21, 32'h429af834};
test_output[4668] = '{32'h429af834};
test_index[4668] = '{7};
test_input[37352:37359] = '{32'h41b750b6, 32'h42b977ba, 32'h42284297, 32'hc2268bfc, 32'hc277b149, 32'h41ad9b1d, 32'hc1db8417, 32'h416f7ac4};
test_output[4669] = '{32'h42b977ba};
test_index[4669] = '{1};
test_input[37360:37367] = '{32'hc2afa3b0, 32'hc289dcc0, 32'h413142ae, 32'hc14bff72, 32'hc2ab81a4, 32'h428d28a5, 32'hc2846c85, 32'h42957f9a};
test_output[4670] = '{32'h42957f9a};
test_index[4670] = '{7};
test_input[37368:37375] = '{32'hc2274d3a, 32'h4203bfec, 32'h42195762, 32'hc2bfbd06, 32'h41a4c768, 32'hc2c7fce5, 32'hc1d19d0b, 32'h4293a8e4};
test_output[4671] = '{32'h4293a8e4};
test_index[4671] = '{7};
test_input[37376:37383] = '{32'hc1d152a1, 32'h41496179, 32'h42a69ca8, 32'h42853c96, 32'h42381515, 32'hc1769f93, 32'h4189064a, 32'h424cef48};
test_output[4672] = '{32'h42a69ca8};
test_index[4672] = '{2};
test_input[37384:37391] = '{32'h429315a1, 32'hc1e3d01e, 32'h41779e33, 32'hc2a5f898, 32'hc256d015, 32'h4188c2d0, 32'h40ec2357, 32'hc2b8fd1b};
test_output[4673] = '{32'h429315a1};
test_index[4673] = '{0};
test_input[37392:37399] = '{32'h42b56f1b, 32'h42ab8705, 32'h4273e256, 32'hc289865c, 32'hc2c05937, 32'hc2a13275, 32'hc23e2f73, 32'h42130561};
test_output[4674] = '{32'h42b56f1b};
test_index[4674] = '{0};
test_input[37400:37407] = '{32'hc23973d5, 32'hc112dfac, 32'h425428e1, 32'hc21561fa, 32'h42871b13, 32'hc213539f, 32'h42bb5a9d, 32'h4276d34d};
test_output[4675] = '{32'h42bb5a9d};
test_index[4675] = '{6};
test_input[37408:37415] = '{32'hc25b63d0, 32'hc2699fbd, 32'hc2bfde2f, 32'hc298e071, 32'hc1c45728, 32'hc27cbf6b, 32'h417e79e4, 32'hc12ea9d2};
test_output[4676] = '{32'h417e79e4};
test_index[4676] = '{6};
test_input[37416:37423] = '{32'h421a126c, 32'hc291de37, 32'h423d5553, 32'h4228156f, 32'hc2138ad9, 32'h4295e6e5, 32'h421a482e, 32'hc1de3cd9};
test_output[4677] = '{32'h4295e6e5};
test_index[4677] = '{5};
test_input[37424:37431] = '{32'hc2b2bd7b, 32'h429ca453, 32'h42b9eda3, 32'hc06a1c41, 32'h4280e1fb, 32'hc2997e51, 32'hc2ab6732, 32'hc25128da};
test_output[4678] = '{32'h42b9eda3};
test_index[4678] = '{2};
test_input[37432:37439] = '{32'h42a03ecc, 32'h422d513d, 32'hc2c5e047, 32'h42b5a5be, 32'h4261b529, 32'h422a4288, 32'h423dfe4b, 32'hc0a93ca8};
test_output[4679] = '{32'h42b5a5be};
test_index[4679] = '{3};
test_input[37440:37447] = '{32'h420fb7ed, 32'h4101d217, 32'hc28dd0c0, 32'hc261192b, 32'h41ab0e7a, 32'h420eb806, 32'h418b5faa, 32'hc19fb636};
test_output[4680] = '{32'h420fb7ed};
test_index[4680] = '{0};
test_input[37448:37455] = '{32'h4278bbed, 32'hc2b6e0d9, 32'hc265c73c, 32'hc2a4dd00, 32'hc24b4f44, 32'h418b6e1d, 32'hc2b61268, 32'hc18f8aa1};
test_output[4681] = '{32'h4278bbed};
test_index[4681] = '{0};
test_input[37456:37463] = '{32'h428f8418, 32'h4253a1a9, 32'hc1ebef92, 32'h41cea9fc, 32'h424cc4cc, 32'hc23d0ce8, 32'hc2ad619b, 32'hc15b7346};
test_output[4682] = '{32'h428f8418};
test_index[4682] = '{0};
test_input[37464:37471] = '{32'h42b93cac, 32'h422e8727, 32'hc27b3140, 32'hc20803e8, 32'h425f97f2, 32'h42831a73, 32'hc2994717, 32'h42c52233};
test_output[4683] = '{32'h42c52233};
test_index[4683] = '{7};
test_input[37472:37479] = '{32'h423cdb0f, 32'h42773728, 32'h41d7c898, 32'hc2aeada3, 32'h42a9a1df, 32'hc18d86ce, 32'hc1f25a2b, 32'h42c3c520};
test_output[4684] = '{32'h42c3c520};
test_index[4684] = '{7};
test_input[37480:37487] = '{32'h4291ed0c, 32'h42a39d50, 32'h42098a54, 32'h426ab2ca, 32'hc0d32fc3, 32'hc18964fa, 32'hc2a07c9a, 32'h42c70ea0};
test_output[4685] = '{32'h42c70ea0};
test_index[4685] = '{7};
test_input[37488:37495] = '{32'h423415e6, 32'h40ae36fd, 32'h42732805, 32'h42b5901c, 32'hc260e802, 32'h427e33cf, 32'hc22621f8, 32'h423a5b05};
test_output[4686] = '{32'h42b5901c};
test_index[4686] = '{3};
test_input[37496:37503] = '{32'h425c59b7, 32'hc2414089, 32'h42093abe, 32'hbff0496e, 32'h4163a3e3, 32'hc1909769, 32'hc2c74c38, 32'h41a5110c};
test_output[4687] = '{32'h425c59b7};
test_index[4687] = '{0};
test_input[37504:37511] = '{32'hc293e573, 32'h4280e52a, 32'h42a0e601, 32'h42965164, 32'h42c655e2, 32'h428abf85, 32'hc24be25f, 32'h42c30f54};
test_output[4688] = '{32'h42c655e2};
test_index[4688] = '{4};
test_input[37512:37519] = '{32'hc21cb681, 32'h416315f5, 32'h41890d68, 32'hc196c462, 32'h42a44c29, 32'h41d195d4, 32'h42295642, 32'h42a9c1c0};
test_output[4689] = '{32'h42a9c1c0};
test_index[4689] = '{7};
test_input[37520:37527] = '{32'h420a54b6, 32'hc255d4c5, 32'h42b46297, 32'h42bfb98f, 32'h41a01859, 32'hc217f140, 32'hc2452c0f, 32'hc2700bf5};
test_output[4690] = '{32'h42bfb98f};
test_index[4690] = '{3};
test_input[37528:37535] = '{32'hc2662a4b, 32'h426ada68, 32'hc2ae710b, 32'hc2021bf2, 32'hc24b9775, 32'hc0e0b771, 32'h42474953, 32'hc21f207e};
test_output[4691] = '{32'h426ada68};
test_index[4691] = '{1};
test_input[37536:37543] = '{32'hc11e8381, 32'hc0a1ac96, 32'h42ab3870, 32'h41fe66ef, 32'h42a4e3a1, 32'h41a2b1ef, 32'hc27e9955, 32'hc2881977};
test_output[4692] = '{32'h42ab3870};
test_index[4692] = '{2};
test_input[37544:37551] = '{32'hc278245f, 32'h42a72199, 32'h42288a56, 32'h42b3ddff, 32'hc1e7c1f6, 32'h42a34758, 32'hc28e0fe7, 32'hc11d8731};
test_output[4693] = '{32'h42b3ddff};
test_index[4693] = '{3};
test_input[37552:37559] = '{32'hc1ea1cff, 32'h42bb1dbb, 32'hc213720c, 32'hc295b489, 32'h42332d48, 32'h4220dd08, 32'h411d2116, 32'h428a57b2};
test_output[4694] = '{32'h42bb1dbb};
test_index[4694] = '{1};
test_input[37560:37567] = '{32'h418519c7, 32'h413d05b4, 32'hc2a15726, 32'h411cad25, 32'h42224285, 32'h41c291cc, 32'hc1ad8e93, 32'h4250f68c};
test_output[4695] = '{32'h4250f68c};
test_index[4695] = '{7};
test_input[37568:37575] = '{32'hc2912baf, 32'h42130832, 32'hc2846067, 32'h42033db6, 32'hc226ee75, 32'hc1e79ec5, 32'h4168c6f3, 32'h41b29789};
test_output[4696] = '{32'h42130832};
test_index[4696] = '{1};
test_input[37576:37583] = '{32'hc2759466, 32'hc291743b, 32'hc26b9073, 32'hc2852a28, 32'h426de66e, 32'hc0c6de6f, 32'hc1d5b64a, 32'h4215a919};
test_output[4697] = '{32'h426de66e};
test_index[4697] = '{4};
test_input[37584:37591] = '{32'h42b84814, 32'hc13b8583, 32'hc2935373, 32'h415ebe30, 32'h42bca689, 32'h41e58778, 32'h42a54e33, 32'hc26f314f};
test_output[4698] = '{32'h42bca689};
test_index[4698] = '{4};
test_input[37592:37599] = '{32'hc2b26d3c, 32'h42103329, 32'hc2796d5b, 32'h41dbc280, 32'hc2c16d86, 32'h42bc02e1, 32'h427b9095, 32'hc2aab05f};
test_output[4699] = '{32'h42bc02e1};
test_index[4699] = '{5};
test_input[37600:37607] = '{32'hc08763f9, 32'h42a9fea7, 32'h428aff89, 32'h427fe106, 32'hc0c0ca45, 32'h422b8a1d, 32'hc28b801a, 32'h40f39cc1};
test_output[4700] = '{32'h42a9fea7};
test_index[4700] = '{1};
test_input[37608:37615] = '{32'h40ffe25f, 32'hc1e3a91f, 32'hc285c372, 32'h41385060, 32'h4243ed1f, 32'hc2683200, 32'hc199f388, 32'h41a57ef6};
test_output[4701] = '{32'h4243ed1f};
test_index[4701] = '{4};
test_input[37616:37623] = '{32'h4119e110, 32'h41debc15, 32'h429c0d2f, 32'hc2143d05, 32'hc1f44a80, 32'hc2c29fce, 32'h428021a4, 32'hc29132dc};
test_output[4702] = '{32'h429c0d2f};
test_index[4702] = '{2};
test_input[37624:37631] = '{32'h40ccde19, 32'hc256417c, 32'h42194827, 32'h42a0e5aa, 32'hc13dbe0b, 32'hc29062d6, 32'h4156fa00, 32'h418ce684};
test_output[4703] = '{32'h42a0e5aa};
test_index[4703] = '{3};
test_input[37632:37639] = '{32'h423f748e, 32'h42042666, 32'h4282b407, 32'hc190c092, 32'hc24616ff, 32'hc29d6ae1, 32'hc21ba6b5, 32'h4237482b};
test_output[4704] = '{32'h4282b407};
test_index[4704] = '{2};
test_input[37640:37647] = '{32'h420b9228, 32'h41caeb55, 32'hc23ceb7a, 32'h422b3acf, 32'h428cee15, 32'hc2af272b, 32'h41d722ea, 32'h42858d51};
test_output[4705] = '{32'h428cee15};
test_index[4705] = '{4};
test_input[37648:37655] = '{32'h401f4bfc, 32'h41a96ece, 32'hc260eeb2, 32'h428766da, 32'h42b4fa02, 32'h429f0cd7, 32'hc040eca5, 32'hc2bf89f2};
test_output[4706] = '{32'h42b4fa02};
test_index[4706] = '{4};
test_input[37656:37663] = '{32'h425d9ec5, 32'hc2a24889, 32'hc280babb, 32'hc080e800, 32'h41b191b4, 32'h42869f34, 32'h41999854, 32'hc2453afa};
test_output[4707] = '{32'h42869f34};
test_index[4707] = '{5};
test_input[37664:37671] = '{32'h3e1e7f0c, 32'hc1db3bbc, 32'h42bf6968, 32'hc1b60367, 32'h4220386e, 32'h427a6195, 32'hc1815c0b, 32'hc266c38a};
test_output[4708] = '{32'h42bf6968};
test_index[4708] = '{2};
test_input[37672:37679] = '{32'hc1be24f0, 32'hc2adf69d, 32'h42bd6f45, 32'h423590a8, 32'hc2c525a4, 32'h41796015, 32'h4266a41a, 32'hc2a0b225};
test_output[4709] = '{32'h42bd6f45};
test_index[4709] = '{2};
test_input[37680:37687] = '{32'h42ace71d, 32'h4018f2b0, 32'hc112a9e7, 32'h42391ff5, 32'hc1924d84, 32'hc193a1ad, 32'hc1a25257, 32'h41bd67ce};
test_output[4710] = '{32'h42ace71d};
test_index[4710] = '{0};
test_input[37688:37695] = '{32'h42b46963, 32'h41944a89, 32'h3f02807f, 32'h421a7f5b, 32'hc1493b0f, 32'h428154af, 32'h414290dc, 32'h42887fe5};
test_output[4711] = '{32'h42b46963};
test_index[4711] = '{0};
test_input[37696:37703] = '{32'h42429ea6, 32'hc25b2446, 32'hc2546028, 32'h4297f46b, 32'h42593daf, 32'h3e20560e, 32'hc109f48e, 32'hc1e9b505};
test_output[4712] = '{32'h4297f46b};
test_index[4712] = '{3};
test_input[37704:37711] = '{32'hc1b6dcb4, 32'hc2958efa, 32'hc28fbb0a, 32'hc223333a, 32'hc286f3b2, 32'h4062b419, 32'h42a99314, 32'hc258461b};
test_output[4713] = '{32'h42a99314};
test_index[4713] = '{6};
test_input[37712:37719] = '{32'h423414d9, 32'h41f9338e, 32'hc28d3550, 32'h40a5a34c, 32'h4276a6a2, 32'hc1d4cf54, 32'hc17fa9f9, 32'h42c0f674};
test_output[4714] = '{32'h42c0f674};
test_index[4714] = '{7};
test_input[37720:37727] = '{32'h4286818c, 32'h422846b1, 32'hc297fe39, 32'hc1b9dc71, 32'hc1f6c051, 32'h4299e3d7, 32'hc15105f9, 32'h41ae5bd8};
test_output[4715] = '{32'h4299e3d7};
test_index[4715] = '{5};
test_input[37728:37735] = '{32'hc2008fd1, 32'h429fcef4, 32'hc1fb8fa7, 32'h40df1b65, 32'hc0f6dea5, 32'h42acee95, 32'h422c2b35, 32'h41014969};
test_output[4716] = '{32'h42acee95};
test_index[4716] = '{5};
test_input[37736:37743] = '{32'h42a1d576, 32'h42bcd8df, 32'hc1606f6d, 32'hc2ba690c, 32'h429a4072, 32'hc1ec0c42, 32'hc23f2e94, 32'hc2b50686};
test_output[4717] = '{32'h42bcd8df};
test_index[4717] = '{1};
test_input[37744:37751] = '{32'hc27c9b25, 32'h42217e2d, 32'hc2079432, 32'h429c6d81, 32'h40a0a817, 32'h428d1580, 32'hc280027d, 32'h4252e630};
test_output[4718] = '{32'h429c6d81};
test_index[4718] = '{3};
test_input[37752:37759] = '{32'hc2a2daa7, 32'hc224f315, 32'hc266bbc7, 32'hc2366c8c, 32'h429dea55, 32'h416634ab, 32'hc286ab09, 32'hc2855b45};
test_output[4719] = '{32'h429dea55};
test_index[4719] = '{4};
test_input[37760:37767] = '{32'hc075086b, 32'h4227b50e, 32'h428c4b3b, 32'h4291781b, 32'h42ab19d5, 32'hc119268d, 32'h4246bbeb, 32'hc0f674d0};
test_output[4720] = '{32'h42ab19d5};
test_index[4720] = '{4};
test_input[37768:37775] = '{32'h42b47518, 32'h42728e39, 32'h40c819bb, 32'hc1b7954c, 32'h3fb66112, 32'hc28f1d1b, 32'h4238a0a1, 32'h42a3dec9};
test_output[4721] = '{32'h42b47518};
test_index[4721] = '{0};
test_input[37776:37783] = '{32'hc299120a, 32'h4262cc95, 32'h42c5f646, 32'hc2abf944, 32'hc24e1bc0, 32'hc2b2e233, 32'hc098ae1f, 32'hc1f4844f};
test_output[4722] = '{32'h42c5f646};
test_index[4722] = '{2};
test_input[37784:37791] = '{32'hc12af797, 32'h4273c885, 32'h41a95c1a, 32'h42a207ff, 32'h428dcf80, 32'hc191dcb4, 32'h429402e2, 32'h42855f73};
test_output[4723] = '{32'h42a207ff};
test_index[4723] = '{3};
test_input[37792:37799] = '{32'hc1073c1e, 32'h41e3f0e5, 32'hc2646799, 32'hc1548c99, 32'h41cb566e, 32'hc2166647, 32'h4292f16d, 32'hc281d6fe};
test_output[4724] = '{32'h4292f16d};
test_index[4724] = '{6};
test_input[37800:37807] = '{32'hc11006ba, 32'h40c6b62d, 32'h4277f804, 32'h42419809, 32'h4296e63e, 32'h41c32433, 32'hc212b7cf, 32'h4270c515};
test_output[4725] = '{32'h4296e63e};
test_index[4725] = '{4};
test_input[37808:37815] = '{32'h4043f8b2, 32'h42c499a4, 32'h402356a5, 32'h41a630fd, 32'hc2828dcd, 32'h42144591, 32'hc095fe2f, 32'hc22f1836};
test_output[4726] = '{32'h42c499a4};
test_index[4726] = '{1};
test_input[37816:37823] = '{32'h42a8885e, 32'hc1ef72db, 32'h42a4a359, 32'h427adc01, 32'hc187b580, 32'h41128876, 32'hc0ce86c1, 32'hc1d5e2be};
test_output[4727] = '{32'h42a8885e};
test_index[4727] = '{0};
test_input[37824:37831] = '{32'hc1aaa79b, 32'h42aca59e, 32'h41a0ec08, 32'hc1a5d4a6, 32'hc0c35902, 32'hc1ed28a3, 32'h42498240, 32'h42a42ea9};
test_output[4728] = '{32'h42aca59e};
test_index[4728] = '{1};
test_input[37832:37839] = '{32'h427ea9aa, 32'h41121aec, 32'hc26463e9, 32'hc1dba614, 32'h42346987, 32'h420d8bf2, 32'hc2a039b4, 32'h42074da3};
test_output[4729] = '{32'h427ea9aa};
test_index[4729] = '{0};
test_input[37840:37847] = '{32'hbf95ae83, 32'hc25c2c19, 32'h420a8c06, 32'hbe8a454f, 32'h42a83e44, 32'hc2bc195d, 32'h42044c65, 32'hc1e6dec6};
test_output[4730] = '{32'h42a83e44};
test_index[4730] = '{4};
test_input[37848:37855] = '{32'hc256ab35, 32'h41e8aea8, 32'h42c13d43, 32'h4246bff8, 32'h421e8671, 32'h42bac154, 32'hc0197289, 32'h4067dc42};
test_output[4731] = '{32'h42c13d43};
test_index[4731] = '{2};
test_input[37856:37863] = '{32'h40f29d4d, 32'hc1ba8ee4, 32'hc2aca322, 32'hc2b20db9, 32'hc267df54, 32'hc2c554df, 32'h42999edf, 32'h428edd63};
test_output[4732] = '{32'h42999edf};
test_index[4732] = '{6};
test_input[37864:37871] = '{32'h42b140a4, 32'hc29af68d, 32'hc21ddfe7, 32'hc28f4326, 32'hc2bfa8b9, 32'h41a4a449, 32'hc26e0164, 32'hc29d53a1};
test_output[4733] = '{32'h42b140a4};
test_index[4733] = '{0};
test_input[37872:37879] = '{32'h41b96e6d, 32'h41e035c7, 32'hc284204f, 32'h422d96fc, 32'h40edae92, 32'hc2ba166f, 32'h421f0705, 32'hc290b582};
test_output[4734] = '{32'h422d96fc};
test_index[4734] = '{3};
test_input[37880:37887] = '{32'h4297da9f, 32'hc1606ad1, 32'h4286d8cf, 32'h426c0e3e, 32'hc25bcc9d, 32'hc02c79a1, 32'h40a5d29e, 32'h42842370};
test_output[4735] = '{32'h4297da9f};
test_index[4735] = '{0};
test_input[37888:37895] = '{32'h417f2f08, 32'h429f8126, 32'hc28569a9, 32'h423bae7a, 32'h4289cb8f, 32'h4236d79f, 32'h41bb08ff, 32'h416ef465};
test_output[4736] = '{32'h429f8126};
test_index[4736] = '{1};
test_input[37896:37903] = '{32'hc1d77906, 32'hc2964d9f, 32'hc2b5ffec, 32'h42521691, 32'hc2c745a6, 32'hc04f240f, 32'hc10c3628, 32'hc2907695};
test_output[4737] = '{32'h42521691};
test_index[4737] = '{3};
test_input[37904:37911] = '{32'hc185f265, 32'hc2238ca6, 32'h42bda500, 32'h41dafd60, 32'h41a44838, 32'h429f0538, 32'h4197e8e6, 32'hc2c22733};
test_output[4738] = '{32'h42bda500};
test_index[4738] = '{2};
test_input[37912:37919] = '{32'hc22fac48, 32'hc1f54ae4, 32'h421f3f7f, 32'h42a0d854, 32'hc22428d0, 32'h42a0a150, 32'h41ca64ad, 32'hc2be6bdd};
test_output[4739] = '{32'h42a0d854};
test_index[4739] = '{3};
test_input[37920:37927] = '{32'hc2b5ca7d, 32'h42bdf296, 32'hc19b926c, 32'hc1eeb3db, 32'hc2674d5a, 32'h40f951b8, 32'hc271ff93, 32'hc23195c4};
test_output[4740] = '{32'h42bdf296};
test_index[4740] = '{1};
test_input[37928:37935] = '{32'h42a10c82, 32'h42886dec, 32'h420dd263, 32'hc2bcbcc2, 32'hc248cca7, 32'h4270fced, 32'h4294743f, 32'hc2bf1883};
test_output[4741] = '{32'h42a10c82};
test_index[4741] = '{0};
test_input[37936:37943] = '{32'hc22f6928, 32'h42c32c7f, 32'h41c9bbcb, 32'h4197621c, 32'h42522ddb, 32'hc2c49933, 32'hc2337d73, 32'hc109e261};
test_output[4742] = '{32'h42c32c7f};
test_index[4742] = '{1};
test_input[37944:37951] = '{32'h3fcec598, 32'hc2c150ff, 32'h409d7b4c, 32'hc1dbd4e0, 32'h41aa67b7, 32'h4289a511, 32'hc289732b, 32'hc102ff5f};
test_output[4743] = '{32'h4289a511};
test_index[4743] = '{5};
test_input[37952:37959] = '{32'hc2997262, 32'hc0c114a7, 32'hc2ad3ded, 32'h42bfb933, 32'hc1ca5e0a, 32'h4260178b, 32'h424c2726, 32'hc1a52ddc};
test_output[4744] = '{32'h42bfb933};
test_index[4744] = '{3};
test_input[37960:37967] = '{32'h423170ff, 32'hc1920c57, 32'h42b37803, 32'hc268c87e, 32'hc2922aca, 32'hc1c53f5d, 32'h423e9437, 32'h42ab8351};
test_output[4745] = '{32'h42b37803};
test_index[4745] = '{2};
test_input[37968:37975] = '{32'hc26804ff, 32'h4199eb05, 32'h42a87802, 32'hc2892a81, 32'hc1aabd70, 32'hc2845e4e, 32'hc1cf2106, 32'hc2658047};
test_output[4746] = '{32'h42a87802};
test_index[4746] = '{2};
test_input[37976:37983] = '{32'h42c75ab9, 32'hc10891b0, 32'h42074609, 32'hc01b19f3, 32'h414d6f71, 32'h40a69634, 32'h426accdf, 32'h40aa8abf};
test_output[4747] = '{32'h42c75ab9};
test_index[4747] = '{0};
test_input[37984:37991] = '{32'hc2bb099a, 32'h429b3f16, 32'hc2c5f3a6, 32'h422be4cb, 32'hc1a220d6, 32'hc24e5b76, 32'hc29a8771, 32'hc26a2ca8};
test_output[4748] = '{32'h429b3f16};
test_index[4748] = '{1};
test_input[37992:37999] = '{32'hc2834944, 32'h42292214, 32'hc257ae1c, 32'hc2b4cca4, 32'h42aca22e, 32'h42abf6ac, 32'hc2afa2d6, 32'hc1f5cfe1};
test_output[4749] = '{32'h42aca22e};
test_index[4749] = '{4};
test_input[38000:38007] = '{32'hc2892029, 32'hc28be2f6, 32'hc2610a56, 32'h422d9faa, 32'hc1d47df7, 32'h4267de95, 32'hc21ba865, 32'hc1105523};
test_output[4750] = '{32'h4267de95};
test_index[4750] = '{5};
test_input[38008:38015] = '{32'h42a38e36, 32'h428ab8b4, 32'h42a1de46, 32'hc1d30e08, 32'hc29e8812, 32'hc2aefa57, 32'h413a97f4, 32'h426e84e7};
test_output[4751] = '{32'h42a38e36};
test_index[4751] = '{0};
test_input[38016:38023] = '{32'hbfd81f70, 32'hc18db34a, 32'h40f9621a, 32'h429fa8fb, 32'h4294adb1, 32'hc276041b, 32'hc0ebb790, 32'h4240c794};
test_output[4752] = '{32'h429fa8fb};
test_index[4752] = '{3};
test_input[38024:38031] = '{32'h429a7b91, 32'hc200e962, 32'h4246dffc, 32'h41b0a5e1, 32'h42b247fe, 32'hc29d8886, 32'hc2363a0c, 32'h421067db};
test_output[4753] = '{32'h42b247fe};
test_index[4753] = '{4};
test_input[38032:38039] = '{32'h415253f5, 32'hc1596a00, 32'h4127c4ec, 32'hc27303b1, 32'h41b26e21, 32'hc2230dec, 32'h42832832, 32'h4271cea9};
test_output[4754] = '{32'h42832832};
test_index[4754] = '{6};
test_input[38040:38047] = '{32'hc28914a0, 32'h4253d3c9, 32'h421f171b, 32'hc29a8be4, 32'hc185030c, 32'h42aa0409, 32'hc1806617, 32'hc13be0d9};
test_output[4755] = '{32'h42aa0409};
test_index[4755] = '{5};
test_input[38048:38055] = '{32'h425e8af7, 32'hc2c43a1c, 32'hc22b9789, 32'hc2839287, 32'hc1c31e8f, 32'hc285065f, 32'hc2a5fb8f, 32'h4285129e};
test_output[4756] = '{32'h4285129e};
test_index[4756] = '{7};
test_input[38056:38063] = '{32'h400a1ace, 32'h42680fc4, 32'h42762649, 32'hc1f78a9c, 32'h411cd966, 32'h41d838e1, 32'h428b4a48, 32'hc27cb162};
test_output[4757] = '{32'h428b4a48};
test_index[4757] = '{6};
test_input[38064:38071] = '{32'hc2c0ff68, 32'h41eeef13, 32'h42afa1ef, 32'h42bdb2cc, 32'hc2b25763, 32'hc2a03970, 32'h42c3ffb1, 32'h4284babf};
test_output[4758] = '{32'h42c3ffb1};
test_index[4758] = '{6};
test_input[38072:38079] = '{32'h40ab999a, 32'hc281d0f8, 32'h412c0933, 32'hc2bebe20, 32'hc2bcb9df, 32'hc281d908, 32'hc284b953, 32'hc2aa2b03};
test_output[4759] = '{32'h412c0933};
test_index[4759] = '{2};
test_input[38080:38087] = '{32'hc2a5c933, 32'h42b37ccb, 32'h41801da7, 32'h424b9292, 32'hc2b549dc, 32'hc2a138fe, 32'h41ce99de, 32'h42703fe0};
test_output[4760] = '{32'h42b37ccb};
test_index[4760] = '{1};
test_input[38088:38095] = '{32'hc2b06973, 32'h424892d1, 32'h42acaa5c, 32'h429fb8e4, 32'h415b473d, 32'h40b5e007, 32'hc28be99a, 32'h41ecc5f1};
test_output[4761] = '{32'h42acaa5c};
test_index[4761] = '{2};
test_input[38096:38103] = '{32'h41c70cc6, 32'h4158447f, 32'hc2809df9, 32'hc2c25062, 32'hc2b47edf, 32'h42b31ebd, 32'hc1ef8d80, 32'hc2c6b42c};
test_output[4762] = '{32'h42b31ebd};
test_index[4762] = '{5};
test_input[38104:38111] = '{32'h40c9c122, 32'h41fa4b19, 32'hc29cb728, 32'h4298e3db, 32'hc2b8019c, 32'h424eac61, 32'hc294ff04, 32'hc2084e04};
test_output[4763] = '{32'h4298e3db};
test_index[4763] = '{3};
test_input[38112:38119] = '{32'h421c90fb, 32'h42480bff, 32'h42773d28, 32'hc28e44c0, 32'hc2c3970d, 32'hc1cf3763, 32'hc24f37e2, 32'hc2bd5f0a};
test_output[4764] = '{32'h42773d28};
test_index[4764] = '{2};
test_input[38120:38127] = '{32'h42689cc3, 32'hc2018dfc, 32'h4292642a, 32'h4282648a, 32'h423e866f, 32'hc2335662, 32'hc2bb3fec, 32'hc217b062};
test_output[4765] = '{32'h4292642a};
test_index[4765] = '{2};
test_input[38128:38135] = '{32'h40bcde7f, 32'h42476787, 32'h416b4e2d, 32'hc23c6a3c, 32'hc23501ff, 32'h4271707a, 32'hc1e0042a, 32'h40adc4a5};
test_output[4766] = '{32'h4271707a};
test_index[4766] = '{5};
test_input[38136:38143] = '{32'h412e8da5, 32'h428e30d4, 32'h4283a7c4, 32'h4202dd01, 32'h4290a4f0, 32'h42ad3967, 32'h42a85a45, 32'h411e7b30};
test_output[4767] = '{32'h42ad3967};
test_index[4767] = '{5};
test_input[38144:38151] = '{32'h423cb41c, 32'hc1c2c58e, 32'h42c1fff6, 32'h4195afe6, 32'h42427b65, 32'hc15577e7, 32'h41a3100d, 32'h42c41716};
test_output[4768] = '{32'h42c41716};
test_index[4768] = '{7};
test_input[38152:38159] = '{32'h4184f119, 32'hc25f1d3f, 32'hc2261238, 32'h424cce97, 32'h420c8d30, 32'h424e65e8, 32'hc2c3ece5, 32'h4191e002};
test_output[4769] = '{32'h424e65e8};
test_index[4769] = '{5};
test_input[38160:38167] = '{32'h4180b465, 32'h42a8d9e3, 32'h4288fe8c, 32'hc1b04f8d, 32'h411fe4e0, 32'hc146b8f5, 32'hc2924fdc, 32'h40e422af};
test_output[4770] = '{32'h42a8d9e3};
test_index[4770] = '{1};
test_input[38168:38175] = '{32'hc2723658, 32'h42b16533, 32'hc29be719, 32'hc2abbc29, 32'hc176d1cd, 32'h40547fcb, 32'h41a4fd6c, 32'hc1be2141};
test_output[4771] = '{32'h42b16533};
test_index[4771] = '{1};
test_input[38176:38183] = '{32'hc14c674b, 32'hc2c6ac52, 32'hc06c2384, 32'h42a91009, 32'h42be6251, 32'h41773a04, 32'hc2b86f33, 32'h42860019};
test_output[4772] = '{32'h42be6251};
test_index[4772] = '{4};
test_input[38184:38191] = '{32'hc2111b1d, 32'h429ee581, 32'hc2902b16, 32'h40b956e3, 32'h42a3e7f4, 32'h4293338b, 32'h4290a24f, 32'hc29c83b3};
test_output[4773] = '{32'h42a3e7f4};
test_index[4773] = '{4};
test_input[38192:38199] = '{32'hc2863939, 32'h42272d8c, 32'h4222989d, 32'hc28bd577, 32'hc22bde77, 32'h429a92a9, 32'h4209b49b, 32'hc265d598};
test_output[4774] = '{32'h429a92a9};
test_index[4774] = '{5};
test_input[38200:38207] = '{32'hc1c4908b, 32'hc225fa7b, 32'hc1a5a952, 32'hc299961f, 32'hc285e1fa, 32'hc299d700, 32'h429ecda4, 32'hc1be247d};
test_output[4775] = '{32'h429ecda4};
test_index[4775] = '{6};
test_input[38208:38215] = '{32'h42c00bf6, 32'h422fb8a1, 32'hc22a2343, 32'hc0a9954e, 32'hc0946259, 32'h4215b22d, 32'hc2a53d9b, 32'hc254f1fb};
test_output[4776] = '{32'h42c00bf6};
test_index[4776] = '{0};
test_input[38216:38223] = '{32'h4260df16, 32'hc1859000, 32'hc1820c89, 32'hc0751726, 32'hc1d80301, 32'h41ded2f1, 32'hc29b75df, 32'hc2993c63};
test_output[4777] = '{32'h4260df16};
test_index[4777] = '{0};
test_input[38224:38231] = '{32'h4285dc91, 32'h427c6d01, 32'h415ba4fb, 32'h4225e694, 32'h42c02b23, 32'hc2bf90b2, 32'h423db3ae, 32'hc000e40d};
test_output[4778] = '{32'h42c02b23};
test_index[4778] = '{4};
test_input[38232:38239] = '{32'hc20208fe, 32'hc2a04868, 32'h42aa50ed, 32'h402b7637, 32'hc264dfc8, 32'hc1442cdf, 32'hc1f324aa, 32'hc19b9782};
test_output[4779] = '{32'h42aa50ed};
test_index[4779] = '{2};
test_input[38240:38247] = '{32'hc0e15c7e, 32'hc23578da, 32'h42af7385, 32'hc2096147, 32'hc02faa88, 32'h423218de, 32'h419a2e56, 32'hc2b62c13};
test_output[4780] = '{32'h42af7385};
test_index[4780] = '{2};
test_input[38248:38255] = '{32'hc29bd65b, 32'hc29835a1, 32'hc228ae4b, 32'h423bcd02, 32'hc2983c4e, 32'hc18c6d41, 32'h42053592, 32'hc1e463aa};
test_output[4781] = '{32'h423bcd02};
test_index[4781] = '{3};
test_input[38256:38263] = '{32'h41cf5738, 32'h423c97dd, 32'hc2630321, 32'h42a10900, 32'h41cd9f21, 32'h42c44dc5, 32'h42c57203, 32'hc29b4a38};
test_output[4782] = '{32'h42c57203};
test_index[4782] = '{6};
test_input[38264:38271] = '{32'h42a6aad4, 32'h4156f300, 32'hc292055f, 32'h4278ecfa, 32'hc29ff685, 32'hc27c960c, 32'h410f6216, 32'hc2b557a2};
test_output[4783] = '{32'h42a6aad4};
test_index[4783] = '{0};
test_input[38272:38279] = '{32'h41796a3d, 32'h42810b35, 32'hc2528347, 32'h42a307c8, 32'h421dafa0, 32'hc25b2043, 32'h4176256d, 32'hc159412c};
test_output[4784] = '{32'h42a307c8};
test_index[4784] = '{3};
test_input[38280:38287] = '{32'h429b8def, 32'h42388b71, 32'h42c22da6, 32'h4120a561, 32'h42ba84a8, 32'hc21e0a22, 32'h42b85f75, 32'h41bb8d6e};
test_output[4785] = '{32'h42c22da6};
test_index[4785] = '{2};
test_input[38288:38295] = '{32'hc2c7dd89, 32'hc2c33b37, 32'h42a3c738, 32'hc212d271, 32'hc21a8d56, 32'h41b40d63, 32'hc29ed705, 32'hc1d06694};
test_output[4786] = '{32'h42a3c738};
test_index[4786] = '{2};
test_input[38296:38303] = '{32'hc136ba66, 32'h41b30e2b, 32'h4240d1c7, 32'hc0b3d46a, 32'hc22af68b, 32'hc2794240, 32'hc28dc1d6, 32'hc23c84bf};
test_output[4787] = '{32'h4240d1c7};
test_index[4787] = '{2};
test_input[38304:38311] = '{32'h42585af1, 32'h42a9419f, 32'hc19b31db, 32'hc1a35084, 32'h4204055a, 32'hc2175595, 32'h418cef75, 32'hc259df84};
test_output[4788] = '{32'h42a9419f};
test_index[4788] = '{1};
test_input[38312:38319] = '{32'hc28aa663, 32'hc29f9bbb, 32'h41ccc52a, 32'h4232409c, 32'h42be33f4, 32'h3ff7a73c, 32'hc1d5acde, 32'h42030400};
test_output[4789] = '{32'h42be33f4};
test_index[4789] = '{4};
test_input[38320:38327] = '{32'h404dc621, 32'h4134e997, 32'hc28a60e7, 32'hc2bdc822, 32'h41c7b188, 32'hc1b4f98b, 32'hc244d287, 32'h42c4b2cd};
test_output[4790] = '{32'h42c4b2cd};
test_index[4790] = '{7};
test_input[38328:38335] = '{32'h42b8182d, 32'h42875bb2, 32'hc284f41f, 32'hc2a7713b, 32'hc2b76212, 32'hc1fac9e1, 32'h41f19c81, 32'h40cef65a};
test_output[4791] = '{32'h42b8182d};
test_index[4791] = '{0};
test_input[38336:38343] = '{32'h41376247, 32'h4263d307, 32'hc24da7ad, 32'h41b1a95d, 32'h4214b37a, 32'h425abe94, 32'h400c894f, 32'hc1cd4284};
test_output[4792] = '{32'h4263d307};
test_index[4792] = '{1};
test_input[38344:38351] = '{32'hc1d85d8e, 32'hc2389a06, 32'h41819122, 32'h4222d855, 32'h41655286, 32'h4206678f, 32'hc2b02791, 32'hc27ec90b};
test_output[4793] = '{32'h4222d855};
test_index[4793] = '{3};
test_input[38352:38359] = '{32'h42678d60, 32'h428a1e85, 32'h401dcc0b, 32'h4244acba, 32'hc2a39e97, 32'hc2202a77, 32'hc23ac548, 32'hc2b1675e};
test_output[4794] = '{32'h428a1e85};
test_index[4794] = '{1};
test_input[38360:38367] = '{32'h42476e43, 32'hc1f18b0c, 32'hc22e1cb2, 32'h42b9b0fe, 32'h410d4fca, 32'hc2051224, 32'h41d9c6d7, 32'h4291b900};
test_output[4795] = '{32'h42b9b0fe};
test_index[4795] = '{3};
test_input[38368:38375] = '{32'hc2b10e59, 32'h41537c8d, 32'hc2b3ea82, 32'hc26ba9c9, 32'h42bb8982, 32'h42aad34f, 32'h42757d78, 32'h419267c7};
test_output[4796] = '{32'h42bb8982};
test_index[4796] = '{4};
test_input[38376:38383] = '{32'h4268331d, 32'hc20f2255, 32'hc27ec617, 32'h4230b174, 32'hc1f0f8b2, 32'h4215a2a6, 32'h42c25a24, 32'h41024494};
test_output[4797] = '{32'h42c25a24};
test_index[4797] = '{6};
test_input[38384:38391] = '{32'h425140eb, 32'hc20d0f2a, 32'h418edebc, 32'hc27a7da0, 32'h42017276, 32'h40be20b7, 32'hc294b6e7, 32'h4110a0e2};
test_output[4798] = '{32'h425140eb};
test_index[4798] = '{0};
test_input[38392:38399] = '{32'hc2baa74a, 32'h421954ec, 32'hc2433bd3, 32'hc19ec835, 32'hc1c989a4, 32'h4209f73f, 32'h429634b9, 32'h42220393};
test_output[4799] = '{32'h429634b9};
test_index[4799] = '{6};
test_input[38400:38407] = '{32'h4267692e, 32'hc2145eb6, 32'hc1ed4b69, 32'h40117627, 32'h41cd666a, 32'hc193f79d, 32'h41dd5529, 32'h42231b1b};
test_output[4800] = '{32'h4267692e};
test_index[4800] = '{0};
test_input[38408:38415] = '{32'h4202ad31, 32'h420cd56e, 32'hc0bd44e4, 32'h42b72984, 32'h42bbd4e3, 32'hc1c45882, 32'h42ad5c94, 32'hc23ca369};
test_output[4801] = '{32'h42bbd4e3};
test_index[4801] = '{4};
test_input[38416:38423] = '{32'hc23abd1c, 32'h42bd5484, 32'hc20e5070, 32'h4281a3fd, 32'hc284eba2, 32'hc2adf4a5, 32'h425ee58d, 32'hc1ca61ea};
test_output[4802] = '{32'h42bd5484};
test_index[4802] = '{1};
test_input[38424:38431] = '{32'hc29932c4, 32'hc268a649, 32'hc263573d, 32'h42355130, 32'h41e6fd3e, 32'h423936f7, 32'hc0ca35d4, 32'hc28fecf8};
test_output[4803] = '{32'h423936f7};
test_index[4803] = '{5};
test_input[38432:38439] = '{32'hc030a5da, 32'h4200b8b5, 32'hc2279265, 32'h4140165c, 32'h429a157e, 32'hc2aa44a3, 32'hc2696925, 32'h3fac3fad};
test_output[4804] = '{32'h429a157e};
test_index[4804] = '{4};
test_input[38440:38447] = '{32'hc2c2ccc5, 32'hc22d3b2c, 32'hc28479f9, 32'h40b338d1, 32'hc2b33e18, 32'hc1fc86f3, 32'hc0a5ae8a, 32'hc26746ac};
test_output[4805] = '{32'h40b338d1};
test_index[4805] = '{3};
test_input[38448:38455] = '{32'hc081d88c, 32'hc2912a17, 32'h41a8ba1a, 32'h428ba753, 32'hc2942cf3, 32'h429b9651, 32'h42633013, 32'h424f1313};
test_output[4806] = '{32'h429b9651};
test_index[4806] = '{5};
test_input[38456:38463] = '{32'h42979277, 32'hc28b195b, 32'hc2491c54, 32'h41efc6b8, 32'h4209b3ab, 32'h42b24a1f, 32'hc23e51b0, 32'h400e37fd};
test_output[4807] = '{32'h42b24a1f};
test_index[4807] = '{5};
test_input[38464:38471] = '{32'h41e7f35c, 32'h42417f30, 32'h429c1ade, 32'h40cdfdca, 32'hc21f1d0c, 32'hc29e8b9f, 32'hc24596e2, 32'hc15d9e1a};
test_output[4808] = '{32'h429c1ade};
test_index[4808] = '{2};
test_input[38472:38479] = '{32'h41211ff3, 32'hc1f962d2, 32'hc153636c, 32'h41779aa3, 32'h423b2128, 32'hc190cbbb, 32'hc2bd943d, 32'hc2c60507};
test_output[4809] = '{32'h423b2128};
test_index[4809] = '{4};
test_input[38480:38487] = '{32'h42ac9552, 32'h423cc532, 32'hc0ac67b1, 32'h41b18de8, 32'hc16b2348, 32'hc209bbad, 32'h423c4efc, 32'h42bdade8};
test_output[4810] = '{32'h42bdade8};
test_index[4810] = '{7};
test_input[38488:38495] = '{32'hc2a48a5c, 32'hc2a2fe47, 32'h42c09dc7, 32'h429d2329, 32'h4231dce7, 32'hc26eb93c, 32'h419290e8, 32'h41901957};
test_output[4811] = '{32'h42c09dc7};
test_index[4811] = '{2};
test_input[38496:38503] = '{32'h42a4989e, 32'h42221583, 32'hc2a55264, 32'h425078ab, 32'hbff623f8, 32'hc01dc826, 32'h427b5e20, 32'hc299c547};
test_output[4812] = '{32'h42a4989e};
test_index[4812] = '{0};
test_input[38504:38511] = '{32'hc2427915, 32'hc2913021, 32'hc2357683, 32'hc26230f6, 32'h41c8fdd3, 32'h42086847, 32'h42370e32, 32'h426382e6};
test_output[4813] = '{32'h426382e6};
test_index[4813] = '{7};
test_input[38512:38519] = '{32'h42c33fc7, 32'h4184d508, 32'h42bef0f0, 32'h41a9acd9, 32'h4209363b, 32'h410bfdcc, 32'h42c36aa0, 32'hc29b30cc};
test_output[4814] = '{32'h42c36aa0};
test_index[4814] = '{6};
test_input[38520:38527] = '{32'hc1bf9cc0, 32'hc2850f14, 32'hc2324735, 32'h41daf3c1, 32'h42b10850, 32'h42769dc7, 32'hc2786d87, 32'hc2633596};
test_output[4815] = '{32'h42b10850};
test_index[4815] = '{4};
test_input[38528:38535] = '{32'hc1a389ad, 32'hc2196229, 32'hc157342e, 32'hc298e4e8, 32'hc2814b59, 32'hc1d4ba62, 32'h42703dfc, 32'hc23147b5};
test_output[4816] = '{32'h42703dfc};
test_index[4816] = '{6};
test_input[38536:38543] = '{32'h424805dd, 32'h40cf59ca, 32'hc1e76adf, 32'h42b768a5, 32'h42b0bd56, 32'hc2ae1767, 32'hc1ada16f, 32'h4291a5ab};
test_output[4817] = '{32'h42b768a5};
test_index[4817] = '{3};
test_input[38544:38551] = '{32'h42a48e29, 32'h426279ab, 32'hc0df16e6, 32'h4126de14, 32'h42be9cf3, 32'hc2943a56, 32'h4267def3, 32'h419e3223};
test_output[4818] = '{32'h42be9cf3};
test_index[4818] = '{4};
test_input[38552:38559] = '{32'hbfbe8736, 32'hc2bc1643, 32'hc28592a3, 32'h420bb615, 32'h41a16ada, 32'hbfa184f3, 32'hc272c335, 32'h408c2805};
test_output[4819] = '{32'h420bb615};
test_index[4819] = '{3};
test_input[38560:38567] = '{32'h42a846fd, 32'h42c19ba2, 32'h419f9199, 32'h42015352, 32'hc1d4338c, 32'hc27bac34, 32'hc28f4e03, 32'h428f8917};
test_output[4820] = '{32'h42c19ba2};
test_index[4820] = '{1};
test_input[38568:38575] = '{32'hc2ae7ee0, 32'hc2aef0ab, 32'hc1dce977, 32'h4245b839, 32'hc2812980, 32'h42465655, 32'hc2678a67, 32'h410e9aa1};
test_output[4821] = '{32'h42465655};
test_index[4821] = '{5};
test_input[38576:38583] = '{32'h41cd005d, 32'h421b4776, 32'h423c0227, 32'hc2972ffe, 32'h424fa0b3, 32'hc2814e96, 32'hc10a7807, 32'h41652742};
test_output[4822] = '{32'h424fa0b3};
test_index[4822] = '{4};
test_input[38584:38591] = '{32'h42ada2b8, 32'h42487a0d, 32'h42732403, 32'h42c32484, 32'hc29aa365, 32'h42c669ea, 32'h42c2d446, 32'hc29e3a23};
test_output[4823] = '{32'h42c669ea};
test_index[4823] = '{5};
test_input[38592:38599] = '{32'h424a7889, 32'hc202d458, 32'h40a0b457, 32'hc1318472, 32'h42a3b0bc, 32'h41ef3d87, 32'h41cf089f, 32'hc2c3ab2e};
test_output[4824] = '{32'h42a3b0bc};
test_index[4824] = '{4};
test_input[38600:38607] = '{32'hc27e8387, 32'h42bda142, 32'h4261efac, 32'hc2ac440e, 32'h41c46911, 32'hc2abd1d0, 32'hc25405c3, 32'hc2bbccb5};
test_output[4825] = '{32'h42bda142};
test_index[4825] = '{1};
test_input[38608:38615] = '{32'hc274e46b, 32'h41f9ddb2, 32'hc289def7, 32'hc1cea111, 32'h41a48bba, 32'h4290609f, 32'hc26d4549, 32'h421932f1};
test_output[4826] = '{32'h4290609f};
test_index[4826] = '{5};
test_input[38616:38623] = '{32'hc1dc9c0a, 32'h419e915a, 32'h41915546, 32'hc1a658a1, 32'h4267a351, 32'hc2827ab5, 32'hc14fb54f, 32'h42a2af2c};
test_output[4827] = '{32'h42a2af2c};
test_index[4827] = '{7};
test_input[38624:38631] = '{32'h4252b037, 32'hc2b81e11, 32'hc1bceed6, 32'h414f167f, 32'h42853a4d, 32'h41a74118, 32'h41d5130b, 32'h421a0697};
test_output[4828] = '{32'h42853a4d};
test_index[4828] = '{4};
test_input[38632:38639] = '{32'h41bc0964, 32'hc2a0e20e, 32'h41bc63ba, 32'h42889ad9, 32'h426ddefa, 32'h42311838, 32'h426f2c68, 32'hc2c64e62};
test_output[4829] = '{32'h42889ad9};
test_index[4829] = '{3};
test_input[38640:38647] = '{32'h4237cb56, 32'hc2879356, 32'hc1e6efb5, 32'h42bade7e, 32'hc28f7b0c, 32'h4289e002, 32'hbf98e9f9, 32'h417bb494};
test_output[4830] = '{32'h42bade7e};
test_index[4830] = '{3};
test_input[38648:38655] = '{32'hc26f423d, 32'h42b93181, 32'hc21072e3, 32'hc28ca93d, 32'hc2406ae1, 32'hc2b3ec81, 32'hc20ce703, 32'h421af241};
test_output[4831] = '{32'h42b93181};
test_index[4831] = '{1};
test_input[38656:38663] = '{32'hc21806cc, 32'h41ecc7a1, 32'h424c3002, 32'hc2ac0cf9, 32'hc083c042, 32'hc1b1b993, 32'hc18cdd78, 32'h426bdac9};
test_output[4832] = '{32'h426bdac9};
test_index[4832] = '{7};
test_input[38664:38671] = '{32'hc2c1e65a, 32'h41589613, 32'hc21c341e, 32'h4290826f, 32'h3ff4f5d5, 32'h42b91a15, 32'h428775ad, 32'h42855a85};
test_output[4833] = '{32'h42b91a15};
test_index[4833] = '{5};
test_input[38672:38679] = '{32'hc2843768, 32'h4287632d, 32'hc29da793, 32'hbf635492, 32'hc0b55de8, 32'h3ed295f5, 32'h42a908e9, 32'h429081eb};
test_output[4834] = '{32'h42a908e9};
test_index[4834] = '{6};
test_input[38680:38687] = '{32'hc21b13cd, 32'hc17a0058, 32'hc142cc06, 32'hc29cdcc0, 32'h41fe5e87, 32'h42967d41, 32'hc209b74a, 32'h4262de68};
test_output[4835] = '{32'h42967d41};
test_index[4835] = '{5};
test_input[38688:38695] = '{32'hc28eb217, 32'h42a55bc9, 32'hc005de66, 32'h42b379c1, 32'h426a21f2, 32'h4088c17a, 32'h42857495, 32'h41bd77c6};
test_output[4836] = '{32'h42b379c1};
test_index[4836] = '{3};
test_input[38696:38703] = '{32'hc1fa9d76, 32'hc189ca08, 32'hc2a2f359, 32'hc1f29935, 32'hc20d0ae8, 32'h422c4392, 32'h42a5985c, 32'h40ba0b93};
test_output[4837] = '{32'h42a5985c};
test_index[4837] = '{6};
test_input[38704:38711] = '{32'hc1dc06f2, 32'h42aca550, 32'h41b739d5, 32'hc1d4a4c6, 32'h42aabf73, 32'hc09b1a18, 32'h42880def, 32'hbfc0ed87};
test_output[4838] = '{32'h42aca550};
test_index[4838] = '{1};
test_input[38712:38719] = '{32'h42413d76, 32'hc2b38d50, 32'hc2666e67, 32'hc217224f, 32'hc13e0a9c, 32'hc26d5e5b, 32'hc26fb0de, 32'hc22aebaf};
test_output[4839] = '{32'h42413d76};
test_index[4839] = '{0};
test_input[38720:38727] = '{32'hc22afec5, 32'hc21008ed, 32'hc2beb95d, 32'hc28f51e1, 32'h426ee282, 32'h41833307, 32'h42bde0cd, 32'hc1f1425b};
test_output[4840] = '{32'h42bde0cd};
test_index[4840] = '{6};
test_input[38728:38735] = '{32'hc2117bc5, 32'hc2b882b6, 32'h42ba7cf3, 32'hc28d5345, 32'h42a07b10, 32'h41d91652, 32'h4130c39a, 32'h4186c6b7};
test_output[4841] = '{32'h42ba7cf3};
test_index[4841] = '{2};
test_input[38736:38743] = '{32'hc2c1fd0b, 32'h420c2fbb, 32'hc25810c9, 32'hc268449c, 32'hc21d942b, 32'hc287e761, 32'hc1f08d3e, 32'h42a98da4};
test_output[4842] = '{32'h42a98da4};
test_index[4842] = '{7};
test_input[38744:38751] = '{32'h42158e71, 32'h4217bbaf, 32'h4291606b, 32'hc21d3290, 32'h41d552cc, 32'hc23a07ae, 32'hc292d29a, 32'hc0e0d082};
test_output[4843] = '{32'h4291606b};
test_index[4843] = '{2};
test_input[38752:38759] = '{32'hc278a6d5, 32'hc1bcb4bc, 32'h4296dcf9, 32'hc27447a5, 32'h425c958b, 32'hc2c4b31b, 32'hc2142c9c, 32'hc2b919e6};
test_output[4844] = '{32'h4296dcf9};
test_index[4844] = '{2};
test_input[38760:38767] = '{32'hc283a781, 32'h421cf104, 32'hc285c9c5, 32'h4281f07d, 32'hc19e7e18, 32'hc2af85d1, 32'hc24bf020, 32'hc2aa774f};
test_output[4845] = '{32'h4281f07d};
test_index[4845] = '{3};
test_input[38768:38775] = '{32'h40813640, 32'hc26d777f, 32'h426d0ee8, 32'hc19641ab, 32'h41bf93ca, 32'h428e12a1, 32'h41624dd4, 32'h42c277af};
test_output[4846] = '{32'h42c277af};
test_index[4846] = '{7};
test_input[38776:38783] = '{32'h418f704e, 32'hc1a860d7, 32'hc0f2204f, 32'hc253274d, 32'h42ad1de2, 32'hc2aa1e46, 32'hc0ea1ed7, 32'h42071544};
test_output[4847] = '{32'h42ad1de2};
test_index[4847] = '{4};
test_input[38784:38791] = '{32'h41a93885, 32'h425006c8, 32'h417f266a, 32'h4297cb4f, 32'h41f8c8db, 32'hc1909bc3, 32'hc1a9169e, 32'hc1c226e8};
test_output[4848] = '{32'h4297cb4f};
test_index[4848] = '{3};
test_input[38792:38799] = '{32'hc2245d9a, 32'h42a13960, 32'h41b1112f, 32'h42c78373, 32'h424950c4, 32'hc006e450, 32'h411ee567, 32'h41e574d9};
test_output[4849] = '{32'h42c78373};
test_index[4849] = '{3};
test_input[38800:38807] = '{32'h42b6b532, 32'h41d38860, 32'h4204b348, 32'hc1910983, 32'h4223eee7, 32'h428ecff8, 32'hc2ac618d, 32'h42afe595};
test_output[4850] = '{32'h42b6b532};
test_index[4850] = '{0};
test_input[38808:38815] = '{32'hc2a20517, 32'hc2a8a0ee, 32'hc2649e4f, 32'hbefb631e, 32'hc21a170a, 32'h40d1b4cf, 32'hc240b1c2, 32'h4283eccb};
test_output[4851] = '{32'h4283eccb};
test_index[4851] = '{7};
test_input[38816:38823] = '{32'hc2c0cbe6, 32'hc223f62d, 32'h4255319d, 32'hc2b1926f, 32'hc21d5998, 32'hc1cefc7d, 32'hc249daf1, 32'h42a196c0};
test_output[4852] = '{32'h42a196c0};
test_index[4852] = '{7};
test_input[38824:38831] = '{32'h423fbc9a, 32'h42b34549, 32'h42872f8b, 32'h4284480a, 32'h404a69f9, 32'h4203885c, 32'hc2931200, 32'hc2a6efa6};
test_output[4853] = '{32'h42b34549};
test_index[4853] = '{1};
test_input[38832:38839] = '{32'hc1fba0fe, 32'h422bbf14, 32'hc22f9593, 32'h42649d91, 32'h429eda6f, 32'h3ecca2af, 32'h42c58846, 32'h42146ec7};
test_output[4854] = '{32'h42c58846};
test_index[4854] = '{6};
test_input[38840:38847] = '{32'h424eb08d, 32'h41edd0e3, 32'h427f5e3c, 32'hc2340a66, 32'hc212863e, 32'h42a21c90, 32'hc2ab379b, 32'hc173c85a};
test_output[4855] = '{32'h42a21c90};
test_index[4855] = '{5};
test_input[38848:38855] = '{32'h403ca4de, 32'h41c78b5d, 32'hc1ca3f7e, 32'h421031fd, 32'h419a1088, 32'hc1a6993a, 32'hc2a39f62, 32'hc29055f4};
test_output[4856] = '{32'h421031fd};
test_index[4856] = '{3};
test_input[38856:38863] = '{32'h42277e17, 32'h42c53f3f, 32'h42392572, 32'hc1748b56, 32'hc23707a9, 32'h42813d3f, 32'hc2109a90, 32'h424a4b76};
test_output[4857] = '{32'h42c53f3f};
test_index[4857] = '{1};
test_input[38864:38871] = '{32'hc09f4617, 32'hc25641e4, 32'hc29c0205, 32'hc291c5b5, 32'hc2b6f7f4, 32'hc2497f6f, 32'h423090fe, 32'h4031c6b8};
test_output[4858] = '{32'h423090fe};
test_index[4858] = '{6};
test_input[38872:38879] = '{32'h428570a1, 32'hc18777fa, 32'h42922ed5, 32'hc126990e, 32'hc218336a, 32'h41cd5322, 32'h40c1556c, 32'hc221aaa0};
test_output[4859] = '{32'h42922ed5};
test_index[4859] = '{2};
test_input[38880:38887] = '{32'hc221faba, 32'h423ac532, 32'hc2aa3941, 32'h42a54f2a, 32'h42a20dbc, 32'h42c04965, 32'hbff16982, 32'h425e9eec};
test_output[4860] = '{32'h42c04965};
test_index[4860] = '{5};
test_input[38888:38895] = '{32'hc2b39ed8, 32'hc2ab60a3, 32'h425064a3, 32'hc2a5f8ec, 32'h4201a582, 32'h419af181, 32'h40435f74, 32'h423fdd3d};
test_output[4861] = '{32'h425064a3};
test_index[4861] = '{2};
test_input[38896:38903] = '{32'h420b21c0, 32'h421d6e75, 32'hc23c811f, 32'h4265231d, 32'hc29d2b3b, 32'h42632aa7, 32'hc28cd6d4, 32'hc2bf4279};
test_output[4862] = '{32'h4265231d};
test_index[4862] = '{3};
test_input[38904:38911] = '{32'hc2c55463, 32'h424e6aa2, 32'hc0f5ae8a, 32'hc1f97ac5, 32'hc23bdbca, 32'h41f5ceac, 32'hc2980ca5, 32'h41f990c8};
test_output[4863] = '{32'h424e6aa2};
test_index[4863] = '{1};
test_input[38912:38919] = '{32'hc24fafc7, 32'h429f824e, 32'h4211f2ba, 32'h425f25e1, 32'h42a1545d, 32'h4249a919, 32'hc28b5a25, 32'h42785bf7};
test_output[4864] = '{32'h42a1545d};
test_index[4864] = '{4};
test_input[38920:38927] = '{32'h421e2725, 32'h41c6c252, 32'h4197a8f6, 32'h4183a142, 32'h4282751a, 32'h429a9172, 32'hc1afe236, 32'h42475c4e};
test_output[4865] = '{32'h429a9172};
test_index[4865] = '{5};
test_input[38928:38935] = '{32'h40f9f808, 32'h41d5db2f, 32'h4150202b, 32'h42753af3, 32'hc16131e6, 32'hc21fd14d, 32'hc24bd7e0, 32'hc2bc9d8b};
test_output[4866] = '{32'h42753af3};
test_index[4866] = '{3};
test_input[38936:38943] = '{32'h42954375, 32'hc131de0a, 32'hc24bcf83, 32'hc2a085e0, 32'h407ae994, 32'h41ef1688, 32'h42c5d76d, 32'hc16f892b};
test_output[4867] = '{32'h42c5d76d};
test_index[4867] = '{6};
test_input[38944:38951] = '{32'hc28f4736, 32'hc2017a97, 32'h42b0e0ed, 32'hc2ac81fe, 32'hc2a1d823, 32'h421f2154, 32'h42736fe6, 32'h421e9227};
test_output[4868] = '{32'h42b0e0ed};
test_index[4868] = '{2};
test_input[38952:38959] = '{32'h42b087ca, 32'h42146489, 32'hc12c16c5, 32'hc1af282c, 32'h424e1f42, 32'h41e1fb8d, 32'hc295ff2a, 32'hc24be054};
test_output[4869] = '{32'h42b087ca};
test_index[4869] = '{0};
test_input[38960:38967] = '{32'h42887dae, 32'hc2759682, 32'h41ee3e18, 32'h41804e83, 32'h42a596d3, 32'hc2992f0f, 32'h41df8cc3, 32'hc1820a9a};
test_output[4870] = '{32'h42a596d3};
test_index[4870] = '{4};
test_input[38968:38975] = '{32'h419b93e2, 32'h402e3311, 32'hc12b7919, 32'h4084cb86, 32'h42a17316, 32'h428101ab, 32'hc29df874, 32'h42b744f9};
test_output[4871] = '{32'h42b744f9};
test_index[4871] = '{7};
test_input[38976:38983] = '{32'hc2c26483, 32'h41f3f858, 32'hc1816c3a, 32'h42480a0c, 32'h4279934d, 32'h4154ac90, 32'h42833b9f, 32'hc1a2fd26};
test_output[4872] = '{32'h42833b9f};
test_index[4872] = '{6};
test_input[38984:38991] = '{32'hc294b271, 32'hc0cf8d79, 32'hc2166b4f, 32'h428195a8, 32'h42b50a44, 32'h42864255, 32'hc21403bb, 32'hc29a5cdf};
test_output[4873] = '{32'h42b50a44};
test_index[4873] = '{4};
test_input[38992:38999] = '{32'hc220e50a, 32'h429abb97, 32'h425a4615, 32'hc1b1a289, 32'hc20dd570, 32'h418d7912, 32'h42c67d3f, 32'hc28efeed};
test_output[4874] = '{32'h42c67d3f};
test_index[4874] = '{6};
test_input[39000:39007] = '{32'h4292e4ed, 32'hc2c01e96, 32'h4236dad8, 32'hc17ad82d, 32'h41da9c88, 32'h41c926f5, 32'hc2bd50ec, 32'h4277551b};
test_output[4875] = '{32'h4292e4ed};
test_index[4875] = '{0};
test_input[39008:39015] = '{32'hbfb77559, 32'h421be04b, 32'h429f5fe2, 32'h42b13f1e, 32'h4225928e, 32'h42311a51, 32'hc211aea6, 32'hc23e9c33};
test_output[4876] = '{32'h42b13f1e};
test_index[4876] = '{3};
test_input[39016:39023] = '{32'h41855884, 32'hc229d591, 32'h41b7ea6c, 32'h421b630b, 32'h427fd670, 32'hc177ed8a, 32'hc2a5a462, 32'hc180f01a};
test_output[4877] = '{32'h427fd670};
test_index[4877] = '{4};
test_input[39024:39031] = '{32'hc2aa02c8, 32'hc11a1915, 32'h42ad804a, 32'hc293dfe2, 32'h42c5a014, 32'h4289ca36, 32'hc2bc1498, 32'hc205d67e};
test_output[4878] = '{32'h42c5a014};
test_index[4878] = '{4};
test_input[39032:39039] = '{32'hc1321307, 32'hc2887364, 32'h41bd9902, 32'hc28b08a9, 32'h4200d6b1, 32'h42bc955d, 32'hc28f851e, 32'h428ff1cd};
test_output[4879] = '{32'h42bc955d};
test_index[4879] = '{5};
test_input[39040:39047] = '{32'h41a6fe96, 32'hc2a8f70f, 32'hc1677c2b, 32'h4281c007, 32'h42a8748c, 32'h4117a545, 32'hc28514a0, 32'h418acfe7};
test_output[4880] = '{32'h42a8748c};
test_index[4880] = '{4};
test_input[39048:39055] = '{32'h42bd6cf5, 32'hc23255b8, 32'h42189e5d, 32'hc1f692a4, 32'hc16af090, 32'h4264e8fb, 32'hc18d62aa, 32'h42b7fb31};
test_output[4881] = '{32'h42bd6cf5};
test_index[4881] = '{0};
test_input[39056:39063] = '{32'hc2b0dddc, 32'hc28313f3, 32'h42a1f411, 32'h411d1711, 32'h42164de0, 32'hc289de5a, 32'h424f4d16, 32'h42bf64ba};
test_output[4882] = '{32'h42bf64ba};
test_index[4882] = '{7};
test_input[39064:39071] = '{32'h41773594, 32'hc21ea12a, 32'hc2747edc, 32'h41ea84dc, 32'hc15e8796, 32'hc207c93f, 32'h4297e7fc, 32'h42888b20};
test_output[4883] = '{32'h4297e7fc};
test_index[4883] = '{6};
test_input[39072:39079] = '{32'hc227e0d4, 32'hc01df08d, 32'h42199305, 32'h419ece51, 32'h4288572b, 32'hc2761a5e, 32'hc2934a6e, 32'h42216ac8};
test_output[4884] = '{32'h4288572b};
test_index[4884] = '{4};
test_input[39080:39087] = '{32'hc1a6180f, 32'h416ef29f, 32'hc19e17b6, 32'hc2be2630, 32'h4106900a, 32'hc2288382, 32'h422dceb2, 32'hc1b26632};
test_output[4885] = '{32'h422dceb2};
test_index[4885] = '{6};
test_input[39088:39095] = '{32'hc1b2da34, 32'hc2334808, 32'hc053cbea, 32'h4276365c, 32'hc287711c, 32'h427562da, 32'hc2076ccd, 32'h422d56bc};
test_output[4886] = '{32'h4276365c};
test_index[4886] = '{3};
test_input[39096:39103] = '{32'h4279b4f7, 32'hc2aa6cbd, 32'h428b0fa5, 32'hc244a16d, 32'hc28917dd, 32'h42869101, 32'h424cd92f, 32'h42478ae6};
test_output[4887] = '{32'h428b0fa5};
test_index[4887] = '{2};
test_input[39104:39111] = '{32'h4207d4cd, 32'hc0b6b7f9, 32'hc231e571, 32'hc2b3bb6a, 32'h42c5e377, 32'hc2443558, 32'h403d07a7, 32'h4109ea31};
test_output[4888] = '{32'h42c5e377};
test_index[4888] = '{4};
test_input[39112:39119] = '{32'h3f4a9eca, 32'h423c02d2, 32'hc1d01020, 32'h428d8e84, 32'hc163074d, 32'h42a66242, 32'hc291b0c0, 32'hc22903dd};
test_output[4889] = '{32'h42a66242};
test_index[4889] = '{5};
test_input[39120:39127] = '{32'h42222a65, 32'hc27f9419, 32'h420c46e8, 32'h41226815, 32'h41e0a56c, 32'h4299fe5e, 32'h42c6317d, 32'h3fded87e};
test_output[4890] = '{32'h42c6317d};
test_index[4890] = '{6};
test_input[39128:39135] = '{32'h41230e43, 32'hc2009454, 32'hc2960bf5, 32'hc2ac098a, 32'h41cf8001, 32'h41bb9b84, 32'hc2c21937, 32'hc29281cf};
test_output[4891] = '{32'h41cf8001};
test_index[4891] = '{4};
test_input[39136:39143] = '{32'h415a1f53, 32'h42716f7a, 32'h42b520c6, 32'hc102bfbe, 32'hc2a7fb00, 32'hc1808788, 32'h41410dd5, 32'hc17ce8e9};
test_output[4892] = '{32'h42b520c6};
test_index[4892] = '{2};
test_input[39144:39151] = '{32'hc289bfee, 32'h42a76c77, 32'hc2657b0f, 32'hc25b401e, 32'hc2a3c469, 32'hc19e48f8, 32'h42bbc993, 32'h41b2050b};
test_output[4893] = '{32'h42bbc993};
test_index[4893] = '{6};
test_input[39152:39159] = '{32'hc2c07f7d, 32'h417120a7, 32'hc18bb66f, 32'hc2abe0bf, 32'h428c0e28, 32'hc1660786, 32'h42bd2bcd, 32'hc2ba3735};
test_output[4894] = '{32'h42bd2bcd};
test_index[4894] = '{6};
test_input[39160:39167] = '{32'h41a655b1, 32'hc29bd5f0, 32'hc291f67d, 32'hc19d8748, 32'hc1a30bce, 32'hc29f0288, 32'hc15f0bdb, 32'h42bced5f};
test_output[4895] = '{32'h42bced5f};
test_index[4895] = '{7};
test_input[39168:39175] = '{32'hc185befb, 32'hc20100a3, 32'h42834507, 32'hc293ad75, 32'h41c649fc, 32'hc2aaf24f, 32'hc2811560, 32'h4289631a};
test_output[4896] = '{32'h4289631a};
test_index[4896] = '{7};
test_input[39176:39183] = '{32'h419daf88, 32'hc2812825, 32'h4110a6b4, 32'hc2898fa2, 32'h4291c3e6, 32'h423b5c12, 32'h42a82bc6, 32'h42a48eed};
test_output[4897] = '{32'h42a82bc6};
test_index[4897] = '{6};
test_input[39184:39191] = '{32'h4290f061, 32'hc28dbc0e, 32'h429dd6af, 32'hc2430a77, 32'hbd75c554, 32'h4298bc19, 32'h428ad52a, 32'h42b39137};
test_output[4898] = '{32'h42b39137};
test_index[4898] = '{7};
test_input[39192:39199] = '{32'hc27b4dcd, 32'hc208b530, 32'hc1b0d127, 32'h42b35944, 32'h42bf2535, 32'h42927c82, 32'h42b13d5c, 32'h429dda3c};
test_output[4899] = '{32'h42bf2535};
test_index[4899] = '{4};
test_input[39200:39207] = '{32'h41805df8, 32'hc2b830ce, 32'hc107b2e4, 32'h4183fb23, 32'h42a907fb, 32'h41ac4509, 32'hc298277e, 32'hc1528275};
test_output[4900] = '{32'h42a907fb};
test_index[4900] = '{4};
test_input[39208:39215] = '{32'hc296a4f1, 32'h414674d9, 32'hc0b47353, 32'hc13906d5, 32'hc23c4112, 32'h42265a5c, 32'h41300606, 32'h42b7f9b2};
test_output[4901] = '{32'h42b7f9b2};
test_index[4901] = '{7};
test_input[39216:39223] = '{32'hc21f8aff, 32'hc29f04d8, 32'h42bf0cc8, 32'h42c115a9, 32'hc287ea64, 32'h42c34d3f, 32'hc2663363, 32'hc1a47bf4};
test_output[4902] = '{32'h42c34d3f};
test_index[4902] = '{5};
test_input[39224:39231] = '{32'hc250f5fa, 32'h4226ca8c, 32'hc22b7a85, 32'h428ffc46, 32'hc2960a3e, 32'hc2926a4c, 32'hc18dd554, 32'hc27344aa};
test_output[4903] = '{32'h428ffc46};
test_index[4903] = '{3};
test_input[39232:39239] = '{32'h42bad1ed, 32'hc297934c, 32'hc1a46e92, 32'hc220dd9b, 32'h42765b2c, 32'h413498c9, 32'h429dae71, 32'hc24925e3};
test_output[4904] = '{32'h42bad1ed};
test_index[4904] = '{0};
test_input[39240:39247] = '{32'h429fb059, 32'hc2ad989f, 32'h3ec62732, 32'h408c0e94, 32'h42247836, 32'hc1e202ef, 32'hc25a7872, 32'h41b4a6ea};
test_output[4905] = '{32'h429fb059};
test_index[4905] = '{0};
test_input[39248:39255] = '{32'h42b02a26, 32'h426ab009, 32'hc2af72a2, 32'hc2c1a199, 32'hc21a74de, 32'hc1473e8a, 32'hc26ea667, 32'h41f89900};
test_output[4906] = '{32'h42b02a26};
test_index[4906] = '{0};
test_input[39256:39263] = '{32'hc0a8b008, 32'h42bf569e, 32'hc286673f, 32'hc279f4cf, 32'h41207f48, 32'h42c7213d, 32'hc2b0cdf7, 32'h40829560};
test_output[4907] = '{32'h42c7213d};
test_index[4907] = '{5};
test_input[39264:39271] = '{32'h42891894, 32'h41b6971b, 32'hc0cf38d7, 32'hc0d8a1a8, 32'hc2360faf, 32'h4208844c, 32'h41b4474d, 32'hc1e90446};
test_output[4908] = '{32'h42891894};
test_index[4908] = '{0};
test_input[39272:39279] = '{32'h426a933b, 32'hc1125e27, 32'hc269700e, 32'h428ded19, 32'h4295fe01, 32'h41f6a228, 32'hc287f52e, 32'h428ff03e};
test_output[4909] = '{32'h4295fe01};
test_index[4909] = '{4};
test_input[39280:39287] = '{32'h42a032c5, 32'h41c866bc, 32'h42a6732c, 32'h40d14630, 32'hc28dd529, 32'hc171a607, 32'h4235a16b, 32'h41cbe2fb};
test_output[4910] = '{32'h42a6732c};
test_index[4910] = '{2};
test_input[39288:39295] = '{32'hc29da595, 32'h4261d524, 32'hc22360a8, 32'hc24b3dd8, 32'hc2938c84, 32'h429e0696, 32'hc2a5900d, 32'h428d3e40};
test_output[4911] = '{32'h429e0696};
test_index[4911] = '{5};
test_input[39296:39303] = '{32'h40f05f61, 32'h424cf3b0, 32'h42ae795d, 32'hc2b0f43f, 32'h3fcc53ca, 32'h420f7e4f, 32'hc266a862, 32'h42a6c331};
test_output[4912] = '{32'h42ae795d};
test_index[4912] = '{2};
test_input[39304:39311] = '{32'hbf7ceb9f, 32'h42702121, 32'h4295c348, 32'h3f894fb1, 32'h41daec9f, 32'h414054d0, 32'h4222aa3e, 32'hc20a464a};
test_output[4913] = '{32'h4295c348};
test_index[4913] = '{2};
test_input[39312:39319] = '{32'h41aa8b25, 32'h424514e9, 32'h42b92b0c, 32'h4161367a, 32'h42806881, 32'h424d5d17, 32'h42bbc26c, 32'hc2a5986b};
test_output[4914] = '{32'h42bbc26c};
test_index[4914] = '{6};
test_input[39320:39327] = '{32'h42b9f2cc, 32'hc2057462, 32'h426ecf8d, 32'h429c39e1, 32'hc1a1065a, 32'hc1e1bdc6, 32'h420ea524, 32'h3ff41956};
test_output[4915] = '{32'h42b9f2cc};
test_index[4915] = '{0};
test_input[39328:39335] = '{32'h40b2efac, 32'h424208cf, 32'hbe5ba213, 32'hc27fb689, 32'h42b4a5e8, 32'h41ea58c9, 32'hc1bd1ff1, 32'hc28d98f8};
test_output[4916] = '{32'h42b4a5e8};
test_index[4916] = '{4};
test_input[39336:39343] = '{32'h4250684c, 32'hc243d1d4, 32'hc229e0c8, 32'h420d8971, 32'h42afa8fc, 32'h42968ecd, 32'hc254fce9, 32'h42c0c551};
test_output[4917] = '{32'h42c0c551};
test_index[4917] = '{7};
test_input[39344:39351] = '{32'h4205d33d, 32'h42bf6305, 32'hc19ffd58, 32'h4284b0f2, 32'h424196be, 32'hc2a95419, 32'hc1593a6f, 32'h420a4ca3};
test_output[4918] = '{32'h42bf6305};
test_index[4918] = '{1};
test_input[39352:39359] = '{32'hc1b28cda, 32'hc252be84, 32'h41e07360, 32'hc2aaa68e, 32'h42b0d39f, 32'h41958769, 32'h42530f6d, 32'h4285c427};
test_output[4919] = '{32'h42b0d39f};
test_index[4919] = '{4};
test_input[39360:39367] = '{32'h4175a9fc, 32'hc252deb7, 32'hc2bb2ce3, 32'h42a7fca5, 32'h429d4c22, 32'h42ad920c, 32'h429f2b45, 32'hc22f4fd4};
test_output[4920] = '{32'h42ad920c};
test_index[4920] = '{5};
test_input[39368:39375] = '{32'h42242010, 32'hc1f8971a, 32'h4216c078, 32'h42b87228, 32'hc28ef985, 32'hc21cb450, 32'hc2b9ec94, 32'h420146e1};
test_output[4921] = '{32'h42b87228};
test_index[4921] = '{3};
test_input[39376:39383] = '{32'hc262345a, 32'h420bb058, 32'h419d0efc, 32'hc110b111, 32'hc29baafe, 32'hc21eca59, 32'hc0a81bc4, 32'h4235e502};
test_output[4922] = '{32'h4235e502};
test_index[4922] = '{7};
test_input[39384:39391] = '{32'hc2a3e7be, 32'hc20745b7, 32'h42a4d5c5, 32'hc2354579, 32'hc21417f7, 32'h40b8bded, 32'hc241f4ea, 32'h42357f52};
test_output[4923] = '{32'h42a4d5c5};
test_index[4923] = '{2};
test_input[39392:39399] = '{32'hc241e2b4, 32'h42b72e46, 32'hc24ea440, 32'h429bc1a8, 32'h41295b21, 32'hc23e2ef4, 32'h4284abc8, 32'h429699d5};
test_output[4924] = '{32'h42b72e46};
test_index[4924] = '{1};
test_input[39400:39407] = '{32'h429a4e40, 32'hc28d8399, 32'hc1dda074, 32'h41a5dd13, 32'h3fc90c96, 32'h424d1355, 32'h426dde0e, 32'hc2bc8caa};
test_output[4925] = '{32'h429a4e40};
test_index[4925] = '{0};
test_input[39408:39415] = '{32'hc2a15b9f, 32'hc2913505, 32'hc26a2951, 32'hc2aa1a9a, 32'h4021c377, 32'h4271fbd3, 32'h429502f7, 32'h4298a7ee};
test_output[4926] = '{32'h4298a7ee};
test_index[4926] = '{7};
test_input[39416:39423] = '{32'h4211df6d, 32'h4296cf5f, 32'h41718ad8, 32'hc1c2815e, 32'h41bc9ead, 32'h412b00bf, 32'h40c1a9bf, 32'hc2c12bda};
test_output[4927] = '{32'h4296cf5f};
test_index[4927] = '{1};
test_input[39424:39431] = '{32'h41e396ee, 32'hc196d7bc, 32'h42b37ae7, 32'h4207feb4, 32'h4286702e, 32'h429e0395, 32'h428c55f1, 32'h423c5b75};
test_output[4928] = '{32'h42b37ae7};
test_index[4928] = '{2};
test_input[39432:39439] = '{32'hc19c0fa9, 32'hc2813fef, 32'hc2132d0c, 32'h42ba2241, 32'h41cf82b1, 32'hc1896d98, 32'h42ab7ca8, 32'h4277fe2f};
test_output[4929] = '{32'h42ba2241};
test_index[4929] = '{3};
test_input[39440:39447] = '{32'hc28a4a3a, 32'hc03e195a, 32'hc1914f3d, 32'h40dc6f30, 32'hc2550e8c, 32'hc202c5bb, 32'h42515eb0, 32'h4222ad4d};
test_output[4930] = '{32'h42515eb0};
test_index[4930] = '{6};
test_input[39448:39455] = '{32'hc20d2e50, 32'hc1dfd71c, 32'hc1a0d1a0, 32'h412e225e, 32'hc2aa3f41, 32'h429a4cd3, 32'hc2a63b9a, 32'hc2bebe1f};
test_output[4931] = '{32'h429a4cd3};
test_index[4931] = '{5};
test_input[39456:39463] = '{32'hc1f44f90, 32'h42b431f0, 32'hc23a4c6a, 32'h3ecb092d, 32'hc13651b0, 32'h41a8b399, 32'h424f1bf5, 32'h420e200b};
test_output[4932] = '{32'h42b431f0};
test_index[4932] = '{1};
test_input[39464:39471] = '{32'h3f578bb5, 32'h42917f79, 32'hc2ba42e1, 32'hc20bf29d, 32'hc26f3baf, 32'hc2572ffb, 32'h42b47c3e, 32'h429cedb4};
test_output[4933] = '{32'h42b47c3e};
test_index[4933] = '{6};
test_input[39472:39479] = '{32'hc27dfaac, 32'hc21df9cd, 32'h42216404, 32'h41df66d9, 32'hc2a6a6a4, 32'hc2b7a958, 32'hc2a2d93b, 32'hc236842e};
test_output[4934] = '{32'h42216404};
test_index[4934] = '{2};
test_input[39480:39487] = '{32'h42acef4b, 32'hc0827b85, 32'hc2b5367f, 32'h413ecd04, 32'h40da355f, 32'h3f8a0b95, 32'h4207246c, 32'h412c97ab};
test_output[4935] = '{32'h42acef4b};
test_index[4935] = '{0};
test_input[39488:39495] = '{32'hc29df2a4, 32'h41e2bdd6, 32'hc20e8231, 32'hc28b833c, 32'hc1889242, 32'h419ffd93, 32'h42bdae9c, 32'hc2c0ab36};
test_output[4936] = '{32'h42bdae9c};
test_index[4936] = '{6};
test_input[39496:39503] = '{32'h4193e2cf, 32'h422dedf0, 32'h42b157ca, 32'hc270ee6d, 32'hc2c12ed7, 32'h41da4983, 32'hc280ec1c, 32'hc27a2a33};
test_output[4937] = '{32'h42b157ca};
test_index[4937] = '{2};
test_input[39504:39511] = '{32'hc264794b, 32'h4101a25b, 32'hc240a417, 32'h41fa3890, 32'hc2127413, 32'hc1b9e742, 32'h423dd286, 32'h42093bb1};
test_output[4938] = '{32'h423dd286};
test_index[4938] = '{6};
test_input[39512:39519] = '{32'h410ef5d6, 32'hc25428b1, 32'h428ae490, 32'h428c203c, 32'hc28aee3e, 32'hc2a71ea1, 32'h42c3f837, 32'hc1e463b8};
test_output[4939] = '{32'h42c3f837};
test_index[4939] = '{6};
test_input[39520:39527] = '{32'h4201b8a8, 32'h42c49939, 32'hc236ef3d, 32'hc2778c63, 32'hc2b07889, 32'hc2aba217, 32'hc2ab02b8, 32'hc2b2066e};
test_output[4940] = '{32'h42c49939};
test_index[4940] = '{1};
test_input[39528:39535] = '{32'h40d48860, 32'h41321ea0, 32'h41880ff7, 32'h41d88a66, 32'hc22ee14b, 32'h42b2690a, 32'h4056d8a8, 32'hc2ac4c6c};
test_output[4941] = '{32'h42b2690a};
test_index[4941] = '{5};
test_input[39536:39543] = '{32'hc2b0c4d6, 32'hc2b0e7f8, 32'h42b2068f, 32'h42058997, 32'h42357da8, 32'h42a2f235, 32'h427c86bb, 32'h4290d194};
test_output[4942] = '{32'h42b2068f};
test_index[4942] = '{2};
test_input[39544:39551] = '{32'hc1abf9d9, 32'hc2bd1942, 32'hc28630e7, 32'h42acd818, 32'h424ee292, 32'h42b4de5b, 32'hc1ed0a23, 32'h4224cff9};
test_output[4943] = '{32'h42b4de5b};
test_index[4943] = '{5};
test_input[39552:39559] = '{32'hc2c6ce59, 32'hc28d7ca1, 32'h429deec9, 32'hc202f873, 32'hc18fea10, 32'hc297eac1, 32'hbf26d22b, 32'h425e2b6d};
test_output[4944] = '{32'h429deec9};
test_index[4944] = '{2};
test_input[39560:39567] = '{32'h4162c30b, 32'hc28e61da, 32'hc1b1164b, 32'h3e478757, 32'h42a2ae92, 32'h429b89d6, 32'hc13cbe4b, 32'h42430b15};
test_output[4945] = '{32'h42a2ae92};
test_index[4945] = '{4};
test_input[39568:39575] = '{32'hc2252ce2, 32'hc23501c1, 32'hc2bd3dc7, 32'h42a2a620, 32'hc285e7f7, 32'h429b800b, 32'h41493060, 32'hc03957b7};
test_output[4946] = '{32'h42a2a620};
test_index[4946] = '{3};
test_input[39576:39583] = '{32'h42a14a52, 32'hc2ba52c2, 32'h428db32e, 32'h429d442d, 32'h426a99ba, 32'h4202e70d, 32'h42c4868a, 32'h42aca0f5};
test_output[4947] = '{32'h42c4868a};
test_index[4947] = '{6};
test_input[39584:39591] = '{32'h42b60130, 32'h415a7246, 32'hc2c6700c, 32'h4082cf3c, 32'hc19a17fc, 32'h41acc256, 32'h42bc0875, 32'h428f14ed};
test_output[4948] = '{32'h42bc0875};
test_index[4948] = '{6};
test_input[39592:39599] = '{32'h427ec030, 32'hc127ffb3, 32'h4206409a, 32'hc29a34b1, 32'h425b4e5e, 32'h40b0d18f, 32'h41fbc937, 32'hc2b6bb7a};
test_output[4949] = '{32'h427ec030};
test_index[4949] = '{0};
test_input[39600:39607] = '{32'hc2c5a964, 32'h42be3991, 32'h42ad33dc, 32'hc26ed853, 32'hc2b19586, 32'hc1e58152, 32'hc0f1eb14, 32'hc22898b1};
test_output[4950] = '{32'h42be3991};
test_index[4950] = '{1};
test_input[39608:39615] = '{32'hc248f081, 32'hc27313b8, 32'hc2bff452, 32'h42b89e49, 32'h41f820ec, 32'hc12b45b7, 32'h42a48171, 32'h42893c5f};
test_output[4951] = '{32'h42b89e49};
test_index[4951] = '{3};
test_input[39616:39623] = '{32'hc1c14648, 32'h4251e666, 32'h40f74c7d, 32'hc2b9aa12, 32'hc1b18095, 32'h41a9de5d, 32'h42171283, 32'hc2290d34};
test_output[4952] = '{32'h4251e666};
test_index[4952] = '{1};
test_input[39624:39631] = '{32'h40814c3a, 32'hc234a291, 32'hc1293e59, 32'h40d1c87c, 32'hc1d9db88, 32'hc22518ff, 32'h41a44a6b, 32'hc1274851};
test_output[4953] = '{32'h41a44a6b};
test_index[4953] = '{6};
test_input[39632:39639] = '{32'h42a58d0e, 32'hc0067694, 32'hc1dbb665, 32'hc1bae144, 32'h4181cead, 32'hc2905c11, 32'h42958a91, 32'h42b75818};
test_output[4954] = '{32'h42b75818};
test_index[4954] = '{7};
test_input[39640:39647] = '{32'h418af2af, 32'hc1f0346b, 32'hc2849fdf, 32'hc28f9d33, 32'h420abdde, 32'hc23d3c11, 32'h40c8e803, 32'hc20a01c5};
test_output[4955] = '{32'h420abdde};
test_index[4955] = '{4};
test_input[39648:39655] = '{32'h42c11fb3, 32'h422cadb5, 32'hbf1fc353, 32'h425edf2e, 32'hc0143f9b, 32'h419a0073, 32'hc2348393, 32'hc2244788};
test_output[4956] = '{32'h42c11fb3};
test_index[4956] = '{0};
test_input[39656:39663] = '{32'h429ba0d7, 32'h4236b136, 32'h425128e3, 32'h413c171d, 32'h4298fa57, 32'h40ce5fb2, 32'h40cceeb1, 32'hc2903977};
test_output[4957] = '{32'h429ba0d7};
test_index[4957] = '{0};
test_input[39664:39671] = '{32'h41e0c943, 32'h42ac6e73, 32'h427ce106, 32'hc2bfebd5, 32'hc1f7d511, 32'hc1f101e2, 32'h41398d54, 32'hc2bc1f27};
test_output[4958] = '{32'h42ac6e73};
test_index[4958] = '{1};
test_input[39672:39679] = '{32'h42126f41, 32'h41a3032e, 32'hc0910353, 32'hc21be0ec, 32'h426006c1, 32'h4263ccca, 32'h424f7af0, 32'hc270e840};
test_output[4959] = '{32'h4263ccca};
test_index[4959] = '{5};
test_input[39680:39687] = '{32'h42ac7eb4, 32'h40ff1516, 32'h42a9b42e, 32'h42ab004e, 32'hc2651be4, 32'h42b7d367, 32'hc28ffa3f, 32'h425ed803};
test_output[4960] = '{32'h42b7d367};
test_index[4960] = '{5};
test_input[39688:39695] = '{32'h42a7ae5b, 32'hc10b9374, 32'h42b31884, 32'h42a3467c, 32'hbf8de4cb, 32'h4260afd6, 32'hc218b9b9, 32'h429487c3};
test_output[4961] = '{32'h42b31884};
test_index[4961] = '{2};
test_input[39696:39703] = '{32'h41ca8215, 32'h4188b1d6, 32'hc20b0f4d, 32'h4259aa55, 32'h41970f56, 32'h42adaa71, 32'h42615c43, 32'h428ccf15};
test_output[4962] = '{32'h42adaa71};
test_index[4962] = '{5};
test_input[39704:39711] = '{32'h4283a76c, 32'hc2609588, 32'h42331283, 32'h42b0c15e, 32'h42596e51, 32'hc1c337ee, 32'hc2825022, 32'hc0832b01};
test_output[4963] = '{32'h42b0c15e};
test_index[4963] = '{3};
test_input[39712:39719] = '{32'h428867cc, 32'h414924f6, 32'hc28b1328, 32'hc23aa680, 32'hc2c52b8c, 32'h427b3a0f, 32'hc2a9b784, 32'hc19ebc2a};
test_output[4964] = '{32'h428867cc};
test_index[4964] = '{0};
test_input[39720:39727] = '{32'hc200baec, 32'h42bd852d, 32'h417541e7, 32'h423439b6, 32'hc22b3ce1, 32'hc2b94871, 32'hbf275c17, 32'hc204a488};
test_output[4965] = '{32'h42bd852d};
test_index[4965] = '{1};
test_input[39728:39735] = '{32'h3ec46a8f, 32'h428ac88c, 32'h42b5bce7, 32'hc2c6e6d9, 32'h4272e47a, 32'hc22a854e, 32'hc2b216b4, 32'h42bbe310};
test_output[4966] = '{32'h42bbe310};
test_index[4966] = '{7};
test_input[39736:39743] = '{32'hc083325e, 32'h42952ba8, 32'h42a58664, 32'h40ed7cbe, 32'h414a6160, 32'hc1ae9e76, 32'h424c9f4a, 32'hc1abcd9a};
test_output[4967] = '{32'h42a58664};
test_index[4967] = '{2};
test_input[39744:39751] = '{32'h42bed948, 32'h42536d99, 32'h42aa0ae6, 32'h40931d0b, 32'h4146b015, 32'h4139899d, 32'h41c277d0, 32'hc21d44da};
test_output[4968] = '{32'h42bed948};
test_index[4968] = '{0};
test_input[39752:39759] = '{32'h4225af2c, 32'h429302b8, 32'hc2b2688d, 32'h41172c5b, 32'h423a9306, 32'h423fbb7c, 32'hc2592c29, 32'hc0e25113};
test_output[4969] = '{32'h429302b8};
test_index[4969] = '{1};
test_input[39760:39767] = '{32'hc1d65426, 32'hc21e865a, 32'hbfb37bea, 32'h42afd434, 32'h42357f90, 32'hc06dcb6c, 32'h41be022d, 32'h4122e985};
test_output[4970] = '{32'h42afd434};
test_index[4970] = '{3};
test_input[39768:39775] = '{32'h4283d975, 32'hc11dd368, 32'hc1ae3369, 32'h42a9d215, 32'hc286606b, 32'h4156d823, 32'hc1d23278, 32'hc23b8982};
test_output[4971] = '{32'h42a9d215};
test_index[4971] = '{3};
test_input[39776:39783] = '{32'hc29d490a, 32'hc25f4fbc, 32'hc1ea5bca, 32'h41d3276d, 32'h4290b04c, 32'h41dd3955, 32'h3f9507e6, 32'hc15fd0ad};
test_output[4972] = '{32'h4290b04c};
test_index[4972] = '{4};
test_input[39784:39791] = '{32'h41d2c74b, 32'h41a86a4c, 32'hc29a4e10, 32'hc21a9462, 32'hc09f9299, 32'h42a381cf, 32'h42bafc58, 32'hc1263259};
test_output[4973] = '{32'h42bafc58};
test_index[4973] = '{6};
test_input[39792:39799] = '{32'h3f4ff1a2, 32'hc169365b, 32'h421a0458, 32'hc28e15f6, 32'hc2975c1d, 32'h42a1e5b1, 32'h425119de, 32'h4257e8ba};
test_output[4974] = '{32'h42a1e5b1};
test_index[4974] = '{5};
test_input[39800:39807] = '{32'h421708e4, 32'hc24418d7, 32'hc17dcc79, 32'h4261f622, 32'hc28e8bdf, 32'hc1ddc17a, 32'hc22b52d9, 32'hc2162422};
test_output[4975] = '{32'h4261f622};
test_index[4975] = '{3};
test_input[39808:39815] = '{32'hc0ac456f, 32'hc1be8ead, 32'hc287d6d8, 32'h4231af45, 32'h42065e77, 32'hc22b4bd1, 32'hc28661d5, 32'h42665e37};
test_output[4976] = '{32'h42665e37};
test_index[4976] = '{7};
test_input[39816:39823] = '{32'hc291fe63, 32'h42bfa8ca, 32'h42bcae6c, 32'h42b3de6e, 32'hbff173f5, 32'hc2441cd4, 32'h4126c240, 32'h41898430};
test_output[4977] = '{32'h42bfa8ca};
test_index[4977] = '{1};
test_input[39824:39831] = '{32'hc2521c8b, 32'hc280ee72, 32'h42328645, 32'h42626a50, 32'h41ae172e, 32'h41be539a, 32'h4279990e, 32'h4260bee3};
test_output[4978] = '{32'h4279990e};
test_index[4978] = '{6};
test_input[39832:39839] = '{32'hc0cb6789, 32'h4123956a, 32'h4214486d, 32'hc25b3507, 32'hc2a6bf63, 32'hc2715805, 32'h41b01a50, 32'hc1b2392f};
test_output[4979] = '{32'h4214486d};
test_index[4979] = '{2};
test_input[39840:39847] = '{32'hc206a20a, 32'h4182be35, 32'hc16959b0, 32'hc2afd133, 32'hc29d87cd, 32'h426c339d, 32'hc2963ac5, 32'hc233a9c6};
test_output[4980] = '{32'h426c339d};
test_index[4980] = '{5};
test_input[39848:39855] = '{32'h426c9272, 32'hc0e10cbb, 32'hc20fe8cc, 32'h41ad3210, 32'hc283e043, 32'h41fc1486, 32'hc2b7d9d4, 32'hc09d112d};
test_output[4981] = '{32'h426c9272};
test_index[4981] = '{0};
test_input[39856:39863] = '{32'hc23dffb3, 32'hc153571a, 32'h40b6d008, 32'hc113cb0c, 32'h4201b03f, 32'h4245b563, 32'h41b146c6, 32'h42b11fff};
test_output[4982] = '{32'h42b11fff};
test_index[4982] = '{7};
test_input[39864:39871] = '{32'h42baa96b, 32'h415ffb27, 32'hc1c60af0, 32'hc2659c8d, 32'h42a3a870, 32'hc0be3d16, 32'hc28a1bf9, 32'h42967862};
test_output[4983] = '{32'h42baa96b};
test_index[4983] = '{0};
test_input[39872:39879] = '{32'h40aa5627, 32'h423e503b, 32'hc21ae926, 32'hc1ff1f88, 32'h42ada5b0, 32'hc281c9db, 32'hc2a62c05, 32'hc196840d};
test_output[4984] = '{32'h42ada5b0};
test_index[4984] = '{4};
test_input[39880:39887] = '{32'h42808871, 32'h428d0265, 32'hc2948e6b, 32'h42a267ed, 32'h41bfc280, 32'h42550993, 32'hc2855f74, 32'h42945d62};
test_output[4985] = '{32'h42a267ed};
test_index[4985] = '{3};
test_input[39888:39895] = '{32'h421c1a24, 32'hc2906cc3, 32'hc2c76623, 32'hc2617962, 32'h420859e7, 32'h42703abf, 32'h426b0d2f, 32'hc2aaaff0};
test_output[4986] = '{32'h42703abf};
test_index[4986] = '{5};
test_input[39896:39903] = '{32'hc26319ec, 32'h42775779, 32'hc1006bab, 32'hc0a6062f, 32'h40d539cd, 32'hc13096d4, 32'hc293d1a8, 32'h42b64f36};
test_output[4987] = '{32'h42b64f36};
test_index[4987] = '{7};
test_input[39904:39911] = '{32'h42c3a032, 32'hc2367d41, 32'hc2867422, 32'hc1a3194c, 32'h41fe476a, 32'hc2c5173a, 32'h42896985, 32'h4227ffdc};
test_output[4988] = '{32'h42c3a032};
test_index[4988] = '{0};
test_input[39912:39919] = '{32'hc2b804a3, 32'h42b21b16, 32'hc1cf00dc, 32'h41935e44, 32'h422f967c, 32'h41e4dead, 32'h418500af, 32'hc20894ae};
test_output[4989] = '{32'h42b21b16};
test_index[4989] = '{1};
test_input[39920:39927] = '{32'h42419d41, 32'hc23b1baa, 32'h42ab5a6d, 32'hc13e0275, 32'hc110d2d9, 32'hc2b78155, 32'hc2a90ad4, 32'hc197302a};
test_output[4990] = '{32'h42ab5a6d};
test_index[4990] = '{2};
test_input[39928:39935] = '{32'h41bdde0e, 32'hc1c84eb2, 32'hc257a370, 32'hc2896b38, 32'hc1f9d16c, 32'h42a5f0b9, 32'h4243c90b, 32'hc10d1547};
test_output[4991] = '{32'h42a5f0b9};
test_index[4991] = '{5};
test_input[39936:39943] = '{32'h4259705c, 32'h422f9235, 32'hc2a743e0, 32'h41c404fd, 32'h42c3c193, 32'hc2b3c1c8, 32'hc16aa931, 32'h42788a8f};
test_output[4992] = '{32'h42c3c193};
test_index[4992] = '{4};
test_input[39944:39951] = '{32'h42c62d97, 32'hc0a96c53, 32'h42c183f7, 32'h421099f9, 32'h42905f1d, 32'h40a5ce70, 32'h428c8297, 32'hbfd58417};
test_output[4993] = '{32'h42c62d97};
test_index[4993] = '{0};
test_input[39952:39959] = '{32'hc13310eb, 32'h41b6b3f0, 32'hc1df6465, 32'h422a7548, 32'h41ea22bf, 32'h4227d94f, 32'hc1647420, 32'hc28703f7};
test_output[4994] = '{32'h422a7548};
test_index[4994] = '{3};
test_input[39960:39967] = '{32'h4195062f, 32'h421d0179, 32'hc045f66a, 32'hc226eb3d, 32'hc235affd, 32'hc2beec2f, 32'h41cfb029, 32'h41564a74};
test_output[4995] = '{32'h421d0179};
test_index[4995] = '{1};
test_input[39968:39975] = '{32'hc19417a7, 32'h40d9ccd9, 32'h42c690eb, 32'h42b648e0, 32'hc1429941, 32'h41d9094d, 32'hc17af69c, 32'h422df9c5};
test_output[4996] = '{32'h42c690eb};
test_index[4996] = '{2};
test_input[39976:39983] = '{32'h42b8ddb1, 32'hc2436d4d, 32'hc2919084, 32'h42a14749, 32'h425cc536, 32'hbe75cd25, 32'h40a0759f, 32'hc277eba4};
test_output[4997] = '{32'h42b8ddb1};
test_index[4997] = '{0};
test_input[39984:39991] = '{32'h4053d57e, 32'h4225ddbe, 32'h42b2ba72, 32'hc1df52ad, 32'h42899c1d, 32'hc1a82857, 32'hc28d2473, 32'h41026880};
test_output[4998] = '{32'h42b2ba72};
test_index[4998] = '{2};
test_input[39992:39999] = '{32'hc2bff55f, 32'h414ff998, 32'hc26a433b, 32'hc20f2137, 32'h423031fa, 32'h425df90e, 32'h42389bf4, 32'hc22e7eb1};
test_output[4999] = '{32'h425df90e};
test_index[4999] = '{5};
test_input[40000:40007] = '{32'hc2a49cba, 32'h425b494c, 32'h429dd28c, 32'hc2ba998a, 32'hc288acd7, 32'hc23595cf, 32'hc05f44ea, 32'hc2b164cf};
test_output[5000] = '{32'h429dd28c};
test_index[5000] = '{2};
test_input[40008:40015] = '{32'hc2b39407, 32'hc0d67991, 32'h42822833, 32'h41c750ec, 32'h42321d8e, 32'hc2946156, 32'h4294059c, 32'h41ff2df2};
test_output[5001] = '{32'h4294059c};
test_index[5001] = '{6};
test_input[40016:40023] = '{32'hc1ea614d, 32'hc1c67e5b, 32'h42b4f0a7, 32'h422be2ee, 32'hc2bdc9dd, 32'h423b1183, 32'h420a4086, 32'h42878d43};
test_output[5002] = '{32'h42b4f0a7};
test_index[5002] = '{2};
test_input[40024:40031] = '{32'hc26dc781, 32'hc1b913b9, 32'h40c879f6, 32'h4284c695, 32'hc2c45723, 32'hc24fe4ac, 32'hc2925496, 32'hc26dd4b1};
test_output[5003] = '{32'h4284c695};
test_index[5003] = '{3};
test_input[40032:40039] = '{32'hc294cd8a, 32'h4268c796, 32'h4266c96e, 32'h429835ce, 32'h4220913e, 32'h423c417c, 32'hc219015d, 32'h4129579b};
test_output[5004] = '{32'h429835ce};
test_index[5004] = '{3};
test_input[40040:40047] = '{32'h41aabd08, 32'h41f231c3, 32'hc27e92d4, 32'hc282d789, 32'h42474135, 32'h42b434f6, 32'hc284357d, 32'hc26ba8f1};
test_output[5005] = '{32'h42b434f6};
test_index[5005] = '{5};
test_input[40048:40055] = '{32'hc2c1e96a, 32'h426b5485, 32'h424fb407, 32'hc29977b0, 32'hc142514a, 32'hc1ed36a7, 32'hbfac6baf, 32'hc20bfdce};
test_output[5006] = '{32'h426b5485};
test_index[5006] = '{1};
test_input[40056:40063] = '{32'hc101b2b6, 32'h42916913, 32'hc29317b1, 32'hc27d907d, 32'h4125bc78, 32'h429dc19f, 32'h422a661a, 32'h42749a04};
test_output[5007] = '{32'h429dc19f};
test_index[5007] = '{5};
test_input[40064:40071] = '{32'h407ee4c8, 32'h42adff3e, 32'hc218b533, 32'h42c4e572, 32'hc1d70c6f, 32'hc29cddc2, 32'hc28b8bcf, 32'hc295a339};
test_output[5008] = '{32'h42c4e572};
test_index[5008] = '{3};
test_input[40072:40079] = '{32'hc218ea46, 32'hc25f5079, 32'hc29425f2, 32'h4290a234, 32'hc24eaabe, 32'hc296ba1f, 32'hc2828e82, 32'hc2bd902d};
test_output[5009] = '{32'h4290a234};
test_index[5009] = '{3};
test_input[40080:40087] = '{32'hbf13f48e, 32'hc2ab12e4, 32'h4287c6e6, 32'hc0874442, 32'h419765ac, 32'h4298de23, 32'h419e1c6f, 32'hc28f72f0};
test_output[5010] = '{32'h4298de23};
test_index[5010] = '{5};
test_input[40088:40095] = '{32'hc2bdd821, 32'hc2bcdb46, 32'h42b301b1, 32'hc12d538c, 32'hc188590b, 32'h41b44407, 32'hc276e1d4, 32'hc20dda82};
test_output[5011] = '{32'h42b301b1};
test_index[5011] = '{2};
test_input[40096:40103] = '{32'hc233bac4, 32'h42a7c1c6, 32'h420096be, 32'h4258b278, 32'h42b23de0, 32'h3f5d7091, 32'h41812599, 32'h4235fb26};
test_output[5012] = '{32'h42b23de0};
test_index[5012] = '{4};
test_input[40104:40111] = '{32'hc2adcb41, 32'h42702cbc, 32'h41dd48ce, 32'hc2bd358f, 32'hc28b2fe5, 32'h403f20ab, 32'hc2c579da, 32'hc2bc603a};
test_output[5013] = '{32'h42702cbc};
test_index[5013] = '{1};
test_input[40112:40119] = '{32'h3fc64485, 32'h42900a79, 32'hc2950dfb, 32'hc28f7d84, 32'h40f12492, 32'h4150f8cf, 32'hc2c1f86c, 32'h42b7ec3e};
test_output[5014] = '{32'h42b7ec3e};
test_index[5014] = '{7};
test_input[40120:40127] = '{32'hc24b5b88, 32'hc2aea13a, 32'hc2a79d7b, 32'h42207405, 32'hc28ead33, 32'h42b3e474, 32'hc2c54489, 32'h4224da47};
test_output[5015] = '{32'h42b3e474};
test_index[5015] = '{5};
test_input[40128:40135] = '{32'hc1ff7c05, 32'hc1ed0faa, 32'hc265660c, 32'h41611bcf, 32'h403b84b5, 32'h42852a9b, 32'hbf3cadb1, 32'hc23be6d4};
test_output[5016] = '{32'h42852a9b};
test_index[5016] = '{5};
test_input[40136:40143] = '{32'h4176ee94, 32'h420f705b, 32'h4238b647, 32'hc29c9ae5, 32'hc253334b, 32'hc2b95f00, 32'h429182bf, 32'h429259bd};
test_output[5017] = '{32'h429259bd};
test_index[5017] = '{7};
test_input[40144:40151] = '{32'hc1d8afb1, 32'hc2b86067, 32'h4138d6d9, 32'h42a158f6, 32'h42a43723, 32'h40f86343, 32'h42add375, 32'hbfbf1ad7};
test_output[5018] = '{32'h42add375};
test_index[5018] = '{6};
test_input[40152:40159] = '{32'h41a5be0f, 32'hc2043782, 32'hc2049d87, 32'h42a8c005, 32'h429c68e1, 32'hc0f5759d, 32'hc2b5c690, 32'h420befce};
test_output[5019] = '{32'h42a8c005};
test_index[5019] = '{3};
test_input[40160:40167] = '{32'h42113cca, 32'h416c8cd2, 32'h41f96382, 32'h428bf713, 32'h40ea59ed, 32'h42b282d8, 32'h41b82bce, 32'hc1a3c9ed};
test_output[5020] = '{32'h42b282d8};
test_index[5020] = '{5};
test_input[40168:40175] = '{32'h4248ef0e, 32'h4282981c, 32'hc20f2fc4, 32'hc25b9c4d, 32'hc2c4c18c, 32'h42a6898e, 32'hc2b294d7, 32'hc2a716d6};
test_output[5021] = '{32'h42a6898e};
test_index[5021] = '{5};
test_input[40176:40183] = '{32'h429e27c3, 32'hc25237fa, 32'h4116fc72, 32'h42bede84, 32'hc2c21f23, 32'h4235d908, 32'hc27db5f9, 32'h40a19813};
test_output[5022] = '{32'h42bede84};
test_index[5022] = '{3};
test_input[40184:40191] = '{32'hc1db9121, 32'h420d188e, 32'h4204a5f5, 32'hc242d501, 32'h42ba8d52, 32'h42c40e24, 32'hc1cb1bf0, 32'hc26ad042};
test_output[5023] = '{32'h42c40e24};
test_index[5023] = '{5};
test_input[40192:40199] = '{32'h42a5ca00, 32'hc10b8b23, 32'h3e2e2d0f, 32'h411c3b5f, 32'hc2269b98, 32'hc1abca77, 32'hc2b623e3, 32'hc1f22425};
test_output[5024] = '{32'h42a5ca00};
test_index[5024] = '{0};
test_input[40200:40207] = '{32'hc2af5372, 32'hc171e3c7, 32'h41560eb8, 32'h422f0e82, 32'hc2aa137d, 32'h4276cd2a, 32'hc2ad2b04, 32'h42b9e7a3};
test_output[5025] = '{32'h42b9e7a3};
test_index[5025] = '{7};
test_input[40208:40215] = '{32'hc1c919a0, 32'h42b4b9e9, 32'hc0efd75c, 32'hc25d2ef3, 32'hc25e93f2, 32'h422b6edc, 32'hc114d5fc, 32'hc29c5550};
test_output[5026] = '{32'h42b4b9e9};
test_index[5026] = '{1};
test_input[40216:40223] = '{32'h41a3f4ec, 32'h427ab2a7, 32'h412bf26b, 32'h4206922f, 32'h4203f768, 32'hc28ae9cc, 32'hc1b70369, 32'h428273fe};
test_output[5027] = '{32'h428273fe};
test_index[5027] = '{7};
test_input[40224:40231] = '{32'h4071c2ac, 32'hc2710731, 32'hc2c21a0c, 32'h4218c863, 32'hc26fae88, 32'hc254178b, 32'h42c2df01, 32'hc2678409};
test_output[5028] = '{32'h42c2df01};
test_index[5028] = '{6};
test_input[40232:40239] = '{32'h42829c4e, 32'h42814467, 32'h4210b357, 32'hc23f6a9f, 32'h421e2be1, 32'h42600a10, 32'hc1ebacfa, 32'hc29ef7e7};
test_output[5029] = '{32'h42829c4e};
test_index[5029] = '{0};
test_input[40240:40247] = '{32'h429e0337, 32'hc2b47bc0, 32'h42acf820, 32'hc1327799, 32'h42b124a7, 32'hc1ddb056, 32'h42a9b928, 32'hc12d5bf1};
test_output[5030] = '{32'h42b124a7};
test_index[5030] = '{4};
test_input[40248:40255] = '{32'hc1e099d6, 32'hc24f4eeb, 32'hc29770d7, 32'h408cc0b0, 32'hc1e5171e, 32'hc09abb42, 32'hc21ba8e1, 32'h42188006};
test_output[5031] = '{32'h42188006};
test_index[5031] = '{7};
test_input[40256:40263] = '{32'hc21371e2, 32'hc2b9e15b, 32'hc1b8a1bd, 32'hc29fc96e, 32'h42330cf9, 32'h42301210, 32'h42363940, 32'hc29f688e};
test_output[5032] = '{32'h42363940};
test_index[5032] = '{6};
test_input[40264:40271] = '{32'h422f35d7, 32'hc28ac973, 32'hc2b1c09d, 32'h423ac003, 32'hc28e5f88, 32'h414730bd, 32'h428e749a, 32'h42b8a5d0};
test_output[5033] = '{32'h42b8a5d0};
test_index[5033] = '{7};
test_input[40272:40279] = '{32'hc005bb88, 32'hc2882254, 32'h42a1d149, 32'h429c9cf3, 32'hc25b035e, 32'h42b6ea44, 32'h4233c3d1, 32'h42964922};
test_output[5034] = '{32'h42b6ea44};
test_index[5034] = '{5};
test_input[40280:40287] = '{32'hc2a5f48d, 32'h42ae3e7d, 32'hc29843cd, 32'h41b68519, 32'hc2c50079, 32'h42637dba, 32'h41718f98, 32'h426c253f};
test_output[5035] = '{32'h42ae3e7d};
test_index[5035] = '{1};
test_input[40288:40295] = '{32'hc24d87d4, 32'h425bb39b, 32'h41d6c67c, 32'hc17839ab, 32'h429e369d, 32'hc29d6441, 32'h4156f9ad, 32'hc232f409};
test_output[5036] = '{32'h429e369d};
test_index[5036] = '{4};
test_input[40296:40303] = '{32'hc202529c, 32'hc1b5ae88, 32'h41a782ff, 32'hc20e1587, 32'hc0075664, 32'hc01e0bd2, 32'h428d4847, 32'hc2c5145d};
test_output[5037] = '{32'h428d4847};
test_index[5037] = '{6};
test_input[40304:40311] = '{32'hc2bd1147, 32'h41f1e95e, 32'h4276468e, 32'h42b66fd3, 32'hc132d6e8, 32'hc223e9f0, 32'h42131fc8, 32'h4285c30a};
test_output[5038] = '{32'h42b66fd3};
test_index[5038] = '{3};
test_input[40312:40319] = '{32'h42a7e17f, 32'h4280690a, 32'hc22d7dfe, 32'h42af363f, 32'hc1f97d62, 32'hc2c00121, 32'hc20fbfb0, 32'hc290213c};
test_output[5039] = '{32'h42af363f};
test_index[5039] = '{3};
test_input[40320:40327] = '{32'hc2acd159, 32'h41fa32c0, 32'h40c91f76, 32'hc0be0e74, 32'hc2a11bf1, 32'hc27e7f98, 32'hc2c26166, 32'h3f577939};
test_output[5040] = '{32'h41fa32c0};
test_index[5040] = '{1};
test_input[40328:40335] = '{32'h42613b20, 32'h417fd25c, 32'h4207994e, 32'hc1ee6f7b, 32'hc2975489, 32'hc1acf2c5, 32'h41422349, 32'hc24fe319};
test_output[5041] = '{32'h42613b20};
test_index[5041] = '{0};
test_input[40336:40343] = '{32'h429f8b72, 32'hc15d128d, 32'hc23b884e, 32'hc294b44b, 32'hc1b7bd74, 32'h4298245b, 32'hc24d132f, 32'hc2aeaffc};
test_output[5042] = '{32'h429f8b72};
test_index[5042] = '{0};
test_input[40344:40351] = '{32'h418f28cf, 32'h41b3bde9, 32'hc244c490, 32'h424fa450, 32'h42183b5a, 32'hc238b459, 32'hc03f4b54, 32'h416c6db3};
test_output[5043] = '{32'h424fa450};
test_index[5043] = '{3};
test_input[40352:40359] = '{32'h4277f677, 32'hc149f659, 32'hc2859cd6, 32'hc298adab, 32'h42c725a2, 32'h411fd54e, 32'h415f6847, 32'h429dea66};
test_output[5044] = '{32'h42c725a2};
test_index[5044] = '{4};
test_input[40360:40367] = '{32'hc2491119, 32'hc2a4694c, 32'hc28882ff, 32'hc2595fc3, 32'h4244d7ed, 32'hc1f98793, 32'h426d181e, 32'hc19155c5};
test_output[5045] = '{32'h426d181e};
test_index[5045] = '{6};
test_input[40368:40375] = '{32'hc210232f, 32'h40a32329, 32'h4255e7ae, 32'h41cf3cb7, 32'h42876146, 32'h4292e57e, 32'h42acf90d, 32'hc2b24699};
test_output[5046] = '{32'h42acf90d};
test_index[5046] = '{6};
test_input[40376:40383] = '{32'h4292e258, 32'hc285dce0, 32'h4295fc12, 32'h41b1dbee, 32'h428e28c2, 32'h41b780e7, 32'h41d96cac, 32'hc29aff36};
test_output[5047] = '{32'h4295fc12};
test_index[5047] = '{2};
test_input[40384:40391] = '{32'hc277dd9d, 32'h42106181, 32'h4248ec57, 32'hc1eebbde, 32'hc1d1048f, 32'hc2a03038, 32'hc2c5638b, 32'h42c178a2};
test_output[5048] = '{32'h42c178a2};
test_index[5048] = '{7};
test_input[40392:40399] = '{32'h41978de1, 32'hc2c1d25e, 32'hc1f5fe38, 32'hc2266741, 32'h41b4a0f2, 32'hc23efeb7, 32'hc2950369, 32'h41dfeeea};
test_output[5049] = '{32'h41dfeeea};
test_index[5049] = '{7};
test_input[40400:40407] = '{32'hc239b7b0, 32'h421d2fc6, 32'h41594c70, 32'hc1d39f39, 32'h4298ae61, 32'hc294d275, 32'hc2c53e89, 32'h42b58b49};
test_output[5050] = '{32'h42b58b49};
test_index[5050] = '{7};
test_input[40408:40415] = '{32'hc26ee57e, 32'h420a2745, 32'hc28e41c1, 32'hc1b24151, 32'h42c49687, 32'h40d2e8a0, 32'hc20428b8, 32'hc2c30555};
test_output[5051] = '{32'h42c49687};
test_index[5051] = '{4};
test_input[40416:40423] = '{32'hc225d257, 32'h429ffa16, 32'hc233af8b, 32'h41c175f2, 32'h42c2b7ba, 32'h42336308, 32'hc2bb34e3, 32'hc093f626};
test_output[5052] = '{32'h42c2b7ba};
test_index[5052] = '{4};
test_input[40424:40431] = '{32'hc2ba93eb, 32'hc18b69d6, 32'h42997b57, 32'hc2b28c0c, 32'h42258a2d, 32'hc2a93061, 32'hc261863b, 32'hc2068569};
test_output[5053] = '{32'h42997b57};
test_index[5053] = '{2};
test_input[40432:40439] = '{32'h41854c06, 32'hc2c6a612, 32'hc0108e25, 32'h420a67d6, 32'h42785cfe, 32'h4103fca1, 32'h42af3566, 32'h42250037};
test_output[5054] = '{32'h42af3566};
test_index[5054] = '{6};
test_input[40440:40447] = '{32'h404abe6c, 32'hc2a68183, 32'hc26368c7, 32'hc2c4187b, 32'h428c1272, 32'h417ae3c4, 32'h42a36397, 32'h419974ea};
test_output[5055] = '{32'h42a36397};
test_index[5055] = '{6};
test_input[40448:40455] = '{32'hc2bcfa7e, 32'hc28fac8c, 32'h42a8fa65, 32'hc2c25a4b, 32'h41c5fc05, 32'hc0748403, 32'hc251ebbb, 32'h423c4a12};
test_output[5056] = '{32'h42a8fa65};
test_index[5056] = '{2};
test_input[40456:40463] = '{32'h429c32c9, 32'h4000e6cf, 32'hc29e8da9, 32'hc29fbe1d, 32'hc1e215fa, 32'h42baaa85, 32'h429502af, 32'h42c044bf};
test_output[5057] = '{32'h42c044bf};
test_index[5057] = '{7};
test_input[40464:40471] = '{32'hc18fa8fe, 32'hc2ae2aef, 32'h4021154e, 32'h425a6c95, 32'h419e3bde, 32'hc2917217, 32'h428d4850, 32'hc29c3140};
test_output[5058] = '{32'h428d4850};
test_index[5058] = '{6};
test_input[40472:40479] = '{32'hc1c9b646, 32'h4190b10f, 32'h41cbfa84, 32'h4248fd9c, 32'h41a15e28, 32'h429600ac, 32'h422f6c5f, 32'hc2c2129a};
test_output[5059] = '{32'h429600ac};
test_index[5059] = '{5};
test_input[40480:40487] = '{32'h40dd4ab1, 32'hc1d956ae, 32'hc299d1d8, 32'hc2108703, 32'h428cce5a, 32'hc2968b3d, 32'h414f8427, 32'hc202099f};
test_output[5060] = '{32'h428cce5a};
test_index[5060] = '{4};
test_input[40488:40495] = '{32'h429080d8, 32'h42bc34a8, 32'h42730797, 32'h41d2eb7a, 32'hc18f7318, 32'h414ca561, 32'hc21f0c8c, 32'hc284a6ed};
test_output[5061] = '{32'h42bc34a8};
test_index[5061] = '{1};
test_input[40496:40503] = '{32'hc28ba2b9, 32'h42023b43, 32'hbfd5a6b2, 32'hbfa17ef7, 32'hc1669333, 32'hc26e11c7, 32'hc1f94092, 32'h42393090};
test_output[5062] = '{32'h42393090};
test_index[5062] = '{7};
test_input[40504:40511] = '{32'hc22150a9, 32'h426b66fb, 32'h4209adb9, 32'h42a504b7, 32'hc204e7fb, 32'hc165e347, 32'hc155387b, 32'h42a5e715};
test_output[5063] = '{32'h42a5e715};
test_index[5063] = '{7};
test_input[40512:40519] = '{32'hc2223e65, 32'hc26aea0a, 32'h4256c095, 32'hc296ed55, 32'hc25553cc, 32'h42086528, 32'h41b64684, 32'hc2c0139f};
test_output[5064] = '{32'h4256c095};
test_index[5064] = '{2};
test_input[40520:40527] = '{32'hc1eb02fd, 32'hc23a3742, 32'h429d73ce, 32'hc2215a99, 32'h4239383d, 32'h42b2854a, 32'h42aee547, 32'h42940bef};
test_output[5065] = '{32'h42b2854a};
test_index[5065] = '{5};
test_input[40528:40535] = '{32'hc2927bfa, 32'hc2975e5c, 32'h42a169ff, 32'hc2bc13d5, 32'h41358626, 32'h429df229, 32'h41b7c0af, 32'hc20b85a0};
test_output[5066] = '{32'h42a169ff};
test_index[5066] = '{2};
test_input[40536:40543] = '{32'hc215319c, 32'hc24194cf, 32'h4252d977, 32'h428d9ba3, 32'hc262b97d, 32'h3fb3091e, 32'hc28951c6, 32'hc2801888};
test_output[5067] = '{32'h428d9ba3};
test_index[5067] = '{3};
test_input[40544:40551] = '{32'h4284bbcb, 32'h4209b174, 32'h42c1a1a6, 32'hc255e4e6, 32'hc064cbcc, 32'hc2c1084f, 32'h4107ba34, 32'hc2c239c1};
test_output[5068] = '{32'h42c1a1a6};
test_index[5068] = '{2};
test_input[40552:40559] = '{32'hc20e41fa, 32'h41415e3a, 32'h4232e1d1, 32'h42bc7404, 32'hc22d8dfa, 32'h429e15cf, 32'h40e763b1, 32'hc19971b9};
test_output[5069] = '{32'h42bc7404};
test_index[5069] = '{3};
test_input[40560:40567] = '{32'h4276da14, 32'h42513a7e, 32'hc220bb6f, 32'hc18cbbbb, 32'hc298f034, 32'h423aa679, 32'hc28b4a2f, 32'h41465f61};
test_output[5070] = '{32'h4276da14};
test_index[5070] = '{0};
test_input[40568:40575] = '{32'hc28065ea, 32'hc28fd982, 32'h425a2855, 32'h42c1b3d9, 32'h425393a1, 32'h429ce922, 32'hc21c61bd, 32'hc275ea9a};
test_output[5071] = '{32'h42c1b3d9};
test_index[5071] = '{3};
test_input[40576:40583] = '{32'hc08a42f7, 32'hc2ab4e58, 32'h4292208c, 32'h42b39dd4, 32'h42bb98eb, 32'hc015b9b0, 32'hc28d32f1, 32'h420f3876};
test_output[5072] = '{32'h42bb98eb};
test_index[5072] = '{4};
test_input[40584:40591] = '{32'hc217f9d6, 32'h421d2897, 32'h40bafb96, 32'hc230930f, 32'hc292d9fe, 32'h426b19de, 32'h407add34, 32'hc29ef4f6};
test_output[5073] = '{32'h426b19de};
test_index[5073] = '{5};
test_input[40592:40599] = '{32'hc22d92d8, 32'h41a46941, 32'hc26d9247, 32'hc19fa67b, 32'hc281dd3b, 32'h428ee61b, 32'h428a7b68, 32'h413d1ecd};
test_output[5074] = '{32'h428ee61b};
test_index[5074] = '{5};
test_input[40600:40607] = '{32'hc1764c37, 32'h42c488c9, 32'h41883667, 32'hc2b7e329, 32'h4290f645, 32'h42a1d074, 32'hc2890a99, 32'h42101b56};
test_output[5075] = '{32'h42c488c9};
test_index[5075] = '{1};
test_input[40608:40615] = '{32'hc22b5e29, 32'hc15571cd, 32'h42868b7f, 32'h4286c4fa, 32'hc28daeee, 32'h4285ed73, 32'h41daafd7, 32'hc25d10b6};
test_output[5076] = '{32'h4286c4fa};
test_index[5076] = '{3};
test_input[40616:40623] = '{32'hc2ae9aa2, 32'h41815af6, 32'h42abd418, 32'hc0e1f062, 32'hc26cced0, 32'h42014061, 32'hc26817ab, 32'hc2adeae7};
test_output[5077] = '{32'h42abd418};
test_index[5077] = '{2};
test_input[40624:40631] = '{32'h421132cc, 32'h418dd037, 32'h4296810c, 32'h4118bb39, 32'hc24cc7c7, 32'h4268e96a, 32'hc14bea4d, 32'h40dec53a};
test_output[5078] = '{32'h4296810c};
test_index[5078] = '{2};
test_input[40632:40639] = '{32'hc200a6da, 32'hc21931cd, 32'hc2b5c023, 32'h42c13920, 32'hc282f7e5, 32'h42590fd5, 32'h42551244, 32'hc2751fde};
test_output[5079] = '{32'h42c13920};
test_index[5079] = '{3};
test_input[40640:40647] = '{32'hc1f4c4fb, 32'h42b4e93e, 32'hc29e63a9, 32'h42bcae21, 32'hc23ccee8, 32'h41ce0a41, 32'h42a302ec, 32'hc19452d3};
test_output[5080] = '{32'h42bcae21};
test_index[5080] = '{3};
test_input[40648:40655] = '{32'h42a3ff5b, 32'hc1666bff, 32'h41ce4a03, 32'hc2899c4d, 32'h40016766, 32'hc2aef47e, 32'h41e3da27, 32'h42aa3bb2};
test_output[5081] = '{32'h42aa3bb2};
test_index[5081] = '{7};
test_input[40656:40663] = '{32'hc21b11a8, 32'hc2a41241, 32'h413059fc, 32'h42254c11, 32'h422e53e7, 32'h4298a148, 32'hc2a0741d, 32'hc2b386f7};
test_output[5082] = '{32'h4298a148};
test_index[5082] = '{5};
test_input[40664:40671] = '{32'hbfd85878, 32'hc21b56fe, 32'hc274f04e, 32'hc28ecd64, 32'h4292b532, 32'h42a08deb, 32'hc2b45a21, 32'hc0e5685a};
test_output[5083] = '{32'h42a08deb};
test_index[5083] = '{5};
test_input[40672:40679] = '{32'h41754207, 32'h41616276, 32'hc0cc6941, 32'h4225e48f, 32'h413696b3, 32'hc1fb4c66, 32'hc1f6c14a, 32'hc2058d30};
test_output[5084] = '{32'h4225e48f};
test_index[5084] = '{3};
test_input[40680:40687] = '{32'hc2c66b3e, 32'hc2b2da48, 32'hc2384f6d, 32'hc2a44bf1, 32'hc28fda9a, 32'hc07bbfe5, 32'h42b8b1a9, 32'h42815366};
test_output[5085] = '{32'h42b8b1a9};
test_index[5085] = '{6};
test_input[40688:40695] = '{32'h42983012, 32'hc1a61483, 32'h423aaa23, 32'h42a45379, 32'h41c8deec, 32'h42973711, 32'h4196db15, 32'hbf4b977e};
test_output[5086] = '{32'h42a45379};
test_index[5086] = '{3};
test_input[40696:40703] = '{32'hc2694567, 32'h42be5fc6, 32'h4179d0df, 32'h4163c0e4, 32'h4217a969, 32'h41a37408, 32'hc2c74560, 32'hc2be8447};
test_output[5087] = '{32'h42be5fc6};
test_index[5087] = '{1};
test_input[40704:40711] = '{32'hc221e5d9, 32'hbfdd4afb, 32'h41ea1949, 32'hc2aa1a2f, 32'h41c69f07, 32'hc1a5c72b, 32'h42b37a09, 32'h410bdb88};
test_output[5088] = '{32'h42b37a09};
test_index[5088] = '{6};
test_input[40712:40719] = '{32'hc1d2035c, 32'h41b9ba7c, 32'h42af8631, 32'hc1e1a8b1, 32'h42a783dd, 32'hc29eafc1, 32'h41a74809, 32'h42935945};
test_output[5089] = '{32'h42af8631};
test_index[5089] = '{2};
test_input[40720:40727] = '{32'h42275d22, 32'h41b65dc2, 32'hc279e7e6, 32'hc186308a, 32'h42c6169c, 32'hc2901f63, 32'h4297f72d, 32'h420b1b08};
test_output[5090] = '{32'h42c6169c};
test_index[5090] = '{4};
test_input[40728:40735] = '{32'hc2988809, 32'hc275caa3, 32'hc27bcbaf, 32'h427843ca, 32'hc2c7b635, 32'h4234380a, 32'hc24d99b1, 32'h416b89df};
test_output[5091] = '{32'h427843ca};
test_index[5091] = '{3};
test_input[40736:40743] = '{32'hc19d8aa1, 32'hc20d0853, 32'hc149cea8, 32'h42c44304, 32'hc1cbc902, 32'hc1c20efc, 32'hc2886947, 32'h422725d2};
test_output[5092] = '{32'h42c44304};
test_index[5092] = '{3};
test_input[40744:40751] = '{32'h41bd61a2, 32'hc1f91577, 32'hc2b99b09, 32'h42baf285, 32'h42526a4b, 32'h426923fa, 32'hc2694e42, 32'hc28ea7e2};
test_output[5093] = '{32'h42baf285};
test_index[5093] = '{3};
test_input[40752:40759] = '{32'hc21a5b8d, 32'hc2c1dbc6, 32'h4211ec25, 32'hc229a804, 32'hc1ad20e4, 32'hc1dd8dd5, 32'h42983ada, 32'hc2a99f9c};
test_output[5094] = '{32'h42983ada};
test_index[5094] = '{6};
test_input[40760:40767] = '{32'hc19f46a3, 32'hc185fb49, 32'hc283f5d2, 32'hc209f5b8, 32'hc2b22c21, 32'hc297ae44, 32'hc1293401, 32'h4261f9cc};
test_output[5095] = '{32'h4261f9cc};
test_index[5095] = '{7};
test_input[40768:40775] = '{32'hc272f417, 32'hc2bc035a, 32'hc1fcf8d1, 32'hc2a9dc05, 32'hc2b0c0f1, 32'hc05619a1, 32'hc2b2cba4, 32'h41d20f22};
test_output[5096] = '{32'h41d20f22};
test_index[5096] = '{7};
test_input[40776:40783] = '{32'h40b9f8bd, 32'hc2ac6406, 32'h428dbbd4, 32'h4200d6e2, 32'hc2bbc94f, 32'hc2a25c0c, 32'hc2ac799a, 32'h429dca1f};
test_output[5097] = '{32'h429dca1f};
test_index[5097] = '{7};
test_input[40784:40791] = '{32'h3ffae74a, 32'h4105c80a, 32'h429e8393, 32'hc215f74c, 32'h428c6282, 32'hc1a57f60, 32'h4289edb7, 32'h42aa110b};
test_output[5098] = '{32'h42aa110b};
test_index[5098] = '{7};
test_input[40792:40799] = '{32'hc0d65c1c, 32'h41ef8b3d, 32'hc27a472b, 32'h42c6655b, 32'hbf75938a, 32'hc2a71cc6, 32'h41d22f7b, 32'hc24b8747};
test_output[5099] = '{32'h42c6655b};
test_index[5099] = '{3};
test_input[40800:40807] = '{32'h42704284, 32'h42c3084c, 32'hc29fb567, 32'h4233276a, 32'hc28b6bcb, 32'h42235035, 32'hbf28b3b9, 32'hc187b3ab};
test_output[5100] = '{32'h42c3084c};
test_index[5100] = '{1};
test_input[40808:40815] = '{32'hc222f065, 32'h41c982de, 32'h42b0cb34, 32'hc2b114bc, 32'h41b34477, 32'hc16e8e2e, 32'h42a1304a, 32'hc0ce8b98};
test_output[5101] = '{32'h42b0cb34};
test_index[5101] = '{2};
test_input[40816:40823] = '{32'hc2411287, 32'h422ad736, 32'h419acaf1, 32'hc2a8ea7c, 32'hc1d72d26, 32'h42532af9, 32'h42acb974, 32'h41adac21};
test_output[5102] = '{32'h42acb974};
test_index[5102] = '{6};
test_input[40824:40831] = '{32'hc1358b49, 32'h4189ff49, 32'hc232072c, 32'h4269a9fb, 32'h415a9ac6, 32'h42c23fd9, 32'h42c39d57, 32'hc2a80abc};
test_output[5103] = '{32'h42c39d57};
test_index[5103] = '{6};
test_input[40832:40839] = '{32'h4219d41f, 32'hc2223b90, 32'h42b5a0fd, 32'h418fc586, 32'hbf061b89, 32'h42302313, 32'h419b2c03, 32'hc1801421};
test_output[5104] = '{32'h42b5a0fd};
test_index[5104] = '{2};
test_input[40840:40847] = '{32'hc1fd5c64, 32'h41a0694b, 32'h4271b2ec, 32'h4281d0a0, 32'hc22e3acb, 32'h41ab6fc7, 32'h429fe9ad, 32'h4227289d};
test_output[5105] = '{32'h429fe9ad};
test_index[5105] = '{6};
test_input[40848:40855] = '{32'h41136b9c, 32'h421ca071, 32'h42bc6ac9, 32'h426811ef, 32'h41bfdad9, 32'hc244dcd6, 32'hc2965a1a, 32'hc12ff109};
test_output[5106] = '{32'h42bc6ac9};
test_index[5106] = '{2};
test_input[40856:40863] = '{32'h42a899ad, 32'h42bf88d7, 32'h426557a8, 32'hc22df0c2, 32'hc25b4d3b, 32'h4019ef06, 32'h4204ff03, 32'h4246a8de};
test_output[5107] = '{32'h42bf88d7};
test_index[5107] = '{1};
test_input[40864:40871] = '{32'h428628a9, 32'hc22bd16b, 32'h42a3884e, 32'h42990a46, 32'h420372f6, 32'hc258e693, 32'h4274d2f7, 32'hc17cae67};
test_output[5108] = '{32'h42a3884e};
test_index[5108] = '{2};
test_input[40872:40879] = '{32'h42308b4b, 32'hc23405cd, 32'h4296b42f, 32'hbffc7a6a, 32'hc282a9e8, 32'hc142c4b5, 32'h42035122, 32'hc2bcb38d};
test_output[5109] = '{32'h4296b42f};
test_index[5109] = '{2};
test_input[40880:40887] = '{32'hc10ae2b1, 32'hc2b1fce4, 32'h426e8636, 32'hc225c288, 32'h421d3343, 32'hc2603790, 32'hc24fec2a, 32'h426118ec};
test_output[5110] = '{32'h426e8636};
test_index[5110] = '{2};
test_input[40888:40895] = '{32'h41d47dd5, 32'h423f1fc2, 32'h42999d15, 32'h4165711c, 32'h422f2a9f, 32'h425274d9, 32'h4283564e, 32'h41f182b1};
test_output[5111] = '{32'h42999d15};
test_index[5111] = '{2};
test_input[40896:40903] = '{32'hc094d4e1, 32'h42021b02, 32'h42248e44, 32'hc1339ed7, 32'hc2bcc1f2, 32'hc2a0c4ee, 32'h4004495d, 32'h428f76c2};
test_output[5112] = '{32'h428f76c2};
test_index[5112] = '{7};
test_input[40904:40911] = '{32'hc2276c18, 32'h42011044, 32'hc089e09b, 32'hc236512a, 32'h42159f9a, 32'hc2ae24bc, 32'hc1e55706, 32'hc2867a0c};
test_output[5113] = '{32'h42159f9a};
test_index[5113] = '{4};
test_input[40912:40919] = '{32'h42b1367c, 32'hc222b18c, 32'hc159fdb0, 32'hc2a3ba36, 32'h42916be8, 32'hc2b19349, 32'hc2a389fb, 32'hc1d6f2d7};
test_output[5114] = '{32'h42b1367c};
test_index[5114] = '{0};
test_input[40920:40927] = '{32'hc28e4846, 32'h411aefe2, 32'hc1cb37d6, 32'h42715b11, 32'h41aa51c1, 32'h421b6a14, 32'hbfc5a009, 32'hc1e99e00};
test_output[5115] = '{32'h42715b11};
test_index[5115] = '{3};
test_input[40928:40935] = '{32'hc1e782e6, 32'hc23562d8, 32'hc1eb700e, 32'hc2996cc4, 32'h420a01e3, 32'h4295fcd2, 32'hc26fad80, 32'hbeaa9dd0};
test_output[5116] = '{32'h4295fcd2};
test_index[5116] = '{5};
test_input[40936:40943] = '{32'hc29cc0ca, 32'hc1dcf5e0, 32'hc1cb8568, 32'h41d42ef4, 32'h427ed34a, 32'hc2c20120, 32'h42bfbe7d, 32'h419900e4};
test_output[5117] = '{32'h42bfbe7d};
test_index[5117] = '{6};
test_input[40944:40951] = '{32'h40a2213a, 32'hc24dca4c, 32'hc198f701, 32'h41e542b3, 32'h42524566, 32'h418c01e4, 32'hc23fef67, 32'hc2a89944};
test_output[5118] = '{32'h42524566};
test_index[5118] = '{4};
test_input[40952:40959] = '{32'hc2b834c5, 32'h422bcee0, 32'h42918d9e, 32'h4280cfc5, 32'h40bc1a37, 32'h424b5b39, 32'hc2578b52, 32'hc2a5741a};
test_output[5119] = '{32'h42918d9e};
test_index[5119] = '{2};
test_input[40960:40967] = '{32'h40e97f41, 32'hc256ec95, 32'hc1677581, 32'hc29bf6ce, 32'hc149eb1b, 32'hc28c1760, 32'h41a0ac06, 32'hc25858f8};
test_output[5120] = '{32'h41a0ac06};
test_index[5120] = '{6};
test_input[40968:40975] = '{32'hc2b2a00b, 32'hc27c85cb, 32'h40df1749, 32'hc294255b, 32'h4244fa5e, 32'hc1a3a3cd, 32'h401c4b67, 32'h42bf19be};
test_output[5121] = '{32'h42bf19be};
test_index[5121] = '{7};
test_input[40976:40983] = '{32'h4244845e, 32'h426c342f, 32'h416d496c, 32'hc206208f, 32'hc0e2a9a8, 32'hc1fb8fa7, 32'hc296561f, 32'h42091d8c};
test_output[5122] = '{32'h426c342f};
test_index[5122] = '{1};
test_input[40984:40991] = '{32'h41b246e0, 32'hc2ab54c1, 32'h41cfddc6, 32'h41b57e09, 32'hc202c53f, 32'h419a3f6a, 32'hc2bd31fa, 32'hc283d7ad};
test_output[5123] = '{32'h41cfddc6};
test_index[5123] = '{2};
test_input[40992:40999] = '{32'h427dc7c3, 32'hc215b7b8, 32'h4207ef06, 32'hc198e9e4, 32'hc1f66a81, 32'h425f4ce4, 32'h4237905e, 32'hc29f8ac2};
test_output[5124] = '{32'h427dc7c3};
test_index[5124] = '{0};
test_input[41000:41007] = '{32'h42a31f03, 32'h41b04a14, 32'hc245605f, 32'hc2c60e73, 32'h42b73521, 32'h428a5c70, 32'h41b02e21, 32'hc27e0b72};
test_output[5125] = '{32'h42b73521};
test_index[5125] = '{4};
test_input[41008:41015] = '{32'hc26c1351, 32'hc220737a, 32'hc2ac795f, 32'hc251ce0c, 32'h4219eb86, 32'h41d83827, 32'hc16b40b4, 32'h41b040a2};
test_output[5126] = '{32'h4219eb86};
test_index[5126] = '{4};
test_input[41016:41023] = '{32'h419495fb, 32'h42448374, 32'hc243fef4, 32'h3fedab54, 32'h407f9d95, 32'hc2b02e31, 32'h424d759e, 32'hc1d91264};
test_output[5127] = '{32'h424d759e};
test_index[5127] = '{6};
test_input[41024:41031] = '{32'hc22afbe7, 32'hc21c6868, 32'h42a59615, 32'h42a15b30, 32'hc2148bfe, 32'h42ae1123, 32'h41cbca6f, 32'h429a70da};
test_output[5128] = '{32'h42ae1123};
test_index[5128] = '{5};
test_input[41032:41039] = '{32'hc2b5a222, 32'hc29568e9, 32'hc107b6fe, 32'h42156621, 32'h41cee497, 32'hc15c5fb2, 32'hc1541f44, 32'hc27f5595};
test_output[5129] = '{32'h42156621};
test_index[5129] = '{3};
test_input[41040:41047] = '{32'h4263a158, 32'h427d9297, 32'hc28f69b7, 32'hc1a72a15, 32'h4019c2f1, 32'hc2800e1c, 32'h4210a072, 32'h40febd40};
test_output[5130] = '{32'h427d9297};
test_index[5130] = '{1};
test_input[41048:41055] = '{32'h41e517d9, 32'h42210262, 32'h42ab21bb, 32'hc209cb5e, 32'hc26d47ec, 32'hc2a66ea7, 32'h425598d3, 32'hc2a27430};
test_output[5131] = '{32'h42ab21bb};
test_index[5131] = '{2};
test_input[41056:41063] = '{32'hc18cb611, 32'hc18f7cdb, 32'hc2c400f0, 32'h427383f2, 32'hc290aebf, 32'h429a32ce, 32'h423d8d4d, 32'h4105af79};
test_output[5132] = '{32'h429a32ce};
test_index[5132] = '{5};
test_input[41064:41071] = '{32'h42851087, 32'hc291e6ac, 32'hc20d174c, 32'hc1e70f0a, 32'hc23df628, 32'h41311fdd, 32'h421a30ec, 32'hc29bbdf0};
test_output[5133] = '{32'h42851087};
test_index[5133] = '{0};
test_input[41072:41079] = '{32'h42b8a8bf, 32'hc1f1b807, 32'hc1992612, 32'h42b0bbf5, 32'h41d494fe, 32'hc1738b72, 32'h414d3993, 32'h42662faa};
test_output[5134] = '{32'h42b8a8bf};
test_index[5134] = '{0};
test_input[41080:41087] = '{32'h427080c1, 32'h42865510, 32'hc21d3367, 32'hbfba23b8, 32'h4094c174, 32'h4230b1b9, 32'hc28007b7, 32'hc2869084};
test_output[5135] = '{32'h42865510};
test_index[5135] = '{1};
test_input[41088:41095] = '{32'h425a4448, 32'hc29c8b4e, 32'h41b5dee0, 32'hc28b1e38, 32'hc022c257, 32'hc2ade6cf, 32'hc2c104a3, 32'h41b3a60e};
test_output[5136] = '{32'h425a4448};
test_index[5136] = '{0};
test_input[41096:41103] = '{32'hc27ae89f, 32'h429b963e, 32'h40e4f992, 32'h4137c41a, 32'h4293481c, 32'hc290aee6, 32'h42459561, 32'hc1c6b757};
test_output[5137] = '{32'h429b963e};
test_index[5137] = '{1};
test_input[41104:41111] = '{32'hc19f181d, 32'hc21ceee4, 32'h4258be07, 32'hc1b5d339, 32'hc08d59a9, 32'h425cd0ea, 32'hc226f3f1, 32'h413f8881};
test_output[5138] = '{32'h425cd0ea};
test_index[5138] = '{5};
test_input[41112:41119] = '{32'hc223d388, 32'hc1dac0e2, 32'h408051e1, 32'hc297a22a, 32'h42668cd1, 32'hc2b23d9f, 32'hc222e957, 32'h4272f7ee};
test_output[5139] = '{32'h4272f7ee};
test_index[5139] = '{7};
test_input[41120:41127] = '{32'hc18d982f, 32'hc0a45649, 32'hc292c429, 32'hbfe59542, 32'h415b1d28, 32'h41cff8ec, 32'hc28e96ee, 32'hc2a79f78};
test_output[5140] = '{32'h41cff8ec};
test_index[5140] = '{5};
test_input[41128:41135] = '{32'hc2bbff4e, 32'h42239612, 32'hc245051e, 32'hc26adfed, 32'hc1f65295, 32'h41bc6c5d, 32'h4109fc1e, 32'h407d8456};
test_output[5141] = '{32'h42239612};
test_index[5141] = '{1};
test_input[41136:41143] = '{32'h42bed269, 32'hc1bd1d56, 32'h4291ca14, 32'h4267c38f, 32'h42a92a06, 32'h42ad4fe5, 32'h4158b101, 32'h422f58d6};
test_output[5142] = '{32'h42bed269};
test_index[5142] = '{0};
test_input[41144:41151] = '{32'h42095292, 32'hc1d006c1, 32'hc2685cf4, 32'h426a45ac, 32'hc22bf1b0, 32'h426d83e1, 32'hc11a4b65, 32'h42076140};
test_output[5143] = '{32'h426d83e1};
test_index[5143] = '{5};
test_input[41152:41159] = '{32'hc217138b, 32'h42ac3a0a, 32'hc0170ec6, 32'hc272816d, 32'h418a96a4, 32'h4159c498, 32'hc2b0bec3, 32'h42aa53f1};
test_output[5144] = '{32'h42ac3a0a};
test_index[5144] = '{1};
test_input[41160:41167] = '{32'h42a509cd, 32'hc2a5885e, 32'h42179f6f, 32'h405006bb, 32'h4263618b, 32'h41aeba1f, 32'hc297f5d2, 32'h41bf5734};
test_output[5145] = '{32'h42a509cd};
test_index[5145] = '{0};
test_input[41168:41175] = '{32'hc23f650c, 32'hc2865822, 32'hc2a8d818, 32'h4161c66a, 32'h4281461e, 32'h423d0612, 32'hc29aecb6, 32'h42477faf};
test_output[5146] = '{32'h4281461e};
test_index[5146] = '{4};
test_input[41176:41183] = '{32'h428db910, 32'h426dd0a4, 32'h418e811e, 32'hc22154f9, 32'hc20da7bb, 32'h41f82f3d, 32'h428d3172, 32'h41f56eee};
test_output[5147] = '{32'h428db910};
test_index[5147] = '{0};
test_input[41184:41191] = '{32'h42bdd995, 32'h4296bccd, 32'h41949583, 32'h42bac7f6, 32'hc205a0d5, 32'hc1ceb9ba, 32'hc207405f, 32'hc25a4d70};
test_output[5148] = '{32'h42bdd995};
test_index[5148] = '{0};
test_input[41192:41199] = '{32'h41e6c5af, 32'hc2a1fadb, 32'h424a179c, 32'h4260eba6, 32'hc150d912, 32'hc0fb2f6d, 32'hbfe984b6, 32'hc2930fe8};
test_output[5149] = '{32'h4260eba6};
test_index[5149] = '{3};
test_input[41200:41207] = '{32'h42335828, 32'h4227fb9b, 32'h42511648, 32'hc2be940d, 32'h423a7853, 32'h41a22c13, 32'h412384bc, 32'hc2286fe9};
test_output[5150] = '{32'h42511648};
test_index[5150] = '{2};
test_input[41208:41215] = '{32'h42c41d08, 32'hc22f143f, 32'h423c59f3, 32'h418a9857, 32'h42b7edc4, 32'hc1edbf6b, 32'hc1a4e2f8, 32'h424f13ea};
test_output[5151] = '{32'h42c41d08};
test_index[5151] = '{0};
test_input[41216:41223] = '{32'hc0985c6a, 32'hc217c4db, 32'hc1c10588, 32'h41afb7ff, 32'h4272354f, 32'h42a8aa47, 32'hc22b905f, 32'hc23e01c9};
test_output[5152] = '{32'h42a8aa47};
test_index[5152] = '{5};
test_input[41224:41231] = '{32'h4211ef7b, 32'h422440c5, 32'hc2b9b4f2, 32'h426880cc, 32'hc292be50, 32'hc26f52b4, 32'hc2aec136, 32'h424602df};
test_output[5153] = '{32'h426880cc};
test_index[5153] = '{3};
test_input[41232:41239] = '{32'hc222fb58, 32'hc1b4e078, 32'hc01cea31, 32'h4099640f, 32'hc2ade27f, 32'h42b799d3, 32'h4275c024, 32'hc22e5814};
test_output[5154] = '{32'h42b799d3};
test_index[5154] = '{5};
test_input[41240:41247] = '{32'h420b101f, 32'hc161c77e, 32'h428b58cc, 32'hc20ca705, 32'hc1d66275, 32'h42bf6d2e, 32'hc2a36f5a, 32'h42a84996};
test_output[5155] = '{32'h42bf6d2e};
test_index[5155] = '{5};
test_input[41248:41255] = '{32'hc28c3a76, 32'hc2a5ce8b, 32'hc28a2472, 32'hc1029afc, 32'hc19da9d1, 32'hc25e7942, 32'h426e9e12, 32'h42c4c028};
test_output[5156] = '{32'h42c4c028};
test_index[5156] = '{7};
test_input[41256:41263] = '{32'hc1a05341, 32'hc2b758a9, 32'h4112b2f7, 32'hc21d6c45, 32'hc26eeefe, 32'h429e3ac7, 32'h4061d56e, 32'hc2221b87};
test_output[5157] = '{32'h429e3ac7};
test_index[5157] = '{5};
test_input[41264:41271] = '{32'hc1a67633, 32'hc295e146, 32'hc04edd9d, 32'hc2b2cbef, 32'hc13466fd, 32'h42549cdf, 32'hc26af5a5, 32'h41521f14};
test_output[5158] = '{32'h42549cdf};
test_index[5158] = '{5};
test_input[41272:41279] = '{32'h42985d6b, 32'h42bafb10, 32'hc2a26a60, 32'hc14b62f2, 32'h41b6ad40, 32'hc2be9b14, 32'hc2ab2b27, 32'hc289eb05};
test_output[5159] = '{32'h42bafb10};
test_index[5159] = '{1};
test_input[41280:41287] = '{32'hc27b0edb, 32'hc27ea104, 32'h423dce53, 32'hc22a9b74, 32'h4112db88, 32'hc225a613, 32'h4266dd1d, 32'h41457d52};
test_output[5160] = '{32'h4266dd1d};
test_index[5160] = '{6};
test_input[41288:41295] = '{32'h421d1746, 32'h423bdf21, 32'hc13dbac4, 32'hc2a33d5f, 32'hc19f5b38, 32'hc27dd9d1, 32'h4282e82a, 32'hc2067b8b};
test_output[5161] = '{32'h4282e82a};
test_index[5161] = '{6};
test_input[41296:41303] = '{32'hc282c9f1, 32'hc2bf50c7, 32'h411af022, 32'h41fabdc0, 32'hc278464a, 32'hc2ab1b97, 32'h42c19107, 32'h3f8f35e5};
test_output[5162] = '{32'h42c19107};
test_index[5162] = '{6};
test_input[41304:41311] = '{32'h428bdbbf, 32'h4162c01c, 32'h41588951, 32'hc284fe62, 32'h41460744, 32'h429d2a36, 32'hc0e199ac, 32'h4264c9de};
test_output[5163] = '{32'h429d2a36};
test_index[5163] = '{5};
test_input[41312:41319] = '{32'hc2370577, 32'hc21074b4, 32'hc2c05468, 32'hc21b27df, 32'h427b51e6, 32'hc02f530f, 32'hc27eb017, 32'h42b5f6f6};
test_output[5164] = '{32'h42b5f6f6};
test_index[5164] = '{7};
test_input[41320:41327] = '{32'hc225c898, 32'hc24859e6, 32'h421f6cff, 32'h426d3031, 32'hc24f6b3b, 32'hc182eb0f, 32'h4245ef99, 32'h42436d70};
test_output[5165] = '{32'h426d3031};
test_index[5165] = '{3};
test_input[41328:41335] = '{32'hc23acd89, 32'hc2ab898c, 32'h4218467d, 32'hc26841d7, 32'hc28af7f7, 32'h421ac7c9, 32'hc22736a0, 32'hbf66e2ad};
test_output[5166] = '{32'h421ac7c9};
test_index[5166] = '{5};
test_input[41336:41343] = '{32'hc2319141, 32'h42ae7c9d, 32'hc2a394a9, 32'h42af87ba, 32'hc214cb92, 32'hc182853b, 32'h41c8fdb9, 32'hc27650fe};
test_output[5167] = '{32'h42af87ba};
test_index[5167] = '{3};
test_input[41344:41351] = '{32'hc0b420b6, 32'hc2a35c02, 32'hc2c4c405, 32'h42be4825, 32'hc2b47b6a, 32'hc2a50735, 32'hc1a600ec, 32'h42c7f4a4};
test_output[5168] = '{32'h42c7f4a4};
test_index[5168] = '{7};
test_input[41352:41359] = '{32'h415a3ea9, 32'h42c30b37, 32'hc1a990e2, 32'hc23c47b0, 32'h41a4a82f, 32'hc2a39b7d, 32'hc177bb27, 32'hc1036f83};
test_output[5169] = '{32'h42c30b37};
test_index[5169] = '{1};
test_input[41360:41367] = '{32'h42b1d6e0, 32'hc2105ebb, 32'hc23d5c59, 32'h4232b29c, 32'h4187482c, 32'hc255536d, 32'h42b2254f, 32'hc23e4e55};
test_output[5170] = '{32'h42b2254f};
test_index[5170] = '{6};
test_input[41368:41375] = '{32'hc2c64aa4, 32'hc0abcf2d, 32'hc281e1da, 32'hc2228955, 32'h428709c0, 32'hc2c6a919, 32'hc1d441d4, 32'hc2ac9600};
test_output[5171] = '{32'h428709c0};
test_index[5171] = '{4};
test_input[41376:41383] = '{32'hc2484585, 32'hc2a9065a, 32'hc2187f80, 32'h41ab8436, 32'h42563bb6, 32'h424bbe80, 32'h41de0ebd, 32'h421365fb};
test_output[5172] = '{32'h42563bb6};
test_index[5172] = '{4};
test_input[41384:41391] = '{32'h3e8e2a6b, 32'h41d24167, 32'h41472908, 32'hc26fc6fe, 32'h4276c84b, 32'h42947259, 32'h41e449b2, 32'hc2c5c373};
test_output[5173] = '{32'h42947259};
test_index[5173] = '{5};
test_input[41392:41399] = '{32'h42b22c5d, 32'h420eee41, 32'h423a26f4, 32'h42c7244a, 32'h42654b74, 32'hc2c1954c, 32'hc23ea4ed, 32'hc26cd177};
test_output[5174] = '{32'h42c7244a};
test_index[5174] = '{3};
test_input[41400:41407] = '{32'h405d2bb9, 32'h4256fbd2, 32'h42c1a581, 32'h42299839, 32'hc2b525fb, 32'h42a98231, 32'h4286233b, 32'hc206566c};
test_output[5175] = '{32'h42c1a581};
test_index[5175] = '{2};
test_input[41408:41415] = '{32'hc18a3600, 32'hc0ab6138, 32'h4269728e, 32'h4212fa42, 32'h428af70f, 32'hc21b42f9, 32'hc2912e95, 32'hc23599b9};
test_output[5176] = '{32'h428af70f};
test_index[5176] = '{4};
test_input[41416:41423] = '{32'hc288f9a3, 32'hc19800d2, 32'h4231a808, 32'hc18ab243, 32'h4172408c, 32'hc289c372, 32'hc004d0f6, 32'h41260be3};
test_output[5177] = '{32'h4231a808};
test_index[5177] = '{2};
test_input[41424:41431] = '{32'hc2c6c50e, 32'h41e354fa, 32'h416a36d5, 32'h41f7c0d9, 32'hc27fcaea, 32'h429185c7, 32'hc0b4a7ed, 32'h41902ab3};
test_output[5178] = '{32'h429185c7};
test_index[5178] = '{5};
test_input[41432:41439] = '{32'hc29b6134, 32'hc238e3f7, 32'h42aa4cef, 32'h41a5cbd5, 32'hc2a0a038, 32'hc20aefc9, 32'h41192b3d, 32'hc288a49f};
test_output[5179] = '{32'h42aa4cef};
test_index[5179] = '{2};
test_input[41440:41447] = '{32'hc097fea9, 32'h41f6b7ae, 32'hc21f2cf2, 32'hc22e86e0, 32'hc1e351d6, 32'hc24f16bc, 32'hc2aadba0, 32'h42a84b39};
test_output[5180] = '{32'h42a84b39};
test_index[5180] = '{7};
test_input[41448:41455] = '{32'h42875edd, 32'h42a5ca91, 32'hc0274594, 32'hc29bae5e, 32'hc1ea082a, 32'hc20772c0, 32'h42bc7dcf, 32'hc2805be3};
test_output[5181] = '{32'h42bc7dcf};
test_index[5181] = '{6};
test_input[41456:41463] = '{32'h42bd9bb2, 32'h41635ca4, 32'hc18dbec0, 32'hbf9177db, 32'h421430a4, 32'h428f5393, 32'hc2838f15, 32'hc2b3db8d};
test_output[5182] = '{32'h42bd9bb2};
test_index[5182] = '{0};
test_input[41464:41471] = '{32'h425cbf88, 32'h427f4bca, 32'hc20af60d, 32'h42b9a50f, 32'hc1e78c05, 32'hc2bc6828, 32'hc23ef16d, 32'h424260be};
test_output[5183] = '{32'h42b9a50f};
test_index[5183] = '{3};
test_input[41472:41479] = '{32'h4286c770, 32'hc2632457, 32'hc29d1265, 32'h42860ba8, 32'h427da669, 32'h40a7aaab, 32'hc1de8242, 32'hc28efb7b};
test_output[5184] = '{32'h4286c770};
test_index[5184] = '{0};
test_input[41480:41487] = '{32'hc29bee18, 32'hc2786c8a, 32'hc2b7b6d6, 32'h423dd368, 32'hc250eb36, 32'hc12c2cc1, 32'hc281156d, 32'h4201a518};
test_output[5185] = '{32'h423dd368};
test_index[5185] = '{3};
test_input[41488:41495] = '{32'h42b5dfb0, 32'hc28ddd35, 32'h42287ad6, 32'h422a054f, 32'h41c17876, 32'hc2427e1b, 32'h422f6ce1, 32'hc2174eeb};
test_output[5186] = '{32'h42b5dfb0};
test_index[5186] = '{0};
test_input[41496:41503] = '{32'h4246639f, 32'hc229a94e, 32'h42925d11, 32'h414c203d, 32'h40fe29a5, 32'hc2c24825, 32'hc2970af8, 32'hc2988387};
test_output[5187] = '{32'h42925d11};
test_index[5187] = '{2};
test_input[41504:41511] = '{32'hc2570957, 32'hc1863ecd, 32'hc1d6b5f5, 32'h420b5a87, 32'hc2b7afa7, 32'hc107227b, 32'h426f1270, 32'h423163d6};
test_output[5188] = '{32'h426f1270};
test_index[5188] = '{6};
test_input[41512:41519] = '{32'h42c28fe2, 32'h421be187, 32'h41bfca19, 32'hc2a0ae13, 32'hc25e6109, 32'hc211d92d, 32'hc22fee43, 32'h42212f4f};
test_output[5189] = '{32'h42c28fe2};
test_index[5189] = '{0};
test_input[41520:41527] = '{32'hc2b50ebf, 32'h42532851, 32'hc2822153, 32'hc1b2748d, 32'h40bcf2b9, 32'h42bd5305, 32'hc27c5dd9, 32'h424a80b3};
test_output[5190] = '{32'h42bd5305};
test_index[5190] = '{5};
test_input[41528:41535] = '{32'hc271b81d, 32'hc205ca66, 32'hc2472433, 32'hc0a66bd1, 32'h427a12de, 32'h423fde73, 32'hc27d8953, 32'h41ae6514};
test_output[5191] = '{32'h427a12de};
test_index[5191] = '{4};
test_input[41536:41543] = '{32'h41854b35, 32'h421d280b, 32'h421c684c, 32'h428517d5, 32'hc2a68256, 32'hc231b715, 32'h423275e5, 32'hc25c9bac};
test_output[5192] = '{32'h428517d5};
test_index[5192] = '{3};
test_input[41544:41551] = '{32'hc1d65f95, 32'hc22cc36d, 32'hc2aa8fef, 32'hc1859fa2, 32'hc263a690, 32'h42b5c8ef, 32'h40c0eeb3, 32'hc23ae970};
test_output[5193] = '{32'h42b5c8ef};
test_index[5193] = '{5};
test_input[41552:41559] = '{32'hc2349e5a, 32'h42bdc71b, 32'h4246927f, 32'hc182ccfa, 32'h401a9bcf, 32'hc2856eba, 32'h4224af17, 32'h41bf2afd};
test_output[5194] = '{32'h42bdc71b};
test_index[5194] = '{1};
test_input[41560:41567] = '{32'h428d2ba6, 32'hc28a96e3, 32'h4281d7dd, 32'h415e9f2d, 32'h42395435, 32'hc265dffe, 32'hc241c69a, 32'h4084096b};
test_output[5195] = '{32'h428d2ba6};
test_index[5195] = '{0};
test_input[41568:41575] = '{32'h420cc4a5, 32'hc133eaeb, 32'hc23e0561, 32'hc2b535f2, 32'hc273e94e, 32'hc1a6bd3d, 32'hc2551fcb, 32'h42c63836};
test_output[5196] = '{32'h42c63836};
test_index[5196] = '{7};
test_input[41576:41583] = '{32'hc1b9512b, 32'h42b919ad, 32'hc280e837, 32'hc263179a, 32'hc2044f35, 32'hc1202c00, 32'hc22696c1, 32'h41e4f7e9};
test_output[5197] = '{32'h42b919ad};
test_index[5197] = '{1};
test_input[41584:41591] = '{32'h428498d2, 32'h41d587ee, 32'hc286ddff, 32'h4252935e, 32'hc2086d02, 32'h41096cd3, 32'h41a27e98, 32'hc2151661};
test_output[5198] = '{32'h428498d2};
test_index[5198] = '{0};
test_input[41592:41599] = '{32'h428c1bda, 32'h42132d28, 32'h41f28ece, 32'hc108c527, 32'h42b8a54d, 32'h424a273b, 32'h42c6118b, 32'h410557be};
test_output[5199] = '{32'h42c6118b};
test_index[5199] = '{6};
test_input[41600:41607] = '{32'hc2c161c8, 32'h429adc68, 32'h401d10bd, 32'hc2be088b, 32'hc292543c, 32'h3f8d8607, 32'h416e4f26, 32'hc1f28587};
test_output[5200] = '{32'h429adc68};
test_index[5200] = '{1};
test_input[41608:41615] = '{32'hc234ff97, 32'h42bdeb23, 32'h42944ab9, 32'hc1150542, 32'hc1f563f7, 32'hc04b2112, 32'h4232f92e, 32'h425d8997};
test_output[5201] = '{32'h42bdeb23};
test_index[5201] = '{1};
test_input[41616:41623] = '{32'hc2606d53, 32'h428ae3fa, 32'h424bc0c4, 32'hc2aefc3a, 32'hc1968547, 32'h40d500bd, 32'hc17a0ad4, 32'hc2a894e9};
test_output[5202] = '{32'h428ae3fa};
test_index[5202] = '{1};
test_input[41624:41631] = '{32'hbf729904, 32'h4244f00f, 32'h41e1a073, 32'h40bab8db, 32'h42a84dd5, 32'hc1e1c044, 32'hc23121a3, 32'h40b19b63};
test_output[5203] = '{32'h42a84dd5};
test_index[5203] = '{4};
test_input[41632:41639] = '{32'h428f55b1, 32'hc1574d77, 32'hc2a585fd, 32'h42c768f3, 32'h42071034, 32'hc0667d81, 32'hc27d15c4, 32'hc1c408bf};
test_output[5204] = '{32'h42c768f3};
test_index[5204] = '{3};
test_input[41640:41647] = '{32'hc2642ee8, 32'h42bde832, 32'hc2808782, 32'h42b18eea, 32'h42538104, 32'h4266dab2, 32'hc0950b54, 32'h40808f74};
test_output[5205] = '{32'h42bde832};
test_index[5205] = '{1};
test_input[41648:41655] = '{32'h42c3f263, 32'hc294e0c8, 32'h41758e94, 32'h4154a427, 32'hc2523c91, 32'hc2c0df45, 32'hc177f656, 32'hc2c5f24b};
test_output[5206] = '{32'h42c3f263};
test_index[5206] = '{0};
test_input[41656:41663] = '{32'h42488023, 32'hc14d31ad, 32'h3e997320, 32'hc14a1288, 32'h4223d349, 32'h428406a4, 32'hc198efe3, 32'h4188279e};
test_output[5207] = '{32'h428406a4};
test_index[5207] = '{5};
test_input[41664:41671] = '{32'hc28fdeee, 32'h4291dee5, 32'hc1b9a1d4, 32'hc281114a, 32'h424cc9e4, 32'h423b9774, 32'h426f37f8, 32'h4246a51a};
test_output[5208] = '{32'h4291dee5};
test_index[5208] = '{1};
test_input[41672:41679] = '{32'hc242ef76, 32'h426ec78d, 32'h42c78c59, 32'h424aab41, 32'hc2920306, 32'hc1767c4c, 32'h429f0d30, 32'hc22546b6};
test_output[5209] = '{32'h42c78c59};
test_index[5209] = '{2};
test_input[41680:41687] = '{32'h42496919, 32'hc2908f75, 32'hc024334f, 32'hc2893ad0, 32'hc23aab6d, 32'hc207312b, 32'h42598ebd, 32'h415a3672};
test_output[5210] = '{32'h42598ebd};
test_index[5210] = '{6};
test_input[41688:41695] = '{32'h41cafbdf, 32'hc265d0c4, 32'h42212ef6, 32'h420132f1, 32'hc1bba096, 32'h42884fb1, 32'hc26f14ca, 32'h42601cb9};
test_output[5211] = '{32'h42884fb1};
test_index[5211] = '{5};
test_input[41696:41703] = '{32'h42986b9f, 32'hc1962c10, 32'h42468401, 32'hc21a88d1, 32'hc1fb642b, 32'hc19994d5, 32'h40bfb744, 32'h4288f963};
test_output[5212] = '{32'h42986b9f};
test_index[5212] = '{0};
test_input[41704:41711] = '{32'hc2c3b902, 32'h42a4801a, 32'h41c172e4, 32'h42bb5330, 32'hc228fa13, 32'h4239c623, 32'hc27e223c, 32'h4276f5a9};
test_output[5213] = '{32'h42bb5330};
test_index[5213] = '{3};
test_input[41712:41719] = '{32'hc2a7c6e3, 32'h428ddc8c, 32'h42c73b77, 32'hc230b5cd, 32'hc1d52558, 32'h428c007d, 32'hc1d25763, 32'hc18ea69e};
test_output[5214] = '{32'h42c73b77};
test_index[5214] = '{2};
test_input[41720:41727] = '{32'hc177ddef, 32'h4266191a, 32'hc1dac1e2, 32'h42c49be1, 32'hc202e237, 32'hc1a95bf6, 32'h423c2fd3, 32'h42b1274b};
test_output[5215] = '{32'h42c49be1};
test_index[5215] = '{3};
test_input[41728:41735] = '{32'h419002ab, 32'hc2120602, 32'hc2b54136, 32'h41a76c51, 32'hc29e945b, 32'hc2ac1ef8, 32'h42275f79, 32'hc050ba5f};
test_output[5216] = '{32'h42275f79};
test_index[5216] = '{6};
test_input[41736:41743] = '{32'h429d8e5e, 32'h428f3930, 32'hc29f50d0, 32'h40f48586, 32'hc11877d5, 32'h42b4333c, 32'h41b2834c, 32'h42890962};
test_output[5217] = '{32'h42b4333c};
test_index[5217] = '{5};
test_input[41744:41751] = '{32'hc1f27621, 32'hc1c559f3, 32'hc2138bf8, 32'hc29de12f, 32'hc286a264, 32'h428a1947, 32'hc2c4bc06, 32'hc1d3328c};
test_output[5218] = '{32'h428a1947};
test_index[5218] = '{5};
test_input[41752:41759] = '{32'h42a62353, 32'hc274628c, 32'h4197eb43, 32'hc0b29150, 32'h4284e152, 32'h42a19a10, 32'hc2222ab9, 32'h42b318e0};
test_output[5219] = '{32'h42b318e0};
test_index[5219] = '{7};
test_input[41760:41767] = '{32'hc247d8f3, 32'h41399dfb, 32'hc2b0279e, 32'h40ecda60, 32'h4287137a, 32'hc0b566b2, 32'h42717c19, 32'h4264b3b5};
test_output[5220] = '{32'h4287137a};
test_index[5220] = '{4};
test_input[41768:41775] = '{32'h42b206d4, 32'hc2227aa5, 32'hc22fe512, 32'hc0421e23, 32'h42b9d19f, 32'h42b9a2f5, 32'h42c130a2, 32'hc1ab7fe1};
test_output[5221] = '{32'h42c130a2};
test_index[5221] = '{6};
test_input[41776:41783] = '{32'hc2959637, 32'h41e6bb5c, 32'h4090d253, 32'h42463c28, 32'h4149b8ec, 32'h419895aa, 32'h42b924b1, 32'hc1385f2e};
test_output[5222] = '{32'h42b924b1};
test_index[5222] = '{6};
test_input[41784:41791] = '{32'h42a58d71, 32'h4299936d, 32'h421806a3, 32'h42a4f361, 32'h3f7b60f8, 32'hc2a9296f, 32'hc23e92f1, 32'hc21773f5};
test_output[5223] = '{32'h42a58d71};
test_index[5223] = '{0};
test_input[41792:41799] = '{32'h403660b8, 32'h429c0809, 32'h42c6bfe6, 32'hc292c2af, 32'hc26d6639, 32'hc2bf15a6, 32'h42797f0d, 32'hc231df4c};
test_output[5224] = '{32'h42c6bfe6};
test_index[5224] = '{2};
test_input[41800:41807] = '{32'hc2b78b39, 32'h429153f1, 32'hc1b5cd6a, 32'h42b75c0c, 32'h42083c55, 32'h425ad1e4, 32'h42b2feb0, 32'h427a4f19};
test_output[5225] = '{32'h42b75c0c};
test_index[5225] = '{3};
test_input[41808:41815] = '{32'hc241c95c, 32'h42901514, 32'h419ddbb7, 32'hc2ba7c14, 32'hc2966a69, 32'h41de4b8f, 32'h42584ad9, 32'hc1918768};
test_output[5226] = '{32'h42901514};
test_index[5226] = '{1};
test_input[41816:41823] = '{32'h417bf97b, 32'h42a39514, 32'hc185e477, 32'h42822bd7, 32'hc247687f, 32'hc2877cfd, 32'hc2b1db5c, 32'h428c6e98};
test_output[5227] = '{32'h42a39514};
test_index[5227] = '{1};
test_input[41824:41831] = '{32'hc2a7c06d, 32'h42a29409, 32'hc292e55a, 32'h42c5fd98, 32'hc26c18f3, 32'h4245ed9c, 32'h428e8006, 32'h42318bbd};
test_output[5228] = '{32'h42c5fd98};
test_index[5228] = '{3};
test_input[41832:41839] = '{32'h41d2600c, 32'h417a189b, 32'hc199ad10, 32'h42b6131e, 32'hc235714a, 32'hc2b45d08, 32'h4224d1d6, 32'hc19c7893};
test_output[5229] = '{32'h42b6131e};
test_index[5229] = '{3};
test_input[41840:41847] = '{32'hc1dc1524, 32'h4105e767, 32'h421fd885, 32'hc1214f72, 32'hc19f5f31, 32'hc28de3b7, 32'h418f2d16, 32'h42ad7c86};
test_output[5230] = '{32'h42ad7c86};
test_index[5230] = '{7};
test_input[41848:41855] = '{32'h429554f8, 32'h41a7f29e, 32'hc203badf, 32'hc1a022d3, 32'h4235db9d, 32'hc1b7e700, 32'hc28f8187, 32'h42a1065f};
test_output[5231] = '{32'h42a1065f};
test_index[5231] = '{7};
test_input[41856:41863] = '{32'hc19a6bd6, 32'hc10318f8, 32'hc2c3513d, 32'h42aae2f3, 32'hc233eb31, 32'hc182fb31, 32'h429e6ce8, 32'h41b2722e};
test_output[5232] = '{32'h42aae2f3};
test_index[5232] = '{3};
test_input[41864:41871] = '{32'hc10453aa, 32'h4095bdfd, 32'hc1c30335, 32'hc298a657, 32'h42935fd2, 32'hc256283e, 32'hc297e05a, 32'hc15289ef};
test_output[5233] = '{32'h42935fd2};
test_index[5233] = '{4};
test_input[41872:41879] = '{32'hc2959526, 32'h42ad0505, 32'hc244f4ea, 32'hbde0ecd3, 32'hc2a39ec4, 32'hc25af1c4, 32'hc2bf0d62, 32'h40f4a835};
test_output[5234] = '{32'h42ad0505};
test_index[5234] = '{1};
test_input[41880:41887] = '{32'h42a4fc82, 32'h41241d57, 32'h425c44e1, 32'h41b00c82, 32'hc2997b8c, 32'hc2aba600, 32'hc2befb00, 32'h429193e7};
test_output[5235] = '{32'h42a4fc82};
test_index[5235] = '{0};
test_input[41888:41895] = '{32'h413aea5f, 32'h421653ff, 32'hc2b8cc37, 32'hc280a29f, 32'h42b3bd36, 32'hc17f7a94, 32'h42c4f55c, 32'hc211bf41};
test_output[5236] = '{32'h42c4f55c};
test_index[5236] = '{6};
test_input[41896:41903] = '{32'h42c7ccb1, 32'h4227f575, 32'hc26f80a8, 32'h40b17eec, 32'h4196454f, 32'hc2aca553, 32'h4279ed9b, 32'h423d9e48};
test_output[5237] = '{32'h42c7ccb1};
test_index[5237] = '{0};
test_input[41904:41911] = '{32'h42307468, 32'h4266de67, 32'hc2aad0b4, 32'hc20f2044, 32'hc2ac18cd, 32'h42a0f303, 32'h42a116d3, 32'h428175fb};
test_output[5238] = '{32'h42a116d3};
test_index[5238] = '{6};
test_input[41912:41919] = '{32'hc2c6c18b, 32'hc1334f5c, 32'h429b0620, 32'hc28ace28, 32'hc14cbdfe, 32'h4158d5af, 32'hc268a29e, 32'h42167c54};
test_output[5239] = '{32'h429b0620};
test_index[5239] = '{2};
test_input[41920:41927] = '{32'h426adb96, 32'h4252122e, 32'hc2256a72, 32'hc20b19be, 32'hc2a8cf7d, 32'hbfd9641e, 32'h41fb1e69, 32'hc1269f68};
test_output[5240] = '{32'h426adb96};
test_index[5240] = '{0};
test_input[41928:41935] = '{32'h42b809d3, 32'hc2a02f87, 32'hc1d1264d, 32'h423112d3, 32'h422d29c3, 32'hc1573662, 32'h42c62aee, 32'hc26ae70e};
test_output[5241] = '{32'h42c62aee};
test_index[5241] = '{6};
test_input[41936:41943] = '{32'hc294f0ed, 32'hc1d35f5d, 32'h42424806, 32'h42c5af11, 32'hc2ab66a2, 32'hc2967cbe, 32'h41a8af1e, 32'hc09f270a};
test_output[5242] = '{32'h42c5af11};
test_index[5242] = '{3};
test_input[41944:41951] = '{32'h428ffad7, 32'h4287a765, 32'h420233d9, 32'h42a98684, 32'h41ce7be4, 32'h42c55825, 32'hc19eb221, 32'h42651933};
test_output[5243] = '{32'h42c55825};
test_index[5243] = '{5};
test_input[41952:41959] = '{32'hc2ac9cee, 32'h40e578d2, 32'h41ae47c5, 32'h428ce6ea, 32'hc276fac4, 32'hc29cd6a0, 32'hc26e169c, 32'hc2971bc6};
test_output[5244] = '{32'h428ce6ea};
test_index[5244] = '{3};
test_input[41960:41967] = '{32'hc205d249, 32'hc178bb32, 32'hc128f222, 32'h41657f8f, 32'hc24a6c9f, 32'h42a6c738, 32'hc086d6c3, 32'hc116965b};
test_output[5245] = '{32'h42a6c738};
test_index[5245] = '{5};
test_input[41968:41975] = '{32'hbeec26ab, 32'h420361c2, 32'hc2a8b741, 32'h419c0e12, 32'hc2511ed8, 32'hc2bab488, 32'hc2c5e449, 32'h42c305ca};
test_output[5246] = '{32'h42c305ca};
test_index[5246] = '{7};
test_input[41976:41983] = '{32'hc2524270, 32'h4257c9aa, 32'h42537bd0, 32'hc1abbf3e, 32'h428bf5a6, 32'h427e4d29, 32'h42807162, 32'h423103f1};
test_output[5247] = '{32'h428bf5a6};
test_index[5247] = '{4};
test_input[41984:41991] = '{32'hc24e6331, 32'hc2accbb8, 32'hc2a9e2dc, 32'h42c4951b, 32'hc0bd26d0, 32'hbfcdbed9, 32'hc2652e54, 32'h40e7daf4};
test_output[5248] = '{32'h42c4951b};
test_index[5248] = '{3};
test_input[41992:41999] = '{32'hc18d11c5, 32'hc27f7c8c, 32'hc23f0743, 32'h42363a05, 32'hc29b4559, 32'hc2761ba8, 32'h42168b51, 32'hc2552d1b};
test_output[5249] = '{32'h42363a05};
test_index[5249] = '{3};
test_input[42000:42007] = '{32'h42b861b9, 32'hc286ec25, 32'h41c59bd0, 32'hc0da9e56, 32'hc2916d45, 32'h415a38ea, 32'hc2c081d1, 32'h4212d9bf};
test_output[5250] = '{32'h42b861b9};
test_index[5250] = '{0};
test_input[42008:42015] = '{32'hc18ef871, 32'hc210ae8e, 32'h422e1bb9, 32'h42bfef4e, 32'hc26a4ad5, 32'h42836e8f, 32'hc0d736a8, 32'hc291cc1c};
test_output[5251] = '{32'h42bfef4e};
test_index[5251] = '{3};
test_input[42016:42023] = '{32'hc128bdb2, 32'hc297e253, 32'hc10f9b00, 32'h429767ac, 32'hc208d262, 32'h41e04bb8, 32'h417ac1d5, 32'hc1cb2575};
test_output[5252] = '{32'h429767ac};
test_index[5252] = '{3};
test_input[42024:42031] = '{32'hc2c2cff3, 32'hc2aaf201, 32'hc20c36c4, 32'hc0344319, 32'hc199913d, 32'h3f1e914c, 32'hc1f69e20, 32'h40cbfae9};
test_output[5253] = '{32'h40cbfae9};
test_index[5253] = '{7};
test_input[42032:42039] = '{32'h423c53af, 32'h4090c937, 32'hc2a374fc, 32'h420560f4, 32'h4190a4b6, 32'hc2af740e, 32'h4281385e, 32'h41826fb6};
test_output[5254] = '{32'h4281385e};
test_index[5254] = '{6};
test_input[42040:42047] = '{32'h4275af78, 32'hc2c7287e, 32'h4292be9b, 32'hc29af123, 32'hc2855b65, 32'h4206cd87, 32'hc1e2d78a, 32'hc1c3a0b5};
test_output[5255] = '{32'h4292be9b};
test_index[5255] = '{2};
test_input[42048:42055] = '{32'h42b200cd, 32'h4281a498, 32'h42ad6ee8, 32'h424291d9, 32'h41e7df6e, 32'hc2a364ba, 32'hc1d231d3, 32'hc185896a};
test_output[5256] = '{32'h42b200cd};
test_index[5256] = '{0};
test_input[42056:42063] = '{32'hc2c7b8df, 32'h424ab963, 32'hc21dfd8b, 32'hc27d2f9f, 32'hc2a9ab76, 32'h42223e0b, 32'hc28d42ab, 32'hbd30f4f5};
test_output[5257] = '{32'h424ab963};
test_index[5257] = '{1};
test_input[42064:42071] = '{32'hc2a86337, 32'hc2aea90d, 32'h42944053, 32'h41800852, 32'h426dfa0a, 32'h41e6b49c, 32'hc1c83c82, 32'hc16b0f19};
test_output[5258] = '{32'h42944053};
test_index[5258] = '{2};
test_input[42072:42079] = '{32'h428631d9, 32'h4241d6f7, 32'h41c76d78, 32'h421ebbf2, 32'hc2847793, 32'hc2c15262, 32'h42bb7ede, 32'hc1179088};
test_output[5259] = '{32'h42bb7ede};
test_index[5259] = '{6};
test_input[42080:42087] = '{32'h42c22b67, 32'hc29a1112, 32'h423173d2, 32'h425e3b16, 32'hc0308719, 32'hc26fba71, 32'h42523892, 32'h424ebed1};
test_output[5260] = '{32'h42c22b67};
test_index[5260] = '{0};
test_input[42088:42095] = '{32'h423f8da7, 32'h411465a5, 32'h412b6f37, 32'h42c52c83, 32'h42954107, 32'h42459254, 32'h420a1f46, 32'hc2a75fbf};
test_output[5261] = '{32'h42c52c83};
test_index[5261] = '{3};
test_input[42096:42103] = '{32'hc2891ad3, 32'h418c8343, 32'hc2c45f1c, 32'h42541f22, 32'h42779fe0, 32'hc0e1da1b, 32'hc0795d8d, 32'h421f7aaa};
test_output[5262] = '{32'h42779fe0};
test_index[5262] = '{4};
test_input[42104:42111] = '{32'hc27f533a, 32'h4298ab5f, 32'hc20c1679, 32'h41d9bb1f, 32'h410afbc4, 32'hc20832a0, 32'hc2b351e5, 32'hc272849e};
test_output[5263] = '{32'h4298ab5f};
test_index[5263] = '{1};
test_input[42112:42119] = '{32'h4203d090, 32'hc210a787, 32'h4110d1a0, 32'h423e159b, 32'hc2047779, 32'hc23ba7b4, 32'h423f8582, 32'hc2821114};
test_output[5264] = '{32'h423f8582};
test_index[5264] = '{6};
test_input[42120:42127] = '{32'hc18ad0ee, 32'hc12465f5, 32'hc2322ef7, 32'hc2391b0e, 32'h4253f525, 32'hc29a0486, 32'hc2c297b9, 32'hc2bd0b11};
test_output[5265] = '{32'h4253f525};
test_index[5265] = '{4};
test_input[42128:42135] = '{32'hc222d3bc, 32'h423154e1, 32'hc2b0ca72, 32'h4236a90f, 32'h42aada6e, 32'hc2ab6ea7, 32'hc298cba9, 32'hc24a72a1};
test_output[5266] = '{32'h42aada6e};
test_index[5266] = '{4};
test_input[42136:42143] = '{32'h41133e68, 32'h424e8c78, 32'hc257d525, 32'hc230a18f, 32'hc2bd9ad2, 32'hc2bc4d0d, 32'hc2a73916, 32'h42b4e74e};
test_output[5267] = '{32'h42b4e74e};
test_index[5267] = '{7};
test_input[42144:42151] = '{32'hc2c2d0c3, 32'h42b56ff6, 32'hc1f83d08, 32'h4273254e, 32'hc2463f77, 32'hc2868287, 32'h424e88c5, 32'h42b60ee9};
test_output[5268] = '{32'h42b60ee9};
test_index[5268] = '{7};
test_input[42152:42159] = '{32'hc29f9c17, 32'h41574617, 32'h4052da78, 32'hc2bcdb47, 32'hc20868c2, 32'hc2151205, 32'h4226c6cc, 32'h427e7557};
test_output[5269] = '{32'h427e7557};
test_index[5269] = '{7};
test_input[42160:42167] = '{32'hc2b0fc58, 32'h3ef4cb18, 32'hc1fb9b5e, 32'h42a39459, 32'hc273e962, 32'h424b9b7c, 32'h42580af5, 32'h42306386};
test_output[5270] = '{32'h42a39459};
test_index[5270] = '{3};
test_input[42168:42175] = '{32'hc21bf6b4, 32'h4298f976, 32'h4299fd3e, 32'hc25ebf76, 32'hc153661a, 32'hbee1c9c3, 32'hc20e86ef, 32'hc054c75f};
test_output[5271] = '{32'h4299fd3e};
test_index[5271] = '{2};
test_input[42176:42183] = '{32'hc2638aaa, 32'h41b3a4f8, 32'h42b458b8, 32'h41def83c, 32'h3ff1bef9, 32'h42a3feab, 32'hc25594ff, 32'hc1df2e93};
test_output[5272] = '{32'h42b458b8};
test_index[5272] = '{2};
test_input[42184:42191] = '{32'hc1c6c815, 32'h420e0245, 32'h42717548, 32'h42240ca5, 32'hc292b4d7, 32'h4233d54f, 32'hc22f10cb, 32'hc2b40767};
test_output[5273] = '{32'h42717548};
test_index[5273] = '{2};
test_input[42192:42199] = '{32'hc285eacf, 32'hc2baf2ca, 32'hc1104e04, 32'h429fc814, 32'h41a48dc5, 32'hc1b1babd, 32'h42532259, 32'h42497d1b};
test_output[5274] = '{32'h429fc814};
test_index[5274] = '{3};
test_input[42200:42207] = '{32'h4290b32b, 32'h4266c2c9, 32'h42519801, 32'h42c5f93c, 32'hbe1a5a82, 32'hc18e420d, 32'hc1ed6360, 32'h4154beb0};
test_output[5275] = '{32'h42c5f93c};
test_index[5275] = '{3};
test_input[42208:42215] = '{32'hc1b25441, 32'hc298588b, 32'h419950ad, 32'h4235f3ac, 32'hc2ada14c, 32'h41e38d38, 32'hc159dde9, 32'hc2894d37};
test_output[5276] = '{32'h4235f3ac};
test_index[5276] = '{3};
test_input[42216:42223] = '{32'h418545b0, 32'h427513de, 32'hc2904352, 32'h42a492ce, 32'h4293a016, 32'hc2a97f02, 32'h417f618d, 32'hc1b0d971};
test_output[5277] = '{32'h42a492ce};
test_index[5277] = '{3};
test_input[42224:42231] = '{32'hc16da451, 32'hc212cfb9, 32'h424a9783, 32'h42aac97e, 32'hc11c4e8d, 32'h41d23442, 32'hc2ae683f, 32'h425c10ef};
test_output[5278] = '{32'h42aac97e};
test_index[5278] = '{3};
test_input[42232:42239] = '{32'hc22f4bb6, 32'h418cde82, 32'h4112fc1f, 32'hc09692fd, 32'hc25f25ba, 32'h424b9842, 32'h41ea780f, 32'hc289062f};
test_output[5279] = '{32'h424b9842};
test_index[5279] = '{5};
test_input[42240:42247] = '{32'h4092bf2a, 32'hc23db780, 32'hc289b9b6, 32'hc2880c5b, 32'hc286ebb1, 32'hc2c3f5b4, 32'h429afabd, 32'h41949d46};
test_output[5280] = '{32'h429afabd};
test_index[5280] = '{6};
test_input[42248:42255] = '{32'hc1ed69c3, 32'hc2c2ce22, 32'h41c30ee1, 32'h41ec340a, 32'hc28b8cd7, 32'h41d0cdb3, 32'hc20e4077, 32'h42bfbc4e};
test_output[5281] = '{32'h42bfbc4e};
test_index[5281] = '{7};
test_input[42256:42263] = '{32'hc104d657, 32'h414c078e, 32'hc1e39f00, 32'h41b3a9b8, 32'hc18ee4cf, 32'hc1ea35ff, 32'hc2684e1e, 32'h42b76472};
test_output[5282] = '{32'h42b76472};
test_index[5282] = '{7};
test_input[42264:42271] = '{32'hc2303886, 32'hbfc16373, 32'h42a3c9f6, 32'hc24c193f, 32'h42b9646e, 32'h42b7dc08, 32'h424ffae8, 32'h42a5576d};
test_output[5283] = '{32'h42b9646e};
test_index[5283] = '{4};
test_input[42272:42279] = '{32'hc198dc1f, 32'h41ad6624, 32'h426bffab, 32'hc2b8eb91, 32'hbe8aca62, 32'hc1161e7a, 32'hc282032a, 32'hc2bb8e23};
test_output[5284] = '{32'h426bffab};
test_index[5284] = '{2};
test_input[42280:42287] = '{32'hc287b451, 32'hc0accf33, 32'hc283eda0, 32'hc1ca5539, 32'h42368efa, 32'hc1ceda4f, 32'h426f66d0, 32'h423032b4};
test_output[5285] = '{32'h426f66d0};
test_index[5285] = '{6};
test_input[42288:42295] = '{32'hc22f49fd, 32'hc2b05f23, 32'hc15905bb, 32'h3e898107, 32'h42a621ff, 32'h41b0db38, 32'h42541c54, 32'hc24679c8};
test_output[5286] = '{32'h42a621ff};
test_index[5286] = '{4};
test_input[42296:42303] = '{32'h418a88bf, 32'h42b0ab5f, 32'h42025935, 32'h4280e4d5, 32'hc2aef621, 32'hc199af16, 32'h3fa3b9a0, 32'hc26bed34};
test_output[5287] = '{32'h42b0ab5f};
test_index[5287] = '{1};
test_input[42304:42311] = '{32'h418f5faf, 32'hc2398471, 32'hc28cbc33, 32'h418086f9, 32'h42bd1ab3, 32'hc0a13213, 32'hc101bfad, 32'hc2c19705};
test_output[5288] = '{32'h42bd1ab3};
test_index[5288] = '{4};
test_input[42312:42319] = '{32'h41c14d65, 32'h411940ce, 32'hc1ef0349, 32'h425a78a5, 32'hc093ae21, 32'h405df488, 32'hc10df0fd, 32'h42adcff2};
test_output[5289] = '{32'h42adcff2};
test_index[5289] = '{7};
test_input[42320:42327] = '{32'h42578dcd, 32'h423502ed, 32'hc240d59f, 32'hc18c4b1a, 32'hc0f079b2, 32'h42ba0906, 32'hc25ff241, 32'hc29abcae};
test_output[5290] = '{32'h42ba0906};
test_index[5290] = '{5};
test_input[42328:42335] = '{32'hc2c34401, 32'hc0f6efc6, 32'h4264abe3, 32'hc1aa706c, 32'h4275af2a, 32'h41e5aac9, 32'h42c366a1, 32'hc287c0af};
test_output[5291] = '{32'h42c366a1};
test_index[5291] = '{6};
test_input[42336:42343] = '{32'h42677bc6, 32'hc1b17fcd, 32'hc27fa694, 32'h4207faaa, 32'h42b6b80d, 32'hc29f3f6d, 32'hc22ed329, 32'hc2932ddc};
test_output[5292] = '{32'h42b6b80d};
test_index[5292] = '{4};
test_input[42344:42351] = '{32'hc20de5cf, 32'hc1d6a844, 32'hc2b90642, 32'h42848c55, 32'h429dd558, 32'h42bb9b07, 32'hc29cc71d, 32'hc2539024};
test_output[5293] = '{32'h42bb9b07};
test_index[5293] = '{5};
test_input[42352:42359] = '{32'h42b53036, 32'h42a6a00d, 32'hc2a43d4b, 32'h424d6de4, 32'h4099e77f, 32'h42b11001, 32'hc2ba497b, 32'h42bb9290};
test_output[5294] = '{32'h42bb9290};
test_index[5294] = '{7};
test_input[42360:42367] = '{32'h42bb3444, 32'hc2bf320a, 32'h419d01a1, 32'h419a8cc6, 32'hc23c7fc3, 32'h4199fbad, 32'hc1e8c6c2, 32'h42a4fac2};
test_output[5295] = '{32'h42bb3444};
test_index[5295] = '{0};
test_input[42368:42375] = '{32'hc1c8140d, 32'hc0f83b80, 32'h42b6a3c7, 32'h425ae327, 32'hc2a1b13c, 32'h42aa9230, 32'hc2c6e77c, 32'h422f6c3b};
test_output[5296] = '{32'h42b6a3c7};
test_index[5296] = '{2};
test_input[42376:42383] = '{32'hc287940b, 32'hc1f92311, 32'h420ab439, 32'h4247ec6f, 32'h4235dc18, 32'hc2c36669, 32'h4291bd84, 32'hc1871c63};
test_output[5297] = '{32'h4291bd84};
test_index[5297] = '{6};
test_input[42384:42391] = '{32'h4278ced9, 32'hc2a86a70, 32'hc2575eed, 32'hc2aa7db0, 32'hc2b6733d, 32'h429fdf58, 32'h41c9d042, 32'h40a2b995};
test_output[5298] = '{32'h429fdf58};
test_index[5298] = '{5};
test_input[42392:42399] = '{32'hc2bebe00, 32'hbfe3abd1, 32'hc2aea1ec, 32'h415c1143, 32'h41dccc9f, 32'hc164087e, 32'h42233928, 32'hc2a14614};
test_output[5299] = '{32'h42233928};
test_index[5299] = '{6};
test_input[42400:42407] = '{32'h42983d53, 32'h42bf81b1, 32'h42a5a62c, 32'hc2026774, 32'hc2c0e5c7, 32'hc21fbe1b, 32'h4236da44, 32'h42a4e1ca};
test_output[5300] = '{32'h42bf81b1};
test_index[5300] = '{1};
test_input[42408:42415] = '{32'hc15d43dd, 32'h4256e1b3, 32'h41aec407, 32'hc28e0b83, 32'h41a95d3f, 32'hc1fb1e9d, 32'hc2b5ef70, 32'h422856ca};
test_output[5301] = '{32'h4256e1b3};
test_index[5301] = '{1};
test_input[42416:42423] = '{32'h428f2284, 32'hc2c21d7a, 32'hc22bea89, 32'h4222b069, 32'hc18f3998, 32'hc15ee286, 32'h425b977a, 32'h42add0ec};
test_output[5302] = '{32'h42add0ec};
test_index[5302] = '{7};
test_input[42424:42431] = '{32'hc2aa28d0, 32'h42633204, 32'h41d56616, 32'hc0a21948, 32'h423aa0a8, 32'hc2be600c, 32'hc1805324, 32'h428f5eb5};
test_output[5303] = '{32'h428f5eb5};
test_index[5303] = '{7};
test_input[42432:42439] = '{32'hc2a000de, 32'hc00d8288, 32'hc2886284, 32'hc2c2bfb3, 32'h427bc496, 32'hc2bae673, 32'h428f0e2e, 32'hc1bf60e6};
test_output[5304] = '{32'h428f0e2e};
test_index[5304] = '{6};
test_input[42440:42447] = '{32'h4298711f, 32'hc2c65143, 32'h4258b615, 32'hc2669f66, 32'hc1eb3bf2, 32'hc2a7bffb, 32'hc1bcbfd1, 32'h42548e19};
test_output[5305] = '{32'h4298711f};
test_index[5305] = '{0};
test_input[42448:42455] = '{32'hc1f8f522, 32'h425f45dd, 32'h42946051, 32'hc2218c95, 32'h420ad27f, 32'h4103ba80, 32'h42945a6f, 32'h42995784};
test_output[5306] = '{32'h42995784};
test_index[5306] = '{7};
test_input[42456:42463] = '{32'h41dd1b6f, 32'hc19d5747, 32'h4026e881, 32'h400fe146, 32'hc23ab45c, 32'hc214551e, 32'hc1d21a61, 32'h42254461};
test_output[5307] = '{32'h42254461};
test_index[5307] = '{7};
test_input[42464:42471] = '{32'hc28c3a5e, 32'h42a1d859, 32'hc2b7ad96, 32'hc2966f9e, 32'h4244eb54, 32'h425f5777, 32'h41585793, 32'h42395802};
test_output[5308] = '{32'h42a1d859};
test_index[5308] = '{1};
test_input[42472:42479] = '{32'hc0fdbf42, 32'h41c3e70e, 32'hc117fab4, 32'h4202bc53, 32'h42c7266b, 32'hc2a7fd6c, 32'hc22464ff, 32'hc2a05daa};
test_output[5309] = '{32'h42c7266b};
test_index[5309] = '{4};
test_input[42480:42487] = '{32'hc11ab72c, 32'hc2839b6b, 32'h41e8c136, 32'h428d7322, 32'h4250a18a, 32'hc1d76245, 32'hc1adf927, 32'h428a0d30};
test_output[5310] = '{32'h428d7322};
test_index[5310] = '{3};
test_input[42488:42495] = '{32'h4141e0cf, 32'hc1cc7f1e, 32'hc18a3dd8, 32'hc2b82675, 32'hc21ca2c8, 32'hc1553962, 32'hc1b72b35, 32'hc2428e15};
test_output[5311] = '{32'h4141e0cf};
test_index[5311] = '{0};
test_input[42496:42503] = '{32'hc1887de0, 32'hbd250692, 32'hc1e5978c, 32'h42b9089a, 32'h429ef7e7, 32'h429ade0c, 32'h410a3336, 32'hc25060b8};
test_output[5312] = '{32'h42b9089a};
test_index[5312] = '{3};
test_input[42504:42511] = '{32'h4146ec67, 32'h41cf8344, 32'hc1c05ba4, 32'h421bdb84, 32'h429be885, 32'h4239d3c3, 32'hc207a8fa, 32'hc2304f12};
test_output[5313] = '{32'h429be885};
test_index[5313] = '{4};
test_input[42512:42519] = '{32'hc170df3e, 32'h418b3cfc, 32'h423ee15f, 32'h3e821302, 32'hc2bb76c1, 32'h412572f6, 32'h4259ede4, 32'hc2073e5f};
test_output[5314] = '{32'h4259ede4};
test_index[5314] = '{6};
test_input[42520:42527] = '{32'hc285433d, 32'h40f46d5e, 32'hc1af4fbe, 32'h41a233a9, 32'h40faf0b0, 32'hc16c0aab, 32'h41561fba, 32'hc283315a};
test_output[5315] = '{32'h41a233a9};
test_index[5315] = '{3};
test_input[42528:42535] = '{32'hc2acd0ce, 32'hc25d8103, 32'h4259ba8c, 32'h419afd72, 32'h41ae4eca, 32'h429841ab, 32'hc2c5ee04, 32'h415eb73b};
test_output[5316] = '{32'h429841ab};
test_index[5316] = '{5};
test_input[42536:42543] = '{32'hc1538c77, 32'hc2ad2b49, 32'h417759f0, 32'hc2a78042, 32'h42028aab, 32'h41b418bd, 32'h42644a49, 32'hc104637d};
test_output[5317] = '{32'h42644a49};
test_index[5317] = '{6};
test_input[42544:42551] = '{32'h4283061d, 32'hc29925ab, 32'hc21fe1f7, 32'h424d045f, 32'h3ede7c05, 32'hc0cb41fa, 32'hc0df9c22, 32'hc241dd2d};
test_output[5318] = '{32'h4283061d};
test_index[5318] = '{0};
test_input[42552:42559] = '{32'h42a35805, 32'hc2b36471, 32'hc253a534, 32'h418d2c82, 32'hc1ba8895, 32'hbfcbe12a, 32'h4287c909, 32'hc24c80e5};
test_output[5319] = '{32'h42a35805};
test_index[5319] = '{0};
test_input[42560:42567] = '{32'h424e8faf, 32'hc22413e9, 32'h426e0f19, 32'h41caa4b1, 32'hc21d65dd, 32'h423968cf, 32'h42084809, 32'h4219c762};
test_output[5320] = '{32'h426e0f19};
test_index[5320] = '{2};
test_input[42568:42575] = '{32'hc1b0392f, 32'hc295b930, 32'hc282a99f, 32'h42bf0306, 32'hc23e3732, 32'h418c6e7f, 32'hc2c7155d, 32'hc280ea8d};
test_output[5321] = '{32'h42bf0306};
test_index[5321] = '{3};
test_input[42576:42583] = '{32'h42910f79, 32'hc2444567, 32'h426c6b30, 32'hc21a56e1, 32'hc05ef945, 32'h3db45915, 32'hc2bea796, 32'h42886018};
test_output[5322] = '{32'h42910f79};
test_index[5322] = '{0};
test_input[42584:42591] = '{32'hc0e34c38, 32'h42613a4b, 32'hc290c35a, 32'hc2b6905f, 32'hc253ee1b, 32'hc28d7c22, 32'hc214218d, 32'hc2833873};
test_output[5323] = '{32'h42613a4b};
test_index[5323] = '{1};
test_input[42592:42599] = '{32'h4294efd5, 32'h40f3f1c1, 32'h429922b6, 32'h42103217, 32'h41e4de83, 32'h421e9fbd, 32'hbfc34151, 32'hc2c768ec};
test_output[5324] = '{32'h429922b6};
test_index[5324] = '{2};
test_input[42600:42607] = '{32'h42354443, 32'h42630e12, 32'hc29c1b20, 32'h42972cca, 32'h426d8256, 32'hc12f0ba1, 32'hc2c07710, 32'h42c547fc};
test_output[5325] = '{32'h42c547fc};
test_index[5325] = '{7};
test_input[42608:42615] = '{32'hc15441e3, 32'h417cfc80, 32'hc2038b8c, 32'h423030c0, 32'h42ab9797, 32'hc117be7c, 32'h4181f649, 32'hc16e9d61};
test_output[5326] = '{32'h42ab9797};
test_index[5326] = '{4};
test_input[42616:42623] = '{32'hc2933777, 32'hc2397c22, 32'h428d74f3, 32'hc1873d5f, 32'h4291569e, 32'hc2c04c52, 32'h4105c0bd, 32'hc2be9364};
test_output[5327] = '{32'h4291569e};
test_index[5327] = '{4};
test_input[42624:42631] = '{32'h3f9b7ab9, 32'hc187ab8c, 32'h41f700e1, 32'h421aef22, 32'hc2495aa5, 32'h42bbe667, 32'hc1264691, 32'h42b84e58};
test_output[5328] = '{32'h42bbe667};
test_index[5328] = '{5};
test_input[42632:42639] = '{32'hc1d6bd49, 32'hc26c9589, 32'h42860d2d, 32'h42be2f1c, 32'hc0caa144, 32'hc2469ab3, 32'h429effaa, 32'hc2b5be68};
test_output[5329] = '{32'h42be2f1c};
test_index[5329] = '{3};
test_input[42640:42647] = '{32'hc177f79f, 32'hc1ab8673, 32'hc1b91bc1, 32'hc236620d, 32'hc23be76b, 32'hc10e0913, 32'h42747fcd, 32'h41e081fe};
test_output[5330] = '{32'h42747fcd};
test_index[5330] = '{6};
test_input[42648:42655] = '{32'h41c2cac7, 32'hc2bc69b3, 32'hc29919d6, 32'h428223a2, 32'h4137a675, 32'h42b6a7bb, 32'hc20d204c, 32'hc2b5274b};
test_output[5331] = '{32'h42b6a7bb};
test_index[5331] = '{5};
test_input[42656:42663] = '{32'h42538108, 32'hc29c1a5e, 32'h422a1b53, 32'hc2b353db, 32'h415bb989, 32'h40496389, 32'h40ba3091, 32'h42155723};
test_output[5332] = '{32'h42538108};
test_index[5332] = '{0};
test_input[42664:42671] = '{32'h4235ad73, 32'hc1b7182a, 32'hc2b586b9, 32'hc2949e4d, 32'hc19f0c37, 32'hc24aabe1, 32'h42be24b4, 32'h4243713b};
test_output[5333] = '{32'h42be24b4};
test_index[5333] = '{6};
test_input[42672:42679] = '{32'hc2a3a3fd, 32'h42b40112, 32'h416b38be, 32'h42b32412, 32'h40e76f84, 32'hc28c6c4f, 32'h42588427, 32'h42b3692b};
test_output[5334] = '{32'h42b40112};
test_index[5334] = '{1};
test_input[42680:42687] = '{32'h425e3891, 32'hc24c6d6a, 32'hc2842b41, 32'h42302781, 32'hc2c211d4, 32'h410758a7, 32'hc2a99f12, 32'hc2b35ceb};
test_output[5335] = '{32'h425e3891};
test_index[5335] = '{0};
test_input[42688:42695] = '{32'hc24d8e0d, 32'hbfc40b57, 32'h42131f0e, 32'h42856b6d, 32'hc28f22ac, 32'hc0314289, 32'h42368484, 32'hc1b7013c};
test_output[5336] = '{32'h42856b6d};
test_index[5336] = '{3};
test_input[42696:42703] = '{32'h429f45b3, 32'hc1ed802f, 32'hc235da58, 32'hc21326f2, 32'hc29c48d4, 32'h3f3a9708, 32'h429a9a75, 32'h40922b09};
test_output[5337] = '{32'h429f45b3};
test_index[5337] = '{0};
test_input[42704:42711] = '{32'hc2b98653, 32'h4022beb9, 32'hc222921d, 32'h42b1a24f, 32'hc20cf25d, 32'h4296efcb, 32'h4238d50f, 32'h4284c44b};
test_output[5338] = '{32'h42b1a24f};
test_index[5338] = '{3};
test_input[42712:42719] = '{32'h4180b7d0, 32'hc17f4fce, 32'h42264ba7, 32'hc2b60392, 32'h425e6859, 32'hc25380db, 32'hc2a290bf, 32'h4264bcb5};
test_output[5339] = '{32'h4264bcb5};
test_index[5339] = '{7};
test_input[42720:42727] = '{32'h42760617, 32'h4215545c, 32'hc286afab, 32'h42bcef10, 32'hc222158f, 32'hc2b6103e, 32'h425cb2c6, 32'h427ff83d};
test_output[5340] = '{32'h42bcef10};
test_index[5340] = '{3};
test_input[42728:42735] = '{32'hc2111e88, 32'h42a9084c, 32'h4234ff8a, 32'h428da5fe, 32'hc1f44e90, 32'hc2a6df75, 32'hc2876eaa, 32'hc1c68ffb};
test_output[5341] = '{32'h42a9084c};
test_index[5341] = '{1};
test_input[42736:42743] = '{32'hc1a15f4d, 32'hc1cb95fe, 32'h4296d99c, 32'hc294f9a9, 32'h42c59a97, 32'hc1cf74ae, 32'hc24deec5, 32'h42c56d87};
test_output[5342] = '{32'h42c59a97};
test_index[5342] = '{4};
test_input[42744:42751] = '{32'hbf46f27e, 32'h42b8f34f, 32'h41bbb481, 32'hc2797a31, 32'hc2aede7e, 32'h42afb08e, 32'hc293cd36, 32'hbfc44979};
test_output[5343] = '{32'h42b8f34f};
test_index[5343] = '{1};
test_input[42752:42759] = '{32'hc100de35, 32'hc1cdaaef, 32'hc22eae30, 32'hc2974686, 32'h425bff52, 32'h4200e262, 32'hc201499a, 32'hc26f3050};
test_output[5344] = '{32'h425bff52};
test_index[5344] = '{4};
test_input[42760:42767] = '{32'h4247c3a8, 32'hc2791f9c, 32'hc273d296, 32'h422c4848, 32'hc2c4fbbb, 32'h42a52324, 32'hc29ae1a8, 32'hc252d2fb};
test_output[5345] = '{32'h42a52324};
test_index[5345] = '{5};
test_input[42768:42775] = '{32'hc28ea8b3, 32'h42ad3e7b, 32'hc237edf4, 32'h42a1d767, 32'h4219e35b, 32'h419ce48f, 32'hc260b8a8, 32'hc2488fd5};
test_output[5346] = '{32'h42ad3e7b};
test_index[5346] = '{1};
test_input[42776:42783] = '{32'h420a4887, 32'hc2a8e550, 32'h417520ef, 32'hbfc276ad, 32'hc2933626, 32'h42829011, 32'hc1ba1884, 32'h41fddb8c};
test_output[5347] = '{32'h42829011};
test_index[5347] = '{5};
test_input[42784:42791] = '{32'h426e97cc, 32'h42b295a0, 32'h422e6894, 32'hc29b2430, 32'hc2b4add4, 32'h42aff89e, 32'hc11158d8, 32'hc28d393a};
test_output[5348] = '{32'h42b295a0};
test_index[5348] = '{1};
test_input[42792:42799] = '{32'hc1b72a29, 32'h42457342, 32'h41926205, 32'hc1b0b7f5, 32'hc2be715b, 32'hc2331877, 32'hc1efc2cc, 32'h41a4fc7a};
test_output[5349] = '{32'h42457342};
test_index[5349] = '{1};
test_input[42800:42807] = '{32'hc22e7c1f, 32'h41e2dc11, 32'hc2b9b25b, 32'hc2985943, 32'h41154a12, 32'hc1d7c4da, 32'hc09a7c4f, 32'h428373a1};
test_output[5350] = '{32'h428373a1};
test_index[5350] = '{7};
test_input[42808:42815] = '{32'hc16c811c, 32'h42a89ef4, 32'h3f7714f5, 32'hc275deaf, 32'hc29bfbc9, 32'h42c6e8cc, 32'hc252268d, 32'h42bf83e9};
test_output[5351] = '{32'h42c6e8cc};
test_index[5351] = '{5};
test_input[42816:42823] = '{32'hc2b43520, 32'hc2298804, 32'h42b58726, 32'h41f7bb86, 32'hc26fab29, 32'hc2b89d38, 32'h424a3186, 32'hc1ada722};
test_output[5352] = '{32'h42b58726};
test_index[5352] = '{2};
test_input[42824:42831] = '{32'h421b2f5d, 32'h4289730d, 32'hc1ddac24, 32'hc08da63f, 32'h423cf73e, 32'h42a8e409, 32'h429fce54, 32'h4257cb07};
test_output[5353] = '{32'h42a8e409};
test_index[5353] = '{5};
test_input[42832:42839] = '{32'hbf88259f, 32'hc29387a0, 32'h420e26f4, 32'hc2a24129, 32'h4200bd31, 32'hc256665b, 32'h427853c8, 32'h401f23e5};
test_output[5354] = '{32'h427853c8};
test_index[5354] = '{6};
test_input[42840:42847] = '{32'hc2c5e171, 32'h41ef749d, 32'hc1a49780, 32'h429678ba, 32'h42549bad, 32'hc234a33d, 32'hc184abd8, 32'h42a492c0};
test_output[5355] = '{32'h42a492c0};
test_index[5355] = '{7};
test_input[42848:42855] = '{32'h42458d38, 32'h421f0fd7, 32'hc1c889fb, 32'h426ba68d, 32'h42c4d172, 32'hc23af06a, 32'hc20544af, 32'h42c46b5a};
test_output[5356] = '{32'h42c4d172};
test_index[5356] = '{4};
test_input[42856:42863] = '{32'hc2b75098, 32'hc2a185b4, 32'hc28c593e, 32'h41813f9e, 32'hc278b547, 32'hc1baeed9, 32'hc1dd80b1, 32'hc2847a93};
test_output[5357] = '{32'h41813f9e};
test_index[5357] = '{3};
test_input[42864:42871] = '{32'hc21c1b3a, 32'h41b1b7ce, 32'hc28862fe, 32'h41807583, 32'hc293408a, 32'h411f8e87, 32'hc2c7fa2f, 32'h428e423a};
test_output[5358] = '{32'h428e423a};
test_index[5358] = '{7};
test_input[42872:42879] = '{32'hc2543426, 32'hc228689c, 32'h41c032cc, 32'h41d940a0, 32'h42288f31, 32'hc18fa95f, 32'h413d3ec2, 32'h418faaec};
test_output[5359] = '{32'h42288f31};
test_index[5359] = '{4};
test_input[42880:42887] = '{32'h4219ecda, 32'hc20f8826, 32'h42b6f7e4, 32'hc28b5261, 32'h4250341f, 32'hc283ff91, 32'hc18df019, 32'h4242973b};
test_output[5360] = '{32'h42b6f7e4};
test_index[5360] = '{2};
test_input[42888:42895] = '{32'h422ff07f, 32'hc216f030, 32'h418efc6e, 32'h4221cdcd, 32'h421801b5, 32'h42c27916, 32'hc2890cd8, 32'h42bbc0d6};
test_output[5361] = '{32'h42c27916};
test_index[5361] = '{5};
test_input[42896:42903] = '{32'hc196ff2d, 32'hc232e36a, 32'h418d2d33, 32'hc2a3275c, 32'hc1827842, 32'hc28fb0b3, 32'h41dfcaeb, 32'h42a5ee00};
test_output[5362] = '{32'h42a5ee00};
test_index[5362] = '{7};
test_input[42904:42911] = '{32'h42b94715, 32'h42af5f9a, 32'h4225e0c7, 32'h42993723, 32'h429b47c6, 32'hc2b34603, 32'hc20418c8, 32'h42900cac};
test_output[5363] = '{32'h42b94715};
test_index[5363] = '{0};
test_input[42912:42919] = '{32'hc2a78df7, 32'hc1f414c1, 32'hc2a68ebb, 32'h4186f023, 32'hc202a181, 32'h41b6a115, 32'h421d1245, 32'h41bb70fe};
test_output[5364] = '{32'h421d1245};
test_index[5364] = '{6};
test_input[42920:42927] = '{32'h42c5a836, 32'hc21ea70a, 32'hc209ae4e, 32'h40367441, 32'h408f388e, 32'h429faa30, 32'hbfeaceb0, 32'hc24946bc};
test_output[5365] = '{32'h42c5a836};
test_index[5365] = '{0};
test_input[42928:42935] = '{32'h3f9b185c, 32'h428444ab, 32'hc1e6452f, 32'hc2ad59ac, 32'h428b2675, 32'h42663723, 32'hc1a22abb, 32'h42bdf153};
test_output[5366] = '{32'h42bdf153};
test_index[5366] = '{7};
test_input[42936:42943] = '{32'h42869093, 32'h428aec5c, 32'hc28e6f50, 32'hc29f3c64, 32'h3fc063b9, 32'hc22ac35e, 32'hc0cd7d89, 32'h4280ba31};
test_output[5367] = '{32'h428aec5c};
test_index[5367] = '{1};
test_input[42944:42951] = '{32'hc2330a9e, 32'h42be78e9, 32'h428af00b, 32'hc26f3908, 32'h410fa848, 32'hc1b8f0e4, 32'h41a6b000, 32'h40d84ae4};
test_output[5368] = '{32'h42be78e9};
test_index[5368] = '{1};
test_input[42952:42959] = '{32'hc1733157, 32'h42258949, 32'hc28e76a2, 32'hc13f8693, 32'h423e2317, 32'h4234ca0e, 32'h426f4b3b, 32'hc1fb9b19};
test_output[5369] = '{32'h426f4b3b};
test_index[5369] = '{6};
test_input[42960:42967] = '{32'hbf962495, 32'h41b87a1d, 32'h42124b95, 32'h408f155e, 32'hc2ad4d4b, 32'hc25c740c, 32'h428780b4, 32'h428b6f09};
test_output[5370] = '{32'h428b6f09};
test_index[5370] = '{7};
test_input[42968:42975] = '{32'hc0f41ece, 32'hbf7ce151, 32'hc294f919, 32'h41516922, 32'h420766c8, 32'h42508662, 32'hc1d92a06, 32'h41e690ee};
test_output[5371] = '{32'h42508662};
test_index[5371] = '{5};
test_input[42976:42983] = '{32'hc1633c54, 32'h4252a373, 32'h415b94c4, 32'h4133e945, 32'h425af785, 32'hc2b3c101, 32'hc1a4b610, 32'hc16d0443};
test_output[5372] = '{32'h425af785};
test_index[5372] = '{4};
test_input[42984:42991] = '{32'hc27cd759, 32'hc2aa4ab8, 32'hc289155e, 32'hc15278ca, 32'h4244dbdb, 32'hc1bd6560, 32'hc2bb46f9, 32'h42739f48};
test_output[5373] = '{32'h42739f48};
test_index[5373] = '{7};
test_input[42992:42999] = '{32'hc22dbff5, 32'h427a2798, 32'h4202e84a, 32'h41fb07f5, 32'hc245ec46, 32'hc08de969, 32'hc28c5a0c, 32'hc2aa6a83};
test_output[5374] = '{32'h427a2798};
test_index[5374] = '{1};
test_input[43000:43007] = '{32'hc29742a9, 32'h426cdda5, 32'h4264ee21, 32'hc288be05, 32'hc216d30f, 32'hc2883c02, 32'hc22ddb9c, 32'hc29d3f6d};
test_output[5375] = '{32'h426cdda5};
test_index[5375] = '{1};
test_input[43008:43015] = '{32'h41ba7270, 32'hc1c3dbaa, 32'hc24a621c, 32'h42916be2, 32'hc20c4b5f, 32'h42115ca9, 32'h40ccef1f, 32'h3feefe22};
test_output[5376] = '{32'h42916be2};
test_index[5376] = '{3};
test_input[43016:43023] = '{32'hc29ae66f, 32'h427c3d60, 32'h42642c61, 32'h419fd8eb, 32'h428023da, 32'h426f26b1, 32'hc2418360, 32'h421cca51};
test_output[5377] = '{32'h428023da};
test_index[5377] = '{4};
test_input[43024:43031] = '{32'h412b21f3, 32'h415e527c, 32'h4204ff11, 32'h418c6922, 32'h41d6da0f, 32'h421f73e1, 32'h41951f16, 32'hc25f456d};
test_output[5378] = '{32'h421f73e1};
test_index[5378] = '{5};
test_input[43032:43039] = '{32'hc228cc4f, 32'hc2095cbe, 32'hc2ae4680, 32'hc26ee05f, 32'hc29c3b66, 32'hc2b0b24c, 32'hc1f7d7b1, 32'hc0f0ce26};
test_output[5379] = '{32'hc0f0ce26};
test_index[5379] = '{7};
test_input[43040:43047] = '{32'h428b144e, 32'h422e22b3, 32'hc1ae615d, 32'hc207d5c2, 32'hc085fcbd, 32'h42901a88, 32'hc1c08ad5, 32'hc0361d0f};
test_output[5380] = '{32'h42901a88};
test_index[5380] = '{5};
test_input[43048:43055] = '{32'hc28b2d66, 32'h422370c2, 32'hc262c78a, 32'hc2a48bb2, 32'h41c0612c, 32'h41e75140, 32'hc2ac64db, 32'h42bdd7c5};
test_output[5381] = '{32'h42bdd7c5};
test_index[5381] = '{7};
test_input[43056:43063] = '{32'hc24123d3, 32'hc2b9ebe9, 32'h423b01b1, 32'h413aad6a, 32'h420df053, 32'hc299ec54, 32'hc2c65704, 32'hc1eba8e3};
test_output[5382] = '{32'h423b01b1};
test_index[5382] = '{2};
test_input[43064:43071] = '{32'hc22b5f3e, 32'h42b03ba9, 32'hc26748ac, 32'hc0eb72df, 32'h420b8e81, 32'h4205b8e7, 32'h41bfe1d6, 32'hc2af0de7};
test_output[5383] = '{32'h42b03ba9};
test_index[5383] = '{1};
test_input[43072:43079] = '{32'hc207a9a9, 32'hc2ace31e, 32'hc293d9b9, 32'hc28c1141, 32'hc2ae20d7, 32'hc251bc92, 32'h411d7c56, 32'hc2ab2ff4};
test_output[5384] = '{32'h411d7c56};
test_index[5384] = '{6};
test_input[43080:43087] = '{32'h411f9b96, 32'hc2975991, 32'hc2c49d87, 32'hc290d126, 32'h426126c2, 32'hbfffa3b9, 32'h41ea4672, 32'hc15be838};
test_output[5385] = '{32'h426126c2};
test_index[5385] = '{4};
test_input[43088:43095] = '{32'hc291078c, 32'h42811067, 32'h42821ffb, 32'h40da5d46, 32'hc19fb349, 32'hc27228af, 32'hc2a96cfe, 32'h420be8fb};
test_output[5386] = '{32'h42821ffb};
test_index[5386] = '{2};
test_input[43096:43103] = '{32'h4174fda4, 32'hc1b72b54, 32'hc185cf70, 32'h41f118d4, 32'hc2b6b67d, 32'h42a80d94, 32'h41b4f1f6, 32'h40a32139};
test_output[5387] = '{32'h42a80d94};
test_index[5387] = '{5};
test_input[43104:43111] = '{32'h42b48e1a, 32'hc1a55376, 32'hbf88c5f0, 32'hc29cbbd9, 32'hc28a90bd, 32'h41b1e9e9, 32'hc29659ba, 32'hc29e170c};
test_output[5388] = '{32'h42b48e1a};
test_index[5388] = '{0};
test_input[43112:43119] = '{32'hc1dab018, 32'h42c31041, 32'h4233c104, 32'hc28d3a48, 32'h4260d5fe, 32'hc226b3a5, 32'h42a3db86, 32'hc2264a34};
test_output[5389] = '{32'h42c31041};
test_index[5389] = '{1};
test_input[43120:43127] = '{32'h42ade85e, 32'h42b97d5e, 32'hc214b59f, 32'h42a7ef1a, 32'hc2ae1049, 32'hbfcec55d, 32'h424a6e70, 32'hc25874fb};
test_output[5390] = '{32'h42b97d5e};
test_index[5390] = '{1};
test_input[43128:43135] = '{32'hc2a9f39d, 32'h415d473f, 32'hc0def96c, 32'hc2b6ad17, 32'h41a79f4a, 32'hc201db29, 32'h42522f08, 32'hc1de7cf4};
test_output[5391] = '{32'h42522f08};
test_index[5391] = '{6};
test_input[43136:43143] = '{32'h42afe7ed, 32'h421de8a9, 32'h40c25245, 32'h410f175b, 32'h427bbff3, 32'h4212ba76, 32'h40aa7f1b, 32'hc2b4e826};
test_output[5392] = '{32'h42afe7ed};
test_index[5392] = '{0};
test_input[43144:43151] = '{32'hc25bf419, 32'h41e8c539, 32'hc1e6c91a, 32'hc1904a20, 32'hc2aa889f, 32'h420cc1f6, 32'hc2bfa0d9, 32'h41830db0};
test_output[5393] = '{32'h420cc1f6};
test_index[5393] = '{5};
test_input[43152:43159] = '{32'h42b3d4f5, 32'hc2865b55, 32'hc1aad82c, 32'h418b2411, 32'hc23e08f2, 32'h42a0193d, 32'h42a3114f, 32'hc1e36386};
test_output[5394] = '{32'h42b3d4f5};
test_index[5394] = '{0};
test_input[43160:43167] = '{32'h41df3e8e, 32'hc28762fb, 32'hc1fb7adf, 32'hbd309341, 32'hc08bf1f3, 32'h4230af3d, 32'hc20661ed, 32'hc2844fd5};
test_output[5395] = '{32'h4230af3d};
test_index[5395] = '{5};
test_input[43168:43175] = '{32'hc2aebcaf, 32'h42973de1, 32'h42bdfba1, 32'hc160c57c, 32'h42893377, 32'h41b2b4fa, 32'hc15dd4a7, 32'hc28200f8};
test_output[5396] = '{32'h42bdfba1};
test_index[5396] = '{2};
test_input[43176:43183] = '{32'hc215d04a, 32'h4227b8e3, 32'h420b9d7a, 32'h42b9389a, 32'hc206424b, 32'h40cb5744, 32'h42991802, 32'hc1a585b1};
test_output[5397] = '{32'h42b9389a};
test_index[5397] = '{3};
test_input[43184:43191] = '{32'hc2c0ec7b, 32'h40d05aae, 32'h41b69b90, 32'h414cc285, 32'hc2b1fefb, 32'h41b64cce, 32'hc24fe2c3, 32'h4229b2de};
test_output[5398] = '{32'h4229b2de};
test_index[5398] = '{7};
test_input[43192:43199] = '{32'h40df2690, 32'hc28c68b7, 32'hc2abbb79, 32'h41d9da4e, 32'h42628c9c, 32'hc0756f74, 32'h41df1fec, 32'h42c68f35};
test_output[5399] = '{32'h42c68f35};
test_index[5399] = '{7};
test_input[43200:43207] = '{32'h4250768c, 32'hc187c161, 32'hc29e4756, 32'hc264f71a, 32'h42573e03, 32'h427d0be7, 32'hbfed7d05, 32'hc2b486a4};
test_output[5400] = '{32'h427d0be7};
test_index[5400] = '{5};
test_input[43208:43215] = '{32'hc2be2e6e, 32'h42bb6eea, 32'h42a21986, 32'hc23ddbdf, 32'hc1452e4c, 32'h40c38423, 32'hc15fdae2, 32'hc0c9e834};
test_output[5401] = '{32'h42bb6eea};
test_index[5401] = '{1};
test_input[43216:43223] = '{32'h4247b84d, 32'hc27677df, 32'hc207904f, 32'h421f64b1, 32'hc106659a, 32'h40e9e6e3, 32'hc26cdce8, 32'h42028257};
test_output[5402] = '{32'h4247b84d};
test_index[5402] = '{0};
test_input[43224:43231] = '{32'hc24d9ba8, 32'h41e9e814, 32'hc1169310, 32'h42910b2e, 32'hc17c39ab, 32'h42c4511d, 32'h42c042bb, 32'h41f90b8f};
test_output[5403] = '{32'h42c4511d};
test_index[5403] = '{5};
test_input[43232:43239] = '{32'hc19137c9, 32'hc2132656, 32'h425bc451, 32'hc28370d2, 32'h420ca4da, 32'hc2481edd, 32'hc1cbbb19, 32'hc255bf61};
test_output[5404] = '{32'h425bc451};
test_index[5404] = '{2};
test_input[43240:43247] = '{32'h419ae8cc, 32'hc1a7d131, 32'h429acf90, 32'h425c537f, 32'hc26a2734, 32'h4284fd2b, 32'hc2c27432, 32'h42046353};
test_output[5405] = '{32'h429acf90};
test_index[5405] = '{2};
test_input[43248:43255] = '{32'h42439fa6, 32'h42aebce6, 32'h42068030, 32'h41f80f8b, 32'hc2bcbda0, 32'h414e74a3, 32'h41ad36b3, 32'hc2a7e1c9};
test_output[5406] = '{32'h42aebce6};
test_index[5406] = '{1};
test_input[43256:43263] = '{32'hc21e7445, 32'hc2bbbece, 32'hc23dd44c, 32'hc20a0012, 32'h4185ea2f, 32'h41cd0fda, 32'hc26cf75f, 32'h420c31d1};
test_output[5407] = '{32'h420c31d1};
test_index[5407] = '{7};
test_input[43264:43271] = '{32'h42a4d468, 32'h42a45286, 32'hc261cddb, 32'hc229e70c, 32'h42930629, 32'h426f740e, 32'h422401e3, 32'h4239a68b};
test_output[5408] = '{32'h42a4d468};
test_index[5408] = '{0};
test_input[43272:43279] = '{32'hc08d1ae1, 32'h4217784f, 32'hc1d40f62, 32'hc2a8449e, 32'h429dc57d, 32'h4294bed7, 32'hc2a56f43, 32'h423f074f};
test_output[5409] = '{32'h429dc57d};
test_index[5409] = '{4};
test_input[43280:43287] = '{32'hc2a972ed, 32'hc24dc28d, 32'hc2b25fa7, 32'hc29ca0be, 32'h41eeebd9, 32'hc1755bea, 32'hc2926bb6, 32'h42039571};
test_output[5410] = '{32'h42039571};
test_index[5410] = '{7};
test_input[43288:43295] = '{32'h41e18a1a, 32'hc2753ce0, 32'hc2a4f809, 32'h42982a54, 32'h410068ae, 32'hc2ab7065, 32'h3fbcf9cf, 32'h410bcdd7};
test_output[5411] = '{32'h42982a54};
test_index[5411] = '{3};
test_input[43296:43303] = '{32'h4237d280, 32'h41a88465, 32'hc2b2a2af, 32'hc28b8996, 32'h42aae35f, 32'h4281e33e, 32'h40ed1d87, 32'hc2065b24};
test_output[5412] = '{32'h42aae35f};
test_index[5412] = '{4};
test_input[43304:43311] = '{32'h42860bb2, 32'hc28d4ebd, 32'h4255c363, 32'hc29bcbe0, 32'hbf79e374, 32'hc28ee07b, 32'hc2624493, 32'hc2923375};
test_output[5413] = '{32'h42860bb2};
test_index[5413] = '{0};
test_input[43312:43319] = '{32'h4258bda1, 32'hc1c90db0, 32'h42a69ac2, 32'hc2b7eb3c, 32'hc217fc30, 32'hc173bb24, 32'hbeb68b75, 32'h41f650d8};
test_output[5414] = '{32'h42a69ac2};
test_index[5414] = '{2};
test_input[43320:43327] = '{32'hc2ac3c45, 32'hc238dd3f, 32'h41e87632, 32'hc2b3fed2, 32'h4125fcbd, 32'h420e9753, 32'hc2123bd4, 32'hc1ffe721};
test_output[5415] = '{32'h420e9753};
test_index[5415] = '{5};
test_input[43328:43335] = '{32'hc1acddd6, 32'hc25d7d27, 32'h42bae99c, 32'h4284a136, 32'h41277b2c, 32'hc2888bd0, 32'hc2173dd4, 32'hc248a8d6};
test_output[5416] = '{32'h42bae99c};
test_index[5416] = '{2};
test_input[43336:43343] = '{32'hc2813cca, 32'h42a4cbed, 32'h421cd005, 32'hc284eb7f, 32'hc2b533e5, 32'h420f6531, 32'h423a002d, 32'h412636b4};
test_output[5417] = '{32'h42a4cbed};
test_index[5417] = '{1};
test_input[43344:43351] = '{32'h422419c6, 32'h42b82217, 32'hc2657e1c, 32'h4208c94e, 32'hc2aaeeaa, 32'h425f3483, 32'hc270f561, 32'hc2a9f090};
test_output[5418] = '{32'h42b82217};
test_index[5418] = '{1};
test_input[43352:43359] = '{32'h423772dc, 32'h419e9930, 32'hc0cccbc0, 32'h42183288, 32'h42ab1f5b, 32'hc25b495c, 32'h42bfb137, 32'h4219dac2};
test_output[5419] = '{32'h42bfb137};
test_index[5419] = '{6};
test_input[43360:43367] = '{32'hc1d5fdcf, 32'h4259299f, 32'h42726c25, 32'hc20b4a7f, 32'hc25e5005, 32'h42bd7f99, 32'hc18c57fa, 32'h42c0325d};
test_output[5420] = '{32'h42c0325d};
test_index[5420] = '{7};
test_input[43368:43375] = '{32'hc289688e, 32'hc2be523d, 32'h412e2af2, 32'hc28f1b51, 32'h42235c4a, 32'h4135e0f4, 32'hc185e932, 32'h4136c3da};
test_output[5421] = '{32'h42235c4a};
test_index[5421] = '{4};
test_input[43376:43383] = '{32'h41ffd3c7, 32'hc2284783, 32'h41897f60, 32'h41e8b965, 32'hc2567774, 32'h4265f303, 32'hc28fc8fe, 32'hc2b1ccd9};
test_output[5422] = '{32'h4265f303};
test_index[5422] = '{5};
test_input[43384:43391] = '{32'h42b8a6e7, 32'hc267ab6e, 32'hc2a23dbb, 32'h42a42646, 32'h41809f88, 32'h42351b77, 32'h4245afa0, 32'hc2018e63};
test_output[5423] = '{32'h42b8a6e7};
test_index[5423] = '{0};
test_input[43392:43399] = '{32'h42692454, 32'hc0208ece, 32'h415f3c8a, 32'hc20c553d, 32'h428e505a, 32'h41fe43e7, 32'hc1d7bec6, 32'h41586915};
test_output[5424] = '{32'h428e505a};
test_index[5424] = '{4};
test_input[43400:43407] = '{32'hc280c6f4, 32'hc226a5e0, 32'h427607e7, 32'h41be3ace, 32'hc20f52d4, 32'hc1dac43d, 32'h420b3086, 32'hc2c02ede};
test_output[5425] = '{32'h427607e7};
test_index[5425] = '{2};
test_input[43408:43415] = '{32'hc1fd1497, 32'hc2a58833, 32'hc2bb2b70, 32'hc2be9205, 32'h40cf6cf6, 32'hc2617864, 32'hc2b39bd5, 32'h4179e96e};
test_output[5426] = '{32'h4179e96e};
test_index[5426] = '{7};
test_input[43416:43423] = '{32'h42568e0c, 32'hc2bf3321, 32'hc14f631c, 32'h42af531d, 32'hc24cbf05, 32'hc1863924, 32'h417cf4f1, 32'hc2b708e9};
test_output[5427] = '{32'h42af531d};
test_index[5427] = '{3};
test_input[43424:43431] = '{32'hc16a1456, 32'hc1aff688, 32'h41cc35e8, 32'hc122e18b, 32'h415746c4, 32'hc2a7ff19, 32'hc25b8121, 32'h420ebbc1};
test_output[5428] = '{32'h420ebbc1};
test_index[5428] = '{7};
test_input[43432:43439] = '{32'hc261c19f, 32'hc1af1f38, 32'h429c647c, 32'hc2c6ef8a, 32'h4293421e, 32'h420e2586, 32'hc259a213, 32'hc219b8ce};
test_output[5429] = '{32'h429c647c};
test_index[5429] = '{2};
test_input[43440:43447] = '{32'h41c38176, 32'h42be510b, 32'hc14f2e36, 32'hc028cd2f, 32'hc29d3a93, 32'h4241777b, 32'hc242a1f1, 32'h4237e003};
test_output[5430] = '{32'h42be510b};
test_index[5430] = '{1};
test_input[43448:43455] = '{32'h41b5fa3f, 32'h425b1463, 32'h420a9146, 32'hc2b37c0b, 32'h42b3d09d, 32'hc27b4fec, 32'h41aafc34, 32'hc2b79188};
test_output[5431] = '{32'h42b3d09d};
test_index[5431] = '{4};
test_input[43456:43463] = '{32'h4280ba98, 32'h41ab04f0, 32'h3fddda75, 32'h4212ba28, 32'hc29b9685, 32'hc28145b1, 32'hc18f8d09, 32'hc2a8a27c};
test_output[5432] = '{32'h4280ba98};
test_index[5432] = '{0};
test_input[43464:43471] = '{32'h42b5d39d, 32'hc2c7e8f6, 32'hc2830d75, 32'h40022c39, 32'hc0da4590, 32'h426ea797, 32'h429347e3, 32'hc2bf5eb5};
test_output[5433] = '{32'h42b5d39d};
test_index[5433] = '{0};
test_input[43472:43479] = '{32'h41d7ced9, 32'h429457b2, 32'h41916561, 32'h42aff42b, 32'h424a6119, 32'hc235cf6a, 32'hc2c151e9, 32'hc19ded99};
test_output[5434] = '{32'h42aff42b};
test_index[5434] = '{3};
test_input[43480:43487] = '{32'hc251d01f, 32'hc29881d2, 32'hc29a64c5, 32'h421b2cb1, 32'h41e52f95, 32'h4288272c, 32'h41cc3c8e, 32'hc1d7349f};
test_output[5435] = '{32'h4288272c};
test_index[5435] = '{5};
test_input[43488:43495] = '{32'hc1c8f8b4, 32'hc25ef67e, 32'hc26d69b0, 32'hc2098df9, 32'hc29eeac1, 32'h42a61207, 32'h4232f59b, 32'h429d00f8};
test_output[5436] = '{32'h42a61207};
test_index[5436] = '{5};
test_input[43496:43503] = '{32'h42a5b703, 32'hc2498405, 32'h429ac852, 32'hc2aaf96c, 32'hc165ff32, 32'hc2b87077, 32'h42ad6948, 32'h41e6cf71};
test_output[5437] = '{32'h42ad6948};
test_index[5437] = '{6};
test_input[43504:43511] = '{32'h42c06010, 32'hc26c8b50, 32'hc003f950, 32'h4230648b, 32'h42ad6772, 32'h4284f0b9, 32'hc26fb29f, 32'h406e30a2};
test_output[5438] = '{32'h42c06010};
test_index[5438] = '{0};
test_input[43512:43519] = '{32'hc200e492, 32'h4232cd60, 32'hbf91c3f4, 32'h427790a8, 32'hc2a79718, 32'h415475ec, 32'h42b9bd57, 32'hc208ad40};
test_output[5439] = '{32'h42b9bd57};
test_index[5439] = '{6};
test_input[43520:43527] = '{32'h41e2c579, 32'hbfd99276, 32'h4177c78c, 32'hc13a6b17, 32'h42bc869b, 32'h429e6e56, 32'hc298c4da, 32'h4150f4c8};
test_output[5440] = '{32'h42bc869b};
test_index[5440] = '{4};
test_input[43528:43535] = '{32'h428a1de8, 32'h42783d9d, 32'h41f50b57, 32'h42a54fb2, 32'h425faa45, 32'h426db781, 32'h419f9e54, 32'h42ac2640};
test_output[5441] = '{32'h42ac2640};
test_index[5441] = '{7};
test_input[43536:43543] = '{32'h4201351e, 32'h42b7c8e1, 32'h42bc13b9, 32'h4292bd48, 32'hc2ac3829, 32'hc2babdcd, 32'hc0409290, 32'hbff82e19};
test_output[5442] = '{32'h42bc13b9};
test_index[5442] = '{2};
test_input[43544:43551] = '{32'h420aafec, 32'hc2b04a89, 32'h4243e9ff, 32'hc2a4c0e8, 32'h4200004c, 32'h41ba6147, 32'h42bb5884, 32'hc2292239};
test_output[5443] = '{32'h42bb5884};
test_index[5443] = '{6};
test_input[43552:43559] = '{32'hc2b65dcc, 32'hc0643470, 32'hc129cd17, 32'hc1af2be3, 32'h428cc2ea, 32'hc2069c06, 32'hc0e4fcec, 32'h42925ba2};
test_output[5444] = '{32'h42925ba2};
test_index[5444] = '{7};
test_input[43560:43567] = '{32'hc1337315, 32'hc088f430, 32'hc28fcb35, 32'h42c74017, 32'hc23a511b, 32'hc27691b1, 32'hc19bd0d8, 32'h4299e1f5};
test_output[5445] = '{32'h42c74017};
test_index[5445] = '{3};
test_input[43568:43575] = '{32'hc233aa22, 32'hc29cd498, 32'hc29e4c94, 32'hc21b2842, 32'h422ad44a, 32'h4282adcf, 32'h4275c984, 32'hc2a6ec1e};
test_output[5446] = '{32'h4282adcf};
test_index[5446] = '{5};
test_input[43576:43583] = '{32'hc1d155d7, 32'hc24faf98, 32'hc221655d, 32'hc14d9bd5, 32'h42b7169c, 32'hc0cccdb0, 32'hc2c6b218, 32'hc2a77f12};
test_output[5447] = '{32'h42b7169c};
test_index[5447] = '{4};
test_input[43584:43591] = '{32'hc0043591, 32'hc2abd759, 32'h41cb13bd, 32'hc28e653d, 32'hc2a393ab, 32'hc27ba3ec, 32'h4228ec19, 32'h4276abc8};
test_output[5448] = '{32'h4276abc8};
test_index[5448] = '{7};
test_input[43592:43599] = '{32'hc26541d2, 32'hc2b96ab7, 32'h41dc222d, 32'hc129e4bf, 32'hc244ec37, 32'hc1c94201, 32'hc07f5bc0, 32'h41689059};
test_output[5449] = '{32'h41dc222d};
test_index[5449] = '{2};
test_input[43600:43607] = '{32'hc2c6a7e4, 32'hc27213a9, 32'hc2989cbe, 32'hc1ff9aa9, 32'h4297b2a8, 32'h41743f2b, 32'h428dc0b2, 32'hc272b817};
test_output[5450] = '{32'h4297b2a8};
test_index[5450] = '{4};
test_input[43608:43615] = '{32'h4225558e, 32'h4175f30b, 32'h416edf9d, 32'hc278dc9b, 32'hc2089404, 32'h42be0cbc, 32'hc1db6050, 32'h41451e60};
test_output[5451] = '{32'h42be0cbc};
test_index[5451] = '{5};
test_input[43616:43623] = '{32'hc2c62bd6, 32'h4279e415, 32'h41a350af, 32'h428ef71e, 32'h42a1c728, 32'h428f505d, 32'h423cba62, 32'h428f8425};
test_output[5452] = '{32'h42a1c728};
test_index[5452] = '{4};
test_input[43624:43631] = '{32'hc179f64c, 32'hc27088a5, 32'hc270800e, 32'hc13f9ddd, 32'h4211b2ae, 32'hc14ccb29, 32'h41b40b75, 32'hc299342b};
test_output[5453] = '{32'h4211b2ae};
test_index[5453] = '{4};
test_input[43632:43639] = '{32'h4205536b, 32'h42af3991, 32'h417ec8f4, 32'h428df246, 32'hc1ab7ab3, 32'hbffcdddd, 32'hc22d77b5, 32'h41f14980};
test_output[5454] = '{32'h42af3991};
test_index[5454] = '{1};
test_input[43640:43647] = '{32'h429bdaf1, 32'hc2ae06ae, 32'h426a26e6, 32'hc229fa64, 32'h428deec1, 32'hc285968e, 32'h4292095e, 32'h42bafee8};
test_output[5455] = '{32'h42bafee8};
test_index[5455] = '{7};
test_input[43648:43655] = '{32'h424bc8f5, 32'h41a71626, 32'h4226d1e4, 32'h429d45fb, 32'hc2bda1fc, 32'hc1e2a546, 32'h428f57a1, 32'h4239a513};
test_output[5456] = '{32'h429d45fb};
test_index[5456] = '{3};
test_input[43656:43663] = '{32'hc26b54cf, 32'hc2afc71f, 32'hc1adf289, 32'h421fc834, 32'h4119d3ba, 32'h4224c236, 32'h4245aad3, 32'h42bfc548};
test_output[5457] = '{32'h42bfc548};
test_index[5457] = '{7};
test_input[43664:43671] = '{32'hc1b27d74, 32'h40d7ff2b, 32'hc29a7df4, 32'hc18cf184, 32'hc2c0d60e, 32'hc29c4b1d, 32'hc21e81e2, 32'hc09c03f8};
test_output[5458] = '{32'h40d7ff2b};
test_index[5458] = '{1};
test_input[43672:43679] = '{32'hc24bb183, 32'hc2518bd7, 32'h4134c1a5, 32'h413cb46f, 32'hc25d3d4d, 32'h41dc8f18, 32'hc22ad1f9, 32'h4293aa4c};
test_output[5459] = '{32'h4293aa4c};
test_index[5459] = '{7};
test_input[43680:43687] = '{32'hc1f18760, 32'h42388e9e, 32'hc1d7792c, 32'hc27361a0, 32'hc2b74a43, 32'h409e5bb2, 32'hc226287f, 32'h418ecf83};
test_output[5460] = '{32'h42388e9e};
test_index[5460] = '{1};
test_input[43688:43695] = '{32'h42126527, 32'hc1178d53, 32'hc20194c7, 32'hc2082676, 32'h3f2bc855, 32'hbf835102, 32'hc2a207f6, 32'h42835170};
test_output[5461] = '{32'h42835170};
test_index[5461] = '{7};
test_input[43696:43703] = '{32'hc1a179ee, 32'h40bf586e, 32'h4274fca9, 32'hc2843a13, 32'hc2af90dc, 32'h428db912, 32'hc28d157f, 32'h429793fd};
test_output[5462] = '{32'h429793fd};
test_index[5462] = '{7};
test_input[43704:43711] = '{32'h425d4fc0, 32'hc2798d21, 32'hc025844e, 32'hc0b256d0, 32'hc2043a7c, 32'hc17b6675, 32'h42239f7f, 32'hc2b3134d};
test_output[5463] = '{32'h425d4fc0};
test_index[5463] = '{0};
test_input[43712:43719] = '{32'h42070233, 32'hc22d9d46, 32'h42a2657a, 32'h422e7644, 32'h41b69d22, 32'h428e7d65, 32'hbfbbab1c, 32'h42a77a85};
test_output[5464] = '{32'h42a77a85};
test_index[5464] = '{7};
test_input[43720:43727] = '{32'hc0c53b59, 32'hc221d784, 32'hc2b90edd, 32'h42c67b3f, 32'hc1ba81da, 32'hc217a5c3, 32'h4261e307, 32'hc2bc7e7a};
test_output[5465] = '{32'h42c67b3f};
test_index[5465] = '{3};
test_input[43728:43735] = '{32'hc2388fc9, 32'h426551b6, 32'h428dbad0, 32'hc1ea2244, 32'hc0f5de92, 32'hc2509c18, 32'h41a92b78, 32'hc20b0c0d};
test_output[5466] = '{32'h428dbad0};
test_index[5466] = '{2};
test_input[43736:43743] = '{32'h42bd33e9, 32'hc1860580, 32'h42a0d8f4, 32'hc2326657, 32'h417465f1, 32'hbfaf9522, 32'hc2a77f9d, 32'hc2aa9d9f};
test_output[5467] = '{32'h42bd33e9};
test_index[5467] = '{0};
test_input[43744:43751] = '{32'h4090c999, 32'hc286c39b, 32'h422970e0, 32'h40552469, 32'hc2662790, 32'hc2bcb651, 32'hc1edd2c7, 32'h429ee830};
test_output[5468] = '{32'h429ee830};
test_index[5468] = '{7};
test_input[43752:43759] = '{32'h424c1781, 32'h422a2620, 32'h42bee88c, 32'hc2330ca4, 32'hc0c81820, 32'h42a64ac4, 32'hc23d2d66, 32'hc20f42f6};
test_output[5469] = '{32'h42bee88c};
test_index[5469] = '{2};
test_input[43760:43767] = '{32'hc26f212a, 32'h4216a5e3, 32'h42947e22, 32'h42a2ac5c, 32'hc28ccda4, 32'h4212533b, 32'hc28beed6, 32'h42448528};
test_output[5470] = '{32'h42a2ac5c};
test_index[5470] = '{3};
test_input[43768:43775] = '{32'hc29df2b1, 32'h41c68ecf, 32'h427d981e, 32'h41bbddaf, 32'hc2a0665c, 32'h417583e4, 32'hc1f7360b, 32'hc1cfc2e2};
test_output[5471] = '{32'h427d981e};
test_index[5471] = '{2};
test_input[43776:43783] = '{32'h424a428b, 32'hc2b6c03f, 32'h42bea42e, 32'h42839ae4, 32'h4253565e, 32'hc2bb98e7, 32'h420625c4, 32'h429d01e8};
test_output[5472] = '{32'h42bea42e};
test_index[5472] = '{2};
test_input[43784:43791] = '{32'hc2bbc264, 32'h421e2156, 32'hc2a5399e, 32'h404cb497, 32'h4196b453, 32'h423d970f, 32'hc1e5d010, 32'h4181d283};
test_output[5473] = '{32'h423d970f};
test_index[5473] = '{5};
test_input[43792:43799] = '{32'hc16af57e, 32'h421bec91, 32'hc1122eee, 32'hc1c19661, 32'hc2859521, 32'hc2c5db92, 32'h42878276, 32'hc00ade84};
test_output[5474] = '{32'h42878276};
test_index[5474] = '{6};
test_input[43800:43807] = '{32'hc166c109, 32'hc2927034, 32'hc15a3c78, 32'h42b2a45a, 32'hc2bd8c77, 32'hc243dc7d, 32'h421676e5, 32'h41e9fa17};
test_output[5475] = '{32'h42b2a45a};
test_index[5475] = '{3};
test_input[43808:43815] = '{32'hc2a8123f, 32'hc244e20e, 32'h42aa4d01, 32'hc28e5ec5, 32'h428dbdeb, 32'h4285e1bb, 32'hc27913cc, 32'hc2761333};
test_output[5476] = '{32'h42aa4d01};
test_index[5476] = '{2};
test_input[43816:43823] = '{32'hc1c8906a, 32'h4290863c, 32'h42b266c9, 32'h429503cc, 32'h4212ff28, 32'hc272db8f, 32'h4176507b, 32'hc236e11a};
test_output[5477] = '{32'h42b266c9};
test_index[5477] = '{2};
test_input[43824:43831] = '{32'hc0bbd8c0, 32'hc0cf4d64, 32'hc1d6e5ce, 32'hc1c6bd68, 32'hc2853ac5, 32'hc23da1bb, 32'h4186ee12, 32'hc2b69646};
test_output[5478] = '{32'h4186ee12};
test_index[5478] = '{6};
test_input[43832:43839] = '{32'hc295508a, 32'hc2aa21a9, 32'h42b953b8, 32'h422014d7, 32'h42825884, 32'hc2c4799c, 32'h424bfa4d, 32'h42667d18};
test_output[5479] = '{32'h42b953b8};
test_index[5479] = '{2};
test_input[43840:43847] = '{32'hc2070be4, 32'hc2226fc4, 32'h4297cd7c, 32'hc2b68b0a, 32'h41a97149, 32'h416f7297, 32'h4199f5f8, 32'hc2b94770};
test_output[5480] = '{32'h4297cd7c};
test_index[5480] = '{2};
test_input[43848:43855] = '{32'hc23e4dde, 32'hc2626b71, 32'hc29556fe, 32'h4212af40, 32'hc12c7522, 32'hc2928021, 32'h4263c055, 32'hc2c09e1b};
test_output[5481] = '{32'h4263c055};
test_index[5481] = '{6};
test_input[43856:43863] = '{32'h41e6babc, 32'h4102749e, 32'h4225e721, 32'h42b1eea7, 32'h42c6143e, 32'h42503fb6, 32'hc2a96349, 32'h424617fa};
test_output[5482] = '{32'h42c6143e};
test_index[5482] = '{4};
test_input[43864:43871] = '{32'h40cedcee, 32'h415258d8, 32'h42c0a7b4, 32'hc2b5b7a2, 32'hc23d969f, 32'hc21f5c1b, 32'hc2af8665, 32'hc18fbe3b};
test_output[5483] = '{32'h42c0a7b4};
test_index[5483] = '{2};
test_input[43872:43879] = '{32'hc1901502, 32'h42017090, 32'hc2041ac8, 32'hc216a85f, 32'hc20c234a, 32'hc27f92ae, 32'h42a721d0, 32'hc1e9be84};
test_output[5484] = '{32'h42a721d0};
test_index[5484] = '{6};
test_input[43880:43887] = '{32'h4191a7d8, 32'h40ddd73d, 32'hc2776a5e, 32'h4117b8da, 32'h4238aaa8, 32'h41c12aa2, 32'hc08bfb50, 32'h4198f1de};
test_output[5485] = '{32'h4238aaa8};
test_index[5485] = '{4};
test_input[43888:43895] = '{32'hc10b05ce, 32'h41ed895a, 32'h417f503b, 32'hc1822e83, 32'h42a2c217, 32'h4192433f, 32'hc1d9e3da, 32'h423795f4};
test_output[5486] = '{32'h42a2c217};
test_index[5486] = '{4};
test_input[43896:43903] = '{32'hc281dd7a, 32'h40cb9a98, 32'hc248bcb3, 32'h4283c4de, 32'hc24b35e1, 32'h4245f6b7, 32'hc28e6f25, 32'hc2b4e308};
test_output[5487] = '{32'h4283c4de};
test_index[5487] = '{3};
test_input[43904:43911] = '{32'hc2a05619, 32'hc2266b43, 32'hc21bd89e, 32'h4084d2d9, 32'hc07a627d, 32'hc29dd40b, 32'h403d03e6, 32'hc289ed50};
test_output[5488] = '{32'h4084d2d9};
test_index[5488] = '{3};
test_input[43912:43919] = '{32'h42210849, 32'hc26c22b8, 32'hc29966f3, 32'hc268cf68, 32'hc1dc9393, 32'h42850514, 32'h41999e27, 32'hc18a8efb};
test_output[5489] = '{32'h42850514};
test_index[5489] = '{5};
test_input[43920:43927] = '{32'hc2c208e0, 32'h418c887c, 32'hc2b08304, 32'hc2abaede, 32'h420210e5, 32'hc1e63270, 32'h41e83076, 32'hc2b84dff};
test_output[5490] = '{32'h420210e5};
test_index[5490] = '{4};
test_input[43928:43935] = '{32'hc1f68e54, 32'hc2b653c3, 32'hc2913c36, 32'hc20595b1, 32'hc264ae0a, 32'h419352f2, 32'hc2566041, 32'h4201a4be};
test_output[5491] = '{32'h4201a4be};
test_index[5491] = '{7};
test_input[43936:43943] = '{32'h40e447b2, 32'hc1188cec, 32'h41163593, 32'h41c4abf4, 32'hc2a1e096, 32'hc261881e, 32'hc2aca12c, 32'hc283b723};
test_output[5492] = '{32'h41c4abf4};
test_index[5492] = '{3};
test_input[43944:43951] = '{32'hc193c597, 32'h422b1140, 32'h4277d961, 32'hc2222867, 32'hc2a27b76, 32'hc24e6355, 32'hc2a55115, 32'hc271cdc9};
test_output[5493] = '{32'h4277d961};
test_index[5493] = '{2};
test_input[43952:43959] = '{32'hc2048868, 32'hc269d838, 32'hc298862b, 32'hc28bb2e6, 32'h40cd2ed6, 32'h428ee878, 32'h4270d650, 32'h4223df05};
test_output[5494] = '{32'h428ee878};
test_index[5494] = '{5};
test_input[43960:43967] = '{32'hc27d0d41, 32'h425cea6e, 32'hc24b83c0, 32'h4233f28a, 32'hc27bb2f0, 32'hc0837402, 32'h423bc5ab, 32'hc1e3f968};
test_output[5495] = '{32'h425cea6e};
test_index[5495] = '{1};
test_input[43968:43975] = '{32'hc1a52f39, 32'hc20b7436, 32'h41aa9554, 32'hc2befb82, 32'hc22789de, 32'hc016147f, 32'hc23d4203, 32'hc2a2e277};
test_output[5496] = '{32'h41aa9554};
test_index[5496] = '{2};
test_input[43976:43983] = '{32'hc24ab1e9, 32'h420a0b62, 32'hc265f28c, 32'hc236e49d, 32'hc246a937, 32'h41593a19, 32'hc2bacd96, 32'h422013cc};
test_output[5497] = '{32'h422013cc};
test_index[5497] = '{7};
test_input[43984:43991] = '{32'h4298760d, 32'h425be96a, 32'hc2357f3a, 32'h4209e088, 32'hc231b2eb, 32'hbf9b416e, 32'hc2bed228, 32'hc288b08d};
test_output[5498] = '{32'h4298760d};
test_index[5498] = '{0};
test_input[43992:43999] = '{32'h41bd8f52, 32'hc138f2bf, 32'h41e77611, 32'h4286aa13, 32'hc248adcd, 32'hc2756d81, 32'h429f7d8c, 32'hc2a714d8};
test_output[5499] = '{32'h429f7d8c};
test_index[5499] = '{6};
test_input[44000:44007] = '{32'h4154fe38, 32'h42916ed9, 32'hc2c6359e, 32'hc115eb16, 32'hc2b43003, 32'hc2561ec0, 32'hc10b15a1, 32'hc26c76b4};
test_output[5500] = '{32'h42916ed9};
test_index[5500] = '{1};
test_input[44008:44015] = '{32'h42932f59, 32'hc2085be8, 32'hc27c75e6, 32'h42898894, 32'hc134b1bc, 32'h4296b13e, 32'hc106cbd9, 32'hc28dc850};
test_output[5501] = '{32'h4296b13e};
test_index[5501] = '{5};
test_input[44016:44023] = '{32'hc2415207, 32'hc284461e, 32'h42c7bebd, 32'hc1fd18ba, 32'h42573ad9, 32'h41c57396, 32'hc2090737, 32'hc1a27f7e};
test_output[5502] = '{32'h42c7bebd};
test_index[5502] = '{2};
test_input[44024:44031] = '{32'h4236ec72, 32'h421174c1, 32'hc2b19e26, 32'hc2b178aa, 32'hc1e853f3, 32'hc2950186, 32'hc23d18cc, 32'h4246a16c};
test_output[5503] = '{32'h4246a16c};
test_index[5503] = '{7};
test_input[44032:44039] = '{32'hc25786c0, 32'hc1abbdcc, 32'h425740d8, 32'h425d256b, 32'hc12699bc, 32'hc14a1efe, 32'hc15ff7f9, 32'h4194bc57};
test_output[5504] = '{32'h425d256b};
test_index[5504] = '{3};
test_input[44040:44047] = '{32'hc1c8c85c, 32'hc132c902, 32'hc2c61616, 32'hc1a94880, 32'hc09c08f9, 32'hc2b70e69, 32'h42bd41f1, 32'hc208ef24};
test_output[5505] = '{32'h42bd41f1};
test_index[5505] = '{6};
test_input[44048:44055] = '{32'h42003f42, 32'h4298bccc, 32'h42a5c5b9, 32'hc17de458, 32'h428b7542, 32'hc2528a4c, 32'hc2000be9, 32'h42c352da};
test_output[5506] = '{32'h42c352da};
test_index[5506] = '{7};
test_input[44056:44063] = '{32'hc23cfaa2, 32'hc2911d23, 32'hc01458e8, 32'h4209eff9, 32'h4205ccc9, 32'hc2b5edaa, 32'hc295d8fa, 32'h420aa0ed};
test_output[5507] = '{32'h420aa0ed};
test_index[5507] = '{7};
test_input[44064:44071] = '{32'h41609e72, 32'hc153ca4d, 32'h42432124, 32'h40b5ceba, 32'hc27588fc, 32'h429f3736, 32'h4291a865, 32'hc2b44d47};
test_output[5508] = '{32'h429f3736};
test_index[5508] = '{5};
test_input[44072:44079] = '{32'h420a1e7f, 32'h3fa35944, 32'hc1185243, 32'h42760872, 32'hc20100e4, 32'hc1e22552, 32'h42a29f18, 32'hc0f75767};
test_output[5509] = '{32'h42a29f18};
test_index[5509] = '{6};
test_input[44080:44087] = '{32'h41f6cdc7, 32'h426b4dab, 32'hc29d5189, 32'h42901ee0, 32'hc29cecef, 32'h420a2e94, 32'h4285d3da, 32'hc21336bc};
test_output[5510] = '{32'h42901ee0};
test_index[5510] = '{3};
test_input[44088:44095] = '{32'h41e3a6d0, 32'hc2be2f22, 32'hc24bcd94, 32'h421f845f, 32'h4259d9c8, 32'h422662d8, 32'h40d96821, 32'hc1a595c0};
test_output[5511] = '{32'h4259d9c8};
test_index[5511] = '{4};
test_input[44096:44103] = '{32'h41e7a459, 32'hc1f6aff5, 32'hc1477816, 32'h41c6f735, 32'hc23d28cc, 32'hc2418a5f, 32'h42427f50, 32'hc29f1cd3};
test_output[5512] = '{32'h42427f50};
test_index[5512] = '{6};
test_input[44104:44111] = '{32'h429a2907, 32'hc2c1db94, 32'hc1c38f17, 32'h4085bf4c, 32'hc1538243, 32'h42ab45b3, 32'hc1f83c7e, 32'h41d32917};
test_output[5513] = '{32'h42ab45b3};
test_index[5513] = '{5};
test_input[44112:44119] = '{32'h42b8a9b7, 32'hc2c630a1, 32'h41ccc1fd, 32'hc24ec30f, 32'h42b3068e, 32'h4295143c, 32'hc268b55a, 32'h42aae3a0};
test_output[5514] = '{32'h42b8a9b7};
test_index[5514] = '{0};
test_input[44120:44127] = '{32'hc025b161, 32'hc283d766, 32'h41845a87, 32'h42c68e54, 32'hc1e0ae32, 32'h4299ba67, 32'h429fcb45, 32'hc1c11ce7};
test_output[5515] = '{32'h42c68e54};
test_index[5515] = '{3};
test_input[44128:44135] = '{32'hc29c00ef, 32'hc1156f3e, 32'h42b1b21d, 32'h428b9720, 32'hc280b723, 32'hc21b3b37, 32'hc0a20daf, 32'hc0b570ee};
test_output[5516] = '{32'h42b1b21d};
test_index[5516] = '{2};
test_input[44136:44143] = '{32'hc2bfd570, 32'hc2ac4b47, 32'hc2c2027a, 32'h42bf8da9, 32'h42a3ab95, 32'h41862fff, 32'h41028827, 32'h41f83d7b};
test_output[5517] = '{32'h42bf8da9};
test_index[5517] = '{3};
test_input[44144:44151] = '{32'hc23b82f6, 32'hc1e6bec8, 32'h423f1487, 32'hc22f368c, 32'hc118daed, 32'hc2b75c9b, 32'h4239a1f2, 32'h4147b36b};
test_output[5518] = '{32'h423f1487};
test_index[5518] = '{2};
test_input[44152:44159] = '{32'hc2a9f672, 32'h427a4962, 32'hc276d90e, 32'h42a7dada, 32'h421f955d, 32'h42b5241b, 32'hc1a8fc90, 32'hc2aa9d5c};
test_output[5519] = '{32'h42b5241b};
test_index[5519] = '{5};
test_input[44160:44167] = '{32'h424c6c9d, 32'h42bb2909, 32'hc0504216, 32'hc2c3f91a, 32'hc29fcae2, 32'hc2a53a90, 32'hc1a04926, 32'h41bdc6cd};
test_output[5520] = '{32'h42bb2909};
test_index[5520] = '{1};
test_input[44168:44175] = '{32'hc241c98a, 32'hc2bee6b0, 32'h42bd61b6, 32'h41ad7b70, 32'h419fae4e, 32'hc188eb74, 32'h421313c9, 32'hc2852fd0};
test_output[5521] = '{32'h42bd61b6};
test_index[5521] = '{2};
test_input[44176:44183] = '{32'h41ba2e49, 32'hc1e6c44a, 32'h4221672b, 32'hc2a2839e, 32'hc0d0ecde, 32'hc1ee65e9, 32'hc1cd6d5d, 32'hc287252a};
test_output[5522] = '{32'h4221672b};
test_index[5522] = '{2};
test_input[44184:44191] = '{32'h4285589e, 32'hc1b7f65f, 32'hc0f57831, 32'h4299e266, 32'h429a5ea5, 32'h424b3913, 32'h41ceaf1d, 32'h426788ec};
test_output[5523] = '{32'h429a5ea5};
test_index[5523] = '{4};
test_input[44192:44199] = '{32'h42abfbf1, 32'hc22a5693, 32'h4233794a, 32'hc277f874, 32'hc2bedb86, 32'hc28ff74d, 32'h42a368ea, 32'h3d8f02d0};
test_output[5524] = '{32'h42abfbf1};
test_index[5524] = '{0};
test_input[44200:44207] = '{32'h424bc974, 32'hc1a40124, 32'h42474a2e, 32'h420bcc62, 32'hc28e2ded, 32'h415e9a84, 32'h428a7ce3, 32'hc1907243};
test_output[5525] = '{32'h428a7ce3};
test_index[5525] = '{6};
test_input[44208:44215] = '{32'h42a1f781, 32'hc0e7c01d, 32'hc1ddec40, 32'hc2c0d30c, 32'hc1110c94, 32'h4267c610, 32'hc1c62820, 32'h4243bfd9};
test_output[5526] = '{32'h42a1f781};
test_index[5526] = '{0};
test_input[44216:44223] = '{32'hc1b0579b, 32'hc2523355, 32'h41909c76, 32'h42c6c662, 32'hc27504ec, 32'h42711a00, 32'h41b2a9bc, 32'hc2b9457e};
test_output[5527] = '{32'h42c6c662};
test_index[5527] = '{3};
test_input[44224:44231] = '{32'hc23dc53b, 32'hc1b1b262, 32'h42552f4c, 32'hc1342aa7, 32'hc2587e6a, 32'hc295c0d8, 32'h420820d3, 32'h41967809};
test_output[5528] = '{32'h42552f4c};
test_index[5528] = '{2};
test_input[44232:44239] = '{32'hc2b4b918, 32'hc26d2e8d, 32'h42bdc755, 32'hc28eefc6, 32'hc2229335, 32'hc2a2d553, 32'hc2bee21d, 32'hc1b8d355};
test_output[5529] = '{32'h42bdc755};
test_index[5529] = '{2};
test_input[44240:44247] = '{32'hc07e476c, 32'hc0007f16, 32'h42933a97, 32'hc2a93bca, 32'h42c39f8d, 32'h42a0d9c3, 32'h421fd051, 32'h42a2e349};
test_output[5530] = '{32'h42c39f8d};
test_index[5530] = '{4};
test_input[44248:44255] = '{32'hc276abaa, 32'h42a0b515, 32'hc262f446, 32'h42b90857, 32'h4288fd15, 32'h41532ed2, 32'hc2592293, 32'hc285b54a};
test_output[5531] = '{32'h42b90857};
test_index[5531] = '{3};
test_input[44256:44263] = '{32'hc2b5d5c9, 32'hc24dc74e, 32'h420020e9, 32'hc2280b3e, 32'h42c60ef7, 32'h429e7724, 32'hc2aa205a, 32'h41afcc04};
test_output[5532] = '{32'h42c60ef7};
test_index[5532] = '{4};
test_input[44264:44271] = '{32'h41cb4dfd, 32'hc2c3d03f, 32'hc24fde97, 32'h41d7dee2, 32'h42bffab3, 32'h42851b64, 32'h42489d4a, 32'hc1e0ef77};
test_output[5533] = '{32'h42bffab3};
test_index[5533] = '{4};
test_input[44272:44279] = '{32'h4209b55f, 32'h421778bd, 32'h41fa46f7, 32'h40edb76c, 32'h417dbb0c, 32'h4258f3c4, 32'hc28a8098, 32'h420fb74d};
test_output[5534] = '{32'h4258f3c4};
test_index[5534] = '{5};
test_input[44280:44287] = '{32'hc1b5591a, 32'hc224ced1, 32'h419f0c2b, 32'h4115e593, 32'hc2a26d8b, 32'h419d79c3, 32'hc190a0d6, 32'h4155d0ee};
test_output[5535] = '{32'h419f0c2b};
test_index[5535] = '{2};
test_input[44288:44295] = '{32'hc24473ab, 32'hc15464f2, 32'hc23d11ec, 32'hc28e7335, 32'hc2c41889, 32'hc18c0271, 32'h42894428, 32'hc292e9f9};
test_output[5536] = '{32'h42894428};
test_index[5536] = '{6};
test_input[44296:44303] = '{32'h42a012a5, 32'hc1f3c4a1, 32'hc2ba9c5d, 32'hbf9dc3b8, 32'h41637699, 32'h41f8f0dc, 32'h427d3937, 32'h40f80169};
test_output[5537] = '{32'h42a012a5};
test_index[5537] = '{0};
test_input[44304:44311] = '{32'hc1e8009e, 32'h42548870, 32'h4298c4a5, 32'hc2331426, 32'hc2b36747, 32'h41a7c38d, 32'hc2ab0d80, 32'hc25f3e46};
test_output[5538] = '{32'h4298c4a5};
test_index[5538] = '{2};
test_input[44312:44319] = '{32'h40e4cf73, 32'h42bc4335, 32'h425a7f97, 32'hc12a2d9f, 32'h3fb7ab32, 32'h410e5223, 32'hc259bee4, 32'h42ac6ce9};
test_output[5539] = '{32'h42bc4335};
test_index[5539] = '{1};
test_input[44320:44327] = '{32'h4132a427, 32'h42a09ca4, 32'hc2c6e371, 32'h4208013d, 32'hc2b9b4e3, 32'h40883bbc, 32'h4212aae3, 32'h41438299};
test_output[5540] = '{32'h42a09ca4};
test_index[5540] = '{1};
test_input[44328:44335] = '{32'h4237097e, 32'h421245a7, 32'h42904651, 32'h3ff28c4c, 32'hbebd4cf6, 32'hc2946c59, 32'h4231672c, 32'h421aac27};
test_output[5541] = '{32'h42904651};
test_index[5541] = '{2};
test_input[44336:44343] = '{32'h426a317d, 32'h4280b800, 32'h422c3b8f, 32'h421d956a, 32'h42885dc7, 32'hc21d6125, 32'h42750777, 32'h42bd0142};
test_output[5542] = '{32'h42bd0142};
test_index[5542] = '{7};
test_input[44344:44351] = '{32'hc2b7907c, 32'h41a7282d, 32'h417b5a38, 32'hc238aaa3, 32'h3f224986, 32'h41ccf084, 32'h4258295c, 32'h41066713};
test_output[5543] = '{32'h4258295c};
test_index[5543] = '{6};
test_input[44352:44359] = '{32'hc1811532, 32'h42107be9, 32'h40de4be9, 32'hc23d441a, 32'h4206035e, 32'h41c5abee, 32'hc1e86c00, 32'hc2acaf74};
test_output[5544] = '{32'h42107be9};
test_index[5544] = '{1};
test_input[44360:44367] = '{32'hc1d1511b, 32'hc240e101, 32'h42082b1a, 32'hc28998b2, 32'h4080d6a2, 32'h42acad98, 32'h423e1dc1, 32'h4125628f};
test_output[5545] = '{32'h42acad98};
test_index[5545] = '{5};
test_input[44368:44375] = '{32'hc219873d, 32'hc2a61468, 32'h428fc82c, 32'h42541e87, 32'h421508b8, 32'h42afef01, 32'h41d10b22, 32'h42886bb9};
test_output[5546] = '{32'h42afef01};
test_index[5546] = '{5};
test_input[44376:44383] = '{32'h42900b8d, 32'h416df1a3, 32'hc276c63e, 32'hc1e842e4, 32'h42a9ab86, 32'hc216224b, 32'h41d6a64c, 32'h42269762};
test_output[5547] = '{32'h42a9ab86};
test_index[5547] = '{4};
test_input[44384:44391] = '{32'hc2029954, 32'hc1c2158d, 32'hc2789cbe, 32'hc15c1948, 32'h42a76b5b, 32'hc2a8fc59, 32'h42a18f00, 32'h41d2fb23};
test_output[5548] = '{32'h42a76b5b};
test_index[5548] = '{4};
test_input[44392:44399] = '{32'hc2a19ab2, 32'hc2009630, 32'h42bec26c, 32'hc25003bc, 32'hc2a74893, 32'h4252f2af, 32'hc2c3ca0a, 32'hc243b52a};
test_output[5549] = '{32'h42bec26c};
test_index[5549] = '{2};
test_input[44400:44407] = '{32'hc16c3ad0, 32'hc29febad, 32'hc208d075, 32'hc29e58bc, 32'h3d24638d, 32'h425db592, 32'hc28d25ba, 32'hc2869d6f};
test_output[5550] = '{32'h425db592};
test_index[5550] = '{5};
test_input[44408:44415] = '{32'hc2bd2410, 32'hc1cea838, 32'h427aa316, 32'h41cd60e9, 32'hc2ad36bf, 32'h418b5165, 32'hc234fc38, 32'h4284bb99};
test_output[5551] = '{32'h4284bb99};
test_index[5551] = '{7};
test_input[44416:44423] = '{32'h428ea35e, 32'hc2986f87, 32'h4137301b, 32'h42637221, 32'hc2942990, 32'h42a0745b, 32'hc24fce02, 32'h42c18654};
test_output[5552] = '{32'h42c18654};
test_index[5552] = '{7};
test_input[44424:44431] = '{32'h42b4c05c, 32'h40d25f9a, 32'h42bb9a9e, 32'h4190463d, 32'hc2174794, 32'hc2090fa1, 32'hc2769036, 32'h42a15e1d};
test_output[5553] = '{32'h42bb9a9e};
test_index[5553] = '{2};
test_input[44432:44439] = '{32'hc29b2770, 32'h41d7d8e5, 32'hc2a2514d, 32'h4118a32c, 32'hc0a75c8e, 32'hc205c3fe, 32'h3f7ab363, 32'h4086c8ce};
test_output[5554] = '{32'h41d7d8e5};
test_index[5554] = '{1};
test_input[44440:44447] = '{32'h41caff68, 32'hc2963189, 32'hc2c620f1, 32'hc2c4e208, 32'h420f74f9, 32'hc2af17cb, 32'hc2b13bb4, 32'hc28631c6};
test_output[5555] = '{32'h420f74f9};
test_index[5555] = '{4};
test_input[44448:44455] = '{32'hc105fd60, 32'hc2a7b568, 32'h42a43e06, 32'hc2a7120f, 32'h42890f14, 32'h4289ebb5, 32'hc28305b6, 32'h42357052};
test_output[5556] = '{32'h42a43e06};
test_index[5556] = '{2};
test_input[44456:44463] = '{32'h42812dc2, 32'hc1f350a8, 32'hc2251fe1, 32'h427c03ab, 32'hc290be79, 32'h41c85217, 32'h42acfed5, 32'h42b03565};
test_output[5557] = '{32'h42b03565};
test_index[5557] = '{7};
test_input[44464:44471] = '{32'h4261c081, 32'hbf8a2230, 32'h4244cf4b, 32'h42ac7aa0, 32'h4205ba9a, 32'h4200055d, 32'hc22ff169, 32'h42a15560};
test_output[5558] = '{32'h42ac7aa0};
test_index[5558] = '{3};
test_input[44472:44479] = '{32'hc23b65f4, 32'h418d5af7, 32'h429e96ff, 32'hc242c514, 32'h4283dde2, 32'h42b7bad7, 32'hc28fbfc1, 32'hc2810893};
test_output[5559] = '{32'h42b7bad7};
test_index[5559] = '{5};
test_input[44480:44487] = '{32'h427d8eee, 32'h403d3950, 32'h429d7c48, 32'h42b55649, 32'h4172fbc4, 32'hc19d1176, 32'h427afed8, 32'h42c29862};
test_output[5560] = '{32'h42c29862};
test_index[5560] = '{7};
test_input[44488:44495] = '{32'hc136a7a0, 32'hc2444ea8, 32'hc26836b2, 32'hc1c58409, 32'hc2b73bed, 32'hc225cf14, 32'hc29c019f, 32'h41d36de5};
test_output[5561] = '{32'h41d36de5};
test_index[5561] = '{7};
test_input[44496:44503] = '{32'hc2b86251, 32'h4261d99c, 32'hc2443a85, 32'h424bfc0d, 32'hc2bfc2cb, 32'h40ef4595, 32'h42b81780, 32'h42365cdf};
test_output[5562] = '{32'h42b81780};
test_index[5562] = '{6};
test_input[44504:44511] = '{32'hc2831577, 32'h428827a4, 32'h42aa0e4c, 32'h42acd4d8, 32'h426a000d, 32'hc2bb3eb9, 32'hc2727b5f, 32'h410770b1};
test_output[5563] = '{32'h42acd4d8};
test_index[5563] = '{3};
test_input[44512:44519] = '{32'h429c343a, 32'hc1dc6b05, 32'hc2b965dc, 32'hc1aa922b, 32'hc245100c, 32'h42addd80, 32'hc2ae05ae, 32'hc1c61526};
test_output[5564] = '{32'h42addd80};
test_index[5564] = '{5};
test_input[44520:44527] = '{32'hc21abd1b, 32'hc27f8666, 32'hc254bfdf, 32'hc2be5b94, 32'h429d327b, 32'hc1904ae8, 32'hc293b99a, 32'hc170541b};
test_output[5565] = '{32'h429d327b};
test_index[5565] = '{4};
test_input[44528:44535] = '{32'h42295a52, 32'hc2199ae0, 32'hc19d2bf9, 32'hc2b6e83d, 32'hc2ab0526, 32'hc29363e1, 32'hc257ac35, 32'hbfe27b79};
test_output[5566] = '{32'h42295a52};
test_index[5566] = '{0};
test_input[44536:44543] = '{32'hc27a9cad, 32'h42b95a3d, 32'h41da0673, 32'h42411043, 32'hc2a2cfd2, 32'h41d19dbf, 32'h42108f55, 32'hc2b41060};
test_output[5567] = '{32'h42b95a3d};
test_index[5567] = '{1};
test_input[44544:44551] = '{32'h42b081e7, 32'h4284dd2f, 32'hc2c5d02a, 32'hc14bb75f, 32'hc2709fe5, 32'h420139f1, 32'h4127a642, 32'hc28e9831};
test_output[5568] = '{32'h42b081e7};
test_index[5568] = '{0};
test_input[44552:44559] = '{32'hc2c1f427, 32'hc18ff65d, 32'hc197dbd2, 32'hc292e38b, 32'hc25792c9, 32'h424ef1d3, 32'h41a68cc1, 32'h4229e8fc};
test_output[5569] = '{32'h424ef1d3};
test_index[5569] = '{5};
test_input[44560:44567] = '{32'hc2906cba, 32'h41bd32a4, 32'h421716e4, 32'hc2a8de18, 32'h420d23a3, 32'hc23c4b6e, 32'h4244330f, 32'h4065c069};
test_output[5570] = '{32'h4244330f};
test_index[5570] = '{6};
test_input[44568:44575] = '{32'h42b4dd0c, 32'h40e8c0e4, 32'hc28a77c5, 32'h42bf1667, 32'h40f814b8, 32'hc24898bb, 32'hc2b733dc, 32'h42af96ed};
test_output[5571] = '{32'h42bf1667};
test_index[5571] = '{3};
test_input[44576:44583] = '{32'h40e13b56, 32'h415acf08, 32'h415b73d9, 32'h42604151, 32'h41999fe3, 32'hc29b9a67, 32'hc28caacc, 32'hc2b647e6};
test_output[5572] = '{32'h42604151};
test_index[5572] = '{3};
test_input[44584:44591] = '{32'hc2a3eec8, 32'hc146f28c, 32'hc29430d2, 32'hc2a7f655, 32'hc0462a26, 32'h419a3a78, 32'hc2c0d3bd, 32'hc180aeb3};
test_output[5573] = '{32'h419a3a78};
test_index[5573] = '{5};
test_input[44592:44599] = '{32'hc1e9865c, 32'h42c316be, 32'h42b73c47, 32'hc1c9edf4, 32'h42580c12, 32'h420c51f0, 32'hc21ab941, 32'h41554b7f};
test_output[5574] = '{32'h42c316be};
test_index[5574] = '{1};
test_input[44600:44607] = '{32'h424df43e, 32'hc2652e89, 32'hc20ae897, 32'hc238aea1, 32'h4289de0c, 32'h420cdb84, 32'hc2490f3b, 32'h41781507};
test_output[5575] = '{32'h4289de0c};
test_index[5575] = '{4};
test_input[44608:44615] = '{32'h420b507a, 32'hc2b01866, 32'hc2c12df6, 32'hc2ab7dfd, 32'h424b2826, 32'h42b82dec, 32'h41bf56ad, 32'h413db223};
test_output[5576] = '{32'h42b82dec};
test_index[5576] = '{5};
test_input[44616:44623] = '{32'h42c66579, 32'hc22ff44a, 32'hc264e12b, 32'h4266353d, 32'h417a6901, 32'hc252c9b5, 32'h42c587fb, 32'hc1f2ac59};
test_output[5577] = '{32'h42c66579};
test_index[5577] = '{0};
test_input[44624:44631] = '{32'hc2882fec, 32'hc2a8c394, 32'h429c14e7, 32'h42401adc, 32'h418e5663, 32'h3fafd7ee, 32'hc21d38fe, 32'h429a8dc5};
test_output[5578] = '{32'h429c14e7};
test_index[5578] = '{2};
test_input[44632:44639] = '{32'h42736f67, 32'h4234dcf2, 32'hc13e1ced, 32'hc168f2a5, 32'hc28bc38f, 32'hc15ca376, 32'hc22301ee, 32'hc1c83895};
test_output[5579] = '{32'h42736f67};
test_index[5579] = '{0};
test_input[44640:44647] = '{32'hc1798873, 32'hc02bbd7f, 32'hc2afe4bb, 32'h426d8d24, 32'hc2bac533, 32'h42717fbf, 32'h429560c4, 32'h420bfb08};
test_output[5580] = '{32'h429560c4};
test_index[5580] = '{6};
test_input[44648:44655] = '{32'hc23c9231, 32'h428da059, 32'hc20d36fd, 32'h41fac7ec, 32'h42af0a9f, 32'h41c6607f, 32'h42621a29, 32'h41cc7038};
test_output[5581] = '{32'h42af0a9f};
test_index[5581] = '{4};
test_input[44656:44663] = '{32'hc1cbc979, 32'h421bc744, 32'hc2407dee, 32'hc1902e6b, 32'hbfaedf4b, 32'hc1180107, 32'hc2930987, 32'hc281749d};
test_output[5582] = '{32'h421bc744};
test_index[5582] = '{1};
test_input[44664:44671] = '{32'h42001455, 32'h421929c1, 32'h424bd207, 32'hc2b90ba4, 32'h42528a57, 32'h420e06e9, 32'hc2643899, 32'h3ffbd147};
test_output[5583] = '{32'h42528a57};
test_index[5583] = '{4};
test_input[44672:44679] = '{32'hc08285a4, 32'hc29c5aed, 32'hc28ae419, 32'h4250b4a4, 32'h40c94cc6, 32'hc2be2b2d, 32'hc1cdca26, 32'hc2ae474d};
test_output[5584] = '{32'h4250b4a4};
test_index[5584] = '{3};
test_input[44680:44687] = '{32'hc2268cbb, 32'h42325980, 32'hc1f968c0, 32'h42c7d4af, 32'h424a5a60, 32'hc0dd43a5, 32'hc12dcba2, 32'hc25b5936};
test_output[5585] = '{32'h42c7d4af};
test_index[5585] = '{3};
test_input[44688:44695] = '{32'hc1b1777e, 32'hc0c0b564, 32'h428127a2, 32'h42571975, 32'hc2abf1f6, 32'hc2926a2a, 32'hc2ba51e8, 32'hc25c53cf};
test_output[5586] = '{32'h428127a2};
test_index[5586] = '{2};
test_input[44696:44703] = '{32'hc1da3ca3, 32'hc2167638, 32'h425fd4c6, 32'hc1549df7, 32'h426c0a40, 32'hc2b96c37, 32'h42731b47, 32'hc2ab19aa};
test_output[5587] = '{32'h42731b47};
test_index[5587] = '{6};
test_input[44704:44711] = '{32'h405e076d, 32'h427e7b7d, 32'hc29a6ea6, 32'hc1a3ee71, 32'h42b2e5f8, 32'hc11f1cf7, 32'hc2ae294d, 32'h42673cc8};
test_output[5588] = '{32'h42b2e5f8};
test_index[5588] = '{4};
test_input[44712:44719] = '{32'hc21bd0a3, 32'hc24d1a82, 32'h428bd3c9, 32'h4231503f, 32'h41972bf1, 32'h418a07b3, 32'h4213c908, 32'hc2aff82f};
test_output[5589] = '{32'h428bd3c9};
test_index[5589] = '{2};
test_input[44720:44727] = '{32'hc246c27b, 32'h42aa81d2, 32'h428647f3, 32'h428835d9, 32'h425db03b, 32'hc2853b6d, 32'h424ded7e, 32'h41241569};
test_output[5590] = '{32'h42aa81d2};
test_index[5590] = '{1};
test_input[44728:44735] = '{32'hc12d24d3, 32'hc264cf9e, 32'hc2114f39, 32'h4298d50a, 32'h426ec51a, 32'hc2b703cc, 32'h428ca3e5, 32'h4296d9b0};
test_output[5591] = '{32'h4298d50a};
test_index[5591] = '{3};
test_input[44736:44743] = '{32'hc223de10, 32'h424500a7, 32'hc21c7c4a, 32'hc216d72a, 32'hc235eb52, 32'h42c04571, 32'h40d46fa1, 32'h3fa44a88};
test_output[5592] = '{32'h42c04571};
test_index[5592] = '{5};
test_input[44744:44751] = '{32'hc282afe9, 32'hc2c5a4fd, 32'hc2829b6b, 32'hc2988cfe, 32'hc2893bea, 32'h4204651e, 32'h427b6ff7, 32'hc296b21d};
test_output[5593] = '{32'h427b6ff7};
test_index[5593] = '{6};
test_input[44752:44759] = '{32'h423bdb8d, 32'h42a25c5c, 32'hc1b0bcfe, 32'h42c2e937, 32'hc20a1c86, 32'h4204a81b, 32'h410ff029, 32'hc0ec8039};
test_output[5594] = '{32'h42c2e937};
test_index[5594] = '{3};
test_input[44760:44767] = '{32'h427aceba, 32'hc2c53f84, 32'h41825d8e, 32'h42180300, 32'h421865df, 32'hc17a8fe2, 32'h42bd7196, 32'hc282f39f};
test_output[5595] = '{32'h42bd7196};
test_index[5595] = '{6};
test_input[44768:44775] = '{32'h41e76dab, 32'hc2af7bfe, 32'hc0c47180, 32'h41ce8219, 32'h41aa3975, 32'hc2aa1eff, 32'h419d95f8, 32'hc17a4330};
test_output[5596] = '{32'h41e76dab};
test_index[5596] = '{0};
test_input[44776:44783] = '{32'hc0bb9da2, 32'hc272719c, 32'h426ee75b, 32'hc2aef105, 32'h42c2cd0a, 32'h424c5099, 32'hc23888a1, 32'hc2c5e700};
test_output[5597] = '{32'h42c2cd0a};
test_index[5597] = '{4};
test_input[44784:44791] = '{32'h423e90ef, 32'hc29583de, 32'hc2500e7e, 32'hc1986c43, 32'hc23eb0d3, 32'hc2679b00, 32'h424468b0, 32'h41fbe58f};
test_output[5598] = '{32'h424468b0};
test_index[5598] = '{6};
test_input[44792:44799] = '{32'h409f518a, 32'h40f61734, 32'h41d81aa9, 32'h3f171142, 32'hbfa560d1, 32'hc2bc4e88, 32'hc2b6d763, 32'h429a0b0d};
test_output[5599] = '{32'h429a0b0d};
test_index[5599] = '{7};
test_input[44800:44807] = '{32'h423425e5, 32'hc29ddfe8, 32'h416ca410, 32'hbf39dffb, 32'hc26d5e31, 32'hc2b89bf2, 32'h41cedb34, 32'hc2c30eb9};
test_output[5600] = '{32'h423425e5};
test_index[5600] = '{0};
test_input[44808:44815] = '{32'h41094120, 32'h42980911, 32'h4186eda5, 32'hc290d497, 32'hc2977a6d, 32'h4140bfbf, 32'h42a6653c, 32'h41fa6b2d};
test_output[5601] = '{32'h42a6653c};
test_index[5601] = '{6};
test_input[44816:44823] = '{32'h421cec1e, 32'h42c34b0a, 32'h41d66e24, 32'h42a0ecfd, 32'h427b19a6, 32'h413a2c38, 32'hc10de706, 32'hc1f55e19};
test_output[5602] = '{32'h42c34b0a};
test_index[5602] = '{1};
test_input[44824:44831] = '{32'hc216f7c1, 32'hc2c7e63d, 32'hc1b108c4, 32'h42bfb069, 32'hc253c9d9, 32'h41031494, 32'h42919b00, 32'hc2bdec5e};
test_output[5603] = '{32'h42bfb069};
test_index[5603] = '{3};
test_input[44832:44839] = '{32'hc2b5a307, 32'h42a9c30d, 32'hc20113e5, 32'h40801eea, 32'hc23945c9, 32'h3efca4e8, 32'hc202d247, 32'hc27d73c5};
test_output[5604] = '{32'h42a9c30d};
test_index[5604] = '{1};
test_input[44840:44847] = '{32'hc28e8067, 32'h4232632d, 32'hc25a10cc, 32'h42c13120, 32'hc29dcc11, 32'h42084964, 32'h429a4acd, 32'hc231b5bb};
test_output[5605] = '{32'h42c13120};
test_index[5605] = '{3};
test_input[44848:44855] = '{32'h422ccea5, 32'h42a1458c, 32'hc20ede02, 32'hc1002401, 32'hc2a68cea, 32'hc2539ff3, 32'hc28417ea, 32'h423258ea};
test_output[5606] = '{32'h42a1458c};
test_index[5606] = '{1};
test_input[44856:44863] = '{32'h41e344b8, 32'h420d288a, 32'h42272f95, 32'h413a2521, 32'h42bbe854, 32'h42837cd4, 32'hc2c5e4c3, 32'h42c1d039};
test_output[5607] = '{32'h42c1d039};
test_index[5607] = '{7};
test_input[44864:44871] = '{32'hc230bb7f, 32'h4261b385, 32'h4267d67d, 32'h41e9ee4a, 32'h41e19f24, 32'hc2b67f43, 32'h4170c8ab, 32'h4273deac};
test_output[5608] = '{32'h4273deac};
test_index[5608] = '{7};
test_input[44872:44879] = '{32'hc1bc0272, 32'h422c1cde, 32'hc22fb232, 32'hc24ae2fc, 32'h42246c5e, 32'hc23f6e5d, 32'hc28937b8, 32'hc0abe7e5};
test_output[5609] = '{32'h422c1cde};
test_index[5609] = '{1};
test_input[44880:44887] = '{32'h40e1a8b3, 32'hc141d69a, 32'hc2a77ae7, 32'hc26670f2, 32'hc282ac3b, 32'h4123cae1, 32'h4222dae4, 32'h423a9597};
test_output[5610] = '{32'h423a9597};
test_index[5610] = '{7};
test_input[44888:44895] = '{32'h42bdea2d, 32'hc1f6d071, 32'h4090fe51, 32'h429c0a61, 32'hc21fc815, 32'hc1f545da, 32'h426bc955, 32'hc2444ff2};
test_output[5611] = '{32'h42bdea2d};
test_index[5611] = '{0};
test_input[44896:44903] = '{32'h428ed06e, 32'hc2b646ab, 32'h420ee6a5, 32'h420b8e29, 32'hc2369635, 32'hc289ddeb, 32'h4286ea8b, 32'h427f26a5};
test_output[5612] = '{32'h428ed06e};
test_index[5612] = '{0};
test_input[44904:44911] = '{32'hc1e53f96, 32'hc2c44877, 32'hc29a12f1, 32'hbfe4dcdb, 32'h4056274c, 32'hc140827b, 32'h42731308, 32'h3efc9332};
test_output[5613] = '{32'h42731308};
test_index[5613] = '{6};
test_input[44912:44919] = '{32'h417e8d12, 32'hc281ac20, 32'h428ad671, 32'h41117801, 32'hc2a36e03, 32'hc086c44d, 32'hc29d7910, 32'hc271cb16};
test_output[5614] = '{32'h428ad671};
test_index[5614] = '{2};
test_input[44920:44927] = '{32'hc2aeca7f, 32'h4206d3ab, 32'h4252817f, 32'hc2581126, 32'h427f6c3b, 32'h417abe1e, 32'hc1d87e07, 32'h422967e1};
test_output[5615] = '{32'h427f6c3b};
test_index[5615] = '{4};
test_input[44928:44935] = '{32'hc192717e, 32'h4274dcfd, 32'h428145b8, 32'hc2bb0b28, 32'hc2aa4647, 32'hc284e903, 32'h4189ed69, 32'h40ab2fb1};
test_output[5616] = '{32'h428145b8};
test_index[5616] = '{2};
test_input[44936:44943] = '{32'hc1fd2b21, 32'h42b67d3c, 32'hc1c73cb7, 32'hc072c6b2, 32'hc290e61b, 32'h42a6a689, 32'h42a04d82, 32'hc28de192};
test_output[5617] = '{32'h42b67d3c};
test_index[5617] = '{1};
test_input[44944:44951] = '{32'hc24c1104, 32'hc2912f3b, 32'hc1642b36, 32'h42518e5c, 32'hc2afcbcc, 32'hc17b947d, 32'h41f5655c, 32'hc20ffd71};
test_output[5618] = '{32'h42518e5c};
test_index[5618] = '{3};
test_input[44952:44959] = '{32'hc2a99466, 32'hc1f63b61, 32'h42c48cf2, 32'hc1b7cd46, 32'h42435f8a, 32'hc23a789b, 32'h41abd35b, 32'h42acace1};
test_output[5619] = '{32'h42c48cf2};
test_index[5619] = '{2};
test_input[44960:44967] = '{32'h3fe2ea3f, 32'h421e57bf, 32'h42c707b7, 32'h412dfab6, 32'h42bddfc8, 32'h4294881c, 32'h42a8ff87, 32'h4201aeef};
test_output[5620] = '{32'h42c707b7};
test_index[5620] = '{2};
test_input[44968:44975] = '{32'h4278df15, 32'h4290d684, 32'hc1a57002, 32'hc23b528c, 32'h4234a495, 32'h428be7a3, 32'hc27cd126, 32'hc2ba2405};
test_output[5621] = '{32'h4290d684};
test_index[5621] = '{1};
test_input[44976:44983] = '{32'h41afd986, 32'h41d686bd, 32'h420bf316, 32'hc1ebea2a, 32'h4227b41d, 32'h42c2bbc5, 32'h4246b3b6, 32'h422ebb4a};
test_output[5622] = '{32'h42c2bbc5};
test_index[5622] = '{5};
test_input[44984:44991] = '{32'h425da605, 32'h41725e5c, 32'hc29e8189, 32'hc2989c35, 32'hc2c48638, 32'hc2a781ae, 32'hc28bfece, 32'h41b8047e};
test_output[5623] = '{32'h425da605};
test_index[5623] = '{0};
test_input[44992:44999] = '{32'h42999a23, 32'hc216d096, 32'h42827e25, 32'hc29a79a9, 32'hc2a5a43e, 32'h4299c5a7, 32'hc04fc593, 32'hc25f231a};
test_output[5624] = '{32'h4299c5a7};
test_index[5624] = '{5};
test_input[45000:45007] = '{32'hc203b811, 32'h410ec81e, 32'hc2a1f444, 32'hc2b76478, 32'hc2a75edd, 32'h428c7dd9, 32'hc224b898, 32'h412fc045};
test_output[5625] = '{32'h428c7dd9};
test_index[5625] = '{5};
test_input[45008:45015] = '{32'h42974fd0, 32'hbf98899a, 32'h422f4cc9, 32'hc26706fb, 32'h42024ac0, 32'hc2aad4ff, 32'hc1dc62dc, 32'h42807023};
test_output[5626] = '{32'h42974fd0};
test_index[5626] = '{0};
test_input[45016:45023] = '{32'h429c1ef3, 32'h3f9fb716, 32'hc1b2bb89, 32'hc2b71ff1, 32'h420ce65d, 32'h41e273e8, 32'hc24f12d4, 32'hc274f1d8};
test_output[5627] = '{32'h429c1ef3};
test_index[5627] = '{0};
test_input[45024:45031] = '{32'h40fb7991, 32'h41e5390f, 32'h42bb7a81, 32'hc2ae1af9, 32'h42a97341, 32'h429a499c, 32'h418fad5e, 32'h428de751};
test_output[5628] = '{32'h42bb7a81};
test_index[5628] = '{2};
test_input[45032:45039] = '{32'h4213dbdc, 32'h417d0a8e, 32'h413729ff, 32'hc238522b, 32'hc0a02c6d, 32'h425c9d97, 32'h423e7fba, 32'h4270c58a};
test_output[5629] = '{32'h4270c58a};
test_index[5629] = '{7};
test_input[45040:45047] = '{32'h428f9f52, 32'h40ff78dd, 32'h4210640f, 32'h41aee71c, 32'h42311258, 32'hc282d4f3, 32'h422fc14e, 32'h40ec0144};
test_output[5630] = '{32'h428f9f52};
test_index[5630] = '{0};
test_input[45048:45055] = '{32'hc283ef24, 32'h42386d47, 32'hc230c93e, 32'h42c60188, 32'hc2c70da1, 32'hc25e3c2b, 32'h42313280, 32'h429b222b};
test_output[5631] = '{32'h42c60188};
test_index[5631] = '{3};
test_input[45056:45063] = '{32'h42bffeeb, 32'hc2336dce, 32'h4153d4cd, 32'h42c4fe51, 32'hc1e355d1, 32'h4271e655, 32'hc2b40e05, 32'h41f16ab4};
test_output[5632] = '{32'h42c4fe51};
test_index[5632] = '{3};
test_input[45064:45071] = '{32'hc1b3acce, 32'hc2b60fff, 32'hc13d53d1, 32'h4211b8c3, 32'hc2841c54, 32'h42715ea0, 32'h42c08568, 32'h42aacd74};
test_output[5633] = '{32'h42c08568};
test_index[5633] = '{6};
test_input[45072:45079] = '{32'hc200d78e, 32'h420f4906, 32'h4255b6c8, 32'h4201f57b, 32'hc24e2c47, 32'hc2a735c0, 32'hc18b59d2, 32'hc09d1172};
test_output[5634] = '{32'h4255b6c8};
test_index[5634] = '{2};
test_input[45080:45087] = '{32'hc2244ff6, 32'hc2926302, 32'hc2722e25, 32'h425507cb, 32'hc2c1aabd, 32'h427f188e, 32'hc1c584d0, 32'hc23c5c08};
test_output[5635] = '{32'h427f188e};
test_index[5635] = '{5};
test_input[45088:45095] = '{32'hc165a511, 32'hc2b3bedb, 32'h42872d3e, 32'hc2766d15, 32'hc1c963c1, 32'hc01c695d, 32'h412abfbc, 32'h429ad80e};
test_output[5636] = '{32'h429ad80e};
test_index[5636] = '{7};
test_input[45096:45103] = '{32'h421a658b, 32'h421d60a5, 32'h41de5887, 32'h42c2e1f1, 32'hc2bb279e, 32'h424630e7, 32'h4260eb59, 32'hc2a6422b};
test_output[5637] = '{32'h42c2e1f1};
test_index[5637] = '{3};
test_input[45104:45111] = '{32'hc2461614, 32'hc1c56409, 32'h41cd5442, 32'hc298e756, 32'hc21ab505, 32'hc2b40162, 32'h42a3803f, 32'h421bc760};
test_output[5638] = '{32'h42a3803f};
test_index[5638] = '{6};
test_input[45112:45119] = '{32'hc246b73c, 32'h4287cdb7, 32'hc2b68bcc, 32'h4296bb8c, 32'h40a1407c, 32'h429becf6, 32'hc01ec6db, 32'h41a9eecc};
test_output[5639] = '{32'h429becf6};
test_index[5639] = '{5};
test_input[45120:45127] = '{32'hbf232166, 32'hc2b47d99, 32'h42083958, 32'hc28e6d7b, 32'hc16ca5f8, 32'hc22e137e, 32'hc22d8069, 32'h4262d5a2};
test_output[5640] = '{32'h4262d5a2};
test_index[5640] = '{7};
test_input[45128:45135] = '{32'hc2be9224, 32'hc290b5b8, 32'h429716eb, 32'hc2c0e1d7, 32'hc23aa920, 32'hc251cd9d, 32'h41534592, 32'hc2c77fc6};
test_output[5641] = '{32'h429716eb};
test_index[5641] = '{2};
test_input[45136:45143] = '{32'h41e8b33c, 32'h422b0ff6, 32'hc1f3609d, 32'h42654e89, 32'h41b35a49, 32'h41e38b75, 32'hbf800c94, 32'h429fa6f0};
test_output[5642] = '{32'h429fa6f0};
test_index[5642] = '{7};
test_input[45144:45151] = '{32'h42b10de4, 32'h41202385, 32'hc29536ea, 32'hc17cc9e1, 32'h429b1da3, 32'hc2affa86, 32'hc0ee45ee, 32'h41a95f30};
test_output[5643] = '{32'h42b10de4};
test_index[5643] = '{0};
test_input[45152:45159] = '{32'hc13e30f8, 32'h42b2084c, 32'h42b3a3d5, 32'hc0254bb9, 32'hc2a5a8b4, 32'hc16a9e3f, 32'h41d8c6c5, 32'h425ee32c};
test_output[5644] = '{32'h42b3a3d5};
test_index[5644] = '{2};
test_input[45160:45167] = '{32'h42777c8c, 32'hc21d1736, 32'h428f20b1, 32'hc2bc48a7, 32'hc0deab90, 32'hc2aadab1, 32'hc2b1e728, 32'hc26a666b};
test_output[5645] = '{32'h428f20b1};
test_index[5645] = '{2};
test_input[45168:45175] = '{32'hc281a978, 32'hc2711b73, 32'h42516e00, 32'hc2817323, 32'h42b7342e, 32'hc27e153b, 32'h42bddd8f, 32'hc277a476};
test_output[5646] = '{32'h42bddd8f};
test_index[5646] = '{6};
test_input[45176:45183] = '{32'h41c6cb25, 32'hc094f64d, 32'hc2135ece, 32'h41b80ebc, 32'hc24f33fb, 32'h42be8120, 32'hc2824736, 32'h42c6575d};
test_output[5647] = '{32'h42c6575d};
test_index[5647] = '{7};
test_input[45184:45191] = '{32'h42048f32, 32'h42a71489, 32'h421d4a17, 32'h41ebca62, 32'h40935f9c, 32'hc26e8ec0, 32'hc111600b, 32'hc21125f5};
test_output[5648] = '{32'h42a71489};
test_index[5648] = '{1};
test_input[45192:45199] = '{32'hc293232c, 32'h428ec4b1, 32'h4282a6fc, 32'h42c19903, 32'hc21e058b, 32'hc042a271, 32'hc25dc1dc, 32'h424edc55};
test_output[5649] = '{32'h42c19903};
test_index[5649] = '{3};
test_input[45200:45207] = '{32'hc15db258, 32'h42b84332, 32'h428a0b4f, 32'hc2b3d4e2, 32'h42848638, 32'h4251ebbf, 32'hc20c6275, 32'hc2159122};
test_output[5650] = '{32'h42b84332};
test_index[5650] = '{1};
test_input[45208:45215] = '{32'hc2b2c74a, 32'h4274eee3, 32'hc1f8a5b1, 32'h42865d2d, 32'hc2929d16, 32'hc20863f6, 32'h412d7be9, 32'hc21549dd};
test_output[5651] = '{32'h42865d2d};
test_index[5651] = '{3};
test_input[45216:45223] = '{32'hc27c567f, 32'hc2975a49, 32'h42b9947b, 32'h42c2ebad, 32'h40b3c748, 32'hc21c43e4, 32'hc1f167eb, 32'hc2225c27};
test_output[5652] = '{32'h42c2ebad};
test_index[5652] = '{3};
test_input[45224:45231] = '{32'h4292f58c, 32'h41ba5ca6, 32'h419673ab, 32'h420ad6c9, 32'h426c90aa, 32'hc2b24b0e, 32'h41c8c318, 32'h42053402};
test_output[5653] = '{32'h4292f58c};
test_index[5653] = '{0};
test_input[45232:45239] = '{32'hc2925584, 32'hc2c74c4a, 32'h4183a5da, 32'hc28405ae, 32'hc1264d1a, 32'hc285d3c5, 32'h42af7ec7, 32'h41bd5ec5};
test_output[5654] = '{32'h42af7ec7};
test_index[5654] = '{6};
test_input[45240:45247] = '{32'h42588990, 32'hc22200e6, 32'hc2015831, 32'hc247db6c, 32'h41f0d53e, 32'h42497a28, 32'h412f721f, 32'hc2b53848};
test_output[5655] = '{32'h42588990};
test_index[5655] = '{0};
test_input[45248:45255] = '{32'hc24a4c2c, 32'h4290bac6, 32'h42959960, 32'hc273c58d, 32'h4185cfc7, 32'h4150d222, 32'hc24661c7, 32'h42286503};
test_output[5656] = '{32'h42959960};
test_index[5656] = '{2};
test_input[45256:45263] = '{32'hc1eb3792, 32'h42808dd8, 32'h41c73c93, 32'hc1c2089f, 32'h41361bb7, 32'h4224b3da, 32'h428dc1d5, 32'hc25cf29b};
test_output[5657] = '{32'h428dc1d5};
test_index[5657] = '{6};
test_input[45264:45271] = '{32'hc2bd6256, 32'h4228e4f3, 32'h425e34b6, 32'h41686bf6, 32'hc1a48207, 32'h429d49f0, 32'hc28d173f, 32'h4181a64c};
test_output[5658] = '{32'h429d49f0};
test_index[5658] = '{5};
test_input[45272:45279] = '{32'h429aa056, 32'h41b508ac, 32'h428bde5a, 32'h428fb6e0, 32'hc1212fc3, 32'h412d6758, 32'h4241d80a, 32'h40d23d05};
test_output[5659] = '{32'h429aa056};
test_index[5659] = '{0};
test_input[45280:45287] = '{32'hc2b2fe78, 32'h42254d42, 32'h428469ca, 32'h42a472d7, 32'hc22cb1f7, 32'h41aeed42, 32'h42316c34, 32'hc2b8422e};
test_output[5660] = '{32'h42a472d7};
test_index[5660] = '{3};
test_input[45288:45295] = '{32'h42746585, 32'h420e3332, 32'h423af0ac, 32'hc10c3b46, 32'hc2b95287, 32'hc265ef10, 32'hc2ba18da, 32'hc2bf422c};
test_output[5661] = '{32'h42746585};
test_index[5661] = '{0};
test_input[45296:45303] = '{32'h42741167, 32'hc239948e, 32'h427077ba, 32'hc26158de, 32'hc273377b, 32'hc1202858, 32'hc205cddb, 32'hc026a178};
test_output[5662] = '{32'h42741167};
test_index[5662] = '{0};
test_input[45304:45311] = '{32'h42ad9694, 32'h42885ef6, 32'hc18e0238, 32'h42972382, 32'h421f5d26, 32'h424a9ac7, 32'hc21b4af1, 32'hc1fb19aa};
test_output[5663] = '{32'h42ad9694};
test_index[5663] = '{0};
test_input[45312:45319] = '{32'hc2215383, 32'hc1c861c1, 32'hc22d54b1, 32'h428d1157, 32'h4248411e, 32'h429be129, 32'hc29acf69, 32'hc2aa96ae};
test_output[5664] = '{32'h429be129};
test_index[5664] = '{5};
test_input[45320:45327] = '{32'h428b6b16, 32'hc29dcda8, 32'h4276d39f, 32'hc1eb298c, 32'hc1f4857b, 32'hc28da7bd, 32'h3b8a2d4a, 32'h42365cbb};
test_output[5665] = '{32'h428b6b16};
test_index[5665] = '{0};
test_input[45328:45335] = '{32'h41db405c, 32'hc13a82e4, 32'h412ea8b0, 32'h424c5b16, 32'h4269b64a, 32'hc18569d0, 32'hc251ab21, 32'hc24b4f53};
test_output[5666] = '{32'h4269b64a};
test_index[5666] = '{4};
test_input[45336:45343] = '{32'hc221c432, 32'h429ebcaf, 32'hc15b3103, 32'h4204630a, 32'h42a1305f, 32'h40b5c0a6, 32'h42540eca, 32'h42498f99};
test_output[5667] = '{32'h42a1305f};
test_index[5667] = '{4};
test_input[45344:45351] = '{32'hc21e6695, 32'h427b4901, 32'hc296fc7c, 32'hc27bc73a, 32'h40ce6004, 32'h41ba6a51, 32'hc24435c4, 32'hc1a37a75};
test_output[5668] = '{32'h427b4901};
test_index[5668] = '{1};
test_input[45352:45359] = '{32'hc1be916e, 32'hc21609b8, 32'hc2066024, 32'h42b35d04, 32'h42c73478, 32'h428a1f16, 32'hc2b3d59a, 32'h4190c3ee};
test_output[5669] = '{32'h42c73478};
test_index[5669] = '{4};
test_input[45360:45367] = '{32'hc1a13077, 32'h4144ad35, 32'h428cb577, 32'h4271d2df, 32'h42bebf5e, 32'h427b89b9, 32'h42a8a56f, 32'hc102122b};
test_output[5670] = '{32'h42bebf5e};
test_index[5670] = '{4};
test_input[45368:45375] = '{32'h42ac0b01, 32'h41d8d620, 32'hc2a62268, 32'hc2c7f419, 32'h410d68f9, 32'h41fd1376, 32'h41f6d21d, 32'hc2bd4b41};
test_output[5671] = '{32'h42ac0b01};
test_index[5671] = '{0};
test_input[45376:45383] = '{32'hc28dfee1, 32'h414ec021, 32'h41c5c260, 32'h41b29cf0, 32'h4298d44b, 32'hc1ddaaff, 32'hc231c3dc, 32'h40456a0e};
test_output[5672] = '{32'h4298d44b};
test_index[5672] = '{4};
test_input[45384:45391] = '{32'h420bd07b, 32'h4213f319, 32'h42bcaa24, 32'hc2c5134f, 32'hc224b5c5, 32'hc146f7ab, 32'h42b906e8, 32'h40a9e5ab};
test_output[5673] = '{32'h42bcaa24};
test_index[5673] = '{2};
test_input[45392:45399] = '{32'hc255c951, 32'h42895127, 32'h42a136f0, 32'h411dff84, 32'hc286b802, 32'hc0b5d231, 32'h420fa92f, 32'hc2c26725};
test_output[5674] = '{32'h42a136f0};
test_index[5674] = '{2};
test_input[45400:45407] = '{32'hc2b4c4f3, 32'h41c20757, 32'hc281c76e, 32'h418397ba, 32'h4218419a, 32'h424eee06, 32'h429a85ec, 32'hc29717d0};
test_output[5675] = '{32'h429a85ec};
test_index[5675] = '{6};
test_input[45408:45415] = '{32'h423664f0, 32'h4282cba1, 32'h424173c8, 32'h42422df7, 32'h42ad6f4d, 32'h42892ba1, 32'h42b4af94, 32'hc2ae2de4};
test_output[5676] = '{32'h42b4af94};
test_index[5676] = '{6};
test_input[45416:45423] = '{32'h424ff118, 32'h42202a0c, 32'h41561dca, 32'hc2959835, 32'h3f1a5a7a, 32'hc1b18f24, 32'h42917d06, 32'h41983d7d};
test_output[5677] = '{32'h42917d06};
test_index[5677] = '{6};
test_input[45424:45431] = '{32'hc2c53fa5, 32'hc2743549, 32'h427851eb, 32'h4238a535, 32'h41307c16, 32'h426f2191, 32'h42c0664b, 32'hc1035ace};
test_output[5678] = '{32'h42c0664b};
test_index[5678] = '{6};
test_input[45432:45439] = '{32'h4150a00b, 32'hc29a7c6b, 32'h4152dccf, 32'hc28c92f7, 32'hc2c7b41c, 32'hc17064cf, 32'h41eaa93c, 32'hc1a1fcb9};
test_output[5679] = '{32'h41eaa93c};
test_index[5679] = '{6};
test_input[45440:45447] = '{32'h41addc9e, 32'hc28fb03e, 32'h427c5890, 32'h42be12b6, 32'h40ae8ea2, 32'h4127cd3a, 32'hc236bdc7, 32'hc20dd7e4};
test_output[5680] = '{32'h42be12b6};
test_index[5680] = '{3};
test_input[45448:45455] = '{32'h40c24eb4, 32'hc2535821, 32'h41fb3c31, 32'hc28f858b, 32'hc1c7a40e, 32'hc1255727, 32'h42361d56, 32'hc251ccdd};
test_output[5681] = '{32'h42361d56};
test_index[5681] = '{6};
test_input[45456:45463] = '{32'hc21627c8, 32'hc2a676e6, 32'hc28e9764, 32'hc179a620, 32'hc2108b67, 32'h42a79466, 32'hc28adae3, 32'h4214be9f};
test_output[5682] = '{32'h42a79466};
test_index[5682] = '{5};
test_input[45464:45471] = '{32'h4193811c, 32'hc250fd4f, 32'h425037ab, 32'hc29e047d, 32'h423a9895, 32'hc29e42a6, 32'hc1b2b32a, 32'hc231bdf2};
test_output[5683] = '{32'h425037ab};
test_index[5683] = '{2};
test_input[45472:45479] = '{32'hc2805c6d, 32'h4204ed4e, 32'h41e5b0d2, 32'hc2527f73, 32'h429c8a46, 32'h4130e660, 32'h429bc26a, 32'hc22af419};
test_output[5684] = '{32'h429c8a46};
test_index[5684] = '{4};
test_input[45480:45487] = '{32'hc217ad1d, 32'h42990909, 32'h422d8327, 32'hc2897326, 32'hbfd87587, 32'hc29c3b82, 32'h4272252c, 32'hc297a5ac};
test_output[5685] = '{32'h42990909};
test_index[5685] = '{1};
test_input[45488:45495] = '{32'hc28e96b7, 32'hc2901e5c, 32'h42929d23, 32'h42a07ca7, 32'h42a2e370, 32'hc278d814, 32'hc20220e2, 32'h427872f4};
test_output[5686] = '{32'h42a2e370};
test_index[5686] = '{4};
test_input[45496:45503] = '{32'h42a99fb2, 32'h42454921, 32'h4204a2cc, 32'h42b1c38d, 32'hc112419f, 32'h4298916f, 32'h4240b8d3, 32'h4219d6a3};
test_output[5687] = '{32'h42b1c38d};
test_index[5687] = '{3};
test_input[45504:45511] = '{32'hc21503b4, 32'h42b37740, 32'hc26785b3, 32'h42723664, 32'h4255b5a4, 32'hc189a0f8, 32'hc1b7d458, 32'hc1389fa5};
test_output[5688] = '{32'h42b37740};
test_index[5688] = '{1};
test_input[45512:45519] = '{32'h421d8450, 32'hc1b570cf, 32'h428ce34b, 32'hc24323bf, 32'h4285ed6f, 32'hc296d9ae, 32'hc27029ca, 32'h41e09c1c};
test_output[5689] = '{32'h428ce34b};
test_index[5689] = '{2};
test_input[45520:45527] = '{32'h4224f2f2, 32'hc1a5756c, 32'h3ffa038d, 32'h41978d7d, 32'h4269e27b, 32'h4188c2c0, 32'h41921ea3, 32'hc29c4b4d};
test_output[5690] = '{32'h4269e27b};
test_index[5690] = '{4};
test_input[45528:45535] = '{32'h41cb2275, 32'h421f6a8a, 32'hc273404a, 32'hc23dd198, 32'hc21af8cc, 32'hc19f85fb, 32'h42bc52e3, 32'h41a6a868};
test_output[5691] = '{32'h42bc52e3};
test_index[5691] = '{6};
test_input[45536:45543] = '{32'hc0d14251, 32'h40894892, 32'h40adce91, 32'hc26fdeec, 32'h41ddbb31, 32'h427256f1, 32'hc1b124b9, 32'h41bc8e61};
test_output[5692] = '{32'h427256f1};
test_index[5692] = '{5};
test_input[45544:45551] = '{32'hc00cba53, 32'h42330992, 32'hc2896595, 32'hc1ddff42, 32'h42b4a9d6, 32'h40835a32, 32'hc27fbcde, 32'h408cb8f3};
test_output[5693] = '{32'h42b4a9d6};
test_index[5693] = '{4};
test_input[45552:45559] = '{32'h424626e9, 32'hc21e6237, 32'hc21441bc, 32'h41f20040, 32'h423a3237, 32'h416d9511, 32'hc2575e55, 32'h42ba72d0};
test_output[5694] = '{32'h42ba72d0};
test_index[5694] = '{7};
test_input[45560:45567] = '{32'hc2bc092b, 32'hc2a88ae9, 32'hc2c28eac, 32'h42bf7cc6, 32'h41c62dfe, 32'hc1fbdcc0, 32'hc2a89d11, 32'hc2bb7706};
test_output[5695] = '{32'h42bf7cc6};
test_index[5695] = '{3};
test_input[45568:45575] = '{32'h42bce536, 32'hc1c8d189, 32'hc2af2d8b, 32'hc27ee215, 32'hc18d632f, 32'h427639be, 32'h42a7d1fc, 32'h4291bdc6};
test_output[5696] = '{32'h42bce536};
test_index[5696] = '{0};
test_input[45576:45583] = '{32'hc284d456, 32'h40aa090b, 32'hc1aaffbb, 32'h42479db7, 32'h4214b658, 32'h404d69df, 32'h427d5eeb, 32'hc2464782};
test_output[5697] = '{32'h427d5eeb};
test_index[5697] = '{6};
test_input[45584:45591] = '{32'hc2890071, 32'hc275f39e, 32'hc156c8ff, 32'hc1840c78, 32'hc28afae0, 32'h41a4d511, 32'h4132f8a5, 32'hc1615454};
test_output[5698] = '{32'h41a4d511};
test_index[5698] = '{5};
test_input[45592:45599] = '{32'h41f86f93, 32'hc2986118, 32'hc135f409, 32'hc23f6c43, 32'h4291332c, 32'hc22f79ce, 32'hc1f882c1, 32'hc1410685};
test_output[5699] = '{32'h4291332c};
test_index[5699] = '{4};
test_input[45600:45607] = '{32'h421a8513, 32'h42a1f19e, 32'h427b0a6d, 32'h429832b1, 32'hc12db4f2, 32'h41983c2f, 32'h428f70f8, 32'hc20633bc};
test_output[5700] = '{32'h42a1f19e};
test_index[5700] = '{1};
test_input[45608:45615] = '{32'hc2bc5fca, 32'h418010d1, 32'hc1dcdb43, 32'hc24805d4, 32'hc2a792b6, 32'h424ca144, 32'hbfc5b245, 32'h42c1e667};
test_output[5701] = '{32'h42c1e667};
test_index[5701] = '{7};
test_input[45616:45623] = '{32'hc28dad8d, 32'h414b44ce, 32'hc274d3d7, 32'h401f5dba, 32'h42122af0, 32'hbf73801c, 32'hc2279ead, 32'h41b63b56};
test_output[5702] = '{32'h42122af0};
test_index[5702] = '{4};
test_input[45624:45631] = '{32'hc26caef8, 32'h40315486, 32'hc28eca07, 32'h424b58dc, 32'hc146d669, 32'hc16da556, 32'hc0f24999, 32'h42c0eeeb};
test_output[5703] = '{32'h42c0eeeb};
test_index[5703] = '{7};
test_input[45632:45639] = '{32'h426bc789, 32'hc2971401, 32'h42563662, 32'h429ba066, 32'hc2be4bf2, 32'h4191b6fe, 32'hc0fa8026, 32'hc01c19ae};
test_output[5704] = '{32'h429ba066};
test_index[5704] = '{3};
test_input[45640:45647] = '{32'h429139bb, 32'hbebfec5b, 32'hc281c878, 32'hc2b65fc1, 32'hc22c2f13, 32'h42c775aa, 32'h4285ebba, 32'h42b03573};
test_output[5705] = '{32'h42c775aa};
test_index[5705] = '{5};
test_input[45648:45655] = '{32'h428cd0c5, 32'hc16be6e4, 32'h423c7dd7, 32'h3f2e0d27, 32'hc1fdae3b, 32'hc1cb59e2, 32'h428a6710, 32'h425f47aa};
test_output[5706] = '{32'h428cd0c5};
test_index[5706] = '{0};
test_input[45656:45663] = '{32'h416200af, 32'h4298b87b, 32'hc2bfd8bb, 32'h4296735a, 32'h420a491b, 32'h41bdab5a, 32'h4276c9ec, 32'hc2a54fe0};
test_output[5707] = '{32'h4298b87b};
test_index[5707] = '{1};
test_input[45664:45671] = '{32'h421cdad7, 32'h41ffb1a5, 32'h41fbe745, 32'h419285c7, 32'hc20d8f3f, 32'h427ea9df, 32'h422d5799, 32'h41fb5e19};
test_output[5708] = '{32'h427ea9df};
test_index[5708] = '{5};
test_input[45672:45679] = '{32'h42ba298f, 32'h42419633, 32'hc2b1f3a7, 32'hc2ad5b8d, 32'hc27fb964, 32'hc26af229, 32'hc2954c19, 32'hc2954071};
test_output[5709] = '{32'h42ba298f};
test_index[5709] = '{0};
test_input[45680:45687] = '{32'hc1ec300d, 32'h423172a9, 32'h413bfd5a, 32'h427ee02a, 32'hc2775bc4, 32'h41af2715, 32'h4297fb0d, 32'h42afae73};
test_output[5710] = '{32'h42afae73};
test_index[5710] = '{7};
test_input[45688:45695] = '{32'hc2c64481, 32'hc2c550c2, 32'h428b7535, 32'h424215af, 32'hc22437f9, 32'hc2080c36, 32'h423183e0, 32'hc25818b6};
test_output[5711] = '{32'h428b7535};
test_index[5711] = '{2};
test_input[45696:45703] = '{32'h41e7d4c4, 32'h41be889d, 32'h42a25c94, 32'hc0389dc1, 32'hc1bdfd51, 32'hc2aa2ad7, 32'h42af172f, 32'h41e08703};
test_output[5712] = '{32'h42af172f};
test_index[5712] = '{6};
test_input[45704:45711] = '{32'h41a60dc7, 32'hbfb5b1fc, 32'h4195a135, 32'h422a5ad3, 32'hc2afeffa, 32'hc2bd277b, 32'hc1ec886e, 32'h420539c8};
test_output[5713] = '{32'h422a5ad3};
test_index[5713] = '{3};
test_input[45712:45719] = '{32'h40c970a4, 32'hc1f341b5, 32'hc1ee45ef, 32'h4281dedd, 32'hc2b47714, 32'hc2a69681, 32'hc16355e9, 32'hc2a57488};
test_output[5714] = '{32'h4281dedd};
test_index[5714] = '{3};
test_input[45720:45727] = '{32'hc2401360, 32'hc2b360c6, 32'hc23f63b2, 32'h425b77b3, 32'hc2554e69, 32'hc1a24021, 32'h412516e7, 32'hc2525119};
test_output[5715] = '{32'h425b77b3};
test_index[5715] = '{3};
test_input[45728:45735] = '{32'h42500292, 32'hc261c6ba, 32'h42aaf957, 32'h428bdcd9, 32'h4194353e, 32'h418b9da0, 32'hc24398c5, 32'hc234ac84};
test_output[5716] = '{32'h42aaf957};
test_index[5716] = '{2};
test_input[45736:45743] = '{32'h4285ade4, 32'hc290bbab, 32'h4247e0e6, 32'hc28d5ddb, 32'h42883586, 32'hc2a78b77, 32'hc1aa22ee, 32'hc25e59c7};
test_output[5717] = '{32'h42883586};
test_index[5717] = '{4};
test_input[45744:45751] = '{32'h42679e88, 32'hc2541713, 32'h41f98144, 32'h420d74d5, 32'hc2bdc8f0, 32'h420e746f, 32'h4043dc9c, 32'hc2afca39};
test_output[5718] = '{32'h42679e88};
test_index[5718] = '{0};
test_input[45752:45759] = '{32'hc205b1d2, 32'h4143c61b, 32'h420c17dc, 32'hc222ec1d, 32'hc0b0d23b, 32'h429ea354, 32'h42c5317f, 32'hc280f5d4};
test_output[5719] = '{32'h42c5317f};
test_index[5719] = '{6};
test_input[45760:45767] = '{32'hc291d21c, 32'h41a51a7a, 32'h40e59562, 32'hc24e5df7, 32'hc20d5ad8, 32'hc2ac95b8, 32'h4173d4f2, 32'hc29bbcfa};
test_output[5720] = '{32'h41a51a7a};
test_index[5720] = '{1};
test_input[45768:45775] = '{32'h421cdc5c, 32'hc209462f, 32'hc29bed67, 32'hc18500a4, 32'h425a43fb, 32'h422e23ef, 32'h4274e229, 32'hc2c602b5};
test_output[5721] = '{32'h4274e229};
test_index[5721] = '{6};
test_input[45776:45783] = '{32'h41a81d2e, 32'hc2bf8577, 32'hc2c28ecd, 32'h42ade68b, 32'h42a87393, 32'hc1de566d, 32'hc23ac5da, 32'h420e1399};
test_output[5722] = '{32'h42ade68b};
test_index[5722] = '{3};
test_input[45784:45791] = '{32'h42c1b15f, 32'h4237d72f, 32'hc24ee76a, 32'hc0ede810, 32'hc29c466f, 32'h42200207, 32'h42b99429, 32'hc236d2dd};
test_output[5723] = '{32'h42c1b15f};
test_index[5723] = '{0};
test_input[45792:45799] = '{32'h424f195d, 32'h419a453a, 32'hc2c7b8d3, 32'hc1cc3fe4, 32'h423d93ee, 32'h427ecadc, 32'hc2960644, 32'hc268357e};
test_output[5724] = '{32'h427ecadc};
test_index[5724] = '{5};
test_input[45800:45807] = '{32'hc1a2f964, 32'hbec3883e, 32'hc247ab69, 32'h41a08bd8, 32'h428c75a7, 32'h42794d37, 32'hc20f35eb, 32'hc180cfac};
test_output[5725] = '{32'h428c75a7};
test_index[5725] = '{4};
test_input[45808:45815] = '{32'hc28441b2, 32'h41cc133c, 32'hc28654ea, 32'h40d30ffd, 32'h41e2487e, 32'h426191d5, 32'h427b9f5c, 32'h419d0f77};
test_output[5726] = '{32'h427b9f5c};
test_index[5726] = '{6};
test_input[45816:45823] = '{32'hc16fc014, 32'hc23e242b, 32'hc25c384c, 32'h4254b323, 32'hc2579d2e, 32'hc24a6287, 32'h418226ce, 32'hc21d7395};
test_output[5727] = '{32'h4254b323};
test_index[5727] = '{3};
test_input[45824:45831] = '{32'h40c25040, 32'hbe65b2fd, 32'h41392a1d, 32'hc29f82fd, 32'h420b439d, 32'h41d99ea8, 32'h415ae079, 32'h42b4cef4};
test_output[5728] = '{32'h42b4cef4};
test_index[5728] = '{7};
test_input[45832:45839] = '{32'hc275f47b, 32'hc197b667, 32'hc0f55902, 32'hc1b9d145, 32'hc1a0f477, 32'hc29322be, 32'h4236cb5b, 32'h423745f2};
test_output[5729] = '{32'h423745f2};
test_index[5729] = '{7};
test_input[45840:45847] = '{32'hc29efafb, 32'h421d1ead, 32'h41c07271, 32'hc2b72ccb, 32'hc166570e, 32'hc2bfc200, 32'h4124030e, 32'hc22af184};
test_output[5730] = '{32'h421d1ead};
test_index[5730] = '{1};
test_input[45848:45855] = '{32'h42014f84, 32'hc1dd3dc1, 32'h42adf163, 32'h428f57da, 32'hc0e8f540, 32'h41e43808, 32'hc1a587e1, 32'hc29cdb3d};
test_output[5731] = '{32'h42adf163};
test_index[5731] = '{2};
test_input[45856:45863] = '{32'hc2980a77, 32'hc2308e7f, 32'h42a31c1e, 32'h41a9b5fa, 32'hc2b3549b, 32'h424e9eb7, 32'h42944bf6, 32'h4103b158};
test_output[5732] = '{32'h42a31c1e};
test_index[5732] = '{2};
test_input[45864:45871] = '{32'hc1c356cc, 32'h429312af, 32'hc2c3edf7, 32'hc246f06a, 32'h411c4fac, 32'hc2907907, 32'h4249155d, 32'h42288dba};
test_output[5733] = '{32'h429312af};
test_index[5733] = '{1};
test_input[45872:45879] = '{32'h41a73db8, 32'h42a5e2e2, 32'h41fec463, 32'h3e566d7e, 32'hc2311c6c, 32'h42541db7, 32'h42aef93e, 32'h42626a55};
test_output[5734] = '{32'h42aef93e};
test_index[5734] = '{6};
test_input[45880:45887] = '{32'hc23cf577, 32'h424728c0, 32'hc2a75e7f, 32'hc2b36f73, 32'h428a384e, 32'hc2b34413, 32'h42a26949, 32'h4206ca4f};
test_output[5735] = '{32'h42a26949};
test_index[5735] = '{6};
test_input[45888:45895] = '{32'h426f1b67, 32'hc28b9645, 32'hc209ecb6, 32'h42ac9b66, 32'hc0903696, 32'hc121d1c2, 32'hc1d92a37, 32'h4240d091};
test_output[5736] = '{32'h42ac9b66};
test_index[5736] = '{3};
test_input[45896:45903] = '{32'h407d785c, 32'hc215c3ce, 32'hc2c4d601, 32'hc22399ca, 32'h429b5bab, 32'h429fc0bc, 32'h404a3f61, 32'h42abe79d};
test_output[5737] = '{32'h42abe79d};
test_index[5737] = '{7};
test_input[45904:45911] = '{32'hc292c9b8, 32'h42a44573, 32'h424a1fbc, 32'hc2bac7ad, 32'h411b6c8b, 32'hc1317178, 32'h41c01b53, 32'h41b8afa6};
test_output[5738] = '{32'h42a44573};
test_index[5738] = '{1};
test_input[45912:45919] = '{32'h4276c710, 32'hc1024947, 32'h40dad02c, 32'h42424052, 32'h4220b99c, 32'h423095ec, 32'h42c6ffb9, 32'hc228688f};
test_output[5739] = '{32'h42c6ffb9};
test_index[5739] = '{6};
test_input[45920:45927] = '{32'h40cec54b, 32'h428787c7, 32'h42961bed, 32'hc1208a99, 32'h41658709, 32'h420d4e2c, 32'h42037fa0, 32'h421b418a};
test_output[5740] = '{32'h42961bed};
test_index[5740] = '{2};
test_input[45928:45935] = '{32'h4225eaa5, 32'hc2205b14, 32'h42845e61, 32'h41cc9a56, 32'h410cf3dc, 32'hc1a6943c, 32'h41ec1c3f, 32'hc1e3f98d};
test_output[5741] = '{32'h42845e61};
test_index[5741] = '{2};
test_input[45936:45943] = '{32'hc1847746, 32'hc28c157e, 32'h42285406, 32'hc18659c7, 32'hc2c5a92d, 32'h40737973, 32'h41198556, 32'h42b46bb4};
test_output[5742] = '{32'h42b46bb4};
test_index[5742] = '{7};
test_input[45944:45951] = '{32'h4184f03c, 32'h4296a60f, 32'h42c77134, 32'hc2a039a0, 32'hc121b4e6, 32'hc1d31139, 32'h429dd193, 32'h41554a5b};
test_output[5743] = '{32'h42c77134};
test_index[5743] = '{2};
test_input[45952:45959] = '{32'h41a78c45, 32'h41b28963, 32'hc282eb40, 32'hc293bf82, 32'hc0e139ae, 32'h427a13e2, 32'h4181f287, 32'h41ad89a7};
test_output[5744] = '{32'h427a13e2};
test_index[5744] = '{5};
test_input[45960:45967] = '{32'h414bc887, 32'h429cc01b, 32'hc16b9959, 32'hc217cf8f, 32'hc29125e1, 32'hc26b0954, 32'h428fbddb, 32'h426efa3b};
test_output[5745] = '{32'h429cc01b};
test_index[5745] = '{1};
test_input[45968:45975] = '{32'hc218e671, 32'h41ef6346, 32'hc28dadd7, 32'hc1b696d2, 32'h41cede70, 32'hc2a53aac, 32'hc28d03e2, 32'hc23160f1};
test_output[5746] = '{32'h41ef6346};
test_index[5746] = '{1};
test_input[45976:45983] = '{32'h4101379b, 32'hc28dead4, 32'hc155fa34, 32'h42a1fe4f, 32'h42810b38, 32'hc148ac04, 32'h42a6b67d, 32'h42018d03};
test_output[5747] = '{32'h42a6b67d};
test_index[5747] = '{6};
test_input[45984:45991] = '{32'h3f1bcbbb, 32'hc28c9d02, 32'h417bd81f, 32'hc249e611, 32'h42a8f855, 32'hc1f250d4, 32'h42489ed8, 32'hc2a14c63};
test_output[5748] = '{32'h42a8f855};
test_index[5748] = '{4};
test_input[45992:45999] = '{32'hc2c4ee51, 32'hbff23b63, 32'h4208246e, 32'hc2150009, 32'hc245a079, 32'h429a0dab, 32'hc148384f, 32'hc230de64};
test_output[5749] = '{32'h429a0dab};
test_index[5749] = '{5};
test_input[46000:46007] = '{32'hc233b4f0, 32'hc23a3128, 32'h42377870, 32'h4268011a, 32'hc1d6523b, 32'h42bb69de, 32'h42934b46, 32'hc280bbd5};
test_output[5750] = '{32'h42bb69de};
test_index[5750] = '{5};
test_input[46008:46015] = '{32'hc2a0640f, 32'h41cc2575, 32'hc2118cb8, 32'h42bdd56d, 32'h41e0f95e, 32'hc2c7beff, 32'hc2ab59b6, 32'h42972164};
test_output[5751] = '{32'h42bdd56d};
test_index[5751] = '{3};
test_input[46016:46023] = '{32'h42ad0ee8, 32'hc29f25b3, 32'hc22fdbc2, 32'hc265b467, 32'h42c2ebd5, 32'hc25e8f01, 32'h42867777, 32'h429f4921};
test_output[5752] = '{32'h42c2ebd5};
test_index[5752] = '{4};
test_input[46024:46031] = '{32'hc10c9a2f, 32'h422f17c2, 32'hc26c1b06, 32'hc1e3cd4a, 32'hc222c836, 32'h4184fb77, 32'hc23c6054, 32'hc2c2e051};
test_output[5753] = '{32'h422f17c2};
test_index[5753] = '{1};
test_input[46032:46039] = '{32'h41fd3ea1, 32'h424af500, 32'hc1f661ad, 32'hc28d6b33, 32'h423f502f, 32'h42c2849b, 32'hc24f125d, 32'hc0def037};
test_output[5754] = '{32'h42c2849b};
test_index[5754] = '{5};
test_input[46040:46047] = '{32'h42703b55, 32'h4275b305, 32'hc2b29cdf, 32'hc21ea68d, 32'hc1b4b871, 32'hc2b2d480, 32'h42513281, 32'hc2068bbf};
test_output[5755] = '{32'h4275b305};
test_index[5755] = '{1};
test_input[46048:46055] = '{32'h42ae7457, 32'hc2b3da59, 32'hc28c0b88, 32'h429c51fc, 32'hc13fe12c, 32'hc0407c9d, 32'h3f2f96cd, 32'h424145ed};
test_output[5756] = '{32'h42ae7457};
test_index[5756] = '{0};
test_input[46056:46063] = '{32'h429dc54d, 32'hc1d48e93, 32'hc24939c4, 32'hc1dbe605, 32'h41bcf2f2, 32'hc191ce0f, 32'h427c992f, 32'hc29357bb};
test_output[5757] = '{32'h429dc54d};
test_index[5757] = '{0};
test_input[46064:46071] = '{32'hc1ad36fa, 32'hc2b6abc1, 32'hc2758c62, 32'h4265d594, 32'h3ff30d27, 32'h42aa2406, 32'h41e1b7c3, 32'h42a53682};
test_output[5758] = '{32'h42aa2406};
test_index[5758] = '{5};
test_input[46072:46079] = '{32'hc1d6c6c1, 32'h42947191, 32'hc05d6d6e, 32'hc1e841f6, 32'h41afd443, 32'h4117d3b0, 32'h428b4dc3, 32'h42a363b9};
test_output[5759] = '{32'h42a363b9};
test_index[5759] = '{7};
test_input[46080:46087] = '{32'h426b6c56, 32'hc2c13811, 32'hc1b9ffad, 32'h41de3464, 32'h42022339, 32'hc1771f02, 32'h40ed627f, 32'hc292a875};
test_output[5760] = '{32'h426b6c56};
test_index[5760] = '{0};
test_input[46088:46095] = '{32'h42bca1b5, 32'h4248a1a9, 32'hc07e1b9c, 32'h4255b47e, 32'h4153b8b3, 32'h428dfc1d, 32'hc1ee2412, 32'hc1838712};
test_output[5761] = '{32'h42bca1b5};
test_index[5761] = '{0};
test_input[46096:46103] = '{32'hc1dd0cff, 32'hc2914a32, 32'hc09569f4, 32'h426b5a1c, 32'h42887319, 32'h41c2411e, 32'hc26b6b7c, 32'h41b26896};
test_output[5762] = '{32'h42887319};
test_index[5762] = '{4};
test_input[46104:46111] = '{32'h410b845f, 32'h4291f8af, 32'hc2954601, 32'h422251a5, 32'h41a3090c, 32'hc2499f59, 32'h421727ce, 32'hc23312a2};
test_output[5763] = '{32'h4291f8af};
test_index[5763] = '{1};
test_input[46112:46119] = '{32'hc2c502e2, 32'h42a35edc, 32'hc2c09166, 32'hc1dc500f, 32'hc22d6242, 32'h42710f9d, 32'hc25bed0a, 32'hc259f0ed};
test_output[5764] = '{32'h42a35edc};
test_index[5764] = '{1};
test_input[46120:46127] = '{32'h4214987a, 32'hc14cf036, 32'h428ac397, 32'h420a190e, 32'h42af3e30, 32'h4135e80e, 32'h429ac255, 32'hc28886fa};
test_output[5765] = '{32'h42af3e30};
test_index[5765] = '{4};
test_input[46128:46135] = '{32'hc09f9387, 32'h428521ff, 32'h424b029e, 32'hc16dba9e, 32'h4258eb88, 32'h419de0c4, 32'hc21907c5, 32'hc2709fd2};
test_output[5766] = '{32'h428521ff};
test_index[5766] = '{1};
test_input[46136:46143] = '{32'hc2b8901a, 32'hc2038e04, 32'hc2877978, 32'hc27b4fc1, 32'hc1cc9b70, 32'hc1cb7e55, 32'h3f19302f, 32'hc2a484c4};
test_output[5767] = '{32'h3f19302f};
test_index[5767] = '{6};
test_input[46144:46151] = '{32'h4281f7ad, 32'hc1fd1f52, 32'hc2acc46f, 32'hc2028dae, 32'hc27dbbf8, 32'hc26168e9, 32'hc29dd919, 32'hc1d86db4};
test_output[5768] = '{32'h4281f7ad};
test_index[5768] = '{0};
test_input[46152:46159] = '{32'h419c74dd, 32'h42c225dd, 32'h426e8b68, 32'h42121b5f, 32'hc2a33138, 32'hc175c8ab, 32'hc29d0351, 32'h4230c970};
test_output[5769] = '{32'h42c225dd};
test_index[5769] = '{1};
test_input[46160:46167] = '{32'h427635a9, 32'hc1614d92, 32'hc1e8f3ea, 32'h42c1abd2, 32'hc2b659c4, 32'hc13e703d, 32'h41f22bf3, 32'hc1ea98ca};
test_output[5770] = '{32'h42c1abd2};
test_index[5770] = '{3};
test_input[46168:46175] = '{32'hc2033431, 32'hc2adc583, 32'h42816b52, 32'h427e4612, 32'hc23f4134, 32'h42be3401, 32'hc25062d3, 32'hc27b9794};
test_output[5771] = '{32'h42be3401};
test_index[5771] = '{5};
test_input[46176:46183] = '{32'h42882b66, 32'h427eb131, 32'h4280eb80, 32'hc2a7c0a7, 32'hc188de7c, 32'h425bd251, 32'hc1fe823c, 32'hc2977765};
test_output[5772] = '{32'h42882b66};
test_index[5772] = '{0};
test_input[46184:46191] = '{32'h427990e3, 32'h42a6e579, 32'h42963ac2, 32'h42c30994, 32'h42a70463, 32'h410cbd75, 32'hc108ab11, 32'hc1a86b54};
test_output[5773] = '{32'h42c30994};
test_index[5773] = '{3};
test_input[46192:46199] = '{32'h42854c17, 32'hc2a9a755, 32'hc2731192, 32'h42c4c42d, 32'hbefdd1e1, 32'h420baea7, 32'h42953033, 32'h42c66d64};
test_output[5774] = '{32'h42c66d64};
test_index[5774] = '{7};
test_input[46200:46207] = '{32'h42312f5f, 32'hc1218353, 32'h424eb20e, 32'hc2475ef6, 32'hc0760da7, 32'h42304210, 32'h423bd8a7, 32'h40efc232};
test_output[5775] = '{32'h424eb20e};
test_index[5775] = '{2};
test_input[46208:46215] = '{32'h412c6c6e, 32'h424fc2a3, 32'hc18c7f8e, 32'hc1528d31, 32'hc2ac07d2, 32'hc1726544, 32'h42c3d53d, 32'h4282b33f};
test_output[5776] = '{32'h42c3d53d};
test_index[5776] = '{6};
test_input[46216:46223] = '{32'hc229a20a, 32'hc2072406, 32'h4109a93f, 32'hc289fc59, 32'hc11a48f0, 32'h428824f3, 32'h41adfc00, 32'h42b9ae07};
test_output[5777] = '{32'h42b9ae07};
test_index[5777] = '{7};
test_input[46224:46231] = '{32'h42c211de, 32'hc286a417, 32'hc27b19a0, 32'h4227c242, 32'hc2acd3bc, 32'h428e1a5a, 32'h4278b4d1, 32'h4239c8cd};
test_output[5778] = '{32'h42c211de};
test_index[5778] = '{0};
test_input[46232:46239] = '{32'h42bc4eda, 32'h42944636, 32'hc18df0d0, 32'hc27a319a, 32'hc1153bc6, 32'hc28e38fc, 32'h42c1f4a4, 32'hc0a98bd9};
test_output[5779] = '{32'h42c1f4a4};
test_index[5779] = '{6};
test_input[46240:46247] = '{32'hc2446416, 32'h418900e2, 32'hc1d9b51b, 32'hc2b0a6ac, 32'h419c1e95, 32'h40eec922, 32'h422bb438, 32'hc1cb1d01};
test_output[5780] = '{32'h422bb438};
test_index[5780] = '{6};
test_input[46248:46255] = '{32'hc2a7347e, 32'hc29571fc, 32'h42668e33, 32'h426f7e15, 32'hc0a2bf7e, 32'h4275ab41, 32'hc1f284a2, 32'hc20fe340};
test_output[5781] = '{32'h4275ab41};
test_index[5781] = '{5};
test_input[46256:46263] = '{32'hc2a52401, 32'h42b39b54, 32'h3ff49938, 32'hc28d9f1c, 32'h41a9da2b, 32'h425d7740, 32'h42bc76de, 32'h42728e95};
test_output[5782] = '{32'h42bc76de};
test_index[5782] = '{6};
test_input[46264:46271] = '{32'hc2c63f49, 32'hc287755b, 32'h42966094, 32'h4288fa3f, 32'h42636d15, 32'h41fe85d2, 32'hc287bd72, 32'hc2b307a6};
test_output[5783] = '{32'h42966094};
test_index[5783] = '{2};
test_input[46272:46279] = '{32'hc1ec3178, 32'h424cb49a, 32'hc2af5409, 32'hc2272f8b, 32'hc2aa5673, 32'h42bde16f, 32'hc28cc9e6, 32'h40a689c5};
test_output[5784] = '{32'h42bde16f};
test_index[5784] = '{5};
test_input[46280:46287] = '{32'h41c32a3e, 32'h429a6232, 32'hc2ab62bf, 32'hc2482155, 32'h42bb20fe, 32'hc285cfef, 32'h42c1877c, 32'h407d8e2e};
test_output[5785] = '{32'h42c1877c};
test_index[5785] = '{6};
test_input[46288:46295] = '{32'hc273f372, 32'hc1145c70, 32'h423c0ca4, 32'hc2a10369, 32'h4222f54f, 32'h429dc90a, 32'hc1a571bd, 32'h4282f90f};
test_output[5786] = '{32'h429dc90a};
test_index[5786] = '{5};
test_input[46296:46303] = '{32'h4247821a, 32'h42bceeac, 32'hc2a49e23, 32'hc236bcfe, 32'h42235f9d, 32'hc2a9ee34, 32'h429b3274, 32'h41576908};
test_output[5787] = '{32'h42bceeac};
test_index[5787] = '{1};
test_input[46304:46311] = '{32'h42678e58, 32'hc20d7713, 32'hc1112ffe, 32'hc17999ad, 32'hc08b426a, 32'h4286d271, 32'h42bee94e, 32'hc202154a};
test_output[5788] = '{32'h42bee94e};
test_index[5788] = '{6};
test_input[46312:46319] = '{32'h4246b56c, 32'hc2c11c51, 32'h41eed722, 32'hc13fc27a, 32'hc195df47, 32'hc193c8ed, 32'hc2813c9a, 32'hc2b57889};
test_output[5789] = '{32'h4246b56c};
test_index[5789] = '{0};
test_input[46320:46327] = '{32'hc218d085, 32'hc28f45c3, 32'h4241de3a, 32'hc21ad645, 32'h4299b69b, 32'h420bb0fc, 32'h41f4f378, 32'hc2492799};
test_output[5790] = '{32'h4299b69b};
test_index[5790] = '{4};
test_input[46328:46335] = '{32'h4202383a, 32'h421c67bf, 32'hc2a8550e, 32'hc28c11f1, 32'h42c74de2, 32'hc2233d38, 32'h421f8ee7, 32'h40874330};
test_output[5791] = '{32'h42c74de2};
test_index[5791] = '{4};
test_input[46336:46343] = '{32'hc2c6c261, 32'hc22d5f78, 32'hc2abb07d, 32'h424b8c64, 32'hc1f14a41, 32'hc2bc8ec7, 32'h41516b91, 32'h420be715};
test_output[5792] = '{32'h424b8c64};
test_index[5792] = '{3};
test_input[46344:46351] = '{32'hc1bb86c1, 32'hc2ae67ce, 32'h42a3ae11, 32'h429f9848, 32'hc2b56375, 32'h428686b7, 32'h428ecd39, 32'h421d18bc};
test_output[5793] = '{32'h42a3ae11};
test_index[5793] = '{2};
test_input[46352:46359] = '{32'hc28a6bc5, 32'hc2b3fd42, 32'hc2ae5dc1, 32'hc2aa18e0, 32'h42c06401, 32'h42c1a54b, 32'h40ac42ca, 32'hc2bdfeaf};
test_output[5794] = '{32'h42c1a54b};
test_index[5794] = '{5};
test_input[46360:46367] = '{32'h421a4e8f, 32'h424e49e5, 32'hc2a0e80c, 32'h426626ef, 32'h425c16f1, 32'hc1b67844, 32'hc29e618e, 32'hc2502200};
test_output[5795] = '{32'h426626ef};
test_index[5795] = '{3};
test_input[46368:46375] = '{32'hc2804da5, 32'hc26957e2, 32'hc26a2e79, 32'hc27091ad, 32'h42ad47cf, 32'h42aa3712, 32'h42074447, 32'hc0fe02fb};
test_output[5796] = '{32'h42ad47cf};
test_index[5796] = '{4};
test_input[46376:46383] = '{32'h415464b9, 32'hc27e9d67, 32'h422229bc, 32'h40a31b9e, 32'hc054b920, 32'h4163b9e5, 32'hc281e34f, 32'hc02dc989};
test_output[5797] = '{32'h422229bc};
test_index[5797] = '{2};
test_input[46384:46391] = '{32'h4229918c, 32'hc29257fc, 32'hc2b4720e, 32'hc1fd2c4c, 32'hc1eddc86, 32'h41a868fc, 32'hc259a8f8, 32'h42339349};
test_output[5798] = '{32'h42339349};
test_index[5798] = '{7};
test_input[46392:46399] = '{32'hc25ae73d, 32'hc288769c, 32'h42a0e651, 32'hc0f65417, 32'h423c5577, 32'h4237c1e6, 32'hc171b277, 32'h42870e8f};
test_output[5799] = '{32'h42a0e651};
test_index[5799] = '{2};
test_input[46400:46407] = '{32'hc20db44b, 32'h42a556a3, 32'hc2aafd22, 32'hc27ab932, 32'h411236a3, 32'hc203f33a, 32'hc1a7587a, 32'h41e0ff0e};
test_output[5800] = '{32'h42a556a3};
test_index[5800] = '{1};
test_input[46408:46415] = '{32'h42926ba3, 32'hbeb71d52, 32'hc1d41588, 32'hc0f9f3b7, 32'hc286b202, 32'hc15a0eae, 32'hc234b41f, 32'h4212ef5d};
test_output[5801] = '{32'h42926ba3};
test_index[5801] = '{0};
test_input[46416:46423] = '{32'h41ac339d, 32'hc26749b9, 32'hc150934f, 32'h41b16a3a, 32'h425c560b, 32'h42c61377, 32'hc1f0e90a, 32'h425e87fa};
test_output[5802] = '{32'h42c61377};
test_index[5802] = '{5};
test_input[46424:46431] = '{32'h4274a97c, 32'hc210d67a, 32'h4296ce79, 32'hc2556916, 32'hc0e18060, 32'h429966e8, 32'hc233e93d, 32'h428a29a9};
test_output[5803] = '{32'h429966e8};
test_index[5803] = '{5};
test_input[46432:46439] = '{32'hc241bfbe, 32'h404ba1c7, 32'h428a94e5, 32'h4129d654, 32'hc171c95f, 32'h428bbcea, 32'hc2b603c1, 32'h418bd232};
test_output[5804] = '{32'h428bbcea};
test_index[5804] = '{5};
test_input[46440:46447] = '{32'hc1c9c4de, 32'hc2153ea9, 32'h425624e0, 32'h41515ed8, 32'h422ee1da, 32'h40922741, 32'h4138b91c, 32'h420bb9fc};
test_output[5805] = '{32'h425624e0};
test_index[5805] = '{2};
test_input[46448:46455] = '{32'hc119e786, 32'h413e6979, 32'hc2877abb, 32'hbdad8e75, 32'h42bd2496, 32'hc28e3bf2, 32'hc2411c79, 32'h426eaec6};
test_output[5806] = '{32'h42bd2496};
test_index[5806] = '{4};
test_input[46456:46463] = '{32'h4179776c, 32'h40bb2e3f, 32'h42947bc7, 32'h42698cfd, 32'hbea1621a, 32'h40cd6cb2, 32'hc2022105, 32'hc220ae11};
test_output[5807] = '{32'h42947bc7};
test_index[5807] = '{2};
test_input[46464:46471] = '{32'hc27a7e11, 32'hc298d9c3, 32'hc2b05f99, 32'hc29575aa, 32'h4126933d, 32'hc155f3d1, 32'hc28afaa7, 32'h4247c54e};
test_output[5808] = '{32'h4247c54e};
test_index[5808] = '{7};
test_input[46472:46479] = '{32'h42a8931d, 32'h425f976d, 32'h42c585bd, 32'hc2400309, 32'hc2907909, 32'hc1ad2148, 32'h429bce69, 32'h42100f6e};
test_output[5809] = '{32'h42c585bd};
test_index[5809] = '{2};
test_input[46480:46487] = '{32'hc1f4d47f, 32'hc1cc875b, 32'h413b89d4, 32'hc2c4aadb, 32'h42997546, 32'h42342559, 32'hc2a85c82, 32'h425ecd8b};
test_output[5810] = '{32'h42997546};
test_index[5810] = '{4};
test_input[46488:46495] = '{32'h42a7ac89, 32'hc1c569c2, 32'hc23c7f77, 32'h42a763a4, 32'h41de1034, 32'hc228fca5, 32'h4258435f, 32'hc26030bd};
test_output[5811] = '{32'h42a7ac89};
test_index[5811] = '{0};
test_input[46496:46503] = '{32'hc2a85f7a, 32'h413e31e6, 32'h40ebedc7, 32'h42052da0, 32'h425eb0ef, 32'hc2b6d6eb, 32'h419ab2a6, 32'hc2a07549};
test_output[5812] = '{32'h425eb0ef};
test_index[5812] = '{4};
test_input[46504:46511] = '{32'hc183724b, 32'hc190c3e0, 32'h426e20f8, 32'h42b2b66c, 32'h42b7351a, 32'h42659fc3, 32'hc2ac450c, 32'hc1502ad1};
test_output[5813] = '{32'h42b7351a};
test_index[5813] = '{4};
test_input[46512:46519] = '{32'hc29908be, 32'hc2a12992, 32'h429366ef, 32'h419c8dad, 32'hc103b458, 32'hc113a7e5, 32'hc261f374, 32'h42720e57};
test_output[5814] = '{32'h429366ef};
test_index[5814] = '{2};
test_input[46520:46527] = '{32'h428b7ad5, 32'hc17ecce0, 32'hc2a64e35, 32'hc2b5c08c, 32'h419cf89f, 32'h42ae5f40, 32'hc13a226b, 32'hc2849c80};
test_output[5815] = '{32'h42ae5f40};
test_index[5815] = '{5};
test_input[46528:46535] = '{32'hc2c6c962, 32'h42c5db4a, 32'h415a5dea, 32'h424c736c, 32'hc24fe014, 32'h42be6a8b, 32'hbf475fa9, 32'hc2551719};
test_output[5816] = '{32'h42c5db4a};
test_index[5816] = '{1};
test_input[46536:46543] = '{32'h42195c6e, 32'hc266e19a, 32'hc24a6b58, 32'h426027f2, 32'h41ae92f8, 32'hc1999216, 32'h417459de, 32'h42682f44};
test_output[5817] = '{32'h42682f44};
test_index[5817] = '{7};
test_input[46544:46551] = '{32'h426413d5, 32'h42803480, 32'h42b9ddf5, 32'hc2a560a9, 32'hc2aa9a95, 32'hc294650e, 32'h4289f36c, 32'h405f3392};
test_output[5818] = '{32'h42b9ddf5};
test_index[5818] = '{2};
test_input[46552:46559] = '{32'h42b92964, 32'hc2842869, 32'h40b94452, 32'hc2129fa4, 32'h3f561cd6, 32'h4275b909, 32'hc05e6982, 32'h413ccfa8};
test_output[5819] = '{32'h42b92964};
test_index[5819] = '{0};
test_input[46560:46567] = '{32'h42a81972, 32'hc2532ab7, 32'hc2355415, 32'hc2357a4d, 32'h42597cc4, 32'hc1f9ea59, 32'hc10b956e, 32'h3ef6c698};
test_output[5820] = '{32'h42a81972};
test_index[5820] = '{0};
test_input[46568:46575] = '{32'hc2c37150, 32'hc2b40026, 32'h42bb88d7, 32'hc27fa71f, 32'hc29998a4, 32'hc050e6bf, 32'hc1d0e6d7, 32'hc23297cc};
test_output[5821] = '{32'h42bb88d7};
test_index[5821] = '{2};
test_input[46576:46583] = '{32'hc20fc9e7, 32'h41172961, 32'hc0c91071, 32'hc2bd16c3, 32'hc2b1ba6d, 32'hc237eb2a, 32'hc2880421, 32'h419630a8};
test_output[5822] = '{32'h419630a8};
test_index[5822] = '{7};
test_input[46584:46591] = '{32'hc237e4b0, 32'hc27bc88a, 32'hc23855d5, 32'hc2a3bd63, 32'h42c4e330, 32'hc220d4af, 32'hc20cb53f, 32'h41d3bdd0};
test_output[5823] = '{32'h42c4e330};
test_index[5823] = '{4};
test_input[46592:46599] = '{32'h42016d4e, 32'h41dcaef9, 32'h421196c8, 32'hc2c057ca, 32'hc26386e8, 32'hc28e625f, 32'h3f967641, 32'hc21a2cef};
test_output[5824] = '{32'h421196c8};
test_index[5824] = '{2};
test_input[46600:46607] = '{32'hc23171ce, 32'hc1e8540d, 32'hc24cdcf7, 32'h42781dcf, 32'h41f3e0d9, 32'h42a01271, 32'hc2acf191, 32'hc264083a};
test_output[5825] = '{32'h42a01271};
test_index[5825] = '{5};
test_input[46608:46615] = '{32'hc2b7ccad, 32'h4299c20b, 32'h42708656, 32'h42291ecc, 32'hc18a2655, 32'h423cd422, 32'hc2610667, 32'h4172f3f9};
test_output[5826] = '{32'h4299c20b};
test_index[5826] = '{1};
test_input[46616:46623] = '{32'hc1c1dcf6, 32'hc2a6ded3, 32'h41a560ce, 32'h42a136d4, 32'hc2c0f7dd, 32'h42bb2edb, 32'h41deed04, 32'hc2c2bde9};
test_output[5827] = '{32'h42bb2edb};
test_index[5827] = '{5};
test_input[46624:46631] = '{32'hc0dc1021, 32'hc2479a96, 32'h40ca6bd8, 32'h426de2dd, 32'hc0583461, 32'h428be64c, 32'h424ece58, 32'h4284e014};
test_output[5828] = '{32'h428be64c};
test_index[5828] = '{5};
test_input[46632:46639] = '{32'hc18de18f, 32'h414aa316, 32'hc27099cb, 32'hc2a906ae, 32'h40edd15d, 32'hc2812d38, 32'h42947be3, 32'h4248f0e4};
test_output[5829] = '{32'h42947be3};
test_index[5829] = '{6};
test_input[46640:46647] = '{32'h41f51631, 32'hc291389c, 32'hc2857ea7, 32'hc2a56dae, 32'hc151c007, 32'hc2140210, 32'h41f89ec8, 32'h409e852f};
test_output[5830] = '{32'h41f89ec8};
test_index[5830] = '{6};
test_input[46648:46655] = '{32'h41c022df, 32'h3d8a6d84, 32'h42041560, 32'h419dfd73, 32'h42a1644b, 32'hc1c8e5a5, 32'hc1cce3c3, 32'hc2b10277};
test_output[5831] = '{32'h42a1644b};
test_index[5831] = '{4};
test_input[46656:46663] = '{32'h4292d685, 32'h42c30d61, 32'hc0a7214f, 32'h42a29488, 32'hc0da7fb8, 32'hc26955ef, 32'h41eef472, 32'h42769caf};
test_output[5832] = '{32'h42c30d61};
test_index[5832] = '{1};
test_input[46664:46671] = '{32'hc287181d, 32'h425793c4, 32'h4218f49d, 32'hc25078d9, 32'h41a4e41f, 32'hc267fc01, 32'h42ad10f1, 32'hc2a68dbc};
test_output[5833] = '{32'h42ad10f1};
test_index[5833] = '{6};
test_input[46672:46679] = '{32'h42403521, 32'hc295245b, 32'hc290ed94, 32'h42983977, 32'hc24113c1, 32'h42b723c3, 32'hc20fbcdb, 32'hc2a1f2cc};
test_output[5834] = '{32'h42b723c3};
test_index[5834] = '{5};
test_input[46680:46687] = '{32'h405203e2, 32'hc2a9ddb7, 32'h42675476, 32'h420eb047, 32'h426bd40c, 32'hc0c0787f, 32'hc24b7596, 32'hc1f75f0d};
test_output[5835] = '{32'h426bd40c};
test_index[5835] = '{4};
test_input[46688:46695] = '{32'h3fa801fd, 32'hc2aacd1d, 32'hc2a78cdf, 32'hc205e626, 32'h42b12ce6, 32'h41a0f6a0, 32'h421c63bf, 32'h415496bb};
test_output[5836] = '{32'h42b12ce6};
test_index[5836] = '{4};
test_input[46696:46703] = '{32'hc22afc4e, 32'hc26b2e77, 32'hc2290803, 32'hc0d5990f, 32'hc1033500, 32'h427e4be5, 32'hc296c19c, 32'h4252394d};
test_output[5837] = '{32'h427e4be5};
test_index[5837] = '{5};
test_input[46704:46711] = '{32'h40cd5aa3, 32'h4287f408, 32'hc28a28f0, 32'hc253a566, 32'h42550f2a, 32'hc26b906c, 32'h4195ac53, 32'hc2ba904b};
test_output[5838] = '{32'h4287f408};
test_index[5838] = '{1};
test_input[46712:46719] = '{32'hc22764ed, 32'h421d381f, 32'h42604e4a, 32'h4146981a, 32'hc231f8af, 32'hc28cf0ef, 32'hc237ed1a, 32'hc2216bd4};
test_output[5839] = '{32'h42604e4a};
test_index[5839] = '{2};
test_input[46720:46727] = '{32'hc10d9183, 32'hc0e314fc, 32'h41d39ed0, 32'hc223e061, 32'hc2abfc28, 32'hc250a3a8, 32'h422d30ed, 32'hc2524dd2};
test_output[5840] = '{32'h422d30ed};
test_index[5840] = '{6};
test_input[46728:46735] = '{32'hc2c75cc1, 32'hc27fa118, 32'hc2ac4308, 32'hc197731c, 32'h41ef8887, 32'h3ec645ba, 32'h4210d4da, 32'h422c0fb0};
test_output[5841] = '{32'h422c0fb0};
test_index[5841] = '{7};
test_input[46736:46743] = '{32'h42a0498f, 32'h42b40a49, 32'h42709e15, 32'h42c5eff1, 32'hc1ca81d3, 32'hc2c03313, 32'h42a74ce0, 32'hc239d5d7};
test_output[5842] = '{32'h42c5eff1};
test_index[5842] = '{3};
test_input[46744:46751] = '{32'h423f4e3a, 32'hc2b50624, 32'hc2492439, 32'h42a1fa5e, 32'hc23e2f17, 32'h42808d6b, 32'hc1520fdd, 32'hc24e2224};
test_output[5843] = '{32'h42a1fa5e};
test_index[5843] = '{3};
test_input[46752:46759] = '{32'hc229459a, 32'h428e0de6, 32'h428c8cee, 32'h429af3e9, 32'h426dac34, 32'h423ff8b9, 32'h42874189, 32'hc178e8e0};
test_output[5844] = '{32'h429af3e9};
test_index[5844] = '{3};
test_input[46760:46767] = '{32'h4188e5aa, 32'hc2a4c55f, 32'hc08cd092, 32'hc2a4573c, 32'h3fd41ad4, 32'h41890d43, 32'h419b7a33, 32'hc1ddd977};
test_output[5845] = '{32'h419b7a33};
test_index[5845] = '{6};
test_input[46768:46775] = '{32'hc299bf0e, 32'h42727bc4, 32'h424e74ab, 32'hc21ed5e8, 32'hc2578989, 32'hc1a5edd2, 32'h4257564e, 32'h41ca4943};
test_output[5846] = '{32'h42727bc4};
test_index[5846] = '{1};
test_input[46776:46783] = '{32'hc1920ceb, 32'h41d6a885, 32'hc210cd8f, 32'hc23d67a7, 32'h40248bfa, 32'h42a2256f, 32'h42bd9ec9, 32'h426873ef};
test_output[5847] = '{32'h42bd9ec9};
test_index[5847] = '{6};
test_input[46784:46791] = '{32'h4296da3e, 32'hc1c5ea55, 32'hc2c03a53, 32'h41772510, 32'hc2b38c58, 32'h40b99c26, 32'h429fd2fb, 32'h41914473};
test_output[5848] = '{32'h429fd2fb};
test_index[5848] = '{6};
test_input[46792:46799] = '{32'hc2a0a95d, 32'h417ce6a3, 32'hc2932947, 32'hc0becc54, 32'h42218350, 32'hc263f286, 32'h42ab51b8, 32'h4154aa8b};
test_output[5849] = '{32'h42ab51b8};
test_index[5849] = '{6};
test_input[46800:46807] = '{32'h4275f8ef, 32'hc2ac2f77, 32'hc2564927, 32'h42641b59, 32'h429c405a, 32'hc2bfe436, 32'h42c23c36, 32'h4251aed8};
test_output[5850] = '{32'h42c23c36};
test_index[5850] = '{6};
test_input[46808:46815] = '{32'h42316982, 32'h42258d79, 32'h4234cab1, 32'hc14fab71, 32'hc25080b6, 32'hc251c229, 32'hc102b76f, 32'hc243b83a};
test_output[5851] = '{32'h4234cab1};
test_index[5851] = '{2};
test_input[46816:46823] = '{32'h41f54948, 32'hc210bdd0, 32'hc2c20af5, 32'hc27b4d2c, 32'hc1ffd5f9, 32'hc1ff1ff9, 32'hc211dd06, 32'hc2504455};
test_output[5852] = '{32'h41f54948};
test_index[5852] = '{0};
test_input[46824:46831] = '{32'hc28d644c, 32'h422b31c2, 32'hc2a28560, 32'h428e5c36, 32'h428786d6, 32'h3fdf8455, 32'h42b503af, 32'h421b3906};
test_output[5853] = '{32'h42b503af};
test_index[5853] = '{6};
test_input[46832:46839] = '{32'hc0fd2e30, 32'hc0e68b36, 32'h41dda39a, 32'hc294d345, 32'h40662f50, 32'hc19b9002, 32'h423b8490, 32'h4223a23e};
test_output[5854] = '{32'h423b8490};
test_index[5854] = '{6};
test_input[46840:46847] = '{32'h42c47ecd, 32'hc2b78c60, 32'hc0b6d4b9, 32'hc16ddd05, 32'h429ad0b0, 32'h426b27f7, 32'hc23d27f8, 32'h422f23b4};
test_output[5855] = '{32'h42c47ecd};
test_index[5855] = '{0};
test_input[46848:46855] = '{32'h42c03c92, 32'hc2bfade9, 32'hc1838be0, 32'h41d1d4f5, 32'hc27862e1, 32'hc1c57c42, 32'hc26131a5, 32'hc131efaa};
test_output[5856] = '{32'h42c03c92};
test_index[5856] = '{0};
test_input[46856:46863] = '{32'hc28ea77b, 32'h42744841, 32'hc27be558, 32'h428ada8e, 32'hc2b1c7d1, 32'h422dabe0, 32'hc1955ca9, 32'hc23d74a5};
test_output[5857] = '{32'h428ada8e};
test_index[5857] = '{3};
test_input[46864:46871] = '{32'h42389977, 32'h42616892, 32'h42907439, 32'h429ec28e, 32'h413211e1, 32'h4271e7e5, 32'hc2bfcb4c, 32'h42409194};
test_output[5858] = '{32'h429ec28e};
test_index[5858] = '{3};
test_input[46872:46879] = '{32'hc1cd4a5a, 32'h429830ef, 32'hc16cfc66, 32'h41fd43da, 32'hc22c2b96, 32'hc1082fb4, 32'hc2c3b6aa, 32'hc25f36f7};
test_output[5859] = '{32'h429830ef};
test_index[5859] = '{1};
test_input[46880:46887] = '{32'h42047a39, 32'hc23ee1f1, 32'hc294b1de, 32'h42b66e9b, 32'h41dfb0ad, 32'h41668890, 32'hc006bea1, 32'hc06ea758};
test_output[5860] = '{32'h42b66e9b};
test_index[5860] = '{3};
test_input[46888:46895] = '{32'h40d72f9c, 32'hc19f4cb6, 32'hc27d006f, 32'hc29286d4, 32'h4233ed15, 32'h42112f78, 32'hc1ebca25, 32'h4261eb6c};
test_output[5861] = '{32'h4261eb6c};
test_index[5861] = '{7};
test_input[46896:46903] = '{32'hc1def6f7, 32'hc230bdc6, 32'h414d63ca, 32'h425b6b44, 32'hc272469e, 32'h42638ad0, 32'h4224807b, 32'h41c2d642};
test_output[5862] = '{32'h42638ad0};
test_index[5862] = '{5};
test_input[46904:46911] = '{32'h4212de75, 32'hc20f95bb, 32'hc2b87ad2, 32'hc1bdc6e0, 32'h41ba05fe, 32'hc25a22be, 32'h41a5ceff, 32'hc0e7b41e};
test_output[5863] = '{32'h4212de75};
test_index[5863] = '{0};
test_input[46912:46919] = '{32'hc21c6e4c, 32'h41332bcb, 32'hc2843547, 32'h42ae3dd8, 32'hc2c67761, 32'h424746bd, 32'h42b74763, 32'h42b52701};
test_output[5864] = '{32'h42b74763};
test_index[5864] = '{6};
test_input[46920:46927] = '{32'hc228c6ca, 32'hc1fb8625, 32'hc139eacb, 32'hc1663fd8, 32'hc23424ff, 32'h41b90b01, 32'h41d1c7c8, 32'hc2b41dd7};
test_output[5865] = '{32'h41d1c7c8};
test_index[5865] = '{6};
test_input[46928:46935] = '{32'hc26c6f2a, 32'hc29899b5, 32'h42b81f39, 32'h42956fd9, 32'hc202510a, 32'hc2c1584b, 32'hc2035f31, 32'hc13566e4};
test_output[5866] = '{32'h42b81f39};
test_index[5866] = '{2};
test_input[46936:46943] = '{32'h41bbba66, 32'h41f324e9, 32'hc2977751, 32'hc28340b0, 32'h42c41882, 32'hc28972d2, 32'hc12beab1, 32'hc0493727};
test_output[5867] = '{32'h42c41882};
test_index[5867] = '{4};
test_input[46944:46951] = '{32'hc20c5a98, 32'hc2bd7be2, 32'hc212b4cd, 32'hc28f08e6, 32'hc194312e, 32'h4203814d, 32'hc2c6fb1e, 32'hc29bfc46};
test_output[5868] = '{32'h4203814d};
test_index[5868] = '{5};
test_input[46952:46959] = '{32'h42816cef, 32'h4210daf3, 32'hc29bd97e, 32'hc2a69e11, 32'hc25ae38e, 32'hc21504d9, 32'h429cebde, 32'hc20ea96e};
test_output[5869] = '{32'h429cebde};
test_index[5869] = '{6};
test_input[46960:46967] = '{32'h41a1cd31, 32'h429336e4, 32'hc291d0e2, 32'h42ab18e0, 32'hc2badf4a, 32'h42824f24, 32'h4208eaa3, 32'h41b72f67};
test_output[5870] = '{32'h42ab18e0};
test_index[5870] = '{3};
test_input[46968:46975] = '{32'h41d81359, 32'hc297de10, 32'hc2b1e67f, 32'hc290554b, 32'hc2bcf6cc, 32'hc1a410f4, 32'hc23ebc9e, 32'h42195b8f};
test_output[5871] = '{32'h42195b8f};
test_index[5871] = '{7};
test_input[46976:46983] = '{32'h421e5d40, 32'hc288387c, 32'hc276eea3, 32'h423ad2a5, 32'h3f0833f7, 32'hc142bf32, 32'hc2b3b16c, 32'h41d349be};
test_output[5872] = '{32'h423ad2a5};
test_index[5872] = '{3};
test_input[46984:46991] = '{32'h42599380, 32'hc24039b8, 32'hc1a7aae2, 32'hc299ef4c, 32'hc29c3c1a, 32'hc2b1304b, 32'hc292a542, 32'h42c7286a};
test_output[5873] = '{32'h42c7286a};
test_index[5873] = '{7};
test_input[46992:46999] = '{32'hc1667f1d, 32'h3f3855c7, 32'hc28a73ea, 32'h415777c0, 32'hc2b4f68a, 32'hc2bac191, 32'hc21cc095, 32'h4244a621};
test_output[5874] = '{32'h4244a621};
test_index[5874] = '{7};
test_input[47000:47007] = '{32'h426bcd2c, 32'hc2a6d53c, 32'hc1897c24, 32'h4050a788, 32'h421bad2d, 32'h42a47f57, 32'hc248c765, 32'h41e8b39d};
test_output[5875] = '{32'h42a47f57};
test_index[5875] = '{5};
test_input[47008:47015] = '{32'h425a3155, 32'h421ac60d, 32'h4195b89f, 32'hc2b3e554, 32'h418bd05a, 32'hc2671091, 32'hbe8e8c2f, 32'h42ba0f3e};
test_output[5876] = '{32'h42ba0f3e};
test_index[5876] = '{7};
test_input[47016:47023] = '{32'hc0b0f51d, 32'h4214202f, 32'hc216d636, 32'hc28f1a09, 32'h4206bb2e, 32'hc288c65a, 32'hc145b966, 32'h42aeec9a};
test_output[5877] = '{32'h42aeec9a};
test_index[5877] = '{7};
test_input[47024:47031] = '{32'hc12dcfeb, 32'h4103b8ab, 32'h41dc4d95, 32'hc29a5e01, 32'h40872004, 32'h41cbff32, 32'hc1164a7c, 32'hc1508380};
test_output[5878] = '{32'h41dc4d95};
test_index[5878] = '{2};
test_input[47032:47039] = '{32'hc2a62b37, 32'h428ff501, 32'hc296a3eb, 32'h419db346, 32'h424714e8, 32'hc2654b52, 32'h4258129c, 32'h413a906b};
test_output[5879] = '{32'h428ff501};
test_index[5879] = '{1};
test_input[47040:47047] = '{32'h4295c4c2, 32'h428ab9ae, 32'hc19c9214, 32'h42c7df48, 32'hc27cad2f, 32'h4052bcc8, 32'hc1b47660, 32'hc15a2631};
test_output[5880] = '{32'h42c7df48};
test_index[5880] = '{3};
test_input[47048:47055] = '{32'hc272c7d2, 32'hc211a4dc, 32'hc15d2a78, 32'h4236ed20, 32'hc2a2c2c7, 32'hc2a610f2, 32'h42504f17, 32'h4058ef19};
test_output[5881] = '{32'h42504f17};
test_index[5881] = '{6};
test_input[47056:47063] = '{32'h4243c32f, 32'h422c8ada, 32'hc27985bb, 32'hc22d82c3, 32'h41d6fe6d, 32'hc14504e2, 32'h426154a6, 32'hc1cfbcbf};
test_output[5882] = '{32'h426154a6};
test_index[5882] = '{6};
test_input[47064:47071] = '{32'hc28755a5, 32'hc297483c, 32'h4270462b, 32'hc273aa74, 32'hc27f540a, 32'hc22e9597, 32'hc2a70ba9, 32'h42c3e5db};
test_output[5883] = '{32'h42c3e5db};
test_index[5883] = '{7};
test_input[47072:47079] = '{32'hc2bb1e24, 32'hc1112c52, 32'h42b47c95, 32'hc2a40452, 32'h42748732, 32'hc2249896, 32'h42b7f5e6, 32'hc2b707f4};
test_output[5884] = '{32'h42b7f5e6};
test_index[5884] = '{6};
test_input[47080:47087] = '{32'hc2194564, 32'hc15b9efa, 32'hc295bccf, 32'h418f3270, 32'hc1ea41c9, 32'h4179cf93, 32'hc1f7011c, 32'hc1c392df};
test_output[5885] = '{32'h418f3270};
test_index[5885] = '{3};
test_input[47088:47095] = '{32'h428e7269, 32'hbf6b48c8, 32'h42a038ed, 32'hc2c0bafc, 32'h42a2202b, 32'h3f9068e8, 32'h40cae078, 32'hc2bcc06c};
test_output[5886] = '{32'h42a2202b};
test_index[5886] = '{4};
test_input[47096:47103] = '{32'hc29b6d25, 32'hc0a78368, 32'h4235d817, 32'hc24f13be, 32'hc2b84d57, 32'hc26139a8, 32'h42a8b7b4, 32'h42c260b0};
test_output[5887] = '{32'h42c260b0};
test_index[5887] = '{7};
test_input[47104:47111] = '{32'hc152d6a6, 32'hc289914c, 32'hc1eac222, 32'hc292d10e, 32'h41da98c2, 32'h411d02d4, 32'h423852aa, 32'h42b219b2};
test_output[5888] = '{32'h42b219b2};
test_index[5888] = '{7};
test_input[47112:47119] = '{32'h41ef5e0b, 32'h4132b8fc, 32'hc1df5b78, 32'hc2b2ac0f, 32'hc235e800, 32'h429a461d, 32'h40f9301b, 32'hc1eced0e};
test_output[5889] = '{32'h429a461d};
test_index[5889] = '{5};
test_input[47120:47127] = '{32'hc2a129f3, 32'hc0fe855c, 32'h42b70950, 32'hc17ef1b1, 32'h41133883, 32'h42b57a6c, 32'h41ac2a8e, 32'h42a7bc5b};
test_output[5890] = '{32'h42b70950};
test_index[5890] = '{2};
test_input[47128:47135] = '{32'h42bc8c09, 32'h4281872b, 32'h420a3590, 32'h428f6f86, 32'h428b33ac, 32'hc263d969, 32'hc2a0497d, 32'h42a477ce};
test_output[5891] = '{32'h42bc8c09};
test_index[5891] = '{0};
test_input[47136:47143] = '{32'h41c3f6d4, 32'h42184c9f, 32'hc2b4d8bb, 32'h42b218f4, 32'h41d38f32, 32'h4118c117, 32'h4211e452, 32'h42a617c5};
test_output[5892] = '{32'h42b218f4};
test_index[5892] = '{3};
test_input[47144:47151] = '{32'h425b4c24, 32'hc23a335e, 32'hc1360110, 32'h42321d41, 32'hc2169b65, 32'hc141dbd0, 32'hc1d6a566, 32'hc24c28e5};
test_output[5893] = '{32'h425b4c24};
test_index[5893] = '{0};
test_input[47152:47159] = '{32'hc18627b1, 32'h4247529e, 32'hc2b043b9, 32'hc07ca7ea, 32'hc21e76f0, 32'hc2728032, 32'hc2281e9d, 32'hc19e1523};
test_output[5894] = '{32'h4247529e};
test_index[5894] = '{1};
test_input[47160:47167] = '{32'h429b70df, 32'hc2955c09, 32'hc1734e9e, 32'h40bb322e, 32'h42ae3ff1, 32'hc271e6f5, 32'h41c8c82c, 32'hc2c4e4b1};
test_output[5895] = '{32'h42ae3ff1};
test_index[5895] = '{4};
test_input[47168:47175] = '{32'h428aeb71, 32'h4288d057, 32'h429fcb33, 32'h418fa712, 32'hc2c65dae, 32'h41fc05cf, 32'h41dab634, 32'h427d85d4};
test_output[5896] = '{32'h429fcb33};
test_index[5896] = '{2};
test_input[47176:47183] = '{32'hc237516a, 32'hc285e24c, 32'h428e3f57, 32'hc211b7f5, 32'h42664a9b, 32'h41ee79f0, 32'hc2bd162e, 32'hc27309e8};
test_output[5897] = '{32'h428e3f57};
test_index[5897] = '{2};
test_input[47184:47191] = '{32'h425445f2, 32'h42a1b95e, 32'h422c3167, 32'hc2b4fd3b, 32'hc1c61c20, 32'hc1abf75f, 32'hc2b491aa, 32'hc2810961};
test_output[5898] = '{32'h42a1b95e};
test_index[5898] = '{1};
test_input[47192:47199] = '{32'hc12ef5c5, 32'h424c4086, 32'hc1a6d6c7, 32'h42a4b9b0, 32'hc1ec4754, 32'hc28f98db, 32'hc2c02df1, 32'h41590fd5};
test_output[5899] = '{32'h42a4b9b0};
test_index[5899] = '{3};
test_input[47200:47207] = '{32'h429383d3, 32'h42c4739c, 32'h423bea1a, 32'hc23f54f2, 32'h400c68e0, 32'hc1a0de47, 32'h3fc79720, 32'hc1d64f3f};
test_output[5900] = '{32'h42c4739c};
test_index[5900] = '{1};
test_input[47208:47215] = '{32'hc293886e, 32'hc2c20c6f, 32'hc11a3c37, 32'hc1e4623e, 32'h40b14fee, 32'hc2a3a684, 32'h424ee78c, 32'h41461e72};
test_output[5901] = '{32'h424ee78c};
test_index[5901] = '{6};
test_input[47216:47223] = '{32'h40a23647, 32'h42b9563a, 32'hc2bac013, 32'hc2494fde, 32'h42303996, 32'h41d3c362, 32'h42aa31cf, 32'h4287b638};
test_output[5902] = '{32'h42b9563a};
test_index[5902] = '{1};
test_input[47224:47231] = '{32'hc27d9fe1, 32'hc265b4e8, 32'hc0593019, 32'hc0a50cd5, 32'hc2c2a5f6, 32'hc296f827, 32'h42277470, 32'h41fc5eb5};
test_output[5903] = '{32'h42277470};
test_index[5903] = '{6};
test_input[47232:47239] = '{32'h4182a4ae, 32'h4102235d, 32'h4218d8d6, 32'hc11bbd66, 32'h4285f535, 32'h423391f4, 32'h428df2d8, 32'h42a56716};
test_output[5904] = '{32'h42a56716};
test_index[5904] = '{7};
test_input[47240:47247] = '{32'hc15f94a4, 32'h42648e53, 32'h4229fb65, 32'h41efa635, 32'hc1059fd3, 32'h42b4f898, 32'hc16bf3aa, 32'h4230b430};
test_output[5905] = '{32'h42b4f898};
test_index[5905] = '{5};
test_input[47248:47255] = '{32'hc1aac6a9, 32'hc1153ca6, 32'h42847929, 32'h42a77e82, 32'h4191dac2, 32'hc2bcef68, 32'hc1f3d7d6, 32'h42a4dfd9};
test_output[5906] = '{32'h42a77e82};
test_index[5906] = '{3};
test_input[47256:47263] = '{32'h4254a940, 32'h422625b9, 32'hc203eabf, 32'h42a973c8, 32'h42b426e9, 32'h4214690d, 32'h42351a33, 32'h42c3ea9e};
test_output[5907] = '{32'h42c3ea9e};
test_index[5907] = '{7};
test_input[47264:47271] = '{32'h425ddb33, 32'hc1a8f1c1, 32'hc2b8f356, 32'h4218288a, 32'hc1dcd1e2, 32'h42051e12, 32'h42912aa7, 32'hc2618c82};
test_output[5908] = '{32'h42912aa7};
test_index[5908] = '{6};
test_input[47272:47279] = '{32'hc29a6cc3, 32'h42b1e2a8, 32'h41ede53b, 32'h425e120c, 32'h428ad1d5, 32'hc2a5a9eb, 32'hc05f6b8b, 32'hc166baf9};
test_output[5909] = '{32'h42b1e2a8};
test_index[5909] = '{1};
test_input[47280:47287] = '{32'h4218d5de, 32'hc232842c, 32'h423c99d5, 32'hc0a01275, 32'h42c76674, 32'hc1a03701, 32'h41f27a01, 32'hc2284695};
test_output[5910] = '{32'h42c76674};
test_index[5910] = '{4};
test_input[47288:47295] = '{32'hc1ff11e8, 32'hc25e2a7b, 32'h429a8963, 32'h42c099eb, 32'hc2327e42, 32'h40af26ec, 32'hc24ebefc, 32'hc2afd035};
test_output[5911] = '{32'h42c099eb};
test_index[5911] = '{3};
test_input[47296:47303] = '{32'hc2a4a2f7, 32'hc20c0a32, 32'hc291c695, 32'h421f7867, 32'hc179d8c5, 32'h423599ca, 32'h422e5cce, 32'h411daa1a};
test_output[5912] = '{32'h423599ca};
test_index[5912] = '{5};
test_input[47304:47311] = '{32'h42308721, 32'hbef272d8, 32'hc0601709, 32'hc29e0568, 32'h4294a0e6, 32'h4281496e, 32'hc2936891, 32'h42b244a0};
test_output[5913] = '{32'h42b244a0};
test_index[5913] = '{7};
test_input[47312:47319] = '{32'hc2067a1b, 32'h4231ffd2, 32'h4104f5a6, 32'h411dbe66, 32'hc2692ccd, 32'hc1b3b0c0, 32'h420f3fe1, 32'h42930583};
test_output[5914] = '{32'h42930583};
test_index[5914] = '{7};
test_input[47320:47327] = '{32'hc0930670, 32'h42c78448, 32'hc2930439, 32'hc237f56e, 32'hc198848a, 32'hc2c11f4b, 32'hc2b92a8e, 32'hc26a0856};
test_output[5915] = '{32'h42c78448};
test_index[5915] = '{1};
test_input[47328:47335] = '{32'hc206bb98, 32'hc2afed86, 32'h42a190e2, 32'h429d97db, 32'hc259a8c7, 32'hc2c0bdd9, 32'h41f809db, 32'hc2b056cb};
test_output[5916] = '{32'h42a190e2};
test_index[5916] = '{2};
test_input[47336:47343] = '{32'hc1a4c54e, 32'hc2666528, 32'hc2be3cb0, 32'hc18e37ed, 32'hc21f1279, 32'hbec1cc2f, 32'hc24d7494, 32'hc278df79};
test_output[5917] = '{32'hbec1cc2f};
test_index[5917] = '{5};
test_input[47344:47351] = '{32'h42ad3d4f, 32'hc2234443, 32'h42bbabf3, 32'hc2bd696b, 32'hc19a6b7f, 32'hc2a890d2, 32'hc1387548, 32'hc28bdc53};
test_output[5918] = '{32'h42bbabf3};
test_index[5918] = '{2};
test_input[47352:47359] = '{32'hc2398ea5, 32'h42a8c2e2, 32'h420b3c43, 32'hc2afc8e3, 32'h41a3dbf0, 32'h41a07ab1, 32'h42132576, 32'hc2a6db6d};
test_output[5919] = '{32'h42a8c2e2};
test_index[5919] = '{1};
test_input[47360:47367] = '{32'h427df311, 32'h421d6a62, 32'h41851f63, 32'h417d8c47, 32'hc2bf75dc, 32'hc2b7d78e, 32'h41887acf, 32'h4238b3d2};
test_output[5920] = '{32'h427df311};
test_index[5920] = '{0};
test_input[47368:47375] = '{32'hc0b978f0, 32'h42357587, 32'h4291d2cf, 32'h429a520a, 32'hc0b6a587, 32'hc2422340, 32'hc2c079a4, 32'h4202e8e6};
test_output[5921] = '{32'h429a520a};
test_index[5921] = '{3};
test_input[47376:47383] = '{32'hc1a07565, 32'h42a73990, 32'hc2c309b5, 32'h40bdeec0, 32'h42697050, 32'hc11a63c7, 32'hc202e951, 32'hc2362198};
test_output[5922] = '{32'h42a73990};
test_index[5922] = '{1};
test_input[47384:47391] = '{32'h410d6b4a, 32'h4242ef7a, 32'hc1720ea9, 32'hc2aac79a, 32'h4299eefb, 32'h428308e1, 32'hc2a317dd, 32'h4143960a};
test_output[5923] = '{32'h4299eefb};
test_index[5923] = '{4};
test_input[47392:47399] = '{32'hc210f145, 32'hc2a072d2, 32'h413ba06b, 32'hc2549474, 32'hc1a90c78, 32'hc17608b2, 32'h41be5498, 32'h42324c4f};
test_output[5924] = '{32'h42324c4f};
test_index[5924] = '{7};
test_input[47400:47407] = '{32'hc2890904, 32'hc2a5b6cf, 32'h428d94bb, 32'hc281da2e, 32'hc17e0b2e, 32'hc2873429, 32'h427aaaba, 32'hc0c765cf};
test_output[5925] = '{32'h428d94bb};
test_index[5925] = '{2};
test_input[47408:47415] = '{32'h41ea5a91, 32'hc27236d1, 32'hc21e75aa, 32'hc197710f, 32'hc282544c, 32'hc2504cc6, 32'h4246fccd, 32'hc2834cf2};
test_output[5926] = '{32'h4246fccd};
test_index[5926] = '{6};
test_input[47416:47423] = '{32'h423f8012, 32'h42587a7c, 32'h42a06184, 32'hc254d5e9, 32'h41049d7a, 32'hc2993d12, 32'h40221d80, 32'h42a49bc2};
test_output[5927] = '{32'h42a49bc2};
test_index[5927] = '{7};
test_input[47424:47431] = '{32'hc2507e32, 32'hc2bf7c72, 32'hc297150f, 32'h42c30725, 32'h42a82711, 32'hc1ffe55b, 32'hc2afae2c, 32'h4241e74a};
test_output[5928] = '{32'h42c30725};
test_index[5928] = '{3};
test_input[47432:47439] = '{32'hc29c9127, 32'h42735a3d, 32'h4206e7e0, 32'h421a7746, 32'h41dbf458, 32'hc1fbcec8, 32'hc18ca89f, 32'hc18a9ae6};
test_output[5929] = '{32'h42735a3d};
test_index[5929] = '{1};
test_input[47440:47447] = '{32'h423aa489, 32'h41c42533, 32'h426b58f1, 32'hc2789fa0, 32'h423e52c6, 32'h4281e789, 32'hc2c1a2c4, 32'h423e921f};
test_output[5930] = '{32'h4281e789};
test_index[5930] = '{5};
test_input[47448:47455] = '{32'h426d9620, 32'h41006c02, 32'h42475f63, 32'h41c02a52, 32'hc2912d69, 32'h416abad4, 32'h4240d56e, 32'h42c28915};
test_output[5931] = '{32'h42c28915};
test_index[5931] = '{7};
test_input[47456:47463] = '{32'h428732a0, 32'hc1aa10d7, 32'h42c6c7fb, 32'h4294fe61, 32'h429e7e8c, 32'h426df527, 32'hc28c1e2a, 32'h4251c45c};
test_output[5932] = '{32'h42c6c7fb};
test_index[5932] = '{2};
test_input[47464:47471] = '{32'h42a62a30, 32'h419e2b78, 32'hbf873498, 32'h42903b8b, 32'h4273ed22, 32'hc28088ed, 32'hc1e2eaff, 32'hc07ff147};
test_output[5933] = '{32'h42a62a30};
test_index[5933] = '{0};
test_input[47472:47479] = '{32'hc2881788, 32'h4284ed8e, 32'h428d90ef, 32'h4149187a, 32'hc20efd69, 32'hc1323e48, 32'h42a1a2a4, 32'h41760bc3};
test_output[5934] = '{32'h42a1a2a4};
test_index[5934] = '{6};
test_input[47480:47487] = '{32'h428b8088, 32'h42c0a4a9, 32'hc0f19818, 32'h42be2e87, 32'hc290ba75, 32'h417034f3, 32'hc24820a1, 32'hc279a57b};
test_output[5935] = '{32'h42c0a4a9};
test_index[5935] = '{1};
test_input[47488:47495] = '{32'hc19bea68, 32'hc21df9e2, 32'hc240d86d, 32'hc251b85b, 32'h4284f6da, 32'hc28f0f9e, 32'h42c0b353, 32'hc2675c3a};
test_output[5936] = '{32'h42c0b353};
test_index[5936] = '{6};
test_input[47496:47503] = '{32'hc29ebf36, 32'h41fdce8c, 32'hc2243008, 32'hc1ec5764, 32'hc29e05f3, 32'hc26568b3, 32'h4243ff2a, 32'hc2b52e93};
test_output[5937] = '{32'h4243ff2a};
test_index[5937] = '{6};
test_input[47504:47511] = '{32'h4260d4fa, 32'hc20722c9, 32'hc2c7848d, 32'h425084b4, 32'hc2a86978, 32'hc26ac921, 32'hc156eff1, 32'h42854168};
test_output[5938] = '{32'h42854168};
test_index[5938] = '{7};
test_input[47512:47519] = '{32'hc2a3c9a4, 32'h42a418fc, 32'h42af174e, 32'hc28b0f04, 32'hc2537f5e, 32'h429ae3b9, 32'hc2c1d289, 32'hc2664739};
test_output[5939] = '{32'h42af174e};
test_index[5939] = '{2};
test_input[47520:47527] = '{32'h41c17594, 32'hc149a229, 32'hc2b137d7, 32'hc23bfe8e, 32'hc22a571e, 32'hc2477054, 32'h416bf1ae, 32'h42bb5f66};
test_output[5940] = '{32'h42bb5f66};
test_index[5940] = '{7};
test_input[47528:47535] = '{32'h429d6ec4, 32'h41e81f08, 32'hc237417a, 32'h42144a15, 32'h4297f760, 32'hc1db2e77, 32'h42954c4d, 32'h4229adde};
test_output[5941] = '{32'h429d6ec4};
test_index[5941] = '{0};
test_input[47536:47543] = '{32'h40a45bac, 32'h422dbc44, 32'hc08cedba, 32'h429e5679, 32'h428083bd, 32'hc27a30bf, 32'hc2a5a8bb, 32'hc2126ad9};
test_output[5942] = '{32'h429e5679};
test_index[5942] = '{3};
test_input[47544:47551] = '{32'hc1ad0a1a, 32'hc28fc13f, 32'hc28be86c, 32'hc26a4c6e, 32'h42c7b76f, 32'hc0c6e0d1, 32'h42aef593, 32'hc2a12632};
test_output[5943] = '{32'h42c7b76f};
test_index[5943] = '{4};
test_input[47552:47559] = '{32'h420f2fb8, 32'h41b708e3, 32'hc22f787d, 32'hc191749c, 32'hc2a0bc7c, 32'h4113e549, 32'hbf8323c3, 32'hc1e5e7ca};
test_output[5944] = '{32'h420f2fb8};
test_index[5944] = '{0};
test_input[47560:47567] = '{32'h42af51b2, 32'h42033c6a, 32'h422eba98, 32'h4283d312, 32'hc22b799e, 32'hc293c6c9, 32'hc2bd7aa3, 32'h428600f6};
test_output[5945] = '{32'h42af51b2};
test_index[5945] = '{0};
test_input[47568:47575] = '{32'h42803b4f, 32'h42a4b290, 32'h42aaa9d6, 32'h42b8e663, 32'hc1316772, 32'hc1595932, 32'h42b6a750, 32'hc2c79afb};
test_output[5946] = '{32'h42b8e663};
test_index[5946] = '{3};
test_input[47576:47583] = '{32'h42b44af6, 32'h422a430b, 32'h41a76a7e, 32'hc2133655, 32'h428949bf, 32'h4151dae9, 32'hc28c3431, 32'h3fd86253};
test_output[5947] = '{32'h42b44af6};
test_index[5947] = '{0};
test_input[47584:47591] = '{32'h40897589, 32'h4287b596, 32'h42c27023, 32'hc2384211, 32'hc2190003, 32'h40db7937, 32'hc26274a7, 32'h41a64619};
test_output[5948] = '{32'h42c27023};
test_index[5948] = '{2};
test_input[47592:47599] = '{32'hc248776c, 32'hc21165f7, 32'h41825a8e, 32'hc20d9c02, 32'h42a0efb6, 32'h419006d8, 32'h4258c5d4, 32'h42c39ab5};
test_output[5949] = '{32'h42c39ab5};
test_index[5949] = '{7};
test_input[47600:47607] = '{32'h41c8944e, 32'h429cba19, 32'hc2affa2d, 32'hc248b5e0, 32'h422e53e0, 32'hc28b2b7d, 32'h4115fc09, 32'h429fd324};
test_output[5950] = '{32'h429fd324};
test_index[5950] = '{7};
test_input[47608:47615] = '{32'hc1771bae, 32'hc2aa9d1e, 32'hc26af027, 32'h42b6aa86, 32'h42864e7a, 32'h41f93c5c, 32'hc282dcd0, 32'h41d765bf};
test_output[5951] = '{32'h42b6aa86};
test_index[5951] = '{3};
test_input[47616:47623] = '{32'hc2a37d24, 32'hc13b0782, 32'h3f6ea71f, 32'hc29c9add, 32'hc2b2ee0d, 32'h419d31ca, 32'hc2950ca5, 32'hc0c87f1d};
test_output[5952] = '{32'h419d31ca};
test_index[5952] = '{5};
test_input[47624:47631] = '{32'hc226de13, 32'hc1f12fd5, 32'hc1387774, 32'h41c80a05, 32'h42446e0d, 32'hc202f045, 32'h42c3cee7, 32'hc230b04f};
test_output[5953] = '{32'h42c3cee7};
test_index[5953] = '{6};
test_input[47632:47639] = '{32'h4203a8ce, 32'hc24046ed, 32'h426e6a20, 32'h415dcb73, 32'hc29d4086, 32'h4239cf0e, 32'h41dd0307, 32'hc1fad7a6};
test_output[5954] = '{32'h426e6a20};
test_index[5954] = '{2};
test_input[47640:47647] = '{32'hc20043dd, 32'hc29e303e, 32'hc23b9d48, 32'hc1ecfa7c, 32'hc1f6c59d, 32'hc2656bb5, 32'h429ae80a, 32'h429d934b};
test_output[5955] = '{32'h429d934b};
test_index[5955] = '{7};
test_input[47648:47655] = '{32'hc0156818, 32'hc1e07112, 32'h41e84f43, 32'hc2b56678, 32'h41fe4e7d, 32'h42414357, 32'h41985db7, 32'hc2100526};
test_output[5956] = '{32'h42414357};
test_index[5956] = '{5};
test_input[47656:47663] = '{32'h40afb676, 32'hc2494410, 32'hc276ef11, 32'hc29dad53, 32'h420736bc, 32'h42b27738, 32'hc271ac67, 32'hc228b7b8};
test_output[5957] = '{32'h42b27738};
test_index[5957] = '{5};
test_input[47664:47671] = '{32'h415daa7d, 32'h41f6c4a5, 32'hc25452de, 32'hc24bb90e, 32'hc1bef560, 32'h420d4d2d, 32'h41e1ce2a, 32'h42522aa8};
test_output[5958] = '{32'h42522aa8};
test_index[5958] = '{7};
test_input[47672:47679] = '{32'hc24df193, 32'hc25cce76, 32'h41195597, 32'hc24cf6a9, 32'hc2887330, 32'hc2b30b5e, 32'h4273bc92, 32'hc220a700};
test_output[5959] = '{32'h4273bc92};
test_index[5959] = '{6};
test_input[47680:47687] = '{32'h42af19a1, 32'hc18614d1, 32'h406aadb5, 32'hc1f505c4, 32'hc2227fb4, 32'h42765b4b, 32'hbe566e51, 32'hc13d840e};
test_output[5960] = '{32'h42af19a1};
test_index[5960] = '{0};
test_input[47688:47695] = '{32'hc299df6a, 32'h4281d17b, 32'h41f4785a, 32'hc1b59822, 32'hc09e838d, 32'hc263162b, 32'h4297a048, 32'h41131c44};
test_output[5961] = '{32'h4297a048};
test_index[5961] = '{6};
test_input[47696:47703] = '{32'h4210fd41, 32'hc2c35632, 32'h407d6639, 32'h419448a4, 32'hc16a172f, 32'hc29e5785, 32'h428943ab, 32'hc0e1b9e1};
test_output[5962] = '{32'h428943ab};
test_index[5962] = '{6};
test_input[47704:47711] = '{32'hc13063da, 32'h424eb607, 32'hc10f5cd4, 32'hc1e64d7a, 32'hc2617743, 32'h41ee1b41, 32'h41cddd4f, 32'h423a13ae};
test_output[5963] = '{32'h424eb607};
test_index[5963] = '{1};
test_input[47712:47719] = '{32'h42c65e76, 32'h41846f8a, 32'h425e12d6, 32'h3f447682, 32'hc1fffb64, 32'hc28123bf, 32'h413257be, 32'hc1b26434};
test_output[5964] = '{32'h42c65e76};
test_index[5964] = '{0};
test_input[47720:47727] = '{32'h4237f70b, 32'hc1bd4168, 32'hc1d88a7e, 32'h41965e9c, 32'hc1b58eb1, 32'h41d12d80, 32'hc1cf5263, 32'h42b2e236};
test_output[5965] = '{32'h42b2e236};
test_index[5965] = '{7};
test_input[47728:47735] = '{32'h421521ac, 32'hc21a57ba, 32'hc2acffb7, 32'hbe03494e, 32'hc2c4abf2, 32'h429b699a, 32'hc298bc3b, 32'h41a87596};
test_output[5966] = '{32'h429b699a};
test_index[5966] = '{5};
test_input[47736:47743] = '{32'hc220ec9e, 32'h4109cdba, 32'h3fcd013b, 32'hc18b6d05, 32'hc22ccd05, 32'h40f24aff, 32'h428fe2b4, 32'hc12a3a5f};
test_output[5967] = '{32'h428fe2b4};
test_index[5967] = '{6};
test_input[47744:47751] = '{32'h420f8b98, 32'h3fb5081a, 32'hc2a83242, 32'h41e90d4f, 32'hc1b8ba94, 32'hc2c2a560, 32'hc21a01d6, 32'h42921c23};
test_output[5968] = '{32'h42921c23};
test_index[5968] = '{7};
test_input[47752:47759] = '{32'hc2ba35d0, 32'hc29d91cf, 32'hc1d58da7, 32'hc1bf2e0a, 32'hc2b14955, 32'hc2b56b36, 32'h42618f1a, 32'hc2a5cab6};
test_output[5969] = '{32'h42618f1a};
test_index[5969] = '{6};
test_input[47760:47767] = '{32'h4296d079, 32'h428bb122, 32'h42956fe1, 32'h42be9534, 32'h428be3ec, 32'h42b20b67, 32'h42bc679a, 32'h42271f8b};
test_output[5970] = '{32'h42be9534};
test_index[5970] = '{3};
test_input[47768:47775] = '{32'h420e8880, 32'hc2bb2595, 32'hc2ace264, 32'hc2a44eda, 32'hc2951f58, 32'hc19ba605, 32'h42769e18, 32'hc0a19b0d};
test_output[5971] = '{32'h42769e18};
test_index[5971] = '{6};
test_input[47776:47783] = '{32'h42a05b0a, 32'hc200159e, 32'hc2909331, 32'hc287fce4, 32'h4205ef01, 32'h41a06808, 32'hc283f32a, 32'hc22f525e};
test_output[5972] = '{32'h42a05b0a};
test_index[5972] = '{0};
test_input[47784:47791] = '{32'h42c009e8, 32'h40779844, 32'hc11f1639, 32'h41ff1959, 32'hc2404f73, 32'hc28436e3, 32'hc2bc1707, 32'hc284ee8c};
test_output[5973] = '{32'h42c009e8};
test_index[5973] = '{0};
test_input[47792:47799] = '{32'h4215fd2a, 32'hc21a6562, 32'hc1be3ff0, 32'hc2991bdb, 32'hc286709d, 32'h41c3739d, 32'h42b71faf, 32'hc2193b91};
test_output[5974] = '{32'h42b71faf};
test_index[5974] = '{6};
test_input[47800:47807] = '{32'h422daaad, 32'hc2754217, 32'h418e75f7, 32'h41f7b113, 32'h4253da37, 32'hc22b6339, 32'hc2bce47b, 32'hc264a6a2};
test_output[5975] = '{32'h4253da37};
test_index[5975] = '{4};
test_input[47808:47815] = '{32'h42706939, 32'hc01c2c93, 32'hc23e343f, 32'hc2a9b942, 32'h41b365ac, 32'hc29f691c, 32'h41273350, 32'hc2b28db3};
test_output[5976] = '{32'h42706939};
test_index[5976] = '{0};
test_input[47816:47823] = '{32'hc2744241, 32'hc1e4dcaf, 32'hc07f4150, 32'h42209781, 32'h422cbc56, 32'hc206d7a7, 32'hc121ff1a, 32'h4237a1ff};
test_output[5977] = '{32'h4237a1ff};
test_index[5977] = '{7};
test_input[47824:47831] = '{32'h42040873, 32'hc2703724, 32'hc2b68e01, 32'hc2c3ebe9, 32'hc2975aa5, 32'hc25c5bac, 32'hc204ea1b, 32'h4245cc76};
test_output[5978] = '{32'h4245cc76};
test_index[5978] = '{7};
test_input[47832:47839] = '{32'h41f0d3dc, 32'h42c6ddfc, 32'hc29f34f6, 32'hc21fddba, 32'h42c7fbf2, 32'h410ec2f5, 32'hc26340db, 32'h426f9294};
test_output[5979] = '{32'h42c7fbf2};
test_index[5979] = '{4};
test_input[47840:47847] = '{32'h41efb495, 32'hc2bd8f3e, 32'h4130293b, 32'hbf347e4f, 32'h42a5aa6f, 32'h424de631, 32'hc23cb5e9, 32'hc2380327};
test_output[5980] = '{32'h42a5aa6f};
test_index[5980] = '{4};
test_input[47848:47855] = '{32'h41cbef5e, 32'hc25e4d35, 32'hc25d7d77, 32'hc18395ad, 32'h425dcb1d, 32'h4224133d, 32'h421aa5ec, 32'hc1630781};
test_output[5981] = '{32'h425dcb1d};
test_index[5981] = '{4};
test_input[47856:47863] = '{32'h41b9f2a5, 32'hc0ce68ed, 32'h426a4720, 32'h41ed5273, 32'hc240cb0a, 32'hc2c290a9, 32'h420aa632, 32'hc001aa05};
test_output[5982] = '{32'h426a4720};
test_index[5982] = '{2};
test_input[47864:47871] = '{32'hc2b6460c, 32'hc2586a98, 32'h426222bd, 32'h42076700, 32'hc24e4caf, 32'hc201a7eb, 32'h42762167, 32'h42907ac1};
test_output[5983] = '{32'h42907ac1};
test_index[5983] = '{7};
test_input[47872:47879] = '{32'h42c28296, 32'h4253d4eb, 32'hc0afb299, 32'h41a298b9, 32'h42affb3f, 32'h41538e27, 32'h41d62b0d, 32'h429a8c68};
test_output[5984] = '{32'h42c28296};
test_index[5984] = '{0};
test_input[47880:47887] = '{32'hc22f7bfc, 32'hc20f26cf, 32'h41e48b67, 32'h4060e941, 32'hc244943e, 32'h429504c0, 32'hc282cd67, 32'hc2839ed2};
test_output[5985] = '{32'h429504c0};
test_index[5985] = '{5};
test_input[47888:47895] = '{32'hc2969f2c, 32'hc26ab0a8, 32'hc298c666, 32'h4244a623, 32'hc22a5ba8, 32'h413d6b64, 32'hc2ababa7, 32'hc27389c7};
test_output[5986] = '{32'h4244a623};
test_index[5986] = '{3};
test_input[47896:47903] = '{32'hc21219ef, 32'hc2b46982, 32'hc2a78d29, 32'h4120aae4, 32'hc0ecd899, 32'h426003ff, 32'hc17a6cc7, 32'h42288782};
test_output[5987] = '{32'h426003ff};
test_index[5987] = '{5};
test_input[47904:47911] = '{32'hc2a4bd79, 32'hc2c1402f, 32'h429b43b8, 32'hc25b25c9, 32'hc1ad3e05, 32'h4201e71a, 32'h42637878, 32'h41a39d54};
test_output[5988] = '{32'h429b43b8};
test_index[5988] = '{2};
test_input[47912:47919] = '{32'h4108aede, 32'hc2195881, 32'h42be34cf, 32'h4197b54d, 32'h420a1322, 32'hc20264f5, 32'hc22c7cdf, 32'h42094ca1};
test_output[5989] = '{32'h42be34cf};
test_index[5989] = '{2};
test_input[47920:47927] = '{32'h429ff0af, 32'h41b22bdf, 32'hc2848219, 32'h421be1b8, 32'h42a6510b, 32'h415b2a6e, 32'hc2bf44ea, 32'h428bd2c4};
test_output[5990] = '{32'h42a6510b};
test_index[5990] = '{4};
test_input[47928:47935] = '{32'h41417243, 32'h40f2af88, 32'hc2a357a0, 32'hc0f00d92, 32'h42c63442, 32'hc22b7497, 32'h428f766f, 32'h42a9c3e5};
test_output[5991] = '{32'h42c63442};
test_index[5991] = '{4};
test_input[47936:47943] = '{32'h4245f390, 32'h4204dc7b, 32'h429db709, 32'h42662177, 32'h41ee761d, 32'h428b0668, 32'h412f766d, 32'hc1f826d5};
test_output[5992] = '{32'h429db709};
test_index[5992] = '{2};
test_input[47944:47951] = '{32'h420e9bd7, 32'h42bec164, 32'h40478da5, 32'hc239b319, 32'hc163974e, 32'hc25a7e71, 32'hbfb1256d, 32'h42bd7e6c};
test_output[5993] = '{32'h42bec164};
test_index[5993] = '{1};
test_input[47952:47959] = '{32'hc2c1cd4b, 32'hc222cb36, 32'hc2afa9a8, 32'h424b0644, 32'hc20affb7, 32'hc08f0054, 32'hc2535d22, 32'hc282cf93};
test_output[5994] = '{32'h424b0644};
test_index[5994] = '{3};
test_input[47960:47967] = '{32'hc1dbaaf5, 32'hc094644d, 32'h41f5446d, 32'hc2b7297a, 32'hc287feff, 32'h423d2b70, 32'hc2ac8642, 32'hc0f46182};
test_output[5995] = '{32'h423d2b70};
test_index[5995] = '{5};
test_input[47968:47975] = '{32'h420843be, 32'hc2a8cad8, 32'h41ecbad3, 32'h420c8572, 32'h41140f00, 32'hc2b00195, 32'hc233b652, 32'h41ebacbb};
test_output[5996] = '{32'h420c8572};
test_index[5996] = '{3};
test_input[47976:47983] = '{32'h41f9c77f, 32'hc2521a43, 32'h41ced86f, 32'h41270e81, 32'hc234a44f, 32'hc19354be, 32'hc245ee2b, 32'hc2b01d69};
test_output[5997] = '{32'h41f9c77f};
test_index[5997] = '{0};
test_input[47984:47991] = '{32'hc0244aae, 32'hc1df38e2, 32'h4263372a, 32'hc2345557, 32'hc281cf2e, 32'h4281a9cf, 32'hc29ec031, 32'hc2097786};
test_output[5998] = '{32'h4281a9cf};
test_index[5998] = '{5};
test_input[47992:47999] = '{32'hc2c2e6f4, 32'h41e03d5a, 32'h42913831, 32'h42c2f862, 32'hc2764fec, 32'h42bb8955, 32'h41ff27fd, 32'hc28a90aa};
test_output[5999] = '{32'h42c2f862};
test_index[5999] = '{3};
test_input[48000:48007] = '{32'hc29462e5, 32'h41d0692e, 32'hc2aff970, 32'h4260a943, 32'h42bc18ae, 32'h42803a4d, 32'h4271501f, 32'hc1ac7692};
test_output[6000] = '{32'h42bc18ae};
test_index[6000] = '{4};
test_input[48008:48015] = '{32'hc267f74e, 32'hc22b1cc9, 32'h42173d47, 32'h42a107f0, 32'h42921b41, 32'hc255697a, 32'hc2815e5c, 32'h4256b1d0};
test_output[6001] = '{32'h42a107f0};
test_index[6001] = '{3};
test_input[48016:48023] = '{32'h427380e2, 32'hc2a61bff, 32'h42b29020, 32'hc27dcc80, 32'h429e573f, 32'hc2ad2dad, 32'h42b98f3b, 32'h42129353};
test_output[6002] = '{32'h42b98f3b};
test_index[6002] = '{6};
test_input[48024:48031] = '{32'hc0004235, 32'hc20243fc, 32'h41f4ec01, 32'hc2972f94, 32'h42877833, 32'hc275a95e, 32'hc27b627a, 32'hc1d203fd};
test_output[6003] = '{32'h42877833};
test_index[6003] = '{4};
test_input[48032:48039] = '{32'h426b66ec, 32'h42a66d9b, 32'h42850904, 32'hc23a9dab, 32'h42988bba, 32'h4293bf70, 32'h41fbef16, 32'hc1df4b67};
test_output[6004] = '{32'h42a66d9b};
test_index[6004] = '{1};
test_input[48040:48047] = '{32'hc255d5dd, 32'hc226fa89, 32'h42c327ee, 32'hc1192adb, 32'hc0a1256f, 32'h420a7060, 32'h41c8a3dd, 32'hc2bd5034};
test_output[6005] = '{32'h42c327ee};
test_index[6005] = '{2};
test_input[48048:48055] = '{32'h41cb04d1, 32'h41c19e18, 32'h424d4394, 32'hc1a30f51, 32'h41b15249, 32'h42b6cad3, 32'h420f9415, 32'hc2a8c65b};
test_output[6006] = '{32'h42b6cad3};
test_index[6006] = '{5};
test_input[48056:48063] = '{32'h41b11f12, 32'hc23b724c, 32'h41f3c353, 32'h419796f4, 32'h42b1d75f, 32'hc280aa08, 32'hc0bb22d7, 32'hc29fe9a5};
test_output[6007] = '{32'h42b1d75f};
test_index[6007] = '{4};
test_input[48064:48071] = '{32'hc17c9803, 32'hc1c481a3, 32'h420b48d3, 32'hc29b8552, 32'hc295c4ce, 32'hc2b00a39, 32'hc25d7574, 32'hc2bb6d74};
test_output[6008] = '{32'h420b48d3};
test_index[6008] = '{2};
test_input[48072:48079] = '{32'h4214ba5e, 32'hc13c8a8a, 32'h4299d50d, 32'hc2bab7da, 32'hc2298955, 32'h42324be6, 32'hc219bc5e, 32'hc2c365b2};
test_output[6009] = '{32'h4299d50d};
test_index[6009] = '{2};
test_input[48080:48087] = '{32'h412a7a18, 32'h428c8dcf, 32'h428b0aac, 32'h421bf064, 32'hc1bf6ae2, 32'hc10eb05a, 32'hc2894b3b, 32'h42201d58};
test_output[6010] = '{32'h428c8dcf};
test_index[6010] = '{1};
test_input[48088:48095] = '{32'h41b00176, 32'h420d0a8c, 32'hc2c365c7, 32'hc2a7ef39, 32'hc1324da5, 32'hc11bab27, 32'h41cf7bd3, 32'h4187962f};
test_output[6011] = '{32'h420d0a8c};
test_index[6011] = '{1};
test_input[48096:48103] = '{32'h42c0c2e9, 32'hc217110b, 32'hc2471102, 32'h42082624, 32'h42c0c9de, 32'hc2abb1c1, 32'h426ed55c, 32'h41c4d1fb};
test_output[6012] = '{32'h42c0c9de};
test_index[6012] = '{4};
test_input[48104:48111] = '{32'h41d7558c, 32'hc268f1d2, 32'h42c36428, 32'h41539947, 32'h4296ea33, 32'hc1fdafca, 32'hc2090aa7, 32'hc21caa18};
test_output[6013] = '{32'h42c36428};
test_index[6013] = '{2};
test_input[48112:48119] = '{32'h426b877f, 32'hc183c497, 32'hc0940624, 32'hc2bc6fb9, 32'h4246ecd3, 32'hc295a3ad, 32'h427c22f0, 32'hc23effa7};
test_output[6014] = '{32'h427c22f0};
test_index[6014] = '{6};
test_input[48120:48127] = '{32'h426327f7, 32'h42afa8cb, 32'h40bb70a8, 32'hc14a5f8a, 32'hc220389a, 32'h4078a505, 32'h42860d0e, 32'hbfd4ec54};
test_output[6015] = '{32'h42afa8cb};
test_index[6015] = '{1};
test_input[48128:48135] = '{32'h42c1b181, 32'h4199c370, 32'h42c08364, 32'hc213c130, 32'h42c59ce5, 32'hc0515900, 32'h41c4ca03, 32'h4256ebae};
test_output[6016] = '{32'h42c59ce5};
test_index[6016] = '{4};
test_input[48136:48143] = '{32'hc24046f8, 32'h40505f45, 32'h42b4e64c, 32'hc225ce41, 32'hc29f939c, 32'hc25cd706, 32'h40efd98e, 32'hc0fb7e2b};
test_output[6017] = '{32'h42b4e64c};
test_index[6017] = '{2};
test_input[48144:48151] = '{32'h42c00ffd, 32'h41f394fa, 32'h42a6370f, 32'h41d681f1, 32'hc1c5cb1b, 32'hc1c48c72, 32'h423948e7, 32'h41e26bca};
test_output[6018] = '{32'h42c00ffd};
test_index[6018] = '{0};
test_input[48152:48159] = '{32'hc266fcb9, 32'hc2bdb024, 32'hc0ddf52f, 32'hc2252341, 32'h428c0499, 32'hc2c3bba3, 32'h410eac39, 32'hc1f6e230};
test_output[6019] = '{32'h428c0499};
test_index[6019] = '{4};
test_input[48160:48167] = '{32'hc2a3dd36, 32'h4288df97, 32'h426fb03d, 32'hc260b2dd, 32'hc181214a, 32'hc1bed0be, 32'h42a8f80d, 32'h429bca56};
test_output[6020] = '{32'h42a8f80d};
test_index[6020] = '{6};
test_input[48168:48175] = '{32'hc1c21e22, 32'h4244aec2, 32'h42af692c, 32'h4272ca74, 32'hc20f0ad9, 32'hc003e978, 32'h417cc8b6, 32'h421075e8};
test_output[6021] = '{32'h42af692c};
test_index[6021] = '{2};
test_input[48176:48183] = '{32'h41ca6fa7, 32'hc2b67be9, 32'hc185b878, 32'hc153ef2d, 32'hc2c4e99e, 32'hbf86f7f6, 32'hc2191914, 32'hc22f184b};
test_output[6022] = '{32'h41ca6fa7};
test_index[6022] = '{0};
test_input[48184:48191] = '{32'h428e18f3, 32'h42bed660, 32'h41a38e87, 32'h4268c2a1, 32'h429b7035, 32'hc2036351, 32'hc2bcec80, 32'hc262e3de};
test_output[6023] = '{32'h42bed660};
test_index[6023] = '{1};
test_input[48192:48199] = '{32'h415fd7e0, 32'hc2a7f343, 32'hc1d0f42d, 32'hc2a0140f, 32'hc11da450, 32'h4224b4ea, 32'h3fbdbca4, 32'hc2491c1d};
test_output[6024] = '{32'h4224b4ea};
test_index[6024] = '{5};
test_input[48200:48207] = '{32'hc26eda10, 32'h40de2643, 32'hc208dc83, 32'hc1c1140a, 32'hc28ce135, 32'h41014c15, 32'h3d213a15, 32'hc2435965};
test_output[6025] = '{32'h41014c15};
test_index[6025] = '{5};
test_input[48208:48215] = '{32'h42968931, 32'h4134698c, 32'h40650da2, 32'hc296fd83, 32'hc22592a9, 32'h409bb116, 32'hc23aa31b, 32'h4296a6de};
test_output[6026] = '{32'h4296a6de};
test_index[6026] = '{7};
test_input[48216:48223] = '{32'h427812ac, 32'h42abbb17, 32'hc2882de5, 32'h41cea85d, 32'h42a03761, 32'hc28e2ca5, 32'hc29792de, 32'hc27ab2fe};
test_output[6027] = '{32'h42abbb17};
test_index[6027] = '{1};
test_input[48224:48231] = '{32'hc1465bb0, 32'h41f0db8f, 32'h427f8755, 32'hc2b8ee6a, 32'h418c253c, 32'h429bc36b, 32'h418ac216, 32'h426e9912};
test_output[6028] = '{32'h429bc36b};
test_index[6028] = '{5};
test_input[48232:48239] = '{32'hc25b056f, 32'hc2a8f5bd, 32'h426100f4, 32'h42a2a979, 32'hc23d84f5, 32'h42bf108b, 32'hc1ebe7c3, 32'h429fe081};
test_output[6029] = '{32'h42bf108b};
test_index[6029] = '{5};
test_input[48240:48247] = '{32'h426c68a2, 32'h4280be15, 32'hc2805195, 32'hc2c35198, 32'hc257dca9, 32'hc20a657c, 32'hc24de1d2, 32'h4250e98d};
test_output[6030] = '{32'h4280be15};
test_index[6030] = '{1};
test_input[48248:48255] = '{32'h42708396, 32'h41848541, 32'h42667506, 32'h41016ba6, 32'hc2337545, 32'hc0e32174, 32'hc231516c, 32'h42910ca0};
test_output[6031] = '{32'h42910ca0};
test_index[6031] = '{7};
test_input[48256:48263] = '{32'hc2a8272d, 32'hc296bfd0, 32'hc09ba25d, 32'h416e3fdc, 32'hc13aeb19, 32'h428b4d61, 32'h41f66e83, 32'h3ffb4455};
test_output[6032] = '{32'h428b4d61};
test_index[6032] = '{5};
test_input[48264:48271] = '{32'h4206842d, 32'hc275d50f, 32'h42ba0d30, 32'hc2b0d3da, 32'h423fd4d6, 32'h4246c139, 32'hc2be5edf, 32'h4285377f};
test_output[6033] = '{32'h42ba0d30};
test_index[6033] = '{2};
test_input[48272:48279] = '{32'hc1f9b375, 32'hc284d507, 32'h42354fdb, 32'hc2bf2180, 32'hc25fb4d5, 32'h4238af10, 32'h428035a4, 32'h41bda69e};
test_output[6034] = '{32'h428035a4};
test_index[6034] = '{6};
test_input[48280:48287] = '{32'h42a167dd, 32'hc24ef83f, 32'hc208cf78, 32'h41febfb8, 32'hc2348114, 32'h42bb0a92, 32'h41fa1b8e, 32'hc22085b4};
test_output[6035] = '{32'h42bb0a92};
test_index[6035] = '{5};
test_input[48288:48295] = '{32'hc29c4559, 32'h4282acdd, 32'h42a6c38d, 32'hc2ba38be, 32'hc2af62c9, 32'h422e1b33, 32'h429c89aa, 32'h423377c0};
test_output[6036] = '{32'h42a6c38d};
test_index[6036] = '{2};
test_input[48296:48303] = '{32'h429d2626, 32'hc2a32a31, 32'hc26b2597, 32'hc17e49fa, 32'h42943392, 32'h42c7d624, 32'h429aa741, 32'hc015643b};
test_output[6037] = '{32'h42c7d624};
test_index[6037] = '{5};
test_input[48304:48311] = '{32'h427ad174, 32'hc1c2e85d, 32'hc22576a4, 32'h42ac81e5, 32'h421745ab, 32'h420438c2, 32'hc21c969f, 32'h42049515};
test_output[6038] = '{32'h42ac81e5};
test_index[6038] = '{3};
test_input[48312:48319] = '{32'hc2a2884f, 32'hc21930f6, 32'h42aa3c74, 32'hc266bab0, 32'hc1d17cd7, 32'h42509afd, 32'hc20a94b8, 32'hc22604d0};
test_output[6039] = '{32'h42aa3c74};
test_index[6039] = '{2};
test_input[48320:48327] = '{32'h4220aaa4, 32'hc228b889, 32'h42226efc, 32'h429aff21, 32'hc204db0f, 32'hc29f4218, 32'h4202e83b, 32'hc27ec0a7};
test_output[6040] = '{32'h429aff21};
test_index[6040] = '{3};
test_input[48328:48335] = '{32'h42b40a6c, 32'h42a5cbca, 32'hc18ff643, 32'h425d4775, 32'hc2917818, 32'h42809baf, 32'hc2b2af71, 32'h42943c13};
test_output[6041] = '{32'h42b40a6c};
test_index[6041] = '{0};
test_input[48336:48343] = '{32'h406e2ede, 32'hc1c62325, 32'hc054962b, 32'h42b32f74, 32'h423d70e4, 32'h415e3eb2, 32'hc1b7aead, 32'hc24cbc79};
test_output[6042] = '{32'h42b32f74};
test_index[6042] = '{3};
test_input[48344:48351] = '{32'h4208f72e, 32'h42b2c1bb, 32'h42b7ff3e, 32'h4213d485, 32'h411649ab, 32'hc19a325b, 32'h41660539, 32'h4215a6ea};
test_output[6043] = '{32'h42b7ff3e};
test_index[6043] = '{2};
test_input[48352:48359] = '{32'hc2b97a93, 32'h42964158, 32'h4249625b, 32'h424462fe, 32'hc2c06419, 32'h4280c05e, 32'hc296b15f, 32'hc19cdbc1};
test_output[6044] = '{32'h42964158};
test_index[6044] = '{1};
test_input[48360:48367] = '{32'h4280f8d0, 32'hc2434951, 32'hc2117047, 32'h42a9fed4, 32'h42b16379, 32'h42af3cb8, 32'hc27d7025, 32'hc27000bf};
test_output[6045] = '{32'h42b16379};
test_index[6045] = '{4};
test_input[48368:48375] = '{32'hc228e467, 32'h42838ad0, 32'h4237eb4f, 32'hc0f63550, 32'hc263049e, 32'h422aade4, 32'hc2323544, 32'h42354734};
test_output[6046] = '{32'h42838ad0};
test_index[6046] = '{1};
test_input[48376:48383] = '{32'h42338f73, 32'h42927ef3, 32'h42add336, 32'h4261d4f0, 32'hc1d9d8bb, 32'hc2602c12, 32'h4229cc6f, 32'hc203c5a3};
test_output[6047] = '{32'h42add336};
test_index[6047] = '{2};
test_input[48384:48391] = '{32'h4299a2ca, 32'h4180074a, 32'h4211c3ae, 32'h41519bae, 32'hc28b8f8c, 32'h428be1ec, 32'h41f2b78c, 32'hc2bea3dd};
test_output[6048] = '{32'h4299a2ca};
test_index[6048] = '{0};
test_input[48392:48399] = '{32'h42a4aaec, 32'hc29fc050, 32'hc14da768, 32'hc1600b36, 32'hc29a0ad0, 32'hc28aa410, 32'h42bde325, 32'h420d3772};
test_output[6049] = '{32'h42bde325};
test_index[6049] = '{6};
test_input[48400:48407] = '{32'hc2bc3218, 32'h42af98bb, 32'hc2066e4d, 32'hc19b9223, 32'h42af650c, 32'h42be8099, 32'hc1137721, 32'hc1917591};
test_output[6050] = '{32'h42be8099};
test_index[6050] = '{5};
test_input[48408:48415] = '{32'h426a2b4b, 32'h42aeea55, 32'h421c70db, 32'h41d2fe2c, 32'hc28f7660, 32'h42631bfd, 32'hc2c5b074, 32'h420db3fe};
test_output[6051] = '{32'h42aeea55};
test_index[6051] = '{1};
test_input[48416:48423] = '{32'hc14dea76, 32'h428c90e1, 32'hc228c83e, 32'h42c673fd, 32'hc247d2e7, 32'h427e46c3, 32'hc269c10f, 32'h420d27c1};
test_output[6052] = '{32'h42c673fd};
test_index[6052] = '{3};
test_input[48424:48431] = '{32'hc1da5451, 32'h428b0acc, 32'hc0a5c295, 32'hc111fff6, 32'h42298732, 32'hc07784aa, 32'hc2a6efa4, 32'h40d5844a};
test_output[6053] = '{32'h428b0acc};
test_index[6053] = '{1};
test_input[48432:48439] = '{32'h42b3d789, 32'hc2bb5a13, 32'h424eeff9, 32'hc2865d45, 32'h42865ab5, 32'hc1d50713, 32'hc28d2161, 32'h4298a26d};
test_output[6054] = '{32'h42b3d789};
test_index[6054] = '{0};
test_input[48440:48447] = '{32'hc23cb497, 32'h42bb0305, 32'h423caf93, 32'hc1b35940, 32'h41d9a2bc, 32'h41cde5e1, 32'h420bcf53, 32'h42bfdae2};
test_output[6055] = '{32'h42bfdae2};
test_index[6055] = '{7};
test_input[48448:48455] = '{32'hc103fab3, 32'hc2a004da, 32'hc2200c16, 32'h421c59bf, 32'h428ca01e, 32'hc1c71103, 32'h4268c5fa, 32'hc280d1ec};
test_output[6056] = '{32'h428ca01e};
test_index[6056] = '{4};
test_input[48456:48463] = '{32'hc1696060, 32'hc2971792, 32'h42011c65, 32'hc26d6df9, 32'h42349d9c, 32'h414606ac, 32'h41be4ffa, 32'h42b99422};
test_output[6057] = '{32'h42b99422};
test_index[6057] = '{7};
test_input[48464:48471] = '{32'hc21a85a5, 32'h425bc3a3, 32'h410c8a57, 32'hc15cba37, 32'h42a314c2, 32'hc2826442, 32'hc2a7099f, 32'h41aae5ed};
test_output[6058] = '{32'h42a314c2};
test_index[6058] = '{4};
test_input[48472:48479] = '{32'hc2482225, 32'h42394dec, 32'hc24ff37c, 32'hc1868e33, 32'h411d47f4, 32'hc28e6ee1, 32'h412aa90a, 32'h40e16e78};
test_output[6059] = '{32'h42394dec};
test_index[6059] = '{1};
test_input[48480:48487] = '{32'h4229677d, 32'h42bccdea, 32'hc2246085, 32'h42ac5eea, 32'hc2a9098a, 32'hc28dbad0, 32'hc2bd49e8, 32'hc19b2ee4};
test_output[6060] = '{32'h42bccdea};
test_index[6060] = '{1};
test_input[48488:48495] = '{32'h42321c20, 32'h41806eca, 32'hc1b7d96e, 32'h4204acb7, 32'h424fa111, 32'h41beadd4, 32'hc2b84023, 32'h41bb77ed};
test_output[6061] = '{32'h424fa111};
test_index[6061] = '{4};
test_input[48496:48503] = '{32'hc146440d, 32'hc289be6b, 32'h41deb829, 32'hc2c53b50, 32'hc2786a9a, 32'hc2afa3b5, 32'h420119c7, 32'h42c772ff};
test_output[6062] = '{32'h42c772ff};
test_index[6062] = '{7};
test_input[48504:48511] = '{32'hc27ccbb7, 32'hc266f133, 32'hc121e9c0, 32'h4208ed13, 32'hc2bab2bc, 32'hc1bbeddf, 32'hc29ced79, 32'h42bfa5f2};
test_output[6063] = '{32'h42bfa5f2};
test_index[6063] = '{7};
test_input[48512:48519] = '{32'hc261a1c3, 32'h41870b7d, 32'h429e4bbd, 32'hc2abd569, 32'h42692a34, 32'hc2720b42, 32'h42a57525, 32'hc1be248f};
test_output[6064] = '{32'h42a57525};
test_index[6064] = '{6};
test_input[48520:48527] = '{32'hc14a99ee, 32'hc2420b89, 32'hc2c2949c, 32'h41e29a9a, 32'h42610aad, 32'h41d6bcaf, 32'hbf5093a9, 32'h42384c69};
test_output[6065] = '{32'h42610aad};
test_index[6065] = '{4};
test_input[48528:48535] = '{32'hc2002381, 32'hc2786f3c, 32'hc26d13ee, 32'h427643a3, 32'hc2b03ae0, 32'h42a276b9, 32'h4298e5a1, 32'h42accd50};
test_output[6066] = '{32'h42accd50};
test_index[6066] = '{7};
test_input[48536:48543] = '{32'h40abcc96, 32'h41a8718b, 32'h42bb0b4f, 32'h42331f91, 32'h420e2e6b, 32'hc29a5828, 32'h4297acda, 32'h4285ea47};
test_output[6067] = '{32'h42bb0b4f};
test_index[6067] = '{2};
test_input[48544:48551] = '{32'h4212136f, 32'hc12a715b, 32'hc2b1df18, 32'hc214950b, 32'hc2a9313f, 32'h420742e7, 32'h410e760a, 32'h42b349ec};
test_output[6068] = '{32'h42b349ec};
test_index[6068] = '{7};
test_input[48552:48559] = '{32'h4168da15, 32'hc0db8eef, 32'h425389d2, 32'h41bf2fa2, 32'h42a724d3, 32'hc2adf17d, 32'h426f2e3d, 32'h423bae17};
test_output[6069] = '{32'h42a724d3};
test_index[6069] = '{4};
test_input[48560:48567] = '{32'hc136ff52, 32'hc1da0acb, 32'h420d540b, 32'h429a7280, 32'hc2c49c97, 32'hc284e643, 32'h42120943, 32'h423b9765};
test_output[6070] = '{32'h429a7280};
test_index[6070] = '{3};
test_input[48568:48575] = '{32'h426ff5c5, 32'h41c86da0, 32'h42bc74d7, 32'hc27fb10c, 32'hc207aedb, 32'hc21a2bb0, 32'h427e1350, 32'h428cded5};
test_output[6071] = '{32'h42bc74d7};
test_index[6071] = '{2};
test_input[48576:48583] = '{32'hc2bbe92c, 32'h3ff234dc, 32'h426feb0b, 32'h426020ab, 32'h428984e9, 32'hc200bff2, 32'h41979fdf, 32'hc28a8c1a};
test_output[6072] = '{32'h428984e9};
test_index[6072] = '{4};
test_input[48584:48591] = '{32'h4297856a, 32'hc27bf77c, 32'h3efaf17f, 32'hc21a9a6c, 32'h4197d0ef, 32'h422baea9, 32'h429e08e1, 32'h42a76a93};
test_output[6073] = '{32'h42a76a93};
test_index[6073] = '{7};
test_input[48592:48599] = '{32'h42b8d814, 32'hc26e35e4, 32'h42b5e0c3, 32'hc0f339da, 32'hc23b0910, 32'h42ab32fe, 32'h42b78e86, 32'h42a6b67c};
test_output[6074] = '{32'h42b8d814};
test_index[6074] = '{0};
test_input[48600:48607] = '{32'hc29405de, 32'hc151f72c, 32'h41e72a2a, 32'hc0a9ad38, 32'h42a5bc5c, 32'hc2a1993a, 32'hc1cec499, 32'hc2a92026};
test_output[6075] = '{32'h42a5bc5c};
test_index[6075] = '{4};
test_input[48608:48615] = '{32'hbfc6a70f, 32'h42a4b777, 32'h41c5e8ac, 32'hc2173f4b, 32'h41405590, 32'h41de4d66, 32'hc2c17fe2, 32'hc184fe33};
test_output[6076] = '{32'h42a4b777};
test_index[6076] = '{1};
test_input[48616:48623] = '{32'h4063551b, 32'h41ac0bdb, 32'hc217b015, 32'hc2a94396, 32'h42582439, 32'h412212d6, 32'hc2bd5904, 32'h41e2a95d};
test_output[6077] = '{32'h42582439};
test_index[6077] = '{4};
test_input[48624:48631] = '{32'h42742cbc, 32'hc143db5c, 32'hc2af46fb, 32'h42890ec3, 32'hc2ad3007, 32'h4229677f, 32'hc28f8711, 32'h42723b90};
test_output[6078] = '{32'h42890ec3};
test_index[6078] = '{3};
test_input[48632:48639] = '{32'hc122e6ae, 32'hc2c3d32f, 32'h42b828ee, 32'hc10bc3c1, 32'hc250de33, 32'h428580f0, 32'h429679db, 32'h4221bb78};
test_output[6079] = '{32'h42b828ee};
test_index[6079] = '{2};
test_input[48640:48647] = '{32'h42b8c2ba, 32'hc2a58d49, 32'h41e3ec01, 32'hc1dc6de9, 32'h427f3431, 32'h42373864, 32'hc2bc7438, 32'h42ae067d};
test_output[6080] = '{32'h42b8c2ba};
test_index[6080] = '{0};
test_input[48648:48655] = '{32'hc18ae736, 32'hc252293f, 32'hc1b591fa, 32'h42c768e3, 32'h412952de, 32'hc1a99b1a, 32'h427e249c, 32'h426b2e3f};
test_output[6081] = '{32'h42c768e3};
test_index[6081] = '{3};
test_input[48656:48663] = '{32'hc2802ad1, 32'hc2548fa5, 32'h4100d3c4, 32'h4118c98f, 32'h4163413a, 32'h426e8e73, 32'hc236f216, 32'h4214cb42};
test_output[6082] = '{32'h426e8e73};
test_index[6082] = '{5};
test_input[48664:48671] = '{32'hc12dab8a, 32'hc256493c, 32'h409159a5, 32'hc2b06b56, 32'h411b9c8e, 32'h4215d2a8, 32'h42c27ce4, 32'hc2bdc63f};
test_output[6083] = '{32'h42c27ce4};
test_index[6083] = '{6};
test_input[48672:48679] = '{32'hbee865ce, 32'hc28646e7, 32'hc161a68f, 32'hc273c918, 32'hc1b3ee51, 32'hc28a94dd, 32'h41b088b3, 32'h428337ff};
test_output[6084] = '{32'h428337ff};
test_index[6084] = '{7};
test_input[48680:48687] = '{32'hc24cb26b, 32'h42b5936a, 32'hc278df40, 32'hc04b6aee, 32'h4285db4f, 32'hc18582f1, 32'h41c0d621, 32'hc0d619bd};
test_output[6085] = '{32'h42b5936a};
test_index[6085] = '{1};
test_input[48688:48695] = '{32'h42a5456b, 32'h425e1725, 32'hc22b29c0, 32'hc25692a8, 32'hc23373a3, 32'h4259d76c, 32'h426a948e, 32'h4241199c};
test_output[6086] = '{32'h42a5456b};
test_index[6086] = '{0};
test_input[48696:48703] = '{32'h4190c2f4, 32'h4223bd65, 32'h426132a7, 32'hc24dde85, 32'h427c86b8, 32'hc294bc78, 32'hc2828021, 32'h41595fb0};
test_output[6087] = '{32'h427c86b8};
test_index[6087] = '{4};
test_input[48704:48711] = '{32'hc2b14d04, 32'h42898805, 32'hc11a6c4f, 32'hc22c50f1, 32'h42311be0, 32'hc2aba303, 32'h42bb0ec4, 32'h41f2a254};
test_output[6088] = '{32'h42bb0ec4};
test_index[6088] = '{6};
test_input[48712:48719] = '{32'h41a5bc07, 32'h42757b19, 32'h4283bc8c, 32'h425db146, 32'h425855c2, 32'hc29268fd, 32'h428061cc, 32'h41d0d4cf};
test_output[6089] = '{32'h4283bc8c};
test_index[6089] = '{2};
test_input[48720:48727] = '{32'hc2800989, 32'hc0f313f3, 32'hc2bbbd2d, 32'h41179b41, 32'hc1323c2d, 32'h42a9d6f1, 32'h42a03f75, 32'h429e4fe0};
test_output[6090] = '{32'h42a9d6f1};
test_index[6090] = '{5};
test_input[48728:48735] = '{32'h42b976ab, 32'h429469cb, 32'hbf84e5b4, 32'h42502b0b, 32'hc260f05e, 32'hc1520be4, 32'h42581b29, 32'hc2335726};
test_output[6091] = '{32'h42b976ab};
test_index[6091] = '{0};
test_input[48736:48743] = '{32'h42282ff1, 32'h41854a05, 32'hc1b92e56, 32'h429f7a0c, 32'hc1a61600, 32'hc203a0ad, 32'hc22cb47c, 32'h421b9faa};
test_output[6092] = '{32'h429f7a0c};
test_index[6092] = '{3};
test_input[48744:48751] = '{32'h42a88fc6, 32'h421dba60, 32'hc23c8014, 32'hc262fe9e, 32'h4239d6a3, 32'hc1328f9d, 32'hc26e0981, 32'h429cbbd6};
test_output[6093] = '{32'h42a88fc6};
test_index[6093] = '{0};
test_input[48752:48759] = '{32'h42ab1f67, 32'hc240b175, 32'hc1d26b62, 32'hc292a2f5, 32'h41a78c89, 32'hc1500d4e, 32'hc2a38bc8, 32'hc1ca6d84};
test_output[6094] = '{32'h42ab1f67};
test_index[6094] = '{0};
test_input[48760:48767] = '{32'h42bf4019, 32'hc21f87d8, 32'hc23e6f8f, 32'h42a76230, 32'h41b65069, 32'h4242b0db, 32'h4264fccf, 32'hc2c7a965};
test_output[6095] = '{32'h42bf4019};
test_index[6095] = '{0};
test_input[48768:48775] = '{32'h42a7ceaa, 32'h4262d699, 32'h4285a6ce, 32'hc28c14fa, 32'hc1adecac, 32'hc2bf8acf, 32'hc252fc9e, 32'hc1c79dc0};
test_output[6096] = '{32'h42a7ceaa};
test_index[6096] = '{0};
test_input[48776:48783] = '{32'h428a8a42, 32'h42bcf910, 32'h426eba63, 32'h421b9807, 32'hc24a4be0, 32'h42a60d16, 32'h40ddd68a, 32'h412ecd72};
test_output[6097] = '{32'h42bcf910};
test_index[6097] = '{1};
test_input[48784:48791] = '{32'hc2acd114, 32'hc284f2f6, 32'h420cecc8, 32'hc2a49523, 32'hc1cdeda3, 32'hc1e024b7, 32'h420bd11a, 32'hc276f431};
test_output[6098] = '{32'h420cecc8};
test_index[6098] = '{2};
test_input[48792:48799] = '{32'hc1eecf6e, 32'hc26b414f, 32'hc243df97, 32'h419ab8b4, 32'h42a8a8d7, 32'hc2156bf8, 32'h40994712, 32'h411eed7f};
test_output[6099] = '{32'h42a8a8d7};
test_index[6099] = '{4};
test_input[48800:48807] = '{32'h41f1e8be, 32'h4294afac, 32'hc2b2fdab, 32'h426f147d, 32'hc1b3d290, 32'h412a668d, 32'hc2a45424, 32'hc29dbd7e};
test_output[6100] = '{32'h4294afac};
test_index[6100] = '{1};
test_input[48808:48815] = '{32'h42c481e2, 32'hc245c126, 32'h4207fb8c, 32'h42841dd2, 32'h4209c3b9, 32'h42180c1a, 32'hc2a12e2c, 32'h42ac1ad9};
test_output[6101] = '{32'h42c481e2};
test_index[6101] = '{0};
test_input[48816:48823] = '{32'h42617e3a, 32'h422633a1, 32'h42a0ec40, 32'h429193c1, 32'h413dafd3, 32'hc255b42f, 32'hc1a2bfea, 32'hc25726e7};
test_output[6102] = '{32'h42a0ec40};
test_index[6102] = '{2};
test_input[48824:48831] = '{32'h4280f7eb, 32'hc1f4433c, 32'h42ac1591, 32'h42afc166, 32'h42aacdf2, 32'h426d9a51, 32'h4295ca25, 32'hc2c4c3f1};
test_output[6103] = '{32'h42afc166};
test_index[6103] = '{3};
test_input[48832:48839] = '{32'hc24f87e4, 32'h41c89819, 32'h42bece13, 32'hc26e06b9, 32'hc236d6ce, 32'hc1a4ec28, 32'hc220166c, 32'hc293bc62};
test_output[6104] = '{32'h42bece13};
test_index[6104] = '{2};
test_input[48840:48847] = '{32'hc0b924c8, 32'h429820d3, 32'h40ae52ca, 32'h42b72220, 32'h42371ca6, 32'hc2841951, 32'h42991027, 32'h410704f2};
test_output[6105] = '{32'h42b72220};
test_index[6105] = '{3};
test_input[48848:48855] = '{32'hc1d2180e, 32'hc25abf8f, 32'hc27c5df5, 32'hc2176799, 32'h40caf95d, 32'h42024c61, 32'hc1d08045, 32'hc2663176};
test_output[6106] = '{32'h42024c61};
test_index[6106] = '{5};
test_input[48856:48863] = '{32'h42bb6be4, 32'h41740c2f, 32'h420bd08a, 32'h423da26d, 32'hc224645d, 32'h42201c95, 32'hc19da53a, 32'h425efbf3};
test_output[6107] = '{32'h42bb6be4};
test_index[6107] = '{0};
test_input[48864:48871] = '{32'hc0b3c1c3, 32'hc2272b3b, 32'hbfbfc8f7, 32'h4279de84, 32'hbf4f8d7e, 32'h3e10540d, 32'hc220fbd9, 32'hc25aea24};
test_output[6108] = '{32'h4279de84};
test_index[6108] = '{3};
test_input[48872:48879] = '{32'h42887ae2, 32'hc2910830, 32'h41a67f4c, 32'hc1671a85, 32'h422dc1f9, 32'h42ad21e1, 32'hc28bd13d, 32'h4264ec4a};
test_output[6109] = '{32'h42ad21e1};
test_index[6109] = '{5};
test_input[48880:48887] = '{32'hc24b59f7, 32'h42a49713, 32'hc280dcfc, 32'h4251b321, 32'h41208fd1, 32'h3fbb9c53, 32'h4142c4d0, 32'h42b116c7};
test_output[6110] = '{32'h42b116c7};
test_index[6110] = '{7};
test_input[48888:48895] = '{32'hc1944c76, 32'hc225673a, 32'h413e5675, 32'h42876209, 32'hc20b0a36, 32'h429cf3bd, 32'h415e8a33, 32'h422827a8};
test_output[6111] = '{32'h429cf3bd};
test_index[6111] = '{5};
test_input[48896:48903] = '{32'hc1985808, 32'hc20a736b, 32'h4282eabd, 32'h41dc678d, 32'h40be4c5e, 32'h423c22ea, 32'h42ade1df, 32'h405594bb};
test_output[6112] = '{32'h42ade1df};
test_index[6112] = '{6};
test_input[48904:48911] = '{32'h41a683e0, 32'hc0ff3403, 32'h42aae11a, 32'hc27ba0ab, 32'h411e9c13, 32'hc286a996, 32'h4278dc49, 32'h40cd5c3b};
test_output[6113] = '{32'h42aae11a};
test_index[6113] = '{2};
test_input[48912:48919] = '{32'h4299ab16, 32'h428882c6, 32'h40d9dd9e, 32'hc195c937, 32'h402af336, 32'hc13f5b7b, 32'h428c4b40, 32'h4295ef72};
test_output[6114] = '{32'h4299ab16};
test_index[6114] = '{0};
test_input[48920:48927] = '{32'hc2aafb1f, 32'hc21a36de, 32'h427e0f18, 32'hc2b38ca6, 32'h426240a2, 32'hc12dd35d, 32'hc0e12060, 32'hc2a986d3};
test_output[6115] = '{32'h427e0f18};
test_index[6115] = '{2};
test_input[48928:48935] = '{32'h42c54919, 32'h41953ace, 32'h429c2806, 32'hc23d42ad, 32'hc1d63be0, 32'hc2262dbb, 32'h4289197e, 32'hc1e656f7};
test_output[6116] = '{32'h42c54919};
test_index[6116] = '{0};
test_input[48936:48943] = '{32'hc2ab003f, 32'h42216c4a, 32'h4110b618, 32'h422b6202, 32'h420c3f03, 32'hc12bb3cd, 32'h428b8c8d, 32'h423bbddf};
test_output[6117] = '{32'h428b8c8d};
test_index[6117] = '{6};
test_input[48944:48951] = '{32'h42825b47, 32'hc29a3de9, 32'h41d5b7ad, 32'hc1c2aabc, 32'h42c4da2d, 32'h42970d99, 32'h429f7479, 32'hc29361e4};
test_output[6118] = '{32'h42c4da2d};
test_index[6118] = '{4};
test_input[48952:48959] = '{32'h42a73c87, 32'hc2b921e9, 32'hc2b88276, 32'hc2398065, 32'hc10f1a65, 32'h425e7c3d, 32'hc2bdb3ca, 32'h4242892f};
test_output[6119] = '{32'h42a73c87};
test_index[6119] = '{0};
test_input[48960:48967] = '{32'hc012ed5f, 32'hc28a804a, 32'hc245dde1, 32'h42a49aa2, 32'hc176dc36, 32'hc21a4cf1, 32'hc28f7f73, 32'h4292ea82};
test_output[6120] = '{32'h42a49aa2};
test_index[6120] = '{3};
test_input[48968:48975] = '{32'h424233dd, 32'h4192b257, 32'hc2558b0a, 32'h4249742e, 32'h42c212ff, 32'hc004ed05, 32'hc1dafc69, 32'h407abaf6};
test_output[6121] = '{32'h42c212ff};
test_index[6121] = '{4};
test_input[48976:48983] = '{32'h42a1c2b4, 32'hbf54f0b9, 32'hc0eb2102, 32'h4203032b, 32'hc2af7e2c, 32'h42b96c18, 32'h42c0169b, 32'hc25fcd90};
test_output[6122] = '{32'h42c0169b};
test_index[6122] = '{6};
test_input[48984:48991] = '{32'hc05b84c4, 32'hc1be3184, 32'hc2585c1b, 32'hc112aca7, 32'h423f34d6, 32'h424d4e63, 32'h42561b71, 32'hc100e631};
test_output[6123] = '{32'h42561b71};
test_index[6123] = '{6};
test_input[48992:48999] = '{32'hc0798000, 32'h40ecdfdc, 32'h42803106, 32'h421ec297, 32'h42577c31, 32'hc2982f5c, 32'hc1da0848, 32'hc2c0a3a8};
test_output[6124] = '{32'h42803106};
test_index[6124] = '{2};
test_input[49000:49007] = '{32'h4093f279, 32'hc25b5ab2, 32'h40a3129b, 32'hc2aa510f, 32'h3fb717d9, 32'hc19b3e1a, 32'h42c3aa26, 32'h4219505a};
test_output[6125] = '{32'h42c3aa26};
test_index[6125] = '{6};
test_input[49008:49015] = '{32'h40f200b6, 32'h42c2cdb8, 32'h4255002f, 32'h424ee0f6, 32'h42adb87a, 32'h4211d2f9, 32'hc1f6ff5c, 32'h424ba5c1};
test_output[6126] = '{32'h42c2cdb8};
test_index[6126] = '{1};
test_input[49016:49023] = '{32'h41d8e2c1, 32'h428564e6, 32'hc226eba3, 32'hc202247b, 32'hc2c0891e, 32'hc170a522, 32'h42370b3b, 32'hc26405e9};
test_output[6127] = '{32'h428564e6};
test_index[6127] = '{1};
test_input[49024:49031] = '{32'h4266f6e5, 32'hc21945a9, 32'h41833625, 32'hc23b766a, 32'h424f31b5, 32'h4257d96f, 32'hc2c68fce, 32'hbf15d491};
test_output[6128] = '{32'h4266f6e5};
test_index[6128] = '{0};
test_input[49032:49039] = '{32'h42005e82, 32'h42308ce0, 32'h415cc951, 32'h418d6d3d, 32'hc2768d96, 32'h41e56d5b, 32'hc20623bb, 32'hc28043aa};
test_output[6129] = '{32'h42308ce0};
test_index[6129] = '{1};
test_input[49040:49047] = '{32'hc1001541, 32'hc24fdd69, 32'hc0ef369a, 32'h428fd61d, 32'hc29b8c8e, 32'h4209e0d5, 32'hc2a87afb, 32'h429b6183};
test_output[6130] = '{32'h429b6183};
test_index[6130] = '{7};
test_input[49048:49055] = '{32'h42c72396, 32'h4230620c, 32'h42b364a0, 32'h415bef61, 32'h42b26395, 32'hc2bb0508, 32'h42a4af67, 32'h4219c6c3};
test_output[6131] = '{32'h42c72396};
test_index[6131] = '{0};
test_input[49056:49063] = '{32'hc108501d, 32'h42a0fa48, 32'h42383432, 32'hc1ed803c, 32'hc206ddd6, 32'hc2c5ea02, 32'h4167f7e6, 32'hc26c1d26};
test_output[6132] = '{32'h42a0fa48};
test_index[6132] = '{1};
test_input[49064:49071] = '{32'h42a096da, 32'h4262740a, 32'h403c76af, 32'h42564dcc, 32'h42797f5c, 32'hc2bfb9ac, 32'hc260c05e, 32'hc0c07bcd};
test_output[6133] = '{32'h42a096da};
test_index[6133] = '{0};
test_input[49072:49079] = '{32'hc271bfca, 32'h4231c8f9, 32'h41cc1b04, 32'hc21b4816, 32'hc200bf97, 32'h4256253a, 32'hc27a187f, 32'h428c4490};
test_output[6134] = '{32'h428c4490};
test_index[6134] = '{7};
test_input[49080:49087] = '{32'hc277ff0b, 32'h42b70dc8, 32'hc287fa4b, 32'hc2702385, 32'hc21c08fd, 32'hc25d3812, 32'h42027107, 32'hc19ee6dd};
test_output[6135] = '{32'h42b70dc8};
test_index[6135] = '{1};
test_input[49088:49095] = '{32'h4209a9b0, 32'hc154f88b, 32'hc2b92985, 32'h421f6170, 32'h42bc1349, 32'h424d824c, 32'hc1744526, 32'h41d05ab7};
test_output[6136] = '{32'h42bc1349};
test_index[6136] = '{4};
test_input[49096:49103] = '{32'h41576498, 32'hc0a78027, 32'hc2b9429f, 32'h4213bdb4, 32'h42777381, 32'hc1cd5b74, 32'hc238dbbb, 32'h423337fa};
test_output[6137] = '{32'h42777381};
test_index[6137] = '{4};
test_input[49104:49111] = '{32'hc22a70c0, 32'h42019def, 32'hc1d94478, 32'hc2982323, 32'hc1971156, 32'hc1934923, 32'h424385ab, 32'h4257ea30};
test_output[6138] = '{32'h4257ea30};
test_index[6138] = '{7};
test_input[49112:49119] = '{32'hc29d43a0, 32'h41ca419b, 32'h428a439a, 32'h42c51a2a, 32'h4235ee97, 32'h42bc38db, 32'h428d5d9c, 32'hc1eb0740};
test_output[6139] = '{32'h42c51a2a};
test_index[6139] = '{3};
test_input[49120:49127] = '{32'h42c4ff53, 32'h42b271df, 32'h41d3dc8d, 32'h417d4528, 32'hc2a9c035, 32'hc250f11a, 32'h41b09151, 32'hc269e107};
test_output[6140] = '{32'h42c4ff53};
test_index[6140] = '{0};
test_input[49128:49135] = '{32'h40673e4a, 32'hc2038210, 32'h4183a896, 32'h41a60396, 32'h4282d111, 32'hc22a81df, 32'h42b40d4f, 32'h426d8bf9};
test_output[6141] = '{32'h42b40d4f};
test_index[6141] = '{6};
test_input[49136:49143] = '{32'hc1859fea, 32'h42bef95d, 32'hc294bc37, 32'hc275b857, 32'hc2a68237, 32'h424496c1, 32'hc20ce2c0, 32'h4222df04};
test_output[6142] = '{32'h42bef95d};
test_index[6142] = '{1};
test_input[49144:49151] = '{32'hc2ab89b1, 32'h4269b7ba, 32'hc293b507, 32'h42a90222, 32'hc1c23bee, 32'h41809f16, 32'hc27c26cd, 32'h42bf150b};
test_output[6143] = '{32'h42bf150b};
test_index[6143] = '{7};
test_input[49152:49159] = '{32'h429b8993, 32'hc209133d, 32'h4005409b, 32'hc2ae4d93, 32'h4215555f, 32'h425383b9, 32'h411fe985, 32'h4188dc90};
test_output[6144] = '{32'h429b8993};
test_index[6144] = '{0};
test_input[49160:49167] = '{32'h42beeb09, 32'hc269e6d9, 32'h42126a37, 32'h42bc5ad0, 32'h423dd426, 32'hc2975b89, 32'hc27ee580, 32'h4239d4ee};
test_output[6145] = '{32'h42beeb09};
test_index[6145] = '{0};
test_input[49168:49175] = '{32'hc1c75bc2, 32'hc2467194, 32'h42aba0e2, 32'h428c9d44, 32'h406fb2da, 32'h41800c9a, 32'hc29a50a9, 32'h41581247};
test_output[6146] = '{32'h42aba0e2};
test_index[6146] = '{2};
test_input[49176:49183] = '{32'h41cbc8ae, 32'hc28f8af9, 32'h428064e7, 32'h425b27b0, 32'h42afc03d, 32'h423ad939, 32'h42bb73e2, 32'h42060bf5};
test_output[6147] = '{32'h42bb73e2};
test_index[6147] = '{6};
test_input[49184:49191] = '{32'hc2ba50a8, 32'h428cc9ae, 32'h425f98cc, 32'hc2b55c8b, 32'h423fc34f, 32'h427241e1, 32'h4281cde4, 32'hc284c598};
test_output[6148] = '{32'h428cc9ae};
test_index[6148] = '{1};
test_input[49192:49199] = '{32'hc2ae3dc8, 32'h41d8d0ba, 32'h42139616, 32'hc2a6a0e9, 32'h424dd1a1, 32'h417861c2, 32'hc2990901, 32'hc2076c95};
test_output[6149] = '{32'h424dd1a1};
test_index[6149] = '{4};
test_input[49200:49207] = '{32'h42be9856, 32'h4199cfd3, 32'h403e584e, 32'h42afc932, 32'h413a3140, 32'h422a31bb, 32'hc120a843, 32'h42ac735e};
test_output[6150] = '{32'h42be9856};
test_index[6150] = '{0};
test_input[49208:49215] = '{32'h4266f017, 32'h42b9dafb, 32'h4156d906, 32'hc20d4273, 32'hc2848403, 32'hc1aecdfd, 32'hc214e5c7, 32'hc1f336a3};
test_output[6151] = '{32'h42b9dafb};
test_index[6151] = '{1};
test_input[49216:49223] = '{32'h42536313, 32'hc28de053, 32'hc0838b8a, 32'h414c0921, 32'h42a1779c, 32'h41f77f6a, 32'h3e95063c, 32'h42536dc2};
test_output[6152] = '{32'h42a1779c};
test_index[6152] = '{4};
test_input[49224:49231] = '{32'h4166b7e2, 32'h40e8583f, 32'h428dbf1a, 32'h42a86be3, 32'hc00308a0, 32'h42883574, 32'hc1fef27a, 32'h40e0da18};
test_output[6153] = '{32'h42a86be3};
test_index[6153] = '{3};
test_input[49232:49239] = '{32'hc2428bba, 32'hc24957af, 32'hc254a69f, 32'hc27c5687, 32'h42a33a2b, 32'hc2518015, 32'hc274824d, 32'h42788c2e};
test_output[6154] = '{32'h42a33a2b};
test_index[6154] = '{4};
test_input[49240:49247] = '{32'h428368dc, 32'hc2847a0d, 32'hc28d2e25, 32'h41d22187, 32'hc2c329dc, 32'hbede694e, 32'hc2ac9d91, 32'h429b8b72};
test_output[6155] = '{32'h429b8b72};
test_index[6155] = '{7};
test_input[49248:49255] = '{32'h4200f935, 32'hc22f44d9, 32'h42876874, 32'h4179c15f, 32'hc22f7f3c, 32'hc28215e8, 32'h420b67d9, 32'hc2b8b458};
test_output[6156] = '{32'h42876874};
test_index[6156] = '{2};
test_input[49256:49263] = '{32'hc222be41, 32'hc221f668, 32'h42144d7e, 32'hc123216d, 32'h429a27fa, 32'h41996fd5, 32'h41059007, 32'hc1b80021};
test_output[6157] = '{32'h429a27fa};
test_index[6157] = '{4};
test_input[49264:49271] = '{32'hc28177ae, 32'h420c723a, 32'h4210b00e, 32'hc293a583, 32'hc2a3aff8, 32'h4198468a, 32'h42b70453, 32'hc2a08af9};
test_output[6158] = '{32'h42b70453};
test_index[6158] = '{6};
test_input[49272:49279] = '{32'h42ba115f, 32'h42acf228, 32'h4204444f, 32'hc2b7436e, 32'hc19ed33c, 32'h41f23b84, 32'h42043797, 32'hc2ad438b};
test_output[6159] = '{32'h42ba115f};
test_index[6159] = '{0};
test_input[49280:49287] = '{32'hc2c7fd86, 32'hc2aaf5c4, 32'hc2bdbdf9, 32'h429e919c, 32'hc275efd8, 32'h42831870, 32'h41a440c2, 32'h4207ee9d};
test_output[6160] = '{32'h429e919c};
test_index[6160] = '{3};
test_input[49288:49295] = '{32'h417f7500, 32'hc269f7ce, 32'hc1bfb889, 32'h428c02f9, 32'h4224bbf2, 32'hc2a28066, 32'h42c6b7f2, 32'h42305502};
test_output[6161] = '{32'h42c6b7f2};
test_index[6161] = '{6};
test_input[49296:49303] = '{32'h42c45ebd, 32'hc27c498a, 32'hc2c04f47, 32'hc231096d, 32'hc19e93c0, 32'h42625fd4, 32'h414dcd7b, 32'h4287a975};
test_output[6162] = '{32'h42c45ebd};
test_index[6162] = '{0};
test_input[49304:49311] = '{32'hc2b590f7, 32'hc262aa2a, 32'hbff1cea7, 32'h419f427f, 32'hc202e5a7, 32'h426aa877, 32'hc2a80c0f, 32'hc2437c48};
test_output[6163] = '{32'h426aa877};
test_index[6163] = '{5};
test_input[49312:49319] = '{32'h41789dbd, 32'h42471dc8, 32'h402452aa, 32'h41e181fa, 32'hc2c442f9, 32'h414b598d, 32'hc2abf221, 32'hc20324e2};
test_output[6164] = '{32'h42471dc8};
test_index[6164] = '{1};
test_input[49320:49327] = '{32'h42b39993, 32'h4193dc8e, 32'h412bb6f3, 32'h4292c6c9, 32'h42bc15e9, 32'hc21fd0fd, 32'hc25666fd, 32'hc0b20a32};
test_output[6165] = '{32'h42bc15e9};
test_index[6165] = '{4};
test_input[49328:49335] = '{32'hc2a70472, 32'hc1e843fa, 32'hc1f30466, 32'h41570727, 32'h4293d40c, 32'hc2283962, 32'hc1e04772, 32'h429ef59f};
test_output[6166] = '{32'h429ef59f};
test_index[6166] = '{7};
test_input[49336:49343] = '{32'hc1b7d927, 32'hc1eaab3d, 32'h40eb2714, 32'hbea69c56, 32'hbfb51d3a, 32'h4244b64f, 32'h41dc7bf2, 32'h4255e50e};
test_output[6167] = '{32'h4255e50e};
test_index[6167] = '{7};
test_input[49344:49351] = '{32'hc1f47ad1, 32'h428cedb0, 32'hc2c4898a, 32'hc17022f3, 32'hc0a610d6, 32'h42354c12, 32'hc183f901, 32'hc282e5b6};
test_output[6168] = '{32'h428cedb0};
test_index[6168] = '{1};
test_input[49352:49359] = '{32'hc0c7dd92, 32'h42963401, 32'hc1c81c23, 32'h42a030ec, 32'h420b2f19, 32'hc295e3b9, 32'h41292ccc, 32'h411f1e2f};
test_output[6169] = '{32'h42a030ec};
test_index[6169] = '{3};
test_input[49360:49367] = '{32'h42c7fc3a, 32'hc1dd2c57, 32'h42a7eed4, 32'h41f90f9b, 32'h4292d81f, 32'h427a69c8, 32'hbf67725e, 32'hc286bd60};
test_output[6170] = '{32'h42c7fc3a};
test_index[6170] = '{0};
test_input[49368:49375] = '{32'h4284d4d8, 32'hc23fbfde, 32'hc244de96, 32'hc211e9ce, 32'h4294d3e6, 32'hc2292ab4, 32'hc28fe9e2, 32'hc2111223};
test_output[6171] = '{32'h4294d3e6};
test_index[6171] = '{4};
test_input[49376:49383] = '{32'hc24c9c19, 32'hc2b9da9a, 32'h4155469c, 32'hc1c0b0c5, 32'h403eaa63, 32'hc22c6616, 32'hc226c320, 32'hc2bdd4d2};
test_output[6172] = '{32'h4155469c};
test_index[6172] = '{2};
test_input[49384:49391] = '{32'hc1dc7d5e, 32'hc245ca1a, 32'h42141bfe, 32'hc1bbe9b0, 32'hc1dc189f, 32'hc22ec9e4, 32'h4228bab3, 32'hc18595bd};
test_output[6173] = '{32'h4228bab3};
test_index[6173] = '{6};
test_input[49392:49399] = '{32'h42443503, 32'h42c46063, 32'h42b529a0, 32'hc24f7779, 32'h41e944ce, 32'hc29e20c7, 32'h42094005, 32'h41e10cb8};
test_output[6174] = '{32'h42c46063};
test_index[6174] = '{1};
test_input[49400:49407] = '{32'h40ca76a1, 32'h4181d61d, 32'hc2c2927d, 32'hc1a61451, 32'h41329e9f, 32'h42850642, 32'h420ed8ed, 32'hc2a79820};
test_output[6175] = '{32'h42850642};
test_index[6175] = '{5};
test_input[49408:49415] = '{32'h4166602f, 32'hc29c1918, 32'h4298ed8e, 32'hc29ccdf0, 32'hc1d0c217, 32'h41ffb97a, 32'hc2b3bd21, 32'hc1bc3b3c};
test_output[6176] = '{32'h4298ed8e};
test_index[6176] = '{2};
test_input[49416:49423] = '{32'hc25573c7, 32'h42541bcb, 32'h4268e6f1, 32'h422182a9, 32'h42941c17, 32'h428c687f, 32'hc21fa5ec, 32'h41b907d9};
test_output[6177] = '{32'h42941c17};
test_index[6177] = '{4};
test_input[49424:49431] = '{32'hc215a91b, 32'hc29df8ca, 32'hc237fa4b, 32'hc1004913, 32'hc2abcbb7, 32'h40a386f1, 32'hc13b1dc7, 32'h426e8532};
test_output[6178] = '{32'h426e8532};
test_index[6178] = '{7};
test_input[49432:49439] = '{32'h40b49b77, 32'hc183bb2a, 32'h429f9aca, 32'hc099fd83, 32'hc1adeddc, 32'h42b11494, 32'hc2059ea0, 32'hc2c3dacd};
test_output[6179] = '{32'h42b11494};
test_index[6179] = '{5};
test_input[49440:49447] = '{32'h4072a805, 32'h4012bc39, 32'h4201ed15, 32'hc25b4a22, 32'hc11dbd6b, 32'hc2c4b49c, 32'h429b7bfa, 32'hc204318f};
test_output[6180] = '{32'h429b7bfa};
test_index[6180] = '{6};
test_input[49448:49455] = '{32'hc1ebb83d, 32'hc2995562, 32'hc1c079c1, 32'h426cacff, 32'hc266a1ed, 32'hc2c159c0, 32'h42c6db12, 32'hc2956731};
test_output[6181] = '{32'h42c6db12};
test_index[6181] = '{6};
test_input[49456:49463] = '{32'h41eb997d, 32'hc149d492, 32'h424db482, 32'hc1784c0f, 32'h413f623b, 32'h42a87be7, 32'hc2c4aba3, 32'hc2806f26};
test_output[6182] = '{32'h42a87be7};
test_index[6182] = '{5};
test_input[49464:49471] = '{32'h428ce8dc, 32'hc1930b10, 32'h3fb4a776, 32'h4245da04, 32'hc256017f, 32'hc268846b, 32'h421fbcda, 32'h4236096e};
test_output[6183] = '{32'h428ce8dc};
test_index[6183] = '{0};
test_input[49472:49479] = '{32'hc2411111, 32'hc23a1652, 32'h412fe554, 32'h42b9a714, 32'hc20f8bbc, 32'hc1d7ce89, 32'hc2a77b09, 32'hc22b814b};
test_output[6184] = '{32'h42b9a714};
test_index[6184] = '{3};
test_input[49480:49487] = '{32'h42071811, 32'hc19eccd1, 32'hc2bd8d6d, 32'h42af1e0e, 32'h425d28d2, 32'hc2305a6d, 32'hc2207bb1, 32'h42356d4a};
test_output[6185] = '{32'h42af1e0e};
test_index[6185] = '{3};
test_input[49488:49495] = '{32'hc2a69c36, 32'hc20c9c54, 32'h41a4b9de, 32'hc1e795b6, 32'h4252a780, 32'h4128c682, 32'h425e1e06, 32'h4243e424};
test_output[6186] = '{32'h425e1e06};
test_index[6186] = '{6};
test_input[49496:49503] = '{32'h4214a0a2, 32'hc28f788f, 32'h426ca4f1, 32'h429ea73f, 32'hc1b78802, 32'h42888052, 32'hc2945ef0, 32'h4290b6d2};
test_output[6187] = '{32'h429ea73f};
test_index[6187] = '{3};
test_input[49504:49511] = '{32'hc29c8bec, 32'h4181e03c, 32'hc231683f, 32'h4282b225, 32'h428af0e0, 32'hc26b41a2, 32'hc284b182, 32'h42a60fb8};
test_output[6188] = '{32'h42a60fb8};
test_index[6188] = '{7};
test_input[49512:49519] = '{32'hc03cd80e, 32'h42590301, 32'h41fb4209, 32'hc265e8df, 32'h42990ade, 32'hc203b3ee, 32'h41a84530, 32'h429e6767};
test_output[6189] = '{32'h429e6767};
test_index[6189] = '{7};
test_input[49520:49527] = '{32'hc286f357, 32'hc23aca4e, 32'h40dc66b2, 32'hc2c6a88e, 32'hc27af563, 32'hc127b250, 32'h423e6ad5, 32'h3fb24327};
test_output[6190] = '{32'h423e6ad5};
test_index[6190] = '{6};
test_input[49528:49535] = '{32'h42b27ad8, 32'hc2c2dfda, 32'h42b9c04f, 32'hc1d14edb, 32'h427e6d79, 32'h41c9ea9c, 32'hc206a079, 32'hc2b8998e};
test_output[6191] = '{32'h42b9c04f};
test_index[6191] = '{2};
test_input[49536:49543] = '{32'hc2431ec9, 32'hc2a92bbd, 32'hc0ec9a9f, 32'hc216062c, 32'h42ad819a, 32'hc2a6c60e, 32'h4201092c, 32'h4293992b};
test_output[6192] = '{32'h42ad819a};
test_index[6192] = '{4};
test_input[49544:49551] = '{32'hc21625f9, 32'hc27f074b, 32'hc2b03813, 32'h41b979cb, 32'hc184010a, 32'hc1f93688, 32'h429b037e, 32'h425b598c};
test_output[6193] = '{32'h429b037e};
test_index[6193] = '{6};
test_input[49552:49559] = '{32'hc247f506, 32'h4291694a, 32'h42245a8d, 32'hc1b64bad, 32'h41a4a8ff, 32'hc1fb708c, 32'h42463a66, 32'h42c60036};
test_output[6194] = '{32'h42c60036};
test_index[6194] = '{7};
test_input[49560:49567] = '{32'h42a49acf, 32'h426aad8f, 32'hc2873f7e, 32'hc1f88962, 32'hc1f60cdf, 32'hc1d8def3, 32'h428841c8, 32'hc0b5a038};
test_output[6195] = '{32'h42a49acf};
test_index[6195] = '{0};
test_input[49568:49575] = '{32'h42569575, 32'h4150b0c6, 32'hc20d607f, 32'h413059af, 32'hc20422a4, 32'h428bfbc7, 32'h42b35400, 32'hc232ffbe};
test_output[6196] = '{32'h42b35400};
test_index[6196] = '{6};
test_input[49576:49583] = '{32'hc296545c, 32'hc1f2199b, 32'h42358f24, 32'hc28b0bd4, 32'hc2044c6b, 32'hc2408146, 32'h421350e4, 32'h42a625b4};
test_output[6197] = '{32'h42a625b4};
test_index[6197] = '{7};
test_input[49584:49591] = '{32'hc23b4fb9, 32'hc1baf530, 32'h42c1ce13, 32'hc2c74c52, 32'hc241b000, 32'hc2190451, 32'hc2980ee7, 32'h4287a7b2};
test_output[6198] = '{32'h42c1ce13};
test_index[6198] = '{2};
test_input[49592:49599] = '{32'h42afe096, 32'hc2bcdf79, 32'hc294dd28, 32'h42442ec0, 32'hc286e874, 32'hc1ca90c7, 32'hc245dd64, 32'hc21aae98};
test_output[6199] = '{32'h42afe096};
test_index[6199] = '{0};
test_input[49600:49607] = '{32'h42b7e594, 32'h42023f52, 32'h41c27573, 32'h4222543c, 32'h428ebf91, 32'h42b413c5, 32'hc2bab054, 32'h42aeb80f};
test_output[6200] = '{32'h42b7e594};
test_index[6200] = '{0};
test_input[49608:49615] = '{32'hc2135f87, 32'hc236c44e, 32'hc24b58ac, 32'hc295a281, 32'hc1a13b2b, 32'hc1e5562f, 32'hc204f785, 32'h42100774};
test_output[6201] = '{32'h42100774};
test_index[6201] = '{7};
test_input[49616:49623] = '{32'hc213f3dd, 32'hc2839b4b, 32'h426e43a7, 32'hc28ac169, 32'hc2b20c40, 32'h42902cdd, 32'h41f599fd, 32'hc109e1f0};
test_output[6202] = '{32'h42902cdd};
test_index[6202] = '{5};
test_input[49624:49631] = '{32'hc1f0c1b4, 32'hc251b763, 32'h42372bbc, 32'hc238fd1a, 32'hc20f6975, 32'hc0b93139, 32'h41eee187, 32'h42496d4c};
test_output[6203] = '{32'h42496d4c};
test_index[6203] = '{7};
test_input[49632:49639] = '{32'hc265b817, 32'hc2942c35, 32'h428fc915, 32'hc212fc74, 32'h42965052, 32'hc278368d, 32'h42b62b1f, 32'hc1d6d050};
test_output[6204] = '{32'h42b62b1f};
test_index[6204] = '{6};
test_input[49640:49647] = '{32'hc2030a8c, 32'h427979f7, 32'hc17c5530, 32'hc1fb82e2, 32'h425c736a, 32'h42a62e17, 32'hc287df7b, 32'h4214ecdf};
test_output[6205] = '{32'h42a62e17};
test_index[6205] = '{5};
test_input[49648:49655] = '{32'h427ed50b, 32'hc2a015c5, 32'h420e8f78, 32'h41fd38b1, 32'hc209ea74, 32'h41df8639, 32'h402340b6, 32'hc1cd4496};
test_output[6206] = '{32'h427ed50b};
test_index[6206] = '{0};
test_input[49656:49663] = '{32'hc2a5ace0, 32'h4198ed2c, 32'hc2a131d4, 32'hc0b8e934, 32'h408d4e1b, 32'h4208b7b8, 32'hc282085d, 32'hc29713c9};
test_output[6207] = '{32'h4208b7b8};
test_index[6207] = '{5};
test_input[49664:49671] = '{32'h42b4b0d7, 32'h42778f3c, 32'hc2b55204, 32'hc162013b, 32'hc2b7bbe7, 32'h426003ce, 32'hc23091ec, 32'hc1a775ab};
test_output[6208] = '{32'h42b4b0d7};
test_index[6208] = '{0};
test_input[49672:49679] = '{32'h421f7812, 32'h4270478c, 32'hc2874e78, 32'h4250a318, 32'h41175baf, 32'hc1a32f90, 32'hc2a69cad, 32'hc25812b0};
test_output[6209] = '{32'h4270478c};
test_index[6209] = '{1};
test_input[49680:49687] = '{32'hc2a73677, 32'h42b7a8c7, 32'h424f0fe5, 32'h423b4324, 32'hc29cab35, 32'hc2868387, 32'hc20e1229, 32'hbe4b0dbe};
test_output[6210] = '{32'h42b7a8c7};
test_index[6210] = '{1};
test_input[49688:49695] = '{32'h42535c7a, 32'hc20afed2, 32'hc1823376, 32'hc2a1da23, 32'h40d68e92, 32'hc2bea10a, 32'h429df37a, 32'h42c02ec7};
test_output[6211] = '{32'h42c02ec7};
test_index[6211] = '{7};
test_input[49696:49703] = '{32'hc13c90ec, 32'h42a344c6, 32'hc2809d62, 32'h427f116d, 32'hc21d45b4, 32'h411819e2, 32'hc0e23ff5, 32'hc1e8dd10};
test_output[6212] = '{32'h42a344c6};
test_index[6212] = '{1};
test_input[49704:49711] = '{32'hc1d41f94, 32'hc1de571b, 32'hc11fe6a8, 32'h42948a31, 32'hc1917103, 32'hc1b7f5b8, 32'hc2c6386a, 32'hc2297dc9};
test_output[6213] = '{32'h42948a31};
test_index[6213] = '{3};
test_input[49712:49719] = '{32'h427482d0, 32'h4141f56e, 32'h40b64009, 32'h42250920, 32'hc1b4415c, 32'hc2b566ea, 32'h42c70e74, 32'hc26cb455};
test_output[6214] = '{32'h42c70e74};
test_index[6214] = '{6};
test_input[49720:49727] = '{32'hc24bf677, 32'hc2bd1ac6, 32'hc2720382, 32'h40baf178, 32'hc17de77b, 32'hc131d133, 32'h422083fb, 32'h41a32f4c};
test_output[6215] = '{32'h422083fb};
test_index[6215] = '{6};
test_input[49728:49735] = '{32'h42809ad1, 32'hc22d39c2, 32'h427dace1, 32'h3f6cba48, 32'h4241c9fc, 32'h429ac29a, 32'h42c44388, 32'h4294a9b4};
test_output[6216] = '{32'h42c44388};
test_index[6216] = '{6};
test_input[49736:49743] = '{32'hc28f7f77, 32'hc2c2b7f0, 32'h417a89bd, 32'hc2a28266, 32'h41b6aafc, 32'hc222350b, 32'h4284d09d, 32'h42969b5a};
test_output[6217] = '{32'h42969b5a};
test_index[6217] = '{7};
test_input[49744:49751] = '{32'hc2c6ed15, 32'h42aeefcf, 32'hc2473295, 32'hc29423d9, 32'h4286f694, 32'h410c4b15, 32'h42b6474e, 32'h42b3eb41};
test_output[6218] = '{32'h42b6474e};
test_index[6218] = '{6};
test_input[49752:49759] = '{32'h42468939, 32'h425e7ddf, 32'h425684f7, 32'hc10ccb54, 32'hc20e7a07, 32'hc168c3aa, 32'h407f10f6, 32'hc23cbfa3};
test_output[6219] = '{32'h425e7ddf};
test_index[6219] = '{1};
test_input[49760:49767] = '{32'h41e6efa3, 32'h42afbd48, 32'hc088e218, 32'h428090a7, 32'hc225ab06, 32'h4298eea6, 32'hc2028788, 32'hc165852b};
test_output[6220] = '{32'h42afbd48};
test_index[6220] = '{1};
test_input[49768:49775] = '{32'hc1b2b0f9, 32'h423d6285, 32'hc259215b, 32'h420bf7ad, 32'hc2898bb5, 32'h4281cf5b, 32'h429c8180, 32'h41c25eae};
test_output[6221] = '{32'h429c8180};
test_index[6221] = '{6};
test_input[49776:49783] = '{32'h41405ac0, 32'hc287d8db, 32'h42843786, 32'hc2a6aabd, 32'h41cb5cb6, 32'h42c5ebfd, 32'hc25b7121, 32'hc18eac39};
test_output[6222] = '{32'h42c5ebfd};
test_index[6222] = '{5};
test_input[49784:49791] = '{32'hc272972e, 32'hc28fa71f, 32'h428009fd, 32'hc15f69b7, 32'h404301e6, 32'h41764ba3, 32'hc181572f, 32'hc20f4470};
test_output[6223] = '{32'h428009fd};
test_index[6223] = '{2};
test_input[49792:49799] = '{32'h4285e582, 32'h428eb278, 32'hc20e2f90, 32'h42a5f69f, 32'h426bfe1e, 32'hc2a15408, 32'h429ffc3c, 32'hc1804d41};
test_output[6224] = '{32'h42a5f69f};
test_index[6224] = '{3};
test_input[49800:49807] = '{32'hc21a3bc9, 32'hc29a1d2c, 32'hc26eb7c3, 32'hc220bc6d, 32'h423e24e0, 32'hc28d76f6, 32'h40f1c6f4, 32'hc21dd258};
test_output[6225] = '{32'h423e24e0};
test_index[6225] = '{4};
test_input[49808:49815] = '{32'hc2bc4460, 32'hc11b3b4f, 32'h41dbd46f, 32'h4228a41d, 32'h42b47009, 32'h40e1976d, 32'h3f89d7fa, 32'h41e9e104};
test_output[6226] = '{32'h42b47009};
test_index[6226] = '{4};
test_input[49816:49823] = '{32'h4219e861, 32'h42ad3c52, 32'h428f0692, 32'h42bcd073, 32'hc2bed66f, 32'h426d9f31, 32'h42aa31f1, 32'hc2c0e16d};
test_output[6227] = '{32'h42bcd073};
test_index[6227] = '{3};
test_input[49824:49831] = '{32'h42ab9db6, 32'h4123f051, 32'hc2853e79, 32'h42ba1b2e, 32'hc164e511, 32'h42a8a419, 32'hc118667b, 32'h4209d73b};
test_output[6228] = '{32'h42ba1b2e};
test_index[6228] = '{3};
test_input[49832:49839] = '{32'h41aed838, 32'hc1b16309, 32'h42b63cef, 32'h41a40782, 32'hc1cdfa11, 32'hc22f17e5, 32'hc1e71cb3, 32'hc264b42d};
test_output[6229] = '{32'h42b63cef};
test_index[6229] = '{2};
test_input[49840:49847] = '{32'hc27a01d6, 32'hc2c0b4ef, 32'h421262b7, 32'hc1963fa8, 32'h42c72c4b, 32'h425f9730, 32'h42878b85, 32'h4271cf7e};
test_output[6230] = '{32'h42c72c4b};
test_index[6230] = '{4};
test_input[49848:49855] = '{32'h415d68ab, 32'h407a2d96, 32'h42873680, 32'h424f667d, 32'h42c5e7ab, 32'h4243495b, 32'h4239c563, 32'hc265cb34};
test_output[6231] = '{32'h42c5e7ab};
test_index[6231] = '{4};
test_input[49856:49863] = '{32'h418a40c0, 32'hc1385ccb, 32'h41955ed0, 32'hc236b57b, 32'hc281d2b1, 32'h413ac933, 32'h423e5a0c, 32'hc284b810};
test_output[6232] = '{32'h423e5a0c};
test_index[6232] = '{6};
test_input[49864:49871] = '{32'hc126eb68, 32'h416b17e6, 32'hbeda2e96, 32'h410b8669, 32'h4195310c, 32'hc1e60d94, 32'hc28649fd, 32'hc2a445b7};
test_output[6233] = '{32'h4195310c};
test_index[6233] = '{4};
test_input[49872:49879] = '{32'h412d6094, 32'hc27f7349, 32'hc0ae3358, 32'h414e9208, 32'hc01005dc, 32'h42491356, 32'hc294a93e, 32'h412f3319};
test_output[6234] = '{32'h42491356};
test_index[6234] = '{5};
test_input[49880:49887] = '{32'h409721c9, 32'h41ed7f7d, 32'h42242c72, 32'h425b2692, 32'hc29b52d2, 32'hc2ae2775, 32'h4211e42a, 32'hc29ad708};
test_output[6235] = '{32'h425b2692};
test_index[6235] = '{3};
test_input[49888:49895] = '{32'h4227e2dd, 32'hc1694fba, 32'h4028e567, 32'h42a71e5d, 32'h421b8b1c, 32'hc1322e0f, 32'h422e91a4, 32'h4196aa37};
test_output[6236] = '{32'h42a71e5d};
test_index[6236] = '{3};
test_input[49896:49903] = '{32'hc189f6f6, 32'hc2174515, 32'h41e0b305, 32'hc20e9e8c, 32'h41fe5450, 32'h427f2d47, 32'h41b382d9, 32'h408db131};
test_output[6237] = '{32'h427f2d47};
test_index[6237] = '{5};
test_input[49904:49911] = '{32'hc2c1db46, 32'hc26a0d3b, 32'hc255df04, 32'hc2c4a598, 32'h428a32f8, 32'h42c0be6a, 32'hc2a7e19d, 32'hc295ede1};
test_output[6238] = '{32'h42c0be6a};
test_index[6238] = '{5};
test_input[49912:49919] = '{32'hc261fd8b, 32'hc14dc83b, 32'hc26d0e29, 32'hc26bbb5b, 32'hc2b3c5d4, 32'h42b70f14, 32'hc27b3567, 32'hc27e4691};
test_output[6239] = '{32'h42b70f14};
test_index[6239] = '{5};
test_input[49920:49927] = '{32'h428c5e91, 32'hc2890436, 32'hc2af47cf, 32'hc13a171d, 32'hc030911a, 32'hc1abf92c, 32'h4214735d, 32'h42201e62};
test_output[6240] = '{32'h428c5e91};
test_index[6240] = '{0};
test_input[49928:49935] = '{32'h42ad8a0e, 32'hc21a199c, 32'hc1531cfb, 32'hc2795704, 32'h429e2ef5, 32'hc2afb22a, 32'h421740d9, 32'hc2477877};
test_output[6241] = '{32'h42ad8a0e};
test_index[6241] = '{0};
test_input[49936:49943] = '{32'h42a9216a, 32'hc1845708, 32'hc2958f94, 32'h42a2a85e, 32'h424b5e4c, 32'hc1cb3073, 32'hc291427a, 32'hc2483387};
test_output[6242] = '{32'h42a9216a};
test_index[6242] = '{0};
test_input[49944:49951] = '{32'h42116da0, 32'hc295d32f, 32'hc0e6626c, 32'h42080d25, 32'hc2b2816d, 32'h42c079ef, 32'h3fb102a5, 32'h421ba7c3};
test_output[6243] = '{32'h42c079ef};
test_index[6243] = '{5};
test_input[49952:49959] = '{32'hc246bd45, 32'hbfdeedbe, 32'h4142e161, 32'hc254383a, 32'hc26d4f5c, 32'h414604fb, 32'h4259034a, 32'h42bc6f9f};
test_output[6244] = '{32'h42bc6f9f};
test_index[6244] = '{7};
test_input[49960:49967] = '{32'h42910aa9, 32'hc205115a, 32'h41f59efd, 32'h42ae7678, 32'h42ab4c22, 32'hc23cd64d, 32'hc2c77d98, 32'hc10e0dbd};
test_output[6245] = '{32'h42ae7678};
test_index[6245] = '{3};
test_input[49968:49975] = '{32'hbfa2a5d5, 32'hc1ed8579, 32'hc28b4945, 32'hc2c458d8, 32'h427a5499, 32'h41313398, 32'h41de0ec5, 32'hc236f19d};
test_output[6246] = '{32'h427a5499};
test_index[6246] = '{4};
test_input[49976:49983] = '{32'h4200f2cb, 32'hc2a1bed5, 32'h410e3401, 32'hc2511420, 32'hc2603c3e, 32'h4286ff79, 32'h42bf0e90, 32'h41b231cf};
test_output[6247] = '{32'h42bf0e90};
test_index[6247] = '{6};
test_input[49984:49991] = '{32'hc2375e19, 32'h41926a36, 32'hc0f019aa, 32'hc292c59f, 32'hc2944f3e, 32'hc2b589fd, 32'hc25c422c, 32'hc1be7c89};
test_output[6248] = '{32'h41926a36};
test_index[6248] = '{1};
test_input[49992:49999] = '{32'hc24c09cc, 32'hc0527aef, 32'h428ea4c4, 32'hc10f40ef, 32'hc222f4b4, 32'h40ad07fa, 32'h42bd7a57, 32'h4249b6f5};
test_output[6249] = '{32'h42bd7a57};
test_index[6249] = '{6};
test_input[50000:50007] = '{32'hc2a1476d, 32'h41d26e85, 32'hbe2b05e4, 32'h4286f015, 32'hc2316677, 32'hc1e55260, 32'hc2821050, 32'hc0aff615};
test_output[6250] = '{32'h4286f015};
test_index[6250] = '{3};
test_input[50008:50015] = '{32'h41b16cf9, 32'hc03792f4, 32'h419d8b19, 32'hc2a01e38, 32'hc234015a, 32'hc284d93d, 32'hc295c21f, 32'h4220d9dc};
test_output[6251] = '{32'h4220d9dc};
test_index[6251] = '{7};
test_input[50016:50023] = '{32'hc26d6e96, 32'h421ac97d, 32'h42beb81b, 32'h42032217, 32'h423537f3, 32'h42b0e3f5, 32'hc2938442, 32'hc1261d6f};
test_output[6252] = '{32'h42beb81b};
test_index[6252] = '{2};
test_input[50024:50031] = '{32'hc2451aab, 32'hc23c200c, 32'hc20994ff, 32'h41194d1d, 32'hc1539aff, 32'h428d61e5, 32'h4142aa5b, 32'h41d54bd3};
test_output[6253] = '{32'h428d61e5};
test_index[6253] = '{5};
test_input[50032:50039] = '{32'h40e23e88, 32'h42b4bf01, 32'hc28dbf53, 32'h40a0d09e, 32'hc23e9017, 32'h41338818, 32'h41e07292, 32'h4267e120};
test_output[6254] = '{32'h42b4bf01};
test_index[6254] = '{1};
test_input[50040:50047] = '{32'h4190866d, 32'h42c0baea, 32'hc1c516f1, 32'hc1a0b035, 32'h4231924d, 32'h4218561b, 32'h41da4413, 32'h42af4d47};
test_output[6255] = '{32'h42c0baea};
test_index[6255] = '{1};
test_input[50048:50055] = '{32'h41b0f282, 32'h4256549b, 32'h42bda89c, 32'h420b497f, 32'hc1ee488e, 32'hbf25afda, 32'hc0851d3d, 32'hc23cfa71};
test_output[6256] = '{32'h42bda89c};
test_index[6256] = '{2};
test_input[50056:50063] = '{32'hc1802df4, 32'h42a21767, 32'hc274b3b7, 32'h42ae1cbe, 32'h429be4d8, 32'hc17446e5, 32'hc1827aed, 32'h427c98e3};
test_output[6257] = '{32'h42ae1cbe};
test_index[6257] = '{3};
test_input[50064:50071] = '{32'hbf8fd0d5, 32'hc2792812, 32'hc21d9d71, 32'h42c6453a, 32'h422c0eba, 32'hc2278fa6, 32'h42b6681e, 32'h41f7d9f8};
test_output[6258] = '{32'h42c6453a};
test_index[6258] = '{3};
test_input[50072:50079] = '{32'hc0802ba5, 32'h41d4d0f3, 32'hc2b8f3d2, 32'h42b767be, 32'hc23c1752, 32'hc298e297, 32'h4278c6de, 32'h427dad48};
test_output[6259] = '{32'h42b767be};
test_index[6259] = '{3};
test_input[50080:50087] = '{32'hc2239ccd, 32'h40a6db71, 32'hc2a3ce14, 32'hc22b58b5, 32'hc28429d9, 32'hc25893c8, 32'hc23feb71, 32'h428071bd};
test_output[6260] = '{32'h428071bd};
test_index[6260] = '{7};
test_input[50088:50095] = '{32'hc25ab1c5, 32'h4240b296, 32'hc1db8f56, 32'hc20602ac, 32'hc1ca0c5f, 32'hc286871d, 32'h418692fd, 32'hc104dcd8};
test_output[6261] = '{32'h4240b296};
test_index[6261] = '{1};
test_input[50096:50103] = '{32'h42626cf3, 32'h41bef455, 32'h4245edf3, 32'h429dd2b1, 32'hc2b85209, 32'h429350d2, 32'h42c5974d, 32'h41aa6924};
test_output[6262] = '{32'h42c5974d};
test_index[6262] = '{6};
test_input[50104:50111] = '{32'hc15e8484, 32'hc1b3417b, 32'hc21758d1, 32'hc22824cb, 32'hc286f5ee, 32'hc25f1954, 32'h4237b6b7, 32'hc1563951};
test_output[6263] = '{32'h4237b6b7};
test_index[6263] = '{6};
test_input[50112:50119] = '{32'h4295fd3f, 32'hc20e9ec6, 32'hc22e7a55, 32'hc2bcf026, 32'hc2790c4e, 32'h42780225, 32'h4187099d, 32'h42535189};
test_output[6264] = '{32'h4295fd3f};
test_index[6264] = '{0};
test_input[50120:50127] = '{32'hc2b093dc, 32'hc19a2560, 32'h42874c56, 32'hc22a7f55, 32'h40098101, 32'h410dd08d, 32'h403eccd2, 32'hc1948e30};
test_output[6265] = '{32'h42874c56};
test_index[6265] = '{2};
test_input[50128:50135] = '{32'h427b3470, 32'h42816365, 32'hc1e5d6b8, 32'hc2b28824, 32'hc27a0493, 32'hc226dab9, 32'h427310fa, 32'h41523ae0};
test_output[6266] = '{32'h42816365};
test_index[6266] = '{1};
test_input[50136:50143] = '{32'hc1ed9b3b, 32'h42585c79, 32'h424508f2, 32'hc287af7a, 32'h42738d8d, 32'h4237d82a, 32'h42c477bb, 32'h3f0c73e5};
test_output[6267] = '{32'h42c477bb};
test_index[6267] = '{6};
test_input[50144:50151] = '{32'h42383f7d, 32'hc1b76862, 32'h3f941b79, 32'hbfc79c9a, 32'hc2765c9c, 32'h42aff03c, 32'hc2acb866, 32'h4213adb2};
test_output[6268] = '{32'h42aff03c};
test_index[6268] = '{5};
test_input[50152:50159] = '{32'h42b7f102, 32'hc2482f33, 32'h42922106, 32'hc24eb249, 32'h41cbb55d, 32'h4129d95b, 32'hc26301c7, 32'h42637c67};
test_output[6269] = '{32'h42b7f102};
test_index[6269] = '{0};
test_input[50160:50167] = '{32'hc22008f0, 32'h42b4a843, 32'hc27983ba, 32'hc2b9e5fa, 32'hc296498f, 32'h421164c6, 32'hc1dad6dc, 32'hc2a67ad6};
test_output[6270] = '{32'h42b4a843};
test_index[6270] = '{1};
test_input[50168:50175] = '{32'hc2b88049, 32'h41a25020, 32'hc1ba262a, 32'hc28517bd, 32'h411ac2dc, 32'hc28c0d75, 32'h40f0d282, 32'hc1979293};
test_output[6271] = '{32'h41a25020};
test_index[6271] = '{1};
test_input[50176:50183] = '{32'hc219bef3, 32'hc138836f, 32'hc28d7ff2, 32'hc167ac24, 32'hc263dc88, 32'hc2ba7987, 32'h42bb1139, 32'h42ac5a53};
test_output[6272] = '{32'h42bb1139};
test_index[6272] = '{6};
test_input[50184:50191] = '{32'hc164aacd, 32'h41e429e4, 32'hc2c2a72e, 32'hc2a3a4f2, 32'hc2223f7a, 32'h4236a0da, 32'hc26aac65, 32'h3f6f2cba};
test_output[6273] = '{32'h4236a0da};
test_index[6273] = '{5};
test_input[50192:50199] = '{32'h42b05171, 32'h420a04d2, 32'hc298959e, 32'hc27d3648, 32'hc20e7124, 32'h4292334f, 32'h418c4754, 32'h41a42aa2};
test_output[6274] = '{32'h42b05171};
test_index[6274] = '{0};
test_input[50200:50207] = '{32'hc14089bf, 32'hc124c12a, 32'h40a602aa, 32'h42649816, 32'hc2a0c3b6, 32'hc23f5ad5, 32'hc2a2b78b, 32'hc2126351};
test_output[6275] = '{32'h42649816};
test_index[6275] = '{3};
test_input[50208:50215] = '{32'hc2bbc6dc, 32'h42815c13, 32'h42acb477, 32'hc2a648b1, 32'hc2747fb6, 32'hc2ba8c65, 32'h423f19da, 32'hc298c354};
test_output[6276] = '{32'h42acb477};
test_index[6276] = '{2};
test_input[50216:50223] = '{32'h42543a04, 32'hc23a4091, 32'h4264434a, 32'hc22e7a12, 32'hc2a323c5, 32'h42761dca, 32'hc086a08d, 32'hc2b278fe};
test_output[6277] = '{32'h42761dca};
test_index[6277] = '{5};
test_input[50224:50231] = '{32'hc24d6071, 32'h41e57fd9, 32'h429a1948, 32'hc1c13404, 32'hc28369ba, 32'h4186219e, 32'hc115dac5, 32'hc2be2281};
test_output[6278] = '{32'h429a1948};
test_index[6278] = '{2};
test_input[50232:50239] = '{32'h3e338989, 32'h41a239eb, 32'hc25f5f41, 32'h42c158b3, 32'h42c3d8b3, 32'h408fc37d, 32'h417889ef, 32'h42bbdd5a};
test_output[6279] = '{32'h42c3d8b3};
test_index[6279] = '{4};
test_input[50240:50247] = '{32'h422bddaf, 32'hc2a9d69b, 32'hc29617a3, 32'hc2bba536, 32'hc27b380d, 32'h41d0265c, 32'hc1ea1e40, 32'h424d2de4};
test_output[6280] = '{32'h424d2de4};
test_index[6280] = '{7};
test_input[50248:50255] = '{32'h4290db94, 32'h41f55ab8, 32'h428f73c7, 32'hc264d434, 32'hc2a0b20e, 32'hc2b066bf, 32'hc2a2b887, 32'hc2399a81};
test_output[6281] = '{32'h4290db94};
test_index[6281] = '{0};
test_input[50256:50263] = '{32'hc00caf0d, 32'hc28e2d5a, 32'hc2b238f3, 32'hc2077e7a, 32'hc1751ff7, 32'h41c2abc8, 32'h429aed88, 32'hc1abd2c8};
test_output[6282] = '{32'h429aed88};
test_index[6282] = '{6};
test_input[50264:50271] = '{32'h41eff7c0, 32'h4194642f, 32'hc2b06ed2, 32'h424c2ec1, 32'h42a9c908, 32'hc29556b7, 32'hc2a444ae, 32'hc25a67fe};
test_output[6283] = '{32'h42a9c908};
test_index[6283] = '{4};
test_input[50272:50279] = '{32'h429d9911, 32'h428137db, 32'h42799461, 32'hc23565f0, 32'h420c3765, 32'hc243c92b, 32'hc1eabbe6, 32'h429f9e0d};
test_output[6284] = '{32'h429f9e0d};
test_index[6284] = '{7};
test_input[50280:50287] = '{32'h42c427d2, 32'h42c5ede9, 32'hc10678fb, 32'hc1222c93, 32'h4285420f, 32'h428e89d3, 32'h40959dcf, 32'h41574e52};
test_output[6285] = '{32'h42c5ede9};
test_index[6285] = '{1};
test_input[50288:50295] = '{32'h4274da5d, 32'h4280f6ab, 32'hc1e85df1, 32'h42c747d5, 32'hc2b968bd, 32'hc23c211c, 32'h428d3459, 32'hc1cf0201};
test_output[6286] = '{32'h42c747d5};
test_index[6286] = '{3};
test_input[50296:50303] = '{32'h428ff814, 32'h41978898, 32'h4248e8e8, 32'hc17436cb, 32'hc14e159d, 32'h42a648d6, 32'hc2bea0de, 32'hc2006433};
test_output[6287] = '{32'h42a648d6};
test_index[6287] = '{5};
test_input[50304:50311] = '{32'hc29de275, 32'hc290ab87, 32'h42c19968, 32'h42a1d918, 32'h42c5ba66, 32'h42be59e2, 32'h42bf8c9a, 32'hc1ae915f};
test_output[6288] = '{32'h42c5ba66};
test_index[6288] = '{4};
test_input[50312:50319] = '{32'h423f3acf, 32'h4283e6b1, 32'hc26886e5, 32'h428401b2, 32'h42a6486a, 32'h42bcf1a1, 32'hc1c7f02c, 32'h4195492f};
test_output[6289] = '{32'h42bcf1a1};
test_index[6289] = '{5};
test_input[50320:50327] = '{32'h425ed468, 32'hc29e873f, 32'hc299d94d, 32'h42aeea35, 32'hc227d898, 32'h425e8a3b, 32'hc193f179, 32'h42801d50};
test_output[6290] = '{32'h42aeea35};
test_index[6290] = '{3};
test_input[50328:50335] = '{32'h4231d52f, 32'h412177c9, 32'hc2a34be6, 32'hc2842b43, 32'hc2174920, 32'h42b8d4c1, 32'h4270eef8, 32'h41934829};
test_output[6291] = '{32'h42b8d4c1};
test_index[6291] = '{5};
test_input[50336:50343] = '{32'h42216a42, 32'h417691f3, 32'h4248fa9b, 32'hc248fbce, 32'hc2c00475, 32'h413e24b7, 32'hc2821482, 32'hc2bde42c};
test_output[6292] = '{32'h4248fa9b};
test_index[6292] = '{2};
test_input[50344:50351] = '{32'h41d936ac, 32'h421f2c44, 32'hc2756806, 32'h4290394f, 32'h42950558, 32'h428253dd, 32'hc1e1e063, 32'h427a8af6};
test_output[6293] = '{32'h42950558};
test_index[6293] = '{4};
test_input[50352:50359] = '{32'hc26407dc, 32'hc1d08189, 32'h42396e55, 32'hc257e60c, 32'h4183ea86, 32'h42003188, 32'h42a50427, 32'hc267b065};
test_output[6294] = '{32'h42a50427};
test_index[6294] = '{6};
test_input[50360:50367] = '{32'h4220ff3e, 32'h42171c15, 32'h42c42620, 32'hc1464bed, 32'hc29fb1e0, 32'h41cd23c0, 32'hc21ba46e, 32'h41c74704};
test_output[6295] = '{32'h42c42620};
test_index[6295] = '{2};
test_input[50368:50375] = '{32'hc1afda23, 32'h42b3eaf0, 32'h418e7936, 32'h42665129, 32'h428a0248, 32'h421bec00, 32'h424d7ba3, 32'hc2a550a0};
test_output[6296] = '{32'h42b3eaf0};
test_index[6296] = '{1};
test_input[50376:50383] = '{32'h41b64437, 32'hc29c37b8, 32'h4264d6af, 32'h41f50025, 32'hc24cef14, 32'h42c79eb1, 32'h42640218, 32'hc2a2333e};
test_output[6297] = '{32'h42c79eb1};
test_index[6297] = '{5};
test_input[50384:50391] = '{32'h42c1d33b, 32'h423d5261, 32'hc2676c6d, 32'hc1b62aa6, 32'hc2ba9149, 32'hc1ba99f7, 32'hc260a1ab, 32'hc13a3722};
test_output[6298] = '{32'h42c1d33b};
test_index[6298] = '{0};
test_input[50392:50399] = '{32'hc297cc8c, 32'h42507a9f, 32'hc29f3a3e, 32'h42b4473a, 32'hc2222f90, 32'h41ed8846, 32'h420978a9, 32'hc24f6525};
test_output[6299] = '{32'h42b4473a};
test_index[6299] = '{3};
test_input[50400:50407] = '{32'hc22f61f0, 32'h41d362a1, 32'hc1d42311, 32'hc2269814, 32'h41a26800, 32'h4206a127, 32'hc2849de7, 32'hc269f6c8};
test_output[6300] = '{32'h4206a127};
test_index[6300] = '{5};
test_input[50408:50415] = '{32'hc01e85e2, 32'hc290f3af, 32'hc2af9a23, 32'h425b8c13, 32'h421bec03, 32'h41e4c390, 32'h41a57909, 32'hc29d1b21};
test_output[6301] = '{32'h425b8c13};
test_index[6301] = '{3};
test_input[50416:50423] = '{32'h42a4f327, 32'h429dd55f, 32'hc10e2f2d, 32'hc2848a2e, 32'h424e861e, 32'hc2bed7fe, 32'hc019ba6b, 32'hc2627695};
test_output[6302] = '{32'h42a4f327};
test_index[6302] = '{0};
test_input[50424:50431] = '{32'h42b8012a, 32'hc087b8fa, 32'h418ae2a9, 32'h42929517, 32'hc11eb3d3, 32'hc1c7ba42, 32'hbf40b084, 32'h421c0880};
test_output[6303] = '{32'h42b8012a};
test_index[6303] = '{0};
test_input[50432:50439] = '{32'h4299a1e7, 32'h41a8917b, 32'h42b571b1, 32'hc28b6630, 32'h429b2b98, 32'hc299df0e, 32'hc2be2fef, 32'h42c77373};
test_output[6304] = '{32'h42c77373};
test_index[6304] = '{7};
test_input[50440:50447] = '{32'h4169f542, 32'hbf889670, 32'h42bb9572, 32'hc2ad6bb6, 32'h41b37f80, 32'hc1d0258b, 32'hc2c587e2, 32'hc1f62878};
test_output[6305] = '{32'h42bb9572};
test_index[6305] = '{2};
test_input[50448:50455] = '{32'h418637af, 32'hc205619e, 32'h421f60cc, 32'hc231b738, 32'hc29ae591, 32'hc154a875, 32'hc2b06ff6, 32'hc1d85463};
test_output[6306] = '{32'h421f60cc};
test_index[6306] = '{2};
test_input[50456:50463] = '{32'hc1fcd830, 32'h42149c6d, 32'h42beb07f, 32'hc27b19d1, 32'h427ada06, 32'hc0fb600f, 32'h425408d1, 32'hc257f02d};
test_output[6307] = '{32'h42beb07f};
test_index[6307] = '{2};
test_input[50464:50471] = '{32'hc2282984, 32'hc196f7b6, 32'h3f5cebf3, 32'h42679f1f, 32'hc2bf665d, 32'h42441423, 32'hc20ce6a2, 32'h40a2ff19};
test_output[6308] = '{32'h42679f1f};
test_index[6308] = '{3};
test_input[50472:50479] = '{32'hc2105f08, 32'h3f40185c, 32'h4258f1e0, 32'h41358e9e, 32'hc209a285, 32'h4252f16f, 32'h40271e23, 32'h42bd86a5};
test_output[6309] = '{32'h42bd86a5};
test_index[6309] = '{7};
test_input[50480:50487] = '{32'hc230b76d, 32'h41455292, 32'hc2c489df, 32'hc2044028, 32'hc28d5228, 32'hc211c791, 32'h415ed69d, 32'hc1e8d8d5};
test_output[6310] = '{32'h415ed69d};
test_index[6310] = '{6};
test_input[50488:50495] = '{32'h42968bfa, 32'hc259e0f7, 32'h41ea6d96, 32'hc29e6e07, 32'hc1a5f306, 32'h41ffdaa9, 32'hc2adb105, 32'h420358ed};
test_output[6311] = '{32'h42968bfa};
test_index[6311] = '{0};
test_input[50496:50503] = '{32'h42afe94a, 32'h4205f637, 32'h3ddf6682, 32'h42904376, 32'hc253a007, 32'h40e786aa, 32'hc28dafaf, 32'hc226f8f8};
test_output[6312] = '{32'h42afe94a};
test_index[6312] = '{0};
test_input[50504:50511] = '{32'h42530728, 32'h42a549ac, 32'hc2727390, 32'hc2515c7b, 32'h429d9575, 32'h42b7addf, 32'h42161141, 32'h4271d458};
test_output[6313] = '{32'h42b7addf};
test_index[6313] = '{5};
test_input[50512:50519] = '{32'h41864a77, 32'h4248b928, 32'hc0ecf0ae, 32'hc11392b4, 32'hc0df31e9, 32'hc2074614, 32'h425f4cb1, 32'h4160fcec};
test_output[6314] = '{32'h425f4cb1};
test_index[6314] = '{6};
test_input[50520:50527] = '{32'h424e05dd, 32'hc019e19d, 32'hbfd1d564, 32'h429f32fd, 32'hc223485d, 32'h419fd94e, 32'hc0e09f45, 32'h42361903};
test_output[6315] = '{32'h429f32fd};
test_index[6315] = '{3};
test_input[50528:50535] = '{32'h41df9dd6, 32'h414bd4a6, 32'h417ef59b, 32'h40d018bf, 32'hc2a644cf, 32'h425f4788, 32'hc2032bb9, 32'h42b89f32};
test_output[6316] = '{32'h42b89f32};
test_index[6316] = '{7};
test_input[50536:50543] = '{32'hc0c802d1, 32'hc088198c, 32'hc12d26f1, 32'h42c15009, 32'hc12f53ff, 32'hc2c46851, 32'h426d5f3e, 32'h4220e16f};
test_output[6317] = '{32'h42c15009};
test_index[6317] = '{3};
test_input[50544:50551] = '{32'hc25cc537, 32'h4145ba91, 32'h427b6add, 32'hc163653b, 32'hc075d719, 32'hc26d6650, 32'h423d7486, 32'hc2b2b7a1};
test_output[6318] = '{32'h427b6add};
test_index[6318] = '{2};
test_input[50552:50559] = '{32'hc23ec640, 32'h3f5edcb2, 32'hc218151f, 32'hc29599e4, 32'h41b4cf23, 32'hc2569128, 32'hc2a3e2c6, 32'hc25261d5};
test_output[6319] = '{32'h41b4cf23};
test_index[6319] = '{4};
test_input[50560:50567] = '{32'hc18eae85, 32'h42803f1e, 32'hc291165b, 32'h41bcb519, 32'hc220c169, 32'h42b350db, 32'h4262d6f1, 32'hc2b7a72a};
test_output[6320] = '{32'h42b350db};
test_index[6320] = '{5};
test_input[50568:50575] = '{32'hc27be2ed, 32'hc0dacfc8, 32'h422a0b63, 32'h42ab0019, 32'h415d4ba8, 32'hc19dfea1, 32'hc237da50, 32'h41b5e654};
test_output[6321] = '{32'h42ab0019};
test_index[6321] = '{3};
test_input[50576:50583] = '{32'h42b63192, 32'hc18f51f4, 32'h408b61a6, 32'hc2b8e94e, 32'h42bfa8d7, 32'hc2078633, 32'h428a95b2, 32'hbf776bc9};
test_output[6322] = '{32'h42bfa8d7};
test_index[6322] = '{4};
test_input[50584:50591] = '{32'hc241efb4, 32'hc283d3df, 32'hbedae51a, 32'h4283a00c, 32'hc2a56ec7, 32'hc2a8c6bd, 32'h3e90769c, 32'hc211a56e};
test_output[6323] = '{32'h4283a00c};
test_index[6323] = '{3};
test_input[50592:50599] = '{32'h4184c099, 32'hc22c1a84, 32'h42c071e5, 32'hc17cef9c, 32'hc26e8c84, 32'h428d6db9, 32'h4251cb54, 32'hc29c6f3b};
test_output[6324] = '{32'h42c071e5};
test_index[6324] = '{2};
test_input[50600:50607] = '{32'hc24c5acf, 32'h428c9a83, 32'hc21c6524, 32'hc2822bfa, 32'hc2386097, 32'hc2c38d81, 32'hc2c5185f, 32'h42ac498f};
test_output[6325] = '{32'h42ac498f};
test_index[6325] = '{7};
test_input[50608:50615] = '{32'h42c07905, 32'hc29b646a, 32'h42135acc, 32'h426e3c01, 32'hc1cb6bb3, 32'h4299f8a6, 32'h40cb060d, 32'hc231806c};
test_output[6326] = '{32'h42c07905};
test_index[6326] = '{0};
test_input[50616:50623] = '{32'h401327f8, 32'h4285d269, 32'hc263f8e0, 32'h4127250f, 32'h3dafd719, 32'h4258a39d, 32'h425ffa8a, 32'h420cfea2};
test_output[6327] = '{32'h4285d269};
test_index[6327] = '{1};
test_input[50624:50631] = '{32'hc091b6b6, 32'hc12754fb, 32'hc2c140c8, 32'hc23649b4, 32'h4226ad7f, 32'h42c446b2, 32'h421c2060, 32'h42222ce3};
test_output[6328] = '{32'h42c446b2};
test_index[6328] = '{5};
test_input[50632:50639] = '{32'hc2a4854a, 32'h42513136, 32'h42260c1b, 32'h42a7e7b9, 32'hc1cfe86f, 32'h42b49e0a, 32'hc252e697, 32'h42845c30};
test_output[6329] = '{32'h42b49e0a};
test_index[6329] = '{5};
test_input[50640:50647] = '{32'hc246459c, 32'hc2507918, 32'hc16cffae, 32'hc1f92ce7, 32'h42a3ea22, 32'h429b0ef2, 32'hc2b4b13b, 32'h422e8871};
test_output[6330] = '{32'h42a3ea22};
test_index[6330] = '{4};
test_input[50648:50655] = '{32'hbf15ee48, 32'hc05a9b28, 32'h41ac675f, 32'h4282656a, 32'h418d6806, 32'hc26eda48, 32'h42c77ef2, 32'h40a70569};
test_output[6331] = '{32'h42c77ef2};
test_index[6331] = '{6};
test_input[50656:50663] = '{32'h4187957c, 32'h407a4926, 32'hc23e79e9, 32'hc2a89ad1, 32'hc2619d6d, 32'hc1d62ddd, 32'h41d4051d, 32'hc2aefcb5};
test_output[6332] = '{32'h41d4051d};
test_index[6332] = '{6};
test_input[50664:50671] = '{32'h418fde79, 32'h42810b44, 32'h41b5af55, 32'hc2051107, 32'h42b4ae37, 32'h4297ce18, 32'h42c102b0, 32'h42384669};
test_output[6333] = '{32'h42c102b0};
test_index[6333] = '{6};
test_input[50672:50679] = '{32'hc2c4a69f, 32'h42446568, 32'hc2108d35, 32'h41dcf1fb, 32'h429ddae5, 32'h42b7e866, 32'h428d5808, 32'hc23cd130};
test_output[6334] = '{32'h42b7e866};
test_index[6334] = '{5};
test_input[50680:50687] = '{32'h4274a0d1, 32'hc033c379, 32'h41ea96ad, 32'h429b9a4f, 32'h41e5cbd3, 32'h41c1812d, 32'hc1c37d5f, 32'h4239b9de};
test_output[6335] = '{32'h429b9a4f};
test_index[6335] = '{3};
test_input[50688:50695] = '{32'hc28aa064, 32'h42b65374, 32'hc26e3fb5, 32'hc18bcb31, 32'hc28b4eb4, 32'h4278c71e, 32'hc2814aec, 32'hc26944bb};
test_output[6336] = '{32'h42b65374};
test_index[6336] = '{1};
test_input[50696:50703] = '{32'hc18f7f60, 32'h42824676, 32'h42a8c64f, 32'h4260c58e, 32'h423ddf8f, 32'h421effb9, 32'hbfdacc2c, 32'hc2c45848};
test_output[6337] = '{32'h42a8c64f};
test_index[6337] = '{2};
test_input[50704:50711] = '{32'h41c922fe, 32'hc2bea675, 32'h429cf336, 32'hc19004d5, 32'hc2420e51, 32'h40c19c1f, 32'h42a300b7, 32'h42a7d965};
test_output[6338] = '{32'h42a7d965};
test_index[6338] = '{7};
test_input[50712:50719] = '{32'h42c666f7, 32'hc24a3446, 32'hc2126ad6, 32'h42918e93, 32'hc1be85b1, 32'h41cd812a, 32'hc257f91e, 32'h41e70ddf};
test_output[6339] = '{32'h42c666f7};
test_index[6339] = '{0};
test_input[50720:50727] = '{32'h42a08902, 32'h428020df, 32'h41c27752, 32'h427261dc, 32'h422eadd6, 32'h42670c56, 32'h429c1d16, 32'h40578f9b};
test_output[6340] = '{32'h42a08902};
test_index[6340] = '{0};
test_input[50728:50735] = '{32'h42a5fd97, 32'hc1ae5a8a, 32'hc2ac647f, 32'hc1bc7225, 32'hc1e53834, 32'h4291202d, 32'hc2a94704, 32'hc2c35644};
test_output[6341] = '{32'h42a5fd97};
test_index[6341] = '{0};
test_input[50736:50743] = '{32'hc227f823, 32'hc21ea6d6, 32'hc294a237, 32'h421929c7, 32'hc25b76df, 32'hc295fc9a, 32'h3fed51df, 32'hc2c6d7d7};
test_output[6342] = '{32'h421929c7};
test_index[6342] = '{3};
test_input[50744:50751] = '{32'hc04b1fc8, 32'h42a2c23d, 32'h41451b08, 32'h42c08cea, 32'h42619304, 32'hc2b68691, 32'h3fa0d62e, 32'h41fb3b60};
test_output[6343] = '{32'h42c08cea};
test_index[6343] = '{3};
test_input[50752:50759] = '{32'hc2492fec, 32'hc28cf733, 32'h422f7675, 32'hc2b1b488, 32'h41ccf780, 32'h429cebc9, 32'hc27fe800, 32'hc2c552e8};
test_output[6344] = '{32'h429cebc9};
test_index[6344] = '{5};
test_input[50760:50767] = '{32'h42519e14, 32'hc259f4e7, 32'h421da712, 32'hc192c9f3, 32'hc2216213, 32'hc2149e13, 32'hc1c9be9e, 32'hc2a81ccf};
test_output[6345] = '{32'h42519e14};
test_index[6345] = '{0};
test_input[50768:50775] = '{32'hc22edda2, 32'hc1b84ae5, 32'h41d3374c, 32'h41a429aa, 32'h4277614b, 32'hc1ab5d98, 32'hc1f02d6c, 32'hc2a21264};
test_output[6346] = '{32'h4277614b};
test_index[6346] = '{4};
test_input[50776:50783] = '{32'hc285933f, 32'h428d42a2, 32'h4111d692, 32'hc2785fd3, 32'hc222c608, 32'h4180b8b8, 32'hc24beb7a, 32'h42940ee7};
test_output[6347] = '{32'h42940ee7};
test_index[6347] = '{7};
test_input[50784:50791] = '{32'h424e830f, 32'hc2300d46, 32'h425ab91f, 32'h419a283f, 32'hc1db8b79, 32'h42307c11, 32'h4268c2d8, 32'h424d47c7};
test_output[6348] = '{32'h4268c2d8};
test_index[6348] = '{6};
test_input[50792:50799] = '{32'hc2460099, 32'hc219e417, 32'h42456bcb, 32'h42bedd54, 32'h418f1fbd, 32'hc2a77b79, 32'hc25ee539, 32'h42855bb7};
test_output[6349] = '{32'h42bedd54};
test_index[6349] = '{3};
test_input[50800:50807] = '{32'hc25cb873, 32'h411ae26d, 32'hc2a447a7, 32'hc28c0607, 32'hc258e861, 32'h42641535, 32'h42889592, 32'h419bfef4};
test_output[6350] = '{32'h42889592};
test_index[6350] = '{6};
test_input[50808:50815] = '{32'h42a26afc, 32'hc2b231d8, 32'hc1ef761a, 32'hc11b6458, 32'h4207d5b2, 32'hc173303f, 32'h42560fb9, 32'h424e08e4};
test_output[6351] = '{32'h42a26afc};
test_index[6351] = '{0};
test_input[50816:50823] = '{32'hc186a42b, 32'h42553ac2, 32'hc2382496, 32'hc28fcfa6, 32'hc237acce, 32'h4240c090, 32'hc29629a7, 32'hc2156306};
test_output[6352] = '{32'h42553ac2};
test_index[6352] = '{1};
test_input[50824:50831] = '{32'h428bd24b, 32'h41abd12a, 32'h42110d6b, 32'h408afb7a, 32'hc203dbf8, 32'h42626e2a, 32'h4271507c, 32'h42368877};
test_output[6353] = '{32'h428bd24b};
test_index[6353] = '{0};
test_input[50832:50839] = '{32'h4287de24, 32'hc035f8a2, 32'hc1b7bcb7, 32'hc2b0a1ad, 32'h42c1f2e6, 32'hc25959e8, 32'h428f5868, 32'hc250a793};
test_output[6354] = '{32'h42c1f2e6};
test_index[6354] = '{4};
test_input[50840:50847] = '{32'hc116ec86, 32'hc1fcd34f, 32'hc1f45601, 32'hc0e8a2d2, 32'h41fc3f69, 32'hc0b74a16, 32'h42ba94ff, 32'hc1fb2c64};
test_output[6355] = '{32'h42ba94ff};
test_index[6355] = '{6};
test_input[50848:50855] = '{32'hc20cdd22, 32'h418172a2, 32'hc2250d56, 32'hc260b6e2, 32'h3d955464, 32'hc29bbb18, 32'h42b03e0c, 32'h4278fec5};
test_output[6356] = '{32'h42b03e0c};
test_index[6356] = '{6};
test_input[50856:50863] = '{32'hc293c8df, 32'h41fdad83, 32'hc121a9ef, 32'h4242764e, 32'hc2826f26, 32'h42adc0a0, 32'hc228af39, 32'hc274976f};
test_output[6357] = '{32'h42adc0a0};
test_index[6357] = '{5};
test_input[50864:50871] = '{32'hc2029277, 32'h4187b0b6, 32'h426f1abd, 32'h42807d43, 32'hc1a238fa, 32'h422fdeb8, 32'hc21b6522, 32'h41e26a87};
test_output[6358] = '{32'h42807d43};
test_index[6358] = '{3};
test_input[50872:50879] = '{32'hc1c65690, 32'h421fe7c9, 32'hc0b689f1, 32'hc25c4226, 32'h421f5300, 32'h42c02079, 32'h42c35f62, 32'h42953bd8};
test_output[6359] = '{32'h42c35f62};
test_index[6359] = '{6};
test_input[50880:50887] = '{32'h42a12497, 32'h416bdc0f, 32'h4139d52a, 32'h425879d6, 32'hc280b73e, 32'h3fcef75e, 32'hc2bc3b7c, 32'h4209245d};
test_output[6360] = '{32'h42a12497};
test_index[6360] = '{0};
test_input[50888:50895] = '{32'hc2b03c10, 32'hc25b3d52, 32'h41d33e44, 32'h41fe3eac, 32'h4157ff1a, 32'h420c79c0, 32'hc282fe66, 32'h41a9908b};
test_output[6361] = '{32'h420c79c0};
test_index[6361] = '{5};
test_input[50896:50903] = '{32'h42614227, 32'hc2c41ce2, 32'hc2ad60a0, 32'h3e8786a7, 32'hc1cffae2, 32'hbff84ffe, 32'h42bb6068, 32'h4292ee5d};
test_output[6362] = '{32'h42bb6068};
test_index[6362] = '{6};
test_input[50904:50911] = '{32'h412400a4, 32'h4145184b, 32'h426a2e29, 32'hc1f2c4f9, 32'h41ffaad5, 32'h41d701ab, 32'hc140b925, 32'h42230eda};
test_output[6363] = '{32'h426a2e29};
test_index[6363] = '{2};
test_input[50912:50919] = '{32'hc005c813, 32'h3fe9671f, 32'hc2b93dd7, 32'hc2acd01e, 32'h41768087, 32'hc19f5f62, 32'h40db77b2, 32'h42ab8179};
test_output[6364] = '{32'h42ab8179};
test_index[6364] = '{7};
test_input[50920:50927] = '{32'h40efa86d, 32'h41af4c0b, 32'h4297c731, 32'h42989b90, 32'h420d2b5d, 32'hc24d0f62, 32'h4260b2f6, 32'hc267a657};
test_output[6365] = '{32'h42989b90};
test_index[6365] = '{3};
test_input[50928:50935] = '{32'hc2769988, 32'h4294c5a0, 32'h42198d3b, 32'h41f6897d, 32'h424955f1, 32'h418bf219, 32'hc0ae568d, 32'h4187a978};
test_output[6366] = '{32'h4294c5a0};
test_index[6366] = '{1};
test_input[50936:50943] = '{32'h42878299, 32'h427a60d2, 32'hc1cf7940, 32'hc29b96fe, 32'hc1031367, 32'hc19710c7, 32'h42b56d21, 32'h424f3249};
test_output[6367] = '{32'h42b56d21};
test_index[6367] = '{6};
test_input[50944:50951] = '{32'hc2c5c95c, 32'hc1eef27d, 32'hc286cfa4, 32'h429a7b70, 32'h4126c962, 32'h41b4c9ba, 32'hc23a5d04, 32'hc2a42426};
test_output[6368] = '{32'h429a7b70};
test_index[6368] = '{3};
test_input[50952:50959] = '{32'hc1a28813, 32'hc2678cd6, 32'hc2c3f653, 32'h41b99574, 32'h427ed093, 32'h42c68905, 32'hc295a754, 32'hc235b636};
test_output[6369] = '{32'h42c68905};
test_index[6369] = '{5};
test_input[50960:50967] = '{32'h427ea7a0, 32'h42b709c1, 32'h42373200, 32'hc2854127, 32'hc23606e9, 32'h4110dd42, 32'h424d3273, 32'hc17a7d8c};
test_output[6370] = '{32'h42b709c1};
test_index[6370] = '{1};
test_input[50968:50975] = '{32'hc1cfc0ea, 32'hc1a3403d, 32'h41376d6b, 32'hc27ff16b, 32'h419f83f6, 32'hc1e4e5db, 32'h426e3102, 32'hc13df07b};
test_output[6371] = '{32'h426e3102};
test_index[6371] = '{6};
test_input[50976:50983] = '{32'hc1c10dbc, 32'hc298bc8a, 32'hbe171cbc, 32'h4293f5d5, 32'h41cf8aad, 32'h42b86f7c, 32'hc1d0d65e, 32'hc270a4db};
test_output[6372] = '{32'h42b86f7c};
test_index[6372] = '{5};
test_input[50984:50991] = '{32'hc0f81f07, 32'hc271e13a, 32'h4294085d, 32'h4218af75, 32'h41925dfb, 32'h4113570e, 32'h3fbade3b, 32'hc2700670};
test_output[6373] = '{32'h4294085d};
test_index[6373] = '{2};
test_input[50992:50999] = '{32'hc180f95a, 32'h426047c4, 32'h41e6b4a7, 32'hc29356e2, 32'h42c5abfa, 32'hc2bb26c0, 32'h425fa5c2, 32'hc202f716};
test_output[6374] = '{32'h42c5abfa};
test_index[6374] = '{4};
test_input[51000:51007] = '{32'hc25854ef, 32'h42327729, 32'hc29cdb7f, 32'h421d34b1, 32'h4232622f, 32'h425b74d4, 32'hc1629fb4, 32'h4280bae5};
test_output[6375] = '{32'h4280bae5};
test_index[6375] = '{7};
test_input[51008:51015] = '{32'hc243f08d, 32'hc1c3a6c4, 32'h41b476a3, 32'h426c54d8, 32'hc1b2f352, 32'hc26cf2f4, 32'hc26e967c, 32'hc231fd19};
test_output[6376] = '{32'h426c54d8};
test_index[6376] = '{3};
test_input[51016:51023] = '{32'h42882ba7, 32'h429f99e1, 32'h41ce8c1e, 32'hc2384864, 32'h42b4463f, 32'h3dd2f1b1, 32'h42a30cf5, 32'h41f24d8f};
test_output[6377] = '{32'h42b4463f};
test_index[6377] = '{4};
test_input[51024:51031] = '{32'hc26e5de2, 32'hc27e2f07, 32'h417adf2a, 32'hc268546d, 32'hc22d8c8b, 32'hc2b6e852, 32'h423b2bf9, 32'hc2924c5a};
test_output[6378] = '{32'h423b2bf9};
test_index[6378] = '{6};
test_input[51032:51039] = '{32'h42539519, 32'hc24cbc79, 32'hc1e83f17, 32'h41350e08, 32'hc2612325, 32'hc0e2174a, 32'hc23106db, 32'h4219779b};
test_output[6379] = '{32'h42539519};
test_index[6379] = '{0};
test_input[51040:51047] = '{32'h41f7b42f, 32'h42161413, 32'hc25dce71, 32'h4208a032, 32'h413ecf05, 32'hc2b32969, 32'h428ba0f7, 32'h41379db8};
test_output[6380] = '{32'h428ba0f7};
test_index[6380] = '{6};
test_input[51048:51055] = '{32'h41240800, 32'h42bd5286, 32'h41ceba47, 32'hc2764078, 32'hc27aad6f, 32'hc29214bf, 32'hc24315e3, 32'hc28ab2f3};
test_output[6381] = '{32'h42bd5286};
test_index[6381] = '{1};
test_input[51056:51063] = '{32'h42c5d0d2, 32'h40a1e52b, 32'hc2adcc86, 32'h41d33ff5, 32'h4090763d, 32'hc20b9dda, 32'h4253a618, 32'h41ae705c};
test_output[6382] = '{32'h42c5d0d2};
test_index[6382] = '{0};
test_input[51064:51071] = '{32'hc27636dd, 32'hc16b2b36, 32'h3f487a3c, 32'hc1ba61d2, 32'hc134c8bf, 32'hc0adfd2f, 32'h42116efc, 32'h42a6e928};
test_output[6383] = '{32'h42a6e928};
test_index[6383] = '{7};
test_input[51072:51079] = '{32'hc292b934, 32'h42a11b03, 32'hc1fd0378, 32'hc1c27c73, 32'hc28831b2, 32'hc26fdd3b, 32'h42908104, 32'h421eeff1};
test_output[6384] = '{32'h42a11b03};
test_index[6384] = '{1};
test_input[51080:51087] = '{32'hc2111201, 32'hc0b4d45a, 32'h424828aa, 32'hc1fa9553, 32'hc29a970c, 32'h41a82356, 32'hc2bed59d, 32'hc16bc1a5};
test_output[6385] = '{32'h424828aa};
test_index[6385] = '{2};
test_input[51088:51095] = '{32'h42b24032, 32'hc085efac, 32'hc2b4d806, 32'h42896ff6, 32'hc2bd0489, 32'hc2ad51bb, 32'hc2ac7efc, 32'hc142f120};
test_output[6386] = '{32'h42b24032};
test_index[6386] = '{0};
test_input[51096:51103] = '{32'h42b1ae3c, 32'hc2680974, 32'hc225d643, 32'h4123cc9f, 32'hc2c3a2af, 32'h41dac6da, 32'hc13d0643, 32'h420733be};
test_output[6387] = '{32'h42b1ae3c};
test_index[6387] = '{0};
test_input[51104:51111] = '{32'hc2a1c7b7, 32'h4156f167, 32'hc177d674, 32'hc266184c, 32'hc116838a, 32'hc16ac592, 32'hc2911aec, 32'hc28070ca};
test_output[6388] = '{32'h4156f167};
test_index[6388] = '{1};
test_input[51112:51119] = '{32'hc09c61f7, 32'hc2bd4af7, 32'h426bbd8a, 32'h428043cd, 32'h42066388, 32'hc2006c20, 32'hc1d6f6a3, 32'h429e8885};
test_output[6389] = '{32'h429e8885};
test_index[6389] = '{7};
test_input[51120:51127] = '{32'h415daefb, 32'hc2a20ef8, 32'hc2c19975, 32'h42b4ce05, 32'h429510b7, 32'hc2a32bc7, 32'h4234896c, 32'h41b04087};
test_output[6390] = '{32'h42b4ce05};
test_index[6390] = '{3};
test_input[51128:51135] = '{32'hc22ba998, 32'h42b826a2, 32'hc2561482, 32'hc21aab02, 32'hc2665157, 32'h41bae186, 32'h4125b88a, 32'h41ed4242};
test_output[6391] = '{32'h42b826a2};
test_index[6391] = '{1};
test_input[51136:51143] = '{32'hc18b2866, 32'hc0e36772, 32'h421a8075, 32'hc0a564a5, 32'hc2820300, 32'hc2c3cdee, 32'h42671525, 32'h42ade6e5};
test_output[6392] = '{32'h42ade6e5};
test_index[6392] = '{7};
test_input[51144:51151] = '{32'hc25ef8ec, 32'hc0946888, 32'hc28025ff, 32'h42afa188, 32'h42c61fdb, 32'hc01ba8db, 32'hc287e107, 32'h3f1cafb3};
test_output[6393] = '{32'h42c61fdb};
test_index[6393] = '{4};
test_input[51152:51159] = '{32'hc27c9391, 32'hc12729ae, 32'h4236f65f, 32'h42479e7e, 32'h4268aab9, 32'h4284e24a, 32'hc2be6cc3, 32'hc24dbc41};
test_output[6394] = '{32'h4284e24a};
test_index[6394] = '{5};
test_input[51160:51167] = '{32'h41d786fb, 32'h41f260ca, 32'hc2a44172, 32'h421cc261, 32'h42263b8f, 32'hc0c410e7, 32'hc2c0191d, 32'h42a9f867};
test_output[6395] = '{32'h42a9f867};
test_index[6395] = '{7};
test_input[51168:51175] = '{32'hc25dd406, 32'h4280ded5, 32'hc1020a40, 32'h41309189, 32'h41c3e004, 32'hc15c0cf2, 32'h41efb839, 32'h42714b83};
test_output[6396] = '{32'h4280ded5};
test_index[6396] = '{1};
test_input[51176:51183] = '{32'h40fe028d, 32'h426fd9f4, 32'hc2c3ff45, 32'h428015d1, 32'h42264a3b, 32'h42b8e087, 32'h4281cbd5, 32'h41f931f2};
test_output[6397] = '{32'h42b8e087};
test_index[6397] = '{5};
test_input[51184:51191] = '{32'hc10464a3, 32'h42056e6c, 32'hc2855741, 32'hc24a9189, 32'h42ba1df6, 32'hc0e04fcf, 32'h428d60ca, 32'hc2624e10};
test_output[6398] = '{32'h42ba1df6};
test_index[6398] = '{4};
test_input[51192:51199] = '{32'h4280b1b5, 32'h41fba407, 32'h42bbba0e, 32'h41547d04, 32'hc1f8e522, 32'h4252857b, 32'hc2bbd565, 32'h424ae6cf};
test_output[6399] = '{32'h42bbba0e};
test_index[6399] = '{2};
test_input[51200:51207] = '{32'h41b5c068, 32'h42a7c3fb, 32'h3f37f920, 32'h40ccce87, 32'h42a6f041, 32'h42816fe3, 32'h4136d382, 32'hbf3c1eaf};
test_output[6400] = '{32'h42a7c3fb};
test_index[6400] = '{1};
test_input[51208:51215] = '{32'hc112117b, 32'h429287cc, 32'h4203ad93, 32'hc26a11b5, 32'hc12d88e3, 32'hc2301e8a, 32'h42c0107e, 32'h40809d97};
test_output[6401] = '{32'h42c0107e};
test_index[6401] = '{6};
test_input[51216:51223] = '{32'hc24758de, 32'hc1fe9376, 32'hc290a64f, 32'h42b11804, 32'h3f6193cc, 32'h41f553f1, 32'h41680a99, 32'hc1fa7a31};
test_output[6402] = '{32'h42b11804};
test_index[6402] = '{3};
test_input[51224:51231] = '{32'h418f48a9, 32'hc2b668b8, 32'h42b8f6e7, 32'h420cb78d, 32'h42b16cc5, 32'hc2af456d, 32'h4235d36c, 32'hc2af24e8};
test_output[6403] = '{32'h42b8f6e7};
test_index[6403] = '{2};
test_input[51232:51239] = '{32'h42a27abf, 32'hc199303e, 32'h40a959ff, 32'h428ccd5e, 32'hc22cd961, 32'hc27208e7, 32'hc11e8cd2, 32'hc2b1b969};
test_output[6404] = '{32'h42a27abf};
test_index[6404] = '{0};
test_input[51240:51247] = '{32'h3ff19ed0, 32'h4290972f, 32'hc292043d, 32'h422870f5, 32'hc2b5e1d5, 32'h42640ab2, 32'h42c42645, 32'hc2748800};
test_output[6405] = '{32'h42c42645};
test_index[6405] = '{6};
test_input[51248:51255] = '{32'hc204dccb, 32'h424eb02a, 32'hc0e0bd2f, 32'hc27a85be, 32'hc2280257, 32'hc241974f, 32'hc03acf0f, 32'hc234d1dd};
test_output[6406] = '{32'h424eb02a};
test_index[6406] = '{1};
test_input[51256:51263] = '{32'hc2321ebb, 32'h4284e555, 32'hc29c17a1, 32'h4216b939, 32'hc1f9ed29, 32'h424ee5fc, 32'hc2c2a4e4, 32'hc114c787};
test_output[6407] = '{32'h4284e555};
test_index[6407] = '{1};
test_input[51264:51271] = '{32'hc281f26f, 32'hc18108e8, 32'hc091ac88, 32'hc287187b, 32'hc15ef452, 32'h4203d13d, 32'h428777c9, 32'h427282f5};
test_output[6408] = '{32'h428777c9};
test_index[6408] = '{6};
test_input[51272:51279] = '{32'h42b91e2d, 32'hc00a5cfc, 32'hc2a5bd85, 32'hc2a6fa31, 32'h4292463f, 32'h42b106c8, 32'h41cd392b, 32'hc2b59fcf};
test_output[6409] = '{32'h42b91e2d};
test_index[6409] = '{0};
test_input[51280:51287] = '{32'h424b4f6e, 32'hc233c580, 32'hbfeae21e, 32'h42c00e37, 32'h425a5a72, 32'h40cef2f3, 32'h401872ca, 32'hc2001da7};
test_output[6410] = '{32'h42c00e37};
test_index[6410] = '{3};
test_input[51288:51295] = '{32'hc122d238, 32'h424fce5c, 32'h4290c2b4, 32'hc22d9a47, 32'hc1d80069, 32'hc1f2a2ed, 32'h4271e3b1, 32'h4237158e};
test_output[6411] = '{32'h4290c2b4};
test_index[6411] = '{2};
test_input[51296:51303] = '{32'hc21255fd, 32'hc29c2e47, 32'hc1b7c268, 32'h4164ccd2, 32'h4213e69d, 32'h42742353, 32'h42870aa6, 32'h4280ed6d};
test_output[6412] = '{32'h42870aa6};
test_index[6412] = '{6};
test_input[51304:51311] = '{32'h428d8810, 32'hc2b84ecd, 32'hc15949f1, 32'hc26fbc63, 32'hc254bb64, 32'h42c45aac, 32'h4015a89d, 32'h4243a32c};
test_output[6413] = '{32'h42c45aac};
test_index[6413] = '{5};
test_input[51312:51319] = '{32'h42395dcf, 32'h42a227f8, 32'hc226e9c2, 32'hc25486eb, 32'h42475b18, 32'h429c1471, 32'hc2a39389, 32'hc108625c};
test_output[6414] = '{32'h42a227f8};
test_index[6414] = '{1};
test_input[51320:51327] = '{32'hc2b147ee, 32'hc2192188, 32'h3fa327f0, 32'hc234cf40, 32'hc2a265c9, 32'h42986603, 32'h428f4406, 32'h410a41f5};
test_output[6415] = '{32'h42986603};
test_index[6415] = '{5};
test_input[51328:51335] = '{32'h41a26329, 32'hc1d13f74, 32'h417419c8, 32'h425a2228, 32'hc1d79925, 32'hc28c310e, 32'h4283aac4, 32'hc21ded00};
test_output[6416] = '{32'h4283aac4};
test_index[6416] = '{6};
test_input[51336:51343] = '{32'hc1cee3c9, 32'h42aa1aea, 32'hc1894c23, 32'hc229de4a, 32'hc2a22b31, 32'hc2701448, 32'hc263f09e, 32'hc1ded4c6};
test_output[6417] = '{32'h42aa1aea};
test_index[6417] = '{1};
test_input[51344:51351] = '{32'h41665251, 32'hc1756888, 32'hc1847543, 32'hc1e4596f, 32'hc212f1f5, 32'hc28f5788, 32'hc257f1af, 32'hc1b15019};
test_output[6418] = '{32'h41665251};
test_index[6418] = '{0};
test_input[51352:51359] = '{32'hc190e84a, 32'hc21a28fa, 32'h41de8de3, 32'hc1367360, 32'h421855f5, 32'h41b5f75e, 32'h4222c71b, 32'h42a3aa78};
test_output[6419] = '{32'h42a3aa78};
test_index[6419] = '{7};
test_input[51360:51367] = '{32'hc21b6075, 32'h424017cf, 32'hc1bf5710, 32'hc1134368, 32'h418fada9, 32'h41c423f6, 32'hc2297547, 32'hc108d4c6};
test_output[6420] = '{32'h424017cf};
test_index[6420] = '{1};
test_input[51368:51375] = '{32'hc251a269, 32'hc0f284ff, 32'hc2b92ae0, 32'hc2021545, 32'h42996011, 32'h42b3b699, 32'h429ee91c, 32'h428c9ab7};
test_output[6421] = '{32'h42b3b699};
test_index[6421] = '{5};
test_input[51376:51383] = '{32'h41c3036e, 32'h41649ddc, 32'h411dbf60, 32'hc19481ec, 32'h42a383ed, 32'h41b35d9c, 32'h4210b02f, 32'h4290a347};
test_output[6422] = '{32'h42a383ed};
test_index[6422] = '{4};
test_input[51384:51391] = '{32'h422b738c, 32'hc2a9347c, 32'h4225cf74, 32'hc244f4de, 32'h4246d293, 32'hc2b31e5a, 32'hc29db421, 32'h425d11b0};
test_output[6423] = '{32'h425d11b0};
test_index[6423] = '{7};
test_input[51392:51399] = '{32'hc27d3b0f, 32'hc26c063d, 32'h4297146c, 32'hc2794c03, 32'h418c3935, 32'h424ab288, 32'hc29c9a41, 32'hbf926d8c};
test_output[6424] = '{32'h4297146c};
test_index[6424] = '{2};
test_input[51400:51407] = '{32'h41e5ae68, 32'hc14cadaa, 32'hc1e266b8, 32'h4287dd2e, 32'h4237442d, 32'hc1986b50, 32'hc25d6ef4, 32'hc1c79865};
test_output[6425] = '{32'h4287dd2e};
test_index[6425] = '{3};
test_input[51408:51415] = '{32'hc211c36f, 32'h428b475f, 32'hc258c833, 32'h412fddb0, 32'hc27d833a, 32'h4224665f, 32'hc0ab581e, 32'hc28c7262};
test_output[6426] = '{32'h428b475f};
test_index[6426] = '{1};
test_input[51416:51423] = '{32'h429dda00, 32'hc1bf6859, 32'h40c3082e, 32'h417f9881, 32'hc25b191a, 32'h42ac9382, 32'hc12e098b, 32'hbffc8d29};
test_output[6427] = '{32'h42ac9382};
test_index[6427] = '{5};
test_input[51424:51431] = '{32'hc21af6d9, 32'hc1e4fc46, 32'h428d4d9a, 32'h40e80d5b, 32'hc1417925, 32'h41dd45b4, 32'hc025006d, 32'hc288828d};
test_output[6428] = '{32'h428d4d9a};
test_index[6428] = '{2};
test_input[51432:51439] = '{32'hc28aec90, 32'hc28cdb5e, 32'h424d9e32, 32'h41d6fadb, 32'h42a3652c, 32'h428f9819, 32'h4202e2c0, 32'hc2b95b1f};
test_output[6429] = '{32'h42a3652c};
test_index[6429] = '{4};
test_input[51440:51447] = '{32'hc2c50460, 32'hc191d9ef, 32'h4276189d, 32'h42c5db5e, 32'h42141486, 32'h428aabe8, 32'h41e7320e, 32'h4152247d};
test_output[6430] = '{32'h42c5db5e};
test_index[6430] = '{3};
test_input[51448:51455] = '{32'hc202d9a9, 32'hc2ba5991, 32'h426b7263, 32'h429766ec, 32'h418acb21, 32'hc2b0cde6, 32'hc239158a, 32'h42188166};
test_output[6431] = '{32'h429766ec};
test_index[6431] = '{3};
test_input[51456:51463] = '{32'h42318434, 32'h42c315b8, 32'hc1d5e0e3, 32'h4269137b, 32'hc218c924, 32'h42b12e37, 32'h4291f3b6, 32'h41f7577a};
test_output[6432] = '{32'h42c315b8};
test_index[6432] = '{1};
test_input[51464:51471] = '{32'h41cf5d4f, 32'hc16049a8, 32'h4255577d, 32'hc1358908, 32'h4276676c, 32'h41650c14, 32'h416458f3, 32'h42ab3a2d};
test_output[6433] = '{32'h42ab3a2d};
test_index[6433] = '{7};
test_input[51472:51479] = '{32'hc2114bff, 32'h41c07030, 32'h429597c5, 32'h412f97ab, 32'hc108bfdc, 32'hc2ac51ef, 32'h419f20c8, 32'h4288764a};
test_output[6434] = '{32'h429597c5};
test_index[6434] = '{2};
test_input[51480:51487] = '{32'hc26b2b58, 32'h42b1c34a, 32'h42c74e5a, 32'hc2311598, 32'hbfe79483, 32'hc188373f, 32'hc0ea1d30, 32'h40854fd2};
test_output[6435] = '{32'h42c74e5a};
test_index[6435] = '{2};
test_input[51488:51495] = '{32'h421c82ff, 32'hc20fb102, 32'h41c5dfa1, 32'h423dd83f, 32'h41a07ae0, 32'h4281cf21, 32'hc23c83b2, 32'h42a070d4};
test_output[6436] = '{32'h42a070d4};
test_index[6436] = '{7};
test_input[51496:51503] = '{32'h416f981b, 32'hc1e2ae9b, 32'hc2c5dcdb, 32'hc2b06190, 32'hc27ef257, 32'hc17ffc7b, 32'h416c3c34, 32'h42938b01};
test_output[6437] = '{32'h42938b01};
test_index[6437] = '{7};
test_input[51504:51511] = '{32'h3ea3534a, 32'h4132c2e5, 32'h4293ef4f, 32'hc2975c07, 32'hc2aaf9f3, 32'hbfd22dcf, 32'hc2c1ad03, 32'h412ad847};
test_output[6438] = '{32'h4293ef4f};
test_index[6438] = '{2};
test_input[51512:51519] = '{32'h42157084, 32'h429753bb, 32'hc0c3e7d3, 32'hc20c4dc2, 32'hc293058d, 32'h42b8ffff, 32'hc2983a0e, 32'hc2a1c34a};
test_output[6439] = '{32'h42b8ffff};
test_index[6439] = '{5};
test_input[51520:51527] = '{32'h42aab54a, 32'h4265bf8d, 32'h41746241, 32'hc13fdfb2, 32'hc074a036, 32'hc26f0af6, 32'hc296e0c7, 32'h41e9ba52};
test_output[6440] = '{32'h42aab54a};
test_index[6440] = '{0};
test_input[51528:51535] = '{32'hc2764d09, 32'h41b8135c, 32'hc243fae0, 32'hc22b4e4a, 32'hc1e84d02, 32'hc2055e35, 32'hc2944f5f, 32'hc1b84f45};
test_output[6441] = '{32'h41b8135c};
test_index[6441] = '{1};
test_input[51536:51543] = '{32'h4240b9e3, 32'hc28874f8, 32'h42536aec, 32'hc2bb1d86, 32'h425bccab, 32'hc1d3c685, 32'hc2adb735, 32'h4022275f};
test_output[6442] = '{32'h425bccab};
test_index[6442] = '{4};
test_input[51544:51551] = '{32'hc2926f8a, 32'h421431d8, 32'h42b3c0ba, 32'hc1613b88, 32'hc2b666e7, 32'h42c43e28, 32'hc297216c, 32'hc211db6a};
test_output[6443] = '{32'h42c43e28};
test_index[6443] = '{5};
test_input[51552:51559] = '{32'h42baf5bc, 32'hc1d5edb1, 32'h42b6b3a7, 32'hc1b1e794, 32'hc2c1c1c0, 32'hc1fbb8af, 32'hc1999d54, 32'h42b5ccc1};
test_output[6444] = '{32'h42baf5bc};
test_index[6444] = '{0};
test_input[51560:51567] = '{32'hc23e129e, 32'hc2c2deed, 32'h42667792, 32'hc01e11bb, 32'hc240ad4e, 32'hc2a5350e, 32'h427111f0, 32'hc28930e1};
test_output[6445] = '{32'h427111f0};
test_index[6445] = '{6};
test_input[51568:51575] = '{32'h42c053e4, 32'h42a56f0a, 32'hc2a9ee8a, 32'h42383150, 32'hc2c69a79, 32'h42282c12, 32'hc18e7942, 32'hc029bbd4};
test_output[6446] = '{32'h42c053e4};
test_index[6446] = '{0};
test_input[51576:51583] = '{32'h41f82792, 32'h406c55b3, 32'hc24fe623, 32'hc246a81e, 32'hc2901f1e, 32'hc2955cf0, 32'h42745c5a, 32'h42abb56d};
test_output[6447] = '{32'h42abb56d};
test_index[6447] = '{7};
test_input[51584:51591] = '{32'hc07701ea, 32'hc2c1b8ab, 32'h41af3b5e, 32'h42a205a5, 32'h417d7715, 32'h42a849d8, 32'hbeab2034, 32'hc290ee72};
test_output[6448] = '{32'h42a849d8};
test_index[6448] = '{5};
test_input[51592:51599] = '{32'hc2a94277, 32'h421c2ad4, 32'hc2adab06, 32'hc2b53ff5, 32'hc29b195a, 32'hc1d7c573, 32'hc2c7038b, 32'h4204d6a5};
test_output[6449] = '{32'h421c2ad4};
test_index[6449] = '{1};
test_input[51600:51607] = '{32'hc29b49ab, 32'hc1b1d286, 32'h414e5255, 32'h4242949a, 32'hc27f483d, 32'h424e0308, 32'h42b3cf6b, 32'h4255ac47};
test_output[6450] = '{32'h42b3cf6b};
test_index[6450] = '{6};
test_input[51608:51615] = '{32'h429e655c, 32'hc24a9360, 32'h41d454ae, 32'h424fa2cb, 32'hc284cac4, 32'h412cee88, 32'hc2c5003c, 32'hc1fe3af6};
test_output[6451] = '{32'h429e655c};
test_index[6451] = '{0};
test_input[51616:51623] = '{32'h40f31781, 32'hc225da27, 32'hc18ff41b, 32'hc240503e, 32'hc2b5fd78, 32'h41f9292c, 32'hc21af7b5, 32'hc2b2e17b};
test_output[6452] = '{32'h41f9292c};
test_index[6452] = '{5};
test_input[51624:51631] = '{32'hc1d9513b, 32'h42b36b06, 32'h41b119bd, 32'h42241cf0, 32'h42c134ef, 32'hc06860eb, 32'h41e3f5a8, 32'h4114afbe};
test_output[6453] = '{32'h42c134ef};
test_index[6453] = '{4};
test_input[51632:51639] = '{32'h420c0acd, 32'hc297c053, 32'hc24c3238, 32'h42b54765, 32'hc1fe5e2a, 32'hc21f70d3, 32'h42001a4e, 32'hc2c03733};
test_output[6454] = '{32'h42b54765};
test_index[6454] = '{3};
test_input[51640:51647] = '{32'hc2939bc7, 32'h411c276d, 32'hc2a674cd, 32'h42a05157, 32'hc2183baf, 32'h40585931, 32'hc1e13797, 32'h42a6f8d0};
test_output[6455] = '{32'h42a6f8d0};
test_index[6455] = '{7};
test_input[51648:51655] = '{32'h42074ed4, 32'hc182e64a, 32'h42858d0d, 32'hc28f984c, 32'h42556e04, 32'hc162ec1b, 32'hc2186929, 32'hc29b591b};
test_output[6456] = '{32'h42858d0d};
test_index[6456] = '{2};
test_input[51656:51663] = '{32'hbfc2478a, 32'hc16acbc4, 32'h42a837ad, 32'h4270199b, 32'h42b73546, 32'hc2bd61c9, 32'hc237ff37, 32'hc265b2aa};
test_output[6457] = '{32'h42b73546};
test_index[6457] = '{4};
test_input[51664:51671] = '{32'h4297c260, 32'hc2b3864b, 32'h4236f83e, 32'hc208a8db, 32'h424b61e0, 32'h414f508f, 32'hc28a4e05, 32'hc1cd1b22};
test_output[6458] = '{32'h4297c260};
test_index[6458] = '{0};
test_input[51672:51679] = '{32'hc0a73f28, 32'hc1c5788f, 32'hc18bcfcc, 32'hc0e17caf, 32'hc20b94fc, 32'h410170ba, 32'hc2a992a3, 32'h42480484};
test_output[6459] = '{32'h42480484};
test_index[6459] = '{7};
test_input[51680:51687] = '{32'h41a7efb2, 32'h41973b58, 32'hc2a0511f, 32'hc104d223, 32'hc0a053d0, 32'hc23f6c92, 32'hc2a5f994, 32'h428b7838};
test_output[6460] = '{32'h428b7838};
test_index[6460] = '{7};
test_input[51688:51695] = '{32'hc181aac6, 32'h4264a303, 32'h4294fa9f, 32'h4290948a, 32'hc10f8176, 32'hc2b29f22, 32'h41bb1d5b, 32'h42b5ca03};
test_output[6461] = '{32'h42b5ca03};
test_index[6461] = '{7};
test_input[51696:51703] = '{32'hc26e42b7, 32'hc20c8511, 32'hc22dcce6, 32'hc214737b, 32'hc2828037, 32'h406f559e, 32'hc2af0c5d, 32'h42b7a4aa};
test_output[6462] = '{32'h42b7a4aa};
test_index[6462] = '{7};
test_input[51704:51711] = '{32'hc0d6e475, 32'h41f33197, 32'h424d4d74, 32'hc2227a84, 32'h4249ae04, 32'hc29bd6c0, 32'hc28224e4, 32'h40da210a};
test_output[6463] = '{32'h424d4d74};
test_index[6463] = '{2};
test_input[51712:51719] = '{32'hc2bad73e, 32'hc241fb54, 32'h42c42dc5, 32'h42adebc1, 32'h423b4e91, 32'hc28245ff, 32'h420cea0c, 32'h41634545};
test_output[6464] = '{32'h42c42dc5};
test_index[6464] = '{2};
test_input[51720:51727] = '{32'h42a18fdc, 32'hc28bf133, 32'hc1f3f7c5, 32'hc26ee7fc, 32'h4272fa08, 32'hc1ab0633, 32'h42b33d76, 32'hc2a0e70c};
test_output[6465] = '{32'h42b33d76};
test_index[6465] = '{6};
test_input[51728:51735] = '{32'hc202864e, 32'h41378bbc, 32'hc2850216, 32'hc21c1dc0, 32'h413c4cb7, 32'hc27d2a36, 32'h41ec1ed9, 32'hc147caca};
test_output[6466] = '{32'h41ec1ed9};
test_index[6466] = '{6};
test_input[51736:51743] = '{32'hc1f6b44f, 32'hc09cd40a, 32'h418c61d0, 32'h429a3a19, 32'hc2349600, 32'hbfdd1b68, 32'h4201aa87, 32'hc21d0ceb};
test_output[6467] = '{32'h429a3a19};
test_index[6467] = '{3};
test_input[51744:51751] = '{32'hc2aec6eb, 32'h428225d0, 32'h42be51b5, 32'hc2ae9d65, 32'hc2bdb9d5, 32'h428e3c2d, 32'h427073ca, 32'hc0c5611a};
test_output[6468] = '{32'h42be51b5};
test_index[6468] = '{2};
test_input[51752:51759] = '{32'h42ad494d, 32'hc11497cf, 32'h41b20629, 32'hc2a14fb4, 32'hc15e6e28, 32'hc1d885f0, 32'h41cd78af, 32'hc1a29b0a};
test_output[6469] = '{32'h42ad494d};
test_index[6469] = '{0};
test_input[51760:51767] = '{32'h41845e39, 32'hc28ba448, 32'hc2a48542, 32'h41bd92c9, 32'hc20bf9ce, 32'hc298bf85, 32'h429de9c0, 32'hc21862d6};
test_output[6470] = '{32'h429de9c0};
test_index[6470] = '{6};
test_input[51768:51775] = '{32'h410d4fc3, 32'hc247ebf0, 32'h42c4db8e, 32'hc08fb72f, 32'hc259942a, 32'h41963a18, 32'hc2b485ee, 32'hc2b34ebd};
test_output[6471] = '{32'h42c4db8e};
test_index[6471] = '{2};
test_input[51776:51783] = '{32'hc28c8143, 32'hc291153b, 32'h42678bbc, 32'hc2bd0529, 32'hc0d60d89, 32'hc22b3024, 32'hc2310f3e, 32'hc2831438};
test_output[6472] = '{32'h42678bbc};
test_index[6472] = '{2};
test_input[51784:51791] = '{32'hc2689ea3, 32'h42b545f2, 32'h42a91a2e, 32'h42067987, 32'h42776af3, 32'h42aeeac6, 32'hc28e95c5, 32'h42b043a9};
test_output[6473] = '{32'h42b545f2};
test_index[6473] = '{1};
test_input[51792:51799] = '{32'h424882cc, 32'hc1d3c517, 32'hc1998d67, 32'hc299f5a6, 32'h412d2ac2, 32'h429a7e30, 32'h427adf54, 32'hc202bee6};
test_output[6474] = '{32'h429a7e30};
test_index[6474] = '{5};
test_input[51800:51807] = '{32'hc258b18b, 32'hc0c31358, 32'hc27b934a, 32'hc0d9ead2, 32'h427ed821, 32'h4136b27e, 32'hc2bb7095, 32'h4297f052};
test_output[6475] = '{32'h4297f052};
test_index[6475] = '{7};
test_input[51808:51815] = '{32'hc24c4141, 32'hc249103b, 32'h41f0d188, 32'hc2bd9f9f, 32'h4255fffb, 32'hc29d8a4c, 32'hc25eca57, 32'hc18041d3};
test_output[6476] = '{32'h4255fffb};
test_index[6476] = '{4};
test_input[51816:51823] = '{32'h42207ff5, 32'hc103da5a, 32'h428ea8ef, 32'hc24c4f04, 32'h415d3828, 32'h42564958, 32'hc25d1208, 32'h4254af21};
test_output[6477] = '{32'h428ea8ef};
test_index[6477] = '{2};
test_input[51824:51831] = '{32'hc1a13b31, 32'h4030345d, 32'hc09c1dd9, 32'hc21e6ed9, 32'h421dfdfb, 32'hc2a1251b, 32'h421c0425, 32'hc2b429e5};
test_output[6478] = '{32'h421dfdfb};
test_index[6478] = '{4};
test_input[51832:51839] = '{32'hc24ad6ad, 32'h420393c3, 32'h4290f440, 32'hc22c6b4a, 32'h40fdfa53, 32'hc1defc52, 32'h421cde32, 32'h42207781};
test_output[6479] = '{32'h4290f440};
test_index[6479] = '{2};
test_input[51840:51847] = '{32'h42084467, 32'hc2899733, 32'h42b03c35, 32'h42223e12, 32'hc1756900, 32'h3ff13f0e, 32'h423ba903, 32'h41da696f};
test_output[6480] = '{32'h42b03c35};
test_index[6480] = '{2};
test_input[51848:51855] = '{32'hc2a1e98a, 32'hc2b96ced, 32'hc2815b11, 32'hc2c384de, 32'h41939f90, 32'hc2ab4ff1, 32'h40bc1457, 32'h420fa67f};
test_output[6481] = '{32'h420fa67f};
test_index[6481] = '{7};
test_input[51856:51863] = '{32'h41dc1ba7, 32'h40d86077, 32'hc242f7e7, 32'hc2c78755, 32'hc2b92e47, 32'h42be5841, 32'h42b9d260, 32'hc00b9a7a};
test_output[6482] = '{32'h42be5841};
test_index[6482] = '{5};
test_input[51864:51871] = '{32'hc2a373e2, 32'hc205adee, 32'hc292d2af, 32'hc255d2be, 32'hc2a5296b, 32'hc2b4bf15, 32'h410f4cab, 32'hc2baab25};
test_output[6483] = '{32'h410f4cab};
test_index[6483] = '{6};
test_input[51872:51879] = '{32'h429c9e4a, 32'h4283c536, 32'hbe80b9e6, 32'hc2abb96c, 32'hc1b483cc, 32'h42478178, 32'h42b5372e, 32'hc27acbe6};
test_output[6484] = '{32'h42b5372e};
test_index[6484] = '{6};
test_input[51880:51887] = '{32'h422bf9bf, 32'hc2acd87d, 32'hc2122d11, 32'h4186ce01, 32'h428b2cf8, 32'hc2738460, 32'hc23c6042, 32'h416ebee8};
test_output[6485] = '{32'h428b2cf8};
test_index[6485] = '{4};
test_input[51888:51895] = '{32'h42b7c146, 32'h42a9767a, 32'hc1097258, 32'h428f64bd, 32'h4202ed7d, 32'hc25394ad, 32'h4280fe08, 32'hc1aef4cf};
test_output[6486] = '{32'h42b7c146};
test_index[6486] = '{0};
test_input[51896:51903] = '{32'h42c02d3b, 32'h42431a25, 32'h42ac7a9c, 32'hc2b6fe72, 32'hbf605bc7, 32'h427a2e2c, 32'h428a5998, 32'hc195b700};
test_output[6487] = '{32'h42c02d3b};
test_index[6487] = '{0};
test_input[51904:51911] = '{32'hc24da83d, 32'hc1433d1b, 32'h40328ce2, 32'hc2bc3cc9, 32'h416f606d, 32'h415f4f85, 32'h4280748e, 32'h411e63b1};
test_output[6488] = '{32'h4280748e};
test_index[6488] = '{6};
test_input[51912:51919] = '{32'hc1621b71, 32'h42adc7bc, 32'h422c7c3f, 32'h422f8435, 32'hc2bd861e, 32'hc2aaa2dc, 32'h42a72f01, 32'hc1b42c4b};
test_output[6489] = '{32'h42adc7bc};
test_index[6489] = '{1};
test_input[51920:51927] = '{32'hc1dd859b, 32'hc26bbdfc, 32'h42048e3e, 32'hc29c95a4, 32'hc28a6b4e, 32'h41a454bc, 32'h420a044e, 32'h42c1b87d};
test_output[6490] = '{32'h42c1b87d};
test_index[6490] = '{7};
test_input[51928:51935] = '{32'h40e69b31, 32'hc2921bf2, 32'hc2a41b2b, 32'hc2092fa2, 32'h41404a07, 32'h4247bd8f, 32'hc221e0d6, 32'h42061909};
test_output[6491] = '{32'h4247bd8f};
test_index[6491] = '{5};
test_input[51936:51943] = '{32'hc23d0d3d, 32'hc29e35b0, 32'h414ad57f, 32'hc28449ef, 32'h42251007, 32'h427eeea7, 32'h42b2f3d2, 32'h42c343c5};
test_output[6492] = '{32'h42c343c5};
test_index[6492] = '{7};
test_input[51944:51951] = '{32'hc1c787f0, 32'h40fc9888, 32'h41ce99a9, 32'h423e8074, 32'h41b88c11, 32'h4213ea79, 32'hc0d11dfd, 32'h404639a2};
test_output[6493] = '{32'h423e8074};
test_index[6493] = '{3};
test_input[51952:51959] = '{32'h414e5dca, 32'h4231bfcd, 32'hc2801398, 32'h420beee1, 32'h423f4748, 32'h42847f4c, 32'h426df35b, 32'hc260b127};
test_output[6494] = '{32'h42847f4c};
test_index[6494] = '{5};
test_input[51960:51967] = '{32'hc294b403, 32'h41261c79, 32'h419f52eb, 32'h42b116cc, 32'hc1879f51, 32'h42aa48b4, 32'h41c697fd, 32'hc280da4c};
test_output[6495] = '{32'h42b116cc};
test_index[6495] = '{3};
test_input[51968:51975] = '{32'hc24ad525, 32'h4243657c, 32'hc25f3878, 32'hc287338b, 32'h42ba0e7a, 32'h408e23d5, 32'hc20a7f3f, 32'hc2113b1e};
test_output[6496] = '{32'h42ba0e7a};
test_index[6496] = '{4};
test_input[51976:51983] = '{32'hc2b78956, 32'hc10ba8cf, 32'hc258b07f, 32'hc19aa65c, 32'h40cece62, 32'h428d06ac, 32'hc24a1005, 32'h428b9bc4};
test_output[6497] = '{32'h428d06ac};
test_index[6497] = '{5};
test_input[51984:51991] = '{32'h40c96473, 32'hc1d8ee10, 32'h41401e1b, 32'h41e84cdb, 32'hc1f3177f, 32'h42135c04, 32'h42ac4d87, 32'h41b35985};
test_output[6498] = '{32'h42ac4d87};
test_index[6498] = '{6};
test_input[51992:51999] = '{32'h41e997e8, 32'hc1dcf4e9, 32'hc1ec38a1, 32'h3fa49615, 32'hc2c1d5f1, 32'h428aae18, 32'hc2c5b707, 32'h427ba3f0};
test_output[6499] = '{32'h428aae18};
test_index[6499] = '{5};
test_input[52000:52007] = '{32'hc06737e9, 32'hc23b6e54, 32'h418f6241, 32'hc271bbef, 32'h425ad17b, 32'h3fe0753a, 32'h42c46b4b, 32'h429f360c};
test_output[6500] = '{32'h42c46b4b};
test_index[6500] = '{6};
test_input[52008:52015] = '{32'hc299623e, 32'hc285ac95, 32'hc28fe313, 32'h426898bd, 32'h4091146d, 32'h42834973, 32'hc2a390b4, 32'h42659554};
test_output[6501] = '{32'h42834973};
test_index[6501] = '{5};
test_input[52016:52023] = '{32'h42b344be, 32'hc224e4ae, 32'h41f1e261, 32'h4299625a, 32'hc2c14403, 32'hc28b7347, 32'h429c3a09, 32'h4092d665};
test_output[6502] = '{32'h42b344be};
test_index[6502] = '{0};
test_input[52024:52031] = '{32'hc2abb8fa, 32'hc225a027, 32'h4209708a, 32'h425bab82, 32'hc2ace8a9, 32'hc0c851e5, 32'h3f862e23, 32'hc2882912};
test_output[6503] = '{32'h425bab82};
test_index[6503] = '{3};
test_input[52032:52039] = '{32'h4234c1e1, 32'h414ed8be, 32'hc1709d40, 32'hc2989455, 32'hc157c24e, 32'h411b7694, 32'h422b4e4c, 32'hc1e42889};
test_output[6504] = '{32'h4234c1e1};
test_index[6504] = '{0};
test_input[52040:52047] = '{32'h428e2ed6, 32'h4186b560, 32'h428bc1e0, 32'h41630067, 32'h42985857, 32'h40caea29, 32'hc1b2ed89, 32'hc209f31f};
test_output[6505] = '{32'h42985857};
test_index[6505] = '{4};
test_input[52048:52055] = '{32'h429a78c9, 32'hc28f9905, 32'hc1b15407, 32'h42abfda3, 32'h415788c5, 32'h427e75e2, 32'hc245770e, 32'hc13c0d90};
test_output[6506] = '{32'h42abfda3};
test_index[6506] = '{3};
test_input[52056:52063] = '{32'h420ad1ee, 32'h4105b57d, 32'h420a4c57, 32'hc26512d8, 32'hc29e4a6d, 32'h41ce8201, 32'hc11bc635, 32'hc28c1d26};
test_output[6507] = '{32'h420ad1ee};
test_index[6507] = '{0};
test_input[52064:52071] = '{32'hc28c1e7f, 32'hc2c7daa3, 32'hc1927021, 32'h424bc1b4, 32'h41eb03ed, 32'h4224c5af, 32'hc243f43c, 32'h416c522c};
test_output[6508] = '{32'h424bc1b4};
test_index[6508] = '{3};
test_input[52072:52079] = '{32'h4210d298, 32'h429725a5, 32'h423c3ecd, 32'h41f92d4f, 32'hc2b486a2, 32'h4248d738, 32'hc1d65397, 32'h42ae614d};
test_output[6509] = '{32'h42ae614d};
test_index[6509] = '{7};
test_input[52080:52087] = '{32'hc289d778, 32'h42a858a8, 32'h42abd9b2, 32'h429fef52, 32'hc29c268d, 32'h42443ed0, 32'h41a41527, 32'hc2b81f68};
test_output[6510] = '{32'h42abd9b2};
test_index[6510] = '{2};
test_input[52088:52095] = '{32'hc2265219, 32'hc2917b3a, 32'hc27c9162, 32'h3fd994c1, 32'hc2abee5c, 32'hc262e93f, 32'hc2a735a2, 32'h4284e4cc};
test_output[6511] = '{32'h4284e4cc};
test_index[6511] = '{7};
test_input[52096:52103] = '{32'h4296984a, 32'hc2c08351, 32'hc1907a32, 32'h42541dbb, 32'hc200469d, 32'h42053b0f, 32'h3d8c035d, 32'h41b9bf99};
test_output[6512] = '{32'h4296984a};
test_index[6512] = '{0};
test_input[52104:52111] = '{32'h42086345, 32'h429d7333, 32'hc2661002, 32'h427e9ea2, 32'hc195bfb0, 32'hc185a686, 32'h41b25076, 32'h429ef8ea};
test_output[6513] = '{32'h429ef8ea};
test_index[6513] = '{7};
test_input[52112:52119] = '{32'h41e26de9, 32'h421043b0, 32'h421ad4cc, 32'h4267689f, 32'h41f1a4b0, 32'h41466061, 32'hc2bf5ed5, 32'h41ab626b};
test_output[6514] = '{32'h4267689f};
test_index[6514] = '{3};
test_input[52120:52127] = '{32'h42abe2a2, 32'hc29f78a3, 32'hc228eca6, 32'hc28cac1d, 32'h40ff338f, 32'h40ebdb3e, 32'h42271a87, 32'hc20cb628};
test_output[6515] = '{32'h42abe2a2};
test_index[6515] = '{0};
test_input[52128:52135] = '{32'h4196b57e, 32'h428c40ff, 32'h40a43252, 32'hc2acff5c, 32'h425dc1d2, 32'hc2c42008, 32'hc1983877, 32'hc25f08c7};
test_output[6516] = '{32'h428c40ff};
test_index[6516] = '{1};
test_input[52136:52143] = '{32'hc26bc015, 32'hc2b9f680, 32'h42bdd8db, 32'h42ad26b9, 32'hc1a9eb3e, 32'hc1ac0851, 32'hc1a3a093, 32'hc244dd67};
test_output[6517] = '{32'h42bdd8db};
test_index[6517] = '{2};
test_input[52144:52151] = '{32'hc1b9036c, 32'h426a368b, 32'hc29094d6, 32'hc25d8396, 32'hc29c132e, 32'h42884db7, 32'hc164df7e, 32'h42bfccd5};
test_output[6518] = '{32'h42bfccd5};
test_index[6518] = '{7};
test_input[52152:52159] = '{32'h425a5165, 32'h416efa6f, 32'h42b63d4c, 32'h416113f8, 32'hc27320eb, 32'h420a9028, 32'h42a5eede, 32'hc1b42284};
test_output[6519] = '{32'h42b63d4c};
test_index[6519] = '{2};
test_input[52160:52167] = '{32'hc0ff471a, 32'hc0966d42, 32'h428581e6, 32'hc28eb3fa, 32'hc28963af, 32'h42387c25, 32'hc1bccaa2, 32'h417ab043};
test_output[6520] = '{32'h428581e6};
test_index[6520] = '{2};
test_input[52168:52175] = '{32'hc2179827, 32'h41ca0e3a, 32'h429377c8, 32'h42b98840, 32'hc2ad1128, 32'h42b4495c, 32'hc0d766a0, 32'h428acb83};
test_output[6521] = '{32'h42b98840};
test_index[6521] = '{3};
test_input[52176:52183] = '{32'hc295576a, 32'h421849ef, 32'h422e516b, 32'h419772d8, 32'h423a0cc7, 32'h422a5dda, 32'hc1cdd024, 32'hc2bd9032};
test_output[6522] = '{32'h423a0cc7};
test_index[6522] = '{4};
test_input[52184:52191] = '{32'hc2b90ba9, 32'h42789b50, 32'h4220047a, 32'hc17adffd, 32'h41f2baaa, 32'hc2a0c73d, 32'h423f5b79, 32'hc18458a1};
test_output[6523] = '{32'h42789b50};
test_index[6523] = '{1};
test_input[52192:52199] = '{32'h42c1716f, 32'h42826916, 32'hc28d3072, 32'h429bb2e2, 32'h4136113f, 32'hc27c9426, 32'h42029f68, 32'hc28d25be};
test_output[6524] = '{32'h42c1716f};
test_index[6524] = '{0};
test_input[52200:52207] = '{32'hc142bb80, 32'hc27068ba, 32'hc1a40d88, 32'h41208723, 32'h413e2af8, 32'h420d3430, 32'hc2aa9976, 32'hc1c7361c};
test_output[6525] = '{32'h420d3430};
test_index[6525] = '{5};
test_input[52208:52215] = '{32'hc217de72, 32'hc2a8b23e, 32'h42861826, 32'h421a3222, 32'h424dfc7b, 32'hc288d181, 32'h41a416ad, 32'hc2c1e6ed};
test_output[6526] = '{32'h42861826};
test_index[6526] = '{2};
test_input[52216:52223] = '{32'h429f353b, 32'h422c9890, 32'h42bc626a, 32'h42c70948, 32'h427fc932, 32'h42664b59, 32'hc1ff9b26, 32'h429e80d2};
test_output[6527] = '{32'h42c70948};
test_index[6527] = '{3};
test_input[52224:52231] = '{32'hc129f634, 32'h41a348b1, 32'hc2b63714, 32'h42b39331, 32'h42c25242, 32'h423399a9, 32'hc22b8cb8, 32'h429ef93b};
test_output[6528] = '{32'h42c25242};
test_index[6528] = '{4};
test_input[52232:52239] = '{32'hc219feba, 32'hc2b4cc82, 32'hc21a72a6, 32'hc0066c06, 32'h418f2bc0, 32'hc2a39a54, 32'hc293ad14, 32'hc1f1cabc};
test_output[6529] = '{32'h418f2bc0};
test_index[6529] = '{4};
test_input[52240:52247] = '{32'h4164a673, 32'hc1c92372, 32'hc1bb6f2c, 32'h42381732, 32'h41a0873a, 32'h42405431, 32'h428f546b, 32'hc250bcc9};
test_output[6530] = '{32'h428f546b};
test_index[6530] = '{6};
test_input[52248:52255] = '{32'h4226a700, 32'hc29061a1, 32'h42063da5, 32'hc205e937, 32'h423adea1, 32'hc2954a70, 32'h41ccbb63, 32'hc18d8417};
test_output[6531] = '{32'h423adea1};
test_index[6531] = '{4};
test_input[52256:52263] = '{32'hc268da43, 32'h41f66c66, 32'hc20e9ad0, 32'h42c052bd, 32'h41bd761d, 32'hc2aaa475, 32'h41d66699, 32'hc0a0fcbd};
test_output[6532] = '{32'h42c052bd};
test_index[6532] = '{3};
test_input[52264:52271] = '{32'h42c26b63, 32'h42bdb691, 32'hc25031d3, 32'hc2c18d5a, 32'hc29e1284, 32'h42b582f8, 32'h42b7f4a9, 32'h4232a0e1};
test_output[6533] = '{32'h42c26b63};
test_index[6533] = '{0};
test_input[52272:52279] = '{32'hc2a98b32, 32'hbfeb6222, 32'h42a00036, 32'h421aea7b, 32'hc09c9cb4, 32'hc29866d7, 32'h4291d11a, 32'h42b38ee9};
test_output[6534] = '{32'h42b38ee9};
test_index[6534] = '{7};
test_input[52280:52287] = '{32'hc217108c, 32'hc229767b, 32'hc25bde8d, 32'h427ebc93, 32'hc1ac631d, 32'hc21d62c3, 32'h421be86b, 32'h426e6815};
test_output[6535] = '{32'h427ebc93};
test_index[6535] = '{3};
test_input[52288:52295] = '{32'hc131c13c, 32'h4252efe0, 32'hc2833a22, 32'h41df5952, 32'hc28e41e0, 32'hc223a439, 32'h419bc9a3, 32'h41bdad71};
test_output[6536] = '{32'h4252efe0};
test_index[6536] = '{1};
test_input[52296:52303] = '{32'h41a47a6f, 32'hc2b5a15c, 32'hc19b0f9a, 32'h428f1178, 32'h427f0f78, 32'hc2a812fa, 32'h42282c79, 32'h426cb490};
test_output[6537] = '{32'h428f1178};
test_index[6537] = '{3};
test_input[52304:52311] = '{32'h422debbf, 32'hc212501e, 32'h3fdbf069, 32'hc2bf4c8f, 32'h41240fb6, 32'h411a7e49, 32'hc2bbed09, 32'h42b2a9e6};
test_output[6538] = '{32'h42b2a9e6};
test_index[6538] = '{7};
test_input[52312:52319] = '{32'h423b864f, 32'h422dab4c, 32'h41dc1bc8, 32'hc2bf59c5, 32'hc1b7409b, 32'h42935302, 32'hc1f511be, 32'hc129886a};
test_output[6539] = '{32'h42935302};
test_index[6539] = '{5};
test_input[52320:52327] = '{32'h429402e2, 32'h422a2122, 32'h42b36490, 32'hc28d0c4a, 32'h42b2928c, 32'h42b8ed2a, 32'h42730c69, 32'hc26a4399};
test_output[6540] = '{32'h42b8ed2a};
test_index[6540] = '{5};
test_input[52328:52335] = '{32'hc27c0e1e, 32'hc007c9f7, 32'h406771a5, 32'h42642121, 32'hc2c09239, 32'hbe40a211, 32'h42183d94, 32'h4295e545};
test_output[6541] = '{32'h4295e545};
test_index[6541] = '{7};
test_input[52336:52343] = '{32'hc2499d49, 32'h41f4da1a, 32'hc1fd8db0, 32'h419e6311, 32'hc1fb5104, 32'h423b334b, 32'h427302f4, 32'h42803c69};
test_output[6542] = '{32'h42803c69};
test_index[6542] = '{7};
test_input[52344:52351] = '{32'h4195c5d0, 32'hc205e9e8, 32'h3fb4ae09, 32'h420303e3, 32'h42beda34, 32'hc292e95b, 32'h41c51519, 32'h424c06c1};
test_output[6543] = '{32'h42beda34};
test_index[6543] = '{4};
test_input[52352:52359] = '{32'h42a6dc5f, 32'h41bc179e, 32'h42246c0a, 32'hc2a3367a, 32'hc1debe81, 32'h4212c0c8, 32'hc27a57f4, 32'hc20f8492};
test_output[6544] = '{32'h42a6dc5f};
test_index[6544] = '{0};
test_input[52360:52367] = '{32'hc2b79f64, 32'hc2a16395, 32'hc25c55ce, 32'hbe5cc254, 32'h41c112d7, 32'hc1abca77, 32'h4207ec5b, 32'h426b973f};
test_output[6545] = '{32'h426b973f};
test_index[6545] = '{7};
test_input[52368:52375] = '{32'hc0a0f360, 32'hc2809470, 32'hc080f7bd, 32'h4122406b, 32'h4267915d, 32'h4138d7f7, 32'h427385c0, 32'h420154c6};
test_output[6546] = '{32'h427385c0};
test_index[6546] = '{6};
test_input[52376:52383] = '{32'hc235a28b, 32'hc25d41ce, 32'h42b0b745, 32'h41de28b9, 32'h424e991b, 32'hc2a10e34, 32'hc27952f7, 32'hc215b88c};
test_output[6547] = '{32'h42b0b745};
test_index[6547] = '{2};
test_input[52384:52391] = '{32'h427cf7a5, 32'hc26b8142, 32'hc2b18d18, 32'h428c55f6, 32'hc1bc1ee5, 32'hc2b227e5, 32'h429f758a, 32'hc2870ed5};
test_output[6548] = '{32'h429f758a};
test_index[6548] = '{6};
test_input[52392:52399] = '{32'h3f290afa, 32'hc1ff8dbc, 32'hc18171ca, 32'h420ca173, 32'hc1a69cc7, 32'h424858f6, 32'hc28939c0, 32'hc2b458a6};
test_output[6549] = '{32'h424858f6};
test_index[6549] = '{5};
test_input[52400:52407] = '{32'h41356a19, 32'h427ba0f9, 32'hc2aba393, 32'hc296c55a, 32'h41c1c12a, 32'hc2a7b146, 32'hc2a96da0, 32'hc241f53f};
test_output[6550] = '{32'h427ba0f9};
test_index[6550] = '{1};
test_input[52408:52415] = '{32'hc127463f, 32'h40d88afa, 32'hc1849c93, 32'h41316ed7, 32'hc0d6d83d, 32'h42adcfc7, 32'h4108ba00, 32'h41849e5c};
test_output[6551] = '{32'h42adcfc7};
test_index[6551] = '{5};
test_input[52416:52423] = '{32'hc19f08b0, 32'hc233d153, 32'hc1930b90, 32'h415a008e, 32'h42701fa2, 32'hc18355cf, 32'hc264c4ae, 32'hc1fa45a1};
test_output[6552] = '{32'h42701fa2};
test_index[6552] = '{4};
test_input[52424:52431] = '{32'h429bbf6f, 32'h4286d4b4, 32'hc1120a77, 32'h42121661, 32'hc2aa2dda, 32'hc27cd9ab, 32'h42aaf070, 32'hc200b027};
test_output[6553] = '{32'h42aaf070};
test_index[6553] = '{6};
test_input[52432:52439] = '{32'h42882aad, 32'h414d6e68, 32'h425d4855, 32'hc1786265, 32'h421bf52b, 32'h41c19355, 32'hc2a5cb19, 32'h429eb9f4};
test_output[6554] = '{32'h429eb9f4};
test_index[6554] = '{7};
test_input[52440:52447] = '{32'h4272cff4, 32'h42a76abd, 32'h427759dd, 32'hc2a693c4, 32'hc1b33c99, 32'hc24357d4, 32'h42881e1a, 32'h423d63c1};
test_output[6555] = '{32'h42a76abd};
test_index[6555] = '{1};
test_input[52448:52455] = '{32'h3fd92768, 32'h42b93953, 32'hc2c742d6, 32'hc1c9643b, 32'hc134245e, 32'h425b3875, 32'hc181b5e3, 32'hc0651e5b};
test_output[6556] = '{32'h42b93953};
test_index[6556] = '{1};
test_input[52456:52463] = '{32'h421091ff, 32'h4277e3b1, 32'hc27553ce, 32'h420daae1, 32'hc14f2a33, 32'hc287ed2c, 32'h402bb7d9, 32'h425b5a38};
test_output[6557] = '{32'h4277e3b1};
test_index[6557] = '{1};
test_input[52464:52471] = '{32'hc268e420, 32'hc2af99b6, 32'h42411c59, 32'hc2ba4ea2, 32'h429e102a, 32'h42c07988, 32'h42963a33, 32'hc2b65354};
test_output[6558] = '{32'h42c07988};
test_index[6558] = '{5};
test_input[52472:52479] = '{32'h427f1256, 32'h4298ec5c, 32'hc205f097, 32'hc27a392b, 32'h4297580c, 32'hc292ac54, 32'hc2b91563, 32'h421ba075};
test_output[6559] = '{32'h4298ec5c};
test_index[6559] = '{1};
test_input[52480:52487] = '{32'h42a5e177, 32'hc1926e06, 32'hc294093d, 32'hc183c625, 32'hc21e31fc, 32'h421271c1, 32'h424af730, 32'hc1cb423c};
test_output[6560] = '{32'h42a5e177};
test_index[6560] = '{0};
test_input[52488:52495] = '{32'h4212bd59, 32'hc1118b59, 32'hc0a98e1b, 32'hc0fdb7f1, 32'hc2862d37, 32'hc28405e3, 32'h42a311c6, 32'hc21aa2f5};
test_output[6561] = '{32'h42a311c6};
test_index[6561] = '{6};
test_input[52496:52503] = '{32'hc211f353, 32'h42167e48, 32'hc26c088e, 32'hc0d350c7, 32'h42943c09, 32'h4256c79e, 32'hc2b3933c, 32'h419ea759};
test_output[6562] = '{32'h42943c09};
test_index[6562] = '{4};
test_input[52504:52511] = '{32'h42c63c79, 32'hc2038591, 32'hc1bb7f6b, 32'h427bf369, 32'h423eede6, 32'hc28cb7bf, 32'hc29cec17, 32'h42368aee};
test_output[6563] = '{32'h42c63c79};
test_index[6563] = '{0};
test_input[52512:52519] = '{32'h42b5dfc2, 32'hc1c11240, 32'hc260d253, 32'h41cca397, 32'hc21f764a, 32'hc24180a7, 32'hc1aad5fe, 32'h40d3e36b};
test_output[6564] = '{32'h42b5dfc2};
test_index[6564] = '{0};
test_input[52520:52527] = '{32'hc297f435, 32'h42870329, 32'h428d1e8a, 32'hc225e940, 32'h410e6173, 32'h42bae872, 32'h42b1e93b, 32'hc2242971};
test_output[6565] = '{32'h42bae872};
test_index[6565] = '{5};
test_input[52528:52535] = '{32'h42be109b, 32'h42368e97, 32'h42b8db05, 32'h41807b1e, 32'h41af9242, 32'hc1e80052, 32'h429ebf9e, 32'hc2191265};
test_output[6566] = '{32'h42be109b};
test_index[6566] = '{0};
test_input[52536:52543] = '{32'h42a4e997, 32'hc2a1ca2e, 32'hc2517477, 32'h42087775, 32'hc266f509, 32'h41f408ca, 32'hc1d35fd9, 32'h42bbdd02};
test_output[6567] = '{32'h42bbdd02};
test_index[6567] = '{7};
test_input[52544:52551] = '{32'hc24d2c6b, 32'h418b6bb1, 32'hc0c991da, 32'hc2bb6873, 32'hc15db332, 32'hc28302f1, 32'hc29a856c, 32'h40dd328e};
test_output[6568] = '{32'h418b6bb1};
test_index[6568] = '{1};
test_input[52552:52559] = '{32'hc281e981, 32'h407882f2, 32'hc244af04, 32'hc0d330b6, 32'hc2b9f4ca, 32'h42413457, 32'h41e2bbf5, 32'hc2992b8e};
test_output[6569] = '{32'h42413457};
test_index[6569] = '{5};
test_input[52560:52567] = '{32'hc299dfe8, 32'h428307c5, 32'hc2a2a543, 32'h42693d14, 32'hc2946d2f, 32'hc2b04bf0, 32'hc2b4c328, 32'h417e1c1d};
test_output[6570] = '{32'h428307c5};
test_index[6570] = '{1};
test_input[52568:52575] = '{32'h418571b5, 32'h428063b4, 32'h4074bb84, 32'h42a24617, 32'hc2171a83, 32'hc1b60f61, 32'h422e9331, 32'h4275c842};
test_output[6571] = '{32'h42a24617};
test_index[6571] = '{3};
test_input[52576:52583] = '{32'h3fd990a9, 32'h428a1108, 32'hc25e7abd, 32'h42961544, 32'h41e751d3, 32'h41e1a7ba, 32'h414df60b, 32'hc19edd3b};
test_output[6572] = '{32'h42961544};
test_index[6572] = '{3};
test_input[52584:52591] = '{32'h42799679, 32'hc2b337c2, 32'h42aa7e6e, 32'h42b3a4cb, 32'h4296e968, 32'h4240d783, 32'hc15761db, 32'hc1c1bcae};
test_output[6573] = '{32'h42b3a4cb};
test_index[6573] = '{3};
test_input[52592:52599] = '{32'hc2858021, 32'h42ab22c4, 32'h42806195, 32'h42391b83, 32'hc0d61458, 32'hc2aada8c, 32'h422751bb, 32'hc23ed77c};
test_output[6574] = '{32'h42ab22c4};
test_index[6574] = '{1};
test_input[52600:52607] = '{32'hc20c3662, 32'h428fb09f, 32'hc28aa35d, 32'hc25cd0e8, 32'h42b15b21, 32'h4246afbe, 32'h42af770b, 32'h429c71ba};
test_output[6575] = '{32'h42b15b21};
test_index[6575] = '{4};
test_input[52608:52615] = '{32'h41816c14, 32'hc26430be, 32'h42b9beb1, 32'hc26d8848, 32'hc2a0b15b, 32'hc216461d, 32'hc24d9b52, 32'hc1d5f7a1};
test_output[6576] = '{32'h42b9beb1};
test_index[6576] = '{2};
test_input[52616:52623] = '{32'h42c6329b, 32'hc26c292b, 32'hc2635006, 32'h41248019, 32'h42ba4175, 32'hc25c3123, 32'h422f0393, 32'h42069a50};
test_output[6577] = '{32'h42c6329b};
test_index[6577] = '{0};
test_input[52624:52631] = '{32'hc2aa278d, 32'h4203b608, 32'h423d33d6, 32'hc22c23d4, 32'hc2a19118, 32'h424a2ed6, 32'h41042df5, 32'hc27e90cc};
test_output[6578] = '{32'h424a2ed6};
test_index[6578] = '{5};
test_input[52632:52639] = '{32'hc284657b, 32'hc213f479, 32'hc28f784e, 32'hc191d8c2, 32'hc0cedff5, 32'h40b53baf, 32'h42a2019b, 32'hc29c5d60};
test_output[6579] = '{32'h42a2019b};
test_index[6579] = '{6};
test_input[52640:52647] = '{32'hc2ba8d68, 32'hc2af6283, 32'h426ee072, 32'hc0ec5c8b, 32'hc205e5d4, 32'h4227707e, 32'h420d1e18, 32'h4101ab16};
test_output[6580] = '{32'h426ee072};
test_index[6580] = '{2};
test_input[52648:52655] = '{32'h41844533, 32'h41e955fc, 32'h42475f76, 32'hc09d474a, 32'hc21dbd90, 32'hc1556142, 32'hc1da6383, 32'h420dbd2f};
test_output[6581] = '{32'h42475f76};
test_index[6581] = '{2};
test_input[52656:52663] = '{32'hc29ce2c5, 32'h429dd747, 32'hc266993a, 32'h4272335b, 32'h42646bfb, 32'h412732ad, 32'h421d64fa, 32'h42c65840};
test_output[6582] = '{32'h42c65840};
test_index[6582] = '{7};
test_input[52664:52671] = '{32'hc29aea7f, 32'hc2a90d8b, 32'h42330155, 32'h41b2258b, 32'hc220cfaf, 32'h429f374e, 32'h41b6a684, 32'h428224ad};
test_output[6583] = '{32'h429f374e};
test_index[6583] = '{5};
test_input[52672:52679] = '{32'h414bd9f2, 32'hc2857e8a, 32'h421bbe44, 32'h4293d6cb, 32'h42413873, 32'hc2b40721, 32'hc29d1185, 32'h4265ef69};
test_output[6584] = '{32'h4293d6cb};
test_index[6584] = '{3};
test_input[52680:52687] = '{32'hc2c36d77, 32'h42c03431, 32'h425bab7f, 32'h41e950ab, 32'h402d6a61, 32'hbe608570, 32'h4274a13a, 32'h4234031b};
test_output[6585] = '{32'h42c03431};
test_index[6585] = '{1};
test_input[52688:52695] = '{32'hc26871c6, 32'hc2381aa6, 32'h42a41add, 32'h4080a81c, 32'h410a0c08, 32'h42c1ca6b, 32'hc28d15f6, 32'hc06081d9};
test_output[6586] = '{32'h42c1ca6b};
test_index[6586] = '{5};
test_input[52696:52703] = '{32'hc2830f70, 32'hc24178b6, 32'hc1e9b08d, 32'hc27a4a57, 32'hc256b450, 32'h4157fddd, 32'hc2b42982, 32'h4295c4e1};
test_output[6587] = '{32'h4295c4e1};
test_index[6587] = '{7};
test_input[52704:52711] = '{32'h411f7feb, 32'h42bba10e, 32'hc2a2f4d8, 32'hc17cf9c5, 32'hc2b406c0, 32'h42c70104, 32'h42b7f168, 32'hc226a22a};
test_output[6588] = '{32'h42c70104};
test_index[6588] = '{5};
test_input[52712:52719] = '{32'hc2104bc2, 32'h418e769c, 32'h421b32e4, 32'h428bd678, 32'h42c175a3, 32'hc1f26c2f, 32'hc23b2039, 32'hc1901eef};
test_output[6589] = '{32'h42c175a3};
test_index[6589] = '{4};
test_input[52720:52727] = '{32'hc22f8754, 32'h423b384d, 32'hc29a3682, 32'h42c0e342, 32'h42c490a7, 32'hbfb6d980, 32'hc2c3a402, 32'hc17b48a0};
test_output[6590] = '{32'h42c490a7};
test_index[6590] = '{4};
test_input[52728:52735] = '{32'h42c3ff64, 32'h429f8988, 32'h422c31d1, 32'h42937a6d, 32'h42ad86ea, 32'hc23e1773, 32'h4274cf27, 32'hc2246c8a};
test_output[6591] = '{32'h42c3ff64};
test_index[6591] = '{0};
test_input[52736:52743] = '{32'h421ad20b, 32'h42098509, 32'h428103e3, 32'hc2c1c39d, 32'h42b78deb, 32'hc2a9a04a, 32'h4280aeda, 32'hc206f194};
test_output[6592] = '{32'h42b78deb};
test_index[6592] = '{4};
test_input[52744:52751] = '{32'hc0c166dd, 32'h428bc1cd, 32'h41a512f2, 32'hc00c91ca, 32'hc18ca948, 32'h423f8b26, 32'h421cf402, 32'hc28301e3};
test_output[6593] = '{32'h428bc1cd};
test_index[6593] = '{1};
test_input[52752:52759] = '{32'h4207f32c, 32'h413150bb, 32'hc11d1414, 32'hc2aa2f05, 32'h42aa2e54, 32'hc2360ac2, 32'h417660ee, 32'h428ed456};
test_output[6594] = '{32'h42aa2e54};
test_index[6594] = '{4};
test_input[52760:52767] = '{32'hc293869c, 32'h40b00b30, 32'hc21cc21b, 32'h42aeecdc, 32'h42929121, 32'h4231d672, 32'hc2bcf28b, 32'hc29d50e0};
test_output[6595] = '{32'h42aeecdc};
test_index[6595] = '{3};
test_input[52768:52775] = '{32'hc20892bc, 32'h411ec424, 32'hc2023600, 32'h4284d683, 32'h4272f079, 32'hc24dadac, 32'hc1ff4fe2, 32'h42176781};
test_output[6596] = '{32'h4284d683};
test_index[6596] = '{3};
test_input[52776:52783] = '{32'hc291f19d, 32'h408b4a14, 32'hc25b335a, 32'hc298b6e0, 32'h4299e858, 32'hc1fb1fca, 32'hc22344c1, 32'h41c89a99};
test_output[6597] = '{32'h4299e858};
test_index[6597] = '{4};
test_input[52784:52791] = '{32'hc0ab9358, 32'hc21e012a, 32'h4229d6f9, 32'h3fb52fbb, 32'h424536d0, 32'h42c4b4c0, 32'h40a86e20, 32'hc2397205};
test_output[6598] = '{32'h42c4b4c0};
test_index[6598] = '{5};
test_input[52792:52799] = '{32'hc2a91074, 32'h422e2953, 32'h427ce752, 32'h4270037d, 32'hc2b219c5, 32'h42a795fa, 32'h423231ba, 32'hc2a8a833};
test_output[6599] = '{32'h42a795fa};
test_index[6599] = '{5};
test_input[52800:52807] = '{32'hc1cb4978, 32'hc29d6ef2, 32'h42a3eadb, 32'hc243d0e1, 32'h427d6590, 32'h41b095ff, 32'h403674ee, 32'h425a7ab2};
test_output[6600] = '{32'h42a3eadb};
test_index[6600] = '{2};
test_input[52808:52815] = '{32'h42a6a6de, 32'hc244da46, 32'h429db6b2, 32'hc1db48bc, 32'h420a491c, 32'h426008b6, 32'h4185e322, 32'h42a75e41};
test_output[6601] = '{32'h42a75e41};
test_index[6601] = '{7};
test_input[52816:52823] = '{32'h4205fab4, 32'hc21d9127, 32'h42a3f63c, 32'h40a167b5, 32'h42c33c15, 32'h42049194, 32'h42b6694b, 32'h40b0fb24};
test_output[6602] = '{32'h42c33c15};
test_index[6602] = '{4};
test_input[52824:52831] = '{32'h3e7a639c, 32'hc21543f5, 32'hc23a41a9, 32'hc27bbcba, 32'h42bc8bd4, 32'h42c764f1, 32'hc23f942e, 32'hc05785e8};
test_output[6603] = '{32'h42c764f1};
test_index[6603] = '{5};
test_input[52832:52839] = '{32'hc29abdc1, 32'h427ebb58, 32'h428fbcd9, 32'h42b6f692, 32'h4096a6e7, 32'hbfa54d6d, 32'h41b3c5b7, 32'h41dfabcf};
test_output[6604] = '{32'h42b6f692};
test_index[6604] = '{3};
test_input[52840:52847] = '{32'h4244c90d, 32'hc1ae8878, 32'h42268044, 32'hc2a66506, 32'hc1c6fb0a, 32'h41df810f, 32'hc180f0f5, 32'h41c7e539};
test_output[6605] = '{32'h4244c90d};
test_index[6605] = '{0};
test_input[52848:52855] = '{32'h4125d96c, 32'h42b016a6, 32'h41407eb7, 32'hc17be33d, 32'h41b39d1a, 32'hc2a1d378, 32'hc2b39291, 32'h41154003};
test_output[6606] = '{32'h42b016a6};
test_index[6606] = '{1};
test_input[52856:52863] = '{32'h4223a8ce, 32'hc1c4dcae, 32'hc0313df3, 32'hc0e513f3, 32'hc2b6497c, 32'hc2bb7d84, 32'h4286b9c5, 32'h42bb1073};
test_output[6607] = '{32'h42bb1073};
test_index[6607] = '{7};
test_input[52864:52871] = '{32'hc26d95fb, 32'h42642220, 32'hc192ec3a, 32'h424acdeb, 32'h403be13e, 32'hc1c80647, 32'hc2c1f3c0, 32'hc1ffa6d3};
test_output[6608] = '{32'h42642220};
test_index[6608] = '{1};
test_input[52872:52879] = '{32'h429d529f, 32'hc12b50e1, 32'hc0306c94, 32'hc26af4bb, 32'hc22b33f3, 32'h42befde1, 32'hc2735e2f, 32'h3f207f6b};
test_output[6609] = '{32'h42befde1};
test_index[6609] = '{5};
test_input[52880:52887] = '{32'hc28418c9, 32'h423ba681, 32'hc2bf7e05, 32'hc25054b1, 32'hc2c7e77e, 32'hc198eb17, 32'hc28d1f83, 32'hc28c1726};
test_output[6610] = '{32'h423ba681};
test_index[6610] = '{1};
test_input[52888:52895] = '{32'h42013948, 32'h42ad8ff7, 32'hc183408f, 32'h4263ffdf, 32'h42a5a89a, 32'h418b6c7f, 32'hc2a61f48, 32'h422216b5};
test_output[6611] = '{32'h42ad8ff7};
test_index[6611] = '{1};
test_input[52896:52903] = '{32'h40fd7c80, 32'hc2858a9d, 32'hc283fb1c, 32'h42059a3c, 32'h41538a13, 32'hc2ac5491, 32'h403a4d46, 32'h4249bc2e};
test_output[6612] = '{32'h4249bc2e};
test_index[6612] = '{7};
test_input[52904:52911] = '{32'hc196db8b, 32'h429bcb52, 32'hc2827de1, 32'h4237aaf1, 32'hc26ba0a3, 32'hc2b881ec, 32'h42b0c027, 32'h424b8d72};
test_output[6613] = '{32'h42b0c027};
test_index[6613] = '{6};
test_input[52912:52919] = '{32'hc1ec2805, 32'hc2628295, 32'hc25330e0, 32'hc1fdd7aa, 32'hc1cb077d, 32'hc275e3a1, 32'h424f3442, 32'hc2a3566d};
test_output[6614] = '{32'h424f3442};
test_index[6614] = '{6};
test_input[52920:52927] = '{32'hc28970ec, 32'hc2831189, 32'hbf23334d, 32'h42b2bb29, 32'hc2af9363, 32'hc1e1c260, 32'hc2819ac3, 32'h42c51129};
test_output[6615] = '{32'h42c51129};
test_index[6615] = '{7};
test_input[52928:52935] = '{32'h40f908a5, 32'h416950e8, 32'h42b2c492, 32'h427362dd, 32'hc2a253bc, 32'h424d60e2, 32'hc2bbd7b2, 32'h429e08d4};
test_output[6616] = '{32'h42b2c492};
test_index[6616] = '{2};
test_input[52936:52943] = '{32'hc27cf120, 32'hc26f575a, 32'h41ea37a6, 32'h41f7bce0, 32'h41820450, 32'h4145e717, 32'h42b5392c, 32'hc1def41b};
test_output[6617] = '{32'h42b5392c};
test_index[6617] = '{6};
test_input[52944:52951] = '{32'h4153c706, 32'h425bb5ef, 32'h4195edfe, 32'h41843f2e, 32'h42076502, 32'h418f5e17, 32'hc268d13d, 32'h428b6c47};
test_output[6618] = '{32'h428b6c47};
test_index[6618] = '{7};
test_input[52952:52959] = '{32'h4244cb79, 32'h4123991f, 32'h42bdb423, 32'h42582c92, 32'h4162f19e, 32'h42bec227, 32'hc2541956, 32'h41e529a3};
test_output[6619] = '{32'h42bec227};
test_index[6619] = '{5};
test_input[52960:52967] = '{32'h423a6ad0, 32'hc237ee18, 32'h42079790, 32'hc1b8dcdc, 32'h4221e327, 32'hc1687b76, 32'hc2b6b89b, 32'h42b5bf8e};
test_output[6620] = '{32'h42b5bf8e};
test_index[6620] = '{7};
test_input[52968:52975] = '{32'hc1d5e382, 32'h424aafac, 32'hc1f65972, 32'h41251e7a, 32'hc23872d9, 32'h422fe0bc, 32'hc29ce0b8, 32'h41b1b819};
test_output[6621] = '{32'h424aafac};
test_index[6621] = '{1};
test_input[52976:52983] = '{32'h428dde47, 32'h4068e9a4, 32'hc12f1dec, 32'hc2c3c98c, 32'hc219f763, 32'h41adce27, 32'h41ad9202, 32'hc29f83c3};
test_output[6622] = '{32'h428dde47};
test_index[6622] = '{0};
test_input[52984:52991] = '{32'h40a4b809, 32'hbedc79f1, 32'h4244c5e3, 32'hc2a38d06, 32'h4292e8f4, 32'hc2623272, 32'h42c26fa9, 32'h4273b64d};
test_output[6623] = '{32'h42c26fa9};
test_index[6623] = '{6};
test_input[52992:52999] = '{32'hc19d71f6, 32'hc0af9fec, 32'h42c728e6, 32'hc23dc717, 32'h420f3bd3, 32'hc194f308, 32'h42055f40, 32'h3f96706a};
test_output[6624] = '{32'h42c728e6};
test_index[6624] = '{2};
test_input[53000:53007] = '{32'hc288efa0, 32'hc13db8c7, 32'hc0a3e803, 32'hc2c2882c, 32'h42029881, 32'h4291681d, 32'h42b4cfa7, 32'hc21fedda};
test_output[6625] = '{32'h42b4cfa7};
test_index[6625] = '{6};
test_input[53008:53015] = '{32'hc1e92686, 32'hc183da06, 32'hc092520d, 32'hc2aebb62, 32'hc25e4b0f, 32'h41316cfe, 32'hc2368b9a, 32'h419daf63};
test_output[6626] = '{32'h419daf63};
test_index[6626] = '{7};
test_input[53016:53023] = '{32'hc1c94c9e, 32'hc0e5d786, 32'hc163da04, 32'hc246816f, 32'h42a26a8d, 32'hc27b7940, 32'hc2bf0d57, 32'hc29883d7};
test_output[6627] = '{32'h42a26a8d};
test_index[6627] = '{4};
test_input[53024:53031] = '{32'h42ad0f9e, 32'hc244ee68, 32'h428599d4, 32'h42301f7b, 32'h4256f25d, 32'h41c5c7f6, 32'h41e7341a, 32'hc2b2c61a};
test_output[6628] = '{32'h42ad0f9e};
test_index[6628] = '{0};
test_input[53032:53039] = '{32'hc181ac35, 32'h418d424b, 32'hc269675c, 32'hc26ab530, 32'hc1cbbaa4, 32'hc1b126b1, 32'hc2bc5649, 32'h4262d9d5};
test_output[6629] = '{32'h4262d9d5};
test_index[6629] = '{7};
test_input[53040:53047] = '{32'h41ace6e2, 32'hc2607dc8, 32'h41cd0590, 32'hc1a0d36e, 32'hc2a1b298, 32'hc2b70807, 32'h42bcee01, 32'hc2ae1834};
test_output[6630] = '{32'h42bcee01};
test_index[6630] = '{6};
test_input[53048:53055] = '{32'hc28ce6fe, 32'hc2bcdd67, 32'h42b906f4, 32'h4106e875, 32'h42c75e23, 32'hc286297e, 32'hc28fab4a, 32'hc27bdbca};
test_output[6631] = '{32'h42c75e23};
test_index[6631] = '{4};
test_input[53056:53063] = '{32'h4275409d, 32'h429940ce, 32'h425f605b, 32'h427eec61, 32'hc1c189b3, 32'hc2bc06b1, 32'h4178a951, 32'hc1f49f2c};
test_output[6632] = '{32'h429940ce};
test_index[6632] = '{1};
test_input[53064:53071] = '{32'hc21c7ded, 32'h426e5dfa, 32'hc297c819, 32'hc18d1514, 32'hc2b49794, 32'hc092e5aa, 32'hc29b3ff7, 32'h3f7c9682};
test_output[6633] = '{32'h426e5dfa};
test_index[6633] = '{1};
test_input[53072:53079] = '{32'h40dbf788, 32'hc261b12a, 32'hc1abc83f, 32'h4236c41f, 32'hc276a146, 32'h416c51ef, 32'h4197b445, 32'hc111d2c2};
test_output[6634] = '{32'h4236c41f};
test_index[6634] = '{3};
test_input[53080:53087] = '{32'h428cb3f6, 32'hc2c5b5ce, 32'hc220ef15, 32'h41a172bd, 32'hc2a77795, 32'hc233480f, 32'h42c7805e, 32'h42a236f8};
test_output[6635] = '{32'h42c7805e};
test_index[6635] = '{6};
test_input[53088:53095] = '{32'hc21e697f, 32'h41b75bc2, 32'hc2036805, 32'h419310d3, 32'hc131c433, 32'hc2399061, 32'hc1e90874, 32'hc29995ee};
test_output[6636] = '{32'h41b75bc2};
test_index[6636] = '{1};
test_input[53096:53103] = '{32'h426006c3, 32'hc1cdeaff, 32'hc28cecb1, 32'hc2782173, 32'h42a3ee74, 32'hbfc89581, 32'h42b7d9e8, 32'hc2a3ee76};
test_output[6637] = '{32'h42b7d9e8};
test_index[6637] = '{6};
test_input[53104:53111] = '{32'hc280820e, 32'hc2998eb9, 32'hc25cf370, 32'h424ed4c7, 32'hc2b28527, 32'h42004aab, 32'h426cfb45, 32'hc2aa2547};
test_output[6638] = '{32'h426cfb45};
test_index[6638] = '{6};
test_input[53112:53119] = '{32'hc0f12af0, 32'h425d5243, 32'hc297f6d0, 32'hc2a540f2, 32'h41b232c0, 32'h414c71dd, 32'hc1a955b7, 32'hc1ddc84d};
test_output[6639] = '{32'h425d5243};
test_index[6639] = '{1};
test_input[53120:53127] = '{32'hc1263c6c, 32'h42a83fb4, 32'h42ab4062, 32'h42719592, 32'hc148ee93, 32'h42251600, 32'hc20de419, 32'h41068cd2};
test_output[6640] = '{32'h42ab4062};
test_index[6640] = '{2};
test_input[53128:53135] = '{32'hc286857a, 32'hc284a646, 32'hc2792193, 32'hc1283aaf, 32'h41e8f840, 32'hc1bfe1cc, 32'hc2929c48, 32'hc2c270ba};
test_output[6641] = '{32'h41e8f840};
test_index[6641] = '{4};
test_input[53136:53143] = '{32'hc2aca0b1, 32'hc193c36f, 32'h41d5119b, 32'h4286cb0d, 32'h419b64d6, 32'hc16622f4, 32'hc1bb5de0, 32'h41b2547f};
test_output[6642] = '{32'h4286cb0d};
test_index[6642] = '{3};
test_input[53144:53151] = '{32'h42852e08, 32'h425ec858, 32'hc267b173, 32'h41734f69, 32'hc2508a4b, 32'h41be862d, 32'hc1046867, 32'h429374ea};
test_output[6643] = '{32'h429374ea};
test_index[6643] = '{7};
test_input[53152:53159] = '{32'hc2bb1cc9, 32'h42873511, 32'h42a61e5a, 32'hc184549c, 32'h429a93fd, 32'hc1f85720, 32'h40fb62dd, 32'hc26ecfe4};
test_output[6644] = '{32'h42a61e5a};
test_index[6644] = '{2};
test_input[53160:53167] = '{32'hc29b1086, 32'h42552276, 32'hc29e51b2, 32'h42bc9310, 32'hc2c4b2a9, 32'h429283d0, 32'h415f42bb, 32'hc14cafa8};
test_output[6645] = '{32'h42bc9310};
test_index[6645] = '{3};
test_input[53168:53175] = '{32'hc22a04e3, 32'hc2b61708, 32'hc083ba11, 32'hc2024b09, 32'h42c5864a, 32'h4248c68c, 32'h426d5ce6, 32'hc1d748ac};
test_output[6646] = '{32'h42c5864a};
test_index[6646] = '{4};
test_input[53176:53183] = '{32'h426db0a2, 32'h423c4c2c, 32'hbfec6fc2, 32'hc25fe9f8, 32'h423f6f90, 32'hc194c1d6, 32'hc2aca74b, 32'hc20fa19b};
test_output[6647] = '{32'h426db0a2};
test_index[6647] = '{0};
test_input[53184:53191] = '{32'hc280219b, 32'hc2b68bf8, 32'h428bf96c, 32'hc2b42b66, 32'h429e6aa1, 32'hc28e6e97, 32'h427091bb, 32'hc2c5978d};
test_output[6648] = '{32'h429e6aa1};
test_index[6648] = '{4};
test_input[53192:53199] = '{32'hc275e05f, 32'hc1cf04f2, 32'h4248cd98, 32'hc296ea7c, 32'hc19e803d, 32'h4281d8ff, 32'hc2b71636, 32'hc2b94c4c};
test_output[6649] = '{32'h4281d8ff};
test_index[6649] = '{5};
test_input[53200:53207] = '{32'h42abc321, 32'h41511505, 32'h4217461f, 32'hc16ad73b, 32'h421965fa, 32'h4215c0a2, 32'hc245ec6b, 32'hc18509bf};
test_output[6650] = '{32'h42abc321};
test_index[6650] = '{0};
test_input[53208:53215] = '{32'h42a1752f, 32'hc286c424, 32'hc1cf19ad, 32'hc25fe8c8, 32'h42b21e46, 32'hc25d097e, 32'h42a2270a, 32'hc2c3da9c};
test_output[6651] = '{32'h42b21e46};
test_index[6651] = '{4};
test_input[53216:53223] = '{32'hc28e7e59, 32'h423406de, 32'hc2578cdf, 32'h423eb842, 32'hc238b2cf, 32'hc22c9d98, 32'hc2125b58, 32'hc1a8af5a};
test_output[6652] = '{32'h423eb842};
test_index[6652] = '{3};
test_input[53224:53231] = '{32'hc288d3b0, 32'h42806a21, 32'h414b0fbc, 32'hc082d0e6, 32'h42b3575a, 32'hc2b50c04, 32'h42b1f545, 32'h42ab5bed};
test_output[6653] = '{32'h42b3575a};
test_index[6653] = '{4};
test_input[53232:53239] = '{32'hc23ed5f9, 32'hc1d34ace, 32'h42ad3e3e, 32'hc1cf4cec, 32'hc282711b, 32'hc22bace2, 32'h4295bca6, 32'h41e33680};
test_output[6654] = '{32'h42ad3e3e};
test_index[6654] = '{2};
test_input[53240:53247] = '{32'hc1f2beea, 32'h429b544a, 32'h42307da8, 32'h3f31af5d, 32'hc1a1f357, 32'hc2230704, 32'hc2c470eb, 32'h42b36d27};
test_output[6655] = '{32'h42b36d27};
test_index[6655] = '{7};
test_input[53248:53255] = '{32'hc0f5e890, 32'hc2a2a5c3, 32'hc295e393, 32'h42af1de8, 32'hc2a60b46, 32'hbffc2159, 32'hc2ad401e, 32'hc1921440};
test_output[6656] = '{32'h42af1de8};
test_index[6656] = '{3};
test_input[53256:53263] = '{32'h42c5aedc, 32'hc2a40e09, 32'h419e2b3f, 32'hc2bb3271, 32'hc2981d07, 32'h42309f92, 32'hc185155d, 32'h400e3bd0};
test_output[6657] = '{32'h42c5aedc};
test_index[6657] = '{0};
test_input[53264:53271] = '{32'h41fc3e8c, 32'hc293b8f9, 32'hbf762600, 32'h4245b289, 32'hc2aba8c4, 32'hc27573e1, 32'h41ba5611, 32'hc212253a};
test_output[6658] = '{32'h4245b289};
test_index[6658] = '{3};
test_input[53272:53279] = '{32'h42c5ba03, 32'h425113a3, 32'h41bf452f, 32'h40339d1b, 32'hc297160e, 32'hc248dce1, 32'hc1ecf19e, 32'h413487cd};
test_output[6659] = '{32'h42c5ba03};
test_index[6659] = '{0};
test_input[53280:53287] = '{32'h42c6fc8c, 32'h417dfa56, 32'h42b634ed, 32'h429527ad, 32'h40fa4306, 32'h4115e854, 32'h4282aea6, 32'hc2364a1d};
test_output[6660] = '{32'h42c6fc8c};
test_index[6660] = '{0};
test_input[53288:53295] = '{32'h41b5ed16, 32'h41ed6751, 32'hc1c4a013, 32'h4274ab8b, 32'h425694be, 32'h4233273a, 32'h414aafd9, 32'hc27750bc};
test_output[6661] = '{32'h4274ab8b};
test_index[6661] = '{3};
test_input[53296:53303] = '{32'h429f5c79, 32'hc2b1bd6f, 32'hc22dd633, 32'hc293968f, 32'hc20383f2, 32'hc1ef5fd1, 32'h411ef7e6, 32'hc2723c3c};
test_output[6662] = '{32'h429f5c79};
test_index[6662] = '{0};
test_input[53304:53311] = '{32'h4198b88f, 32'h41a8f11b, 32'h416aae74, 32'hc0a84ca2, 32'hc28f1df3, 32'h41da7fd7, 32'hc27040be, 32'hc2a65421};
test_output[6663] = '{32'h41da7fd7};
test_index[6663] = '{5};
test_input[53312:53319] = '{32'h428384a3, 32'h41fcc4ed, 32'hc2ac781f, 32'hbf90f41e, 32'hc2b571cf, 32'h41221497, 32'hc2c41dd6, 32'hc1e17f77};
test_output[6664] = '{32'h428384a3};
test_index[6664] = '{0};
test_input[53320:53327] = '{32'hc15a37ec, 32'h421c64df, 32'hc11afa93, 32'hc2402bfc, 32'hbfdfa6a3, 32'h4236598b, 32'h421b5e45, 32'hc28365db};
test_output[6665] = '{32'h4236598b};
test_index[6665] = '{5};
test_input[53328:53335] = '{32'hc299832d, 32'hc2aa6a8a, 32'hc2b80b45, 32'hc26bbd63, 32'h429c0a63, 32'h41b07da0, 32'hc02a86a1, 32'h42a29c7a};
test_output[6666] = '{32'h42a29c7a};
test_index[6666] = '{7};
test_input[53336:53343] = '{32'hc2893bdc, 32'h401a9e77, 32'h42c1012e, 32'h41bfccc0, 32'h404db3ff, 32'h4282e74a, 32'hc2808537, 32'hc1f37712};
test_output[6667] = '{32'h42c1012e};
test_index[6667] = '{2};
test_input[53344:53351] = '{32'hc23d7140, 32'h428e8e39, 32'hc2812a22, 32'hc29bea37, 32'hc1a940e0, 32'hc1df0b33, 32'hc20528e5, 32'h42aa08ef};
test_output[6668] = '{32'h42aa08ef};
test_index[6668] = '{7};
test_input[53352:53359] = '{32'hc232538a, 32'h41d09ae0, 32'h41906d66, 32'h3efe4db1, 32'h425b3412, 32'hc2812ab4, 32'h4204b100, 32'h42bf1bfe};
test_output[6669] = '{32'h42bf1bfe};
test_index[6669] = '{7};
test_input[53360:53367] = '{32'h420fda24, 32'hc205e580, 32'hc24d28e5, 32'hc2c0d147, 32'h42904460, 32'h41a206af, 32'h412b1ba7, 32'h42219cb5};
test_output[6670] = '{32'h42904460};
test_index[6670] = '{4};
test_input[53368:53375] = '{32'hc2654073, 32'hc25551ab, 32'hc290d6ce, 32'h42a2a650, 32'hc1a90058, 32'h42be5b72, 32'hc21672f9, 32'hc0d3953c};
test_output[6671] = '{32'h42be5b72};
test_index[6671] = '{5};
test_input[53376:53383] = '{32'h42683a2d, 32'hc2443d31, 32'h42989b5f, 32'h42acebaa, 32'h4236a9f5, 32'h3fee8c20, 32'hc15ea2a2, 32'h42b68dc3};
test_output[6672] = '{32'h42b68dc3};
test_index[6672] = '{7};
test_input[53384:53391] = '{32'h411e3cf7, 32'h42a8070f, 32'hc23b6e43, 32'hc157898b, 32'h4202bc72, 32'h4222bbc8, 32'hc2901c32, 32'hc12a76d2};
test_output[6673] = '{32'h42a8070f};
test_index[6673] = '{1};
test_input[53392:53399] = '{32'hc10d53f2, 32'h4092103b, 32'h42c688fd, 32'h42c49d4c, 32'hc25d6ff7, 32'h40c6443f, 32'hc290cebf, 32'h421d29db};
test_output[6674] = '{32'h42c688fd};
test_index[6674] = '{2};
test_input[53400:53407] = '{32'hc2b14801, 32'h424288da, 32'hbf14d763, 32'h41fb2f52, 32'hc242ae33, 32'h4298a440, 32'h41b97dd0, 32'hc284709b};
test_output[6675] = '{32'h4298a440};
test_index[6675] = '{5};
test_input[53408:53415] = '{32'h3dfa7b7e, 32'hc245555e, 32'hc237204c, 32'hc2b5618f, 32'hc2976adf, 32'h4062ba8f, 32'h423393cd, 32'hc1c1a287};
test_output[6676] = '{32'h423393cd};
test_index[6676] = '{6};
test_input[53416:53423] = '{32'h424d40e2, 32'h42c4a059, 32'hc2333680, 32'h42afb119, 32'hc2c0e169, 32'h41a9d934, 32'h42bae76b, 32'h42a559f0};
test_output[6677] = '{32'h42c4a059};
test_index[6677] = '{1};
test_input[53424:53431] = '{32'hc2b6ef2a, 32'hbd49c648, 32'h419947ba, 32'h41a8cba7, 32'h42403934, 32'hc17bbd39, 32'hc2aa4951, 32'h4282eca1};
test_output[6678] = '{32'h4282eca1};
test_index[6678] = '{7};
test_input[53432:53439] = '{32'h42c103bf, 32'hc2c6d869, 32'hc1c58e65, 32'hc1b9a7d2, 32'hc25ec8c4, 32'h42a4c41c, 32'h41af5f53, 32'hbf05fdfc};
test_output[6679] = '{32'h42c103bf};
test_index[6679] = '{0};
test_input[53440:53447] = '{32'h4191ded4, 32'h428458b9, 32'hc290d75d, 32'h42ac2a6c, 32'hc1e308ec, 32'h424dfaeb, 32'h4273019d, 32'h42021084};
test_output[6680] = '{32'h42ac2a6c};
test_index[6680] = '{3};
test_input[53448:53455] = '{32'h424748dd, 32'hc1282ce3, 32'h40e51dcc, 32'h41fa716f, 32'h428fa5e7, 32'hc2c4907b, 32'hc0dfead6, 32'h422e4ad3};
test_output[6681] = '{32'h428fa5e7};
test_index[6681] = '{4};
test_input[53456:53463] = '{32'hc2bb19d8, 32'hc21a6793, 32'hc2120934, 32'h424ad271, 32'hc12ddf36, 32'hc2a69cfd, 32'hc1830f84, 32'hc14ce47b};
test_output[6682] = '{32'h424ad271};
test_index[6682] = '{3};
test_input[53464:53471] = '{32'hc29d3281, 32'h425e1783, 32'hc2b2d8dd, 32'hc2c1dd9a, 32'h40b0c481, 32'hc28d74e7, 32'h41a89cb4, 32'hc205a6ec};
test_output[6683] = '{32'h425e1783};
test_index[6683] = '{1};
test_input[53472:53479] = '{32'h42a14c21, 32'hc0ff1fab, 32'h4283e01e, 32'h425a0cd9, 32'hc273927d, 32'h42c646d1, 32'hc2a5ad53, 32'h42a4c3dc};
test_output[6684] = '{32'h42c646d1};
test_index[6684] = '{5};
test_input[53480:53487] = '{32'h4296e946, 32'hc1065ec8, 32'h42a6bd6d, 32'hc219711b, 32'hc2b35cfb, 32'h4121a236, 32'hc18bb4dd, 32'hc1a79fce};
test_output[6685] = '{32'h42a6bd6d};
test_index[6685] = '{2};
test_input[53488:53495] = '{32'hc2c73a5a, 32'hc2b21edc, 32'hc01bac11, 32'h42afa2fa, 32'hc20b3abd, 32'h412343bc, 32'hc1d13d41, 32'hc1b3fe39};
test_output[6686] = '{32'h42afa2fa};
test_index[6686] = '{3};
test_input[53496:53503] = '{32'h4230675b, 32'h41ba29b8, 32'hc2824bc6, 32'hc1497b63, 32'h402195db, 32'h40e21ef2, 32'h41d83532, 32'hc15d01cc};
test_output[6687] = '{32'h4230675b};
test_index[6687] = '{0};
test_input[53504:53511] = '{32'hc29eeeff, 32'hc223c2e5, 32'h420f5f98, 32'h41e5fd2c, 32'hc2063cc9, 32'h42be8e6e, 32'h42a73428, 32'h42ac0450};
test_output[6688] = '{32'h42be8e6e};
test_index[6688] = '{5};
test_input[53512:53519] = '{32'hc293829e, 32'hc2bf77a4, 32'hc096c2c3, 32'hc29a3b56, 32'hc21f38c2, 32'h42261c13, 32'h42b5578b, 32'h427b3978};
test_output[6689] = '{32'h42b5578b};
test_index[6689] = '{6};
test_input[53520:53527] = '{32'hc11fed7d, 32'hc07a8c7a, 32'hc279379d, 32'h426186de, 32'hc29f0b97, 32'hc23af6db, 32'h42ac0e8b, 32'hc1f753b1};
test_output[6690] = '{32'h42ac0e8b};
test_index[6690] = '{6};
test_input[53528:53535] = '{32'hc2abeb56, 32'hc2303ea9, 32'hc2193409, 32'hc205187c, 32'h424a5602, 32'hc2ab8296, 32'h4146d280, 32'h4287d278};
test_output[6691] = '{32'h4287d278};
test_index[6691] = '{7};
test_input[53536:53543] = '{32'hc266cdb0, 32'hc13cad42, 32'h42ac6214, 32'h428e4e2f, 32'h41c2adef, 32'hc2b82db1, 32'h423cd6b3, 32'h410462bc};
test_output[6692] = '{32'h42ac6214};
test_index[6692] = '{2};
test_input[53544:53551] = '{32'hc0d5e5fc, 32'hbb0e6540, 32'h41fea7b9, 32'hc1590c25, 32'hc1e99af4, 32'hc2452389, 32'h4233c4ea, 32'hc182739f};
test_output[6693] = '{32'h4233c4ea};
test_index[6693] = '{6};
test_input[53552:53559] = '{32'hc252b747, 32'h401d0960, 32'h417f7d40, 32'hc29b377c, 32'hc05c93ba, 32'hc2512478, 32'hc2625f93, 32'h42b010f5};
test_output[6694] = '{32'h42b010f5};
test_index[6694] = '{7};
test_input[53560:53567] = '{32'h42bd80ad, 32'h42b631af, 32'h41ddcd10, 32'hc2a6d29c, 32'h428a19cd, 32'hc2a6e7c1, 32'h42b1fab2, 32'hc0bdbc1e};
test_output[6695] = '{32'h42bd80ad};
test_index[6695] = '{0};
test_input[53568:53575] = '{32'h4285d1e9, 32'h41332805, 32'h41db6e60, 32'hc25be1d7, 32'hc1cf440e, 32'h41d5413c, 32'hc243aede, 32'hc209fa25};
test_output[6696] = '{32'h4285d1e9};
test_index[6696] = '{0};
test_input[53576:53583] = '{32'hc1f3e789, 32'h4236d1fa, 32'h41fe699d, 32'h4107c530, 32'h42115a2b, 32'h422f4447, 32'h412f1adf, 32'h419ec64f};
test_output[6697] = '{32'h4236d1fa};
test_index[6697] = '{1};
test_input[53584:53591] = '{32'hc24e6d34, 32'hc1e5a1eb, 32'h428ead18, 32'hc220a7ec, 32'h422063db, 32'hc2a828fe, 32'hc1236856, 32'hc2c37695};
test_output[6698] = '{32'h428ead18};
test_index[6698] = '{2};
test_input[53592:53599] = '{32'hc2a449db, 32'h41fb548e, 32'hc25463a5, 32'hc2a0c4a0, 32'hc28328db, 32'h42966b6b, 32'h42b38af2, 32'hc22e08e2};
test_output[6699] = '{32'h42b38af2};
test_index[6699] = '{6};
test_input[53600:53607] = '{32'hc1dad69e, 32'h40ce9db8, 32'h42118489, 32'hc292ca2e, 32'hc1e7ffcc, 32'hc28d310b, 32'h40b76282, 32'hc2a31078};
test_output[6700] = '{32'h42118489};
test_index[6700] = '{2};
test_input[53608:53615] = '{32'hc2b7509c, 32'h41e281a0, 32'h42040c53, 32'h405a15f6, 32'h4253cbd6, 32'h41d394a8, 32'hc19038dc, 32'h416d2a11};
test_output[6701] = '{32'h4253cbd6};
test_index[6701] = '{4};
test_input[53616:53623] = '{32'hc29d820b, 32'hc2017198, 32'hc288730c, 32'hc1e6d800, 32'hc26f0c16, 32'h418fc094, 32'h42b15e69, 32'hc28510cb};
test_output[6702] = '{32'h42b15e69};
test_index[6702] = '{6};
test_input[53624:53631] = '{32'h42183558, 32'h420147e6, 32'hc291ab39, 32'hc218e0e6, 32'hc2191136, 32'hc262f375, 32'h428450f3, 32'h40f4d8af};
test_output[6703] = '{32'h428450f3};
test_index[6703] = '{6};
test_input[53632:53639] = '{32'hc2c76765, 32'h4289ce9f, 32'h429d3cce, 32'hc29ba7a5, 32'hc227cca5, 32'hc2639e82, 32'hc294d4f6, 32'hc2446e4d};
test_output[6704] = '{32'h429d3cce};
test_index[6704] = '{2};
test_input[53640:53647] = '{32'h416bde00, 32'h427d0fdb, 32'hc2bba1af, 32'hc29b682b, 32'hc2c2ed3e, 32'h40962633, 32'hc29ad2f8, 32'h4195ba2b};
test_output[6705] = '{32'h427d0fdb};
test_index[6705] = '{1};
test_input[53648:53655] = '{32'hc2b883c0, 32'h411ff0cd, 32'hc2bd7864, 32'h42865994, 32'h41c1300e, 32'hc270ec19, 32'h42aa95c0, 32'h42917654};
test_output[6706] = '{32'h42aa95c0};
test_index[6706] = '{6};
test_input[53656:53663] = '{32'hc282e406, 32'h41c117ef, 32'hc2aac474, 32'h408f4455, 32'hc2812aa2, 32'hc1a6f552, 32'h428259b9, 32'hc298cec0};
test_output[6707] = '{32'h428259b9};
test_index[6707] = '{6};
test_input[53664:53671] = '{32'hc1afeb64, 32'hc27ffba8, 32'hc1963dd4, 32'hc289b674, 32'h424b5b13, 32'h42497b18, 32'h42c133fd, 32'h4288cd60};
test_output[6708] = '{32'h42c133fd};
test_index[6708] = '{6};
test_input[53672:53679] = '{32'hc1b9c11c, 32'hc2628f2d, 32'h419d8d07, 32'hc1b5de9d, 32'hc2bfac28, 32'hc294598f, 32'hc1fbb5c5, 32'hc2bbf233};
test_output[6709] = '{32'h419d8d07};
test_index[6709] = '{2};
test_input[53680:53687] = '{32'hc22092a5, 32'h42a2a802, 32'h4214bcbb, 32'h42574e5e, 32'h4282acb0, 32'hc1746eb6, 32'hc298beb8, 32'hc2c29196};
test_output[6710] = '{32'h42a2a802};
test_index[6710] = '{1};
test_input[53688:53695] = '{32'hc23a5ea2, 32'h429477ba, 32'h428b5514, 32'hc2a6133e, 32'hc1a72caa, 32'h41117238, 32'hc21aba99, 32'hc2bc1e66};
test_output[6711] = '{32'h429477ba};
test_index[6711] = '{1};
test_input[53696:53703] = '{32'h428fbab8, 32'hc2c1fb46, 32'hc0f326bb, 32'hc2c15ab7, 32'hc282eb09, 32'hc2831a35, 32'h416ff110, 32'h422fb19e};
test_output[6712] = '{32'h428fbab8};
test_index[6712] = '{0};
test_input[53704:53711] = '{32'h4282cea5, 32'hc26fde4b, 32'h42814f75, 32'hc2afb990, 32'h42557859, 32'hc13d5d87, 32'hc223c2a4, 32'h421ba2ed};
test_output[6713] = '{32'h4282cea5};
test_index[6713] = '{0};
test_input[53712:53719] = '{32'hc19c89f9, 32'h421b57da, 32'hc25686c0, 32'h41ccce73, 32'h409bae64, 32'h422fe0ae, 32'hc287027e, 32'h4263238e};
test_output[6714] = '{32'h4263238e};
test_index[6714] = '{7};
test_input[53720:53727] = '{32'h4153facd, 32'hc2bdfa68, 32'h42679a1b, 32'h4246366b, 32'h41fb5214, 32'hc0f208b8, 32'hc0b09cae, 32'hc2454294};
test_output[6715] = '{32'h42679a1b};
test_index[6715] = '{2};
test_input[53728:53735] = '{32'hc257e247, 32'hc0867d7e, 32'h4293faf8, 32'hc15a5777, 32'hc29dc3cd, 32'h42ad714f, 32'h42a4bf7f, 32'h42afc0ef};
test_output[6716] = '{32'h42afc0ef};
test_index[6716] = '{7};
test_input[53736:53743] = '{32'h4265ab4a, 32'h4271f490, 32'h42c30645, 32'hc2165cee, 32'hc1e4abc6, 32'h4278e0bc, 32'h422da8cd, 32'h42b586a5};
test_output[6717] = '{32'h42c30645};
test_index[6717] = '{2};
test_input[53744:53751] = '{32'hc1da9484, 32'h409ec341, 32'hc255b871, 32'hc2c69f83, 32'h4246379a, 32'h42bd94b3, 32'hc2719673, 32'hc2846682};
test_output[6718] = '{32'h42bd94b3};
test_index[6718] = '{5};
test_input[53752:53759] = '{32'h42a60c76, 32'h41c131f1, 32'hc18cb8d8, 32'h41268e20, 32'hc2baea05, 32'h4289b309, 32'h4288998c, 32'hc285966d};
test_output[6719] = '{32'h42a60c76};
test_index[6719] = '{0};
test_input[53760:53767] = '{32'hc261b409, 32'h42bb5037, 32'h4222f0ef, 32'hc14b55ba, 32'hc293f165, 32'h419d47dd, 32'hc24e68fd, 32'h42993fd0};
test_output[6720] = '{32'h42bb5037};
test_index[6720] = '{1};
test_input[53768:53775] = '{32'h41200c33, 32'hc154d268, 32'hc23d4f2b, 32'hc26efbd8, 32'h42c7ec35, 32'h42699893, 32'h42b07d28, 32'h42758db0};
test_output[6721] = '{32'h42c7ec35};
test_index[6721] = '{4};
test_input[53776:53783] = '{32'h4284dc25, 32'h42c14e04, 32'hc20e6a50, 32'hc2a76ee6, 32'h4293c5aa, 32'hc1b55276, 32'h41f4b89b, 32'h42892832};
test_output[6722] = '{32'h42c14e04};
test_index[6722] = '{1};
test_input[53784:53791] = '{32'hc23d0c72, 32'hc2bc0252, 32'h429ccba8, 32'hc297b670, 32'h42041da8, 32'hc17fdb51, 32'hc2b99f76, 32'hc1214094};
test_output[6723] = '{32'h429ccba8};
test_index[6723] = '{2};
test_input[53792:53799] = '{32'h42988f79, 32'hc14a5db4, 32'hc255a5b2, 32'h422c21a5, 32'hc25c5ec1, 32'h42a3de95, 32'h40f511ad, 32'h427280f6};
test_output[6724] = '{32'h42a3de95};
test_index[6724] = '{5};
test_input[53800:53807] = '{32'h4229b2f4, 32'h4291c9b6, 32'h425cc106, 32'hc28e3c91, 32'hc112bf1a, 32'h42438a51, 32'h428c2744, 32'h42a52332};
test_output[6725] = '{32'h42a52332};
test_index[6725] = '{7};
test_input[53808:53815] = '{32'hc0c617c2, 32'h427bdb96, 32'h42349dec, 32'hc1d20f6c, 32'hc2c21b04, 32'h421b1444, 32'hc05c6b79, 32'hc2160c0e};
test_output[6726] = '{32'h427bdb96};
test_index[6726] = '{1};
test_input[53816:53823] = '{32'hc2b8cdd5, 32'hc2976810, 32'hc28cc586, 32'hc1a27305, 32'hc297a753, 32'h41ab4b32, 32'hc20f57a9, 32'h42ba67fb};
test_output[6727] = '{32'h42ba67fb};
test_index[6727] = '{7};
test_input[53824:53831] = '{32'h41947a96, 32'hc1871f1f, 32'hc1bbf9c8, 32'hbfa1ba53, 32'h428ac7e4, 32'hc0701c2c, 32'hc0538381, 32'h419b4452};
test_output[6728] = '{32'h428ac7e4};
test_index[6728] = '{4};
test_input[53832:53839] = '{32'h4253237b, 32'hc22919f3, 32'h42124765, 32'h42869fe6, 32'h41926e82, 32'h41e857a7, 32'h421295f0, 32'hc1da9839};
test_output[6729] = '{32'h42869fe6};
test_index[6729] = '{3};
test_input[53840:53847] = '{32'h420f9685, 32'h41ef4a02, 32'hc28064d1, 32'h4265223d, 32'hc2148867, 32'hc282fbd3, 32'hc1a35a2f, 32'hc22e0a66};
test_output[6730] = '{32'h4265223d};
test_index[6730] = '{3};
test_input[53848:53855] = '{32'h424a6170, 32'h4105aa80, 32'h42c23509, 32'hc1d40d54, 32'hc2b6e043, 32'hc2c0dca9, 32'hc29ebbfb, 32'hc26f7d18};
test_output[6731] = '{32'h42c23509};
test_index[6731] = '{2};
test_input[53856:53863] = '{32'hc2a363c1, 32'h4287484c, 32'hc25fb689, 32'h42931296, 32'h40c230e2, 32'hc20e73ea, 32'h425f860a, 32'h424e8edf};
test_output[6732] = '{32'h42931296};
test_index[6732] = '{3};
test_input[53864:53871] = '{32'hc294eca4, 32'hc226fbdb, 32'hc29e1795, 32'hc23e277c, 32'hc22f1352, 32'h4280861d, 32'hc10f149e, 32'hc2ad2ba4};
test_output[6733] = '{32'h4280861d};
test_index[6733] = '{5};
test_input[53872:53879] = '{32'h42506075, 32'hc0165680, 32'hc110ca6a, 32'hc269ac36, 32'hc2c63d27, 32'hc1ae4797, 32'h4118f45c, 32'hc21999b9};
test_output[6734] = '{32'h42506075};
test_index[6734] = '{0};
test_input[53880:53887] = '{32'h42131dd6, 32'hc0ba5a69, 32'h42307215, 32'hc200da23, 32'h4246b609, 32'h4274d846, 32'hc286af5d, 32'hc11e3525};
test_output[6735] = '{32'h4274d846};
test_index[6735] = '{5};
test_input[53888:53895] = '{32'h426eaf47, 32'h42be4eab, 32'h42ac23dd, 32'h422c23d3, 32'hc17e7606, 32'hc2c25f57, 32'h426dad24, 32'h422da17f};
test_output[6736] = '{32'h42be4eab};
test_index[6736] = '{1};
test_input[53896:53903] = '{32'h426ad505, 32'hc2af59ca, 32'h42890131, 32'h4245f5c1, 32'hc2b1e81e, 32'hc282232c, 32'hc2085328, 32'hc2a2dec5};
test_output[6737] = '{32'h42890131};
test_index[6737] = '{2};
test_input[53904:53911] = '{32'hc29242ea, 32'hc15841a4, 32'hc2bbb25d, 32'hc20bc3c5, 32'hc26e37bd, 32'hc19fec0f, 32'h41cf2aa3, 32'h42a79153};
test_output[6738] = '{32'h42a79153};
test_index[6738] = '{7};
test_input[53912:53919] = '{32'h42521f1b, 32'hc128cf3b, 32'h4299ddc3, 32'h4275089a, 32'hc137d274, 32'hc148d9d9, 32'hc2956203, 32'hc24a34e1};
test_output[6739] = '{32'h4299ddc3};
test_index[6739] = '{2};
test_input[53920:53927] = '{32'hc29b0645, 32'hc14837ed, 32'hc199dd6c, 32'hc1b29440, 32'h421b0726, 32'hbfcb49be, 32'hc0eee35e, 32'h42a3374e};
test_output[6740] = '{32'h42a3374e};
test_index[6740] = '{7};
test_input[53928:53935] = '{32'hc198e88b, 32'h42b14bfa, 32'hc143588e, 32'hc118f1eb, 32'hc24281b3, 32'h428e77df, 32'hc14bfa2e, 32'hc2c7c698};
test_output[6741] = '{32'h42b14bfa};
test_index[6741] = '{1};
test_input[53936:53943] = '{32'h42866ac0, 32'h42a9a5da, 32'h402885fb, 32'hc1aa7468, 32'hbfeb5533, 32'h428e89dc, 32'h4298a07b, 32'h42821412};
test_output[6742] = '{32'h42a9a5da};
test_index[6742] = '{1};
test_input[53944:53951] = '{32'h41cfdfa8, 32'h4234444d, 32'h4281cd8b, 32'h41b74743, 32'hc22daadc, 32'hc298b8c9, 32'hc22d18e7, 32'h424d8998};
test_output[6743] = '{32'h4281cd8b};
test_index[6743] = '{2};
test_input[53952:53959] = '{32'hc2379eee, 32'hc27e25e7, 32'hc13d1383, 32'h42be64cd, 32'h42bef3f4, 32'h42a9c80e, 32'h427ce2c5, 32'h42581589};
test_output[6744] = '{32'h42bef3f4};
test_index[6744] = '{4};
test_input[53960:53967] = '{32'h42a80159, 32'h41c8895c, 32'h426b53a2, 32'hc2a817a4, 32'h42848ba1, 32'h41bc8706, 32'hc28bdda8, 32'hc2117f74};
test_output[6745] = '{32'h42a80159};
test_index[6745] = '{0};
test_input[53968:53975] = '{32'h4291b4f6, 32'h424270ef, 32'h41dad001, 32'hc1974b92, 32'h42bdbaaf, 32'h429731a0, 32'hc12975d7, 32'h3f707f3a};
test_output[6746] = '{32'h42bdbaaf};
test_index[6746] = '{4};
test_input[53976:53983] = '{32'h423ac689, 32'h429bfe5b, 32'h4294b6da, 32'hc13c2873, 32'h41bcff2b, 32'h42c55c6e, 32'h41e712ee, 32'hc2afe29c};
test_output[6747] = '{32'h42c55c6e};
test_index[6747] = '{5};
test_input[53984:53991] = '{32'h42ba1bbf, 32'hc187abf5, 32'hc234fb41, 32'hc13b0ad6, 32'h422378b3, 32'h41b5d3e9, 32'hc23091a9, 32'h413d0418};
test_output[6748] = '{32'h42ba1bbf};
test_index[6748] = '{0};
test_input[53992:53999] = '{32'hc2478316, 32'h426eac70, 32'hc2950191, 32'hc26d7d7e, 32'h4137124f, 32'h42bc1442, 32'h4051947f, 32'hc2b160c1};
test_output[6749] = '{32'h42bc1442};
test_index[6749] = '{5};
test_input[54000:54007] = '{32'h417306ac, 32'hc28f139c, 32'h41da6cb6, 32'hc2bd21f5, 32'hc2a71931, 32'hc2b08f30, 32'h420522bf, 32'hc2b736c5};
test_output[6750] = '{32'h420522bf};
test_index[6750] = '{6};
test_input[54008:54015] = '{32'h419b5139, 32'hc2537abb, 32'hbf71fa04, 32'hc208dd2b, 32'h418c8cf2, 32'h42575158, 32'hc2319ecc, 32'h42b95fef};
test_output[6751] = '{32'h42b95fef};
test_index[6751] = '{7};
test_input[54016:54023] = '{32'hc27ef817, 32'h428fa4bd, 32'h4288ef49, 32'h40a81590, 32'h42bad278, 32'hc2abdc99, 32'h428f565e, 32'hc249a4f8};
test_output[6752] = '{32'h42bad278};
test_index[6752] = '{4};
test_input[54024:54031] = '{32'h421583f0, 32'hc28e4dd7, 32'hc2a89004, 32'h42886344, 32'hc26a5b83, 32'hc1afa94e, 32'h42186884, 32'hc22a59c4};
test_output[6753] = '{32'h42886344};
test_index[6753] = '{3};
test_input[54032:54039] = '{32'h41e5efdd, 32'hc1ff14f4, 32'hc286d1d6, 32'h4010898a, 32'h4252dda3, 32'hc288ef2b, 32'h4240c6a0, 32'hc156629e};
test_output[6754] = '{32'h4252dda3};
test_index[6754] = '{4};
test_input[54040:54047] = '{32'h41022ab6, 32'h429bdea9, 32'hc28e12ba, 32'h419b39cd, 32'h425a15e1, 32'h41c1ea97, 32'h41658086, 32'h42882a79};
test_output[6755] = '{32'h429bdea9};
test_index[6755] = '{1};
test_input[54048:54055] = '{32'hc0e2d667, 32'h42692956, 32'hc2407930, 32'h420a70bd, 32'hc04f7ca9, 32'h42bc0206, 32'h421a41c7, 32'h42a0b23d};
test_output[6756] = '{32'h42bc0206};
test_index[6756] = '{5};
test_input[54056:54063] = '{32'h42c471f2, 32'hc2c30f18, 32'hc269a62b, 32'hc2011f81, 32'hc2827eb9, 32'hc25dc847, 32'hc0fb0ca8, 32'hc15501ea};
test_output[6757] = '{32'h42c471f2};
test_index[6757] = '{0};
test_input[54064:54071] = '{32'h41cb77ff, 32'h40ccc5b5, 32'h41be9eb0, 32'h41f41643, 32'h426464be, 32'h41f33e81, 32'h42b24c3f, 32'hc2b5bcae};
test_output[6758] = '{32'h42b24c3f};
test_index[6758] = '{6};
test_input[54072:54079] = '{32'h42ac4003, 32'hc22329f3, 32'hc24b9668, 32'h419e557f, 32'hc27e75b8, 32'h42bbacc3, 32'hc229ebae, 32'hc186c263};
test_output[6759] = '{32'h42bbacc3};
test_index[6759] = '{5};
test_input[54080:54087] = '{32'hc271788e, 32'h40e10bbf, 32'hbee264bd, 32'hc247418c, 32'h418b9ab4, 32'h428aca5d, 32'hc2850ae8, 32'hc267fe46};
test_output[6760] = '{32'h428aca5d};
test_index[6760] = '{5};
test_input[54088:54095] = '{32'h42851012, 32'hc216e3dc, 32'h42670d12, 32'hc02d6745, 32'h42099ff2, 32'h427eb67d, 32'h425232b8, 32'h42069231};
test_output[6761] = '{32'h42851012};
test_index[6761] = '{0};
test_input[54096:54103] = '{32'h42497537, 32'hc286708d, 32'hc298c5e8, 32'hc12332b8, 32'hc23b463e, 32'hc1306272, 32'hc2c0b2b8, 32'hc18bb277};
test_output[6762] = '{32'h42497537};
test_index[6762] = '{0};
test_input[54104:54111] = '{32'hc2632f11, 32'hc28e0fd4, 32'hc24bf9f4, 32'h42332dad, 32'h4210f01b, 32'hc2705155, 32'hc2937666, 32'h423e1ef3};
test_output[6763] = '{32'h423e1ef3};
test_index[6763] = '{7};
test_input[54112:54119] = '{32'h4194bb23, 32'h3fbefe9c, 32'hc2407518, 32'h42220e3e, 32'hc0e527bc, 32'h427d78ab, 32'hc1efddae, 32'h42959a67};
test_output[6764] = '{32'h42959a67};
test_index[6764] = '{7};
test_input[54120:54127] = '{32'h41fd500f, 32'hc293a455, 32'hbfce6edd, 32'hc2b14cf6, 32'h4286ee08, 32'hc247b026, 32'hc2175fd8, 32'hc2c06956};
test_output[6765] = '{32'h4286ee08};
test_index[6765] = '{4};
test_input[54128:54135] = '{32'hc2900fc7, 32'h40cc13a4, 32'hc2c45b0a, 32'hc2b1cdd6, 32'hc2081fc8, 32'h42af3e4d, 32'h42bbf7b8, 32'h4277d11b};
test_output[6766] = '{32'h42bbf7b8};
test_index[6766] = '{6};
test_input[54136:54143] = '{32'hc27b50ed, 32'h425bd40d, 32'h41e5d6b1, 32'h41963d7f, 32'hc080916b, 32'hc239c9a1, 32'h429bd40b, 32'h4201173b};
test_output[6767] = '{32'h429bd40b};
test_index[6767] = '{6};
test_input[54144:54151] = '{32'h427852ec, 32'hc2a1751d, 32'hc16bce73, 32'hc20a5e7e, 32'hc26ef8ae, 32'hc2b765e8, 32'hc11d570f, 32'h42029d94};
test_output[6768] = '{32'h427852ec};
test_index[6768] = '{0};
test_input[54152:54159] = '{32'hc123926e, 32'hc2c16d39, 32'h410ab779, 32'hc192772e, 32'h41b96dbd, 32'h4117eea1, 32'h42babe4b, 32'hc2624cfe};
test_output[6769] = '{32'h42babe4b};
test_index[6769] = '{6};
test_input[54160:54167] = '{32'h41012735, 32'h428ee59e, 32'hc194bfb4, 32'h42679a95, 32'hc2ad9b23, 32'h42a1022d, 32'hc1f2b1d7, 32'hc29f6bd3};
test_output[6770] = '{32'h42a1022d};
test_index[6770] = '{5};
test_input[54168:54175] = '{32'hc297844e, 32'h4289b27a, 32'h42a898e9, 32'h42a3dde2, 32'h42485e4c, 32'h418a968f, 32'hc224b3d2, 32'h4282e50c};
test_output[6771] = '{32'h42a898e9};
test_index[6771] = '{2};
test_input[54176:54183] = '{32'hc25dd766, 32'h41ef25a0, 32'h424d42d8, 32'hc2949ee4, 32'h3f7b7047, 32'h41aebed5, 32'hc2acde44, 32'h41c04b7e};
test_output[6772] = '{32'h424d42d8};
test_index[6772] = '{2};
test_input[54184:54191] = '{32'hc2653639, 32'hc2122bd9, 32'h412d432c, 32'hc2148bd0, 32'hc28c6e3b, 32'h42772092, 32'hc1a9c48b, 32'hc2a18571};
test_output[6773] = '{32'h42772092};
test_index[6773] = '{5};
test_input[54192:54199] = '{32'hc2c65468, 32'hc27e7239, 32'hc2243e06, 32'h42a29019, 32'h41a834a2, 32'h4226d921, 32'hc2b3b2a7, 32'h42021fce};
test_output[6774] = '{32'h42a29019};
test_index[6774] = '{3};
test_input[54200:54207] = '{32'h41c1c0f8, 32'h42a9e1d4, 32'h4222b73f, 32'h41829707, 32'hc267f4d9, 32'h42931c49, 32'hc1fed877, 32'hc24304c1};
test_output[6775] = '{32'h42a9e1d4};
test_index[6775] = '{1};
test_input[54208:54215] = '{32'hc1a9048c, 32'hc236d827, 32'hc2820a02, 32'h41fe7f37, 32'hc2a41a10, 32'h42a33e05, 32'hc16dd06f, 32'hc207dada};
test_output[6776] = '{32'h42a33e05};
test_index[6776] = '{5};
test_input[54216:54223] = '{32'h4246d853, 32'hc2aec01a, 32'hc1fde17a, 32'hc213b3aa, 32'hc278b76d, 32'h41a98a99, 32'hc0ce0af9, 32'h42104d6c};
test_output[6777] = '{32'h4246d853};
test_index[6777] = '{0};
test_input[54224:54231] = '{32'hc1d0d565, 32'h422caecb, 32'h42862c43, 32'h427e914a, 32'hc288b5df, 32'h429453a7, 32'h42978149, 32'h40cddeed};
test_output[6778] = '{32'h42978149};
test_index[6778] = '{6};
test_input[54232:54239] = '{32'hc2b136e6, 32'hc1d0614a, 32'hc21ad228, 32'hc1616158, 32'h4216b8f7, 32'h42143fcb, 32'h422fde70, 32'hc28421ca};
test_output[6779] = '{32'h422fde70};
test_index[6779] = '{6};
test_input[54240:54247] = '{32'hc2792212, 32'h41d120fe, 32'hc2c2a7fc, 32'h41fa89e7, 32'h4296e2fa, 32'h4054643f, 32'h419908aa, 32'hc21abfb8};
test_output[6780] = '{32'h4296e2fa};
test_index[6780] = '{4};
test_input[54248:54255] = '{32'hc2598385, 32'h426c6e24, 32'hc291d337, 32'h4282e15d, 32'hc2925e5a, 32'h4272c4e1, 32'hc1646ea6, 32'hc02b9d98};
test_output[6781] = '{32'h4282e15d};
test_index[6781] = '{3};
test_input[54256:54263] = '{32'h4199aec7, 32'hc2938c8f, 32'hc2c18087, 32'h4296a6f2, 32'hc1a5aae1, 32'hc1a39873, 32'h420e6e1a, 32'h42b11ec8};
test_output[6782] = '{32'h42b11ec8};
test_index[6782] = '{7};
test_input[54264:54271] = '{32'h4153b0af, 32'h42013445, 32'h417a9fdd, 32'hc24a9811, 32'h3e98178b, 32'h422d41de, 32'hc2aad903, 32'hc2a976d4};
test_output[6783] = '{32'h422d41de};
test_index[6783] = '{5};
test_input[54272:54279] = '{32'hc1aff018, 32'hc26ae636, 32'h42933929, 32'h42976695, 32'h42519515, 32'h4239a6dc, 32'h429dcdf0, 32'hc24e8e1c};
test_output[6784] = '{32'h429dcdf0};
test_index[6784] = '{6};
test_input[54280:54287] = '{32'h41efe5cc, 32'hc26b584c, 32'h419b8443, 32'h42467e66, 32'h42491a9e, 32'h4077eeb9, 32'hc206b6e1, 32'hc26006f7};
test_output[6785] = '{32'h42491a9e};
test_index[6785] = '{4};
test_input[54288:54295] = '{32'hc27a1d32, 32'hc22bf5d5, 32'hc29c9052, 32'hc2627b4d, 32'hc268ced3, 32'h4252eb60, 32'h420a31cd, 32'hc2a992f9};
test_output[6786] = '{32'h4252eb60};
test_index[6786] = '{5};
test_input[54296:54303] = '{32'h42c4e321, 32'hc29443f3, 32'h41db5ec1, 32'hc2c1297e, 32'h42a8251f, 32'hc2be9219, 32'h42943a5a, 32'h42032302};
test_output[6787] = '{32'h42c4e321};
test_index[6787] = '{0};
test_input[54304:54311] = '{32'h41f06686, 32'h4249b424, 32'hc274de2e, 32'h418001da, 32'h427c7f8f, 32'h40c76e99, 32'h425ea304, 32'hc259252d};
test_output[6788] = '{32'h427c7f8f};
test_index[6788] = '{4};
test_input[54312:54319] = '{32'hc1bf5873, 32'hc2c1ea21, 32'hc2bf306d, 32'h42b3173a, 32'hc26f590a, 32'h42c4e2d7, 32'hc2928747, 32'hc181a582};
test_output[6789] = '{32'h42c4e2d7};
test_index[6789] = '{5};
test_input[54320:54327] = '{32'hc1597c73, 32'h4077ff37, 32'h42266ee0, 32'hc10c05a2, 32'hc21484b4, 32'hc24b2e67, 32'h426d7579, 32'hc286f432};
test_output[6790] = '{32'h426d7579};
test_index[6790] = '{6};
test_input[54328:54335] = '{32'hc1ba122f, 32'hc0cfd5b0, 32'h40ce6b49, 32'hc2b9903b, 32'h420da918, 32'hc262da59, 32'hc2163717, 32'h4227a32a};
test_output[6791] = '{32'h4227a32a};
test_index[6791] = '{7};
test_input[54336:54343] = '{32'hbff36b6b, 32'h41d3fb0b, 32'h42a5155f, 32'hc243e8a1, 32'h4155db47, 32'h42296b2a, 32'h42290a82, 32'hc2b50076};
test_output[6792] = '{32'h42a5155f};
test_index[6792] = '{2};
test_input[54344:54351] = '{32'hc1d3694c, 32'hc20e7982, 32'hc2c1d398, 32'hc199c9a3, 32'hc29ee697, 32'hc29c7d3a, 32'hc2bd2312, 32'hc2a74e3a};
test_output[6793] = '{32'hc199c9a3};
test_index[6793] = '{3};
test_input[54352:54359] = '{32'hc2b7fec6, 32'hc2a6a134, 32'hc296d287, 32'h4283e5ff, 32'hc2bf982e, 32'hc1b76a04, 32'hc292c3b6, 32'h42ab5f8e};
test_output[6794] = '{32'h42ab5f8e};
test_index[6794] = '{7};
test_input[54360:54367] = '{32'h4036e496, 32'hc1e84023, 32'hc22e09c8, 32'hbead4657, 32'hc18ef525, 32'hc2b31985, 32'h427bb7e8, 32'hc25c6375};
test_output[6795] = '{32'h427bb7e8};
test_index[6795] = '{6};
test_input[54368:54375] = '{32'hc2b6800c, 32'h3e6eba05, 32'hc2bbf6b6, 32'hc25e1d4b, 32'hc2c7fc1c, 32'h421e4ba6, 32'hc202bd21, 32'hc0f85d9d};
test_output[6796] = '{32'h421e4ba6};
test_index[6796] = '{5};
test_input[54376:54383] = '{32'hc2a16e77, 32'hc1db6a86, 32'h40b42799, 32'h42a0d3ee, 32'h4280e07e, 32'h40ecf1e4, 32'hc2323297, 32'hc28cc511};
test_output[6797] = '{32'h42a0d3ee};
test_index[6797] = '{3};
test_input[54384:54391] = '{32'hc253e321, 32'hc20f640b, 32'hc2127597, 32'hc1bbcb4a, 32'h424454d1, 32'hc2a26f2e, 32'hc2bde9cf, 32'hc1d6f699};
test_output[6798] = '{32'h424454d1};
test_index[6798] = '{4};
test_input[54392:54399] = '{32'h42577959, 32'hc22e2122, 32'h429b3663, 32'hc2698023, 32'h42b75034, 32'hc283414a, 32'h4147dbca, 32'hc28149bd};
test_output[6799] = '{32'h42b75034};
test_index[6799] = '{4};
test_input[54400:54407] = '{32'h41b71b38, 32'h41152a77, 32'hc2440294, 32'h41130f4a, 32'hc18172bf, 32'h420b1fb0, 32'h42933640, 32'h42920235};
test_output[6800] = '{32'h42933640};
test_index[6800] = '{6};
test_input[54408:54415] = '{32'hc010b97e, 32'h41d64489, 32'h41f5ccf1, 32'hc27884b9, 32'hc282ac7c, 32'h42441114, 32'h4213dca3, 32'h421d170d};
test_output[6801] = '{32'h42441114};
test_index[6801] = '{5};
test_input[54416:54423] = '{32'hc2055132, 32'h3e5e570d, 32'h42a2db3b, 32'hc2780856, 32'h3fcfddee, 32'h429b1de2, 32'h421e152f, 32'hc1ab0d12};
test_output[6802] = '{32'h42a2db3b};
test_index[6802] = '{2};
test_input[54424:54431] = '{32'h4297388c, 32'h41dbaeca, 32'hc20aa0b5, 32'h420b6305, 32'hc2ab60b9, 32'hc2800bb6, 32'hc19a4832, 32'h42bf7c87};
test_output[6803] = '{32'h42bf7c87};
test_index[6803] = '{7};
test_input[54432:54439] = '{32'h41b27483, 32'h4121c369, 32'h42935992, 32'h40a423c3, 32'h41a92916, 32'h42406b63, 32'h42792ce0, 32'hc29fe167};
test_output[6804] = '{32'h42935992};
test_index[6804] = '{2};
test_input[54440:54447] = '{32'h4273f586, 32'hc2c1c197, 32'hc2610ab6, 32'hc18aea5b, 32'hc28b6cb1, 32'hc161668a, 32'hc23bd573, 32'h428b6520};
test_output[6805] = '{32'h428b6520};
test_index[6805] = '{7};
test_input[54448:54455] = '{32'h3ff36b3e, 32'h4077463d, 32'hc17f4c04, 32'h42825401, 32'hc28f6a34, 32'hc173f7f1, 32'h42ba8430, 32'hc26f2f07};
test_output[6806] = '{32'h42ba8430};
test_index[6806] = '{6};
test_input[54456:54463] = '{32'h428dabc4, 32'hc214b735, 32'hc005a036, 32'h42bf4f46, 32'h3e48da1f, 32'h4286c1a0, 32'h424b3134, 32'h4296cf96};
test_output[6807] = '{32'h42bf4f46};
test_index[6807] = '{3};
test_input[54464:54471] = '{32'hc2272b7c, 32'hbad6ac2d, 32'h4275c0e6, 32'hc0304140, 32'hc2b990dc, 32'hc0538e7e, 32'h41c84af7, 32'hc2a0d9de};
test_output[6808] = '{32'h4275c0e6};
test_index[6808] = '{2};
test_input[54472:54479] = '{32'hc2035cb1, 32'hc22fd8d4, 32'hc2af41a6, 32'hc28fcbba, 32'h3fd40dfd, 32'h41c18220, 32'hc26a89f5, 32'h41bde07a};
test_output[6809] = '{32'h41c18220};
test_index[6809] = '{5};
test_input[54480:54487] = '{32'h411cef54, 32'hc2b33dfa, 32'hc2aebd0b, 32'hc10dfa74, 32'hc253eb43, 32'hc18b402b, 32'hc267eb77, 32'hc2ad5cad};
test_output[6810] = '{32'h411cef54};
test_index[6810] = '{0};
test_input[54488:54495] = '{32'hbf959030, 32'h425d97b9, 32'h42b5cc41, 32'h3ffa1ab0, 32'hc2be8d1c, 32'h4257278d, 32'hc2ada75b, 32'hc26a5182};
test_output[6811] = '{32'h42b5cc41};
test_index[6811] = '{2};
test_input[54496:54503] = '{32'hc26faf43, 32'hc237be54, 32'hc291f4d1, 32'hc29003fa, 32'h42958893, 32'hc29c881f, 32'hc2a68712, 32'h412a0f8f};
test_output[6812] = '{32'h42958893};
test_index[6812] = '{4};
test_input[54504:54511] = '{32'h41c9ed4c, 32'hc2853dbf, 32'hc204899b, 32'hc2b9aa72, 32'h41e555af, 32'hc22f5a79, 32'hc19e3d30, 32'h419863df};
test_output[6813] = '{32'h41e555af};
test_index[6813] = '{4};
test_input[54512:54519] = '{32'h42ba0481, 32'hc2c67349, 32'h42c5a282, 32'hc2804ce0, 32'h42a7575e, 32'h41d99cdd, 32'hc184937b, 32'h427cddf7};
test_output[6814] = '{32'h42c5a282};
test_index[6814] = '{2};
test_input[54520:54527] = '{32'hc2417e3d, 32'h42b5400e, 32'hc2a1257a, 32'hc2bab779, 32'hc2827b27, 32'hc293eac5, 32'hc27c1fb5, 32'h4052ce99};
test_output[6815] = '{32'h42b5400e};
test_index[6815] = '{1};
test_input[54528:54535] = '{32'hc14968b2, 32'hc12998e6, 32'hc0d3d0f1, 32'hc248f7f4, 32'h42700126, 32'h425531c5, 32'hc276c9ca, 32'h428d8211};
test_output[6816] = '{32'h428d8211};
test_index[6816] = '{7};
test_input[54536:54543] = '{32'hc26fac51, 32'h41401c95, 32'h42aa5b86, 32'hc1b66a9d, 32'h42b2d0f9, 32'hc0e5364f, 32'hc25385a5, 32'h4210d045};
test_output[6817] = '{32'h42b2d0f9};
test_index[6817] = '{4};
test_input[54544:54551] = '{32'h41aec75a, 32'hc28636c4, 32'hc2aae360, 32'h4284edeb, 32'hc186a51e, 32'h4296ea90, 32'h42ba46a6, 32'hc20fbd94};
test_output[6818] = '{32'h42ba46a6};
test_index[6818] = '{6};
test_input[54552:54559] = '{32'h42149a50, 32'h421c1741, 32'hc1fe811e, 32'h41858003, 32'h42882aaa, 32'h422b8efa, 32'hc247e275, 32'h423660e1};
test_output[6819] = '{32'h42882aaa};
test_index[6819] = '{4};
test_input[54560:54567] = '{32'h42592621, 32'h42aeabac, 32'hc23d8949, 32'hc220bed0, 32'hc2892a8f, 32'h41fb635a, 32'h423afd00, 32'hc277fb7b};
test_output[6820] = '{32'h42aeabac};
test_index[6820] = '{1};
test_input[54568:54575] = '{32'hc23a3f1a, 32'h42049b67, 32'h41dc48cf, 32'hc1c156d0, 32'h42ba5b73, 32'h424d01f9, 32'hc26781eb, 32'hc2a4e851};
test_output[6821] = '{32'h42ba5b73};
test_index[6821] = '{4};
test_input[54576:54583] = '{32'hc267c48b, 32'h42760167, 32'h429038e0, 32'h41a79358, 32'hc282b0fa, 32'h427a8a1d, 32'h4281f58b, 32'hc1d5c2d7};
test_output[6822] = '{32'h429038e0};
test_index[6822] = '{2};
test_input[54584:54591] = '{32'h422fd97c, 32'hc1a9b2e9, 32'h42573a29, 32'h4249f46b, 32'hc27a0a9f, 32'hc0b62b8d, 32'h42c39be7, 32'hc25027ed};
test_output[6823] = '{32'h42c39be7};
test_index[6823] = '{6};
test_input[54592:54599] = '{32'h428092d8, 32'hc29fb841, 32'h40475e4d, 32'h42081f26, 32'hc171849b, 32'hc1e2bc8b, 32'h42769109, 32'hc2996fef};
test_output[6824] = '{32'h428092d8};
test_index[6824] = '{0};
test_input[54600:54607] = '{32'hc24e3e41, 32'hc269f553, 32'h41e74c40, 32'hc2a4286c, 32'hc2b18bc3, 32'hc18d8d47, 32'hc2c537cd, 32'h427f7cb5};
test_output[6825] = '{32'h427f7cb5};
test_index[6825] = '{7};
test_input[54608:54615] = '{32'h427452d4, 32'hc2c61436, 32'h424e2f63, 32'hc21fac3e, 32'hc20038bd, 32'h413e7a31, 32'h42909299, 32'h42018630};
test_output[6826] = '{32'h42909299};
test_index[6826] = '{6};
test_input[54616:54623] = '{32'h42a7cffb, 32'hc207ede6, 32'hc1cea7b8, 32'h426a29c0, 32'hc2549d0d, 32'hc28af1a4, 32'h419e8f1a, 32'hc192d421};
test_output[6827] = '{32'h42a7cffb};
test_index[6827] = '{0};
test_input[54624:54631] = '{32'h42941a7f, 32'h40584e22, 32'h41f612c7, 32'hc11358cf, 32'h427b84a5, 32'hc1ddad8d, 32'hc16d67aa, 32'hc28e634d};
test_output[6828] = '{32'h42941a7f};
test_index[6828] = '{0};
test_input[54632:54639] = '{32'h42415b31, 32'hc1118488, 32'h4284e5e6, 32'hc291afe5, 32'hc25360b4, 32'h42b1b614, 32'hc2050e11, 32'hc2bc1b10};
test_output[6829] = '{32'h42b1b614};
test_index[6829] = '{5};
test_input[54640:54647] = '{32'hc19bead8, 32'hc170e5dc, 32'hc27fdff6, 32'hc2a402aa, 32'hc23e0c33, 32'h42b31f73, 32'hc2099097, 32'hc2910b93};
test_output[6830] = '{32'h42b31f73};
test_index[6830] = '{5};
test_input[54648:54655] = '{32'h41ce2529, 32'h42a3e0bf, 32'hbdd41bf3, 32'hc2953b3f, 32'h42af8d86, 32'h4227d303, 32'hc29d401c, 32'h42247e4e};
test_output[6831] = '{32'h42af8d86};
test_index[6831] = '{4};
test_input[54656:54663] = '{32'h40527b6f, 32'hc22a07f2, 32'hc2b33f1a, 32'hc18b9bbc, 32'hc215b7a1, 32'h42bd3c3b, 32'hc2c0573e, 32'h428c2403};
test_output[6832] = '{32'h42bd3c3b};
test_index[6832] = '{5};
test_input[54664:54671] = '{32'hc1a108ef, 32'h41a35c6c, 32'hc2987698, 32'hc295c0c0, 32'hc2a9ffd6, 32'h42b9e745, 32'h3f566420, 32'hc2ac4f20};
test_output[6833] = '{32'h42b9e745};
test_index[6833] = '{5};
test_input[54672:54679] = '{32'hc21208a4, 32'h428b9375, 32'h42c6788e, 32'hc26fe343, 32'h42bf8f9e, 32'hc2b72d76, 32'h3fd15681, 32'h4293f418};
test_output[6834] = '{32'h42c6788e};
test_index[6834] = '{2};
test_input[54680:54687] = '{32'hc218d05e, 32'h429f7133, 32'hbf5f6150, 32'h42822cde, 32'hc1bea5fb, 32'h42c2684e, 32'h41f03e2b, 32'hc29b0e99};
test_output[6835] = '{32'h42c2684e};
test_index[6835] = '{5};
test_input[54688:54695] = '{32'h40a4d8eb, 32'h4298a2dd, 32'h41310903, 32'h41e62c8b, 32'hc10d26a4, 32'hc258ebca, 32'hc26541d3, 32'hc0f8535f};
test_output[6836] = '{32'h4298a2dd};
test_index[6836] = '{1};
test_input[54696:54703] = '{32'hc2777472, 32'hc2b370a9, 32'hc20ad979, 32'h428d5d89, 32'hc181b1ec, 32'hc2bac8d4, 32'h428dbd4a, 32'hc2bca7ab};
test_output[6837] = '{32'h428dbd4a};
test_index[6837] = '{6};
test_input[54704:54711] = '{32'h423ed89b, 32'h41b5208b, 32'hc28fff44, 32'h42271a21, 32'h420b22cd, 32'hc258cb12, 32'h424f5e99, 32'h42aa876c};
test_output[6838] = '{32'h42aa876c};
test_index[6838] = '{7};
test_input[54712:54719] = '{32'hc228e57b, 32'hc20aeff3, 32'h409de825, 32'h42a3434a, 32'hc0dc509d, 32'hc0460dba, 32'hc1cb07c4, 32'hc2bf5d0c};
test_output[6839] = '{32'h42a3434a};
test_index[6839] = '{3};
test_input[54720:54727] = '{32'hc2b704aa, 32'hc217e3f0, 32'h42abb09b, 32'h4288bd10, 32'hc2a0fd3e, 32'hc11e2f72, 32'h401c9d22, 32'hc26113ac};
test_output[6840] = '{32'h42abb09b};
test_index[6840] = '{2};
test_input[54728:54735] = '{32'hc2902e4d, 32'h429e8c23, 32'h42055e90, 32'h42c5b32b, 32'hbf70650f, 32'hc20ee8a5, 32'h423c436a, 32'hc29fe160};
test_output[6841] = '{32'h42c5b32b};
test_index[6841] = '{3};
test_input[54736:54743] = '{32'hc102f9af, 32'h41e125a8, 32'h401c5d88, 32'hc2a01fd1, 32'hc28619cd, 32'hc27c73e2, 32'hc1e8a803, 32'hc2c6a72f};
test_output[6842] = '{32'h41e125a8};
test_index[6842] = '{1};
test_input[54744:54751] = '{32'hc157da52, 32'h422b45f1, 32'h41fb5cb5, 32'hc27aaa97, 32'hc19e7e84, 32'hc14ff41a, 32'hc298a552, 32'hc130e3eb};
test_output[6843] = '{32'h422b45f1};
test_index[6843] = '{1};
test_input[54752:54759] = '{32'hc05df02f, 32'hc05008d6, 32'h42b825ba, 32'h42ba7441, 32'hc2ac7846, 32'h41f2d2c3, 32'hc2a46720, 32'h423da9de};
test_output[6844] = '{32'h42ba7441};
test_index[6844] = '{3};
test_input[54760:54767] = '{32'hc232aeac, 32'hc28a5c2b, 32'h42c55f7c, 32'h40e78da9, 32'hc2065bb8, 32'h428f4918, 32'h426cfa85, 32'hc239f849};
test_output[6845] = '{32'h42c55f7c};
test_index[6845] = '{2};
test_input[54768:54775] = '{32'h423cba73, 32'hc2b8e996, 32'h42714ce7, 32'h429a9939, 32'hc1a49ec1, 32'h422c7a81, 32'h41d886df, 32'h41e8775e};
test_output[6846] = '{32'h429a9939};
test_index[6846] = '{3};
test_input[54776:54783] = '{32'hc234e523, 32'h42316d69, 32'h42392c07, 32'hc20234df, 32'h42123c50, 32'hc13c34b8, 32'hc0ac7ff6, 32'h42660adc};
test_output[6847] = '{32'h42660adc};
test_index[6847] = '{7};
test_input[54784:54791] = '{32'h424f86b9, 32'h4266a5a8, 32'hc2bfec34, 32'h4279bc0c, 32'hc253125c, 32'hc2816ae6, 32'hc25ce663, 32'h4177189d};
test_output[6848] = '{32'h4279bc0c};
test_index[6848] = '{3};
test_input[54792:54799] = '{32'hc24a085e, 32'hc25dbcc9, 32'h4272bfc5, 32'h428f5a83, 32'h4297ec33, 32'hc02136e3, 32'h426b445f, 32'hc2b365ae};
test_output[6849] = '{32'h4297ec33};
test_index[6849] = '{4};
test_input[54800:54807] = '{32'h4236b45a, 32'hc2a6350b, 32'hc278c92a, 32'h4252dfec, 32'h42c4d433, 32'h41aa9e46, 32'hc1f2122d, 32'hc28f0cc2};
test_output[6850] = '{32'h42c4d433};
test_index[6850] = '{4};
test_input[54808:54815] = '{32'hc2afcd98, 32'hc1b8cc77, 32'hc2aafe27, 32'h41d0d2bf, 32'h429c9fb3, 32'hc0e5c6db, 32'h4139d3d7, 32'hc2679f8d};
test_output[6851] = '{32'h429c9fb3};
test_index[6851] = '{4};
test_input[54816:54823] = '{32'h41bc5cdb, 32'h415310c9, 32'hc1cb3c15, 32'hc2b459da, 32'h409604d0, 32'h426314eb, 32'hc2119166, 32'hc1816570};
test_output[6852] = '{32'h426314eb};
test_index[6852] = '{5};
test_input[54824:54831] = '{32'hc221a079, 32'h41a08e21, 32'h4265b428, 32'hc2739431, 32'hc294bf48, 32'hc1fa97cc, 32'h41007cda, 32'h42a05217};
test_output[6853] = '{32'h42a05217};
test_index[6853] = '{7};
test_input[54832:54839] = '{32'h428bc727, 32'hc2619146, 32'h42b7b756, 32'h4179cc54, 32'h423846e5, 32'hc27339ab, 32'h42aa933b, 32'hc13b56a3};
test_output[6854] = '{32'h42b7b756};
test_index[6854] = '{2};
test_input[54840:54847] = '{32'hc181b890, 32'h41fd53c3, 32'hc29af410, 32'h42344da0, 32'h405d4b55, 32'hc17d65c4, 32'h42733be5, 32'h42b22072};
test_output[6855] = '{32'h42b22072};
test_index[6855] = '{7};
test_input[54848:54855] = '{32'hc2c5c8e8, 32'h419c1ee4, 32'hc2884553, 32'h42693137, 32'h40e521bf, 32'h41e147f6, 32'h428293f5, 32'hc17651a6};
test_output[6856] = '{32'h428293f5};
test_index[6856] = '{6};
test_input[54856:54863] = '{32'h42935470, 32'h4127ba51, 32'hc22284ca, 32'hc262387a, 32'hc0e72818, 32'hc1853f2c, 32'h42560136, 32'hc2774806};
test_output[6857] = '{32'h42935470};
test_index[6857] = '{0};
test_input[54864:54871] = '{32'h418e69fd, 32'hc25ead23, 32'hc2a6b975, 32'hc1557f43, 32'h419a7053, 32'h41dd6b7b, 32'hc289d5b5, 32'h428686f1};
test_output[6858] = '{32'h428686f1};
test_index[6858] = '{7};
test_input[54872:54879] = '{32'hc2020b16, 32'h41c84335, 32'hc2af0233, 32'hc14d1143, 32'hc1497572, 32'h41d73f9e, 32'h4250ba96, 32'h41456c70};
test_output[6859] = '{32'h4250ba96};
test_index[6859] = '{6};
test_input[54880:54887] = '{32'hc2481aca, 32'h42b0d019, 32'h426d32a1, 32'h41ddef5c, 32'hc18f9288, 32'h42568a28, 32'hc2b03328, 32'h42a9c694};
test_output[6860] = '{32'h42b0d019};
test_index[6860] = '{1};
test_input[54888:54895] = '{32'h409ead11, 32'hc1f3ed02, 32'hc2bb75b0, 32'hc2be41ac, 32'h428663b2, 32'hc1df652c, 32'hc1b138a9, 32'hc278bc9a};
test_output[6861] = '{32'h428663b2};
test_index[6861] = '{4};
test_input[54896:54903] = '{32'hc0ec9824, 32'hc152502b, 32'hc2134072, 32'hc20dc109, 32'h4299793b, 32'hc08cf904, 32'hc1eab1d0, 32'h4117e1f0};
test_output[6862] = '{32'h4299793b};
test_index[6862] = '{4};
test_input[54904:54911] = '{32'hc06746a0, 32'hc22bd4a2, 32'h42a5a89f, 32'hc2107259, 32'h4173df60, 32'h41816e2d, 32'hc2ad0d4a, 32'hc2c2516e};
test_output[6863] = '{32'h42a5a89f};
test_index[6863] = '{2};
test_input[54912:54919] = '{32'hc2bad4c6, 32'hc2abb179, 32'hc27c25cb, 32'hc2b5ba69, 32'h4221dc26, 32'h4281c086, 32'hc2462054, 32'hc2221f5b};
test_output[6864] = '{32'h4281c086};
test_index[6864] = '{5};
test_input[54920:54927] = '{32'hc28ce265, 32'h4291542b, 32'h42bbf87f, 32'hc28052a8, 32'hc1a1bd4e, 32'h418888d2, 32'h427c5733, 32'h42bdba9b};
test_output[6865] = '{32'h42bdba9b};
test_index[6865] = '{7};
test_input[54928:54935] = '{32'hc279e241, 32'hc290603e, 32'h42a2e2ce, 32'hc2b9d365, 32'h427f21cf, 32'h427cadac, 32'h427c72ab, 32'h42af1529};
test_output[6866] = '{32'h42af1529};
test_index[6866] = '{7};
test_input[54936:54943] = '{32'hc28f9a52, 32'h421bc4e6, 32'hc26595f8, 32'hc23ccf7e, 32'h422ff986, 32'hc24eba1f, 32'hc2467035, 32'h4271f774};
test_output[6867] = '{32'h4271f774};
test_index[6867] = '{7};
test_input[54944:54951] = '{32'hc2149c5d, 32'hc249fa4c, 32'h42974619, 32'hc2843dcf, 32'hbfd827fe, 32'h424dae45, 32'hc1dceed6, 32'h425dc666};
test_output[6868] = '{32'h42974619};
test_index[6868] = '{2};
test_input[54952:54959] = '{32'h42a65e5e, 32'h42715110, 32'h42bd4200, 32'h42088b41, 32'h3d17f250, 32'h42761f5a, 32'hc2be90eb, 32'hc2bf53c9};
test_output[6869] = '{32'h42bd4200};
test_index[6869] = '{2};
test_input[54960:54967] = '{32'h4286e718, 32'hc1d841b2, 32'h40d7f7c4, 32'h40a60df6, 32'h42bf6ee6, 32'h4233b90c, 32'hc297466e, 32'hc2ba0a84};
test_output[6870] = '{32'h42bf6ee6};
test_index[6870] = '{4};
test_input[54968:54975] = '{32'hc29c5510, 32'hc23b8816, 32'hc23964ac, 32'hc2906f68, 32'hc22c0bfc, 32'h42901ce5, 32'h4111bf79, 32'hc288ca57};
test_output[6871] = '{32'h42901ce5};
test_index[6871] = '{5};
test_input[54976:54983] = '{32'h42659601, 32'hc29d9806, 32'h42a5a228, 32'hc1b9f4da, 32'hc2af27bc, 32'h429bac46, 32'hc1ac79c6, 32'h4198893b};
test_output[6872] = '{32'h42a5a228};
test_index[6872] = '{2};
test_input[54984:54991] = '{32'hc21650ae, 32'h41f30a37, 32'hc1d2cd27, 32'h4284753a, 32'hc2184b64, 32'h42bf8fb8, 32'hc1b1e24c, 32'hc296cb73};
test_output[6873] = '{32'h42bf8fb8};
test_index[6873] = '{5};
test_input[54992:54999] = '{32'h426155e7, 32'h4296df75, 32'hc2c60680, 32'h42221600, 32'h41b4eadf, 32'hc2a09b6f, 32'hc206354d, 32'h41901df9};
test_output[6874] = '{32'h4296df75};
test_index[6874] = '{1};
test_input[55000:55007] = '{32'h420eb02e, 32'h424453b2, 32'h418279fe, 32'h416d2db6, 32'h40a79ab6, 32'h428be55d, 32'hc0bbacd0, 32'h41ec49cf};
test_output[6875] = '{32'h428be55d};
test_index[6875] = '{5};
test_input[55008:55015] = '{32'hc2beb290, 32'hc28bc600, 32'hc2c529be, 32'h4204816f, 32'h41989162, 32'h423d677d, 32'hc2004587, 32'hc2106692};
test_output[6876] = '{32'h423d677d};
test_index[6876] = '{5};
test_input[55016:55023] = '{32'h42be1d97, 32'h4235383a, 32'hc1eb200a, 32'h421bb83d, 32'hc281f7d0, 32'hc2abb6b7, 32'h42a96e04, 32'hc27177f0};
test_output[6877] = '{32'h42be1d97};
test_index[6877] = '{0};
test_input[55024:55031] = '{32'hc26ecc40, 32'hc2a7049c, 32'hc156043c, 32'hc2a183d7, 32'hc2ad3f6a, 32'h42a3fa4b, 32'h416cd10f, 32'hc2918ff8};
test_output[6878] = '{32'h42a3fa4b};
test_index[6878] = '{5};
test_input[55032:55039] = '{32'hc2ac1039, 32'h427866e5, 32'hc2c1d918, 32'h40db633c, 32'h42931ec0, 32'hc1aad994, 32'h42894a32, 32'hc292e7ed};
test_output[6879] = '{32'h42931ec0};
test_index[6879] = '{4};
test_input[55040:55047] = '{32'hc075bdc8, 32'h425fa96e, 32'h42a90928, 32'hc2ab2552, 32'h42a24d50, 32'h428fc378, 32'h4007e65f, 32'h41e3e934};
test_output[6880] = '{32'h42a90928};
test_index[6880] = '{2};
test_input[55048:55055] = '{32'hc1ca98bb, 32'hc29fcca0, 32'hc2a03470, 32'hc249804e, 32'h41e1aea8, 32'h42168162, 32'hc29c64ea, 32'h42b8420a};
test_output[6881] = '{32'h42b8420a};
test_index[6881] = '{7};
test_input[55056:55063] = '{32'hc1949871, 32'hc29690b7, 32'hbfd46f14, 32'h41aaff8c, 32'h42204588, 32'h424b5d27, 32'hc18e15c8, 32'h4294fc28};
test_output[6882] = '{32'h4294fc28};
test_index[6882] = '{7};
test_input[55064:55071] = '{32'h42714023, 32'h42c01c4e, 32'h42183fa9, 32'hc1d9f7bb, 32'h412bc671, 32'hc2a52924, 32'hc1a7a187, 32'hc27c00d9};
test_output[6883] = '{32'h42c01c4e};
test_index[6883] = '{1};
test_input[55072:55079] = '{32'hc1878928, 32'hc277b555, 32'h424b4f50, 32'h42968850, 32'hc28685ef, 32'h4239265e, 32'h41c2c1fb, 32'hc141d2ec};
test_output[6884] = '{32'h42968850};
test_index[6884] = '{3};
test_input[55080:55087] = '{32'hc2a729c5, 32'hc1ec0c62, 32'h42bc0666, 32'hc20478b2, 32'hc2183e68, 32'hc24cc696, 32'h41defb81, 32'hc23b029a};
test_output[6885] = '{32'h42bc0666};
test_index[6885] = '{2};
test_input[55088:55095] = '{32'h423a2e07, 32'hc2a3bed1, 32'h4188d0ec, 32'h4230ddc0, 32'hc2a83e5e, 32'h42c16ef1, 32'h4201b556, 32'hc2847d1f};
test_output[6886] = '{32'h42c16ef1};
test_index[6886] = '{5};
test_input[55096:55103] = '{32'hc291cf36, 32'h4275f333, 32'hc24725e6, 32'h40e666fe, 32'h4290ae5a, 32'hc145579d, 32'hc26f0064, 32'hc2944c42};
test_output[6887] = '{32'h4290ae5a};
test_index[6887] = '{4};
test_input[55104:55111] = '{32'h4197cb5e, 32'hc06ec16b, 32'hc2465091, 32'h419baad1, 32'hc20b22fb, 32'hc21df198, 32'h42be5980, 32'h4298c798};
test_output[6888] = '{32'h42be5980};
test_index[6888] = '{6};
test_input[55112:55119] = '{32'hc269e925, 32'h40f41cd8, 32'h4211de4e, 32'hc2719558, 32'hc13cc3cd, 32'h41af3a52, 32'hc25a85c7, 32'h414097ee};
test_output[6889] = '{32'h4211de4e};
test_index[6889] = '{2};
test_input[55120:55127] = '{32'h42b5d0ce, 32'h429cd53d, 32'hc25d017d, 32'h42ae274d, 32'h42713587, 32'hc28a7379, 32'hc25ffc20, 32'h41dfd248};
test_output[6890] = '{32'h42b5d0ce};
test_index[6890] = '{0};
test_input[55128:55135] = '{32'h4269af57, 32'hc20ffe4f, 32'h4289f5dd, 32'hc0d4c16c, 32'h422f28a2, 32'h4222398f, 32'hc27acd71, 32'hc28fd1be};
test_output[6891] = '{32'h4289f5dd};
test_index[6891] = '{2};
test_input[55136:55143] = '{32'h42323232, 32'h4233a920, 32'hbfd2fb8a, 32'h3e0edead, 32'h42413ae5, 32'hc1b7ae0c, 32'hc2827e83, 32'hc2a0f7f6};
test_output[6892] = '{32'h42413ae5};
test_index[6892] = '{4};
test_input[55144:55151] = '{32'hc2ba4deb, 32'hc0d2a92e, 32'hc1c99000, 32'h42c495e2, 32'h424b34f0, 32'hc250b376, 32'hc18b303c, 32'h421122d6};
test_output[6893] = '{32'h42c495e2};
test_index[6893] = '{3};
test_input[55152:55159] = '{32'h405554f8, 32'hc1fb8e1b, 32'h4274d03c, 32'hc23c1b63, 32'hc1ae6979, 32'hc19fc088, 32'hc23e96bc, 32'h42bfd959};
test_output[6894] = '{32'h42bfd959};
test_index[6894] = '{7};
test_input[55160:55167] = '{32'hc1c88f88, 32'h41f9ef1e, 32'h42a32362, 32'hc1339c0e, 32'h428ee4ba, 32'h42b2b2b2, 32'h41d40cc6, 32'h424bd1ed};
test_output[6895] = '{32'h42b2b2b2};
test_index[6895] = '{5};
test_input[55168:55175] = '{32'h41cb10e2, 32'hc2aa21b9, 32'hc26d9823, 32'hc20692e7, 32'hc2323523, 32'h428fdffd, 32'h424f1d74, 32'hc285f0a0};
test_output[6896] = '{32'h428fdffd};
test_index[6896] = '{5};
test_input[55176:55183] = '{32'hc239841f, 32'h421fb6c8, 32'h42226c86, 32'h42b19be1, 32'hc2aa0302, 32'hc2887479, 32'h42bb67b9, 32'hc144b1b3};
test_output[6897] = '{32'h42bb67b9};
test_index[6897] = '{6};
test_input[55184:55191] = '{32'hc20e0833, 32'h427d400e, 32'h42bf31ee, 32'h425df88c, 32'hc27eb47e, 32'h4283b942, 32'h42ac12b9, 32'h4077ac63};
test_output[6898] = '{32'h42bf31ee};
test_index[6898] = '{2};
test_input[55192:55199] = '{32'hc1991ad5, 32'h4292d6a1, 32'hc29a2429, 32'hc1b3307b, 32'hc2a7dba5, 32'hc2b8b1aa, 32'hc126e4a7, 32'h42c4e485};
test_output[6899] = '{32'h42c4e485};
test_index[6899] = '{7};
test_input[55200:55207] = '{32'hc29a89e0, 32'hc2467954, 32'hc2bfb7c9, 32'h424425a9, 32'hc2b7c01b, 32'h42a04565, 32'hc1f080d5, 32'h41f65728};
test_output[6900] = '{32'h42a04565};
test_index[6900] = '{5};
test_input[55208:55215] = '{32'h4204decc, 32'hc15d0970, 32'h41b86f00, 32'h4208235f, 32'h4230303e, 32'h423a3970, 32'hc29150e7, 32'h4187bfbd};
test_output[6901] = '{32'h423a3970};
test_index[6901] = '{5};
test_input[55216:55223] = '{32'h41033b13, 32'hc2c68f44, 32'h42a57c68, 32'h42909bb7, 32'hc297f848, 32'h42012d94, 32'hc111944a, 32'hc2a319b2};
test_output[6902] = '{32'h42a57c68};
test_index[6902] = '{2};
test_input[55224:55231] = '{32'h40eb4b7b, 32'h408c5ff4, 32'h419a4c24, 32'hc1b4792e, 32'h423ae23d, 32'h41029fe3, 32'hc117db1f, 32'hc1de57ac};
test_output[6903] = '{32'h423ae23d};
test_index[6903] = '{4};
test_input[55232:55239] = '{32'hc2924c26, 32'h41368741, 32'hc1867d57, 32'h42048654, 32'h42822993, 32'h41b304ca, 32'h41940a50, 32'hc17bf599};
test_output[6904] = '{32'h42822993};
test_index[6904] = '{4};
test_input[55240:55247] = '{32'h4198dce0, 32'h41af5948, 32'h3f6890f4, 32'hc211a4e9, 32'h4186c653, 32'hc2a9d178, 32'h427df53c, 32'hc22c5dc3};
test_output[6905] = '{32'h427df53c};
test_index[6905] = '{6};
test_input[55248:55255] = '{32'h41101209, 32'h420a8a6b, 32'hc28ef692, 32'h427fc662, 32'h41d854af, 32'hc2162d09, 32'h40cfeb82, 32'hc2a22a36};
test_output[6906] = '{32'h427fc662};
test_index[6906] = '{3};
test_input[55256:55263] = '{32'h4249c34d, 32'hc27c29f8, 32'h4252b8ea, 32'hc0715886, 32'hc23e3cd8, 32'h426728e0, 32'hc298a476, 32'h416c18a4};
test_output[6907] = '{32'h426728e0};
test_index[6907] = '{5};
test_input[55264:55271] = '{32'hc2b2cf09, 32'hc00a8df7, 32'hc29d5ca1, 32'h41a3315a, 32'hc206a14c, 32'h40db2f7f, 32'hc113eb57, 32'h41932eeb};
test_output[6908] = '{32'h41a3315a};
test_index[6908] = '{3};
test_input[55272:55279] = '{32'h413c8a6f, 32'hc1e10664, 32'hc128149d, 32'hc10d1227, 32'h415d25a9, 32'hc22badac, 32'hc280c325, 32'hc2874dab};
test_output[6909] = '{32'h415d25a9};
test_index[6909] = '{4};
test_input[55280:55287] = '{32'h4251cead, 32'hc27aa7cd, 32'hc269b6f4, 32'hc2ab6a49, 32'h42b1c379, 32'hc065ed78, 32'hc265a584, 32'hc1d4f672};
test_output[6910] = '{32'h42b1c379};
test_index[6910] = '{4};
test_input[55288:55295] = '{32'h4100a02f, 32'h414f3a0a, 32'hc2994890, 32'h42433482, 32'hc2526ada, 32'hc2143ac5, 32'hc2880fd3, 32'hbea2894e};
test_output[6911] = '{32'h42433482};
test_index[6911] = '{3};
test_input[55296:55303] = '{32'hc2101693, 32'h41c8953a, 32'hc23e6026, 32'hc295d1fb, 32'hc21c9b7f, 32'hc2c4310c, 32'h41e1b408, 32'h414df92c};
test_output[6912] = '{32'h41e1b408};
test_index[6912] = '{6};
test_input[55304:55311] = '{32'hc0c67abf, 32'h421e5c2b, 32'h4219cd10, 32'hc15254ff, 32'h42984fc2, 32'hc21540f3, 32'h426cc885, 32'hc158bd9c};
test_output[6913] = '{32'h42984fc2};
test_index[6913] = '{4};
test_input[55312:55319] = '{32'hc28f6630, 32'hc2208e00, 32'hc1d9f33a, 32'h42710fe4, 32'h42b104b1, 32'hc1705aca, 32'hc15f1108, 32'hc129c78d};
test_output[6914] = '{32'h42b104b1};
test_index[6914] = '{4};
test_input[55320:55327] = '{32'hc24313a2, 32'h4113330f, 32'hc2afdaf8, 32'hc2b4cba2, 32'h42a52728, 32'hc1ea95ab, 32'hc2ad9706, 32'h42794592};
test_output[6915] = '{32'h42a52728};
test_index[6915] = '{4};
test_input[55328:55335] = '{32'h429f7d8d, 32'h42c333cf, 32'hc1927866, 32'h4266c536, 32'h4169c352, 32'h42530c63, 32'h42a567f3, 32'h428992c7};
test_output[6916] = '{32'h42c333cf};
test_index[6916] = '{1};
test_input[55336:55343] = '{32'hc0038ab4, 32'hc2151db2, 32'h409478de, 32'hc1f4726e, 32'hc1b13dba, 32'h41fd46d8, 32'h42bb7d65, 32'hc2c2706a};
test_output[6917] = '{32'h42bb7d65};
test_index[6917] = '{6};
test_input[55344:55351] = '{32'hc260198a, 32'hc285c9db, 32'hc101fc64, 32'h41d928b7, 32'h42a5fea4, 32'hc1212416, 32'hc1a13138, 32'h4235e9ec};
test_output[6918] = '{32'h42a5fea4};
test_index[6918] = '{4};
test_input[55352:55359] = '{32'hc23540d5, 32'hc209abb1, 32'hc13c2840, 32'hc1e2d2b4, 32'h40d70451, 32'hc2b674c0, 32'hc26a7a1b, 32'h426b0d23};
test_output[6919] = '{32'h426b0d23};
test_index[6919] = '{7};
test_input[55360:55367] = '{32'hc2b78c2e, 32'hc25fd72c, 32'hc24a4c5c, 32'h41eb2aee, 32'hc2aee59f, 32'h42a0dd07, 32'hc2c21d5d, 32'hc2191321};
test_output[6920] = '{32'h42a0dd07};
test_index[6920] = '{5};
test_input[55368:55375] = '{32'hc02b2020, 32'hbe3d2aff, 32'hc1b7f12e, 32'hc2930471, 32'hc2a568cb, 32'hc235fe98, 32'hc2b117f6, 32'h401fc6c0};
test_output[6921] = '{32'h401fc6c0};
test_index[6921] = '{7};
test_input[55376:55383] = '{32'hc274485f, 32'h42500b76, 32'h426d4dfc, 32'hc273bf12, 32'hc279b957, 32'hc281536e, 32'hc1d8e64a, 32'hc2a969c3};
test_output[6922] = '{32'h426d4dfc};
test_index[6922] = '{2};
test_input[55384:55391] = '{32'hc29d6e93, 32'h42b6b992, 32'hbf890ba7, 32'h42a34c43, 32'hc1e4d1f3, 32'h428ae78b, 32'h420977e4, 32'h4255298e};
test_output[6923] = '{32'h42b6b992};
test_index[6923] = '{1};
test_input[55392:55399] = '{32'h42650da2, 32'h41e12f45, 32'h42a8126d, 32'h4102d732, 32'h416118d3, 32'hc12d31bc, 32'h4289c6ef, 32'hc253edfd};
test_output[6924] = '{32'h42a8126d};
test_index[6924] = '{2};
test_input[55400:55407] = '{32'hbfc76e73, 32'h427f47e5, 32'h41d797a3, 32'hc2008c03, 32'hc200b9ba, 32'h4255c1c4, 32'hc1ce93a9, 32'hc2341b0b};
test_output[6925] = '{32'h427f47e5};
test_index[6925] = '{1};
test_input[55408:55415] = '{32'hc265b56e, 32'hc2430ee6, 32'h421f6eda, 32'hc0cf5a33, 32'hc2a8fe1e, 32'hc21e8c90, 32'hc2b41c1c, 32'h402c2504};
test_output[6926] = '{32'h421f6eda};
test_index[6926] = '{2};
test_input[55416:55423] = '{32'hc280a17d, 32'hc1e4dc6d, 32'hc0d5a0d5, 32'hc29652ab, 32'h42a7abb6, 32'hc13e5fd2, 32'h420e4360, 32'hc2863c9e};
test_output[6927] = '{32'h42a7abb6};
test_index[6927] = '{4};
test_input[55424:55431] = '{32'hc2b7f98f, 32'hc22841f1, 32'hc13b9d78, 32'h41785d4e, 32'hc22d08e8, 32'h422b89ed, 32'hc2b95c90, 32'hc1ba2625};
test_output[6928] = '{32'h422b89ed};
test_index[6928] = '{5};
test_input[55432:55439] = '{32'h3f7ac0e2, 32'h428f9b46, 32'h4240b4db, 32'h42ad9bf2, 32'h41456a4b, 32'hc1ba4321, 32'hc0c77b2b, 32'h41f4ef27};
test_output[6929] = '{32'h42ad9bf2};
test_index[6929] = '{3};
test_input[55440:55447] = '{32'hc2920787, 32'h42189736, 32'h41d05e42, 32'hc2c43937, 32'h41d17ecb, 32'h40392499, 32'h41fa8f5f, 32'h4219ecda};
test_output[6930] = '{32'h4219ecda};
test_index[6930] = '{7};
test_input[55448:55455] = '{32'h428736fc, 32'hc2884e6b, 32'h42c5307a, 32'hc1482ab7, 32'hc2962284, 32'hc240f4f5, 32'hc1dee3d5, 32'h42c7d7d8};
test_output[6931] = '{32'h42c7d7d8};
test_index[6931] = '{7};
test_input[55456:55463] = '{32'hc2356902, 32'h42a2e094, 32'hc29942cb, 32'hc1d33e54, 32'h41d1220c, 32'h4140c8a0, 32'h4240d23e, 32'h41f37ccc};
test_output[6932] = '{32'h42a2e094};
test_index[6932] = '{1};
test_input[55464:55471] = '{32'h429f7288, 32'h42a942cb, 32'h3e4554b1, 32'hc22a6db3, 32'hc288fdf7, 32'hc28447d0, 32'h42b3a6f7, 32'h42393ab8};
test_output[6933] = '{32'h42b3a6f7};
test_index[6933] = '{6};
test_input[55472:55479] = '{32'hc231c795, 32'hc28c4c65, 32'hc233e4c8, 32'h42a13f54, 32'hc29fb87a, 32'h42828387, 32'h41b5ac5e, 32'hc1becf55};
test_output[6934] = '{32'h42a13f54};
test_index[6934] = '{3};
test_input[55480:55487] = '{32'h428c0331, 32'hc14a5290, 32'hc29944dd, 32'h428ccaf8, 32'hc18e8073, 32'hc2a3f9c7, 32'h42064436, 32'hc22d58b3};
test_output[6935] = '{32'h428ccaf8};
test_index[6935] = '{3};
test_input[55488:55495] = '{32'hc1cf953e, 32'hc152bb23, 32'h42bd1e06, 32'hc2839e1d, 32'h41c740d5, 32'h41305a8e, 32'h41b9d2b2, 32'hc29f07c9};
test_output[6936] = '{32'h42bd1e06};
test_index[6936] = '{2};
test_input[55496:55503] = '{32'hc2c282f4, 32'hc2a6631b, 32'h42bddaf5, 32'hc177b5a6, 32'hc2c0a9dd, 32'hc25309dc, 32'hc0cc6f23, 32'hc2a30732};
test_output[6937] = '{32'h42bddaf5};
test_index[6937] = '{2};
test_input[55504:55511] = '{32'hc2804880, 32'h422d315a, 32'h4261fd57, 32'h42c397c1, 32'hc2ba4528, 32'h4183b631, 32'h42c52a1e, 32'h420467bf};
test_output[6938] = '{32'h42c52a1e};
test_index[6938] = '{6};
test_input[55512:55519] = '{32'h41b3124e, 32'h41a270e9, 32'h427c2ce3, 32'h41e7d623, 32'hc2a96d53, 32'hc238fcb8, 32'h428759ef, 32'hc22bec5f};
test_output[6939] = '{32'h428759ef};
test_index[6939] = '{6};
test_input[55520:55527] = '{32'h41680282, 32'h42add795, 32'hc232711d, 32'hc1cf971d, 32'hc2333c2e, 32'h41026b30, 32'h42bc7b86, 32'h42945ea2};
test_output[6940] = '{32'h42bc7b86};
test_index[6940] = '{6};
test_input[55528:55535] = '{32'hc268a2a6, 32'hc2120cd7, 32'hc12f3454, 32'h42a1e055, 32'hc28692df, 32'h42944482, 32'h42b71edb, 32'h41cc8dad};
test_output[6941] = '{32'h42b71edb};
test_index[6941] = '{6};
test_input[55536:55543] = '{32'hc2c57e89, 32'hc2c5fecd, 32'h42a794ba, 32'hc25c15fc, 32'h42b15f6d, 32'h40df246a, 32'hc26519ae, 32'hc29d29b5};
test_output[6942] = '{32'h42b15f6d};
test_index[6942] = '{4};
test_input[55544:55551] = '{32'h421d3df3, 32'h429ea45b, 32'h42a24095, 32'hc14b991b, 32'hc23096c7, 32'h419c3738, 32'h41deb65c, 32'hc28986b6};
test_output[6943] = '{32'h42a24095};
test_index[6943] = '{2};
test_input[55552:55559] = '{32'hc274930d, 32'h4191253d, 32'h42515248, 32'h4282764c, 32'h427128a4, 32'h41f48a27, 32'hc2a742d2, 32'hc2aefcd3};
test_output[6944] = '{32'h4282764c};
test_index[6944] = '{3};
test_input[55560:55567] = '{32'hc1f4fc7e, 32'h426495a7, 32'h421a3550, 32'h429359a0, 32'h41dda483, 32'h41f1e974, 32'h42c6e065, 32'h42ac325d};
test_output[6945] = '{32'h42c6e065};
test_index[6945] = '{6};
test_input[55568:55575] = '{32'hc1d1b941, 32'h42a2573a, 32'h429e8e5b, 32'hbfbc8d5c, 32'h4291e8ff, 32'hc2b94147, 32'h422c2c81, 32'h42bfe0a7};
test_output[6946] = '{32'h42bfe0a7};
test_index[6946] = '{7};
test_input[55576:55583] = '{32'h420ab89f, 32'hc25b5118, 32'h41cde1c3, 32'hc2a14f6a, 32'hbf0b2d8b, 32'hc21414c6, 32'h42045643, 32'hc2a3ff4a};
test_output[6947] = '{32'h420ab89f};
test_index[6947] = '{0};
test_input[55584:55591] = '{32'hc18e6f11, 32'hc28ecfbc, 32'hc1a609c6, 32'h427988e6, 32'hc034f16b, 32'hc2a0142e, 32'h40bc9e20, 32'hc24d67fd};
test_output[6948] = '{32'h427988e6};
test_index[6948] = '{3};
test_input[55592:55599] = '{32'hc2bc1b9a, 32'h42c06003, 32'h42593a82, 32'hc2a58855, 32'h423cd95c, 32'h41a8eb94, 32'h427c2c8c, 32'hc16ae7c7};
test_output[6949] = '{32'h42c06003};
test_index[6949] = '{1};
test_input[55600:55607] = '{32'h418d8102, 32'h42891cea, 32'hc2370b7d, 32'h429ebeb1, 32'hc2273bf0, 32'hc24ae11d, 32'h3e9f16d2, 32'hc207521f};
test_output[6950] = '{32'h429ebeb1};
test_index[6950] = '{3};
test_input[55608:55615] = '{32'hc10b932c, 32'h429d31db, 32'h426c7fca, 32'h4102bf4e, 32'h4087e8ef, 32'hc294cc6a, 32'h41e7fc25, 32'h4077802b};
test_output[6951] = '{32'h429d31db};
test_index[6951] = '{1};
test_input[55616:55623] = '{32'hbb5167e1, 32'hc28aa434, 32'h4255c9bb, 32'hc268340f, 32'hc285a8fc, 32'h41d575d8, 32'h428ad718, 32'h42b08361};
test_output[6952] = '{32'h42b08361};
test_index[6952] = '{7};
test_input[55624:55631] = '{32'h41e48488, 32'h422e1bad, 32'hc00ee286, 32'hc22f1230, 32'h429d23af, 32'h4251d725, 32'hc2c609bc, 32'h4205032c};
test_output[6953] = '{32'h429d23af};
test_index[6953] = '{4};
test_input[55632:55639] = '{32'h404bfa93, 32'h42ad04ac, 32'h41d235e1, 32'h41e0f7ab, 32'hc21d8ec3, 32'h42a49ce9, 32'h3ff86d04, 32'hc1f4186d};
test_output[6954] = '{32'h42ad04ac};
test_index[6954] = '{1};
test_input[55640:55647] = '{32'h42325d6b, 32'hc2952024, 32'hc1cd031e, 32'h4273b244, 32'h40fe10f0, 32'hc290523b, 32'h41b81557, 32'h42895e0f};
test_output[6955] = '{32'h42895e0f};
test_index[6955] = '{7};
test_input[55648:55655] = '{32'h3ffe79c8, 32'h42083beb, 32'hc2914ca1, 32'hbf58cb97, 32'h41e6d6ee, 32'hc2b349ab, 32'hc2999cca, 32'hc2bee67a};
test_output[6956] = '{32'h42083beb};
test_index[6956] = '{1};
test_input[55656:55663] = '{32'h4200c248, 32'hc1aa38bb, 32'hc1870180, 32'h4298d437, 32'h42c6f806, 32'h422bc926, 32'hc224bcff, 32'hc2b47aa9};
test_output[6957] = '{32'h42c6f806};
test_index[6957] = '{4};
test_input[55664:55671] = '{32'h4185886e, 32'hc23b7aae, 32'hc140d342, 32'hc29b9ad8, 32'h42a8d357, 32'hc28b150f, 32'h42a41191, 32'hc28defba};
test_output[6958] = '{32'h42a8d357};
test_index[6958] = '{4};
test_input[55672:55679] = '{32'hc0ab53f6, 32'hc2395f44, 32'hc1821af3, 32'h41a2d2bb, 32'h414e4564, 32'hc2796be2, 32'hc2349153, 32'h42b0f90a};
test_output[6959] = '{32'h42b0f90a};
test_index[6959] = '{7};
test_input[55680:55687] = '{32'h4282b379, 32'hc04cc0ff, 32'h41a3a7fe, 32'hc19dcbad, 32'hc20253da, 32'h42620f55, 32'hc2970354, 32'hc23b4330};
test_output[6960] = '{32'h4282b379};
test_index[6960] = '{0};
test_input[55688:55695] = '{32'hc2b4283d, 32'hc0a57283, 32'hc2768ac7, 32'h42c11fc9, 32'h42c5f7a9, 32'hc073d99a, 32'h41035464, 32'h425e41d9};
test_output[6961] = '{32'h42c5f7a9};
test_index[6961] = '{4};
test_input[55696:55703] = '{32'hc2a20794, 32'hbf13d179, 32'hc1977001, 32'h42a590e4, 32'h42a258ef, 32'hc22632c4, 32'h427c64a0, 32'hc284bdad};
test_output[6962] = '{32'h42a590e4};
test_index[6962] = '{3};
test_input[55704:55711] = '{32'h4258f5ff, 32'h42a69b4a, 32'h41d6c306, 32'hc2b95b07, 32'h4238853e, 32'h4201f58a, 32'h42715986, 32'h41b7f0e3};
test_output[6963] = '{32'h42a69b4a};
test_index[6963] = '{1};
test_input[55712:55719] = '{32'h42a4d088, 32'h4236afd2, 32'hc218c2d1, 32'hc1f5f4ff, 32'hc2125fec, 32'h42c3b3ae, 32'hc1d620e1, 32'h4232dedc};
test_output[6964] = '{32'h42c3b3ae};
test_index[6964] = '{5};
test_input[55720:55727] = '{32'h4231a225, 32'h408a64c9, 32'hc1b3751b, 32'h41c7ece4, 32'h420413f0, 32'hc2849fbf, 32'h4213a013, 32'hc26e75cc};
test_output[6965] = '{32'h4231a225};
test_index[6965] = '{0};
test_input[55728:55735] = '{32'hc290fcad, 32'hc2c0cc90, 32'hc2606967, 32'h424850d6, 32'h429d7e5b, 32'h42bae9fe, 32'hc23572a9, 32'h419901ae};
test_output[6966] = '{32'h42bae9fe};
test_index[6966] = '{5};
test_input[55736:55743] = '{32'h420f1aa9, 32'h41316b5f, 32'hc0f2104a, 32'h413b7d7e, 32'hc28a42f0, 32'hc02f7427, 32'hc2a53c76, 32'hc288f0d5};
test_output[6967] = '{32'h420f1aa9};
test_index[6967] = '{0};
test_input[55744:55751] = '{32'hc28b54d2, 32'h4115ae86, 32'hc237bd42, 32'h42b7a3a7, 32'hc185a855, 32'h42768933, 32'hc26920a1, 32'h429172bb};
test_output[6968] = '{32'h42b7a3a7};
test_index[6968] = '{3};
test_input[55752:55759] = '{32'h4239aca1, 32'h420217ae, 32'h42af870b, 32'h42a45a17, 32'h423df87b, 32'h42b6ae3a, 32'hc251da7a, 32'h41a5db34};
test_output[6969] = '{32'h42b6ae3a};
test_index[6969] = '{5};
test_input[55760:55767] = '{32'hc00c18b4, 32'h40d41850, 32'hc2813c31, 32'hc19b5550, 32'hc2233e37, 32'h42392141, 32'hc286fdee, 32'h4235902e};
test_output[6970] = '{32'h42392141};
test_index[6970] = '{5};
test_input[55768:55775] = '{32'hc24d7805, 32'h425ea471, 32'h41ce6fd7, 32'hc2c49484, 32'h419de29e, 32'hc1dd5d7a, 32'h42a0dfa0, 32'h42c6a89a};
test_output[6971] = '{32'h42c6a89a};
test_index[6971] = '{7};
test_input[55776:55783] = '{32'h42a6c2cc, 32'hc2a33fef, 32'hc14a90ed, 32'hc25174ac, 32'h426354ec, 32'h40ab1c53, 32'hc198c479, 32'hc2aac386};
test_output[6972] = '{32'h42a6c2cc};
test_index[6972] = '{0};
test_input[55784:55791] = '{32'h42619157, 32'h426ea312, 32'hc2935080, 32'h42c3827d, 32'hc267e35e, 32'hc274004f, 32'h4245d082, 32'h42414c9b};
test_output[6973] = '{32'h42c3827d};
test_index[6973] = '{3};
test_input[55792:55799] = '{32'hc0c475e4, 32'h42ba6ceb, 32'h423fa616, 32'hc29d78ff, 32'hc2a5c704, 32'hc22fd51e, 32'h420a75cf, 32'h42661a73};
test_output[6974] = '{32'h42ba6ceb};
test_index[6974] = '{1};
test_input[55800:55807] = '{32'h42b0332f, 32'hc276b7be, 32'hc29ab631, 32'hc240439b, 32'hc297dcdc, 32'h428f43fc, 32'h4044547f, 32'h426c577b};
test_output[6975] = '{32'h42b0332f};
test_index[6975] = '{0};
test_input[55808:55815] = '{32'hc23eb9d2, 32'hc231d232, 32'h41b2e1b6, 32'h402cfa0b, 32'hc2b398f7, 32'hc19a45a9, 32'h429e1072, 32'h42bf22ff};
test_output[6976] = '{32'h42bf22ff};
test_index[6976] = '{7};
test_input[55816:55823] = '{32'hc26f18e7, 32'hc152f584, 32'h41062a8b, 32'h426c6f6f, 32'hc21add6c, 32'hc223fb24, 32'h42a8f6f7, 32'hc24921f2};
test_output[6977] = '{32'h42a8f6f7};
test_index[6977] = '{6};
test_input[55824:55831] = '{32'h42513644, 32'h41c5f574, 32'h421cf31a, 32'hc2bfe5e9, 32'hc2b9b40d, 32'hc24518fd, 32'hc2b198e3, 32'h42b952e0};
test_output[6978] = '{32'h42b952e0};
test_index[6978] = '{7};
test_input[55832:55839] = '{32'hc11e6c10, 32'h403d14f2, 32'hc242bf52, 32'h42863370, 32'hc1ac4b22, 32'h42a71a28, 32'h4291a6eb, 32'h41d3dac9};
test_output[6979] = '{32'h42a71a28};
test_index[6979] = '{5};
test_input[55840:55847] = '{32'hc211a470, 32'h429a95f0, 32'hc29cc691, 32'h420f3d8c, 32'hc1e7d93c, 32'hc0b506f9, 32'hc28c21c2, 32'hc17bfe4b};
test_output[6980] = '{32'h429a95f0};
test_index[6980] = '{1};
test_input[55848:55855] = '{32'h42c6ee30, 32'h417d8e17, 32'hc0ffaaf5, 32'h42af6bcd, 32'hc254cdec, 32'h424b29f5, 32'h42a10de5, 32'hc1b6712e};
test_output[6981] = '{32'h42c6ee30};
test_index[6981] = '{0};
test_input[55856:55863] = '{32'h42248bf6, 32'h400e2530, 32'h42b2d2c6, 32'h4280a334, 32'h42654190, 32'hc2ac7303, 32'hc267da2a, 32'h4175ddf0};
test_output[6982] = '{32'h42b2d2c6};
test_index[6982] = '{2};
test_input[55864:55871] = '{32'h42a8e63c, 32'h42a08881, 32'h420724e5, 32'hc2a72bea, 32'hc2c2dedb, 32'h42be6650, 32'hc191b1bd, 32'h4258020a};
test_output[6983] = '{32'h42be6650};
test_index[6983] = '{5};
test_input[55872:55879] = '{32'h42467670, 32'hc254bfeb, 32'hc20b4a2a, 32'hc282d75e, 32'hc29b5cfb, 32'hc16925df, 32'h420cbbae, 32'h42286525};
test_output[6984] = '{32'h42467670};
test_index[6984] = '{0};
test_input[55880:55887] = '{32'h4265434e, 32'hc291b110, 32'hc1b295c1, 32'h42a72975, 32'h4256e53b, 32'h42ad5343, 32'hc2b673b5, 32'h4265e97b};
test_output[6985] = '{32'h42ad5343};
test_index[6985] = '{5};
test_input[55888:55895] = '{32'hc0f8a271, 32'h41a03a15, 32'h42488c56, 32'h42c70f75, 32'h4253e0af, 32'hc1e42f3f, 32'h428dd091, 32'h42525bfb};
test_output[6986] = '{32'h42c70f75};
test_index[6986] = '{3};
test_input[55896:55903] = '{32'hc26f7ef3, 32'hc22f4d30, 32'h426a0e78, 32'hc122a7e5, 32'hc1aa0908, 32'hc1e74f38, 32'h4126a7bb, 32'hc1cf2a2f};
test_output[6987] = '{32'h426a0e78};
test_index[6987] = '{2};
test_input[55904:55911] = '{32'hc29a9c9a, 32'h425f9a74, 32'h42a5b93b, 32'hc1e0ff61, 32'hc298a08d, 32'hc22d0c3c, 32'hc1d4e10b, 32'h3f4e5e23};
test_output[6988] = '{32'h42a5b93b};
test_index[6988] = '{2};
test_input[55912:55919] = '{32'hc271cb8a, 32'h4277859d, 32'h429e3e8f, 32'h4196ccc1, 32'h4262a29b, 32'h426ab863, 32'hc1d3a771, 32'hc14be458};
test_output[6989] = '{32'h429e3e8f};
test_index[6989] = '{2};
test_input[55920:55927] = '{32'hc2931a33, 32'hc2a1a1f5, 32'h42152171, 32'h42591e0f, 32'h410b80f0, 32'hc2803b65, 32'hc2ba9883, 32'h42852caf};
test_output[6990] = '{32'h42852caf};
test_index[6990] = '{7};
test_input[55928:55935] = '{32'h42c1d601, 32'hc2ad12ca, 32'h428d2362, 32'hc25903b4, 32'hc22719b4, 32'hc182fb15, 32'hc1944d50, 32'h42aad825};
test_output[6991] = '{32'h42c1d601};
test_index[6991] = '{0};
test_input[55936:55943] = '{32'hc1dc80e0, 32'hc1afb9ee, 32'hc227ec87, 32'h429748ef, 32'hc2891455, 32'h427d19f0, 32'h41834b40, 32'h429249c5};
test_output[6992] = '{32'h429748ef};
test_index[6992] = '{3};
test_input[55944:55951] = '{32'hc228837d, 32'h428c3264, 32'hc201f7ff, 32'h422d020a, 32'h42615be6, 32'hc2ab3698, 32'hc2b5bc96, 32'hc2933e7d};
test_output[6993] = '{32'h428c3264};
test_index[6993] = '{1};
test_input[55952:55959] = '{32'hc0c3728b, 32'hc103d03c, 32'h41caf2f0, 32'h42bb36cc, 32'hc233c514, 32'hc23c5d69, 32'hc1abe67d, 32'hc0d7f374};
test_output[6994] = '{32'h42bb36cc};
test_index[6994] = '{3};
test_input[55960:55967] = '{32'h4289f339, 32'hc2313bb6, 32'h40972b4b, 32'h420aaa88, 32'h429940d8, 32'h42bd8e03, 32'h41ab8f17, 32'h406bc4a5};
test_output[6995] = '{32'h42bd8e03};
test_index[6995] = '{5};
test_input[55968:55975] = '{32'h4224ce1c, 32'hc2a43cc0, 32'hc2aa2424, 32'h429ce4cf, 32'hc28b8415, 32'h425808c6, 32'h4288d9df, 32'h42c4a037};
test_output[6996] = '{32'h42c4a037};
test_index[6996] = '{7};
test_input[55976:55983] = '{32'h42951916, 32'h42336105, 32'h420c206b, 32'h422f8358, 32'hc2436b2a, 32'hc264e370, 32'h41e97a06, 32'hc1a52231};
test_output[6997] = '{32'h42951916};
test_index[6997] = '{0};
test_input[55984:55991] = '{32'hc1a5c288, 32'h4279bf89, 32'hc2a4bfb5, 32'hc2aad390, 32'h42833c6a, 32'hc23ae6ab, 32'h424826c3, 32'h400b8b81};
test_output[6998] = '{32'h42833c6a};
test_index[6998] = '{4};
test_input[55992:55999] = '{32'h42092f22, 32'hc269c9b7, 32'h40c6e8cb, 32'hc193aed3, 32'h41ff035b, 32'h428aa322, 32'hc2b23a23, 32'hc217abc9};
test_output[6999] = '{32'h428aa322};
test_index[6999] = '{5};
test_input[56000:56007] = '{32'h429cd73f, 32'h425405f3, 32'hc244570c, 32'hc0401dd7, 32'hc231129e, 32'hc29ef410, 32'hc28b6804, 32'hbec87e51};
test_output[7000] = '{32'h429cd73f};
test_index[7000] = '{0};
test_input[56008:56015] = '{32'h410317c3, 32'h421fa5ad, 32'h421e625c, 32'h41a466f9, 32'h4190acc6, 32'hc2982e46, 32'h3feaf9f0, 32'h428df334};
test_output[7001] = '{32'h428df334};
test_index[7001] = '{7};
test_input[56016:56023] = '{32'hc2c3b81e, 32'h4262dbe7, 32'h4277f218, 32'hc297b0a3, 32'hc1b3c007, 32'h420b7389, 32'h428e958b, 32'hc1d08036};
test_output[7002] = '{32'h428e958b};
test_index[7002] = '{6};
test_input[56024:56031] = '{32'hc28e1535, 32'hc1dd3f39, 32'hc22f77a1, 32'h41a2668b, 32'hc239c26d, 32'hc286aac2, 32'hc2c19a17, 32'h427a134e};
test_output[7003] = '{32'h427a134e};
test_index[7003] = '{7};
test_input[56032:56039] = '{32'hc251c42b, 32'hc2380972, 32'h420c1d6b, 32'h42a272da, 32'hc2675cbf, 32'h41d93b44, 32'h427fc79a, 32'hc26a4a3d};
test_output[7004] = '{32'h42a272da};
test_index[7004] = '{3};
test_input[56040:56047] = '{32'hc1e3474d, 32'hc2a63715, 32'h41ce8354, 32'hc1c55d76, 32'h427cb1c0, 32'hc2253a64, 32'hc27ec1cc, 32'hc24c5166};
test_output[7005] = '{32'h427cb1c0};
test_index[7005] = '{4};
test_input[56048:56055] = '{32'hc0b735f9, 32'hc29f3bd3, 32'h426694db, 32'hc28685a6, 32'h429591a8, 32'hc2c68196, 32'h42a9693a, 32'h4250888b};
test_output[7006] = '{32'h42a9693a};
test_index[7006] = '{6};
test_input[56056:56063] = '{32'h420853b6, 32'h41c50a12, 32'hc17603bb, 32'hc267bf48, 32'h42034492, 32'h428ec8f0, 32'hc28af06b, 32'h42b9a832};
test_output[7007] = '{32'h42b9a832};
test_index[7007] = '{7};
test_input[56064:56071] = '{32'hc28c76c0, 32'h40b829d0, 32'hc2799ae9, 32'h428212d3, 32'hc2446925, 32'h429c228f, 32'hc29ebe9c, 32'hc1f8195c};
test_output[7008] = '{32'h429c228f};
test_index[7008] = '{5};
test_input[56072:56079] = '{32'hc11780b8, 32'hc24e6d6d, 32'h4271849f, 32'hc2904149, 32'h41c26702, 32'hc0e5c321, 32'hc1d8d31d, 32'hc2a08432};
test_output[7009] = '{32'h4271849f};
test_index[7009] = '{2};
test_input[56080:56087] = '{32'h429b435a, 32'hc2491bb8, 32'h42830e30, 32'h42b4d4e9, 32'h42868f5b, 32'hc29ac727, 32'h42b96ac5, 32'hc1df26cf};
test_output[7010] = '{32'h42b96ac5};
test_index[7010] = '{6};
test_input[56088:56095] = '{32'h421424be, 32'h42bd9097, 32'h425638a6, 32'hc24c2705, 32'hc0bf8e35, 32'hc0aa63a1, 32'h41911e70, 32'hc289d10e};
test_output[7011] = '{32'h42bd9097};
test_index[7011] = '{1};
test_input[56096:56103] = '{32'hc1f746df, 32'hc20aa742, 32'h402f93a8, 32'hc2be7e72, 32'hc1a9d460, 32'hc2afab2d, 32'h427c5d00, 32'h4271b98d};
test_output[7012] = '{32'h427c5d00};
test_index[7012] = '{6};
test_input[56104:56111] = '{32'hc24c204a, 32'hc19e2676, 32'hc2bc6a2c, 32'h40baf665, 32'hc280f4ee, 32'h4284ca93, 32'h4068df2b, 32'hc29902a3};
test_output[7013] = '{32'h4284ca93};
test_index[7013] = '{5};
test_input[56112:56119] = '{32'hc23a90fe, 32'hc180a9c2, 32'h41d50851, 32'h41635349, 32'hc297efc3, 32'h41f2f97b, 32'h42c2f633, 32'h42b54139};
test_output[7014] = '{32'h42c2f633};
test_index[7014] = '{6};
test_input[56120:56127] = '{32'h3ff13017, 32'hc25882c4, 32'hc1ba7bc6, 32'hc2b468e9, 32'h42bf6f82, 32'hc2945a41, 32'hc0aaf806, 32'hc2b5c49f};
test_output[7015] = '{32'h42bf6f82};
test_index[7015] = '{4};
test_input[56128:56135] = '{32'hc13d8d3f, 32'hc1282733, 32'h41affeb9, 32'hc26f32db, 32'h42b57444, 32'hc291e6b5, 32'h41121f71, 32'hc1d334fd};
test_output[7016] = '{32'h42b57444};
test_index[7016] = '{4};
test_input[56136:56143] = '{32'h428b01c4, 32'hc2943589, 32'h428fc1d9, 32'h3f04a8c8, 32'hc29da2dc, 32'h42c1dd41, 32'hc2762889, 32'hc1d8d176};
test_output[7017] = '{32'h42c1dd41};
test_index[7017] = '{5};
test_input[56144:56151] = '{32'h4271eea5, 32'hc244efe8, 32'hc016aac6, 32'hc2c4ed26, 32'hc228f48f, 32'h42b8b06a, 32'h42ab2778, 32'hc23f5b35};
test_output[7018] = '{32'h42b8b06a};
test_index[7018] = '{5};
test_input[56152:56159] = '{32'hc29e939e, 32'hc29e5d5a, 32'hc21d71eb, 32'hc1b384f0, 32'hc28af25d, 32'h42a8d45e, 32'h42b83a73, 32'h42ae707c};
test_output[7019] = '{32'h42b83a73};
test_index[7019] = '{6};
test_input[56160:56167] = '{32'h427c5275, 32'hc1cb3289, 32'h422906b2, 32'h42c073e9, 32'h42b44c0c, 32'h42017fbc, 32'hc24630cb, 32'h42aa0cf3};
test_output[7020] = '{32'h42c073e9};
test_index[7020] = '{3};
test_input[56168:56175] = '{32'h4233423d, 32'h42a998e9, 32'hc2ad7068, 32'hc2b19382, 32'hc2a718ed, 32'h42bc54ff, 32'h42444f48, 32'h4254c318};
test_output[7021] = '{32'h42bc54ff};
test_index[7021] = '{5};
test_input[56176:56183] = '{32'h42b2ea89, 32'h4292dab4, 32'h42260835, 32'hc2aafec6, 32'hc24ddd01, 32'h41c5fba1, 32'h426f7471, 32'h426377bf};
test_output[7022] = '{32'h42b2ea89};
test_index[7022] = '{0};
test_input[56184:56191] = '{32'h42c2cb14, 32'hc250a9d4, 32'hc26d94e7, 32'h42c30cb3, 32'h4102056a, 32'h42769c3d, 32'hc290376a, 32'h42bb6b39};
test_output[7023] = '{32'h42c30cb3};
test_index[7023] = '{3};
test_input[56192:56199] = '{32'h412a7364, 32'hc11003b5, 32'hbf207567, 32'h42bc9276, 32'hc1ac447c, 32'h4145b0ed, 32'h4286b24d, 32'hc209dac3};
test_output[7024] = '{32'h42bc9276};
test_index[7024] = '{3};
test_input[56200:56207] = '{32'hc2558725, 32'hc17ba90f, 32'hc2c2a884, 32'hc1a71d8d, 32'hc18006e0, 32'hc26876eb, 32'hc18006bc, 32'h42493af6};
test_output[7025] = '{32'h42493af6};
test_index[7025] = '{7};
test_input[56208:56215] = '{32'h42932374, 32'hc149a87a, 32'h42a5a3ba, 32'hc1191c9a, 32'hc29a0cb6, 32'h42901116, 32'h421030fe, 32'hc29b00d3};
test_output[7026] = '{32'h42a5a3ba};
test_index[7026] = '{2};
test_input[56216:56223] = '{32'hc2943846, 32'h428bf8a2, 32'hc297741f, 32'h415372fb, 32'hc1bb04f5, 32'hbf45e2d7, 32'hc22471ba, 32'hc29d583a};
test_output[7027] = '{32'h428bf8a2};
test_index[7027] = '{1};
test_input[56224:56231] = '{32'h4247ed08, 32'h428ab37b, 32'h42ae0925, 32'h42b1cfb6, 32'hc183a243, 32'h40e71d5e, 32'hc1826909, 32'hc2be0286};
test_output[7028] = '{32'h42b1cfb6};
test_index[7028] = '{3};
test_input[56232:56239] = '{32'h41675937, 32'hc2c31727, 32'h4267959b, 32'h428f7f1a, 32'h428f7f88, 32'hc0d22863, 32'h410888f3, 32'h42c1c0eb};
test_output[7029] = '{32'h42c1c0eb};
test_index[7029] = '{7};
test_input[56240:56247] = '{32'hc22f2f91, 32'h42ac1457, 32'hc2832b3b, 32'hc286aae1, 32'h427e414b, 32'hc265a31c, 32'hc2006e55, 32'hc214be41};
test_output[7030] = '{32'h42ac1457};
test_index[7030] = '{1};
test_input[56248:56255] = '{32'hc251582e, 32'hc2a8ea67, 32'h428689ad, 32'h429cb3d5, 32'hc238bee1, 32'h41b014d4, 32'h420e348a, 32'hc2509a0a};
test_output[7031] = '{32'h429cb3d5};
test_index[7031] = '{3};
test_input[56256:56263] = '{32'h4191d1c5, 32'h4279228c, 32'h4281ab65, 32'h41a01319, 32'h41d3192a, 32'h429c739a, 32'h424a9dee, 32'h41f303ab};
test_output[7032] = '{32'h429c739a};
test_index[7032] = '{5};
test_input[56264:56271] = '{32'h42ac83bf, 32'hc28ffb02, 32'h42094e8a, 32'hc2128cfb, 32'h42863e67, 32'hc2c76872, 32'hc28c6a8a, 32'h41b0aea7};
test_output[7033] = '{32'h42ac83bf};
test_index[7033] = '{0};
test_input[56272:56279] = '{32'hc185bd4e, 32'h42ad787a, 32'hc1b2ebe0, 32'h4299fc7e, 32'hbff0bb80, 32'h42abc34b, 32'h42c4c6d5, 32'hc2c35451};
test_output[7034] = '{32'h42c4c6d5};
test_index[7034] = '{6};
test_input[56280:56287] = '{32'hc227b640, 32'hc2be2ba1, 32'h417475c3, 32'hc296c652, 32'h41a92c15, 32'hc27dfb95, 32'h42141496, 32'hc247bf75};
test_output[7035] = '{32'h42141496};
test_index[7035] = '{6};
test_input[56288:56295] = '{32'h42897142, 32'h41d9fb03, 32'h42a4d984, 32'h4229265f, 32'h418b4327, 32'hc13105ef, 32'hc25e6b04, 32'hc27b6211};
test_output[7036] = '{32'h42a4d984};
test_index[7036] = '{2};
test_input[56296:56303] = '{32'h3f052b3d, 32'h42613e85, 32'h42c713f8, 32'hbfd4fdf6, 32'h42b87c3a, 32'h414afba7, 32'h42c1c05a, 32'hc11ef4da};
test_output[7037] = '{32'h42c713f8};
test_index[7037] = '{2};
test_input[56304:56311] = '{32'hc2c7d3c9, 32'h421bb70c, 32'hbf8c09b4, 32'hc1961723, 32'hc28b1b3b, 32'h4056d952, 32'hc2bb47b1, 32'hc20299cb};
test_output[7038] = '{32'h421bb70c};
test_index[7038] = '{1};
test_input[56312:56319] = '{32'h423ccec7, 32'hc124803c, 32'h425047b4, 32'hc2930cfb, 32'h41e8c391, 32'hc2b98c58, 32'h40d2efac, 32'h427222ce};
test_output[7039] = '{32'h427222ce};
test_index[7039] = '{7};
test_input[56320:56327] = '{32'h42a686b6, 32'hc29fcb0e, 32'h42b121b8, 32'h425767d6, 32'hc056ef16, 32'h42b544fa, 32'h4151b98a, 32'hc2a456ea};
test_output[7040] = '{32'h42b544fa};
test_index[7040] = '{5};
test_input[56328:56335] = '{32'hc0eb1b4e, 32'h424f45b2, 32'h4149b8ae, 32'hc1c3d7e0, 32'hc2708d90, 32'h3e02be4e, 32'hc218b999, 32'hc2915527};
test_output[7041] = '{32'h424f45b2};
test_index[7041] = '{1};
test_input[56336:56343] = '{32'hc15e5249, 32'h41cb3d79, 32'hc22432a4, 32'h428eb8a0, 32'hc27fe5d9, 32'hc1e7f5ed, 32'hc2b07b06, 32'h41af8e2c};
test_output[7042] = '{32'h428eb8a0};
test_index[7042] = '{3};
test_input[56344:56351] = '{32'h42b5b8b2, 32'h424807f8, 32'h42b7d294, 32'hc29e84a1, 32'h42a3b679, 32'h42c77b4e, 32'h424ba7f6, 32'hc28d95c5};
test_output[7043] = '{32'h42c77b4e};
test_index[7043] = '{5};
test_input[56352:56359] = '{32'h424bf6a1, 32'hc23ce5ae, 32'h418ac234, 32'h42c756be, 32'hc25264a1, 32'h4272aa4a, 32'hbf255f8d, 32'hc2bb876c};
test_output[7044] = '{32'h42c756be};
test_index[7044] = '{3};
test_input[56360:56367] = '{32'h42a23d59, 32'hc22bbb9b, 32'h428b2e6d, 32'h422d0816, 32'hc25a46be, 32'h428d3880, 32'h42c3f447, 32'h4244f441};
test_output[7045] = '{32'h42c3f447};
test_index[7045] = '{6};
test_input[56368:56375] = '{32'h42c34fe5, 32'hc2a6d8a1, 32'hc26a4fdb, 32'h42c6ce40, 32'hc2bc49be, 32'hc2579bb8, 32'hbf0bf252, 32'hc2222bd6};
test_output[7046] = '{32'h42c6ce40};
test_index[7046] = '{3};
test_input[56376:56383] = '{32'h4186a2bb, 32'hc2837e56, 32'hc275b891, 32'hc27778d6, 32'hc1502630, 32'h42244883, 32'hc282eb66, 32'hc2bb229f};
test_output[7047] = '{32'h42244883};
test_index[7047] = '{5};
test_input[56384:56391] = '{32'hc278fde4, 32'hc2a1b5de, 32'h40e0aa0e, 32'hc15bb9f8, 32'hc255e076, 32'h41ff72df, 32'h42127432, 32'hc202a07e};
test_output[7048] = '{32'h42127432};
test_index[7048] = '{6};
test_input[56392:56399] = '{32'h422d9230, 32'hc2294868, 32'hc1e6d60f, 32'hc2a0fb06, 32'hc1fbc660, 32'h42adc318, 32'hc2861c8b, 32'h420689f9};
test_output[7049] = '{32'h42adc318};
test_index[7049] = '{5};
test_input[56400:56407] = '{32'h42bb17d4, 32'hc2558237, 32'hc2203159, 32'hc2680519, 32'h4246ce1b, 32'hc1be310d, 32'h42a2819b, 32'hbfe38559};
test_output[7050] = '{32'h42bb17d4};
test_index[7050] = '{0};
test_input[56408:56415] = '{32'h422c3b44, 32'h4244c43a, 32'h3fe2f210, 32'h4260af10, 32'hc21039c6, 32'h42096736, 32'hc100d21a, 32'hc2be5e82};
test_output[7051] = '{32'h4260af10};
test_index[7051] = '{3};
test_input[56416:56423] = '{32'hc2bf58fb, 32'h42a009b9, 32'h423c566b, 32'h42a835e3, 32'h425e211e, 32'h415d86d0, 32'h42bf801f, 32'hc1d201bb};
test_output[7052] = '{32'h42bf801f};
test_index[7052] = '{6};
test_input[56424:56431] = '{32'h426c7529, 32'h4141f1a3, 32'h42b77b60, 32'h4252123b, 32'h40c4e58c, 32'hc26ca0c4, 32'hc1bdb7a7, 32'h4219524d};
test_output[7053] = '{32'h42b77b60};
test_index[7053] = '{2};
test_input[56432:56439] = '{32'h4194129d, 32'hc237a494, 32'hc2a4a33c, 32'h4238641c, 32'hc1f8660a, 32'hc151d243, 32'hc293497b, 32'h428f1ea3};
test_output[7054] = '{32'h428f1ea3};
test_index[7054] = '{7};
test_input[56440:56447] = '{32'h429a0574, 32'hc2ab293a, 32'h420a48ca, 32'h42b5b6cb, 32'h41097e2f, 32'h41e268dc, 32'hc279396e, 32'hc25c87df};
test_output[7055] = '{32'h42b5b6cb};
test_index[7055] = '{3};
test_input[56448:56455] = '{32'hc187e238, 32'hc2870090, 32'h42c3fcb9, 32'hc256a37d, 32'hc1a1cd21, 32'h422ee800, 32'hc2800b7d, 32'hc1d6d6df};
test_output[7056] = '{32'h42c3fcb9};
test_index[7056] = '{2};
test_input[56456:56463] = '{32'h41fa7089, 32'h426cd474, 32'hc225b1d7, 32'h4292e99a, 32'hc28f70cc, 32'h42891d9c, 32'h42003ead, 32'hc28de5d9};
test_output[7057] = '{32'h4292e99a};
test_index[7057] = '{3};
test_input[56464:56471] = '{32'h4292aba9, 32'h42725997, 32'hc2b90d2f, 32'hc1860a0b, 32'hc1828133, 32'hc2c6c293, 32'h426c62b2, 32'h42bfb544};
test_output[7058] = '{32'h42bfb544};
test_index[7058] = '{7};
test_input[56472:56479] = '{32'hc22b357d, 32'h42a4a8ae, 32'h421311e0, 32'h420778e7, 32'hc29863f2, 32'hc2b072a5, 32'h42acbfa6, 32'h4140bf8f};
test_output[7059] = '{32'h42acbfa6};
test_index[7059] = '{6};
test_input[56480:56487] = '{32'hc191437e, 32'hc129a39e, 32'hc2ab04a7, 32'hc2b2a197, 32'h422a6461, 32'hc201fc2f, 32'hc2640df1, 32'h41671c08};
test_output[7060] = '{32'h422a6461};
test_index[7060] = '{4};
test_input[56488:56495] = '{32'h42454ad5, 32'h42c2e4f4, 32'hc18d8ef3, 32'h41935baf, 32'h3fd93187, 32'h422652cb, 32'h42a24a76, 32'hc260d7db};
test_output[7061] = '{32'h42c2e4f4};
test_index[7061] = '{1};
test_input[56496:56503] = '{32'hc2b8b002, 32'hc2c3e30c, 32'h42a74e1c, 32'hc29f4696, 32'h4297704a, 32'hc009b1b9, 32'h419dfbba, 32'h425c15b5};
test_output[7062] = '{32'h42a74e1c};
test_index[7062] = '{2};
test_input[56504:56511] = '{32'hc15f7d73, 32'h40dc7488, 32'h4250be19, 32'h4212db27, 32'hc26815f8, 32'h42273bf2, 32'h42b50d0d, 32'hc296e7ee};
test_output[7063] = '{32'h42b50d0d};
test_index[7063] = '{6};
test_input[56512:56519] = '{32'h41ccc6df, 32'hc27d5f8c, 32'h41c18022, 32'hc28d198f, 32'hc24d904b, 32'h4235d586, 32'h42253e07, 32'hc125d6be};
test_output[7064] = '{32'h4235d586};
test_index[7064] = '{5};
test_input[56520:56527] = '{32'hc2874cfd, 32'h429146a1, 32'hc2a16585, 32'hc2c2f93b, 32'hc15e6f7f, 32'hc2650890, 32'h428df0b3, 32'h41ca40b3};
test_output[7065] = '{32'h429146a1};
test_index[7065] = '{1};
test_input[56528:56535] = '{32'h4257f758, 32'h41880900, 32'h4228cc5d, 32'h422665ba, 32'h42826b27, 32'hc280c1b5, 32'h4151203f, 32'hc2ac6b73};
test_output[7066] = '{32'h42826b27};
test_index[7066] = '{4};
test_input[56536:56543] = '{32'h4287cb2d, 32'hc29b8d3b, 32'h42668cd9, 32'hc212e002, 32'hc23b967e, 32'h429ab4ac, 32'h41de476e, 32'h42a6e8b6};
test_output[7067] = '{32'h42a6e8b6};
test_index[7067] = '{7};
test_input[56544:56551] = '{32'hc29b5bce, 32'hc2c5c4ed, 32'hc234486e, 32'h4286fcf9, 32'hc00d513d, 32'h42abc2c9, 32'h4267153c, 32'h3f3caa32};
test_output[7068] = '{32'h42abc2c9};
test_index[7068] = '{5};
test_input[56552:56559] = '{32'hbecf6de8, 32'h428bf3fd, 32'h417557ff, 32'hc27b063e, 32'hc2347248, 32'h41a2827e, 32'hc23d2a8f, 32'hc1da0393};
test_output[7069] = '{32'h428bf3fd};
test_index[7069] = '{1};
test_input[56560:56567] = '{32'hc272a224, 32'hc182f247, 32'h42b12a3b, 32'h42522608, 32'hc242217c, 32'h409a10ef, 32'h429432c8, 32'h4234cea3};
test_output[7070] = '{32'h42b12a3b};
test_index[7070] = '{2};
test_input[56568:56575] = '{32'hc2bfd811, 32'h428e6eb6, 32'h42833dc7, 32'h42c05acd, 32'h413e6276, 32'h415327d7, 32'h42785156, 32'h42c309b8};
test_output[7071] = '{32'h42c309b8};
test_index[7071] = '{7};
test_input[56576:56583] = '{32'hc1d80293, 32'hc22c3b42, 32'hc28f41fb, 32'h42b95d77, 32'hc2638a7d, 32'hc1c23c91, 32'h4208bbf3, 32'h42080e8b};
test_output[7072] = '{32'h42b95d77};
test_index[7072] = '{3};
test_input[56584:56591] = '{32'hc1b7e704, 32'hc1bf7fe6, 32'h3f31f3b8, 32'h41975012, 32'h421b8fe5, 32'h42c5d0e5, 32'h41454a35, 32'hc2a08e22};
test_output[7073] = '{32'h42c5d0e5};
test_index[7073] = '{5};
test_input[56592:56599] = '{32'h4294520d, 32'h41fed701, 32'h42c1198e, 32'h42981b21, 32'h42b23ba8, 32'h4136cb72, 32'h42a57898, 32'h42b2e2a7};
test_output[7074] = '{32'h42c1198e};
test_index[7074] = '{2};
test_input[56600:56607] = '{32'hc2678664, 32'h42ab0a9b, 32'hc297bb0f, 32'hc23088ad, 32'hc28d1071, 32'hc233a7f9, 32'hc1c766cc, 32'hc203b500};
test_output[7075] = '{32'h42ab0a9b};
test_index[7075] = '{1};
test_input[56608:56615] = '{32'h42a5e487, 32'h4149a222, 32'h428053ae, 32'hc29192d1, 32'hc2aead86, 32'hc2b4eb04, 32'hc236ecad, 32'h42b135ba};
test_output[7076] = '{32'h42b135ba};
test_index[7076] = '{7};
test_input[56616:56623] = '{32'hc29c310d, 32'hc2b16c8b, 32'h424bb22a, 32'hc242293f, 32'hc28a9cae, 32'hc271bc85, 32'hc1a88838, 32'hc1db8bbb};
test_output[7077] = '{32'h424bb22a};
test_index[7077] = '{2};
test_input[56624:56631] = '{32'h41a566c4, 32'h41ce2b2e, 32'hc2639d57, 32'h420f6006, 32'hc151298d, 32'hc1a2b44d, 32'hc0198056, 32'h4288c840};
test_output[7078] = '{32'h4288c840};
test_index[7078] = '{7};
test_input[56632:56639] = '{32'hc1aeefcc, 32'hc208a367, 32'hc13524b9, 32'hc29319df, 32'hc2320845, 32'hc17a6d7e, 32'hc2b28865, 32'hc08f419f};
test_output[7079] = '{32'hc08f419f};
test_index[7079] = '{7};
test_input[56640:56647] = '{32'hc202ba8e, 32'h419b050c, 32'hc2ab0799, 32'hc1f2c0a1, 32'h41dc3e7d, 32'hc1fb9f45, 32'hc06aa4cf, 32'hc26058de};
test_output[7080] = '{32'h41dc3e7d};
test_index[7080] = '{4};
test_input[56648:56655] = '{32'h429eec3d, 32'h41a52e5e, 32'h42539f35, 32'h4281452d, 32'hc19a6658, 32'hc22d1695, 32'hc1af384c, 32'hc21d4b41};
test_output[7081] = '{32'h429eec3d};
test_index[7081] = '{0};
test_input[56656:56663] = '{32'hc2b5e591, 32'h428712a2, 32'h429c1823, 32'hc1563abc, 32'hc1dbe412, 32'hc2ba07c4, 32'h428cf3ec, 32'h408f95c5};
test_output[7082] = '{32'h429c1823};
test_index[7082] = '{2};
test_input[56664:56671] = '{32'h42a0313a, 32'h41d19158, 32'hc2ad51b9, 32'hc1da90be, 32'hc1d03eda, 32'h4275f921, 32'hc1297067, 32'hc2868628};
test_output[7083] = '{32'h42a0313a};
test_index[7083] = '{0};
test_input[56672:56679] = '{32'hc28abfe7, 32'hc23fe19e, 32'h423d6d32, 32'h41f2e419, 32'h42337f36, 32'hc01289d9, 32'hc2bb667b, 32'hc037efec};
test_output[7084] = '{32'h423d6d32};
test_index[7084] = '{2};
test_input[56680:56687] = '{32'h429a6d26, 32'hc2071b48, 32'hc2b19121, 32'h41341bba, 32'h42a8628f, 32'hc03f57c7, 32'hc0a64020, 32'hc1d3cc89};
test_output[7085] = '{32'h42a8628f};
test_index[7085] = '{4};
test_input[56688:56695] = '{32'h41c229a9, 32'h422297be, 32'h42afd9a8, 32'hc28cfa48, 32'h4258d33e, 32'h427bb0d7, 32'hc2a292c7, 32'hc2260213};
test_output[7086] = '{32'h42afd9a8};
test_index[7086] = '{2};
test_input[56696:56703] = '{32'hc22c2f2f, 32'h426560fb, 32'h418c512e, 32'h42a2ddcb, 32'hc2a74acc, 32'h41b6277e, 32'hc043543b, 32'hc2467abd};
test_output[7087] = '{32'h42a2ddcb};
test_index[7087] = '{3};
test_input[56704:56711] = '{32'h421af546, 32'hc292503d, 32'hc2bef696, 32'h428ff23b, 32'h42933aec, 32'h417b379a, 32'hc27875cd, 32'hc1fbd746};
test_output[7088] = '{32'h42933aec};
test_index[7088] = '{4};
test_input[56712:56719] = '{32'hc1b946ad, 32'h4240075f, 32'h410c0380, 32'hc2541d41, 32'hc155e9f7, 32'hc2adc4be, 32'hbf96ebfc, 32'h416a881d};
test_output[7089] = '{32'h4240075f};
test_index[7089] = '{1};
test_input[56720:56727] = '{32'hc281a20f, 32'h41fd605d, 32'h424701cb, 32'hc26faa15, 32'h41f55b4e, 32'hc2125a27, 32'hbfc10c48, 32'hc25a554c};
test_output[7090] = '{32'h424701cb};
test_index[7090] = '{2};
test_input[56728:56735] = '{32'h403ef329, 32'h42793a35, 32'h42a03ec3, 32'h4280d4bf, 32'hc203ebf3, 32'h3fb13b61, 32'hc2850b28, 32'hc0d1d68e};
test_output[7091] = '{32'h42a03ec3};
test_index[7091] = '{2};
test_input[56736:56743] = '{32'h420756a8, 32'h41b2d882, 32'hc2ba82fc, 32'hc296698b, 32'hc2798a0c, 32'h4191e919, 32'hc25b3441, 32'h42b8ff04};
test_output[7092] = '{32'h42b8ff04};
test_index[7092] = '{7};
test_input[56744:56751] = '{32'hc236bcc0, 32'h42a24515, 32'hc1d15d6d, 32'hc1bdd091, 32'h40cfb514, 32'hc2897223, 32'hc0e19316, 32'h42a61035};
test_output[7093] = '{32'h42a61035};
test_index[7093] = '{7};
test_input[56752:56759] = '{32'hc1f26c89, 32'hc2ab131c, 32'hc12cbf96, 32'h424802c1, 32'h418eb8a7, 32'h42c7248a, 32'h422e34b6, 32'hc2a89c55};
test_output[7094] = '{32'h42c7248a};
test_index[7094] = '{5};
test_input[56760:56767] = '{32'hc161cdbc, 32'h41a41160, 32'h41fc0f1e, 32'h4229ac21, 32'h418d0d52, 32'h41f173a0, 32'h42c07a5f, 32'h42891617};
test_output[7095] = '{32'h42c07a5f};
test_index[7095] = '{6};
test_input[56768:56775] = '{32'h41410b61, 32'hc29de5df, 32'hc23259e2, 32'hc1759d7c, 32'h40f0a672, 32'hc1a81040, 32'hc2b28a2a, 32'hc2a7c965};
test_output[7096] = '{32'h41410b61};
test_index[7096] = '{0};
test_input[56776:56783] = '{32'h42acbf5d, 32'hc2ab6da3, 32'hc2112915, 32'hc05a9631, 32'hc2bed3ed, 32'hc2ae115a, 32'h429b1e71, 32'h42580e09};
test_output[7097] = '{32'h42acbf5d};
test_index[7097] = '{0};
test_input[56784:56791] = '{32'h42a98ee6, 32'hc2b0a858, 32'h413a7990, 32'h4168de83, 32'h424d1dc5, 32'hc11a09fc, 32'hc28cc806, 32'hc2b6018a};
test_output[7098] = '{32'h42a98ee6};
test_index[7098] = '{0};
test_input[56792:56799] = '{32'h41cbe520, 32'hc28ef772, 32'h42917f06, 32'h42011103, 32'hc1b51d8a, 32'hc2bd9318, 32'hc23cfab8, 32'hc2bcb4f9};
test_output[7099] = '{32'h42917f06};
test_index[7099] = '{2};
test_input[56800:56807] = '{32'hc2c4aafb, 32'h41c45b13, 32'h418d6b80, 32'h3fba7c9e, 32'h4161f621, 32'h427298ef, 32'h42ad9d1e, 32'h4289e8b2};
test_output[7100] = '{32'h42ad9d1e};
test_index[7100] = '{6};
test_input[56808:56815] = '{32'hc2484a2d, 32'h42a4f44a, 32'hc288b8c0, 32'hc1ebb094, 32'hc2a2164a, 32'hc1912d42, 32'hc14c48bd, 32'hc10c8a3c};
test_output[7101] = '{32'h42a4f44a};
test_index[7101] = '{1};
test_input[56816:56823] = '{32'hc29255d4, 32'hc1174980, 32'hc2492005, 32'hc2adf38f, 32'hc224be5c, 32'hc242725f, 32'h429bdb76, 32'h4295b69b};
test_output[7102] = '{32'h429bdb76};
test_index[7102] = '{6};
test_input[56824:56831] = '{32'hc299163d, 32'h428ed998, 32'hc2c152d9, 32'hc29b709c, 32'hc1102eab, 32'hc15ae3b3, 32'hc0da5c43, 32'h428820bb};
test_output[7103] = '{32'h428ed998};
test_index[7103] = '{1};
test_input[56832:56839] = '{32'h42aa2e52, 32'h42c595e6, 32'hc28f84d4, 32'hc2ae3bde, 32'h4276af29, 32'hc24483ef, 32'hc2856544, 32'h412d37f5};
test_output[7104] = '{32'h42c595e6};
test_index[7104] = '{1};
test_input[56840:56847] = '{32'hc187f62e, 32'h42a67b4c, 32'hc29eae59, 32'hc1d7024f, 32'hc219c8dc, 32'h42904a20, 32'hc15c21b8, 32'h4078578f};
test_output[7105] = '{32'h42a67b4c};
test_index[7105] = '{1};
test_input[56848:56855] = '{32'h429c1b8a, 32'h40c475ef, 32'hc207a40f, 32'h425c20a0, 32'hc2355ec8, 32'h42649433, 32'h423422d1, 32'h41911104};
test_output[7106] = '{32'h429c1b8a};
test_index[7106] = '{0};
test_input[56856:56863] = '{32'h426943fa, 32'h418dec74, 32'h4253d7df, 32'hc2ab984b, 32'hc17967ae, 32'h425f13de, 32'h42018b01, 32'h41f7d8bb};
test_output[7107] = '{32'h426943fa};
test_index[7107] = '{0};
test_input[56864:56871] = '{32'hc114f123, 32'h408bba87, 32'hc2b92db2, 32'hc2773b5f, 32'hc2bcc829, 32'hc239eb45, 32'hc2bf0f0f, 32'h4298f97f};
test_output[7108] = '{32'h4298f97f};
test_index[7108] = '{7};
test_input[56872:56879] = '{32'hc0545d1d, 32'hc2c68607, 32'h41cb8bd9, 32'h421bc70d, 32'hc2c09ca5, 32'h413b2ed7, 32'h4234ab2e, 32'h415658f4};
test_output[7109] = '{32'h4234ab2e};
test_index[7109] = '{6};
test_input[56880:56887] = '{32'h41dbe58c, 32'h42ae5042, 32'hc15ebd9c, 32'h42850103, 32'hc22d8a04, 32'h42c5f526, 32'h415128f8, 32'h424112bb};
test_output[7110] = '{32'h42c5f526};
test_index[7110] = '{5};
test_input[56888:56895] = '{32'hc26ba103, 32'hc02d167f, 32'h426ae334, 32'h42917b4e, 32'hc2afa501, 32'h41877389, 32'h4214ff49, 32'h41e2b82f};
test_output[7111] = '{32'h42917b4e};
test_index[7111] = '{3};
test_input[56896:56903] = '{32'h406bb6da, 32'h42bc134f, 32'h428bd600, 32'h42a4c684, 32'hbf8d9ee7, 32'h42c61ea7, 32'hc0ab44ee, 32'h4271c353};
test_output[7112] = '{32'h42c61ea7};
test_index[7112] = '{5};
test_input[56904:56911] = '{32'hc29e9884, 32'hc242e9dd, 32'hc23261d9, 32'hc0595ea9, 32'h41df2b8f, 32'h4186d804, 32'h425394a0, 32'hc1c38131};
test_output[7113] = '{32'h425394a0};
test_index[7113] = '{6};
test_input[56912:56919] = '{32'hc2847f1c, 32'hc2a7ce9c, 32'hc1cd5a02, 32'hc06a4d5a, 32'h41131a8d, 32'h416a35f0, 32'h428fc487, 32'h40bf579a};
test_output[7114] = '{32'h428fc487};
test_index[7114] = '{6};
test_input[56920:56927] = '{32'h42c2e245, 32'h428d56c1, 32'h428898d1, 32'h425f8903, 32'hc2b9ed38, 32'hc2bf5a89, 32'h429f2cce, 32'hc2bb51e6};
test_output[7115] = '{32'h42c2e245};
test_index[7115] = '{0};
test_input[56928:56935] = '{32'h41b353fd, 32'hc2838d36, 32'hc2976624, 32'h426be241, 32'h42a489ce, 32'hc23afd56, 32'hc130c101, 32'h41d11f79};
test_output[7116] = '{32'h42a489ce};
test_index[7116] = '{4};
test_input[56936:56943] = '{32'h4278a40a, 32'hc28cb51d, 32'h425f7aae, 32'hc2affe3a, 32'h4284b0e5, 32'hc1afb87a, 32'h427344df, 32'hc2b6da47};
test_output[7117] = '{32'h4284b0e5};
test_index[7117] = '{4};
test_input[56944:56951] = '{32'hc24887ee, 32'h42585ad5, 32'h41be821e, 32'h424581a0, 32'h4153449c, 32'h41c3656a, 32'h42b584fe, 32'hc25b7371};
test_output[7118] = '{32'h42b584fe};
test_index[7118] = '{6};
test_input[56952:56959] = '{32'h42aa1a2f, 32'hc2138004, 32'hc1e81b46, 32'h4266cbc2, 32'hc244fdba, 32'hc26d7294, 32'h42bc94ab, 32'h42178339};
test_output[7119] = '{32'h42bc94ab};
test_index[7119] = '{6};
test_input[56960:56967] = '{32'hc0c4707c, 32'h42691e93, 32'hc283c39b, 32'hc1bdb318, 32'h414cde08, 32'hc28cd78e, 32'hc27a8e29, 32'h42330752};
test_output[7120] = '{32'h42691e93};
test_index[7120] = '{1};
test_input[56968:56975] = '{32'h41e27f45, 32'h42318224, 32'hc278af84, 32'h422cebc3, 32'h42917411, 32'h425b5c33, 32'hc28786d6, 32'hc1e7d64b};
test_output[7121] = '{32'h42917411};
test_index[7121] = '{4};
test_input[56976:56983] = '{32'h425387b7, 32'h411df036, 32'hc23bb3f8, 32'h426f8268, 32'h42c5a7aa, 32'hc273c563, 32'h41b12ecc, 32'h42af68dd};
test_output[7122] = '{32'h42c5a7aa};
test_index[7122] = '{4};
test_input[56984:56991] = '{32'hc286a12a, 32'h42629c51, 32'h421c0be8, 32'hc2857ccd, 32'h429629df, 32'hc28bb233, 32'hc2266506, 32'h42948db5};
test_output[7123] = '{32'h429629df};
test_index[7123] = '{4};
test_input[56992:56999] = '{32'hc20babfb, 32'h42544ccd, 32'h427c0518, 32'hc2619a8a, 32'hc2af8053, 32'hc23f8e37, 32'hc277dbe0, 32'hc2a4dd66};
test_output[7124] = '{32'h427c0518};
test_index[7124] = '{2};
test_input[57000:57007] = '{32'hc2b70da1, 32'h41cae696, 32'hc0a5cff5, 32'hc2777e57, 32'hc2a3b7da, 32'hc1ae8836, 32'h42303d7c, 32'h41909b75};
test_output[7125] = '{32'h42303d7c};
test_index[7125] = '{6};
test_input[57008:57015] = '{32'hc2566649, 32'h42870d2a, 32'hc28a4cf9, 32'hc1e2b699, 32'hc29bcad7, 32'h408e07ef, 32'h4137dfcf, 32'h419ed824};
test_output[7126] = '{32'h42870d2a};
test_index[7126] = '{1};
test_input[57016:57023] = '{32'h4231363b, 32'hc29b2838, 32'hc28ca938, 32'hc2a92caf, 32'h425e7a85, 32'hc257fbab, 32'h428418fc, 32'h41b7c31a};
test_output[7127] = '{32'h428418fc};
test_index[7127] = '{6};
test_input[57024:57031] = '{32'hc23cc4c7, 32'hc2b450ce, 32'hc10def74, 32'h42b339ad, 32'h426ea370, 32'hc1b3159c, 32'hc14851b2, 32'h3f679367};
test_output[7128] = '{32'h42b339ad};
test_index[7128] = '{3};
test_input[57032:57039] = '{32'hc2a3a75c, 32'h42ae938c, 32'hc26ad0c0, 32'h410501f8, 32'h4294dcab, 32'h417d0b0e, 32'h4271f9fa, 32'hc2570fe7};
test_output[7129] = '{32'h42ae938c};
test_index[7129] = '{1};
test_input[57040:57047] = '{32'h42458472, 32'hc29958c8, 32'h42bedf9d, 32'h419aba39, 32'h424b3efb, 32'hc295037c, 32'hc2082375, 32'hc25d5038};
test_output[7130] = '{32'h42bedf9d};
test_index[7130] = '{2};
test_input[57048:57055] = '{32'hc21c5d93, 32'h42891d4e, 32'hc0ef9a9a, 32'hc22a990a, 32'h4093e156, 32'h422f283f, 32'h42982dda, 32'h420f04aa};
test_output[7131] = '{32'h42982dda};
test_index[7131] = '{6};
test_input[57056:57063] = '{32'h407c5f09, 32'hc291437c, 32'h40a63a75, 32'hc1b31733, 32'hc286e026, 32'h41beb566, 32'hc2868e95, 32'hc237a214};
test_output[7132] = '{32'h41beb566};
test_index[7132] = '{5};
test_input[57064:57071] = '{32'hc2a20f65, 32'h42a78238, 32'h423cc6ee, 32'h42bc00a5, 32'h4262cf2b, 32'hc0dbacbc, 32'h4138dddc, 32'h4135112a};
test_output[7133] = '{32'h42bc00a5};
test_index[7133] = '{3};
test_input[57072:57079] = '{32'hc01bf46d, 32'h41922a7b, 32'hc080d2d0, 32'hc1f75e96, 32'h42101256, 32'hc215fe3c, 32'h42b56e31, 32'hc27543ad};
test_output[7134] = '{32'h42b56e31};
test_index[7134] = '{6};
test_input[57080:57087] = '{32'hc22f2ae1, 32'hc208d8ad, 32'h4278707f, 32'h40e632b7, 32'hc27171dd, 32'h414f49cb, 32'h42442d55, 32'h4239b6e6};
test_output[7135] = '{32'h4278707f};
test_index[7135] = '{2};
test_input[57088:57095] = '{32'hc2bc3cb1, 32'hc2563177, 32'hc2a13da4, 32'h41a47702, 32'hc1795138, 32'hc2861130, 32'hc2c6ecf8, 32'hc292a164};
test_output[7136] = '{32'h41a47702};
test_index[7136] = '{3};
test_input[57096:57103] = '{32'h40eb4a17, 32'hc1e855ce, 32'hc28f6537, 32'h41ab2f98, 32'h42743117, 32'h42b2bb94, 32'hc2606e0f, 32'h41b67dd2};
test_output[7137] = '{32'h42b2bb94};
test_index[7137] = '{5};
test_input[57104:57111] = '{32'hc1d51be8, 32'hc1e8f4f2, 32'h42796ca4, 32'h426b4b37, 32'h420fe47d, 32'h42825d70, 32'h423292e7, 32'hc29ba56b};
test_output[7138] = '{32'h42825d70};
test_index[7138] = '{5};
test_input[57112:57119] = '{32'h42422aaf, 32'h423f4024, 32'h423b84a2, 32'h429849e5, 32'hc27d3764, 32'hc28d8d86, 32'hc2af8d1f, 32'hc28bf785};
test_output[7139] = '{32'h429849e5};
test_index[7139] = '{3};
test_input[57120:57127] = '{32'hc1d0f0da, 32'h4214abc0, 32'h42b2f4df, 32'h4251ea44, 32'hc1eb267c, 32'hc26453c4, 32'h407bc60c, 32'hc03b7fb5};
test_output[7140] = '{32'h42b2f4df};
test_index[7140] = '{2};
test_input[57128:57135] = '{32'hc1d85acc, 32'hc21b0c60, 32'hc282400d, 32'hc1d51ba3, 32'hc25f59f2, 32'hc2a31d38, 32'h414c0ea9, 32'h42b132c7};
test_output[7141] = '{32'h42b132c7};
test_index[7141] = '{7};
test_input[57136:57143] = '{32'h427e4f7a, 32'h42177697, 32'hc14637e2, 32'h41ed64c1, 32'hc13b3a2a, 32'hc181d7ce, 32'h4294d9e2, 32'hc2b846db};
test_output[7142] = '{32'h4294d9e2};
test_index[7142] = '{6};
test_input[57144:57151] = '{32'h429b2ed4, 32'hc221a3db, 32'hc2c49cb0, 32'h41b0bc93, 32'hc091e6eb, 32'h40878208, 32'h429a0516, 32'hc27c91da};
test_output[7143] = '{32'h429b2ed4};
test_index[7143] = '{0};
test_input[57152:57159] = '{32'hc1c3d0b5, 32'hc16487c8, 32'hc226cb1d, 32'h421b3d1d, 32'hc2896667, 32'h42be91f4, 32'h4241b8e5, 32'h41066569};
test_output[7144] = '{32'h42be91f4};
test_index[7144] = '{5};
test_input[57160:57167] = '{32'h3d36dfaf, 32'hc21ffaf2, 32'hc2688230, 32'h42b9c13b, 32'hc0313ef2, 32'hc1e7c51b, 32'hc2522548, 32'hc2557033};
test_output[7145] = '{32'h42b9c13b};
test_index[7145] = '{3};
test_input[57168:57175] = '{32'hc24cc2ef, 32'h408fe5bd, 32'hc1982795, 32'h423d3dbe, 32'h4156c986, 32'h428e1809, 32'hc230df57, 32'hc26aeb12};
test_output[7146] = '{32'h428e1809};
test_index[7146] = '{5};
test_input[57176:57183] = '{32'hc2b91873, 32'h42568eb1, 32'h41885234, 32'hc2791fa8, 32'h41c00702, 32'h4096ba55, 32'hc27726a0, 32'hc190a19b};
test_output[7147] = '{32'h42568eb1};
test_index[7147] = '{1};
test_input[57184:57191] = '{32'hc22d4752, 32'hc2ba4a25, 32'hc1f3bda8, 32'hc2938130, 32'h4282aa05, 32'h42839f75, 32'hc203d120, 32'h428380a9};
test_output[7148] = '{32'h42839f75};
test_index[7148] = '{5};
test_input[57192:57199] = '{32'hc2beb0e4, 32'hbd3c201f, 32'h42a461ae, 32'h4249c6c1, 32'hc2a17891, 32'h4141409c, 32'hc2aa079f, 32'h41079f18};
test_output[7149] = '{32'h42a461ae};
test_index[7149] = '{2};
test_input[57200:57207] = '{32'h428b772f, 32'h424ac72d, 32'h4287d005, 32'h4297a424, 32'hc203e1c3, 32'hc1d3a814, 32'hc1ff3f18, 32'hc2c51f0f};
test_output[7150] = '{32'h4297a424};
test_index[7150] = '{3};
test_input[57208:57215] = '{32'h42b47d71, 32'hbfa68ba5, 32'hc204544a, 32'h40c16aa7, 32'hc2bc9667, 32'h422f9ec0, 32'h41eaac46, 32'h411dfb72};
test_output[7151] = '{32'h42b47d71};
test_index[7151] = '{0};
test_input[57216:57223] = '{32'h42b300be, 32'hc21f0a4d, 32'hc1b60e74, 32'h429cc9ab, 32'h41224332, 32'hc1bd2142, 32'h4254b2ca, 32'h426e310d};
test_output[7152] = '{32'h42b300be};
test_index[7152] = '{0};
test_input[57224:57231] = '{32'h416e4072, 32'h425c6c31, 32'hc2a53c64, 32'hc0264b97, 32'h42074564, 32'hc2a024a3, 32'h414baa81, 32'hc2a530e3};
test_output[7153] = '{32'h425c6c31};
test_index[7153] = '{1};
test_input[57232:57239] = '{32'h418480e7, 32'hc21b585a, 32'hc29887d2, 32'hc2938c2e, 32'hc1ca7c4a, 32'h42a7f809, 32'h410342b7, 32'h42a5b37c};
test_output[7154] = '{32'h42a7f809};
test_index[7154] = '{5};
test_input[57240:57247] = '{32'h42574426, 32'hc280c0f4, 32'hc18d47eb, 32'h42042c14, 32'h42c2f9b9, 32'hc26c485f, 32'h4296af6a, 32'h42237d32};
test_output[7155] = '{32'h42c2f9b9};
test_index[7155] = '{4};
test_input[57248:57255] = '{32'hc16e309b, 32'hc28725fd, 32'h4241bfa4, 32'h41d56a2c, 32'hc163ee6b, 32'h42b79575, 32'h429ba051, 32'h4209ffc2};
test_output[7156] = '{32'h42b79575};
test_index[7156] = '{5};
test_input[57256:57263] = '{32'hc1102f2c, 32'h42a6d4bf, 32'hc23d8ee2, 32'hc1610565, 32'hc1d36432, 32'h42b37a24, 32'h413e3e9d, 32'h4294e4a4};
test_output[7157] = '{32'h42b37a24};
test_index[7157] = '{5};
test_input[57264:57271] = '{32'hc21b49c6, 32'h422af155, 32'hc2959f98, 32'h42a7a5bc, 32'h4246619d, 32'h4281bdbd, 32'hc2a55f0e, 32'hc26e6366};
test_output[7158] = '{32'h42a7a5bc};
test_index[7158] = '{3};
test_input[57272:57279] = '{32'hc143161b, 32'h4221c2e1, 32'hc23c4cc5, 32'h40ae921b, 32'h42b48867, 32'hc22eec6d, 32'h421fc2d3, 32'hc2b2c0a0};
test_output[7159] = '{32'h42b48867};
test_index[7159] = '{4};
test_input[57280:57287] = '{32'h42b365b0, 32'h41e565bb, 32'h411b7b16, 32'h4210e0f6, 32'h42672d54, 32'h42b02c6c, 32'hc1b97e9a, 32'h4148c4ad};
test_output[7160] = '{32'h42b365b0};
test_index[7160] = '{0};
test_input[57288:57295] = '{32'hc19913a3, 32'h428b8851, 32'h42ace251, 32'hc2570e86, 32'h419a8c2a, 32'h428a35eb, 32'h426ff4a7, 32'h421955cf};
test_output[7161] = '{32'h42ace251};
test_index[7161] = '{2};
test_input[57296:57303] = '{32'hc263013c, 32'hc22dd490, 32'h422fe4a3, 32'hc2652012, 32'hc2c5e82b, 32'h426e47c2, 32'hc29ce74f, 32'h426e7879};
test_output[7162] = '{32'h426e7879};
test_index[7162] = '{7};
test_input[57304:57311] = '{32'h4212d5c2, 32'hc28d4c07, 32'h426662ce, 32'hc280ffca, 32'hc2b13774, 32'h42747498, 32'h423fb8d2, 32'h428c7c1d};
test_output[7163] = '{32'h428c7c1d};
test_index[7163] = '{7};
test_input[57312:57319] = '{32'hc189bafb, 32'hc2bd72df, 32'hc2976371, 32'h428cc665, 32'hc0ffcc34, 32'hc28cb20b, 32'hc13ac602, 32'h4230507d};
test_output[7164] = '{32'h428cc665};
test_index[7164] = '{3};
test_input[57320:57327] = '{32'h421d7e68, 32'hc27e298e, 32'h427a3b41, 32'hc2661ad1, 32'hc275f272, 32'h40b28075, 32'h4205af1b, 32'h41b83759};
test_output[7165] = '{32'h427a3b41};
test_index[7165] = '{2};
test_input[57328:57335] = '{32'hc29b9c13, 32'hc28c40e4, 32'h429f6155, 32'h41b18640, 32'hc2c70105, 32'hc238d492, 32'h42b5322c, 32'h4256f7e4};
test_output[7166] = '{32'h42b5322c};
test_index[7166] = '{6};
test_input[57336:57343] = '{32'hc20fe4ad, 32'h42c47ec2, 32'h41e20e48, 32'h420b6e28, 32'hc2a97a06, 32'hc1ef6021, 32'hc2b9735a, 32'h41a66a2a};
test_output[7167] = '{32'h42c47ec2};
test_index[7167] = '{1};
test_input[57344:57351] = '{32'h429dc0ef, 32'h42a9496e, 32'h42520b79, 32'hc23ba27b, 32'hc09d82c5, 32'hc0b09f35, 32'hc27fda6a, 32'hc256ab3b};
test_output[7168] = '{32'h42a9496e};
test_index[7168] = '{1};
test_input[57352:57359] = '{32'hc00483ec, 32'hc17cf9fa, 32'h41407e37, 32'hc20ba242, 32'hc2861939, 32'h411be150, 32'h4143496e, 32'hc230c786};
test_output[7169] = '{32'h4143496e};
test_index[7169] = '{6};
test_input[57360:57367] = '{32'hc2b37501, 32'hc2b01be3, 32'hc1a60cfe, 32'hc296e982, 32'hc2a796d7, 32'h42b1bbf2, 32'hc2af0922, 32'h4218e458};
test_output[7170] = '{32'h42b1bbf2};
test_index[7170] = '{5};
test_input[57368:57375] = '{32'hc2444332, 32'hc2b07a48, 32'h4230bcf9, 32'h41f5bfa5, 32'h428541f5, 32'hc073994a, 32'h4286d3bb, 32'hc1472fcb};
test_output[7171] = '{32'h4286d3bb};
test_index[7171] = '{6};
test_input[57376:57383] = '{32'hc2b2eff2, 32'hc28f2774, 32'hc0ed85c1, 32'h41ee74ab, 32'h429624b3, 32'h42afd42e, 32'h42b90ec6, 32'hc29fc2ca};
test_output[7172] = '{32'h42b90ec6};
test_index[7172] = '{6};
test_input[57384:57391] = '{32'h41a7f1f2, 32'hc2abea12, 32'h41c648fe, 32'h4202cf39, 32'hc1b03b36, 32'h4017d52e, 32'h4260bb76, 32'h41537d8a};
test_output[7173] = '{32'h4260bb76};
test_index[7173] = '{6};
test_input[57392:57399] = '{32'h41dabef0, 32'h42aaf0d7, 32'hc1adb795, 32'h42aa786b, 32'h4015387c, 32'hc29ddced, 32'h418c48aa, 32'hc262b231};
test_output[7174] = '{32'h42aaf0d7};
test_index[7174] = '{1};
test_input[57400:57407] = '{32'hc20459d4, 32'h425fe394, 32'h419d894f, 32'h4189ecb3, 32'h42c46b0a, 32'hc26d32bc, 32'h426faf44, 32'hc29deb9d};
test_output[7175] = '{32'h42c46b0a};
test_index[7175] = '{4};
test_input[57408:57415] = '{32'hc24d2d74, 32'h42415113, 32'h40619779, 32'hc20b2117, 32'h4225c60e, 32'h42ad5d15, 32'hc2207ced, 32'h4253ed8c};
test_output[7176] = '{32'h42ad5d15};
test_index[7176] = '{5};
test_input[57416:57423] = '{32'h42818a94, 32'h42789f6f, 32'h42081472, 32'h429bb1c7, 32'hc2771a14, 32'hc28db467, 32'h425468ba, 32'hc2a2ed15};
test_output[7177] = '{32'h429bb1c7};
test_index[7177] = '{3};
test_input[57424:57431] = '{32'h425dfcc4, 32'hc23980ab, 32'h421e34f0, 32'h4186f8ca, 32'hc25377b5, 32'hc2bc84e0, 32'hc0364e27, 32'hc2683743};
test_output[7178] = '{32'h425dfcc4};
test_index[7178] = '{0};
test_input[57432:57439] = '{32'hc1edab49, 32'hc10cf789, 32'hc2b20b63, 32'h4289ce25, 32'h4298b813, 32'hc2159fc0, 32'hc05c95bf, 32'h411c83bb};
test_output[7179] = '{32'h4298b813};
test_index[7179] = '{4};
test_input[57440:57447] = '{32'h4233135d, 32'hc23cdbc0, 32'h42110e91, 32'h424990ff, 32'h426f56ec, 32'h41ffe4b0, 32'hc2500fac, 32'h42266e0b};
test_output[7180] = '{32'h426f56ec};
test_index[7180] = '{4};
test_input[57448:57455] = '{32'h42b55b4d, 32'hc2a01388, 32'hc27359ca, 32'h42a99b05, 32'hc1d8465d, 32'hc1c54de2, 32'h42b9445f, 32'hc06e36ff};
test_output[7181] = '{32'h42b9445f};
test_index[7181] = '{6};
test_input[57456:57463] = '{32'hc10c0164, 32'hc26815db, 32'h42420c1f, 32'h418bc59f, 32'h419bc804, 32'h4170aa0b, 32'hc291f5c1, 32'hc2c22b9b};
test_output[7182] = '{32'h42420c1f};
test_index[7182] = '{2};
test_input[57464:57471] = '{32'hc28b63a3, 32'h420f273e, 32'h4191e2a1, 32'hc267fe7d, 32'hc1c56e4d, 32'h4218e9f2, 32'h4233da2f, 32'hc28b2fe5};
test_output[7183] = '{32'h4233da2f};
test_index[7183] = '{6};
test_input[57472:57479] = '{32'hc05063ec, 32'h425bcab8, 32'hc110036a, 32'h421d386f, 32'hc18f9879, 32'hc2862215, 32'hc2ab0630, 32'hc269365c};
test_output[7184] = '{32'h425bcab8};
test_index[7184] = '{1};
test_input[57480:57487] = '{32'hc22466d7, 32'hc2b78175, 32'hc2743212, 32'hc2318d94, 32'h42a8cbaf, 32'h4281f1a2, 32'h42335255, 32'h42746baa};
test_output[7185] = '{32'h42a8cbaf};
test_index[7185] = '{4};
test_input[57488:57495] = '{32'h428ea951, 32'h420f5bfa, 32'hc26f0915, 32'h428a8713, 32'h41151636, 32'hc28299cf, 32'hc2c702fe, 32'hc2b43607};
test_output[7186] = '{32'h428ea951};
test_index[7186] = '{0};
test_input[57496:57503] = '{32'h420da7ec, 32'hc2c48b39, 32'hc2bd0c85, 32'h42101226, 32'h4295649a, 32'hc257c104, 32'hc1764fc5, 32'hc2468093};
test_output[7187] = '{32'h4295649a};
test_index[7187] = '{4};
test_input[57504:57511] = '{32'h42752e95, 32'h428eecd9, 32'h41266ea0, 32'h42630d10, 32'h4184e797, 32'hc02468c5, 32'hc256aaca, 32'h42af5e47};
test_output[7188] = '{32'h42af5e47};
test_index[7188] = '{7};
test_input[57512:57519] = '{32'h425a4529, 32'hc127b1bf, 32'hc26788cf, 32'h40935e30, 32'hc1d20d97, 32'hc07ccf6b, 32'h42b9f5ca, 32'hc2c6a1e2};
test_output[7189] = '{32'h42b9f5ca};
test_index[7189] = '{6};
test_input[57520:57527] = '{32'hc231e179, 32'h4258c837, 32'h4247e691, 32'h418b6bd7, 32'hc2c73a62, 32'h429dd637, 32'hc142d852, 32'hc294a3dc};
test_output[7190] = '{32'h429dd637};
test_index[7190] = '{5};
test_input[57528:57535] = '{32'hc2b4aed2, 32'h40b08dac, 32'hc2c1bc1a, 32'hc2b6c168, 32'h429d905f, 32'hc0f87672, 32'h4265c512, 32'h421110fe};
test_output[7191] = '{32'h429d905f};
test_index[7191] = '{4};
test_input[57536:57543] = '{32'hc28aa7bd, 32'h42be961f, 32'h421b1b5c, 32'hc2492c06, 32'h428e51cc, 32'hc2106472, 32'hc21e36a9, 32'h41bb8451};
test_output[7192] = '{32'h42be961f};
test_index[7192] = '{1};
test_input[57544:57551] = '{32'h4294235d, 32'hc250344e, 32'h422c1f10, 32'h423cfb1e, 32'hc1ae6eba, 32'hc043c91d, 32'h416860be, 32'hc28ee901};
test_output[7193] = '{32'h4294235d};
test_index[7193] = '{0};
test_input[57552:57559] = '{32'h421aff65, 32'h42c230fa, 32'h429d4fed, 32'hc2b2c722, 32'h420b3ee9, 32'h42c7730b, 32'hbfcdafa0, 32'hc2bfe864};
test_output[7194] = '{32'h42c7730b};
test_index[7194] = '{5};
test_input[57560:57567] = '{32'hc2b58aa2, 32'h42a17dbf, 32'hc1addea3, 32'hc2ad42ee, 32'hc28190da, 32'hc2bc2feb, 32'hc23f4241, 32'hc2405f45};
test_output[7195] = '{32'h42a17dbf};
test_index[7195] = '{1};
test_input[57568:57575] = '{32'h41d0275f, 32'hc25021c2, 32'h41a633d8, 32'hc0715980, 32'hc2adbcd1, 32'h41cc2ece, 32'hc296cef8, 32'hbff840dd};
test_output[7196] = '{32'h41d0275f};
test_index[7196] = '{0};
test_input[57576:57583] = '{32'h42a0e02e, 32'h4173690f, 32'h40f80d3c, 32'hc2bf920f, 32'h42077765, 32'h426fb2c0, 32'h4219f21a, 32'hc2b4b073};
test_output[7197] = '{32'h42a0e02e};
test_index[7197] = '{0};
test_input[57584:57591] = '{32'hc20b5631, 32'hc27692b1, 32'h4260956d, 32'h423fdf07, 32'h4147f96d, 32'hc1f546bd, 32'h42c72b69, 32'hc23dc611};
test_output[7198] = '{32'h42c72b69};
test_index[7198] = '{6};
test_input[57592:57599] = '{32'hc2408a79, 32'hc0ebdb4f, 32'h422aa94a, 32'hc20feb07, 32'hc1fdf751, 32'h42c7bba3, 32'hc2804449, 32'hc2b718c4};
test_output[7199] = '{32'h42c7bba3};
test_index[7199] = '{5};
test_input[57600:57607] = '{32'hc2aee2cc, 32'hc24a0dd5, 32'h42a2fb5d, 32'hc2c07566, 32'hc08b22fb, 32'h42285a2d, 32'hc2c1f749, 32'hc2802124};
test_output[7200] = '{32'h42a2fb5d};
test_index[7200] = '{2};
test_input[57608:57615] = '{32'hc2b863c9, 32'h425e8e5a, 32'h424953b2, 32'hc2b68807, 32'h424197d8, 32'h42859c33, 32'h42088ce1, 32'h42b3861a};
test_output[7201] = '{32'h42b3861a};
test_index[7201] = '{7};
test_input[57616:57623] = '{32'h428352dc, 32'hc2c34cff, 32'h42a413d8, 32'h4280e779, 32'h42694191, 32'hc292065a, 32'hc28eefa1, 32'hc27fc453};
test_output[7202] = '{32'h42a413d8};
test_index[7202] = '{2};
test_input[57624:57631] = '{32'hc2a2c2be, 32'h41504ab2, 32'hc13f9566, 32'hc203944e, 32'hc21cdc21, 32'h421832cf, 32'h42957ac0, 32'hbfe0b08b};
test_output[7203] = '{32'h42957ac0};
test_index[7203] = '{6};
test_input[57632:57639] = '{32'hc203c54c, 32'hc22146d3, 32'h412953aa, 32'h41fab09e, 32'h40494650, 32'hc21624a1, 32'hc201cd4d, 32'h428397cc};
test_output[7204] = '{32'h428397cc};
test_index[7204] = '{7};
test_input[57640:57647] = '{32'h42969aff, 32'hc239146d, 32'h41ae51eb, 32'h41b6aae3, 32'h41cf4f13, 32'h414f249b, 32'hc1969abf, 32'hc29d9f5b};
test_output[7205] = '{32'h42969aff};
test_index[7205] = '{0};
test_input[57648:57655] = '{32'hc2b739b5, 32'hc198e4f6, 32'h4118590a, 32'h42a6cacd, 32'h42b43186, 32'hc23ed09e, 32'h41f6caec, 32'hc2325253};
test_output[7206] = '{32'h42b43186};
test_index[7206] = '{4};
test_input[57656:57663] = '{32'h42286887, 32'h41d3b1d4, 32'hc228b427, 32'h42aef1a9, 32'h42b8af4e, 32'hc21c1a54, 32'h4286ed31, 32'h4154d583};
test_output[7207] = '{32'h42b8af4e};
test_index[7207] = '{4};
test_input[57664:57671] = '{32'h42bcbc7e, 32'hc1f527b1, 32'hc219000b, 32'hc2961f54, 32'hc2b7d4dd, 32'hc29ca04e, 32'h42073183, 32'hc1043d81};
test_output[7208] = '{32'h42bcbc7e};
test_index[7208] = '{0};
test_input[57672:57679] = '{32'h42acfa74, 32'hc2408f98, 32'h426f6229, 32'hc282a019, 32'h42860769, 32'h4230ba5a, 32'hc1caa427, 32'hc220d8e1};
test_output[7209] = '{32'h42acfa74};
test_index[7209] = '{0};
test_input[57680:57687] = '{32'hc28748db, 32'hc19876ab, 32'hc2b8c1fe, 32'hc250ef63, 32'h42830688, 32'h419350ef, 32'h41c21d7c, 32'h41050309};
test_output[7210] = '{32'h42830688};
test_index[7210] = '{4};
test_input[57688:57695] = '{32'h42b3041e, 32'hc28f2099, 32'h41a3e4fd, 32'hc1808174, 32'hc0bbf665, 32'h422af09d, 32'h4228ec84, 32'h41608211};
test_output[7211] = '{32'h42b3041e};
test_index[7211] = '{0};
test_input[57696:57703] = '{32'hc1ba8f75, 32'hc2a9a564, 32'h423e0c62, 32'h41bc52b5, 32'h42b14e98, 32'h421f0b31, 32'hc2349bf7, 32'h42122b54};
test_output[7212] = '{32'h42b14e98};
test_index[7212] = '{4};
test_input[57704:57711] = '{32'hc0e5a2ca, 32'hc1e9cf53, 32'hc2341cd7, 32'h428608e2, 32'h4282f9c5, 32'h3f7b4804, 32'h41db7f1b, 32'hc2b309e9};
test_output[7213] = '{32'h428608e2};
test_index[7213] = '{3};
test_input[57712:57719] = '{32'h420eb667, 32'h41e990ec, 32'hc298c477, 32'h42a5fbd3, 32'h41e593ae, 32'h4139beb5, 32'h4063cb54, 32'h42848972};
test_output[7214] = '{32'h42a5fbd3};
test_index[7214] = '{3};
test_input[57720:57727] = '{32'hc26d99f2, 32'h41a3969e, 32'h41c87204, 32'hc29af886, 32'h422b80bd, 32'h429e645d, 32'h41915930, 32'h41c3e039};
test_output[7215] = '{32'h429e645d};
test_index[7215] = '{5};
test_input[57728:57735] = '{32'hc239ef8a, 32'h41906959, 32'h428f6571, 32'hc23dfcb7, 32'hc2a7f61e, 32'hbd5021ce, 32'h42ac8d51, 32'h428cb1b9};
test_output[7216] = '{32'h42ac8d51};
test_index[7216] = '{6};
test_input[57736:57743] = '{32'hc1670628, 32'h42c44307, 32'hc2c24ef7, 32'hc2949155, 32'h416c2b65, 32'hc2be2921, 32'hc18097f5, 32'h429ee85b};
test_output[7217] = '{32'h42c44307};
test_index[7217] = '{1};
test_input[57744:57751] = '{32'hc2a928f6, 32'hbfabdb3e, 32'h41463486, 32'h4269c7a0, 32'h41b992f3, 32'hc1f700df, 32'h421da280, 32'hc19f9226};
test_output[7218] = '{32'h4269c7a0};
test_index[7218] = '{3};
test_input[57752:57759] = '{32'hc2adcb4b, 32'hc2c23cc4, 32'hc1100cf8, 32'h406cd1f0, 32'hc25d42ea, 32'hc18b50a9, 32'h427dfa7a, 32'hc13782be};
test_output[7219] = '{32'h427dfa7a};
test_index[7219] = '{6};
test_input[57760:57767] = '{32'hc0f3eff2, 32'h4249c1f4, 32'hc0c530ff, 32'h42770250, 32'h4298e65e, 32'h4256dd46, 32'hc2b0f5a2, 32'hc22ff456};
test_output[7220] = '{32'h4298e65e};
test_index[7220] = '{4};
test_input[57768:57775] = '{32'hc2550804, 32'h420ce651, 32'h40ba5135, 32'h4214ca2e, 32'h4202524b, 32'hc187383a, 32'hc2bc7d28, 32'h42b4b436};
test_output[7221] = '{32'h42b4b436};
test_index[7221] = '{7};
test_input[57776:57783] = '{32'hc09b301b, 32'h427e3567, 32'hc2991b8e, 32'h428a9cb1, 32'hc23f0076, 32'h40e4382e, 32'hc229a7a9, 32'h41293f66};
test_output[7222] = '{32'h428a9cb1};
test_index[7222] = '{3};
test_input[57784:57791] = '{32'hc132cfd2, 32'h42be3c9f, 32'hc28171cb, 32'h41e61a32, 32'hc18ba389, 32'h425ab138, 32'hc2b4e805, 32'h422c2208};
test_output[7223] = '{32'h42be3c9f};
test_index[7223] = '{1};
test_input[57792:57799] = '{32'hc2c5d5f3, 32'h4288d18c, 32'h42b31ceb, 32'h412ea919, 32'hc19622ae, 32'h41b2b96a, 32'h422d9477, 32'hc27cbc03};
test_output[7224] = '{32'h42b31ceb};
test_index[7224] = '{2};
test_input[57800:57807] = '{32'hc20f5652, 32'h41dee40b, 32'hc1919467, 32'hc2349fc4, 32'hc203b4cc, 32'h4299680b, 32'hbf10a005, 32'h41ff5b72};
test_output[7225] = '{32'h4299680b};
test_index[7225] = '{5};
test_input[57808:57815] = '{32'h4290b503, 32'hc1d26322, 32'hc18c653f, 32'h4208f498, 32'hc234e271, 32'h429b033b, 32'h41bc86aa, 32'h3dd0eff2};
test_output[7226] = '{32'h429b033b};
test_index[7226] = '{5};
test_input[57816:57823] = '{32'hc2969637, 32'h401541d1, 32'h42666c22, 32'h42151cc0, 32'h419944ab, 32'hc16f0d03, 32'h428d9f11, 32'h426b505b};
test_output[7227] = '{32'h428d9f11};
test_index[7227] = '{6};
test_input[57824:57831] = '{32'hc193ff93, 32'h41c79158, 32'hc29fdd48, 32'h42a4486e, 32'h4293a71f, 32'hc2896f2f, 32'hc27f47ac, 32'h426d5a0f};
test_output[7228] = '{32'h42a4486e};
test_index[7228] = '{3};
test_input[57832:57839] = '{32'hc2c72d99, 32'h402ea1ca, 32'h426e2b27, 32'h42b4186f, 32'hc2b4c090, 32'h42b9bdf3, 32'h42a64af7, 32'hc130bfc0};
test_output[7229] = '{32'h42b9bdf3};
test_index[7229] = '{5};
test_input[57840:57847] = '{32'hc214c5aa, 32'h42bab4f1, 32'h42c71cf6, 32'h42ae956b, 32'hc0b47a7a, 32'hc1b88216, 32'h4242b95e, 32'hc16e70d3};
test_output[7230] = '{32'h42c71cf6};
test_index[7230] = '{2};
test_input[57848:57855] = '{32'hc27dffd6, 32'hc14d1a97, 32'h426b6613, 32'hbf4baa10, 32'h4227b2d6, 32'h427a8d0c, 32'hc2a3a33b, 32'hc1ad9e7a};
test_output[7231] = '{32'h427a8d0c};
test_index[7231] = '{5};
test_input[57856:57863] = '{32'h3eb8e727, 32'hc1f5162d, 32'hc189d325, 32'hc2ae125a, 32'h41788368, 32'hc206ecc4, 32'h42473dba, 32'hc260a2ba};
test_output[7232] = '{32'h42473dba};
test_index[7232] = '{6};
test_input[57864:57871] = '{32'hc0baa1cc, 32'h42943dd9, 32'h4249fcb7, 32'hc23c153a, 32'h412ad6a6, 32'h421cd03c, 32'hc22b4a02, 32'hc101f7c7};
test_output[7233] = '{32'h42943dd9};
test_index[7233] = '{1};
test_input[57872:57879] = '{32'h4295c7db, 32'h42c6153c, 32'hc29adfaf, 32'hc28a883b, 32'h42c32782, 32'hc2919776, 32'hc247b7ba, 32'h41e535bd};
test_output[7234] = '{32'h42c6153c};
test_index[7234] = '{1};
test_input[57880:57887] = '{32'hc22cbe9d, 32'h42b4fe37, 32'hc22201ff, 32'h422d2ba1, 32'h40965db9, 32'h42252da1, 32'hc2683a75, 32'h4120f273};
test_output[7235] = '{32'h42b4fe37};
test_index[7235] = '{1};
test_input[57888:57895] = '{32'h428a6632, 32'h4056e45a, 32'hc1fc9fec, 32'hc2a69512, 32'h429e5f50, 32'h4284b757, 32'h415fe0cb, 32'hc1704c1a};
test_output[7236] = '{32'h429e5f50};
test_index[7236] = '{4};
test_input[57896:57903] = '{32'h42aadd5d, 32'h42af1fab, 32'hc2ad25c6, 32'hc297b284, 32'hc22a7446, 32'h400dd64f, 32'hc1f463f5, 32'h428d3cd5};
test_output[7237] = '{32'h42af1fab};
test_index[7237] = '{1};
test_input[57904:57911] = '{32'hc20898e0, 32'h42a597bc, 32'hc281be29, 32'h4257715f, 32'h40d75247, 32'h42933249, 32'hc1427ea5, 32'h427269ed};
test_output[7238] = '{32'h42a597bc};
test_index[7238] = '{1};
test_input[57912:57919] = '{32'h426514c5, 32'hc20ce316, 32'hc1fcf9f7, 32'h42a19f32, 32'hbecd0192, 32'h4280032a, 32'h40c4b073, 32'hc2781585};
test_output[7239] = '{32'h42a19f32};
test_index[7239] = '{3};
test_input[57920:57927] = '{32'h42910248, 32'h42bb120d, 32'h41f96517, 32'hc26d7d84, 32'hc2be9099, 32'h42a2aa13, 32'hc2ac8610, 32'hc23c2785};
test_output[7240] = '{32'h42bb120d};
test_index[7240] = '{1};
test_input[57928:57935] = '{32'h42c4b943, 32'hc238f007, 32'hc2b64bb1, 32'hc2a6cc8a, 32'h429f7379, 32'h426852e1, 32'hc2943a17, 32'h41ed828d};
test_output[7241] = '{32'h42c4b943};
test_index[7241] = '{0};
test_input[57936:57943] = '{32'hc2537aa0, 32'h428a25f9, 32'hc2813d9c, 32'h4112a6bd, 32'h41c0e5ce, 32'hc231cdfe, 32'hc20d3075, 32'h428ef3b8};
test_output[7242] = '{32'h428ef3b8};
test_index[7242] = '{7};
test_input[57944:57951] = '{32'h42271432, 32'h429a62e6, 32'h425ae617, 32'h3e57106c, 32'hc2782bc2, 32'h421c4aa5, 32'h422d36a5, 32'hbf8f8d1d};
test_output[7243] = '{32'h429a62e6};
test_index[7243] = '{1};
test_input[57952:57959] = '{32'h410f7c7d, 32'h42bd54d3, 32'hc2493ae3, 32'h421016cc, 32'hc16052d6, 32'hc2b0a0db, 32'hc1a6bdc2, 32'h41b9d74b};
test_output[7244] = '{32'h42bd54d3};
test_index[7244] = '{1};
test_input[57960:57967] = '{32'h428d34da, 32'hc2447a2a, 32'hc29faabf, 32'h4291f0cb, 32'hc1e914ed, 32'h4291e3b4, 32'h42209710, 32'h4269c0ed};
test_output[7245] = '{32'h4291f0cb};
test_index[7245] = '{3};
test_input[57968:57975] = '{32'h41920d26, 32'hc2245bf4, 32'h428c70d3, 32'h41949fe4, 32'hc2345d54, 32'h42836017, 32'h426bdba4, 32'h420fd64f};
test_output[7246] = '{32'h428c70d3};
test_index[7246] = '{2};
test_input[57976:57983] = '{32'hc29ebb4d, 32'h42bc4b54, 32'hc2b85c7f, 32'h40e7441c, 32'hc171825e, 32'h418c5944, 32'hc1b3c4ff, 32'hc1ba5419};
test_output[7247] = '{32'h42bc4b54};
test_index[7247] = '{1};
test_input[57984:57991] = '{32'hc06a0a9a, 32'h42a0ba9c, 32'hc2b911bb, 32'h41b7b698, 32'hc1513a81, 32'hc06feb1d, 32'h41d33fcd, 32'hc197f12d};
test_output[7248] = '{32'h42a0ba9c};
test_index[7248] = '{1};
test_input[57992:57999] = '{32'hc2543a7c, 32'h4275ce1d, 32'h423e3779, 32'hc212de1a, 32'hc2a709a3, 32'h426fa4fc, 32'hc1e3ed3d, 32'h42360153};
test_output[7249] = '{32'h4275ce1d};
test_index[7249] = '{1};
test_input[58000:58007] = '{32'hc0885e98, 32'hc26dc796, 32'hc298523c, 32'hc151da63, 32'h42c36df5, 32'hc17d854d, 32'h3ea1df5d, 32'h4188ce56};
test_output[7250] = '{32'h42c36df5};
test_index[7250] = '{4};
test_input[58008:58015] = '{32'h4296bd10, 32'h42ae93cc, 32'h42344df8, 32'hc1ee8fb8, 32'hc216be60, 32'h4288abd7, 32'h415ba670, 32'h4275ea82};
test_output[7251] = '{32'h42ae93cc};
test_index[7251] = '{1};
test_input[58016:58023] = '{32'hc21f00a8, 32'hc2a8f412, 32'h42a681de, 32'h42b41562, 32'h418fa6e9, 32'h418a8e53, 32'h42978514, 32'h4158e6fe};
test_output[7252] = '{32'h42b41562};
test_index[7252] = '{3};
test_input[58024:58031] = '{32'hc15fb3da, 32'hc2c1e77d, 32'h42b7d2ff, 32'h41a433e6, 32'hc21481d3, 32'h42903de3, 32'h411e1ca5, 32'hc157ae7e};
test_output[7253] = '{32'h42b7d2ff};
test_index[7253] = '{2};
test_input[58032:58039] = '{32'h4252ea29, 32'h42c45307, 32'h413c4820, 32'hc2ae0a4d, 32'h40f50bdf, 32'h42469631, 32'hc2222a7f, 32'hc2b68e7c};
test_output[7254] = '{32'h42c45307};
test_index[7254] = '{1};
test_input[58040:58047] = '{32'hc28f35d9, 32'hc1c34dcf, 32'hc2159c40, 32'hc2a6d03b, 32'hc2ab97a1, 32'hc1d88f5a, 32'h4031fde1, 32'h425c33ee};
test_output[7255] = '{32'h425c33ee};
test_index[7255] = '{7};
test_input[58048:58055] = '{32'hc2b3db3f, 32'hc0b97689, 32'h4283041f, 32'hc2553aac, 32'hc2885276, 32'h42457711, 32'hc12b6b24, 32'hc2972d8b};
test_output[7256] = '{32'h4283041f};
test_index[7256] = '{2};
test_input[58056:58063] = '{32'hc22a5401, 32'h40a4defe, 32'hc2b76d32, 32'h42bbbc3a, 32'hc2617da8, 32'hc27dd77c, 32'h428eeea2, 32'h429c9032};
test_output[7257] = '{32'h42bbbc3a};
test_index[7257] = '{3};
test_input[58064:58071] = '{32'hc2ba0a59, 32'hc2babe3d, 32'hc0eeb2ea, 32'hc21d0dbf, 32'h41bff6d1, 32'h42bdd059, 32'hc1d133bc, 32'h4081912a};
test_output[7258] = '{32'h42bdd059};
test_index[7258] = '{5};
test_input[58072:58079] = '{32'hc20b7eab, 32'hc28e5246, 32'h41647295, 32'h42542e9b, 32'h420fc990, 32'hc1de8966, 32'hc1a6c3db, 32'h421c180a};
test_output[7259] = '{32'h42542e9b};
test_index[7259] = '{3};
test_input[58080:58087] = '{32'hc2908da8, 32'h424429b9, 32'h42c35555, 32'h420ec378, 32'h414c6f3f, 32'hc2be823f, 32'h4286af80, 32'hc18085d7};
test_output[7260] = '{32'h42c35555};
test_index[7260] = '{2};
test_input[58088:58095] = '{32'h41840820, 32'hc21371ad, 32'hc2a358ff, 32'hc2a25455, 32'hc09b26e5, 32'hc1b167d5, 32'h41e9d4ba, 32'h40e9c61e};
test_output[7261] = '{32'h41e9d4ba};
test_index[7261] = '{6};
test_input[58096:58103] = '{32'hc11b897f, 32'hc2101b37, 32'h42c6fb48, 32'h4288d1e9, 32'h428fa790, 32'hc1bebdbb, 32'h425bb87f, 32'hc13a57e6};
test_output[7262] = '{32'h42c6fb48};
test_index[7262] = '{2};
test_input[58104:58111] = '{32'h429753b5, 32'hc0123e26, 32'h42afa5b3, 32'h428c1208, 32'h42c79f71, 32'hc1f8c105, 32'h42999912, 32'hc1cb61c5};
test_output[7263] = '{32'h42c79f71};
test_index[7263] = '{4};
test_input[58112:58119] = '{32'hbedebaab, 32'h42b94d6d, 32'h418245dd, 32'h40d47aa5, 32'hc29f1d1c, 32'hc24ddb27, 32'hc1ba81c6, 32'hc1a18b97};
test_output[7264] = '{32'h42b94d6d};
test_index[7264] = '{1};
test_input[58120:58127] = '{32'h42965971, 32'hc2b93cc2, 32'hc29535aa, 32'hc09a0333, 32'h41a1a918, 32'h4296b7b7, 32'h427c3c7c, 32'hc2622b61};
test_output[7265] = '{32'h4296b7b7};
test_index[7265] = '{5};
test_input[58128:58135] = '{32'hc2178e76, 32'h42b43419, 32'h421dbff0, 32'hc09a4508, 32'h41ac2935, 32'hc1a36311, 32'h42964861, 32'hc2b64069};
test_output[7266] = '{32'h42b43419};
test_index[7266] = '{1};
test_input[58136:58143] = '{32'hc095339f, 32'h4299f198, 32'h41e689c8, 32'hc2b9de6c, 32'h42a01611, 32'hc214d45d, 32'hc219c560, 32'h41111667};
test_output[7267] = '{32'h42a01611};
test_index[7267] = '{4};
test_input[58144:58151] = '{32'h41fde440, 32'h42385599, 32'hc270b006, 32'h42c2bd21, 32'h41810caa, 32'hc2ba2094, 32'h413d3c83, 32'h421790d1};
test_output[7268] = '{32'h42c2bd21};
test_index[7268] = '{3};
test_input[58152:58159] = '{32'h42c60389, 32'h41cd5f72, 32'h41d0e7e9, 32'hc0bf5877, 32'h42aa3d1b, 32'hc2c08255, 32'h4237179d, 32'h41857daf};
test_output[7269] = '{32'h42c60389};
test_index[7269] = '{0};
test_input[58160:58167] = '{32'h4138fa74, 32'h4227dc46, 32'hc2a38c8d, 32'hc21d1863, 32'h424ee585, 32'h428ff58b, 32'hc20e0159, 32'h424217e5};
test_output[7270] = '{32'h428ff58b};
test_index[7270] = '{5};
test_input[58168:58175] = '{32'h42b9cf70, 32'hc236c3f1, 32'h41be3006, 32'h428f16f9, 32'hc1f5dfd6, 32'hc2b47850, 32'h42865c4e, 32'hc2af4577};
test_output[7271] = '{32'h42b9cf70};
test_index[7271] = '{0};
test_input[58176:58183] = '{32'hc1fcaa36, 32'h4135cfb9, 32'hc26d4f80, 32'hc2617ed1, 32'hc2af049a, 32'h418c5d55, 32'h413b1a86, 32'hc28f34dd};
test_output[7272] = '{32'h418c5d55};
test_index[7272] = '{5};
test_input[58184:58191] = '{32'h417312e7, 32'hc194a324, 32'hc277a60c, 32'hc2c26ee1, 32'h42b1971a, 32'hc24f1e43, 32'h42519fa4, 32'h42a11bf2};
test_output[7273] = '{32'h42b1971a};
test_index[7273] = '{4};
test_input[58192:58199] = '{32'h429f4fe5, 32'h424f8b04, 32'h3fc9dfaf, 32'h41aaa25f, 32'hc1923e12, 32'hc2a01f5c, 32'h42942041, 32'h41914f36};
test_output[7274] = '{32'h429f4fe5};
test_index[7274] = '{0};
test_input[58200:58207] = '{32'h423187d1, 32'h425c6bc8, 32'h428f9607, 32'h4288f1e9, 32'hc2b8ee1b, 32'h411c318b, 32'h41355cee, 32'hc114d2ab};
test_output[7275] = '{32'h428f9607};
test_index[7275] = '{2};
test_input[58208:58215] = '{32'hc1c6f4d5, 32'h42b62c97, 32'h428fd1ba, 32'hc2a880c9, 32'hc24faa13, 32'hc28dcb64, 32'hc2a51cef, 32'h42c716fb};
test_output[7276] = '{32'h42c716fb};
test_index[7276] = '{7};
test_input[58216:58223] = '{32'hc246e335, 32'h42c071dc, 32'h41dcf755, 32'h419c2d34, 32'h4018a49e, 32'h4097a190, 32'hc2a08e39, 32'h4186d745};
test_output[7277] = '{32'h42c071dc};
test_index[7277] = '{1};
test_input[58224:58231] = '{32'hc29a51fb, 32'h429d7074, 32'hc024b06c, 32'h428a9bdb, 32'hc2a050e2, 32'hc1da91fc, 32'hc2c1a6b3, 32'h4270976b};
test_output[7278] = '{32'h429d7074};
test_index[7278] = '{1};
test_input[58232:58239] = '{32'hc1d7c822, 32'h411401ab, 32'hc1ad44e5, 32'hc1c62c06, 32'hc1874e74, 32'hc2836b63, 32'h424a2744, 32'h413d5706};
test_output[7279] = '{32'h424a2744};
test_index[7279] = '{6};
test_input[58240:58247] = '{32'h420a05a7, 32'hc1c8f330, 32'hc2758f88, 32'h411d65a4, 32'h408ad389, 32'h4237aed0, 32'hc2820995, 32'hc1f1169f};
test_output[7280] = '{32'h4237aed0};
test_index[7280] = '{5};
test_input[58248:58255] = '{32'h4295bf7c, 32'hc22997f8, 32'hc276e38f, 32'h42a461f7, 32'hc22d4cde, 32'hc2bf8d6e, 32'h42ba9b1f, 32'hc208e1ea};
test_output[7281] = '{32'h42ba9b1f};
test_index[7281] = '{6};
test_input[58256:58263] = '{32'h425c5125, 32'hc1ea42d3, 32'h419df3e6, 32'hc111e6b0, 32'h423d3ee8, 32'hbe58f28c, 32'h429f2cea, 32'hc188e0f3};
test_output[7282] = '{32'h429f2cea};
test_index[7282] = '{6};
test_input[58264:58271] = '{32'h4166ce3d, 32'hc2c31b87, 32'h429971d3, 32'h42a12c35, 32'hc27c0047, 32'h42b0a783, 32'hc0a522f8, 32'hc19b252c};
test_output[7283] = '{32'h42b0a783};
test_index[7283] = '{5};
test_input[58272:58279] = '{32'h42bb42bf, 32'hc1f28ff9, 32'h4261bf8d, 32'hc0ec8032, 32'hc2ad30f9, 32'h4207e847, 32'h4215c7c4, 32'hc12bb197};
test_output[7284] = '{32'h42bb42bf};
test_index[7284] = '{0};
test_input[58280:58287] = '{32'hc230ad20, 32'h42ac3cc2, 32'h424b7140, 32'h427e40ae, 32'hc2b43438, 32'h42c1b215, 32'h423c72a8, 32'hc1d3e412};
test_output[7285] = '{32'h42c1b215};
test_index[7285] = '{5};
test_input[58288:58295] = '{32'h4284f243, 32'h42aa7c50, 32'h3fe75163, 32'hc2ba45bb, 32'h42241558, 32'h4123e86b, 32'hc2a0458d, 32'h40d49d69};
test_output[7286] = '{32'h42aa7c50};
test_index[7286] = '{1};
test_input[58296:58303] = '{32'hc25de4d0, 32'hc29190b5, 32'hc2a8c46b, 32'hc088602a, 32'h41e30582, 32'hc2890097, 32'hc2b9f22d, 32'h4213a664};
test_output[7287] = '{32'h4213a664};
test_index[7287] = '{7};
test_input[58304:58311] = '{32'h42ab423b, 32'hc20b8b36, 32'h429ca8f8, 32'h42aac1b9, 32'hc191e0ea, 32'h3fd06767, 32'h4299d96e, 32'h42113c59};
test_output[7288] = '{32'h42ab423b};
test_index[7288] = '{0};
test_input[58312:58319] = '{32'hc22b1fa4, 32'h4256b618, 32'h42b92d98, 32'h41f39abd, 32'hc23c997e, 32'h4159db54, 32'hc2427473, 32'hc1ed190a};
test_output[7289] = '{32'h42b92d98};
test_index[7289] = '{2};
test_input[58320:58327] = '{32'h42085fd5, 32'h428e0f61, 32'hc214c76b, 32'h409bcfb6, 32'hc26a8fda, 32'h428692c5, 32'h40cda41d, 32'h3fb93a68};
test_output[7290] = '{32'h428e0f61};
test_index[7290] = '{1};
test_input[58328:58335] = '{32'h42afc683, 32'hc1f16e83, 32'h41a4f2b3, 32'h41d44a1b, 32'h40bfd6ca, 32'hc1d05788, 32'hc1a13df3, 32'h4181081d};
test_output[7291] = '{32'h42afc683};
test_index[7291] = '{0};
test_input[58336:58343] = '{32'h4238192f, 32'h41bcbde8, 32'h42956e23, 32'hc278fb37, 32'h40520b0e, 32'hc2a640ed, 32'h42a0c09b, 32'hc2ac0de6};
test_output[7292] = '{32'h42a0c09b};
test_index[7292] = '{6};
test_input[58344:58351] = '{32'hc2491303, 32'hc2712371, 32'hc290e952, 32'hc28b071b, 32'hc29e9544, 32'hc227b074, 32'h42911526, 32'h4284e608};
test_output[7293] = '{32'h42911526};
test_index[7293] = '{6};
test_input[58352:58359] = '{32'h4171a809, 32'h425135ba, 32'hc2aad927, 32'h427e93e9, 32'hc2903df8, 32'hc20f2e4e, 32'h41e69ce2, 32'h425b2bdb};
test_output[7294] = '{32'h427e93e9};
test_index[7294] = '{3};
test_input[58360:58367] = '{32'hc143008b, 32'hc28866fc, 32'hc19e0dfb, 32'hc2375877, 32'h4190ce37, 32'hc001b9e6, 32'h42bbd99f, 32'hc0c3d107};
test_output[7295] = '{32'h42bbd99f};
test_index[7295] = '{6};
test_input[58368:58375] = '{32'hc2c0f4e6, 32'hc2ba7390, 32'hc2a15d5f, 32'h42365f24, 32'h42b5d62f, 32'hc21513db, 32'hc298fc0d, 32'hc1f1aac1};
test_output[7296] = '{32'h42b5d62f};
test_index[7296] = '{4};
test_input[58376:58383] = '{32'hc281af3b, 32'h41ec1219, 32'hc2845225, 32'h4192105d, 32'h411ee8c6, 32'h4210055c, 32'hc2b55ef0, 32'hc2987e27};
test_output[7297] = '{32'h4210055c};
test_index[7297] = '{5};
test_input[58384:58391] = '{32'hc267d7b6, 32'hc1bd6509, 32'hc29d6085, 32'hc25bf80e, 32'h41c52e2f, 32'hc2a79b51, 32'h41cfe461, 32'h42c1dd8d};
test_output[7298] = '{32'h42c1dd8d};
test_index[7298] = '{7};
test_input[58392:58399] = '{32'hc26c8b32, 32'hc24415a7, 32'h429f5fcc, 32'h410b9194, 32'h41295ef8, 32'h42066b75, 32'h41e721e4, 32'hc1842eaf};
test_output[7299] = '{32'h429f5fcc};
test_index[7299] = '{2};
test_input[58400:58407] = '{32'h4204adee, 32'hc2c7dc85, 32'hc2baf7e2, 32'h4218a2a7, 32'h42bf0eb7, 32'h41ecc7d6, 32'hc1a9002f, 32'hc24a9453};
test_output[7300] = '{32'h42bf0eb7};
test_index[7300] = '{4};
test_input[58408:58415] = '{32'hc16ac0e9, 32'h41d6ca3f, 32'hc2847ec5, 32'h421a64b5, 32'hc23453b8, 32'h4262f161, 32'hc1cff9ac, 32'hc1448393};
test_output[7301] = '{32'h4262f161};
test_index[7301] = '{5};
test_input[58416:58423] = '{32'hc2945722, 32'hc21dd2fe, 32'h42ace7eb, 32'hc13ff163, 32'hc2af0d03, 32'hc2318094, 32'hc2af7029, 32'h414ede27};
test_output[7302] = '{32'h42ace7eb};
test_index[7302] = '{2};
test_input[58424:58431] = '{32'h42299191, 32'hc0e71805, 32'h42a1b5aa, 32'hc129045b, 32'hc150a011, 32'hc2b03ec1, 32'hc2519492, 32'hc24372bc};
test_output[7303] = '{32'h42a1b5aa};
test_index[7303] = '{2};
test_input[58432:58439] = '{32'h41ea87f0, 32'h41fbf432, 32'h4101a016, 32'hc04ff0c7, 32'hc28c36c5, 32'hc268e1fa, 32'hc27ccf88, 32'h427507cc};
test_output[7304] = '{32'h427507cc};
test_index[7304] = '{7};
test_input[58440:58447] = '{32'h418b43fc, 32'h426748db, 32'hc1de379e, 32'h424e10e0, 32'h4292332e, 32'hc2a44c91, 32'hc0230a00, 32'hc2b66740};
test_output[7305] = '{32'h4292332e};
test_index[7305] = '{4};
test_input[58448:58455] = '{32'hc29b914f, 32'hbfe3d9c8, 32'h41ccce6d, 32'hc29fd14a, 32'hc216bbf6, 32'h42b91c2a, 32'h42af3844, 32'h419725f0};
test_output[7306] = '{32'h42b91c2a};
test_index[7306] = '{5};
test_input[58456:58463] = '{32'h41f67d13, 32'hc2be0e46, 32'h41d2ada6, 32'hc1ec1d6c, 32'h42c454b4, 32'hc1198ab9, 32'hc1ba178a, 32'hc2c20b94};
test_output[7307] = '{32'h42c454b4};
test_index[7307] = '{4};
test_input[58464:58471] = '{32'hc277dfa6, 32'hc299c9ed, 32'h4286f734, 32'h4273357b, 32'h4209e9a0, 32'hc28e01c1, 32'hc229813f, 32'hc2b5992e};
test_output[7308] = '{32'h4286f734};
test_index[7308] = '{2};
test_input[58472:58479] = '{32'hc1a626cf, 32'hc1d695cc, 32'hc273fb43, 32'hc1b26ec8, 32'hc2ad58a7, 32'h42a26fc2, 32'hc0e2474d, 32'hc292b578};
test_output[7309] = '{32'h42a26fc2};
test_index[7309] = '{5};
test_input[58480:58487] = '{32'h42b00221, 32'h429943cc, 32'h42a24246, 32'h42b2228f, 32'hc204e4fa, 32'hc2a52a37, 32'h41ed02af, 32'hc20246b4};
test_output[7310] = '{32'h42b2228f};
test_index[7310] = '{3};
test_input[58488:58495] = '{32'h40e95ab0, 32'hc21da7d5, 32'hc2bd04bc, 32'h428a7c7d, 32'h41cb1968, 32'hc146fb6f, 32'hc298b3dd, 32'h414bd1c6};
test_output[7311] = '{32'h428a7c7d};
test_index[7311] = '{3};
test_input[58496:58503] = '{32'h428852c2, 32'h42087230, 32'hc20d29db, 32'hc28ac84f, 32'h423934c6, 32'h421cb6c2, 32'hc28da18a, 32'h41b83da6};
test_output[7312] = '{32'h428852c2};
test_index[7312] = '{0};
test_input[58504:58511] = '{32'h42c138b3, 32'hc2a351da, 32'hc2c7788b, 32'hc26f7dde, 32'hc1a5f315, 32'hc1395ee4, 32'h41be17a0, 32'hc29a9959};
test_output[7313] = '{32'h42c138b3};
test_index[7313] = '{0};
test_input[58512:58519] = '{32'hc2721d4d, 32'h4291b57a, 32'hbed689c1, 32'hc2a1347c, 32'hc10c8dba, 32'h42926271, 32'hc2b097b6, 32'hc19792fc};
test_output[7314] = '{32'h42926271};
test_index[7314] = '{5};
test_input[58520:58527] = '{32'hc2c5db96, 32'hc1f064a3, 32'hc26ad30d, 32'hc292ff5f, 32'h4289b6f8, 32'h4288e13c, 32'h42134edd, 32'h41c38fd3};
test_output[7315] = '{32'h4289b6f8};
test_index[7315] = '{4};
test_input[58528:58535] = '{32'h42c77e6c, 32'h41b3c1dc, 32'h42a66715, 32'hc172615a, 32'hc2a54f8d, 32'h429e52ea, 32'hc2909e3e, 32'hc231052e};
test_output[7316] = '{32'h42c77e6c};
test_index[7316] = '{0};
test_input[58536:58543] = '{32'h40f7bf75, 32'hc28c1c90, 32'h4241dd56, 32'h4122d854, 32'h429d024c, 32'h42371ca7, 32'hc16bf2d4, 32'hc2180d09};
test_output[7317] = '{32'h429d024c};
test_index[7317] = '{4};
test_input[58544:58551] = '{32'h42aece16, 32'h429cc45e, 32'hc1f780c0, 32'h429d5527, 32'hc2a167c7, 32'hc2b45295, 32'hc13a9302, 32'h410ac341};
test_output[7318] = '{32'h42aece16};
test_index[7318] = '{0};
test_input[58552:58559] = '{32'hc272da6d, 32'h41ce4ee0, 32'hc2c63fb4, 32'h42c2a9c8, 32'h41d54dcd, 32'hc1072aa2, 32'h41f0a273, 32'h42935164};
test_output[7319] = '{32'h42c2a9c8};
test_index[7319] = '{3};
test_input[58560:58567] = '{32'hc272351c, 32'hc281b9c3, 32'hc1e03fbd, 32'h426164e6, 32'h417a9720, 32'h4282dae0, 32'h4294b13f, 32'hc262dade};
test_output[7320] = '{32'h4294b13f};
test_index[7320] = '{6};
test_input[58568:58575] = '{32'hc1976954, 32'h4187665f, 32'h42b873cd, 32'h42abf9b4, 32'h41fdace6, 32'hc2a3b0ea, 32'h4250cb5b, 32'hc2bfac1f};
test_output[7321] = '{32'h42b873cd};
test_index[7321] = '{2};
test_input[58576:58583] = '{32'h42137342, 32'h41d86512, 32'hc2ada885, 32'h42c661e6, 32'hc289ec78, 32'h42360ff5, 32'hc27e2483, 32'hc2753d64};
test_output[7322] = '{32'h42c661e6};
test_index[7322] = '{3};
test_input[58584:58591] = '{32'h4272d1e5, 32'h42aa053d, 32'hc260add9, 32'h41e8e34e, 32'h42aba2db, 32'h42beec2f, 32'h41892e27, 32'h419d9d49};
test_output[7323] = '{32'h42beec2f};
test_index[7323] = '{5};
test_input[58592:58599] = '{32'h41b64e88, 32'hc27f195b, 32'hc1574ec5, 32'h41a1b43c, 32'hc291b740, 32'h42a2cdad, 32'h4101b2ec, 32'h42b4afaa};
test_output[7324] = '{32'h42b4afaa};
test_index[7324] = '{7};
test_input[58600:58607] = '{32'h42b0ef38, 32'h421ab77b, 32'h42734118, 32'hc28d86c7, 32'h4278478e, 32'h427d697f, 32'h42b0a3d8, 32'hc2a83af9};
test_output[7325] = '{32'h42b0ef38};
test_index[7325] = '{0};
test_input[58608:58615] = '{32'hc2b9eaf8, 32'h422585b6, 32'hc2c70caf, 32'hc12a6acc, 32'h42457d04, 32'hc162f187, 32'hc2b49aea, 32'hc2abff47};
test_output[7326] = '{32'h42457d04};
test_index[7326] = '{4};
test_input[58616:58623] = '{32'hc1d046b0, 32'h4249d47d, 32'h4263993b, 32'hc2bca950, 32'hc2b674a6, 32'hc1e6270f, 32'h42ae980c, 32'hc291d53a};
test_output[7327] = '{32'h42ae980c};
test_index[7327] = '{6};
test_input[58624:58631] = '{32'hc2ac90dc, 32'hc29d00b1, 32'h42833a73, 32'h41eb0773, 32'hc239662e, 32'hc2c56eb4, 32'h42476938, 32'h42889161};
test_output[7328] = '{32'h42889161};
test_index[7328] = '{7};
test_input[58632:58639] = '{32'hc29e8e7f, 32'h4294c191, 32'hc28aeb93, 32'h41bf522e, 32'h423d79ab, 32'hc22c5181, 32'h419836a7, 32'hc050502b};
test_output[7329] = '{32'h4294c191};
test_index[7329] = '{1};
test_input[58640:58647] = '{32'hc1e44a48, 32'h42794032, 32'h42a6d595, 32'h41898a62, 32'h41159b6f, 32'h408aa353, 32'hc121d2c8, 32'hc1e7c009};
test_output[7330] = '{32'h42a6d595};
test_index[7330] = '{2};
test_input[58648:58655] = '{32'hc29afe3c, 32'h42a146f8, 32'h428c05e0, 32'h4218e4ed, 32'hc29dd39d, 32'hc25afb9c, 32'h428ad7cc, 32'h424c44bf};
test_output[7331] = '{32'h42a146f8};
test_index[7331] = '{1};
test_input[58656:58663] = '{32'hc0e88963, 32'h422d02dd, 32'h4285e560, 32'hc257c182, 32'hc2525a49, 32'h4240ed8f, 32'h4247d137, 32'h400f18cb};
test_output[7332] = '{32'h4285e560};
test_index[7332] = '{2};
test_input[58664:58671] = '{32'hc27085ca, 32'h42b5bbc3, 32'h42189b09, 32'h4289e0e4, 32'h411f8867, 32'hc2834844, 32'h422776f7, 32'hc2556d44};
test_output[7333] = '{32'h42b5bbc3};
test_index[7333] = '{1};
test_input[58672:58679] = '{32'hc20af447, 32'hc2c0850e, 32'hc2aa7ff2, 32'hc256231b, 32'h425197a3, 32'hc16d47d6, 32'h41349b8a, 32'hc29c64e0};
test_output[7334] = '{32'h425197a3};
test_index[7334] = '{4};
test_input[58680:58687] = '{32'h4059065d, 32'h42c5085b, 32'hc102faea, 32'hc28c0053, 32'hc1da1401, 32'hc20df0ab, 32'hc1f10970, 32'hc21c7939};
test_output[7335] = '{32'h42c5085b};
test_index[7335] = '{1};
test_input[58688:58695] = '{32'h42a1a16a, 32'h42ab0f01, 32'hc299b752, 32'h42b7dbd1, 32'hc26a68e3, 32'h428a2fd0, 32'hc2ab731f, 32'h421bc9b3};
test_output[7336] = '{32'h42b7dbd1};
test_index[7336] = '{3};
test_input[58696:58703] = '{32'hc2a9b5eb, 32'h40d53fd6, 32'h41a92249, 32'hc1f79c29, 32'h4280ad1d, 32'hc2782cb7, 32'h42b61ce1, 32'h42b97372};
test_output[7337] = '{32'h42b97372};
test_index[7337] = '{7};
test_input[58704:58711] = '{32'hc1eb57d2, 32'h42c565a5, 32'hc25819fe, 32'hc2b93426, 32'hc26808af, 32'h41cf882b, 32'hc14980ab, 32'hc2799f1c};
test_output[7338] = '{32'h42c565a5};
test_index[7338] = '{1};
test_input[58712:58719] = '{32'h4241a731, 32'hc1b2d2e9, 32'hc2160326, 32'h428a2bae, 32'h424781e6, 32'hc2abc621, 32'hc2c17366, 32'hc26faf70};
test_output[7339] = '{32'h428a2bae};
test_index[7339] = '{3};
test_input[58720:58727] = '{32'hc26b917c, 32'hc10f9bb5, 32'h42ac2ca3, 32'h411675f2, 32'hc28b3057, 32'hc210af04, 32'hc20b7d5f, 32'hc28f807a};
test_output[7340] = '{32'h42ac2ca3};
test_index[7340] = '{2};
test_input[58728:58735] = '{32'h42a41fbe, 32'hc218d087, 32'h42bcd5dc, 32'h4253716f, 32'h426120fd, 32'h41f0a979, 32'hc20cc556, 32'hc20e78c5};
test_output[7341] = '{32'h42bcd5dc};
test_index[7341] = '{2};
test_input[58736:58743] = '{32'h42680f67, 32'h424bd7e2, 32'h421419ba, 32'hc290119f, 32'h418b1451, 32'h42abe24c, 32'hc281a6a0, 32'h42079f92};
test_output[7342] = '{32'h42abe24c};
test_index[7342] = '{5};
test_input[58744:58751] = '{32'hc2735ff4, 32'h42bfa988, 32'h40afe36b, 32'hc2c3c208, 32'h41c0c467, 32'hc18ba4a4, 32'h42b97819, 32'h426077c7};
test_output[7343] = '{32'h42bfa988};
test_index[7343] = '{1};
test_input[58752:58759] = '{32'h4228d0c6, 32'h4214a6d4, 32'h4208a9d1, 32'h42c42271, 32'hc2a75d8b, 32'hc242ac8a, 32'h428d1ddd, 32'hc22caaa4};
test_output[7344] = '{32'h42c42271};
test_index[7344] = '{3};
test_input[58760:58767] = '{32'h42a25f98, 32'hc0e98d79, 32'hc29b41ae, 32'hc2b7704f, 32'h4195173c, 32'hc2b5016b, 32'h42b11a15, 32'h425f208f};
test_output[7345] = '{32'h42b11a15};
test_index[7345] = '{6};
test_input[58768:58775] = '{32'hc132cdba, 32'hc1198814, 32'h425eecd7, 32'hc29a7be1, 32'h41962fa1, 32'hc2b6c5e2, 32'h42acd214, 32'hc2ab9388};
test_output[7346] = '{32'h42acd214};
test_index[7346] = '{6};
test_input[58776:58783] = '{32'h42596b63, 32'h42a827e6, 32'hc23a0977, 32'hc18c5f5a, 32'hc23b501e, 32'h40d391db, 32'h416b0255, 32'hc2b61527};
test_output[7347] = '{32'h42a827e6};
test_index[7347] = '{1};
test_input[58784:58791] = '{32'hc2aac64f, 32'hc157ce77, 32'hc28a92fe, 32'h4200ee5d, 32'h410658e3, 32'h429bec70, 32'hc2bc944a, 32'h425cedec};
test_output[7348] = '{32'h429bec70};
test_index[7348] = '{5};
test_input[58792:58799] = '{32'h417e92bc, 32'h3fcec555, 32'hc25dec08, 32'h42332d76, 32'hc182daa1, 32'h42917d7d, 32'hc265341c, 32'h42b0ff4b};
test_output[7349] = '{32'h42b0ff4b};
test_index[7349] = '{7};
test_input[58800:58807] = '{32'h419365af, 32'hc1a3d853, 32'h41c54aef, 32'h4223a781, 32'hc24a4f6c, 32'hc01f6d6f, 32'h4225e865, 32'hc163729e};
test_output[7350] = '{32'h4225e865};
test_index[7350] = '{6};
test_input[58808:58815] = '{32'h41f6e7bf, 32'h42872c1d, 32'h418349e8, 32'hc1c9fa9e, 32'h41864c5c, 32'hc2223e56, 32'hc2a1e9bd, 32'hc248c71b};
test_output[7351] = '{32'h42872c1d};
test_index[7351] = '{1};
test_input[58816:58823] = '{32'h42a97d0a, 32'hc2ad7ca7, 32'h429f66de, 32'h4200e65b, 32'h41dba022, 32'hc26e5a81, 32'hc2b15b22, 32'h408ffaa2};
test_output[7352] = '{32'h42a97d0a};
test_index[7352] = '{0};
test_input[58824:58831] = '{32'hc0b60e81, 32'hc2c2c2ea, 32'h4219354b, 32'h421e0bc7, 32'hc2c50c40, 32'h3fd543d3, 32'h42467547, 32'h421e30d2};
test_output[7353] = '{32'h42467547};
test_index[7353] = '{6};
test_input[58832:58839] = '{32'h428acaaa, 32'h4287bebf, 32'hc0f5001e, 32'h42b19a0a, 32'h428c5bbb, 32'h42a20a3d, 32'h427f256a, 32'hc1cab1de};
test_output[7354] = '{32'h42b19a0a};
test_index[7354] = '{3};
test_input[58840:58847] = '{32'h42437c93, 32'hc222f690, 32'h423e7ff0, 32'h42909512, 32'hc20def6e, 32'h409109e2, 32'hc285adf5, 32'hbf0004be};
test_output[7355] = '{32'h42909512};
test_index[7355] = '{3};
test_input[58848:58855] = '{32'hc1594ee8, 32'h426a7001, 32'h425ebe47, 32'h42685be2, 32'h4219d958, 32'h4181a7c8, 32'hc211e49d, 32'h40373a1d};
test_output[7356] = '{32'h426a7001};
test_index[7356] = '{1};
test_input[58856:58863] = '{32'hc206f714, 32'h42b2336b, 32'h411b0703, 32'h41cc25ad, 32'hc2b0b296, 32'h4231be42, 32'hc1d71c56, 32'hbf8245ad};
test_output[7357] = '{32'h42b2336b};
test_index[7357] = '{1};
test_input[58864:58871] = '{32'hc2152d41, 32'h42a6de6c, 32'h41b7ff80, 32'h429b4da5, 32'hc1d4df6b, 32'h42b7347c, 32'h42bbe12b, 32'h41ff44aa};
test_output[7358] = '{32'h42bbe12b};
test_index[7358] = '{6};
test_input[58872:58879] = '{32'hc1674ff1, 32'h42a6d1e8, 32'hc18bea7c, 32'h42987565, 32'h42c227b8, 32'hc1bbbcc6, 32'hc28c0991, 32'h41bdced2};
test_output[7359] = '{32'h42c227b8};
test_index[7359] = '{4};
test_input[58880:58887] = '{32'hc2758111, 32'h42523479, 32'h4283541b, 32'hc22620e4, 32'h42b06b38, 32'h41b8106c, 32'h41df54aa, 32'hc27dc4ca};
test_output[7360] = '{32'h42b06b38};
test_index[7360] = '{4};
test_input[58888:58895] = '{32'h42b2008e, 32'h4287b44c, 32'hc121ee00, 32'hc20540ab, 32'h410bb166, 32'h42a09eb4, 32'hc274b7de, 32'h42c126e6};
test_output[7361] = '{32'h42c126e6};
test_index[7361] = '{7};
test_input[58896:58903] = '{32'hc2bbcdab, 32'hc23f20e6, 32'h42991f0a, 32'h4264ce9d, 32'h420d8a9c, 32'h4209aa16, 32'h416d2833, 32'hc2053855};
test_output[7362] = '{32'h42991f0a};
test_index[7362] = '{2};
test_input[58904:58911] = '{32'h4240cc77, 32'hc023597f, 32'h42591ee2, 32'hc0e57664, 32'h42af5599, 32'h42894966, 32'h42876152, 32'h418bfbf1};
test_output[7363] = '{32'h42af5599};
test_index[7363] = '{4};
test_input[58912:58919] = '{32'hc29c7c69, 32'hc2a925a8, 32'h42b6f96e, 32'hc1afa3b0, 32'hc25b3a1e, 32'hc2b4260e, 32'h428766d7, 32'hc23efdef};
test_output[7364] = '{32'h42b6f96e};
test_index[7364] = '{2};
test_input[58920:58927] = '{32'h42212ffe, 32'h42c1a973, 32'h422d3ae8, 32'hc296e6f4, 32'h42180c3f, 32'hc00f78fe, 32'hc287617c, 32'h424a84b0};
test_output[7365] = '{32'h42c1a973};
test_index[7365] = '{1};
test_input[58928:58935] = '{32'hc297ef7d, 32'hc283c3d1, 32'hc20ec6a3, 32'h42c00eef, 32'h401ef92c, 32'hc289fbaa, 32'h42c61865, 32'h4275d8ef};
test_output[7366] = '{32'h42c61865};
test_index[7366] = '{6};
test_input[58936:58943] = '{32'h41c37d8c, 32'h42bd2f73, 32'hc29a82fd, 32'h41a974fa, 32'h40ce1beb, 32'h4244d7a7, 32'h413293de, 32'hc22aede4};
test_output[7367] = '{32'h42bd2f73};
test_index[7367] = '{1};
test_input[58944:58951] = '{32'h41c44e4d, 32'h42a6d423, 32'hc2a25224, 32'hc1d8803f, 32'h42308776, 32'h425ec0ad, 32'h4252d131, 32'hc27944ee};
test_output[7368] = '{32'h42a6d423};
test_index[7368] = '{1};
test_input[58952:58959] = '{32'h4283083d, 32'h40cb49ee, 32'h41a6aefc, 32'hc1c2228d, 32'hc2be6980, 32'h407757d9, 32'hc189bc64, 32'h424b4591};
test_output[7369] = '{32'h4283083d};
test_index[7369] = '{0};
test_input[58960:58967] = '{32'h4296dd12, 32'hc0524f45, 32'hc2a96481, 32'hc1adc827, 32'hc298175a, 32'h4203e849, 32'h42b5497b, 32'hc20668e4};
test_output[7370] = '{32'h42b5497b};
test_index[7370] = '{6};
test_input[58968:58975] = '{32'hc1e52503, 32'hc2357cb2, 32'hc2be6304, 32'h41b3393f, 32'h417df17d, 32'h42910eed, 32'hc1d1ce4c, 32'h416bfc7e};
test_output[7371] = '{32'h42910eed};
test_index[7371] = '{5};
test_input[58976:58983] = '{32'h42899869, 32'h429b3419, 32'hc217786f, 32'hc2ba1c24, 32'h412d6298, 32'h42b2d039, 32'hc1f68a95, 32'hc2182c21};
test_output[7372] = '{32'h42b2d039};
test_index[7372] = '{5};
test_input[58984:58991] = '{32'hc2c470af, 32'hc29b0cbf, 32'hc269031c, 32'hc2bd9111, 32'h4182662d, 32'hc2b57a1a, 32'hc2b44587, 32'h42bc7fc5};
test_output[7373] = '{32'h42bc7fc5};
test_index[7373] = '{7};
test_input[58992:58999] = '{32'h423b9eda, 32'hc24dbb3e, 32'hc282a6c2, 32'h4218793c, 32'h4272c375, 32'h4293c09d, 32'hc1963516, 32'hc1ee84f4};
test_output[7374] = '{32'h4293c09d};
test_index[7374] = '{5};
test_input[59000:59007] = '{32'h428b3c45, 32'hc1263ff9, 32'h428cad9a, 32'h41c744d3, 32'h42971805, 32'h41c4fe7f, 32'hc289c02f, 32'h42c2fef3};
test_output[7375] = '{32'h42c2fef3};
test_index[7375] = '{7};
test_input[59008:59015] = '{32'hc1832c8e, 32'hc25f94b3, 32'h42885385, 32'hc26f1d51, 32'h429f4228, 32'hc204cd84, 32'hc209df28, 32'h426632ee};
test_output[7376] = '{32'h429f4228};
test_index[7376] = '{4};
test_input[59016:59023] = '{32'hc2a8a803, 32'hc22b08cc, 32'h41887ca7, 32'h42c062eb, 32'h42b0c94b, 32'hc1265c55, 32'h42c23b78, 32'hc22c2036};
test_output[7377] = '{32'h42c23b78};
test_index[7377] = '{6};
test_input[59024:59031] = '{32'hc2a1fc38, 32'h413dfb24, 32'hc2845a93, 32'h41cddaed, 32'hc2a11ed6, 32'h42ba4d36, 32'hc21e474f, 32'h425cb9af};
test_output[7378] = '{32'h42ba4d36};
test_index[7378] = '{5};
test_input[59032:59039] = '{32'h4273f9b5, 32'hc2837f0f, 32'hc1f33835, 32'hc2673f4a, 32'hc24fd6e7, 32'hc1b5d644, 32'hc1dd619f, 32'hc2721c1b};
test_output[7379] = '{32'h4273f9b5};
test_index[7379] = '{0};
test_input[59040:59047] = '{32'hc26f4347, 32'h428795b5, 32'hc2a59a7c, 32'hc28c6c2b, 32'hc2899589, 32'hc202d73a, 32'h424b2c8c, 32'hc1b576c0};
test_output[7380] = '{32'h428795b5};
test_index[7380] = '{1};
test_input[59048:59055] = '{32'hc2b581cf, 32'h42c16b6e, 32'hc216be72, 32'hc297e15c, 32'h411687bc, 32'h41327bc1, 32'h422f6fcb, 32'h415bb50c};
test_output[7381] = '{32'h42c16b6e};
test_index[7381] = '{1};
test_input[59056:59063] = '{32'h42c13f74, 32'hc18855bc, 32'h3edbd7c6, 32'h418ea271, 32'h4111eee7, 32'h41399d3a, 32'h422dfd12, 32'h41bb7a59};
test_output[7382] = '{32'h42c13f74};
test_index[7382] = '{0};
test_input[59064:59071] = '{32'hc2343db9, 32'hc1969297, 32'h429afa48, 32'hc238d46b, 32'h429e0ad7, 32'hc2a76d4e, 32'hc299070f, 32'h428175ba};
test_output[7383] = '{32'h429e0ad7};
test_index[7383] = '{4};
test_input[59072:59079] = '{32'h42ae1431, 32'hc2b1b1cf, 32'h425c5357, 32'hc20f2e26, 32'hc2aacd24, 32'h42a28ec4, 32'h42acc872, 32'h42a75033};
test_output[7384] = '{32'h42ae1431};
test_index[7384] = '{0};
test_input[59080:59087] = '{32'h42c7e121, 32'hc1337f2f, 32'h424c1138, 32'h422f6ec5, 32'hc227cce1, 32'hc2ac11af, 32'hc277f536, 32'hc2a23115};
test_output[7385] = '{32'h42c7e121};
test_index[7385] = '{0};
test_input[59088:59095] = '{32'h428d43a1, 32'hc1b9b666, 32'hc2b4e445, 32'h42224e82, 32'h428053d9, 32'hc1b91eb7, 32'hc262c957, 32'hc2bbecfd};
test_output[7386] = '{32'h428d43a1};
test_index[7386] = '{0};
test_input[59096:59103] = '{32'h42691f97, 32'h42899554, 32'h42a01f30, 32'hc264df57, 32'h4288bd5a, 32'h42409cbe, 32'h41d7e81e, 32'hc216d094};
test_output[7387] = '{32'h42a01f30};
test_index[7387] = '{2};
test_input[59104:59111] = '{32'h427274e8, 32'hc27b68a2, 32'hc2a79aa3, 32'hc2342133, 32'hc2a97fb0, 32'h42a732a8, 32'hc29ea169, 32'hc22ae0b1};
test_output[7388] = '{32'h42a732a8};
test_index[7388] = '{5};
test_input[59112:59119] = '{32'h429d7bda, 32'h4219d810, 32'hc297ac32, 32'h428f64cf, 32'h40c5e376, 32'hc2a62e9f, 32'h4210b805, 32'h42b2cf35};
test_output[7389] = '{32'h42b2cf35};
test_index[7389] = '{7};
test_input[59120:59127] = '{32'h420efe5c, 32'hc1070ded, 32'h408f1b2d, 32'h418a0df8, 32'hc2ae0325, 32'hc1ab0ddf, 32'hc2138cc3, 32'hc1980412};
test_output[7390] = '{32'h420efe5c};
test_index[7390] = '{0};
test_input[59128:59135] = '{32'hc1907b8d, 32'h428c44a0, 32'h4280fba4, 32'hc0ab7b77, 32'h42b376d5, 32'hc287aa2a, 32'h426811e8, 32'h42b2f965};
test_output[7391] = '{32'h42b376d5};
test_index[7391] = '{4};
test_input[59136:59143] = '{32'h42b6910f, 32'h415aab55, 32'hc21d7c90, 32'hc1887c31, 32'hc2afe712, 32'hc1daa8c2, 32'hc01b0ae0, 32'h424eaa24};
test_output[7392] = '{32'h42b6910f};
test_index[7392] = '{0};
test_input[59144:59151] = '{32'hc18ff394, 32'hc2bc8a9d, 32'hc2a0d9a0, 32'h42bc7f68, 32'h4247e963, 32'hc23a129f, 32'h422ef3b5, 32'h41da9fc2};
test_output[7393] = '{32'h42bc7f68};
test_index[7393] = '{3};
test_input[59152:59159] = '{32'hc22dd2f8, 32'h42028b8c, 32'hc2221926, 32'h421ca339, 32'h421cd2c1, 32'hc1856301, 32'h42c656fc, 32'h42ba8ad2};
test_output[7394] = '{32'h42c656fc};
test_index[7394] = '{6};
test_input[59160:59167] = '{32'h420950f7, 32'h41d4b799, 32'h4204d8bd, 32'hc087cabc, 32'h418ad564, 32'h41c0430b, 32'h424f77be, 32'hc2b3cb6a};
test_output[7395] = '{32'h424f77be};
test_index[7395] = '{6};
test_input[59168:59175] = '{32'h41bd3b2e, 32'hc266f9d8, 32'hc29d7d3a, 32'h42b3c9c7, 32'hc1a66a31, 32'h42865c88, 32'h41bf4c9d, 32'h41f83e73};
test_output[7396] = '{32'h42b3c9c7};
test_index[7396] = '{3};
test_input[59176:59183] = '{32'h4293e607, 32'hc28f0936, 32'h420372d6, 32'hc2960a78, 32'h427ad013, 32'hc1e821b7, 32'hc129843a, 32'hc0b45497};
test_output[7397] = '{32'h4293e607};
test_index[7397] = '{0};
test_input[59184:59191] = '{32'hc099f6d6, 32'h42a97865, 32'h42b7a5d5, 32'h42c11bc2, 32'h4239b275, 32'hc2021a0e, 32'h427fa24f, 32'hc0554be6};
test_output[7398] = '{32'h42c11bc2};
test_index[7398] = '{3};
test_input[59192:59199] = '{32'hc2204241, 32'hc2bd8a38, 32'h41a8a5dc, 32'hc09f5e4b, 32'h429644e8, 32'hc2a3fae2, 32'h42a771d7, 32'h42638efb};
test_output[7399] = '{32'h42a771d7};
test_index[7399] = '{6};
test_input[59200:59207] = '{32'h4244a85d, 32'h420a54bc, 32'hc28bdb90, 32'hc2af3a20, 32'hc24a1b87, 32'h410f0f5a, 32'h428d5fff, 32'hc189dcbf};
test_output[7400] = '{32'h428d5fff};
test_index[7400] = '{6};
test_input[59208:59215] = '{32'h4278bc14, 32'hc273a672, 32'hc2713a5a, 32'h4053a914, 32'hc289da38, 32'h41220f13, 32'h429896b6, 32'h4207b779};
test_output[7401] = '{32'h429896b6};
test_index[7401] = '{6};
test_input[59216:59223] = '{32'hc28c823e, 32'h427b5c34, 32'h429a372b, 32'h41418377, 32'hc0d778c4, 32'h422efe25, 32'hc23046a5, 32'hc226251f};
test_output[7402] = '{32'h429a372b};
test_index[7402] = '{2};
test_input[59224:59231] = '{32'h427b42b7, 32'hc28a55a2, 32'h412fa019, 32'hc14fe12a, 32'h42bce1be, 32'hc2927aec, 32'h413465d7, 32'h3feae9f7};
test_output[7403] = '{32'h42bce1be};
test_index[7403] = '{4};
test_input[59232:59239] = '{32'h41191a40, 32'h4268ee5b, 32'hc29b7ecf, 32'hc2aa79c2, 32'h4248b9d7, 32'hc1e32320, 32'hc2bb8428, 32'hc2892596};
test_output[7404] = '{32'h4268ee5b};
test_index[7404] = '{1};
test_input[59240:59247] = '{32'hc2229189, 32'hc1fab0cb, 32'h42896f5f, 32'h416651e8, 32'hc21f9228, 32'h429e748d, 32'h424950a9, 32'h412b59ef};
test_output[7405] = '{32'h429e748d};
test_index[7405] = '{5};
test_input[59248:59255] = '{32'hc29357cd, 32'h42bb778a, 32'hc1e1413e, 32'h42b8d524, 32'hc2818314, 32'hc1594c0a, 32'hc2bb2eed, 32'h42ab2531};
test_output[7406] = '{32'h42bb778a};
test_index[7406] = '{1};
test_input[59256:59263] = '{32'hc25c3454, 32'hc1bc5573, 32'h428d5eff, 32'hc21309a6, 32'hc1072aa8, 32'hc2935d96, 32'hc1f8449d, 32'hc2a91f82};
test_output[7407] = '{32'h428d5eff};
test_index[7407] = '{2};
test_input[59264:59271] = '{32'hc284b356, 32'hc26c07b8, 32'h42b7743a, 32'h42aaa5f0, 32'hc11eb425, 32'h40a82b26, 32'h42876f7b, 32'h41ea0361};
test_output[7408] = '{32'h42b7743a};
test_index[7408] = '{2};
test_input[59272:59279] = '{32'hc11f7c29, 32'hc1d0cf3a, 32'h406f3659, 32'h42119217, 32'hc2a7b564, 32'hbe3b51f1, 32'hc11ad22e, 32'h429e9d77};
test_output[7409] = '{32'h429e9d77};
test_index[7409] = '{7};
test_input[59280:59287] = '{32'hc23601e7, 32'h41840789, 32'h41aeea49, 32'h42b4b6fb, 32'h4063479c, 32'h429b105e, 32'h418bbee0, 32'hc2976c03};
test_output[7410] = '{32'h42b4b6fb};
test_index[7410] = '{3};
test_input[59288:59295] = '{32'hc1b3dd48, 32'hc1dcea3d, 32'hc2c723d4, 32'hc2c2cdb2, 32'h4298b31e, 32'h411e3970, 32'h428dc44e, 32'h42b0fa0b};
test_output[7411] = '{32'h42b0fa0b};
test_index[7411] = '{7};
test_input[59296:59303] = '{32'h411fe7d3, 32'hc1d78ac6, 32'hc2bc07f9, 32'h409c3749, 32'h405cfef5, 32'hc1c4b6ee, 32'h3f0033e1, 32'h4239038b};
test_output[7412] = '{32'h4239038b};
test_index[7412] = '{7};
test_input[59304:59311] = '{32'h42503cc0, 32'h4269a07e, 32'h428c81ac, 32'h4234efe8, 32'h4238b39b, 32'h4279ecf0, 32'hc166fb84, 32'hc2451afa};
test_output[7413] = '{32'h428c81ac};
test_index[7413] = '{2};
test_input[59312:59319] = '{32'hc15a20f6, 32'hc21caa32, 32'hc286186e, 32'h42c189a7, 32'hc2c06113, 32'h4291ded4, 32'h418aa545, 32'h42247b18};
test_output[7414] = '{32'h42c189a7};
test_index[7414] = '{3};
test_input[59320:59327] = '{32'h429697f3, 32'hc2ad2a05, 32'h42c71b01, 32'hc1a09e03, 32'h42a49dfa, 32'hc20aa395, 32'h42154f47, 32'h420b4743};
test_output[7415] = '{32'h42c71b01};
test_index[7415] = '{2};
test_input[59328:59335] = '{32'h420e7715, 32'h42140d73, 32'h428ee143, 32'h42b0788b, 32'h428288cf, 32'h42b3ed3d, 32'h42c21063, 32'hc2b71c87};
test_output[7416] = '{32'h42c21063};
test_index[7416] = '{6};
test_input[59336:59343] = '{32'hc283a51b, 32'h429d84e9, 32'h429d50ee, 32'h41c5f1ee, 32'h42ae1301, 32'hc243663a, 32'hc226f7d3, 32'hc1bbb61d};
test_output[7417] = '{32'h42ae1301};
test_index[7417] = '{4};
test_input[59344:59351] = '{32'hc2badd5a, 32'h421875b6, 32'h4289e64e, 32'h425f8624, 32'hc051dfdb, 32'hc18bcf8a, 32'hc1ee9965, 32'h42c7709a};
test_output[7418] = '{32'h42c7709a};
test_index[7418] = '{7};
test_input[59352:59359] = '{32'h418b12cc, 32'h429c6197, 32'hc1e2907a, 32'h4108a750, 32'hc20a9ff1, 32'h42c0b73a, 32'h42b0bd74, 32'hc28e062c};
test_output[7419] = '{32'h42c0b73a};
test_index[7419] = '{5};
test_input[59360:59367] = '{32'hc282023d, 32'hc0050bdf, 32'h428365a4, 32'h409e4d1e, 32'h42a46656, 32'h428d4d4f, 32'h42aef5ae, 32'hc1f10188};
test_output[7420] = '{32'h42aef5ae};
test_index[7420] = '{6};
test_input[59368:59375] = '{32'h4102ea9e, 32'h426e7341, 32'hc0d67e66, 32'hc217a584, 32'hc223055c, 32'h429ed61a, 32'hc24057a9, 32'h42a79fd4};
test_output[7421] = '{32'h42a79fd4};
test_index[7421] = '{7};
test_input[59376:59383] = '{32'hc229b22e, 32'h4236cf97, 32'h42a2d55e, 32'hc2b592d0, 32'hc1d686c3, 32'hc2c23b45, 32'hc2198040, 32'hc2349718};
test_output[7422] = '{32'h42a2d55e};
test_index[7422] = '{2};
test_input[59384:59391] = '{32'hc1bab4e8, 32'h414696f3, 32'h405bb380, 32'h41a3180c, 32'hbf1cf1e9, 32'h411f196c, 32'h42a6b92d, 32'h41a27ea2};
test_output[7423] = '{32'h42a6b92d};
test_index[7423] = '{6};
test_input[59392:59399] = '{32'h42576d01, 32'h42266c05, 32'h42525c8e, 32'hc25732b4, 32'hc2ba1b26, 32'hc23ba4b2, 32'hc2b43f84, 32'hc2c3591d};
test_output[7424] = '{32'h42576d01};
test_index[7424] = '{0};
test_input[59400:59407] = '{32'h425e487e, 32'h42a26354, 32'h42831e85, 32'hc1e55001, 32'hc291e603, 32'h4231ef35, 32'hc2c1a926, 32'hc2ae5835};
test_output[7425] = '{32'h42a26354};
test_index[7425] = '{1};
test_input[59408:59415] = '{32'hc2ad432c, 32'h428bf92e, 32'hc2698479, 32'hc2c0935e, 32'h41b01400, 32'hc2aada0f, 32'hc28f4a9a, 32'hc2a01c17};
test_output[7426] = '{32'h428bf92e};
test_index[7426] = '{1};
test_input[59416:59423] = '{32'h40d880af, 32'hc29e56ea, 32'h3f43834c, 32'hc1aff7ed, 32'hc2225e4d, 32'hc1cb91d1, 32'h42aad0d7, 32'h4273419c};
test_output[7427] = '{32'h42aad0d7};
test_index[7427] = '{6};
test_input[59424:59431] = '{32'hc24dc596, 32'h42441b86, 32'hc20100f6, 32'h42a157b0, 32'h41a63bfa, 32'h42a7202a, 32'h3eb2b3d4, 32'h426c719d};
test_output[7428] = '{32'h42a7202a};
test_index[7428] = '{5};
test_input[59432:59439] = '{32'hc2c04a6f, 32'hc09d8117, 32'h42784112, 32'hc2be5c45, 32'hc29a1b46, 32'h410e1c27, 32'hc2593467, 32'hc123141f};
test_output[7429] = '{32'h42784112};
test_index[7429] = '{2};
test_input[59440:59447] = '{32'h42168b53, 32'hc2285985, 32'h42654258, 32'h42b8ff65, 32'h41f385c3, 32'hc21c1ebb, 32'h42c1f049, 32'hc28ea431};
test_output[7430] = '{32'h42c1f049};
test_index[7430] = '{6};
test_input[59448:59455] = '{32'hc191f82b, 32'hbf6b1ffd, 32'h4108201a, 32'h422f4615, 32'h42801fc5, 32'hc2524408, 32'hc1f75842, 32'h42bdaf7f};
test_output[7431] = '{32'h42bdaf7f};
test_index[7431] = '{7};
test_input[59456:59463] = '{32'h418802d4, 32'h427ced5b, 32'h42b351b0, 32'h429c4e8a, 32'h4269f61f, 32'hc1a33fc9, 32'h410931f3, 32'h42a42d9d};
test_output[7432] = '{32'h42b351b0};
test_index[7432] = '{2};
test_input[59464:59471] = '{32'h415d6409, 32'h4233a853, 32'hc2aef60b, 32'hc0dc797a, 32'hc295c919, 32'hc2a16ae6, 32'h42a31bbe, 32'hc1ef590a};
test_output[7433] = '{32'h42a31bbe};
test_index[7433] = '{6};
test_input[59472:59479] = '{32'h4273b773, 32'hc2a7bb58, 32'h42b614b6, 32'h428cff42, 32'hc2172961, 32'h40bf2154, 32'h408029ec, 32'hc19ff64d};
test_output[7434] = '{32'h42b614b6};
test_index[7434] = '{2};
test_input[59480:59487] = '{32'h4106ef2e, 32'h429f9ce1, 32'h428e8a52, 32'h4229d64e, 32'h427d8be2, 32'h422fc6f9, 32'h4289d379, 32'hc21f08e8};
test_output[7435] = '{32'h429f9ce1};
test_index[7435] = '{1};
test_input[59488:59495] = '{32'hc1c892f1, 32'h429cf13f, 32'hc2644d5e, 32'h41c2f60f, 32'hc086fe8a, 32'hc1005331, 32'h42bd10c4, 32'h4085dc74};
test_output[7436] = '{32'h42bd10c4};
test_index[7436] = '{6};
test_input[59496:59503] = '{32'hbfbd1d11, 32'h4209f051, 32'hc25054e9, 32'h41ed0b8e, 32'hc2b721cb, 32'h42a54f9d, 32'h42243d63, 32'h4122b021};
test_output[7437] = '{32'h42a54f9d};
test_index[7437] = '{5};
test_input[59504:59511] = '{32'hc29058db, 32'h424efbbd, 32'h429c4392, 32'h428c5317, 32'hc2b8e011, 32'hc24ee23b, 32'hc19d1fe6, 32'h4169e020};
test_output[7438] = '{32'h429c4392};
test_index[7438] = '{2};
test_input[59512:59519] = '{32'h408e447d, 32'h42707f70, 32'h41e6782e, 32'hc2b9bc23, 32'h4206a354, 32'h429bc3c1, 32'hc2938f0f, 32'h42b05380};
test_output[7439] = '{32'h42b05380};
test_index[7439] = '{7};
test_input[59520:59527] = '{32'hc11ffc47, 32'hc10ca3fd, 32'hc216015d, 32'h42039913, 32'hc24cd2a1, 32'h41b85aba, 32'hc1959fc9, 32'hc2122a65};
test_output[7440] = '{32'h42039913};
test_index[7440] = '{3};
test_input[59528:59535] = '{32'h421ed5ce, 32'hc2a21d24, 32'hc29c08a0, 32'hbfa935dd, 32'hc25d17a7, 32'hc2a474b0, 32'h41b54aad, 32'hc1316b59};
test_output[7441] = '{32'h421ed5ce};
test_index[7441] = '{0};
test_input[59536:59543] = '{32'h42a59b60, 32'hc227fefb, 32'h42a4137f, 32'h4218d56c, 32'hc2247dde, 32'h427495ed, 32'h3ff3604a, 32'h412c371b};
test_output[7442] = '{32'h42a59b60};
test_index[7442] = '{0};
test_input[59544:59551] = '{32'h42c38404, 32'h4150b99e, 32'hc13c8a0b, 32'hc1233f28, 32'h41da743e, 32'h4299f6ab, 32'hc2bc77e2, 32'hc2133659};
test_output[7443] = '{32'h42c38404};
test_index[7443] = '{0};
test_input[59552:59559] = '{32'h42951143, 32'h421db4f9, 32'h423608e5, 32'h42875e12, 32'h4283b2df, 32'h424ed948, 32'h42337250, 32'h42529321};
test_output[7444] = '{32'h42951143};
test_index[7444] = '{0};
test_input[59560:59567] = '{32'h4180c350, 32'hc2a8125c, 32'hc2bfdd34, 32'h426ef72e, 32'h42829531, 32'hc28df101, 32'h42ac85a9, 32'hc26f122c};
test_output[7445] = '{32'h42ac85a9};
test_index[7445] = '{6};
test_input[59568:59575] = '{32'h41aa32ad, 32'hc22c0ce3, 32'hc2422b6c, 32'hc2377242, 32'h4003ebb4, 32'hc18921d5, 32'h41426bcd, 32'h42c12acd};
test_output[7446] = '{32'h42c12acd};
test_index[7446] = '{7};
test_input[59576:59583] = '{32'hc21114b0, 32'hc1932fb5, 32'h42ab04ca, 32'h413184d7, 32'hc22c2485, 32'hc2394759, 32'hc13a5028, 32'h4297ece4};
test_output[7447] = '{32'h42ab04ca};
test_index[7447] = '{2};
test_input[59584:59591] = '{32'hc28a29b6, 32'hc25f6f9c, 32'hc186bb2b, 32'h4254037a, 32'h41510c76, 32'hc2805bf1, 32'hc2360f5a, 32'hc201a53b};
test_output[7448] = '{32'h4254037a};
test_index[7448] = '{3};
test_input[59592:59599] = '{32'hc140752a, 32'hc230e675, 32'hc263ff0f, 32'hc2476a0d, 32'hc2289b56, 32'h41110434, 32'h42a34439, 32'h40fc9339};
test_output[7449] = '{32'h42a34439};
test_index[7449] = '{6};
test_input[59600:59607] = '{32'hc1ab5726, 32'h4294dacf, 32'h42534768, 32'h41d18755, 32'h4197ad60, 32'h420b461a, 32'hc2bb3d3e, 32'hc1a38a42};
test_output[7450] = '{32'h4294dacf};
test_index[7450] = '{1};
test_input[59608:59615] = '{32'h409e8203, 32'h41ad3aa0, 32'hc2832c11, 32'h4277a0fd, 32'h41b8a493, 32'hc123d28e, 32'hc138b712, 32'hbe7d556a};
test_output[7451] = '{32'h4277a0fd};
test_index[7451] = '{3};
test_input[59616:59623] = '{32'h413bb69f, 32'h4272f877, 32'hc2af2829, 32'hc2b6746d, 32'hc243ae28, 32'h42aefad9, 32'h41b93e3f, 32'hc2b3c992};
test_output[7452] = '{32'h42aefad9};
test_index[7452] = '{5};
test_input[59624:59631] = '{32'h41ba557b, 32'h41b3dce1, 32'hc1377f20, 32'h40e48722, 32'hc2024f93, 32'hc22986ef, 32'h424260a8, 32'hc23e93ca};
test_output[7453] = '{32'h424260a8};
test_index[7453] = '{6};
test_input[59632:59639] = '{32'h428e11c1, 32'h4283a77d, 32'hc257995e, 32'h422752ee, 32'hc1cc01a9, 32'hc209e0b5, 32'h4209504a, 32'h42b436a0};
test_output[7454] = '{32'h42b436a0};
test_index[7454] = '{7};
test_input[59640:59647] = '{32'h42aa1ddb, 32'hc2a8bba6, 32'h42936732, 32'hc22de3cd, 32'hc297a815, 32'hc1506d36, 32'hc278e9d8, 32'hc2b66364};
test_output[7455] = '{32'h42aa1ddb};
test_index[7455] = '{0};
test_input[59648:59655] = '{32'hc14925cc, 32'h42764384, 32'hc18d314b, 32'h41d2be6b, 32'hc14cc910, 32'h421bcbae, 32'h41cf1dc1, 32'hc29ae8ea};
test_output[7456] = '{32'h42764384};
test_index[7456] = '{1};
test_input[59656:59663] = '{32'h42b7c424, 32'hc23abd1c, 32'h429d8221, 32'h420f76bc, 32'h42abe60f, 32'h41aaf8b6, 32'hc2b75329, 32'hc1004500};
test_output[7457] = '{32'h42b7c424};
test_index[7457] = '{0};
test_input[59664:59671] = '{32'h428f7d97, 32'hc21be4dd, 32'hc1e39725, 32'hc284b95b, 32'hc2bbbb01, 32'hc28d8b5b, 32'hc1182625, 32'hbf9110ee};
test_output[7458] = '{32'h428f7d97};
test_index[7458] = '{0};
test_input[59672:59679] = '{32'h42082772, 32'hc28b97d0, 32'h4200f060, 32'h42a3de95, 32'hc25da5ce, 32'hc2193195, 32'hc16301fe, 32'h42112581};
test_output[7459] = '{32'h42a3de95};
test_index[7459] = '{3};
test_input[59680:59687] = '{32'h42b43a78, 32'h41684494, 32'h4206d213, 32'hc29493c4, 32'hc2531017, 32'hc25ab4f6, 32'hc2c184a6, 32'h4291da2e};
test_output[7460] = '{32'h42b43a78};
test_index[7460] = '{0};
test_input[59688:59695] = '{32'hc20fe9c2, 32'h4222cc74, 32'h42a8f0f4, 32'hc29e0eb5, 32'hc250561c, 32'h41a3c5ab, 32'hc2024ee1, 32'hc29ae086};
test_output[7461] = '{32'h42a8f0f4};
test_index[7461] = '{2};
test_input[59696:59703] = '{32'hc25a2275, 32'hc264f537, 32'h426c26f6, 32'h422c6186, 32'h4256057d, 32'hc281a5eb, 32'h42c3e68d, 32'h42a59806};
test_output[7462] = '{32'h42c3e68d};
test_index[7462] = '{6};
test_input[59704:59711] = '{32'h42c1fcf4, 32'h42b70deb, 32'h42b8902d, 32'h4295de6b, 32'h41f8084f, 32'h42252895, 32'hc1b3f009, 32'h4196afdc};
test_output[7463] = '{32'h42c1fcf4};
test_index[7463] = '{0};
test_input[59712:59719] = '{32'h427bcb08, 32'hc18a9992, 32'h42b14c42, 32'h4182e0e0, 32'h428b05a6, 32'hc22182de, 32'h4249bc96, 32'hc2a9dbc6};
test_output[7464] = '{32'h42b14c42};
test_index[7464] = '{2};
test_input[59720:59727] = '{32'hc293ea62, 32'h416f387e, 32'hc287f669, 32'h4278b648, 32'h426e1b8c, 32'h428db238, 32'hc2a9afef, 32'h4282cc06};
test_output[7465] = '{32'h428db238};
test_index[7465] = '{5};
test_input[59728:59735] = '{32'h4227c041, 32'hc183a268, 32'hc0cc2b17, 32'hc295a63f, 32'hc27a0136, 32'hc222f8de, 32'hc29d8fd3, 32'h42ad020f};
test_output[7466] = '{32'h42ad020f};
test_index[7466] = '{7};
test_input[59736:59743] = '{32'hc1b6b754, 32'hc21ae8dd, 32'hc286236e, 32'h42b37c8a, 32'hc20edd4d, 32'hc1f5e4f0, 32'hc2298c12, 32'h429fb9de};
test_output[7467] = '{32'h42b37c8a};
test_index[7467] = '{3};
test_input[59744:59751] = '{32'hc21fd8de, 32'hc252b4d8, 32'hc2b7c9f6, 32'h42afbd4b, 32'hc10f9396, 32'h429ab396, 32'h423e00cc, 32'h4227d0ad};
test_output[7468] = '{32'h42afbd4b};
test_index[7468] = '{3};
test_input[59752:59759] = '{32'hc2b2c8d0, 32'h42a4281d, 32'hc0869c8d, 32'hc24521d3, 32'h42bcb6bd, 32'h426e70ce, 32'h41b83bef, 32'hc13692e5};
test_output[7469] = '{32'h42bcb6bd};
test_index[7469] = '{4};
test_input[59760:59767] = '{32'h427452b9, 32'hc161eef1, 32'hc211bba6, 32'hc1ef248a, 32'hbf33b881, 32'h42892689, 32'hc11a0af3, 32'hc2256fdd};
test_output[7470] = '{32'h42892689};
test_index[7470] = '{5};
test_input[59768:59775] = '{32'h41b9f47e, 32'h4291dddd, 32'hc1cf5451, 32'h42306e51, 32'hc20bf103, 32'hc2b6fcf2, 32'hc2ab645f, 32'hc230fa2b};
test_output[7471] = '{32'h4291dddd};
test_index[7471] = '{1};
test_input[59776:59783] = '{32'hbdbca4b5, 32'h41bc246a, 32'hc1ee0a0d, 32'hc0e08b93, 32'h425fdd9c, 32'h429829db, 32'hc28fd782, 32'hc267711f};
test_output[7472] = '{32'h429829db};
test_index[7472] = '{5};
test_input[59784:59791] = '{32'hc233f63c, 32'hc19b3ac1, 32'h41a2af03, 32'hc27d1319, 32'h420a7eea, 32'hc2c2337f, 32'hc2064ee7, 32'h429bf7ed};
test_output[7473] = '{32'h429bf7ed};
test_index[7473] = '{7};
test_input[59792:59799] = '{32'hc1f375cc, 32'hc13755db, 32'hc27ffef9, 32'hc263213f, 32'hc0867e62, 32'hc24efba4, 32'h4234958b, 32'h41d2f990};
test_output[7474] = '{32'h4234958b};
test_index[7474] = '{6};
test_input[59800:59807] = '{32'h421e3fe1, 32'h4149955a, 32'h42704274, 32'h42611288, 32'hc138425d, 32'h40b6e24e, 32'h41d47396, 32'hc263fe0a};
test_output[7475] = '{32'h42704274};
test_index[7475] = '{2};
test_input[59808:59815] = '{32'h426afd38, 32'hc1b384e5, 32'h42b6afbe, 32'h420c9ce8, 32'hc0b7a3b8, 32'hc208a805, 32'hc26725c5, 32'hc24d6a72};
test_output[7476] = '{32'h42b6afbe};
test_index[7476] = '{2};
test_input[59816:59823] = '{32'h42a664d8, 32'hc21776cf, 32'h42b432f4, 32'h428ba424, 32'h42b25202, 32'h426a0c17, 32'hc1c6420a, 32'h423a9051};
test_output[7477] = '{32'h42b432f4};
test_index[7477] = '{2};
test_input[59824:59831] = '{32'h42a4de39, 32'hc20868ca, 32'hc27ae282, 32'hc2bec477, 32'h4183f38c, 32'h42c29ae1, 32'h418892f8, 32'hc293e356};
test_output[7478] = '{32'h42c29ae1};
test_index[7478] = '{5};
test_input[59832:59839] = '{32'hc1b4aaae, 32'hc29a514e, 32'h429d8ac2, 32'h425f0d9e, 32'h420c234f, 32'h42020e7f, 32'hc1ea5c34, 32'h4244170b};
test_output[7479] = '{32'h429d8ac2};
test_index[7479] = '{2};
test_input[59840:59847] = '{32'h4292c78a, 32'h42063f34, 32'h42761aa5, 32'h42138bc3, 32'hc1de0ba3, 32'hc246f08f, 32'h41f7f28d, 32'h4277975c};
test_output[7480] = '{32'h4292c78a};
test_index[7480] = '{0};
test_input[59848:59855] = '{32'hc25f5227, 32'h429eb803, 32'hc28a6ab1, 32'h42015b76, 32'h42c63131, 32'h42b4cb21, 32'h42c1954e, 32'h4272d185};
test_output[7481] = '{32'h42c63131};
test_index[7481] = '{4};
test_input[59856:59863] = '{32'h42374ba3, 32'hc238c37d, 32'hc29f1256, 32'hc2b023b6, 32'hc23c4022, 32'h421ee2f6, 32'h4205adfc, 32'h41091096};
test_output[7482] = '{32'h42374ba3};
test_index[7482] = '{0};
test_input[59864:59871] = '{32'h42c62f3f, 32'hc12ba34d, 32'h41ca375b, 32'hc0e8f759, 32'hc2008635, 32'h4022e119, 32'hc2b23204, 32'hc23fdb94};
test_output[7483] = '{32'h42c62f3f};
test_index[7483] = '{0};
test_input[59872:59879] = '{32'hc0a8980c, 32'hc2328cbb, 32'h42211fbb, 32'hc299f57a, 32'hc2a9adf5, 32'h42016db3, 32'hc275aae8, 32'h421e7ebe};
test_output[7484] = '{32'h42211fbb};
test_index[7484] = '{2};
test_input[59880:59887] = '{32'hc21e9d1d, 32'hc28ee192, 32'hc1f716db, 32'hc2b19ec0, 32'hc2268c0a, 32'hc29de406, 32'h41051fff, 32'hc274781c};
test_output[7485] = '{32'h41051fff};
test_index[7485] = '{6};
test_input[59888:59895] = '{32'hc25b0c4e, 32'h423b4f65, 32'h4250c36a, 32'h427ac46c, 32'hc28a46e6, 32'h42c46396, 32'h428b300c, 32'h42697493};
test_output[7486] = '{32'h42c46396};
test_index[7486] = '{5};
test_input[59896:59903] = '{32'h41ad51c3, 32'h4284c5a6, 32'hc1e482f0, 32'hc2b8301f, 32'h42af2cea, 32'hc1505913, 32'hc288cde4, 32'hc265e7be};
test_output[7487] = '{32'h42af2cea};
test_index[7487] = '{4};
test_input[59904:59911] = '{32'hc24649d8, 32'h41c4a0c2, 32'hc2c42b79, 32'h41b4b950, 32'hc185f6f1, 32'hc259e98d, 32'h42b68357, 32'hc27fb711};
test_output[7488] = '{32'h42b68357};
test_index[7488] = '{6};
test_input[59912:59919] = '{32'hc266fafc, 32'h4206af5e, 32'hc2b1d029, 32'hc11f5da2, 32'hc29b6732, 32'h426a3e69, 32'h424aaf14, 32'h42c07f74};
test_output[7489] = '{32'h42c07f74};
test_index[7489] = '{7};
test_input[59920:59927] = '{32'h42097250, 32'h420007c7, 32'hc2382224, 32'hc24829bf, 32'hc210c1fd, 32'hc2b845f4, 32'h42c458c4, 32'hc2b78869};
test_output[7490] = '{32'h42c458c4};
test_index[7490] = '{6};
test_input[59928:59935] = '{32'hc2a21423, 32'hc26a7f17, 32'h42b272a6, 32'hc1b78978, 32'h42aebcd9, 32'hc2499e53, 32'hc1e5ab9a, 32'h42ac25b9};
test_output[7491] = '{32'h42b272a6};
test_index[7491] = '{2};
test_input[59936:59943] = '{32'hc21e1693, 32'hc273f780, 32'h42c011cf, 32'hc29094fd, 32'hc2b8ca67, 32'hc2c1ce79, 32'h42b363f1, 32'hc29975de};
test_output[7492] = '{32'h42c011cf};
test_index[7492] = '{2};
test_input[59944:59951] = '{32'hc1c6f1dc, 32'hc2597370, 32'hc2c74c6f, 32'h424e5609, 32'h42a982b5, 32'h42688f5c, 32'h42a04763, 32'h428f2cfe};
test_output[7493] = '{32'h42a982b5};
test_index[7493] = '{4};
test_input[59952:59959] = '{32'h420afdd2, 32'h42929e6c, 32'h41fa82be, 32'h42ac34e4, 32'h422f2ed2, 32'hc165c4ee, 32'h426ce631, 32'hc15dc25e};
test_output[7494] = '{32'h42ac34e4};
test_index[7494] = '{3};
test_input[59960:59967] = '{32'h42c0a41c, 32'h424adf68, 32'h413834b6, 32'hc282c589, 32'hc2ae4f0d, 32'hc203b0b0, 32'h420ef5f0, 32'hc2c4cd8f};
test_output[7495] = '{32'h42c0a41c};
test_index[7495] = '{0};
test_input[59968:59975] = '{32'h41ea8250, 32'h426bc508, 32'hc1b24785, 32'hc287d733, 32'hc243bbef, 32'h422cf7e5, 32'hc2936e66, 32'hc2020e73};
test_output[7496] = '{32'h426bc508};
test_index[7496] = '{1};
test_input[59976:59983] = '{32'h427aaced, 32'h422c9b7a, 32'hc26359bc, 32'hc2a8e68c, 32'hc0442546, 32'hc2260093, 32'h42560595, 32'hc043c12f};
test_output[7497] = '{32'h427aaced};
test_index[7497] = '{0};
test_input[59984:59991] = '{32'h42b3b480, 32'h427e106a, 32'hc2bad0a6, 32'h429a83b6, 32'hc0b0d407, 32'hc28a12d2, 32'hc27f2fba, 32'hc144b281};
test_output[7498] = '{32'h42b3b480};
test_index[7498] = '{0};
test_input[59992:59999] = '{32'h41b45c43, 32'h42227827, 32'h429eeceb, 32'hc22bc22c, 32'hc2997dbd, 32'hc231444c, 32'hc2b62618, 32'h42843853};
test_output[7499] = '{32'h429eeceb};
test_index[7499] = '{2};
test_input[60000:60007] = '{32'h41255a65, 32'h422b0df3, 32'h425f5743, 32'h41a8f222, 32'h4250aa31, 32'hc28dfe16, 32'hc222ee5a, 32'h41a83a61};
test_output[7500] = '{32'h425f5743};
test_index[7500] = '{2};
test_input[60008:60015] = '{32'h4247f348, 32'h42a1212e, 32'hc2c709be, 32'hc2c1d29b, 32'hc13acfca, 32'hc2b9d222, 32'hc295a3bc, 32'h4093f2d2};
test_output[7501] = '{32'h42a1212e};
test_index[7501] = '{1};
test_input[60016:60023] = '{32'hc25c509c, 32'hc23001c3, 32'hc0ef148c, 32'hc1b9327d, 32'hc2198186, 32'hc20a457e, 32'h420795d3, 32'h41740361};
test_output[7502] = '{32'h420795d3};
test_index[7502] = '{6};
test_input[60024:60031] = '{32'h42765880, 32'hc2b4c640, 32'h42151509, 32'hc2689224, 32'h41fbb390, 32'hc220cbbc, 32'h42855263, 32'hc2b617b2};
test_output[7503] = '{32'h42855263};
test_index[7503] = '{6};
test_input[60032:60039] = '{32'h4001a2a7, 32'hc2a29d5d, 32'hc267735d, 32'h4268534d, 32'h42a8bf8d, 32'hc2c54bed, 32'hc1eb54b8, 32'hc1748b6c};
test_output[7504] = '{32'h42a8bf8d};
test_index[7504] = '{4};
test_input[60040:60047] = '{32'hc274059a, 32'h42778a79, 32'h42535f7c, 32'hc13c64e6, 32'hc234f9e5, 32'hc28eec72, 32'hc279f1e5, 32'hc2bfde09};
test_output[7505] = '{32'h42778a79};
test_index[7505] = '{1};
test_input[60048:60055] = '{32'hc2872dd1, 32'hc216159f, 32'h42a3dedb, 32'hc20cbd07, 32'h3fff81c5, 32'hc2abde46, 32'h42b18d3f, 32'h42b244a4};
test_output[7506] = '{32'h42b244a4};
test_index[7506] = '{7};
test_input[60056:60063] = '{32'h4113e133, 32'hc2b6fe6c, 32'h418d0d01, 32'hc2176f31, 32'hc2c59e25, 32'hc2802e1c, 32'h42a34e46, 32'hc18a0965};
test_output[7507] = '{32'h42a34e46};
test_index[7507] = '{6};
test_input[60064:60071] = '{32'h40e709fe, 32'hc24bb945, 32'hc0399848, 32'h427f6697, 32'h424d93eb, 32'h4230dd04, 32'h41c39265, 32'hc2687796};
test_output[7508] = '{32'h427f6697};
test_index[7508] = '{3};
test_input[60072:60079] = '{32'hc1f89b11, 32'hc2ad3c97, 32'h413d24ec, 32'h41ee3be4, 32'h42b09ecd, 32'hc2a8da54, 32'hc29da9a3, 32'hc1f4d4aa};
test_output[7509] = '{32'h42b09ecd};
test_index[7509] = '{4};
test_input[60080:60087] = '{32'hc23a0241, 32'h4294262e, 32'h4249d478, 32'h42483b97, 32'hc11328ca, 32'h429aba76, 32'h425764f0, 32'hc2359364};
test_output[7510] = '{32'h429aba76};
test_index[7510] = '{5};
test_input[60088:60095] = '{32'h420f511d, 32'h428ea10c, 32'hc1ad0300, 32'h419f77b1, 32'hc28af864, 32'h4286041c, 32'h419271cc, 32'hc2474bf8};
test_output[7511] = '{32'h428ea10c};
test_index[7511] = '{1};
test_input[60096:60103] = '{32'h421588bc, 32'h42ad4a3b, 32'hc25c4391, 32'h42943fb6, 32'h42af8812, 32'h424ba350, 32'h41b22b10, 32'hc1cb768b};
test_output[7512] = '{32'h42af8812};
test_index[7512] = '{4};
test_input[60104:60111] = '{32'h423d6202, 32'h41a93fc8, 32'h429551b8, 32'hc2a8be9a, 32'h429810f7, 32'hc274160c, 32'h422936ba, 32'h422d3cd4};
test_output[7513] = '{32'h429810f7};
test_index[7513] = '{4};
test_input[60112:60119] = '{32'h41e25503, 32'hc2045b6f, 32'h4199c927, 32'hc29dd59f, 32'hc2b34adb, 32'h42553776, 32'h41fa23b0, 32'hc28daefc};
test_output[7514] = '{32'h42553776};
test_index[7514] = '{5};
test_input[60120:60127] = '{32'h41c39220, 32'hc2aa24ab, 32'h41375c92, 32'hc2286f96, 32'h42c7ee74, 32'hc1bb9a87, 32'h41349fbc, 32'hc1cb4d21};
test_output[7515] = '{32'h42c7ee74};
test_index[7515] = '{4};
test_input[60128:60135] = '{32'h42ba30c4, 32'hc2b1780a, 32'h425a8aba, 32'h42234dd9, 32'hc2c5588b, 32'hc118ea42, 32'h429c33fb, 32'h4249fa96};
test_output[7516] = '{32'h42ba30c4};
test_index[7516] = '{0};
test_input[60136:60143] = '{32'hc1a45698, 32'h4259f016, 32'hc2a60707, 32'h4242716e, 32'h419df6e1, 32'hc2055fc6, 32'hc2c65465, 32'h424c58e8};
test_output[7517] = '{32'h4259f016};
test_index[7517] = '{1};
test_input[60144:60151] = '{32'h42c0c89d, 32'hc2551cd9, 32'h42514ece, 32'h4209e62d, 32'hc210bf71, 32'h42aa3808, 32'h41cf4b34, 32'h42b858dd};
test_output[7518] = '{32'h42c0c89d};
test_index[7518] = '{0};
test_input[60152:60159] = '{32'h407afcc8, 32'h410a022d, 32'hc2834b98, 32'hc2c1a797, 32'h41c5d6fb, 32'h4293860c, 32'hc29dc6f1, 32'hc189451f};
test_output[7519] = '{32'h4293860c};
test_index[7519] = '{5};
test_input[60160:60167] = '{32'h41693fb4, 32'hc26a43fb, 32'h41eb3612, 32'h41403e69, 32'hc28fb12c, 32'hc2b98beb, 32'h42553dc8, 32'h41e0bed8};
test_output[7520] = '{32'h42553dc8};
test_index[7520] = '{6};
test_input[60168:60175] = '{32'h41eca4e6, 32'hc22c2212, 32'hc262e61b, 32'hc29b7712, 32'hc1488700, 32'hc24b6590, 32'hc291df1f, 32'hc23a453f};
test_output[7521] = '{32'h41eca4e6};
test_index[7521] = '{0};
test_input[60176:60183] = '{32'hc234d11e, 32'hc1f17ada, 32'hc2343907, 32'h41065802, 32'hc2a84c71, 32'hc2b65b0a, 32'hc2939f76, 32'hc1055c66};
test_output[7522] = '{32'h41065802};
test_index[7522] = '{3};
test_input[60184:60191] = '{32'hc2c62df8, 32'hc28c139d, 32'hc1817786, 32'hc2220221, 32'hc28782d1, 32'h42a0475d, 32'hc0bef9b1, 32'hc1137d92};
test_output[7523] = '{32'h42a0475d};
test_index[7523] = '{5};
test_input[60192:60199] = '{32'hc1f52bf5, 32'h42199dc4, 32'hc2a90edb, 32'hc2bafbc9, 32'h4265556b, 32'hc28b7b48, 32'h42a81101, 32'h4296e400};
test_output[7524] = '{32'h42a81101};
test_index[7524] = '{6};
test_input[60200:60207] = '{32'hc2b42b7a, 32'hc23e6b2a, 32'hc297d873, 32'h42805093, 32'h4201c7be, 32'h428cf2dd, 32'h41f607ca, 32'hc222681e};
test_output[7525] = '{32'h428cf2dd};
test_index[7525] = '{5};
test_input[60208:60215] = '{32'hc2ab48a3, 32'h4295528f, 32'h418123b8, 32'hc217f789, 32'h42846719, 32'hc221115a, 32'hc2960b90, 32'h42a63185};
test_output[7526] = '{32'h42a63185};
test_index[7526] = '{7};
test_input[60216:60223] = '{32'h4265a99b, 32'hc25d6070, 32'hc1612b87, 32'h4225c184, 32'h42c458f2, 32'h42261b25, 32'hc08e98b4, 32'h423c2c32};
test_output[7527] = '{32'h42c458f2};
test_index[7527] = '{4};
test_input[60224:60231] = '{32'h410c08ff, 32'h41341d10, 32'hc1dfd212, 32'hc1df895f, 32'hc245a1c7, 32'h42553a56, 32'h4270f311, 32'hc29bece3};
test_output[7528] = '{32'h4270f311};
test_index[7528] = '{6};
test_input[60232:60239] = '{32'hc2373452, 32'hc23c15e4, 32'hc24c3cf1, 32'h42976a96, 32'hc2c631a5, 32'hc116fd15, 32'hc2b4bff6, 32'h42a19a84};
test_output[7529] = '{32'h42a19a84};
test_index[7529] = '{7};
test_input[60240:60247] = '{32'hc27fe2ef, 32'h423bead4, 32'h428cc47d, 32'hc23d4c62, 32'h42886f59, 32'hc2132744, 32'hc2a07431, 32'h42b1bb2b};
test_output[7530] = '{32'h42b1bb2b};
test_index[7530] = '{7};
test_input[60248:60255] = '{32'h41f0d6aa, 32'h428c5c93, 32'h418364d0, 32'h42c3e2e9, 32'h42baada5, 32'hc2b3d2f0, 32'h42913390, 32'h428e9fd4};
test_output[7531] = '{32'h42c3e2e9};
test_index[7531] = '{3};
test_input[60256:60263] = '{32'h424044c4, 32'h41f4d40f, 32'hc286c2e9, 32'hc235cf50, 32'h41417f06, 32'h4280735f, 32'hc29d8d36, 32'h421283f0};
test_output[7532] = '{32'h4280735f};
test_index[7532] = '{5};
test_input[60264:60271] = '{32'h42aa2f8f, 32'hc23bb933, 32'hc1a1c70b, 32'hc07caa7a, 32'h42bcbc1e, 32'h420242a3, 32'hc2684ee6, 32'hc16c5547};
test_output[7533] = '{32'h42bcbc1e};
test_index[7533] = '{4};
test_input[60272:60279] = '{32'hc223c4c8, 32'h3fb6d578, 32'h4283e81f, 32'hbe379f10, 32'hc25dd551, 32'hc13f748d, 32'hc1c08a5e, 32'h41bd1515};
test_output[7534] = '{32'h4283e81f};
test_index[7534] = '{2};
test_input[60280:60287] = '{32'hc1eb6adb, 32'hc27e3339, 32'h41aed304, 32'hc21b0989, 32'hc1c6aed4, 32'h40ea8ac7, 32'hc2139e2f, 32'hc1144d84};
test_output[7535] = '{32'h41aed304};
test_index[7535] = '{2};
test_input[60288:60295] = '{32'hc29f9e8b, 32'h41fae096, 32'hc1909425, 32'hc0a5b4c9, 32'h3e4cb1db, 32'h420fa68e, 32'h3ff32fe5, 32'hc002d4f4};
test_output[7536] = '{32'h420fa68e};
test_index[7536] = '{5};
test_input[60296:60303] = '{32'h413a2e27, 32'h426e9ffe, 32'h4212c9ea, 32'hc20665d0, 32'hc1a17896, 32'h42c66e2f, 32'h40e93466, 32'hc272fbf5};
test_output[7537] = '{32'h42c66e2f};
test_index[7537] = '{5};
test_input[60304:60311] = '{32'h4180f878, 32'h4297876b, 32'h40e1c8f2, 32'h413e6460, 32'hc202a829, 32'h4250f480, 32'h426a6676, 32'h4298ae3f};
test_output[7538] = '{32'h4298ae3f};
test_index[7538] = '{7};
test_input[60312:60319] = '{32'h427b2404, 32'hc2bedfcb, 32'hc2439cdc, 32'hc29412d2, 32'h42918719, 32'h429721e0, 32'hc28d739f, 32'hc232a483};
test_output[7539] = '{32'h429721e0};
test_index[7539] = '{5};
test_input[60320:60327] = '{32'hc1fbd03d, 32'hc160276a, 32'h4240d3ed, 32'hc1f3e20f, 32'h4289507d, 32'h42518ce7, 32'h3f6d72bb, 32'h42ab731f};
test_output[7540] = '{32'h42ab731f};
test_index[7540] = '{7};
test_input[60328:60335] = '{32'hc2c2055c, 32'hc02f15a7, 32'hc24bafab, 32'hc207afc3, 32'h4252de3e, 32'hc2a3bade, 32'h424643c6, 32'h42ad4a56};
test_output[7541] = '{32'h42ad4a56};
test_index[7541] = '{7};
test_input[60336:60343] = '{32'hc0f134dd, 32'hc1a5f875, 32'hc2150669, 32'hc26623c7, 32'h42ac0d30, 32'hc19ff9b9, 32'hc28e7f50, 32'h41dfb794};
test_output[7542] = '{32'h42ac0d30};
test_index[7542] = '{4};
test_input[60344:60351] = '{32'h4252e4b9, 32'h41838246, 32'hc281a3bc, 32'hc2183c45, 32'hc29849b6, 32'h42490ec2, 32'hc2bca3c7, 32'h42be11e0};
test_output[7543] = '{32'h42be11e0};
test_index[7543] = '{7};
test_input[60352:60359] = '{32'h41973b22, 32'h41d865be, 32'hc1bfa7b0, 32'h428b1b00, 32'h410673d5, 32'hc24f2a53, 32'h4254e21f, 32'h4207c94e};
test_output[7544] = '{32'h428b1b00};
test_index[7544] = '{3};
test_input[60360:60367] = '{32'h424f172c, 32'hc2a467c2, 32'hc299b2f8, 32'hc14f70dc, 32'hc2b33ac7, 32'h429ccd0f, 32'hc286ed53, 32'h41e1b536};
test_output[7545] = '{32'h429ccd0f};
test_index[7545] = '{5};
test_input[60368:60375] = '{32'h422bfe2f, 32'hc2a76bcf, 32'hc2a6e302, 32'h41533e80, 32'hc28d2fbe, 32'hc2c6f3dc, 32'hc2ac100b, 32'hc02f277e};
test_output[7546] = '{32'h422bfe2f};
test_index[7546] = '{0};
test_input[60376:60383] = '{32'h40799802, 32'h4265b245, 32'hc27d7555, 32'h426c0d5b, 32'hc2b52d34, 32'hc28ee3a9, 32'h42b72300, 32'h410eb849};
test_output[7547] = '{32'h42b72300};
test_index[7547] = '{6};
test_input[60384:60391] = '{32'hc23fa7ec, 32'hc244e371, 32'hc2a2b386, 32'h42807fe4, 32'h4262ee60, 32'h4292e6ce, 32'hc064b279, 32'hc2be654a};
test_output[7548] = '{32'h4292e6ce};
test_index[7548] = '{5};
test_input[60392:60399] = '{32'h42c42ae1, 32'hc2bf4c47, 32'hc157e7f7, 32'h41beb60a, 32'hc257dcd2, 32'hc25c5cdd, 32'h420df5dd, 32'hc27431e4};
test_output[7549] = '{32'h42c42ae1};
test_index[7549] = '{0};
test_input[60400:60407] = '{32'hc289838e, 32'h42a2acca, 32'hc213529d, 32'h415ad02f, 32'h4153d23e, 32'h41c656da, 32'h40e272cf, 32'h41ce7ffb};
test_output[7550] = '{32'h42a2acca};
test_index[7550] = '{1};
test_input[60408:60415] = '{32'h40caabd0, 32'h425b5144, 32'hc0e60c4a, 32'h420eb34d, 32'hc2852c77, 32'hc007b131, 32'h427f8c82, 32'h429622b5};
test_output[7551] = '{32'h429622b5};
test_index[7551] = '{7};
test_input[60416:60423] = '{32'h423c93e6, 32'h413a823f, 32'hc1b91f90, 32'hc1cf0b34, 32'hc2c1fdd1, 32'h3fb637cc, 32'h42b5f425, 32'hc2a0bfde};
test_output[7552] = '{32'h42b5f425};
test_index[7552] = '{6};
test_input[60424:60431] = '{32'h42c1928b, 32'hc1d6fc86, 32'hc29f7c96, 32'h42b1a320, 32'hc27f00f1, 32'hc21c1f76, 32'h4118a4b1, 32'h41ea5851};
test_output[7553] = '{32'h42c1928b};
test_index[7553] = '{0};
test_input[60432:60439] = '{32'h427a45ef, 32'h429e1389, 32'hc29d1e5e, 32'hc2694a0b, 32'h423c1a80, 32'h422af5d9, 32'h423dda1d, 32'h42b7d4f0};
test_output[7554] = '{32'h42b7d4f0};
test_index[7554] = '{7};
test_input[60440:60447] = '{32'h426b8b13, 32'hc2823681, 32'hc0cdc5ec, 32'hc21edf10, 32'h4252c5a6, 32'hc1894940, 32'h4210a569, 32'h4280ed54};
test_output[7555] = '{32'h4280ed54};
test_index[7555] = '{7};
test_input[60448:60455] = '{32'h40e3cd98, 32'hc0c5a4a9, 32'hc232c937, 32'hc2803770, 32'hc089ab94, 32'h4099cd6f, 32'h4166b36a, 32'hc2c2584b};
test_output[7556] = '{32'h4166b36a};
test_index[7556] = '{6};
test_input[60456:60463] = '{32'hc2894913, 32'hc237c29e, 32'h3ea317df, 32'h42ada1af, 32'hc288efb5, 32'hc2520773, 32'hc22e74e9, 32'h429047ba};
test_output[7557] = '{32'h42ada1af};
test_index[7557] = '{3};
test_input[60464:60471] = '{32'h42b606db, 32'hc25c52ff, 32'h426a2708, 32'h415b26a6, 32'hc21fa032, 32'h42ba3fa9, 32'h418a8c24, 32'h42831b36};
test_output[7558] = '{32'h42ba3fa9};
test_index[7558] = '{5};
test_input[60472:60479] = '{32'hc2374947, 32'hc22ad7e5, 32'h41dad186, 32'hc21fc1c2, 32'hc28e7538, 32'h41b65045, 32'h42973d05, 32'h4102b623};
test_output[7559] = '{32'h42973d05};
test_index[7559] = '{6};
test_input[60480:60487] = '{32'hc2a32795, 32'hc256ce6e, 32'hc288e002, 32'hc2971bc2, 32'h41c390cb, 32'hc29baad4, 32'hc153c227, 32'h42670ba6};
test_output[7560] = '{32'h42670ba6};
test_index[7560] = '{7};
test_input[60488:60495] = '{32'hc2b0a1f1, 32'hc28fb0a9, 32'h42a6ef93, 32'hc21bd10a, 32'h41f7c735, 32'hc1b327dc, 32'h421decd6, 32'h42089342};
test_output[7561] = '{32'h42a6ef93};
test_index[7561] = '{2};
test_input[60496:60503] = '{32'hc288469f, 32'hc1c2c448, 32'h41fa9e7a, 32'hc0f90e74, 32'h41aae5a2, 32'hc2b5fe9f, 32'hc15f8468, 32'h41798dc8};
test_output[7562] = '{32'h41fa9e7a};
test_index[7562] = '{2};
test_input[60504:60511] = '{32'h42ae13d2, 32'hc20dfd2f, 32'h4265daa8, 32'hc13f9907, 32'h42862133, 32'hc2357548, 32'hc24f2587, 32'hc20e2267};
test_output[7563] = '{32'h42ae13d2};
test_index[7563] = '{0};
test_input[60512:60519] = '{32'h42aebf6e, 32'h4263f1b6, 32'hc2576595, 32'h42577f17, 32'hc2b82fc2, 32'hbf018987, 32'hc2914306, 32'h41fc21be};
test_output[7564] = '{32'h42aebf6e};
test_index[7564] = '{0};
test_input[60520:60527] = '{32'hc11a0bd4, 32'hc0bc3058, 32'h4257ed49, 32'hc2ba064d, 32'hc128ee36, 32'h4143ce3b, 32'hc2125787, 32'h429f40eb};
test_output[7565] = '{32'h429f40eb};
test_index[7565] = '{7};
test_input[60528:60535] = '{32'h428c00fd, 32'hc0aa1586, 32'h42298288, 32'h4211d74e, 32'hc25df266, 32'h42b8c7d1, 32'h42be1ff0, 32'hc2c20d4b};
test_output[7566] = '{32'h42be1ff0};
test_index[7566] = '{6};
test_input[60536:60543] = '{32'h3f1737fe, 32'h3fb5c47b, 32'h40fc94a5, 32'h411626d2, 32'hc29d677b, 32'h4231a219, 32'hc1b434a2, 32'h419cdb9e};
test_output[7567] = '{32'h4231a219};
test_index[7567] = '{5};
test_input[60544:60551] = '{32'h40dff5d4, 32'hc2259a22, 32'h41c8fa1c, 32'hc27c921d, 32'hc0a8c845, 32'h42aac1a8, 32'h4262e962, 32'hc283d666};
test_output[7568] = '{32'h42aac1a8};
test_index[7568] = '{5};
test_input[60552:60559] = '{32'hc27a4423, 32'h42629ffc, 32'h42bcbcf8, 32'hc24f1445, 32'h42b88bf9, 32'hc0c56987, 32'h4243fb31, 32'h422cf744};
test_output[7569] = '{32'h42bcbcf8};
test_index[7569] = '{2};
test_input[60560:60567] = '{32'hc1ff2146, 32'h428a8d62, 32'hc20e198d, 32'h42c0ffed, 32'hc1763dba, 32'h426037cc, 32'hc2220fa2, 32'h424bdc42};
test_output[7570] = '{32'h42c0ffed};
test_index[7570] = '{3};
test_input[60568:60575] = '{32'hc1dbf112, 32'hc25f76c6, 32'h42741667, 32'hbfa5f671, 32'hc15df901, 32'hc28d9265, 32'hc27b8566, 32'hbfd728c4};
test_output[7571] = '{32'h42741667};
test_index[7571] = '{2};
test_input[60576:60583] = '{32'h42454790, 32'hc283c6ce, 32'hc269159e, 32'hc2a4b862, 32'hc2859cfa, 32'hc2b91f90, 32'hc2476e31, 32'hc29e3d04};
test_output[7572] = '{32'h42454790};
test_index[7572] = '{0};
test_input[60584:60591] = '{32'h42a8772e, 32'hc280a15a, 32'hc14bf4bb, 32'h428b0db8, 32'h42100bf9, 32'hc1d4b43e, 32'hc1050cb1, 32'h4274c1b6};
test_output[7573] = '{32'h42a8772e};
test_index[7573] = '{0};
test_input[60592:60599] = '{32'hc109a6bf, 32'h41678f25, 32'h4187f064, 32'h4281e326, 32'hc0e2a0ca, 32'hc2936d05, 32'h41924193, 32'hc2ab459d};
test_output[7574] = '{32'h4281e326};
test_index[7574] = '{3};
test_input[60600:60607] = '{32'hbf2e13b4, 32'h3f73b75c, 32'hc24c0474, 32'h41b76b6b, 32'h41a1d690, 32'h423294ed, 32'h42a97d1f, 32'h427c1807};
test_output[7575] = '{32'h42a97d1f};
test_index[7575] = '{6};
test_input[60608:60615] = '{32'hc1a40765, 32'hc1e671fd, 32'hc17f339a, 32'h42124396, 32'hc18c2346, 32'h419be18e, 32'h42b19025, 32'hc2b92d2b};
test_output[7576] = '{32'h42b19025};
test_index[7576] = '{6};
test_input[60616:60623] = '{32'h4287fca9, 32'hc2100535, 32'h42837b63, 32'hc2a76b8d, 32'h4241642e, 32'h424abf8c, 32'h42b5369f, 32'h42a6d0f6};
test_output[7577] = '{32'h42b5369f};
test_index[7577] = '{6};
test_input[60624:60631] = '{32'hc2bd76ff, 32'hc2368bb9, 32'hc2276b0f, 32'h42a41aef, 32'hbf0d7a2d, 32'h41f68f24, 32'hc2369f35, 32'hc2a6277d};
test_output[7578] = '{32'h42a41aef};
test_index[7578] = '{3};
test_input[60632:60639] = '{32'hc2b33b1c, 32'hc1bee596, 32'hc154a4a6, 32'h4289e418, 32'h429533b3, 32'h417c9f67, 32'hc10d06d9, 32'h429a230b};
test_output[7579] = '{32'h429a230b};
test_index[7579] = '{7};
test_input[60640:60647] = '{32'hc1358c54, 32'h40b13c8a, 32'hc1cf0f87, 32'hc2701a58, 32'h428ffeed, 32'hc28ed8ae, 32'hc2c0b09f, 32'h428ce458};
test_output[7580] = '{32'h428ffeed};
test_index[7580] = '{4};
test_input[60648:60655] = '{32'hc2938e5e, 32'hc29b29c4, 32'hc1c297e8, 32'hc1aae333, 32'hc2613eed, 32'h4249f207, 32'h418de818, 32'h424fb652};
test_output[7581] = '{32'h424fb652};
test_index[7581] = '{7};
test_input[60656:60663] = '{32'h42bd16ab, 32'hc29c09bd, 32'hc1f5b773, 32'h42659a82, 32'h42b350dd, 32'h424de944, 32'h41c5838b, 32'hc00d13c1};
test_output[7582] = '{32'h42bd16ab};
test_index[7582] = '{0};
test_input[60664:60671] = '{32'h42c60cb7, 32'hc2a55329, 32'h423a7445, 32'hc1fdc044, 32'h426b6e5e, 32'h42b43334, 32'h42801623, 32'h42019169};
test_output[7583] = '{32'h42c60cb7};
test_index[7583] = '{0};
test_input[60672:60679] = '{32'hc2a96535, 32'hc2a038ec, 32'hc07016fa, 32'h41cd7aa3, 32'hc2516663, 32'hc22e25f8, 32'hc2669066, 32'h428502e3};
test_output[7584] = '{32'h428502e3};
test_index[7584] = '{7};
test_input[60680:60687] = '{32'h42a69603, 32'h413421df, 32'hc2951b76, 32'hc20bed24, 32'h42285d29, 32'h40c8cb34, 32'h42897e8a, 32'hc21ab8e2};
test_output[7585] = '{32'h42a69603};
test_index[7585] = '{0};
test_input[60688:60695] = '{32'hc24e597b, 32'hc2b811e2, 32'hc25cd45f, 32'h41a37e0d, 32'hbfc722dc, 32'h42244e4d, 32'h42624818, 32'h42bcde05};
test_output[7586] = '{32'h42bcde05};
test_index[7586] = '{7};
test_input[60696:60703] = '{32'hc21e2d5a, 32'hc2c4d8ae, 32'h4297b3dd, 32'h40d3e4a2, 32'hc2850edc, 32'h40c53b38, 32'hc2b2dc95, 32'h429fe29c};
test_output[7587] = '{32'h429fe29c};
test_index[7587] = '{7};
test_input[60704:60711] = '{32'hc22a4a34, 32'h41aa24cd, 32'hc2c6630d, 32'hc2bb011c, 32'h42c20bd9, 32'h41fdf33e, 32'h42794667, 32'hc2b6a745};
test_output[7588] = '{32'h42c20bd9};
test_index[7588] = '{4};
test_input[60712:60719] = '{32'hbec80ba1, 32'h408d4fff, 32'h42ad0ceb, 32'h41ee08eb, 32'h42187d4e, 32'hc2c01976, 32'h42a4772e, 32'hc2bbe9fd};
test_output[7589] = '{32'h42ad0ceb};
test_index[7589] = '{2};
test_input[60720:60727] = '{32'h418397d0, 32'hc2bd7e4e, 32'hc260407d, 32'hc230db72, 32'h429571b4, 32'h42b02c9a, 32'hc2346ee4, 32'hc0d2b66f};
test_output[7590] = '{32'h42b02c9a};
test_index[7590] = '{5};
test_input[60728:60735] = '{32'hc2424705, 32'h42255e29, 32'h42507318, 32'h421c0b9a, 32'h41226f31, 32'hc2888fe5, 32'hc29e816d, 32'hc28b6c6a};
test_output[7591] = '{32'h42507318};
test_index[7591] = '{2};
test_input[60736:60743] = '{32'h42c7bc72, 32'hc20dc597, 32'h422c5a4e, 32'hc1de10a9, 32'hc2013fa9, 32'h42be4472, 32'h41f962f6, 32'hc1ac9bff};
test_output[7592] = '{32'h42c7bc72};
test_index[7592] = '{0};
test_input[60744:60751] = '{32'h423fbb64, 32'hc08a0ebb, 32'h42346102, 32'h42b7b1a6, 32'h41ae46fe, 32'hc265b9f2, 32'h420b5e1a, 32'h425f8108};
test_output[7593] = '{32'h42b7b1a6};
test_index[7593] = '{3};
test_input[60752:60759] = '{32'h4216361b, 32'hc2c07ed0, 32'hc17fdb13, 32'hc1d3e588, 32'hc002d6b0, 32'h4260a3fd, 32'hc0f3cde4, 32'h41cddc32};
test_output[7594] = '{32'h4260a3fd};
test_index[7594] = '{5};
test_input[60760:60767] = '{32'h41968637, 32'h4239b8e2, 32'h420984dc, 32'hc24191fd, 32'h424aa457, 32'h42652aa9, 32'hc2367961, 32'h415de607};
test_output[7595] = '{32'h42652aa9};
test_index[7595] = '{5};
test_input[60768:60775] = '{32'hc1b7bf8e, 32'hc2b2069a, 32'h42881e25, 32'h42a97e52, 32'h42425b63, 32'hc27a9fec, 32'hc2253e62, 32'h421d3744};
test_output[7596] = '{32'h42a97e52};
test_index[7596] = '{3};
test_input[60776:60783] = '{32'h3fa23248, 32'h42387e42, 32'hc2441649, 32'hc0fe0bff, 32'hc24e295d, 32'h41972059, 32'h42a47a95, 32'h41b63243};
test_output[7597] = '{32'h42a47a95};
test_index[7597] = '{6};
test_input[60784:60791] = '{32'h420a4bc9, 32'hc266a23b, 32'h427abb8e, 32'hc2a32acf, 32'h42af7e89, 32'hc22e3d5e, 32'hc2370b22, 32'h423cf3ab};
test_output[7598] = '{32'h42af7e89};
test_index[7598] = '{4};
test_input[60792:60799] = '{32'h42373b47, 32'h41531f2e, 32'hc2b9e08b, 32'hc13b22f9, 32'h421dad24, 32'h40cf7bf2, 32'hc13e6777, 32'hc29eac1a};
test_output[7599] = '{32'h42373b47};
test_index[7599] = '{0};
test_input[60800:60807] = '{32'h41078a24, 32'hc2965b87, 32'h428e27db, 32'h41daabb2, 32'hc2122448, 32'h429c96d3, 32'h428859cd, 32'h42b13d3f};
test_output[7600] = '{32'h42b13d3f};
test_index[7600] = '{7};
test_input[60808:60815] = '{32'h416f382e, 32'h4150e9e2, 32'h42b2929e, 32'hc21903f2, 32'h42563e3a, 32'h42bcdd59, 32'hc2937f86, 32'hc2b68216};
test_output[7601] = '{32'h42bcdd59};
test_index[7601] = '{5};
test_input[60816:60823] = '{32'h3fe9d41c, 32'hc14f6b69, 32'hc2b35515, 32'hc1a9db82, 32'h41f6da63, 32'h428baead, 32'h423ebacb, 32'h428fb0ea};
test_output[7602] = '{32'h428fb0ea};
test_index[7602] = '{7};
test_input[60824:60831] = '{32'h42ae5912, 32'h42bc311b, 32'hc2c604f5, 32'hc255ae43, 32'h409f453a, 32'hc0a42f62, 32'hc2a621e7, 32'hc27ab3e9};
test_output[7603] = '{32'h42bc311b};
test_index[7603] = '{1};
test_input[60832:60839] = '{32'hc28f05d2, 32'hc2bd8e07, 32'h424ae9d5, 32'h41237c4a, 32'hc26d2a56, 32'h42920065, 32'hc2785494, 32'hc2bfc03e};
test_output[7604] = '{32'h42920065};
test_index[7604] = '{5};
test_input[60840:60847] = '{32'h41ae6421, 32'hc23ec73c, 32'h4047fa08, 32'hc2ace141, 32'h42b21bac, 32'hc1baeeaa, 32'hc2632ebf, 32'h42761b1a};
test_output[7605] = '{32'h42b21bac};
test_index[7605] = '{4};
test_input[60848:60855] = '{32'h42976083, 32'h41b256b0, 32'hc2b4ce5b, 32'hc1ee33e2, 32'h41ccab8c, 32'h42a48544, 32'h424d033b, 32'hc0ba4643};
test_output[7606] = '{32'h42a48544};
test_index[7606] = '{5};
test_input[60856:60863] = '{32'h42149723, 32'hc2a6480e, 32'hc2225a66, 32'hc1f86079, 32'h40fc6146, 32'hc246c570, 32'hc24bf8b7, 32'h42361ed6};
test_output[7607] = '{32'h42361ed6};
test_index[7607] = '{7};
test_input[60864:60871] = '{32'h423927f8, 32'h42123a09, 32'h420a1b62, 32'h425d4de0, 32'hc20f21e2, 32'hbfb34b47, 32'h42c74a44, 32'hc1b2951b};
test_output[7608] = '{32'h42c74a44};
test_index[7608] = '{6};
test_input[60872:60879] = '{32'h426b4049, 32'hc2a1242f, 32'hc2a19460, 32'hc235e908, 32'h424ac35e, 32'h42a05087, 32'h409a7d81, 32'h425262dc};
test_output[7609] = '{32'h42a05087};
test_index[7609] = '{5};
test_input[60880:60887] = '{32'hc29d6e81, 32'hc230f124, 32'h424aa317, 32'hc1fd592c, 32'hc29d63d4, 32'hc2a76f43, 32'hc20a4953, 32'h42a489e5};
test_output[7610] = '{32'h42a489e5};
test_index[7610] = '{7};
test_input[60888:60895] = '{32'h42790e9a, 32'h427ef8a9, 32'h426e995a, 32'hc1502a6a, 32'h40ac6e96, 32'h426868f7, 32'h42baaf8d, 32'h424279fc};
test_output[7611] = '{32'h42baaf8d};
test_index[7611] = '{6};
test_input[60896:60903] = '{32'h421ce70f, 32'h403b47bf, 32'hc2116276, 32'h42a434ed, 32'h42aa2046, 32'hc2a0dff9, 32'h41f1c933, 32'h41158437};
test_output[7612] = '{32'h42aa2046};
test_index[7612] = '{4};
test_input[60904:60911] = '{32'h42a19553, 32'h41f2a813, 32'hc253769c, 32'h42aa597e, 32'hc2ae3e98, 32'h42867b96, 32'hc225b40e, 32'hc217993c};
test_output[7613] = '{32'h42aa597e};
test_index[7613] = '{3};
test_input[60912:60919] = '{32'h41ef6053, 32'h42c66ce6, 32'hc284c91e, 32'hc16d990b, 32'hc130e38e, 32'hc1f4c7c2, 32'h4251ef90, 32'hc2bfa3f8};
test_output[7614] = '{32'h42c66ce6};
test_index[7614] = '{1};
test_input[60920:60927] = '{32'h42bd2422, 32'hc290773b, 32'h41e66a51, 32'h42529a65, 32'hc2104d24, 32'hc283060f, 32'hc1b3f312, 32'hc190b2e9};
test_output[7615] = '{32'h42bd2422};
test_index[7615] = '{0};
test_input[60928:60935] = '{32'hc2183a82, 32'h42a2c372, 32'h42b29f17, 32'hc1bf6801, 32'h40bf3511, 32'hc10972b1, 32'hc2b17d9a, 32'hc2c3aa04};
test_output[7616] = '{32'h42b29f17};
test_index[7616] = '{2};
test_input[60936:60943] = '{32'hc24d0bcb, 32'hc2054a00, 32'h41f6dcfe, 32'hc2077658, 32'h41865adf, 32'h42ad9427, 32'h418aec7c, 32'hc22ab41b};
test_output[7617] = '{32'h42ad9427};
test_index[7617] = '{5};
test_input[60944:60951] = '{32'hc29f8587, 32'h42620e9a, 32'h418c97dc, 32'hc18d86a7, 32'hc2492396, 32'h41d9658a, 32'h4267d209, 32'hc1ba2264};
test_output[7618] = '{32'h4267d209};
test_index[7618] = '{6};
test_input[60952:60959] = '{32'hc2b7ecdb, 32'h41df37f6, 32'hc23f7269, 32'h41f0898d, 32'h4267f1fc, 32'h42a033e8, 32'h41815a74, 32'h3f841966};
test_output[7619] = '{32'h42a033e8};
test_index[7619] = '{5};
test_input[60960:60967] = '{32'hc288dcfa, 32'h429e8710, 32'h425b806b, 32'hc1766f77, 32'hc1f44eff, 32'hc2840651, 32'h41d5efa7, 32'h41ca69d5};
test_output[7620] = '{32'h429e8710};
test_index[7620] = '{1};
test_input[60968:60975] = '{32'h42ac817a, 32'hc0c3d2d0, 32'hc2a78387, 32'hc29ac2bd, 32'h4206ff8a, 32'h42a0caca, 32'h429ca57e, 32'hc1daa692};
test_output[7621] = '{32'h42ac817a};
test_index[7621] = '{0};
test_input[60976:60983] = '{32'hc2b4b3ca, 32'h429918b8, 32'h421bff92, 32'hc0e23670, 32'hc1fc8fc0, 32'h42aabe63, 32'h42a120ba, 32'h42ac1a50};
test_output[7622] = '{32'h42ac1a50};
test_index[7622] = '{7};
test_input[60984:60991] = '{32'h420aeef7, 32'h42a51e3c, 32'hc28f4482, 32'hc0189373, 32'h42a2fea7, 32'h424d94d5, 32'h42a4257c, 32'hc129e68d};
test_output[7623] = '{32'h42a51e3c};
test_index[7623] = '{1};
test_input[60992:60999] = '{32'h4299c004, 32'hc22af757, 32'h410f4e69, 32'h41a3ba92, 32'hc2ac0216, 32'h42835bd4, 32'h42693ca3, 32'hc23c8b8e};
test_output[7624] = '{32'h4299c004};
test_index[7624] = '{0};
test_input[61000:61007] = '{32'hc292f0ec, 32'hc2a41431, 32'hc1142028, 32'h42c42f59, 32'h429ed9e7, 32'h409850ba, 32'h42bb1bcd, 32'h42098610};
test_output[7625] = '{32'h42c42f59};
test_index[7625] = '{3};
test_input[61008:61015] = '{32'h42bb85fa, 32'hc218b49f, 32'h415aa1e9, 32'hc28b135e, 32'h42baad78, 32'hc21b3b6e, 32'hc1896843, 32'h429e6a1c};
test_output[7626] = '{32'h42bb85fa};
test_index[7626] = '{0};
test_input[61016:61023] = '{32'h429b7f29, 32'hc27d7291, 32'hc102d0fe, 32'h418ca45a, 32'h41a8c73d, 32'hc232c672, 32'hc17fd1e2, 32'hc1126178};
test_output[7627] = '{32'h429b7f29};
test_index[7627] = '{0};
test_input[61024:61031] = '{32'hc2a9e375, 32'hc2880563, 32'hc25a2279, 32'hc29ddf3d, 32'hc2c585f0, 32'hc022982a, 32'hc1f41fb7, 32'hc214ed9e};
test_output[7628] = '{32'hc022982a};
test_index[7628] = '{5};
test_input[61032:61039] = '{32'h40d5125a, 32'hc234eb8a, 32'hc2c06a6e, 32'h4204fb46, 32'hc2044d0c, 32'hc2ba02b6, 32'h423c9957, 32'h4191d6d6};
test_output[7629] = '{32'h423c9957};
test_index[7629] = '{6};
test_input[61040:61047] = '{32'h41e69e7d, 32'hc2c05548, 32'hc123d175, 32'h4281fb8b, 32'h421b53f1, 32'h4291fc5e, 32'hc278977f, 32'hc1b5cdc4};
test_output[7630] = '{32'h4291fc5e};
test_index[7630] = '{5};
test_input[61048:61055] = '{32'h42b1a703, 32'h4281ae6e, 32'hc2800f40, 32'h41a38b24, 32'hc2ac0799, 32'hc2bd91f3, 32'h42670bfb, 32'h425d7109};
test_output[7631] = '{32'h42b1a703};
test_index[7631] = '{0};
test_input[61056:61063] = '{32'hc2be965a, 32'hc1d64c03, 32'h42b2ea98, 32'h417bccd9, 32'hc1d29019, 32'hc2900025, 32'hc2322fb3, 32'hc214fbb9};
test_output[7632] = '{32'h42b2ea98};
test_index[7632] = '{2};
test_input[61064:61071] = '{32'hc2aee2ba, 32'h4234a284, 32'hc210cbdb, 32'h4221369f, 32'hc11ea76d, 32'h4280efb8, 32'h4191d8c4, 32'h42c7aeda};
test_output[7633] = '{32'h42c7aeda};
test_index[7633] = '{7};
test_input[61072:61079] = '{32'h41a49157, 32'h42b57a31, 32'hc1b42d8e, 32'h42363195, 32'h42829945, 32'h42a56fe1, 32'hc292e635, 32'hc29e06c0};
test_output[7634] = '{32'h42b57a31};
test_index[7634] = '{1};
test_input[61080:61087] = '{32'h40c117f7, 32'h423d9ba4, 32'hc282e309, 32'h41b296f3, 32'hc28fa717, 32'hc12fc2a5, 32'hc283c4b5, 32'h419288c1};
test_output[7635] = '{32'h423d9ba4};
test_index[7635] = '{1};
test_input[61088:61095] = '{32'h422d43ce, 32'h42c0bf97, 32'h42a674ee, 32'h421526b2, 32'hc0d3cba7, 32'h415b8661, 32'h4283d50d, 32'h42aedf73};
test_output[7636] = '{32'h42c0bf97};
test_index[7636] = '{1};
test_input[61096:61103] = '{32'hc299ba6e, 32'hc2a93fd0, 32'h413cedfa, 32'h4216f064, 32'h42390748, 32'hc2c13645, 32'h41f7f8b9, 32'hc0ffc1a7};
test_output[7637] = '{32'h42390748};
test_index[7637] = '{4};
test_input[61104:61111] = '{32'hc211f925, 32'h42a70ebd, 32'hbf761f98, 32'h42108292, 32'hc2b4de08, 32'h41debb16, 32'h411b4bb0, 32'h41b980cc};
test_output[7638] = '{32'h42a70ebd};
test_index[7638] = '{1};
test_input[61112:61119] = '{32'h411a143a, 32'hc115eddc, 32'h42b6f438, 32'hc29911c9, 32'hbf7d3b7d, 32'h425fce0f, 32'hc28e305b, 32'h4294b408};
test_output[7639] = '{32'h42b6f438};
test_index[7639] = '{2};
test_input[61120:61127] = '{32'h41cc95bd, 32'h42b7161d, 32'h429db9af, 32'hc272f860, 32'hc2164391, 32'h4215f9a3, 32'hc198f1c0, 32'h424b25b6};
test_output[7640] = '{32'h42b7161d};
test_index[7640] = '{1};
test_input[61128:61135] = '{32'hc19c5579, 32'h40ac7b16, 32'hc1cde8b9, 32'hc20015b6, 32'hc1c2d03e, 32'hc26ae878, 32'h41979bac, 32'hc2b6b1ac};
test_output[7641] = '{32'h41979bac};
test_index[7641] = '{6};
test_input[61136:61143] = '{32'hc2912fed, 32'hc23c5b1c, 32'h42a5f331, 32'h41f96e46, 32'hc26076ca, 32'hc2125227, 32'hc2b6c83f, 32'h41516804};
test_output[7642] = '{32'h42a5f331};
test_index[7642] = '{2};
test_input[61144:61151] = '{32'h41a07545, 32'h42c0b67f, 32'h42748e67, 32'h428d337d, 32'h428fe40f, 32'hc1f06a2a, 32'h42196e6f, 32'hbf24020d};
test_output[7643] = '{32'h42c0b67f};
test_index[7643] = '{1};
test_input[61152:61159] = '{32'hc0c279be, 32'h4205da54, 32'hc27b8d0a, 32'h42a34119, 32'hc21ba538, 32'h41dc7713, 32'h429516a5, 32'hc1c2f296};
test_output[7644] = '{32'h42a34119};
test_index[7644] = '{3};
test_input[61160:61167] = '{32'h428eea2e, 32'hc2104206, 32'h41a3ae3b, 32'hc23a7600, 32'hc273b758, 32'hc2672e90, 32'hc1d33c53, 32'hc2624af6};
test_output[7645] = '{32'h428eea2e};
test_index[7645] = '{0};
test_input[61168:61175] = '{32'h42651af7, 32'h424955bf, 32'h40fe2963, 32'hc296cb81, 32'hc284fccc, 32'h40a4c824, 32'h41f05baf, 32'h421a7758};
test_output[7646] = '{32'h42651af7};
test_index[7646] = '{0};
test_input[61176:61183] = '{32'hc2b805ed, 32'hc1f31978, 32'h41df9967, 32'hc2203665, 32'h419fffa0, 32'hc2a633ff, 32'hc239063c, 32'h4195741d};
test_output[7647] = '{32'h41df9967};
test_index[7647] = '{2};
test_input[61184:61191] = '{32'hc19d9958, 32'hc2890ae6, 32'h42b03f6b, 32'hc27d2b24, 32'hc06c27ce, 32'hc24dd7c3, 32'h42931a25, 32'hc1d67fd1};
test_output[7648] = '{32'h42b03f6b};
test_index[7648] = '{2};
test_input[61192:61199] = '{32'hc2b037ca, 32'h42515a67, 32'h4298a628, 32'h41f2fa8d, 32'h429b5d9a, 32'hc2944b93, 32'hc2c1d747, 32'h42980f26};
test_output[7649] = '{32'h429b5d9a};
test_index[7649] = '{4};
test_input[61200:61207] = '{32'h4214ebd3, 32'h427d04f1, 32'hc2b49541, 32'hc240b319, 32'h428820ff, 32'hc2275f30, 32'hbf729371, 32'h4284847e};
test_output[7650] = '{32'h428820ff};
test_index[7650] = '{4};
test_input[61208:61215] = '{32'h42699162, 32'h42844a93, 32'hc20cbd8e, 32'h41c5c9e6, 32'hc2c7ae60, 32'hc20a704e, 32'h42936cfa, 32'h41859655};
test_output[7651] = '{32'h42936cfa};
test_index[7651] = '{6};
test_input[61216:61223] = '{32'hc2b68177, 32'hc1bf6aab, 32'hc080ba12, 32'h41e4ac90, 32'h42a6eb99, 32'h429952da, 32'h41a27c82, 32'hc281dfb2};
test_output[7652] = '{32'h42a6eb99};
test_index[7652] = '{4};
test_input[61224:61231] = '{32'h42b68a75, 32'h42afd003, 32'h42a3337f, 32'hc2a543b1, 32'hc2bd73e7, 32'hc2c0a4ef, 32'h40c7aac7, 32'hc279b35a};
test_output[7653] = '{32'h42b68a75};
test_index[7653] = '{0};
test_input[61232:61239] = '{32'hc1241792, 32'hc29cae91, 32'hc2814e6b, 32'h4193e671, 32'hc1e3cd8e, 32'h41a49780, 32'hc234e341, 32'hc2c707c1};
test_output[7654] = '{32'h41a49780};
test_index[7654] = '{5};
test_input[61240:61247] = '{32'hc21cac86, 32'h422906f4, 32'hc184f8bb, 32'hc2a6b038, 32'hc276292f, 32'h42a57f68, 32'h42b02b8e, 32'hc2405858};
test_output[7655] = '{32'h42b02b8e};
test_index[7655] = '{6};
test_input[61248:61255] = '{32'hc2a68547, 32'h4296e401, 32'hc218f067, 32'hc2bea3d3, 32'hc14f650b, 32'h4261bc31, 32'h429a1c0d, 32'h407e98f1};
test_output[7656] = '{32'h429a1c0d};
test_index[7656] = '{6};
test_input[61256:61263] = '{32'hc25269e9, 32'hc13d5b1b, 32'hc241c92b, 32'h427558b0, 32'h42c078aa, 32'hc26fc66b, 32'hc23e0e56, 32'hc2c0cb4d};
test_output[7657] = '{32'h42c078aa};
test_index[7657] = '{4};
test_input[61264:61271] = '{32'h421585ba, 32'hc28df864, 32'hc2afdedd, 32'h41ce92aa, 32'hc2b34ae7, 32'h42af12ed, 32'hc24a50ce, 32'hc286d504};
test_output[7658] = '{32'h42af12ed};
test_index[7658] = '{5};
test_input[61272:61279] = '{32'h429226f1, 32'hc2bef391, 32'hc1275ac0, 32'h42920fad, 32'hc2165cb9, 32'h426e01d7, 32'hc2411fe9, 32'hc2502e09};
test_output[7659] = '{32'h429226f1};
test_index[7659] = '{0};
test_input[61280:61287] = '{32'h3f37980b, 32'hc2a26b56, 32'h41149ecd, 32'hc2908eb2, 32'h41ed9fa4, 32'hc27266af, 32'hc2934c15, 32'hc2b6b4ee};
test_output[7660] = '{32'h41ed9fa4};
test_index[7660] = '{4};
test_input[61288:61295] = '{32'h4202fd20, 32'h41cc435d, 32'hc1228b11, 32'hc25222f4, 32'h42ba9b0c, 32'hc286a86d, 32'h420cf0a0, 32'hc2364e00};
test_output[7661] = '{32'h42ba9b0c};
test_index[7661] = '{4};
test_input[61296:61303] = '{32'h42af6f90, 32'h415ea1ff, 32'h420b5bd1, 32'h42a16e3b, 32'hc287d593, 32'h41e1b8c1, 32'hc1c50b02, 32'hc1ad4fe4};
test_output[7662] = '{32'h42af6f90};
test_index[7662] = '{0};
test_input[61304:61311] = '{32'h428d70e3, 32'hc299bd48, 32'hc2964668, 32'h420dc1eb, 32'h4271802f, 32'h42b964b7, 32'hc1f0ae7e, 32'h428a49c4};
test_output[7663] = '{32'h42b964b7};
test_index[7663] = '{5};
test_input[61312:61319] = '{32'hc2386ba8, 32'hc1cc3e88, 32'hc0fb8ed9, 32'hc2ac9161, 32'h41b326ff, 32'h427bd2d3, 32'h425c44eb, 32'hc20977ad};
test_output[7664] = '{32'h427bd2d3};
test_index[7664] = '{5};
test_input[61320:61327] = '{32'hc23ce417, 32'hc28f27d0, 32'hc19dd6a3, 32'h42961e10, 32'hc1b5300f, 32'hc1aae1b6, 32'h423c5584, 32'h429cb4c2};
test_output[7665] = '{32'h429cb4c2};
test_index[7665] = '{7};
test_input[61328:61335] = '{32'hc24c1e10, 32'h425495c6, 32'hc239be9b, 32'h42c2ca06, 32'hc29d1573, 32'hc1d20a43, 32'hc2205321, 32'h41998098};
test_output[7666] = '{32'h42c2ca06};
test_index[7666] = '{3};
test_input[61336:61343] = '{32'hc03e9440, 32'hc2bdcba8, 32'hc23a495d, 32'h4284929f, 32'hc28022bd, 32'h412cc99a, 32'hc1badb4b, 32'h41b8f44c};
test_output[7667] = '{32'h4284929f};
test_index[7667] = '{3};
test_input[61344:61351] = '{32'h4130e2c9, 32'h4295276c, 32'h423623be, 32'hc1132ce4, 32'h42c31e19, 32'h41326e69, 32'h4149db5a, 32'h41ec96ee};
test_output[7668] = '{32'h42c31e19};
test_index[7668] = '{4};
test_input[61352:61359] = '{32'hc1d1e35e, 32'hc2c112f9, 32'hc2823104, 32'hc29b686a, 32'h408e63dd, 32'hc2887ea7, 32'h3f9c73be, 32'hc20f97e7};
test_output[7669] = '{32'h408e63dd};
test_index[7669] = '{4};
test_input[61360:61367] = '{32'h421f4318, 32'hc25e00ea, 32'h4105ff37, 32'hc235088b, 32'h42911d54, 32'hc285c4aa, 32'hc278dc2a, 32'hc11d42a7};
test_output[7670] = '{32'h42911d54};
test_index[7670] = '{4};
test_input[61368:61375] = '{32'h42875329, 32'hc19f1479, 32'hc211177b, 32'hc2232b2d, 32'hc2991822, 32'h42b262ae, 32'hc2a8e293, 32'h42a3e974};
test_output[7671] = '{32'h42b262ae};
test_index[7671] = '{5};
test_input[61376:61383] = '{32'hc269b742, 32'hc254e913, 32'h42845a38, 32'hc2a86405, 32'hc2ae5685, 32'hc2235724, 32'h4251abf4, 32'h4297d0bc};
test_output[7672] = '{32'h4297d0bc};
test_index[7672] = '{7};
test_input[61384:61391] = '{32'hc29f2636, 32'h411a2189, 32'h428b2f88, 32'hc26477ef, 32'hc08c6493, 32'hc246a82c, 32'h426e75d8, 32'hc1f9c38f};
test_output[7673] = '{32'h428b2f88};
test_index[7673] = '{2};
test_input[61392:61399] = '{32'hc2c019f2, 32'hc28e2fcd, 32'hc1f0d6b3, 32'h41b66a5c, 32'h4209478b, 32'hc298ac76, 32'hc2a5e4bd, 32'h4229cded};
test_output[7674] = '{32'h4229cded};
test_index[7674] = '{7};
test_input[61400:61407] = '{32'hc19ce9e7, 32'h419b9855, 32'h42609312, 32'h40322133, 32'hc2615c7d, 32'hc21374cd, 32'h41e06d1d, 32'h42128358};
test_output[7675] = '{32'h42609312};
test_index[7675] = '{2};
test_input[61408:61415] = '{32'h42276b1f, 32'hc28670a8, 32'h40f59f1a, 32'hc2a773e8, 32'h409b20a5, 32'h42bf96ae, 32'hc2c4e063, 32'h418e8303};
test_output[7676] = '{32'h42bf96ae};
test_index[7676] = '{5};
test_input[61416:61423] = '{32'hc16a1b98, 32'h4120104b, 32'h4222a454, 32'hc2b7fbf6, 32'hc1935a79, 32'hc2721b64, 32'hc2a5cf3f, 32'h4249ad9f};
test_output[7677] = '{32'h4249ad9f};
test_index[7677] = '{7};
test_input[61424:61431] = '{32'hc1c88dd0, 32'h410d5398, 32'h42754b15, 32'h42c7141a, 32'h402289a6, 32'h426d2567, 32'hc21a5a25, 32'h420efcd9};
test_output[7678] = '{32'h42c7141a};
test_index[7678] = '{3};
test_input[61432:61439] = '{32'hc2935e7d, 32'h427665e7, 32'hc10431a2, 32'h429a8911, 32'h42800ac9, 32'h41ad1291, 32'hc2937738, 32'h42a8402e};
test_output[7679] = '{32'h42a8402e};
test_index[7679] = '{7};
test_input[61440:61447] = '{32'hc289a121, 32'h42a9771d, 32'hc2844520, 32'hc2135f55, 32'h40df1f9e, 32'h41eae20c, 32'hc1e55343, 32'hc1bd191b};
test_output[7680] = '{32'h42a9771d};
test_index[7680] = '{1};
test_input[61448:61455] = '{32'hc296c240, 32'h42c3a60b, 32'h4210c374, 32'h4208ddd7, 32'hbf87912f, 32'hc2b6a084, 32'hc1e9d649, 32'hc16ef3b8};
test_output[7681] = '{32'h42c3a60b};
test_index[7681] = '{1};
test_input[61456:61463] = '{32'hc186158a, 32'h42a90177, 32'hc2a4a65f, 32'h4184e9b4, 32'h415c5e4e, 32'hc1d1290c, 32'hc22a645b, 32'hc2c3b9e3};
test_output[7682] = '{32'h42a90177};
test_index[7682] = '{1};
test_input[61464:61471] = '{32'h41c4a3db, 32'h42a5a317, 32'hc2a2bbdc, 32'hc298d60d, 32'h42294194, 32'hc2148f62, 32'hc2298118, 32'hc2b1f06f};
test_output[7683] = '{32'h42a5a317};
test_index[7683] = '{1};
test_input[61472:61479] = '{32'h41d6a04a, 32'h42c1c4d1, 32'h42aeabd7, 32'hc1279a3d, 32'h41a7eae2, 32'hc25b1776, 32'h41ff147d, 32'hc23255f7};
test_output[7684] = '{32'h42c1c4d1};
test_index[7684] = '{1};
test_input[61480:61487] = '{32'hc118bb80, 32'hc1a6f7fe, 32'h4253a47e, 32'h422f1de0, 32'hc269c2ab, 32'hc0bc6e96, 32'h42bac835, 32'h4220ba92};
test_output[7685] = '{32'h42bac835};
test_index[7685] = '{6};
test_input[61488:61495] = '{32'hc2a548c1, 32'hc299b093, 32'h426c5c72, 32'h42b4be2a, 32'h419fa960, 32'h42b470a7, 32'h426e746d, 32'hc1eb00e8};
test_output[7686] = '{32'h42b4be2a};
test_index[7686] = '{3};
test_input[61496:61503] = '{32'hc23bb457, 32'hc204f8ea, 32'hc27345a2, 32'h4246da40, 32'h4252d009, 32'h42bab509, 32'hc2c2d459, 32'hc1ab6bf3};
test_output[7687] = '{32'h42bab509};
test_index[7687] = '{5};
test_input[61504:61511] = '{32'h419d2a5f, 32'h429f91bb, 32'hc187b11f, 32'h41482d49, 32'hc2a31d43, 32'h40d1fcb3, 32'h428cd08b, 32'h400c14f0};
test_output[7688] = '{32'h429f91bb};
test_index[7688] = '{1};
test_input[61512:61519] = '{32'h42126c43, 32'h420cced7, 32'hc2a5458e, 32'h42997a0f, 32'h429f0ee7, 32'h4159531d, 32'h424a6a35, 32'hc2ab8560};
test_output[7689] = '{32'h429f0ee7};
test_index[7689] = '{4};
test_input[61520:61527] = '{32'hc28d5e29, 32'h42ad6b1e, 32'hc282fdfd, 32'hc2c48167, 32'h4283ab7e, 32'hc1654bd5, 32'h41eb1134, 32'h4226b910};
test_output[7690] = '{32'h42ad6b1e};
test_index[7690] = '{1};
test_input[61528:61535] = '{32'hc203ff7d, 32'h428154c6, 32'hc24a92e8, 32'h4278d82d, 32'h42825b1b, 32'h41ecd849, 32'h41d61b50, 32'hc246bb58};
test_output[7691] = '{32'h42825b1b};
test_index[7691] = '{4};
test_input[61536:61543] = '{32'hc2aed3a5, 32'h4290c1fb, 32'h411bf304, 32'hc2ad9d2c, 32'hc25d8e66, 32'hc15f3ea6, 32'hc182a4af, 32'hc29c7df4};
test_output[7692] = '{32'h4290c1fb};
test_index[7692] = '{1};
test_input[61544:61551] = '{32'hc24bed8b, 32'h4280bec8, 32'hc24cc5b1, 32'hc2376dd7, 32'h4275d59e, 32'h41a19c8e, 32'hc245773e, 32'hc28fea0e};
test_output[7693] = '{32'h4280bec8};
test_index[7693] = '{1};
test_input[61552:61559] = '{32'hc1ce35b1, 32'hc17a1f55, 32'h41ca0b90, 32'hc2c23065, 32'hc2c651e3, 32'h42b4ae74, 32'hc26e08c3, 32'h42b815b9};
test_output[7694] = '{32'h42b815b9};
test_index[7694] = '{7};
test_input[61560:61567] = '{32'hc2a19f7b, 32'h418659a5, 32'hc2a01f89, 32'h4244600a, 32'h4103a403, 32'hc2b70f5e, 32'h4117cb64, 32'hc294040d};
test_output[7695] = '{32'h4244600a};
test_index[7695] = '{3};
test_input[61568:61575] = '{32'h41dfb714, 32'h42a8c64b, 32'h421e0db4, 32'hc2b22054, 32'h42c1fd76, 32'hc2c18f3c, 32'hc266b469, 32'h424c354c};
test_output[7696] = '{32'h42c1fd76};
test_index[7696] = '{4};
test_input[61576:61583] = '{32'hc2173987, 32'hc2955212, 32'h4288f420, 32'hc0c9833b, 32'h42098d3d, 32'h4180d8d6, 32'hc1a51ea4, 32'hc1cc091f};
test_output[7697] = '{32'h4288f420};
test_index[7697] = '{2};
test_input[61584:61591] = '{32'h423effa0, 32'h426c62d0, 32'hc2a04845, 32'hc152cc2a, 32'h41920448, 32'h4281fdf9, 32'h42702b78, 32'h42431331};
test_output[7698] = '{32'h4281fdf9};
test_index[7698] = '{5};
test_input[61592:61599] = '{32'hc04f772b, 32'hc260fd59, 32'hc1c71cad, 32'h42c20d74, 32'hc250725c, 32'hc2c0e94a, 32'h42285121, 32'h41951d8b};
test_output[7699] = '{32'h42c20d74};
test_index[7699] = '{3};
test_input[61600:61607] = '{32'h4298b984, 32'h3fb73276, 32'hc28666e9, 32'h42506d5d, 32'hc2b821d9, 32'h425c037d, 32'hc28958e7, 32'hc2c41b3c};
test_output[7700] = '{32'h4298b984};
test_index[7700] = '{0};
test_input[61608:61615] = '{32'h4238f07e, 32'h404a4156, 32'hc23355b3, 32'h4115f443, 32'h41dd3c13, 32'hc1354104, 32'hc2810f02, 32'hc2a5bc2b};
test_output[7701] = '{32'h4238f07e};
test_index[7701] = '{0};
test_input[61616:61623] = '{32'h4218130a, 32'hc2971c8c, 32'hc1a06ec1, 32'h42ab673b, 32'h422437bc, 32'h429468c6, 32'h40d20c86, 32'h41bf43fe};
test_output[7702] = '{32'h42ab673b};
test_index[7702] = '{3};
test_input[61624:61631] = '{32'hc2881d67, 32'h421f8906, 32'h4282208b, 32'hc1420c9e, 32'hc22859f9, 32'hc2bd5bd3, 32'h42464be2, 32'hc26ece2c};
test_output[7703] = '{32'h4282208b};
test_index[7703] = '{2};
test_input[61632:61639] = '{32'hc0951bd2, 32'h428d2fc6, 32'hc226145e, 32'hc0d32147, 32'hc2af3d34, 32'hc1896704, 32'hc2ab6841, 32'h41f7dc5b};
test_output[7704] = '{32'h428d2fc6};
test_index[7704] = '{1};
test_input[61640:61647] = '{32'hc2c4f268, 32'h40367bc8, 32'h421b8132, 32'hc2852927, 32'hc1c86b95, 32'h42b958dd, 32'h42bff36a, 32'hc27afad4};
test_output[7705] = '{32'h42bff36a};
test_index[7705] = '{6};
test_input[61648:61655] = '{32'hc2c03baa, 32'hc1b612b2, 32'hc1cf52d9, 32'hc27ddd43, 32'h41d8bf33, 32'h426ab0c9, 32'hc20d216c, 32'h421c53cb};
test_output[7706] = '{32'h426ab0c9};
test_index[7706] = '{5};
test_input[61656:61663] = '{32'h427b6dee, 32'hc1dd2254, 32'hc2bdc964, 32'hc2c46e66, 32'h42b99815, 32'hc27fc998, 32'h4220422f, 32'h425b5079};
test_output[7707] = '{32'h42b99815};
test_index[7707] = '{4};
test_input[61664:61671] = '{32'hc1915076, 32'hc238b46c, 32'hc2a0b4e2, 32'h429c7184, 32'hc2905407, 32'hc0e7a508, 32'hc221e125, 32'hc0a5ef8d};
test_output[7708] = '{32'h429c7184};
test_index[7708] = '{3};
test_input[61672:61679] = '{32'h3fa9f8b0, 32'h42c417b6, 32'hc0644980, 32'h41fb193e, 32'h410604cb, 32'h40da318a, 32'hc0728bb1, 32'h42b78050};
test_output[7709] = '{32'h42c417b6};
test_index[7709] = '{1};
test_input[61680:61687] = '{32'h42407519, 32'h428ba604, 32'hc2b2a53a, 32'h42867af9, 32'hc26af86d, 32'h421fab5d, 32'hc16e0cd8, 32'hc29d82bf};
test_output[7710] = '{32'h428ba604};
test_index[7710] = '{1};
test_input[61688:61695] = '{32'h427f2a44, 32'h42a03d2f, 32'h42044652, 32'hc19047fe, 32'hc23b240e, 32'h421c7fbc, 32'h4128aa05, 32'h423a9fe9};
test_output[7711] = '{32'h42a03d2f};
test_index[7711] = '{1};
test_input[61696:61703] = '{32'h42c7f20d, 32'hc240cbe4, 32'h42934ddf, 32'hc2c0306e, 32'h3fb2daff, 32'h421f719d, 32'hc284f65d, 32'hc1c0a307};
test_output[7712] = '{32'h42c7f20d};
test_index[7712] = '{0};
test_input[61704:61711] = '{32'h42815719, 32'hc2b926e0, 32'h428a799e, 32'h4291bcb3, 32'h42c4e783, 32'hc1a7b838, 32'hc228aff3, 32'hc0af7d79};
test_output[7713] = '{32'h42c4e783};
test_index[7713] = '{4};
test_input[61712:61719] = '{32'h422eea9c, 32'h41b635f7, 32'hc265c800, 32'hc1076931, 32'hc17cf327, 32'hc0db4ca8, 32'hc2bf9bc8, 32'h41b92f91};
test_output[7714] = '{32'h422eea9c};
test_index[7714] = '{0};
test_input[61720:61727] = '{32'h428e6725, 32'h41ce31ba, 32'h4198183e, 32'h42848566, 32'hc2baa28c, 32'h41dab697, 32'hc2a5889f, 32'h418f6313};
test_output[7715] = '{32'h428e6725};
test_index[7715] = '{0};
test_input[61728:61735] = '{32'hc076d07f, 32'h42a38934, 32'hc29d2011, 32'hc2b52972, 32'h42a72344, 32'h42108dec, 32'hc1a226fe, 32'h419923e1};
test_output[7716] = '{32'h42a72344};
test_index[7716] = '{4};
test_input[61736:61743] = '{32'hc28c62b3, 32'h4187188f, 32'hc2b169da, 32'h40a818b8, 32'h41f827ec, 32'h42c27711, 32'h423e6360, 32'h415dcc89};
test_output[7717] = '{32'h42c27711};
test_index[7717] = '{5};
test_input[61744:61751] = '{32'h402009d2, 32'hc1d139f9, 32'h4145c515, 32'h424b9737, 32'h42984388, 32'h429956df, 32'h429c8bf7, 32'hc2c0a8fb};
test_output[7718] = '{32'h429c8bf7};
test_index[7718] = '{6};
test_input[61752:61759] = '{32'hc2705baa, 32'h42aa8458, 32'h427b7a9a, 32'h42c5badd, 32'hc28ba695, 32'h41bf8d77, 32'h42b6f282, 32'h416b56cb};
test_output[7719] = '{32'h42c5badd};
test_index[7719] = '{3};
test_input[61760:61767] = '{32'h4257d07a, 32'hc2a865de, 32'h419445ad, 32'hc15178a6, 32'hc21f9dcb, 32'h428e2704, 32'h4232d0a8, 32'hc23266b8};
test_output[7720] = '{32'h428e2704};
test_index[7720] = '{5};
test_input[61768:61775] = '{32'h421a4c02, 32'h41bd7818, 32'h42a1cef9, 32'h428c09ca, 32'h4147cdcf, 32'h429e946d, 32'h42bf6d30, 32'h425ed53f};
test_output[7721] = '{32'h42bf6d30};
test_index[7721] = '{6};
test_input[61776:61783] = '{32'hc28ae8f5, 32'h41ec6a13, 32'hc2793a7c, 32'hc29f2cb6, 32'hc29bd057, 32'h41eefd1d, 32'hc2a33817, 32'h42bb034e};
test_output[7722] = '{32'h42bb034e};
test_index[7722] = '{7};
test_input[61784:61791] = '{32'hc21a7253, 32'h42074b80, 32'hc2a8c61b, 32'hc2400009, 32'hc27cbc07, 32'h4240b0cd, 32'hc24573df, 32'hc2bddde0};
test_output[7723] = '{32'h4240b0cd};
test_index[7723] = '{5};
test_input[61792:61799] = '{32'hc219eea4, 32'hc2aeb175, 32'hc24c758c, 32'hc038b811, 32'h3f2bf00a, 32'hc203db40, 32'h41590b73, 32'hc23cd82f};
test_output[7724] = '{32'h41590b73};
test_index[7724] = '{6};
test_input[61800:61807] = '{32'hc2855014, 32'hc2c44ef6, 32'h429ff05f, 32'hc2acc840, 32'h3e705af0, 32'h41e6be75, 32'h429221e0, 32'hc282817a};
test_output[7725] = '{32'h429ff05f};
test_index[7725] = '{2};
test_input[61808:61815] = '{32'hc29868b4, 32'h41f4a1a7, 32'hc2c3f3d6, 32'hc16bc2c8, 32'hc2ba6147, 32'hc20ca61b, 32'h42c6afff, 32'h42bdbb26};
test_output[7726] = '{32'h42c6afff};
test_index[7726] = '{6};
test_input[61816:61823] = '{32'h428da415, 32'h42a9f538, 32'h422cad7a, 32'hc276adca, 32'hc2b45331, 32'h42baf2f9, 32'hc2a351dc, 32'h42006d97};
test_output[7727] = '{32'h42baf2f9};
test_index[7727] = '{5};
test_input[61824:61831] = '{32'hc1c19cb7, 32'h41e34143, 32'h42c168f8, 32'h42974b18, 32'h41ea4a8f, 32'hc2a5adbc, 32'h4254dd94, 32'h4229c9af};
test_output[7728] = '{32'h42c168f8};
test_index[7728] = '{2};
test_input[61832:61839] = '{32'hc28d5c45, 32'hc18e7568, 32'hc2b2ad2e, 32'h42b4c59e, 32'h4222fb8c, 32'hc245cc35, 32'h42c3e3fd, 32'hc07a8afc};
test_output[7729] = '{32'h42c3e3fd};
test_index[7729] = '{6};
test_input[61840:61847] = '{32'h41e51b3a, 32'h42b5b875, 32'h415c0c96, 32'hc27dbd76, 32'h419b5990, 32'h4220edef, 32'h41d112fc, 32'h428b8006};
test_output[7730] = '{32'h42b5b875};
test_index[7730] = '{1};
test_input[61848:61855] = '{32'hc04bb39b, 32'hc29303fb, 32'hc28d8341, 32'hc17659a1, 32'h42c08452, 32'h42ac06ed, 32'hc2c50087, 32'h4193c32c};
test_output[7731] = '{32'h42c08452};
test_index[7731] = '{4};
test_input[61856:61863] = '{32'hc0ff5b55, 32'h4095ec58, 32'h421e7216, 32'hc0b441ed, 32'h426b0de9, 32'hc19267bc, 32'hc23c9419, 32'hc2ae5668};
test_output[7732] = '{32'h426b0de9};
test_index[7732] = '{4};
test_input[61864:61871] = '{32'hc2708d34, 32'hc26c6856, 32'hc2af69ed, 32'h423b6617, 32'hc021d50c, 32'h41bac506, 32'h42b49cd3, 32'hc2ac12c1};
test_output[7733] = '{32'h42b49cd3};
test_index[7733] = '{6};
test_input[61872:61879] = '{32'hc20ce099, 32'h42562a41, 32'h4286bf3d, 32'h41a7ce07, 32'h42463c21, 32'hc2c03b4b, 32'h41121483, 32'hc284bca3};
test_output[7734] = '{32'h4286bf3d};
test_index[7734] = '{2};
test_input[61880:61887] = '{32'hc249708e, 32'h427abd9e, 32'h428d8869, 32'h425d2456, 32'hc294b598, 32'h428a3ab9, 32'h4287d29b, 32'h3ec42db2};
test_output[7735] = '{32'h428d8869};
test_index[7735] = '{2};
test_input[61888:61895] = '{32'hc12a1433, 32'h42c4372b, 32'hc2aa688a, 32'hbed02b01, 32'hc21090c0, 32'h428e2cd0, 32'hc290b6ce, 32'h41d64b6a};
test_output[7736] = '{32'h42c4372b};
test_index[7736] = '{1};
test_input[61896:61903] = '{32'h42519ee9, 32'h42c71797, 32'h429d0bf5, 32'hc11f7b62, 32'h42bd0b93, 32'h420984fb, 32'hc2c2b88e, 32'h42031c7c};
test_output[7737] = '{32'h42c71797};
test_index[7737] = '{1};
test_input[61904:61911] = '{32'h41a636c5, 32'hc0a7ef9f, 32'hc29e9ab9, 32'h4218264a, 32'h3f8a1263, 32'hc29711b0, 32'h42ac7fc7, 32'hc25bbb41};
test_output[7738] = '{32'h42ac7fc7};
test_index[7738] = '{6};
test_input[61912:61919] = '{32'h41cd91df, 32'h4282455c, 32'hc2310376, 32'h4289846d, 32'h42c00b7e, 32'hc2257aaf, 32'h42a5e5c7, 32'h41841b0f};
test_output[7739] = '{32'h42c00b7e};
test_index[7739] = '{4};
test_input[61920:61927] = '{32'h427f07d5, 32'h4264a95d, 32'h429fabb7, 32'hc0e10462, 32'hc1d80901, 32'hc2ab6aeb, 32'hc215df8f, 32'h41ddf9fe};
test_output[7740] = '{32'h429fabb7};
test_index[7740] = '{2};
test_input[61928:61935] = '{32'h425c5dcd, 32'h4245cd58, 32'hc2491633, 32'hc23157c3, 32'h4154fcd9, 32'h42834ff3, 32'hc289bd05, 32'hc2149e44};
test_output[7741] = '{32'h42834ff3};
test_index[7741] = '{5};
test_input[61936:61943] = '{32'hc02f1901, 32'hc2933d86, 32'hc2a48f6d, 32'hc227e9a3, 32'h42552440, 32'hc2ae0cf7, 32'h41a65bbc, 32'hc1266116};
test_output[7742] = '{32'h42552440};
test_index[7742] = '{4};
test_input[61944:61951] = '{32'hc25f7ecc, 32'hc29a9452, 32'hc28246a3, 32'hc11f4270, 32'hc204bfe4, 32'h41bc8e8a, 32'h4240dabd, 32'hc2100861};
test_output[7743] = '{32'h4240dabd};
test_index[7743] = '{6};
test_input[61952:61959] = '{32'hc109cf10, 32'hc0d961e7, 32'hc1b698cb, 32'h3f484f93, 32'h42c0a736, 32'hc2bdf911, 32'hc1d1395d, 32'h42909d29};
test_output[7744] = '{32'h42c0a736};
test_index[7744] = '{4};
test_input[61960:61967] = '{32'h42ba85bb, 32'h41e80b3c, 32'hc17e4280, 32'h41bba943, 32'h42ba104d, 32'hc0b4007f, 32'h4209ad2f, 32'hc09791f3};
test_output[7745] = '{32'h42ba85bb};
test_index[7745] = '{0};
test_input[61968:61975] = '{32'h424e582e, 32'h410161ca, 32'h41aede3d, 32'h426bcb06, 32'h42b82c4a, 32'h41ad161e, 32'h41f9083d, 32'h4252758a};
test_output[7746] = '{32'h42b82c4a};
test_index[7746] = '{4};
test_input[61976:61983] = '{32'h41d88ee1, 32'hc275a209, 32'hc2a63d97, 32'hc24b7132, 32'hc28c6892, 32'h42aa5920, 32'h42beea30, 32'h427e4c6c};
test_output[7747] = '{32'h42beea30};
test_index[7747] = '{6};
test_input[61984:61991] = '{32'hc2819351, 32'h42b851ac, 32'hc2c5486f, 32'hc2247dc6, 32'hc1fcd737, 32'h42385d9e, 32'hc2559686, 32'hc2a2efac};
test_output[7748] = '{32'h42b851ac};
test_index[7748] = '{1};
test_input[61992:61999] = '{32'hc20108c0, 32'hc25eae70, 32'h4224146b, 32'hc2bbb1ba, 32'hc2699e45, 32'h4293d0bb, 32'h40c838d1, 32'hc133eea4};
test_output[7749] = '{32'h4293d0bb};
test_index[7749] = '{5};
test_input[62000:62007] = '{32'hc2c4cff7, 32'h426c5967, 32'hc29617f0, 32'h42c108e2, 32'h420802e1, 32'h426b902d, 32'hc28dea46, 32'h425e9742};
test_output[7750] = '{32'h42c108e2};
test_index[7750] = '{3};
test_input[62008:62015] = '{32'h4228ac09, 32'h42c1281d, 32'hc0366205, 32'hc230596f, 32'hc16892c9, 32'h41b864ec, 32'hc2be8716, 32'hc27d363d};
test_output[7751] = '{32'h42c1281d};
test_index[7751] = '{1};
test_input[62016:62023] = '{32'hc2872c48, 32'hc2956ded, 32'hc2296f94, 32'h42b49729, 32'h4125c988, 32'h418fde2b, 32'h4290ad8f, 32'hbf05bf7f};
test_output[7752] = '{32'h42b49729};
test_index[7752] = '{3};
test_input[62024:62031] = '{32'hc2854890, 32'hc211e261, 32'h403f0c1b, 32'h419317f2, 32'hc194eaf2, 32'hc28b3df0, 32'h4213af91, 32'hc27d04ec};
test_output[7753] = '{32'h4213af91};
test_index[7753] = '{6};
test_input[62032:62039] = '{32'h424e73a9, 32'hc29aa57a, 32'hc20ae41b, 32'hc29ea4fa, 32'h4261e597, 32'h429cf788, 32'hc21dca58, 32'hc1b86319};
test_output[7754] = '{32'h429cf788};
test_index[7754] = '{5};
test_input[62040:62047] = '{32'h422fd815, 32'hc2672e0f, 32'h42c6733b, 32'hc19b6cbd, 32'h412ec8f7, 32'hc28e5490, 32'hc291b649, 32'h4107efb9};
test_output[7755] = '{32'h42c6733b};
test_index[7755] = '{2};
test_input[62048:62055] = '{32'h42b1f5a1, 32'h42a1d8d1, 32'h419bc9ed, 32'h42a65c05, 32'h42be7a8d, 32'hc26f9c24, 32'h42c50025, 32'hc25ac4cc};
test_output[7756] = '{32'h42c50025};
test_index[7756] = '{6};
test_input[62056:62063] = '{32'hc2896c64, 32'h4293703c, 32'h40d07ace, 32'h42bb233c, 32'hc25bf42d, 32'hc0878768, 32'hc10972ca, 32'hc282c550};
test_output[7757] = '{32'h42bb233c};
test_index[7757] = '{3};
test_input[62064:62071] = '{32'h425ed80c, 32'hc2b7c577, 32'h42920d1c, 32'h40c2f8b3, 32'hc289f52c, 32'hc24236a0, 32'h42421b85, 32'h4232667e};
test_output[7758] = '{32'h42920d1c};
test_index[7758] = '{2};
test_input[62072:62079] = '{32'h42b20129, 32'h41f65f7d, 32'h4245f11c, 32'h42b05e21, 32'hc110dd2c, 32'hc24de9c4, 32'h4137b1e5, 32'hc2793b78};
test_output[7759] = '{32'h42b20129};
test_index[7759] = '{0};
test_input[62080:62087] = '{32'h422cf7c0, 32'h42057195, 32'hc23ee405, 32'hc229a9bf, 32'h4250976d, 32'h428bb490, 32'hc2984be4, 32'h3f8d14db};
test_output[7760] = '{32'h428bb490};
test_index[7760] = '{5};
test_input[62088:62095] = '{32'h415f2813, 32'h41974134, 32'h42869572, 32'h42aabae9, 32'hc13da905, 32'h42a19ebb, 32'hc2739a45, 32'hc265f736};
test_output[7761] = '{32'h42aabae9};
test_index[7761] = '{3};
test_input[62096:62103] = '{32'h409cde9e, 32'h4252a52b, 32'hc25eab6d, 32'hc294927d, 32'h42999f3b, 32'h41afc4cf, 32'hc21c0860, 32'hc1772385};
test_output[7762] = '{32'h42999f3b};
test_index[7762] = '{4};
test_input[62104:62111] = '{32'h4184deaa, 32'hc2aea339, 32'h424aecfc, 32'h4295bfdc, 32'hc16f4e75, 32'hc2579371, 32'h42b349ca, 32'h4216b04e};
test_output[7763] = '{32'h42b349ca};
test_index[7763] = '{6};
test_input[62112:62119] = '{32'h4287c63e, 32'h4283419f, 32'h41900dbe, 32'hc21d9c03, 32'hc0ade03a, 32'hc1fa332f, 32'hc19e74fe, 32'h4219b8ba};
test_output[7764] = '{32'h4287c63e};
test_index[7764] = '{0};
test_input[62120:62127] = '{32'h41c238ac, 32'hc1b6d2e8, 32'h429ec7d3, 32'h426ae379, 32'h42b63d3e, 32'h419cb779, 32'hc286615c, 32'h41a0a322};
test_output[7765] = '{32'h42b63d3e};
test_index[7765] = '{4};
test_input[62128:62135] = '{32'h42be9fe1, 32'h42c70ad9, 32'hc21e4ae1, 32'hc218d788, 32'h4296530b, 32'hc1fa9ba3, 32'hc2bea384, 32'h42115d60};
test_output[7766] = '{32'h42c70ad9};
test_index[7766] = '{1};
test_input[62136:62143] = '{32'hc2bf4d97, 32'hc2878415, 32'h42234a95, 32'h4250076f, 32'hc2474fd8, 32'h419a07c4, 32'h42aa584a, 32'hc2659e79};
test_output[7767] = '{32'h42aa584a};
test_index[7767] = '{6};
test_input[62144:62151] = '{32'h425956be, 32'hc08156f6, 32'hc238ba5c, 32'h428be83d, 32'h41bb4a51, 32'hc2a9401e, 32'h4292d0db, 32'h42473c97};
test_output[7768] = '{32'h4292d0db};
test_index[7768] = '{6};
test_input[62152:62159] = '{32'hc288054d, 32'h401aa984, 32'hc0627550, 32'h425d3164, 32'h4241fa54, 32'hc2b99857, 32'hc2b8d355, 32'hc24fe0dd};
test_output[7769] = '{32'h425d3164};
test_index[7769] = '{3};
test_input[62160:62167] = '{32'h429edcbf, 32'h41e4af0a, 32'hc1d8e854, 32'hc1b0d6ce, 32'h42c745f0, 32'h428422ce, 32'h42169dc8, 32'h42bcd06d};
test_output[7770] = '{32'h42c745f0};
test_index[7770] = '{4};
test_input[62168:62175] = '{32'hc1f54271, 32'h4271ec22, 32'h42bd4e11, 32'hc276d23a, 32'h421f6f9b, 32'hc2b641f0, 32'h421f49d6, 32'hc2b1c8dc};
test_output[7771] = '{32'h42bd4e11};
test_index[7771] = '{2};
test_input[62176:62183] = '{32'h4288629a, 32'hc29e59f9, 32'h3e75d0af, 32'hc2af5278, 32'hc24b7492, 32'hc2b729c0, 32'hc264a2e9, 32'h4282f91a};
test_output[7772] = '{32'h4288629a};
test_index[7772] = '{0};
test_input[62184:62191] = '{32'hc101332e, 32'h42c71b9b, 32'hc2b4b62f, 32'h4191f2e2, 32'h4148551e, 32'hc2014df0, 32'h4263fec4, 32'h429402fa};
test_output[7773] = '{32'h42c71b9b};
test_index[7773] = '{1};
test_input[62192:62199] = '{32'hc1ec4dab, 32'hc2be0451, 32'h40a4c35f, 32'hc2b147d1, 32'h3c9a1c9b, 32'hc2b6fd92, 32'hc28f7965, 32'h41c51e99};
test_output[7774] = '{32'h41c51e99};
test_index[7774] = '{7};
test_input[62200:62207] = '{32'h41707849, 32'h4282fdbb, 32'h424c1510, 32'h42412927, 32'h42ad669c, 32'h41ff442d, 32'h429e59a4, 32'h4281a5b7};
test_output[7775] = '{32'h42ad669c};
test_index[7775] = '{4};
test_input[62208:62215] = '{32'hc29b7577, 32'h42bea6d8, 32'hc2565503, 32'hc2b1a11e, 32'h427003aa, 32'hc21707d1, 32'hbe8cbd58, 32'h41f5b9d9};
test_output[7776] = '{32'h42bea6d8};
test_index[7776] = '{1};
test_input[62216:62223] = '{32'hc2ade9e9, 32'h42620884, 32'h426132f5, 32'hc2afdf01, 32'h425f1d7f, 32'hc22201b3, 32'hc2745677, 32'hc2014222};
test_output[7777] = '{32'h42620884};
test_index[7777] = '{1};
test_input[62224:62231] = '{32'hc284d4fb, 32'hc28354ec, 32'h42182d57, 32'hc11d516f, 32'h4236dbf5, 32'h421ae791, 32'h4109d11d, 32'h41e6ac26};
test_output[7778] = '{32'h4236dbf5};
test_index[7778] = '{4};
test_input[62232:62239] = '{32'hc18fa6f1, 32'h42c18399, 32'hc14bffa0, 32'h411109e5, 32'h42bad6ab, 32'h41d28f8e, 32'hc285f8c2, 32'hc22d8009};
test_output[7779] = '{32'h42c18399};
test_index[7779] = '{1};
test_input[62240:62247] = '{32'hc29a06d1, 32'h3da271c3, 32'hc21ce95e, 32'hc2507420, 32'hc135a0fd, 32'h4292e51f, 32'h42682eb2, 32'hc2377710};
test_output[7780] = '{32'h4292e51f};
test_index[7780] = '{5};
test_input[62248:62255] = '{32'h4258a37b, 32'h4289d20f, 32'hc208e31a, 32'h42c12295, 32'hc05ffdb6, 32'hc223d9e6, 32'h426e49f6, 32'hc2824cd8};
test_output[7781] = '{32'h42c12295};
test_index[7781] = '{3};
test_input[62256:62263] = '{32'h410abea5, 32'hc2130fdb, 32'h42b5e7ac, 32'h41c98141, 32'h42b1031e, 32'hc11bc088, 32'h41be055b, 32'hc1652c5c};
test_output[7782] = '{32'h42b5e7ac};
test_index[7782] = '{2};
test_input[62264:62271] = '{32'hc2068398, 32'h425deb21, 32'h40af138e, 32'h426bf430, 32'hc25cf790, 32'h42101586, 32'h41861399, 32'h4241a7b3};
test_output[7783] = '{32'h426bf430};
test_index[7783] = '{3};
test_input[62272:62279] = '{32'hc2b31535, 32'h41733b43, 32'h425cfb15, 32'h426d8052, 32'h40cc56c2, 32'h40e52457, 32'h4298dfbb, 32'h42b7b183};
test_output[7784] = '{32'h42b7b183};
test_index[7784] = '{7};
test_input[62280:62287] = '{32'h42890442, 32'h427e53dc, 32'h41d17857, 32'hc2ac0fb0, 32'hc1ae3b19, 32'hc2b37cd8, 32'h41012335, 32'hc2688a68};
test_output[7785] = '{32'h42890442};
test_index[7785] = '{0};
test_input[62288:62295] = '{32'hc2bb5473, 32'h428f864b, 32'h42b96e62, 32'h428fd584, 32'h423f3696, 32'hc20850a0, 32'h42a47ff5, 32'hc13bef70};
test_output[7786] = '{32'h42b96e62};
test_index[7786] = '{2};
test_input[62296:62303] = '{32'h4240e582, 32'h4232a919, 32'h429e00a4, 32'hc28c05eb, 32'h41e040e2, 32'hc2c15d00, 32'hc27d0c2a, 32'hc291e670};
test_output[7787] = '{32'h429e00a4};
test_index[7787] = '{2};
test_input[62304:62311] = '{32'h426f5608, 32'hc1d8ca02, 32'h426b50a5, 32'hc2914912, 32'hc21853cd, 32'hc21ce97a, 32'h427c84c0, 32'h42c19a33};
test_output[7788] = '{32'h42c19a33};
test_index[7788] = '{7};
test_input[62312:62319] = '{32'h427d966b, 32'h4172b28c, 32'h41be04b4, 32'h4287840d, 32'hc2257373, 32'hc0e2d89b, 32'h41db16f8, 32'hc201ef01};
test_output[7789] = '{32'h4287840d};
test_index[7789] = '{3};
test_input[62320:62327] = '{32'h428c094a, 32'hc28700da, 32'h410fa59b, 32'hc29ac8eb, 32'h423a5b8a, 32'hc29bfe28, 32'h4168bcbb, 32'h4294b2aa};
test_output[7790] = '{32'h4294b2aa};
test_index[7790] = '{7};
test_input[62328:62335] = '{32'hc280b6df, 32'h4278b41d, 32'h41b05003, 32'hc180b3d7, 32'hc2affb9c, 32'hc28325bb, 32'hc24622bb, 32'hc1c86694};
test_output[7791] = '{32'h4278b41d};
test_index[7791] = '{1};
test_input[62336:62343] = '{32'h42c6eb6b, 32'h42a87639, 32'h42933b17, 32'h42b42d38, 32'hc2ac57b2, 32'h41f23991, 32'hc264d2fe, 32'h4273dca6};
test_output[7792] = '{32'h42c6eb6b};
test_index[7792] = '{0};
test_input[62344:62351] = '{32'hc2c6cdc1, 32'h42391e07, 32'hc06d120f, 32'h42b7da3b, 32'hc2127344, 32'h42c51a88, 32'hc284cd09, 32'hc158ec2b};
test_output[7793] = '{32'h42c51a88};
test_index[7793] = '{5};
test_input[62352:62359] = '{32'hc1082755, 32'h420ba9df, 32'hc2434be0, 32'h419ee836, 32'hc29bebea, 32'h42776b31, 32'h41c4d509, 32'hc29eff5d};
test_output[7794] = '{32'h42776b31};
test_index[7794] = '{5};
test_input[62360:62367] = '{32'hc279e280, 32'h420675e0, 32'hc2147c98, 32'h4257b547, 32'hc2bd3f34, 32'h429e20da, 32'hc2c15d2b, 32'hc29d953f};
test_output[7795] = '{32'h429e20da};
test_index[7795] = '{5};
test_input[62368:62375] = '{32'hc2475526, 32'hc10cb992, 32'h41db8f14, 32'h420421ea, 32'h40f7df25, 32'h4294a330, 32'h424e88c0, 32'h42ae4fd4};
test_output[7796] = '{32'h42ae4fd4};
test_index[7796] = '{7};
test_input[62376:62383] = '{32'h425736fc, 32'h427716e1, 32'hc0ec190e, 32'hc295b186, 32'h421bade7, 32'h418af81d, 32'hc28cc875, 32'h4236a38a};
test_output[7797] = '{32'h427716e1};
test_index[7797] = '{1};
test_input[62384:62391] = '{32'hc129ef87, 32'hc09621de, 32'hc2833da5, 32'hc25641fa, 32'h42c44e91, 32'hc1ee6ef6, 32'hc2c74dfd, 32'h42017f7c};
test_output[7798] = '{32'h42c44e91};
test_index[7798] = '{4};
test_input[62392:62399] = '{32'h420a00ef, 32'h422dd43e, 32'hc1f334c0, 32'hc20bf270, 32'hc2aa078c, 32'h42910fea, 32'h418389ab, 32'h423865bd};
test_output[7799] = '{32'h42910fea};
test_index[7799] = '{5};
test_input[62400:62407] = '{32'h428b174d, 32'h4292dac4, 32'h41c1bd77, 32'h42a299d9, 32'hc2bdf342, 32'h41c40354, 32'h42c759a6, 32'hc29d3412};
test_output[7800] = '{32'h42c759a6};
test_index[7800] = '{6};
test_input[62408:62415] = '{32'hc244b89c, 32'hc29bd346, 32'hc208e21e, 32'h4201d3d0, 32'hc23a9e94, 32'hc11a1363, 32'hc2acbeae, 32'h424ebd97};
test_output[7801] = '{32'h424ebd97};
test_index[7801] = '{7};
test_input[62416:62423] = '{32'h4143632b, 32'hc2c3bb49, 32'h422024de, 32'h42b38674, 32'h424192e2, 32'h4250d30a, 32'h4228b4a1, 32'hc2191588};
test_output[7802] = '{32'h42b38674};
test_index[7802] = '{3};
test_input[62424:62431] = '{32'hc2b2a2e5, 32'h421d4e9c, 32'hc203bdea, 32'hc2a38cbd, 32'h4283e0f0, 32'h4115bcfe, 32'hc2b386a8, 32'hbff129f8};
test_output[7803] = '{32'h4283e0f0};
test_index[7803] = '{4};
test_input[62432:62439] = '{32'hc2250ffe, 32'hc2aabaae, 32'h42012903, 32'hc19f9403, 32'h41ea5f78, 32'h425f3d07, 32'hc2a1e60f, 32'hbf9008bf};
test_output[7804] = '{32'h425f3d07};
test_index[7804] = '{5};
test_input[62440:62447] = '{32'hc296132f, 32'hc235df1a, 32'hc2910fc2, 32'h40d82d11, 32'hc164ec12, 32'h41b211c2, 32'hc12931c5, 32'hbf9c99d3};
test_output[7805] = '{32'h41b211c2};
test_index[7805] = '{5};
test_input[62448:62455] = '{32'h416b1569, 32'h4155737d, 32'h41c98c2e, 32'hc2a7a86f, 32'h4230e105, 32'h4252ccb3, 32'hc294d5f6, 32'h42334682};
test_output[7806] = '{32'h4252ccb3};
test_index[7806] = '{5};
test_input[62456:62463] = '{32'hc0dd6da5, 32'hc21ed683, 32'hc25c317c, 32'h42b31dea, 32'hc2c6c218, 32'h426ddb74, 32'hc2a0176c, 32'hc29d793d};
test_output[7807] = '{32'h42b31dea};
test_index[7807] = '{3};
test_input[62464:62471] = '{32'hc1f3fd05, 32'h42916775, 32'h424c1a27, 32'h41134399, 32'h42a196c3, 32'h42bdc93d, 32'h42128764, 32'hbf82c5c8};
test_output[7808] = '{32'h42bdc93d};
test_index[7808] = '{5};
test_input[62472:62479] = '{32'hc21bfc6e, 32'h410d7e58, 32'hc20fdad9, 32'hc134b236, 32'hc2545593, 32'h42968b20, 32'h41f65212, 32'hc209d6d8};
test_output[7809] = '{32'h42968b20};
test_index[7809] = '{5};
test_input[62480:62487] = '{32'hc11753bc, 32'h422418de, 32'hc261db5c, 32'h4138039a, 32'hc299c558, 32'hc2ab6a47, 32'hc25cf422, 32'h4201c89f};
test_output[7810] = '{32'h422418de};
test_index[7810] = '{1};
test_input[62488:62495] = '{32'hbe21c70e, 32'h42c3625f, 32'hc2c4056e, 32'hc1fea471, 32'h42996a67, 32'h42ab53bb, 32'hc229d07b, 32'h425e3bbf};
test_output[7811] = '{32'h42c3625f};
test_index[7811] = '{1};
test_input[62496:62503] = '{32'hc2a8ea9a, 32'h421034cf, 32'hc1bc477e, 32'hc08a322b, 32'h42ab7fa5, 32'h424b658f, 32'h423ce9ee, 32'hc2854783};
test_output[7812] = '{32'h42ab7fa5};
test_index[7812] = '{4};
test_input[62504:62511] = '{32'h42810f9d, 32'h42c62419, 32'hc00f5b10, 32'hc2bcda3a, 32'h42a8a7a9, 32'h4222a249, 32'h42640d0f, 32'h42bfbfaf};
test_output[7813] = '{32'h42c62419};
test_index[7813] = '{1};
test_input[62512:62519] = '{32'h41a8a7f8, 32'hc2b223c7, 32'hc20396e7, 32'hbdd73425, 32'hc121fbc7, 32'h404746dd, 32'hc09cf25b, 32'h41cf179f};
test_output[7814] = '{32'h41cf179f};
test_index[7814] = '{7};
test_input[62520:62527] = '{32'hc29fe1f3, 32'hc29eaeae, 32'hc2506477, 32'h40eda21d, 32'hc2288608, 32'hc2c3289a, 32'hc1404f54, 32'h403ce871};
test_output[7815] = '{32'h40eda21d};
test_index[7815] = '{3};
test_input[62528:62535] = '{32'hc2adcdf4, 32'h40d860d5, 32'hc1c59ea7, 32'hc288f7e3, 32'hc20705a5, 32'h42c2467f, 32'hc0b186f7, 32'h428a70de};
test_output[7816] = '{32'h42c2467f};
test_index[7816] = '{5};
test_input[62536:62543] = '{32'hc2bbbcb4, 32'hc2a1cb9f, 32'h422bb8ac, 32'hc2176177, 32'h42679d12, 32'h428a3432, 32'hc21432e4, 32'hc0bd9ce6};
test_output[7817] = '{32'h428a3432};
test_index[7817] = '{5};
test_input[62544:62551] = '{32'h41dba627, 32'hc27f7258, 32'hc2a4f066, 32'hc2904bda, 32'hc13630fd, 32'h42691c56, 32'hc1c756cb, 32'h4206612e};
test_output[7818] = '{32'h42691c56};
test_index[7818] = '{5};
test_input[62552:62559] = '{32'hc2523057, 32'hc1cf40ba, 32'h41f45ef1, 32'h4205cc11, 32'h42907311, 32'h42116985, 32'h427560fe, 32'hc2bb7722};
test_output[7819] = '{32'h42907311};
test_index[7819] = '{4};
test_input[62560:62567] = '{32'hc161ff8e, 32'h42c549a7, 32'h4114ee03, 32'h429c0379, 32'h40bcabbb, 32'h41c71779, 32'hc1a0e3c1, 32'hc22ccc4e};
test_output[7820] = '{32'h42c549a7};
test_index[7820] = '{1};
test_input[62568:62575] = '{32'h4287bfe4, 32'hc293556f, 32'hc0b06a2a, 32'h42b864d7, 32'h42071be3, 32'hc2b6b044, 32'hc1d3ef15, 32'hc2c7789a};
test_output[7821] = '{32'h42b864d7};
test_index[7821] = '{3};
test_input[62576:62583] = '{32'hc2556ebf, 32'hc2408353, 32'hc261e12c, 32'h3f8f8496, 32'h42ab10fa, 32'h41e1eb6e, 32'hc2b39f89, 32'h4249076d};
test_output[7822] = '{32'h42ab10fa};
test_index[7822] = '{4};
test_input[62584:62591] = '{32'hc1869fa4, 32'hc05a0531, 32'h42840a64, 32'h41d4fc7b, 32'hc1ed0ea1, 32'hc2660164, 32'hc18b9447, 32'h40c237c6};
test_output[7823] = '{32'h42840a64};
test_index[7823] = '{2};
test_input[62592:62599] = '{32'hc224c58e, 32'h42b653e6, 32'h400fba0f, 32'h4296cdb3, 32'h40be6bad, 32'h42b71f9a, 32'hc279044d, 32'hc2c2138c};
test_output[7824] = '{32'h42b71f9a};
test_index[7824] = '{5};
test_input[62600:62607] = '{32'h42b9cf0a, 32'hc28044c9, 32'hc22e6641, 32'hc1aeb00d, 32'h41a02b05, 32'h41658d89, 32'h41406858, 32'h428bc9cf};
test_output[7825] = '{32'h42b9cf0a};
test_index[7825] = '{0};
test_input[62608:62615] = '{32'hc19c0d12, 32'h420395c4, 32'h40fba891, 32'h428538ae, 32'h412468e7, 32'h41a59ce5, 32'h42af36c2, 32'hc2c35266};
test_output[7826] = '{32'h42af36c2};
test_index[7826] = '{6};
test_input[62616:62623] = '{32'hc1e0c016, 32'hc26abb93, 32'h42befbb8, 32'h42a02b12, 32'h421ec34b, 32'h42bcd048, 32'h4250b855, 32'hc0a35e96};
test_output[7827] = '{32'h42befbb8};
test_index[7827] = '{2};
test_input[62624:62631] = '{32'h4217bcbb, 32'hc096b8e1, 32'hc2b450c4, 32'hc2a61d5f, 32'hc1561bb1, 32'hc26a0441, 32'h41a3444b, 32'hc2a7d5c9};
test_output[7828] = '{32'h4217bcbb};
test_index[7828] = '{0};
test_input[62632:62639] = '{32'hc28ba66d, 32'h426d4289, 32'h405181e4, 32'hc14554ee, 32'hc2b4f7c2, 32'h429062a6, 32'hc21ac845, 32'h411ae860};
test_output[7829] = '{32'h429062a6};
test_index[7829] = '{5};
test_input[62640:62647] = '{32'h3ee6d75b, 32'h42be4ad5, 32'h42bc50b8, 32'h428a7f16, 32'hc121007c, 32'h42c00dfb, 32'hbe940f1d, 32'hc2b401ec};
test_output[7830] = '{32'h42c00dfb};
test_index[7830] = '{5};
test_input[62648:62655] = '{32'hc2270110, 32'h4209f627, 32'hc1d9e9f1, 32'hc2216933, 32'h42b2669a, 32'h41632063, 32'hc27bb1c7, 32'hc23dca95};
test_output[7831] = '{32'h42b2669a};
test_index[7831] = '{4};
test_input[62656:62663] = '{32'hc26923fb, 32'hc2923d8e, 32'h42124c8c, 32'h427c4d02, 32'h4194a138, 32'hbea1a4fa, 32'h429aefa8, 32'h3f33dad7};
test_output[7832] = '{32'h429aefa8};
test_index[7832] = '{6};
test_input[62664:62671] = '{32'hc1e71f5f, 32'h4212d7d1, 32'hc2c54300, 32'hc204b6c5, 32'hc294a2dd, 32'hc0c0f977, 32'h426e147c, 32'h42c7540c};
test_output[7833] = '{32'h42c7540c};
test_index[7833] = '{7};
test_input[62672:62679] = '{32'hc2905c7d, 32'h42197895, 32'hc2118975, 32'hc2a76787, 32'h42be3662, 32'hc0126354, 32'h4201efa9, 32'h42877d4c};
test_output[7834] = '{32'h42be3662};
test_index[7834] = '{4};
test_input[62680:62687] = '{32'hc26430e7, 32'hc21fa7db, 32'hc28dd68e, 32'h426add7a, 32'h425f7da4, 32'hc23f4bb4, 32'hc28dd2e5, 32'hc2923884};
test_output[7835] = '{32'h426add7a};
test_index[7835] = '{3};
test_input[62688:62695] = '{32'hc20e2644, 32'h40cecddf, 32'hc2786df1, 32'hc25978b1, 32'hc2b47289, 32'hc2bebd74, 32'hc2420842, 32'hc2717515};
test_output[7836] = '{32'h40cecddf};
test_index[7836] = '{1};
test_input[62696:62703] = '{32'h42c58360, 32'h428a4773, 32'h42b2d166, 32'h42ab4aac, 32'hc2782648, 32'hc2a11e89, 32'hc2a47b15, 32'h42c3a428};
test_output[7837] = '{32'h42c58360};
test_index[7837] = '{0};
test_input[62704:62711] = '{32'h420e2712, 32'hbefe6730, 32'h422fb7b6, 32'hc25b52f4, 32'hc12a225a, 32'h42147d63, 32'h4120e47f, 32'h410db730};
test_output[7838] = '{32'h422fb7b6};
test_index[7838] = '{2};
test_input[62712:62719] = '{32'hc116df9f, 32'h420353c1, 32'h4213a656, 32'h4263a757, 32'h41ef1d51, 32'h41427587, 32'h421a4993, 32'h4168e321};
test_output[7839] = '{32'h4263a757};
test_index[7839] = '{3};
test_input[62720:62727] = '{32'h424b0e82, 32'h42b777bd, 32'h423afec4, 32'h4260d77e, 32'h42a60a16, 32'hc2076394, 32'hc281d9cf, 32'hc1d6d0dd};
test_output[7840] = '{32'h42b777bd};
test_index[7840] = '{1};
test_input[62728:62735] = '{32'hc20661d7, 32'h422cb921, 32'h41b539f7, 32'h415956b9, 32'h42062f75, 32'h42b8a3ac, 32'h3ef5b915, 32'h41d16f5b};
test_output[7841] = '{32'h42b8a3ac};
test_index[7841] = '{5};
test_input[62736:62743] = '{32'hbed84cbc, 32'h42af6da0, 32'hc2a9b542, 32'hc0075b1c, 32'h428d222d, 32'hc2aa8d41, 32'h4204e6f1, 32'h41b21509};
test_output[7842] = '{32'h42af6da0};
test_index[7842] = '{1};
test_input[62744:62751] = '{32'hc2c6d38a, 32'hc213a8f1, 32'h4084006a, 32'hc21537d5, 32'h42bd9d08, 32'h428c545b, 32'h41b7d988, 32'hc242fbd9};
test_output[7843] = '{32'h42bd9d08};
test_index[7843] = '{4};
test_input[62752:62759] = '{32'h4190af8e, 32'h414bf698, 32'hc28bd2ca, 32'h4289704d, 32'hc22e2be9, 32'hc291480a, 32'hc21ed01c, 32'h42797df0};
test_output[7844] = '{32'h4289704d};
test_index[7844] = '{3};
test_input[62760:62767] = '{32'h42743149, 32'h41fd8f4f, 32'hc134ebf0, 32'hc24ef9fe, 32'hc1a949f0, 32'hc1dd3b64, 32'hc23e1e01, 32'h42c44644};
test_output[7845] = '{32'h42c44644};
test_index[7845] = '{7};
test_input[62768:62775] = '{32'hc19d0ad1, 32'h42adeafd, 32'h41762688, 32'hc1c227ca, 32'h4285be20, 32'hc19d2f2f, 32'hc2ad1268, 32'h4293e2a6};
test_output[7846] = '{32'h42adeafd};
test_index[7846] = '{1};
test_input[62776:62783] = '{32'hc23c7ca3, 32'hc2563294, 32'hc29c2c68, 32'h429157e5, 32'hc29cb435, 32'h426637b2, 32'h4269431d, 32'hc2c58662};
test_output[7847] = '{32'h429157e5};
test_index[7847] = '{3};
test_input[62784:62791] = '{32'hc292676b, 32'h428b55d8, 32'hc292abee, 32'hc2a9a86d, 32'h42ace4a5, 32'hc2ad5dcb, 32'hc1d3f704, 32'hc23e7652};
test_output[7848] = '{32'h42ace4a5};
test_index[7848] = '{4};
test_input[62792:62799] = '{32'hc2860519, 32'h423b2793, 32'hc1d08f25, 32'h42bb93f7, 32'hc256012e, 32'h42b3394d, 32'h421fd408, 32'h429a2c1c};
test_output[7849] = '{32'h42bb93f7};
test_index[7849] = '{3};
test_input[62800:62807] = '{32'h40556171, 32'hc2720413, 32'h4225f224, 32'hc28db0b2, 32'h42bc0089, 32'hc1a475b5, 32'hc2b363f1, 32'hc246e367};
test_output[7850] = '{32'h42bc0089};
test_index[7850] = '{4};
test_input[62808:62815] = '{32'hc23d3fd6, 32'hc13d193a, 32'h4267538a, 32'hc218d179, 32'h4267d0d7, 32'hc2627358, 32'hc292578d, 32'h40e6d88f};
test_output[7851] = '{32'h4267d0d7};
test_index[7851] = '{4};
test_input[62816:62823] = '{32'h429a31be, 32'h4212e90c, 32'hc27bfcab, 32'hc225eeeb, 32'h42afbfb9, 32'h41c3d123, 32'h4269cc02, 32'h42838b2a};
test_output[7852] = '{32'h42afbfb9};
test_index[7852] = '{4};
test_input[62824:62831] = '{32'hc2be51a5, 32'hc1846d5f, 32'h42042367, 32'hc1893265, 32'h4250c09e, 32'hc260230f, 32'h42ad68d0, 32'hc29eb8d6};
test_output[7853] = '{32'h42ad68d0};
test_index[7853] = '{6};
test_input[62832:62839] = '{32'hc2019930, 32'h423f5a7b, 32'h420d4651, 32'hc2914235, 32'h41a57f77, 32'hc23ff1d9, 32'h426cd82a, 32'h42b02280};
test_output[7854] = '{32'h42b02280};
test_index[7854] = '{7};
test_input[62840:62847] = '{32'h4198e40b, 32'h42495a64, 32'hc2997bdd, 32'h4290cab6, 32'h423b7f7d, 32'h42450fce, 32'hc256faf9, 32'h42608f5f};
test_output[7855] = '{32'h4290cab6};
test_index[7855] = '{3};
test_input[62848:62855] = '{32'h42091c60, 32'h4280af7c, 32'h41a506af, 32'hc1da6962, 32'h42bb3eec, 32'h40caad1b, 32'hc22e2136, 32'h42acb133};
test_output[7856] = '{32'h42bb3eec};
test_index[7856] = '{4};
test_input[62856:62863] = '{32'hc20b555e, 32'h422c7ff0, 32'hc0e7efa2, 32'hc28ec3df, 32'hc25d881f, 32'hc293d2e5, 32'hc1b40122, 32'h42c71ac2};
test_output[7857] = '{32'h42c71ac2};
test_index[7857] = '{7};
test_input[62864:62871] = '{32'hc16a3082, 32'h413fc50d, 32'hc27266da, 32'hc27604f6, 32'h42a143d1, 32'h42bab1c2, 32'hbf93858b, 32'h42245bfd};
test_output[7858] = '{32'h42bab1c2};
test_index[7858] = '{5};
test_input[62872:62879] = '{32'h405ec67e, 32'h418ea6cb, 32'hc1e9b6e5, 32'h42a566c9, 32'h40b7e9a7, 32'h427e84ee, 32'hc23c5ab2, 32'h40a93025};
test_output[7859] = '{32'h42a566c9};
test_index[7859] = '{3};
test_input[62880:62887] = '{32'h4268c641, 32'hc248a770, 32'hc00f2ec4, 32'h4299e091, 32'h41854b97, 32'h42595be2, 32'hc1d31710, 32'hc0b90e60};
test_output[7860] = '{32'h4299e091};
test_index[7860] = '{3};
test_input[62888:62895] = '{32'hc1eb29e0, 32'h420953a5, 32'hc24344f5, 32'h42a4c878, 32'hc2c67ed8, 32'h409c90d1, 32'hc1bbc8d8, 32'h4216596a};
test_output[7861] = '{32'h42a4c878};
test_index[7861] = '{3};
test_input[62896:62903] = '{32'hc19ad590, 32'hc27be028, 32'hc22f5525, 32'h42c5df64, 32'h426ac8ef, 32'h423e47ee, 32'h421757e4, 32'h42a9a49e};
test_output[7862] = '{32'h42c5df64};
test_index[7862] = '{3};
test_input[62904:62911] = '{32'h42b4beee, 32'h42103840, 32'h4298bbad, 32'h41ef245e, 32'hc286b0e4, 32'hc0b83f94, 32'hc285cf51, 32'h42777cd6};
test_output[7863] = '{32'h42b4beee};
test_index[7863] = '{0};
test_input[62912:62919] = '{32'h4157fc86, 32'h428e86a4, 32'h4296d79f, 32'hc18587d2, 32'hc1bbbb08, 32'h429d8876, 32'h42581715, 32'h42ae8391};
test_output[7864] = '{32'h42ae8391};
test_index[7864] = '{7};
test_input[62920:62927] = '{32'hc138ebbe, 32'h4236956a, 32'h419275e3, 32'h42464de2, 32'h42266b91, 32'hc0ce2f7f, 32'h41842a94, 32'hc2b40578};
test_output[7865] = '{32'h42464de2};
test_index[7865] = '{3};
test_input[62928:62935] = '{32'h422ab01f, 32'h423bec07, 32'h422b510b, 32'hc1fb2ee2, 32'hc27a9533, 32'h415cec46, 32'hc2a242a8, 32'h429dd994};
test_output[7866] = '{32'h429dd994};
test_index[7866] = '{7};
test_input[62936:62943] = '{32'hc2bae57e, 32'hc2af6410, 32'hc29a1c8d, 32'h4216f3ae, 32'hc0914c72, 32'hc295d1fb, 32'hc2a7f056, 32'hc1f34adb};
test_output[7867] = '{32'h4216f3ae};
test_index[7867] = '{3};
test_input[62944:62951] = '{32'h42b6d5ff, 32'h42afb802, 32'hc1f95674, 32'h42166654, 32'h429087bd, 32'h4188e176, 32'h423eb427, 32'h418f0604};
test_output[7868] = '{32'h42b6d5ff};
test_index[7868] = '{0};
test_input[62952:62959] = '{32'hc2439931, 32'hc2330d48, 32'hc1b51b38, 32'hc2182e88, 32'hc19e08df, 32'hc26cf351, 32'h420a2e27, 32'hc25b07ee};
test_output[7869] = '{32'h420a2e27};
test_index[7869] = '{6};
test_input[62960:62967] = '{32'h41491614, 32'h4203d19f, 32'h429aad14, 32'hc2bbaa69, 32'hc2a648c7, 32'hc2be45f6, 32'hc2984313, 32'hc1ba6794};
test_output[7870] = '{32'h429aad14};
test_index[7870] = '{2};
test_input[62968:62975] = '{32'hc207dca8, 32'hc23e8669, 32'hc21f3cc9, 32'hc1f98e44, 32'hc2043fb2, 32'hc2855b1a, 32'hc22e6f2b, 32'hc2177091};
test_output[7871] = '{32'hc1f98e44};
test_index[7871] = '{3};
test_input[62976:62983] = '{32'h42445488, 32'hc1c77615, 32'hc2a746f0, 32'h42825b68, 32'h42a02315, 32'hc2c6a0bf, 32'hc04c1d7c, 32'h42aa7f31};
test_output[7872] = '{32'h42aa7f31};
test_index[7872] = '{7};
test_input[62984:62991] = '{32'h42b9ac91, 32'hc2a184f4, 32'h40f972bc, 32'h429d5f73, 32'h4297ad29, 32'h426984d8, 32'hc1af0dd1, 32'hc1f7b470};
test_output[7873] = '{32'h42b9ac91};
test_index[7873] = '{0};
test_input[62992:62999] = '{32'hc2a42135, 32'hc2c641dd, 32'h429e5f1b, 32'h426ba0f6, 32'h413f3452, 32'hc2240a5a, 32'h42b953ed, 32'hc297e1e1};
test_output[7874] = '{32'h42b953ed};
test_index[7874] = '{6};
test_input[63000:63007] = '{32'h42c26a26, 32'hc29b4de2, 32'hc22cb55e, 32'hc2868cb9, 32'h428ac8fb, 32'hc2a94ed2, 32'h4233ef11, 32'hc1068535};
test_output[7875] = '{32'h42c26a26};
test_index[7875] = '{0};
test_input[63008:63015] = '{32'h420e2adc, 32'hc1f584d5, 32'h4217fddf, 32'hc22bb119, 32'h42484512, 32'h422c596b, 32'h41891c2c, 32'hc14e4fa8};
test_output[7876] = '{32'h42484512};
test_index[7876] = '{4};
test_input[63016:63023] = '{32'hc2b2d16b, 32'hc2885ab3, 32'h40e0e71e, 32'hc23022fc, 32'h412dfe0c, 32'hc2a6ff09, 32'h42a65fc7, 32'hc292c435};
test_output[7877] = '{32'h42a65fc7};
test_index[7877] = '{6};
test_input[63024:63031] = '{32'h424d7585, 32'hc2c3ce34, 32'hc24d57d1, 32'h429c5487, 32'hc1b9e6ae, 32'hc255c0e4, 32'h3fe0b29e, 32'h426ef9e4};
test_output[7878] = '{32'h429c5487};
test_index[7878] = '{3};
test_input[63032:63039] = '{32'hc0cb1fd0, 32'hc1b996a9, 32'h3ff0e6c0, 32'hc19c998d, 32'hc274d1a4, 32'hc29b09f7, 32'h42ba28c7, 32'h423d8060};
test_output[7879] = '{32'h42ba28c7};
test_index[7879] = '{6};
test_input[63040:63047] = '{32'h4264d8ad, 32'hc2933f56, 32'hc168bdf4, 32'h42625cc1, 32'hc0b6f199, 32'h428e6c4c, 32'h42534193, 32'hc26127af};
test_output[7880] = '{32'h428e6c4c};
test_index[7880] = '{5};
test_input[63048:63055] = '{32'hc1a45250, 32'h42af00ca, 32'hc1a532c4, 32'h4214ffcb, 32'hc2a47f21, 32'h424ed7dd, 32'h42a7555f, 32'hc2b3528c};
test_output[7881] = '{32'h42af00ca};
test_index[7881] = '{1};
test_input[63056:63063] = '{32'h4225f434, 32'hc1bac93f, 32'h41b445ae, 32'hc27703f5, 32'h42bafa75, 32'hc204a148, 32'hc1952030, 32'hc23f5764};
test_output[7882] = '{32'h42bafa75};
test_index[7882] = '{4};
test_input[63064:63071] = '{32'h4247b7b5, 32'hbf65c784, 32'hc25989ee, 32'h41ab2e95, 32'h42953205, 32'h42b106bc, 32'h42221d4d, 32'hc215932b};
test_output[7883] = '{32'h42b106bc};
test_index[7883] = '{5};
test_input[63072:63079] = '{32'h42a80358, 32'h4235b1cc, 32'hc275b4f5, 32'hc2b4b3aa, 32'h4226545a, 32'hc28a6f21, 32'h42c60bcf, 32'hc1faa568};
test_output[7884] = '{32'h42c60bcf};
test_index[7884] = '{6};
test_input[63080:63087] = '{32'h420c9f8e, 32'hc29cab87, 32'h413fe94b, 32'h4281ed95, 32'h417ded67, 32'h4182f366, 32'hc2aa7c4d, 32'hc2a234d1};
test_output[7885] = '{32'h4281ed95};
test_index[7885] = '{3};
test_input[63088:63095] = '{32'hc16ae80e, 32'hc27b0975, 32'h41cec5dc, 32'hc16ab7f8, 32'h4262c13f, 32'h42c265d4, 32'h422dcf1f, 32'h42ad7776};
test_output[7886] = '{32'h42c265d4};
test_index[7886] = '{5};
test_input[63096:63103] = '{32'h41cdfc9e, 32'h42a0a61b, 32'h429d744d, 32'hc247de0f, 32'h408df8e3, 32'hc2085afd, 32'h427c0464, 32'h41ece4cf};
test_output[7887] = '{32'h42a0a61b};
test_index[7887] = '{1};
test_input[63104:63111] = '{32'hc11e9bfb, 32'h417a5476, 32'hc2bd0d00, 32'hc2287275, 32'hc2311f57, 32'h424391bd, 32'h42c11b92, 32'h42bece2b};
test_output[7888] = '{32'h42c11b92};
test_index[7888] = '{6};
test_input[63112:63119] = '{32'h428a5992, 32'h42292715, 32'h419e3482, 32'h41c5c205, 32'h42ab22ba, 32'h42872b23, 32'h42476c5f, 32'h4242af55};
test_output[7889] = '{32'h42ab22ba};
test_index[7889] = '{4};
test_input[63120:63127] = '{32'h41d5f9b5, 32'hc22b8dc5, 32'hc1a40ff3, 32'h428fac1f, 32'hc291b63d, 32'h42b4cdff, 32'hc267fd32, 32'hc1a2a30f};
test_output[7890] = '{32'h42b4cdff};
test_index[7890] = '{5};
test_input[63128:63135] = '{32'hc1967d7f, 32'h42871491, 32'hc2a42e1c, 32'h42373640, 32'hc21b8fad, 32'hc0aec10f, 32'h42603063, 32'hc2362b3d};
test_output[7891] = '{32'h42871491};
test_index[7891] = '{1};
test_input[63136:63143] = '{32'h4219d404, 32'h4232d34e, 32'hc22e0d0c, 32'hc0d4c0ac, 32'hc2a345f5, 32'h429e4ddd, 32'hc256daf5, 32'h4286897e};
test_output[7892] = '{32'h429e4ddd};
test_index[7892] = '{5};
test_input[63144:63151] = '{32'hc2525dd3, 32'hc20df40e, 32'hc20ba9ff, 32'h421bc100, 32'h425d60bb, 32'hc240a4b3, 32'h42bfc00e, 32'h41805c02};
test_output[7893] = '{32'h42bfc00e};
test_index[7893] = '{6};
test_input[63152:63159] = '{32'h41b391d9, 32'hc2aacc9e, 32'hc28cf0b5, 32'hc1a90e07, 32'hc235f09c, 32'h406856f4, 32'h42835127, 32'h42550ae7};
test_output[7894] = '{32'h42835127};
test_index[7894] = '{6};
test_input[63160:63167] = '{32'h42217345, 32'hc1223497, 32'h42834329, 32'hc1d05641, 32'h41afbd39, 32'h40d37a59, 32'hc281cbfa, 32'hc25cf97a};
test_output[7895] = '{32'h42834329};
test_index[7895] = '{2};
test_input[63168:63175] = '{32'hc2c72c40, 32'h41b5c9ee, 32'h429dcc2f, 32'hc299a11e, 32'h418b9348, 32'h42278703, 32'h41cb0880, 32'h40a143e3};
test_output[7896] = '{32'h429dcc2f};
test_index[7896] = '{2};
test_input[63176:63183] = '{32'h42859cd3, 32'h42b7d6e2, 32'h4133cd57, 32'h41de2397, 32'hc16c69c0, 32'h425a21c6, 32'h423e3cfe, 32'hc2c6c94e};
test_output[7897] = '{32'h42b7d6e2};
test_index[7897] = '{1};
test_input[63184:63191] = '{32'hc28397f9, 32'hc288ca96, 32'h41f716c8, 32'h42347b27, 32'h42bc7cb2, 32'h4292ce94, 32'h41dfc713, 32'h429158ab};
test_output[7898] = '{32'h42bc7cb2};
test_index[7898] = '{4};
test_input[63192:63199] = '{32'hc2785630, 32'hc1cda1f7, 32'hc195f9af, 32'hc2b27d0f, 32'h40d930c1, 32'h4196d798, 32'hc2946757, 32'h426a2de7};
test_output[7899] = '{32'h426a2de7};
test_index[7899] = '{7};
test_input[63200:63207] = '{32'h41a5efd0, 32'h3ffca8b4, 32'h4246ecf1, 32'h429d2e88, 32'hc1b46c28, 32'hc29b355f, 32'hc2b1cc47, 32'hc29c7445};
test_output[7900] = '{32'h429d2e88};
test_index[7900] = '{3};
test_input[63208:63215] = '{32'h41950069, 32'hc1dcbb0d, 32'hc2b413ae, 32'h426ecc09, 32'hc20977d2, 32'hc12f0956, 32'hc2675080, 32'hc2b36721};
test_output[7901] = '{32'h426ecc09};
test_index[7901] = '{3};
test_input[63216:63223] = '{32'h421767f9, 32'h42c3566f, 32'hc1a1c836, 32'h42a293d8, 32'h42949287, 32'h42a1ea55, 32'hc2c4e20a, 32'hc29c57c1};
test_output[7902] = '{32'h42c3566f};
test_index[7902] = '{1};
test_input[63224:63231] = '{32'h41da529b, 32'h4180953b, 32'h42a8a847, 32'hc221b312, 32'hc2c66900, 32'hc2b28a84, 32'h42b69ab2, 32'hc23d3bef};
test_output[7903] = '{32'h42b69ab2};
test_index[7903] = '{6};
test_input[63232:63239] = '{32'hc277ba8b, 32'h41f88b07, 32'h41acbc5d, 32'hc2aadab3, 32'hc24dee2b, 32'hc1f512e7, 32'hc26fdb20, 32'hbf9d2b2e};
test_output[7904] = '{32'h41f88b07};
test_index[7904] = '{1};
test_input[63240:63247] = '{32'h42507b98, 32'hc24c576d, 32'hc1a049fc, 32'h424b375f, 32'hc1a9b6f2, 32'hc24213be, 32'h42356cea, 32'hc26971f3};
test_output[7905] = '{32'h42507b98};
test_index[7905] = '{0};
test_input[63248:63255] = '{32'hc2ab694b, 32'h414e61bc, 32'h41f2f584, 32'hc27460d3, 32'h42c773f0, 32'hc2891985, 32'h4212ccb4, 32'hc2ba43ed};
test_output[7906] = '{32'h42c773f0};
test_index[7906] = '{4};
test_input[63256:63263] = '{32'hc206580d, 32'h429c038a, 32'hc2a481ca, 32'h42934314, 32'h420c9a56, 32'h41a96fd2, 32'h3dc4d882, 32'h425b3754};
test_output[7907] = '{32'h429c038a};
test_index[7907] = '{1};
test_input[63264:63271] = '{32'hc0bf1873, 32'hc22db2fa, 32'hc0fe2553, 32'hc227c82c, 32'h4223def4, 32'hc24b843b, 32'hc2693c67, 32'hc24c42c9};
test_output[7908] = '{32'h4223def4};
test_index[7908] = '{4};
test_input[63272:63279] = '{32'hc234d244, 32'h41bafd74, 32'h426c5917, 32'h41e80a21, 32'h42a00a22, 32'hc10951c7, 32'h41822a2c, 32'hc1a1aeeb};
test_output[7909] = '{32'h42a00a22};
test_index[7909] = '{4};
test_input[63280:63287] = '{32'h41122410, 32'hc24a4d6c, 32'h41fb732f, 32'h42bbe686, 32'hc0312f52, 32'hc244314f, 32'h41c5fa06, 32'hc2866fbe};
test_output[7910] = '{32'h42bbe686};
test_index[7910] = '{3};
test_input[63288:63295] = '{32'hc295cf95, 32'h4230566d, 32'h3fa57f31, 32'hc29d4af3, 32'hc20c46dd, 32'h427757fe, 32'h417144c7, 32'hc20d09b2};
test_output[7911] = '{32'h427757fe};
test_index[7911] = '{5};
test_input[63296:63303] = '{32'hc2c6b832, 32'h42273e1d, 32'hc12d2b00, 32'hc2c68930, 32'hc2a55d94, 32'h42c40ea9, 32'h412d422f, 32'hc1a59d35};
test_output[7912] = '{32'h42c40ea9};
test_index[7912] = '{5};
test_input[63304:63311] = '{32'hc29da32b, 32'hc20b85d7, 32'hc1b5ab75, 32'h420209db, 32'hc0bc73e9, 32'hc238f39c, 32'h4229eb30, 32'h42baa95f};
test_output[7913] = '{32'h42baa95f};
test_index[7913] = '{7};
test_input[63312:63319] = '{32'hc2bd4eee, 32'h4270460a, 32'h4280e4a2, 32'h41c645be, 32'h4260967d, 32'h4225231d, 32'hc2253349, 32'hc0b8c1ea};
test_output[7914] = '{32'h4280e4a2};
test_index[7914] = '{2};
test_input[63320:63327] = '{32'hc280741d, 32'hc0d69c8f, 32'hc27e083b, 32'hc2321ce8, 32'hbf121191, 32'h417712c4, 32'hc1f45e00, 32'hc279b377};
test_output[7915] = '{32'h417712c4};
test_index[7915] = '{5};
test_input[63328:63335] = '{32'hc102a361, 32'h42b0e806, 32'h42350ca7, 32'h42816938, 32'h4237a965, 32'h415b3123, 32'h41770d56, 32'h427525d3};
test_output[7916] = '{32'h42b0e806};
test_index[7916] = '{1};
test_input[63336:63343] = '{32'h42900992, 32'h42ab26fe, 32'hc2c3a6ba, 32'hc283543d, 32'hc2193ae7, 32'hc2acee12, 32'hc2253468, 32'hc287af39};
test_output[7917] = '{32'h42ab26fe};
test_index[7917] = '{1};
test_input[63344:63351] = '{32'hc2874121, 32'h4290901a, 32'hc28bec64, 32'h42998aad, 32'h42c4a3ff, 32'hc29f4f19, 32'hc2869bd5, 32'h421e27f6};
test_output[7918] = '{32'h42c4a3ff};
test_index[7918] = '{4};
test_input[63352:63359] = '{32'h3f7f57dd, 32'h42abffab, 32'h41ba143e, 32'hc2257f68, 32'hc2a030b7, 32'h41157709, 32'h42708459, 32'h426034bc};
test_output[7919] = '{32'h42abffab};
test_index[7919] = '{1};
test_input[63360:63367] = '{32'h41b1c3af, 32'h412d80a4, 32'hc19197b4, 32'hc197bf86, 32'hc24dea40, 32'h4215297a, 32'hc0bd7d33, 32'hc2727623};
test_output[7920] = '{32'h4215297a};
test_index[7920] = '{5};
test_input[63368:63375] = '{32'h424b712d, 32'hc270e694, 32'hc1fd6eaa, 32'hc2b90718, 32'h41ced5d6, 32'h42b38206, 32'hc1bd63b9, 32'hc1ab4ba6};
test_output[7921] = '{32'h42b38206};
test_index[7921] = '{5};
test_input[63376:63383] = '{32'hc2354437, 32'h41f44fd5, 32'h42aeffe4, 32'hc1fb4ba9, 32'h42032fec, 32'hc2446475, 32'hc23825cf, 32'h42ac2c3c};
test_output[7922] = '{32'h42aeffe4};
test_index[7922] = '{2};
test_input[63384:63391] = '{32'hc25f6441, 32'h42b0e5f3, 32'hc298d880, 32'h41febda4, 32'hc2929b1e, 32'hc22bac64, 32'hc200bd46, 32'hc1c42597};
test_output[7923] = '{32'h42b0e5f3};
test_index[7923] = '{1};
test_input[63392:63399] = '{32'hc202df86, 32'h42067757, 32'h42b7d410, 32'hc24ba9ef, 32'hc29713c3, 32'h41fdfd4e, 32'hc1cc9953, 32'h423ff59d};
test_output[7924] = '{32'h42b7d410};
test_index[7924] = '{2};
test_input[63400:63407] = '{32'hc2505170, 32'h4289f80f, 32'hc1df4053, 32'hc268416e, 32'hc22b42bd, 32'hc2a89fee, 32'hc256926f, 32'h408f47d8};
test_output[7925] = '{32'h4289f80f};
test_index[7925] = '{1};
test_input[63408:63415] = '{32'hc26583f4, 32'hc27a874c, 32'hc21381ac, 32'h416df918, 32'h42627270, 32'hc1915628, 32'hc2577e6b, 32'hc16c0e17};
test_output[7926] = '{32'h42627270};
test_index[7926] = '{4};
test_input[63416:63423] = '{32'h420e5614, 32'hc2b075b3, 32'hc1df8119, 32'hc192b93a, 32'h40ae41c7, 32'hc2c2a5f2, 32'h413e4e5a, 32'hc2c02f87};
test_output[7927] = '{32'h420e5614};
test_index[7927] = '{0};
test_input[63424:63431] = '{32'hc1921ca1, 32'hc2aa9a2c, 32'hc28cc0c6, 32'h4244bea5, 32'hc2862d84, 32'h42856477, 32'h429548c7, 32'hc22355ee};
test_output[7928] = '{32'h429548c7};
test_index[7928] = '{6};
test_input[63432:63439] = '{32'hc27d50c0, 32'hc2be2fd9, 32'h4062744b, 32'h42305aff, 32'hc220f3b4, 32'h4259533f, 32'hc2845796, 32'h4203d432};
test_output[7929] = '{32'h4259533f};
test_index[7929] = '{5};
test_input[63440:63447] = '{32'hc2a1ffa7, 32'h410c1783, 32'hc277b44a, 32'hc10317ea, 32'hbf2e2b36, 32'h41e93707, 32'h4045aee4, 32'h42b66cf2};
test_output[7930] = '{32'h42b66cf2};
test_index[7930] = '{7};
test_input[63448:63455] = '{32'hc1bb9ac0, 32'h412e3b1e, 32'hc1e4e141, 32'hc01d1627, 32'h418ca60c, 32'hc0d2eca2, 32'h429db711, 32'h41072832};
test_output[7931] = '{32'h429db711};
test_index[7931] = '{6};
test_input[63456:63463] = '{32'h41166497, 32'h40558547, 32'h426aa3a4, 32'hc143b766, 32'hc2a59629, 32'h42a64041, 32'hc1964efc, 32'hc2810045};
test_output[7932] = '{32'h42a64041};
test_index[7932] = '{5};
test_input[63464:63471] = '{32'h42848789, 32'h41946afd, 32'h41c444f6, 32'hc26c2dbb, 32'h422ceca4, 32'h424b39cc, 32'hc2805f0b, 32'hc0cce3c2};
test_output[7933] = '{32'h42848789};
test_index[7933] = '{0};
test_input[63472:63479] = '{32'h42ae6520, 32'h409c0991, 32'hc2937074, 32'h42054194, 32'h4247e395, 32'hc2b0bfbd, 32'h41d108d3, 32'hc1423e95};
test_output[7934] = '{32'h42ae6520};
test_index[7934] = '{0};
test_input[63480:63487] = '{32'hc1c8e6fb, 32'hc106e620, 32'hc2ae9409, 32'hc13784f1, 32'hc28694ad, 32'hc2b22715, 32'hc292ec62, 32'h42b26d0f};
test_output[7935] = '{32'h42b26d0f};
test_index[7935] = '{7};
test_input[63488:63495] = '{32'hc2bafe86, 32'h41fe6c7d, 32'h425529fb, 32'hc2a873a8, 32'h4287a215, 32'h41b4428e, 32'hc282bf6b, 32'h41d440ee};
test_output[7936] = '{32'h4287a215};
test_index[7936] = '{4};
test_input[63496:63503] = '{32'hc1e4ed3f, 32'hc18337e9, 32'hc29502ee, 32'hc2678793, 32'h429eba1f, 32'h412d916d, 32'hc2c5f313, 32'h41bbe5cc};
test_output[7937] = '{32'h429eba1f};
test_index[7937] = '{4};
test_input[63504:63511] = '{32'h4277b033, 32'hc22173cb, 32'hc234a7d6, 32'h42c7be8e, 32'h41a99c81, 32'hc0e9b8a6, 32'h41834c8e, 32'hc17449b0};
test_output[7938] = '{32'h42c7be8e};
test_index[7938] = '{3};
test_input[63512:63519] = '{32'hc272d255, 32'hc2348520, 32'hc28751d6, 32'hc211bad8, 32'h42a672b1, 32'h41b65f4b, 32'hc20abb76, 32'hc228113e};
test_output[7939] = '{32'h42a672b1};
test_index[7939] = '{4};
test_input[63520:63527] = '{32'hc20ae710, 32'hc2c7e720, 32'h421d77eb, 32'hc18975cf, 32'h41912ea5, 32'h4097a162, 32'h42a64a73, 32'h429acdf3};
test_output[7940] = '{32'h42a64a73};
test_index[7940] = '{6};
test_input[63528:63535] = '{32'hc1dbedfe, 32'hc1a85728, 32'h42607d09, 32'h41bdf911, 32'h42910d96, 32'hc27ddf7f, 32'h42bfcb9e, 32'hc1a21da1};
test_output[7941] = '{32'h42bfcb9e};
test_index[7941] = '{6};
test_input[63536:63543] = '{32'h41ffb945, 32'hc271b7ed, 32'hc1221014, 32'h4224321a, 32'h427f1bcf, 32'h423f8bfe, 32'hc29c6b8f, 32'hc22a09ed};
test_output[7942] = '{32'h427f1bcf};
test_index[7942] = '{4};
test_input[63544:63551] = '{32'h42ba232c, 32'h4250e8e7, 32'hc2af6197, 32'h41d7aa21, 32'h420a520d, 32'hc20ff4f0, 32'h423ce204, 32'h42b2efd8};
test_output[7943] = '{32'h42ba232c};
test_index[7943] = '{0};
test_input[63552:63559] = '{32'h41bca23b, 32'hc24feaaa, 32'h4229bf3a, 32'hc298e4d9, 32'h40adeb6a, 32'h4296b3d6, 32'h42174a1e, 32'hbe90654b};
test_output[7944] = '{32'h4296b3d6};
test_index[7944] = '{5};
test_input[63560:63567] = '{32'hc15fcf8d, 32'hc26f5af3, 32'h429783cf, 32'hc222442e, 32'hc1c1a440, 32'hc2b642cf, 32'h427b5bd9, 32'h42b941a8};
test_output[7945] = '{32'h42b941a8};
test_index[7945] = '{7};
test_input[63568:63575] = '{32'h413c79fc, 32'hc280a9f5, 32'hc25e4ec1, 32'hc1e3e407, 32'hc24a265a, 32'h415cb1b6, 32'hc23cfe49, 32'hc2b15d04};
test_output[7946] = '{32'h415cb1b6};
test_index[7946] = '{5};
test_input[63576:63583] = '{32'h4289eb00, 32'h4246706c, 32'h42576e92, 32'hc2b171ab, 32'hc1e636b6, 32'hc03ccfdc, 32'hc2b67869, 32'hc142df8b};
test_output[7947] = '{32'h4289eb00};
test_index[7947] = '{0};
test_input[63584:63591] = '{32'h4266e079, 32'hc1266110, 32'hc1577236, 32'hc0d78d45, 32'hc1efcabf, 32'h422480fc, 32'hc19c2b5e, 32'h40b2efaf};
test_output[7948] = '{32'h4266e079};
test_index[7948] = '{0};
test_input[63592:63599] = '{32'h428060f0, 32'hc2b39e33, 32'hc2792137, 32'h42b37817, 32'hc0e750ea, 32'hc12c329a, 32'h41f1c9b9, 32'hc061a186};
test_output[7949] = '{32'h42b37817};
test_index[7949] = '{3};
test_input[63600:63607] = '{32'hc2c2f5f0, 32'hc2addd30, 32'h40e555d7, 32'hc239e745, 32'h41ca4c77, 32'hc10eef07, 32'hc2912af8, 32'hc242ae07};
test_output[7950] = '{32'h41ca4c77};
test_index[7950] = '{4};
test_input[63608:63615] = '{32'h42a42c27, 32'h4263e488, 32'hc02beaf3, 32'h4131d8a4, 32'h425981d0, 32'h42c0ea16, 32'hc28b4bfc, 32'h41f62b88};
test_output[7951] = '{32'h42c0ea16};
test_index[7951] = '{5};
test_input[63616:63623] = '{32'h4188b8a1, 32'h423620c0, 32'h4161fe49, 32'hc0e77863, 32'h42be142c, 32'h426ce6a6, 32'hc242e163, 32'h428b33fa};
test_output[7952] = '{32'h42be142c};
test_index[7952] = '{4};
test_input[63624:63631] = '{32'h415bc6b1, 32'h42a07b96, 32'hc218cd66, 32'h4074a59c, 32'hc15233ea, 32'h4255cc1d, 32'h423d795a, 32'hc26a0f4e};
test_output[7953] = '{32'h42a07b96};
test_index[7953] = '{1};
test_input[63632:63639] = '{32'h428c82cf, 32'h42a794bb, 32'hc2a34c3c, 32'hc243f962, 32'h41b3103c, 32'hc2a58867, 32'hc25903a0, 32'hc15e7952};
test_output[7954] = '{32'h42a794bb};
test_index[7954] = '{1};
test_input[63640:63647] = '{32'hc1adb39c, 32'hc28753e7, 32'h42a4001b, 32'h42716a57, 32'hc199e143, 32'hc2bd10f9, 32'h403c9f03, 32'h420ea4f7};
test_output[7955] = '{32'h42a4001b};
test_index[7955] = '{2};
test_input[63648:63655] = '{32'hc21b93e6, 32'h4033a0d1, 32'h40be6b6f, 32'h428748a1, 32'h42a78a90, 32'h418f1ea9, 32'h417d38ac, 32'hc21a6014};
test_output[7956] = '{32'h42a78a90};
test_index[7956] = '{4};
test_input[63656:63663] = '{32'hc24f700e, 32'h41a9e2d7, 32'hbeb7ff64, 32'h42409cbe, 32'hc2b09c0f, 32'h4236ea4b, 32'hc1a7c3bf, 32'hc17d5092};
test_output[7957] = '{32'h42409cbe};
test_index[7957] = '{3};
test_input[63664:63671] = '{32'h4296beeb, 32'hc13f8c14, 32'h409c3c45, 32'h4241d4bf, 32'h42b767ed, 32'h4119697c, 32'hc207a44b, 32'hc299f5f0};
test_output[7958] = '{32'h42b767ed};
test_index[7958] = '{4};
test_input[63672:63679] = '{32'hc2a21f87, 32'hc23e2480, 32'hc25cb0ff, 32'h429d573b, 32'h415de7bd, 32'hc2b95b5b, 32'hc1899764, 32'h42bfac7b};
test_output[7959] = '{32'h42bfac7b};
test_index[7959] = '{7};
test_input[63680:63687] = '{32'hc2923882, 32'h42852bab, 32'hc0a154c1, 32'hc0f8e5eb, 32'h42adfd29, 32'hc26836fd, 32'h42c1ce1d, 32'hc1849a17};
test_output[7960] = '{32'h42c1ce1d};
test_index[7960] = '{6};
test_input[63688:63695] = '{32'h42580623, 32'hc09dbaf1, 32'hc12867e9, 32'hc28430b4, 32'h4279e421, 32'h3fff3ba5, 32'hc2bf58c4, 32'hc222813e};
test_output[7961] = '{32'h4279e421};
test_index[7961] = '{4};
test_input[63696:63703] = '{32'h3fe04256, 32'h4040d928, 32'hc2a9afb1, 32'hc26ebf0f, 32'h4237d66c, 32'hc11b1140, 32'h423117ce, 32'hc282f9d2};
test_output[7962] = '{32'h4237d66c};
test_index[7962] = '{4};
test_input[63704:63711] = '{32'h42b24290, 32'h42a386e8, 32'h42b6f698, 32'hc209d5c9, 32'h4211be54, 32'h42b9a120, 32'h420618cf, 32'h423f9086};
test_output[7963] = '{32'h42b9a120};
test_index[7963] = '{5};
test_input[63712:63719] = '{32'hc2b9583c, 32'h41a0a2aa, 32'h41840985, 32'h41aa3f8e, 32'h429f15a9, 32'h429a4c99, 32'hc1f57d52, 32'h429cf8af};
test_output[7964] = '{32'h429f15a9};
test_index[7964] = '{4};
test_input[63720:63727] = '{32'h4230fe59, 32'h42934cf8, 32'hc2bfd63b, 32'hc1fd1305, 32'h42670033, 32'hc22d25e6, 32'h4258a67c, 32'hc26e3854};
test_output[7965] = '{32'h42934cf8};
test_index[7965] = '{1};
test_input[63728:63735] = '{32'hc13093d8, 32'h42aeb948, 32'h422a5d20, 32'hc1856318, 32'hc1de8586, 32'h41776608, 32'h41cdee65, 32'hc0aaa7c1};
test_output[7966] = '{32'h42aeb948};
test_index[7966] = '{1};
test_input[63736:63743] = '{32'h426e698f, 32'hc2097772, 32'h3fbd5eae, 32'hc2b88717, 32'hc291f95e, 32'hc208ff87, 32'hc0426289, 32'h428f4c67};
test_output[7967] = '{32'h428f4c67};
test_index[7967] = '{7};
test_input[63744:63751] = '{32'hc2bb4c70, 32'hc19b535d, 32'h3f4d5719, 32'h3f856a56, 32'hbeea6802, 32'hc28a511d, 32'hc0c2e27d, 32'hc2bc02f0};
test_output[7968] = '{32'h3f856a56};
test_index[7968] = '{3};
test_input[63752:63759] = '{32'h4202f220, 32'h40eefb61, 32'h41bd74c2, 32'hc26a7309, 32'h41b11ff8, 32'hc20dfb60, 32'h412dc753, 32'h415dc1d7};
test_output[7969] = '{32'h4202f220};
test_index[7969] = '{0};
test_input[63760:63767] = '{32'h4223635b, 32'hc2352c43, 32'hc2239c63, 32'h415a3efb, 32'hc2147844, 32'h41586c5a, 32'h422c0a47, 32'h4253ebcb};
test_output[7970] = '{32'h4253ebcb};
test_index[7970] = '{7};
test_input[63768:63775] = '{32'hc24a32c1, 32'h42b36e1d, 32'h42991661, 32'h429790f3, 32'h42bd46b4, 32'h429a886d, 32'hc13198c7, 32'h42450c7c};
test_output[7971] = '{32'h42bd46b4};
test_index[7971] = '{4};
test_input[63776:63783] = '{32'hc2c4df13, 32'hc1704032, 32'h4273653c, 32'hc2a081d6, 32'hc20dc1ae, 32'hc28b7e33, 32'h42649da0, 32'hc15c8e24};
test_output[7972] = '{32'h4273653c};
test_index[7972] = '{2};
test_input[63784:63791] = '{32'hc207e93e, 32'hc1617265, 32'h40265bf6, 32'h428839b7, 32'h429277dc, 32'hc13c7ce2, 32'h428268b0, 32'h422307a1};
test_output[7973] = '{32'h429277dc};
test_index[7973] = '{4};
test_input[63792:63799] = '{32'hc2992617, 32'hc1ea2487, 32'hc124b83c, 32'h422a69a7, 32'h42acc4bb, 32'h42858900, 32'hc24b5fd3, 32'hc20369b9};
test_output[7974] = '{32'h42acc4bb};
test_index[7974] = '{4};
test_input[63800:63807] = '{32'hc1c2ba49, 32'hc1a265cc, 32'hc1a1f237, 32'h41e08a33, 32'hc2515bcf, 32'hc281902d, 32'hc2348c82, 32'h419bdeb4};
test_output[7975] = '{32'h41e08a33};
test_index[7975] = '{3};
test_input[63808:63815] = '{32'h42ae50d8, 32'h42bbf177, 32'hbfdcb66b, 32'h42be02b9, 32'hc28618f2, 32'hc27a2226, 32'h428b99da, 32'h4162e6c5};
test_output[7976] = '{32'h42be02b9};
test_index[7976] = '{3};
test_input[63816:63823] = '{32'h421d2d35, 32'h4216b5fe, 32'h41f3f88d, 32'hc2587eb0, 32'h425b765f, 32'h428e0f9c, 32'hc08eb47e, 32'h422e7aa9};
test_output[7977] = '{32'h428e0f9c};
test_index[7977] = '{5};
test_input[63824:63831] = '{32'h42ba1644, 32'hc28dd7c6, 32'h41cefbff, 32'hc18a9da7, 32'h41100e95, 32'h42021e4b, 32'hc2943a91, 32'h42b6fba9};
test_output[7978] = '{32'h42ba1644};
test_index[7978] = '{0};
test_input[63832:63839] = '{32'h4290fc9a, 32'hc1e71f6b, 32'hc187e368, 32'h429e0712, 32'hc2a0cb8a, 32'h4214b907, 32'hc253c522, 32'hc2ba269d};
test_output[7979] = '{32'h429e0712};
test_index[7979] = '{3};
test_input[63840:63847] = '{32'hc0e590ce, 32'hc197443c, 32'h40200da5, 32'h42a84ebd, 32'hc2a6814c, 32'h429f8115, 32'h426d8f83, 32'hc26be6a6};
test_output[7980] = '{32'h42a84ebd};
test_index[7980] = '{3};
test_input[63848:63855] = '{32'h3f77de8e, 32'h420b3af2, 32'h42986908, 32'hc2c3fcc1, 32'hc191dd3c, 32'hc2b2dcf2, 32'hc281b04a, 32'hc2c6c7cf};
test_output[7981] = '{32'h42986908};
test_index[7981] = '{2};
test_input[63856:63863] = '{32'h42608329, 32'h42417039, 32'h4279c09d, 32'h42ad02a3, 32'hc1f9c836, 32'hc2a5f1f8, 32'hc1e03221, 32'hc2ab587a};
test_output[7982] = '{32'h42ad02a3};
test_index[7982] = '{3};
test_input[63864:63871] = '{32'hc20b7b77, 32'h42c46558, 32'h4164b3be, 32'h429a20b8, 32'hc2526db5, 32'hc298a829, 32'h4229acaf, 32'hc25c6f86};
test_output[7983] = '{32'h42c46558};
test_index[7983] = '{1};
test_input[63872:63879] = '{32'h4205b579, 32'hc24efc9f, 32'hc2a1c896, 32'hc1b7bb92, 32'h426a4fce, 32'h426a3152, 32'hc2a018c0, 32'hc2111ef3};
test_output[7984] = '{32'h426a4fce};
test_index[7984] = '{4};
test_input[63880:63887] = '{32'h428bada4, 32'hc1908c9a, 32'hc10abe85, 32'hc25282dc, 32'h427ca64b, 32'hc2a6a065, 32'hc1e31256, 32'hc280830f};
test_output[7985] = '{32'h428bada4};
test_index[7985] = '{0};
test_input[63888:63895] = '{32'hc1c2c0e0, 32'h429097a5, 32'hc2bc2f5e, 32'hc2b25f3d, 32'hc29163b0, 32'hc2657e2b, 32'hc2599da4, 32'h40ec473c};
test_output[7986] = '{32'h429097a5};
test_index[7986] = '{1};
test_input[63896:63903] = '{32'hc0fb0601, 32'h429ba3ad, 32'hc267d033, 32'hc1c60b77, 32'h426f8c84, 32'hc1f5bd29, 32'hc0909deb, 32'h42b8735d};
test_output[7987] = '{32'h42b8735d};
test_index[7987] = '{7};
test_input[63904:63911] = '{32'hc271e45d, 32'h4252df5b, 32'h42647356, 32'hc20b1f88, 32'hc2c71102, 32'h42257a9e, 32'hc2489e33, 32'hc2522164};
test_output[7988] = '{32'h42647356};
test_index[7988] = '{2};
test_input[63912:63919] = '{32'hc2972fcc, 32'hc25e886b, 32'h41a1e246, 32'h426bc074, 32'h42167669, 32'h42439085, 32'hbfdac5ef, 32'h4289e392};
test_output[7989] = '{32'h4289e392};
test_index[7989] = '{7};
test_input[63920:63927] = '{32'h42bfb2ad, 32'h42b04bca, 32'hc2b44b3d, 32'hc2be4feb, 32'hc2338369, 32'h42c4a60b, 32'h415cf0b5, 32'hc2b48ff1};
test_output[7990] = '{32'h42c4a60b};
test_index[7990] = '{5};
test_input[63928:63935] = '{32'h422c7a25, 32'h41d180f5, 32'hc2b8929e, 32'hc2a035d8, 32'h42c14089, 32'h41dfce5e, 32'hc2a179ef, 32'hc22aaeff};
test_output[7991] = '{32'h42c14089};
test_index[7991] = '{4};
test_input[63936:63943] = '{32'h408d57ab, 32'hc2c0ce57, 32'hc2941de4, 32'hc053bd3f, 32'h4276fb58, 32'h42c435bb, 32'h42349855, 32'h42739507};
test_output[7992] = '{32'h42c435bb};
test_index[7992] = '{5};
test_input[63944:63951] = '{32'hbfd15b39, 32'hc2add908, 32'hc2bf0b83, 32'hc1fcee8d, 32'h420df384, 32'h408c4cef, 32'h42982594, 32'h41b126f7};
test_output[7993] = '{32'h42982594};
test_index[7993] = '{6};
test_input[63952:63959] = '{32'hc2b78825, 32'hc29e429d, 32'hc219f956, 32'h426de2ed, 32'hc27ee1f3, 32'h42b252f2, 32'h4281acc6, 32'hc1a2c29e};
test_output[7994] = '{32'h42b252f2};
test_index[7994] = '{5};
test_input[63960:63967] = '{32'h41b3369c, 32'h42c44d57, 32'h429ddedd, 32'h42342aa0, 32'hc25235a3, 32'hc22fa209, 32'h4264db84, 32'h41c0af32};
test_output[7995] = '{32'h42c44d57};
test_index[7995] = '{1};
test_input[63968:63975] = '{32'h41665acb, 32'hc0c3b28f, 32'h423a83fd, 32'h41d64bb1, 32'hc20a7bd5, 32'hc1371fb1, 32'hc2095228, 32'h42afe656};
test_output[7996] = '{32'h42afe656};
test_index[7996] = '{7};
test_input[63976:63983] = '{32'h42a5fd8d, 32'h42146a6e, 32'h41d94df9, 32'hc255fb36, 32'hc2277b78, 32'h42168cb4, 32'hc249843c, 32'h42666abe};
test_output[7997] = '{32'h42a5fd8d};
test_index[7997] = '{0};
test_input[63984:63991] = '{32'h426c764a, 32'h41f24930, 32'h4175da71, 32'hc23ac3d0, 32'hc0b2116a, 32'hc149c420, 32'h42b4f3d7, 32'h4224cac7};
test_output[7998] = '{32'h42b4f3d7};
test_index[7998] = '{6};
test_input[63992:63999] = '{32'hc1742eb0, 32'hc286cc9b, 32'hc1df3fbc, 32'h42a854d0, 32'hc2587cd4, 32'h42879d88, 32'hc2ac8eff, 32'hc242ee26};
test_output[7999] = '{32'h42a854d0};
test_index[7999] = '{3};
test_input[64000:64007] = '{32'h41c3a0b9, 32'hc29fc042, 32'h4203acae, 32'h42a60e35, 32'h428e136c, 32'h4278dffb, 32'h422174d5, 32'hc1f42be8};
test_output[8000] = '{32'h42a60e35};
test_index[8000] = '{3};
test_input[64008:64015] = '{32'hc28e5656, 32'h4205513b, 32'hc20351d4, 32'hc18e1ef4, 32'h42b13798, 32'hc233b458, 32'hc2bde574, 32'hc2aaa654};
test_output[8001] = '{32'h42b13798};
test_index[8001] = '{4};
test_input[64016:64023] = '{32'hc2b3717f, 32'hc2751e82, 32'h422e8c76, 32'h42157f59, 32'h4123d036, 32'hc18fa17e, 32'h4212a48f, 32'h42b0878a};
test_output[8002] = '{32'h42b0878a};
test_index[8002] = '{7};
test_input[64024:64031] = '{32'hc29e1dc9, 32'h42bb0772, 32'hc23c9522, 32'h3f87f290, 32'h406a10c1, 32'h429b204b, 32'hc2c33951, 32'h425122ad};
test_output[8003] = '{32'h42bb0772};
test_index[8003] = '{1};
test_input[64032:64039] = '{32'h4277add6, 32'hc20aba62, 32'hc2969f64, 32'hc0344bca, 32'hc22c69b4, 32'hc02568b6, 32'hc1ddbd85, 32'h4284775c};
test_output[8004] = '{32'h4284775c};
test_index[8004] = '{7};
test_input[64040:64047] = '{32'hc2a9aae6, 32'h41cdd24f, 32'h41988c64, 32'hc1859900, 32'h419b9975, 32'h429b29fd, 32'h4236b8b9, 32'hc2097d35};
test_output[8005] = '{32'h429b29fd};
test_index[8005] = '{5};
test_input[64048:64055] = '{32'hc298e94f, 32'hc1a718b0, 32'hc107c4cb, 32'h423907b5, 32'hbff92a1c, 32'h423fe115, 32'hc1d7eb29, 32'h42516a2f};
test_output[8006] = '{32'h42516a2f};
test_index[8006] = '{7};
test_input[64056:64063] = '{32'hc25a9ef2, 32'h424bffc9, 32'hc1091847, 32'hc2b2b3d3, 32'h4297dca0, 32'hc28eeb04, 32'hc2929049, 32'hc28c30a5};
test_output[8007] = '{32'h4297dca0};
test_index[8007] = '{4};
test_input[64064:64071] = '{32'h427659d6, 32'h41fa53b0, 32'h42be4fc0, 32'h42107d20, 32'hc2b5bee8, 32'hc2c014a7, 32'h425785fc, 32'h40003db8};
test_output[8008] = '{32'h42be4fc0};
test_index[8008] = '{2};
test_input[64072:64079] = '{32'hc26361db, 32'hc2c6e579, 32'hc2bb091a, 32'hbef03b8b, 32'h429c44a0, 32'h41eca33a, 32'h426c7fef, 32'hc2c5491c};
test_output[8009] = '{32'h429c44a0};
test_index[8009] = '{4};
test_input[64080:64087] = '{32'hc26e0c5d, 32'hc2aaa479, 32'h428998cc, 32'hc1c5ece0, 32'h415f7727, 32'h40b95993, 32'hc2b5c9a6, 32'hc104eaee};
test_output[8010] = '{32'h428998cc};
test_index[8010] = '{2};
test_input[64088:64095] = '{32'h421ca6d0, 32'h4261c8df, 32'hc156b628, 32'hc283ae94, 32'hc2bba8ea, 32'hc26d49bd, 32'hc227e74c, 32'h420afc61};
test_output[8011] = '{32'h4261c8df};
test_index[8011] = '{1};
test_input[64096:64103] = '{32'hc2c35ae6, 32'hc1a9b55d, 32'h422390ab, 32'hc27b5cc1, 32'hc28f8e77, 32'hc1492393, 32'h429c190c, 32'h42235944};
test_output[8012] = '{32'h429c190c};
test_index[8012] = '{6};
test_input[64104:64111] = '{32'hc20fe596, 32'hc08801ab, 32'h41945979, 32'h4187787e, 32'hc19bf1ae, 32'h42b89003, 32'hc294915d, 32'hc1b34209};
test_output[8013] = '{32'h42b89003};
test_index[8013] = '{5};
test_input[64112:64119] = '{32'hc1c54492, 32'h42ae110f, 32'h422466d0, 32'hc26d3dbc, 32'h4290ee6d, 32'h424851c0, 32'h4198ad17, 32'hc1dab536};
test_output[8014] = '{32'h42ae110f};
test_index[8014] = '{1};
test_input[64120:64127] = '{32'h4155a34b, 32'hc1d7454e, 32'hc296c6c3, 32'h41c265ce, 32'h4278e251, 32'h42b567f8, 32'hc0645db3, 32'h428c82eb};
test_output[8015] = '{32'h42b567f8};
test_index[8015] = '{5};
test_input[64128:64135] = '{32'hc2788148, 32'hc2ac6de9, 32'hc1cb9b42, 32'hc1e6f435, 32'h41e69308, 32'hc1b9d6e5, 32'hc2917394, 32'hc2162291};
test_output[8016] = '{32'h41e69308};
test_index[8016] = '{4};
test_input[64136:64143] = '{32'h42bbf62e, 32'h4201e2e5, 32'hc1f753a7, 32'hc26c71c5, 32'hc1f6ae2d, 32'h42a805d2, 32'hc2a1b97c, 32'h4296aa30};
test_output[8017] = '{32'h42bbf62e};
test_index[8017] = '{0};
test_input[64144:64151] = '{32'h41a3ceba, 32'hc28ef2e7, 32'h42b052c5, 32'hc18c4e37, 32'hc0bdc382, 32'hc26428f9, 32'hc2bd5e6a, 32'h42a8e73a};
test_output[8018] = '{32'h42b052c5};
test_index[8018] = '{2};
test_input[64152:64159] = '{32'hc234e5a6, 32'hc26e9812, 32'h42562475, 32'h425fbb5e, 32'hc0eee3c2, 32'hc28dd067, 32'hc2903329, 32'h41b386c3};
test_output[8019] = '{32'h425fbb5e};
test_index[8019] = '{3};
test_input[64160:64167] = '{32'hc26f2e04, 32'hc29be4f6, 32'h41901633, 32'hc1f557d6, 32'h40c34d38, 32'hc25daec8, 32'h42981102, 32'hc28ead80};
test_output[8020] = '{32'h42981102};
test_index[8020] = '{6};
test_input[64168:64175] = '{32'h422cb3a3, 32'hc25f0336, 32'h41c74fec, 32'h42802ac1, 32'h4281a0be, 32'h42bf83c1, 32'hc249f06d, 32'hc2b1d980};
test_output[8021] = '{32'h42bf83c1};
test_index[8021] = '{5};
test_input[64176:64183] = '{32'hc265e436, 32'h413cac1e, 32'hc2ae8624, 32'hc2591148, 32'h422e129d, 32'hc21829c7, 32'h42adb3a7, 32'h42441f91};
test_output[8022] = '{32'h42adb3a7};
test_index[8022] = '{6};
test_input[64184:64191] = '{32'h404b476e, 32'hc20962ef, 32'h41cba799, 32'hc2818ecd, 32'h427f6e9d, 32'h3f6d32aa, 32'hc29679b5, 32'h42882362};
test_output[8023] = '{32'h42882362};
test_index[8023] = '{7};
test_input[64192:64199] = '{32'hc2b2a01f, 32'hc23b98b9, 32'hc295f48a, 32'h42bae2c6, 32'h42bada6b, 32'h420f5f16, 32'hc291793b, 32'hc23dbdaf};
test_output[8024] = '{32'h42bae2c6};
test_index[8024] = '{3};
test_input[64200:64207] = '{32'h4244645c, 32'hc29070a8, 32'hc1953257, 32'h40ffb798, 32'hc2c398f0, 32'h423d01f8, 32'h42b6e4e7, 32'hc2c0d5fb};
test_output[8025] = '{32'h42b6e4e7};
test_index[8025] = '{6};
test_input[64208:64215] = '{32'hc2921ce4, 32'h4175e688, 32'h421e2a8a, 32'h428e3a6a, 32'h426627aa, 32'hc28fc270, 32'h427886eb, 32'h4298544a};
test_output[8026] = '{32'h4298544a};
test_index[8026] = '{7};
test_input[64216:64223] = '{32'h42a5c31e, 32'hc22b5917, 32'h428a0936, 32'hc171a3b3, 32'h3f14d97f, 32'h4295c0ab, 32'h42103c42, 32'hc1f0a3b7};
test_output[8027] = '{32'h42a5c31e};
test_index[8027] = '{0};
test_input[64224:64231] = '{32'h42299375, 32'hc1d201e9, 32'h42b02325, 32'hc2939c7c, 32'hc2052b48, 32'h411ba556, 32'h42864bf6, 32'h428fdae7};
test_output[8028] = '{32'h42b02325};
test_index[8028] = '{2};
test_input[64232:64239] = '{32'h42b148ac, 32'hc24e3014, 32'hc2a5714c, 32'hc2821f7f, 32'hc2b4f126, 32'h426aa0fb, 32'hc2aa3e2e, 32'h42384a5e};
test_output[8029] = '{32'h42b148ac};
test_index[8029] = '{0};
test_input[64240:64247] = '{32'h42c5d053, 32'hc2b76227, 32'hc0014e82, 32'h42b2c5b2, 32'h42b26084, 32'h429b6684, 32'h41aaf463, 32'hc292a627};
test_output[8030] = '{32'h42c5d053};
test_index[8030] = '{0};
test_input[64248:64255] = '{32'h42665c0c, 32'h4111bfee, 32'h413761b8, 32'h41c82d76, 32'hc261eb5e, 32'h4183374a, 32'hc2145475, 32'hc0495962};
test_output[8031] = '{32'h42665c0c};
test_index[8031] = '{0};
test_input[64256:64263] = '{32'h4297ab79, 32'hc228d690, 32'h4142adcd, 32'hc2b24614, 32'hc1902d8b, 32'hc1b3daf3, 32'h42b4df5b, 32'hc2154bcc};
test_output[8032] = '{32'h42b4df5b};
test_index[8032] = '{6};
test_input[64264:64271] = '{32'h429b7702, 32'h42248605, 32'hc0f62ee3, 32'hc28f3d49, 32'hc2241946, 32'h42430f33, 32'hc2539310, 32'h42c3b42a};
test_output[8033] = '{32'h42c3b42a};
test_index[8033] = '{7};
test_input[64272:64279] = '{32'h4271af0d, 32'h41969a40, 32'hc291aec7, 32'h4230e251, 32'h4003f347, 32'hc194b8b8, 32'h42a106b4, 32'h42c4013e};
test_output[8034] = '{32'h42c4013e};
test_index[8034] = '{7};
test_input[64280:64287] = '{32'h4268d8d2, 32'h421e96ae, 32'h429b2f91, 32'hc18df94c, 32'hc2b7b63d, 32'hc1df6323, 32'h41d57a9b, 32'h42b8fa01};
test_output[8035] = '{32'h42b8fa01};
test_index[8035] = '{7};
test_input[64288:64295] = '{32'h429aaeb3, 32'hc2681661, 32'hc2a702d2, 32'h4265b50a, 32'h42a8743d, 32'h426e11e8, 32'hc2620607, 32'hc1ca2065};
test_output[8036] = '{32'h42a8743d};
test_index[8036] = '{4};
test_input[64296:64303] = '{32'h42bcb00e, 32'h42622b94, 32'h429236cb, 32'h42498cee, 32'hc2b85b8f, 32'h42772091, 32'h41898e68, 32'h4211d15b};
test_output[8037] = '{32'h42bcb00e};
test_index[8037] = '{0};
test_input[64304:64311] = '{32'hc1a1d8ed, 32'hc1145bf6, 32'hc2b2bc4d, 32'hc17d775e, 32'h4244269b, 32'hc2b35008, 32'hc1e29416, 32'hc2ba8965};
test_output[8038] = '{32'h4244269b};
test_index[8038] = '{4};
test_input[64312:64319] = '{32'h41f6c70c, 32'h421a4ea7, 32'hc2512711, 32'hc27f188c, 32'hc296ef22, 32'hc1c02661, 32'hc29d1c2f, 32'h42b324dd};
test_output[8039] = '{32'h42b324dd};
test_index[8039] = '{7};
test_input[64320:64327] = '{32'h42915cb4, 32'hc2856113, 32'hc23c77b6, 32'hc28ccd62, 32'hc1da41b4, 32'h428cc98a, 32'h429e1ec9, 32'h428cf428};
test_output[8040] = '{32'h429e1ec9};
test_index[8040] = '{6};
test_input[64328:64335] = '{32'hc29cd66a, 32'hc1902cf8, 32'h41268396, 32'h427a8e71, 32'hc2bdce47, 32'h422df26e, 32'hc2270f46, 32'hc2be3b85};
test_output[8041] = '{32'h427a8e71};
test_index[8041] = '{3};
test_input[64336:64343] = '{32'h41637575, 32'hc149c356, 32'h4207b866, 32'hc2b054a3, 32'hc2930d7e, 32'h4289c760, 32'h4281b537, 32'hc0568d59};
test_output[8042] = '{32'h4289c760};
test_index[8042] = '{5};
test_input[64344:64351] = '{32'hc21158a9, 32'hc12d7375, 32'hc28a5a0e, 32'h424c3871, 32'hc261d6e2, 32'h42a55442, 32'hbf9f7918, 32'hc20b0808};
test_output[8043] = '{32'h42a55442};
test_index[8043] = '{5};
test_input[64352:64359] = '{32'hc1fb63d9, 32'h42a814bf, 32'h42b7452e, 32'hc2795336, 32'hc1b9d3db, 32'h42b8dc59, 32'hc2856bfe, 32'h42a8bf0b};
test_output[8044] = '{32'h42b8dc59};
test_index[8044] = '{5};
test_input[64360:64367] = '{32'h40750526, 32'hc1ece847, 32'hc253ded8, 32'h42ab7b4b, 32'hc280b751, 32'hc1ed841d, 32'hc2abece6, 32'h42964b05};
test_output[8045] = '{32'h42ab7b4b};
test_index[8045] = '{3};
test_input[64368:64375] = '{32'hc28925a4, 32'hc1486ec8, 32'h427ffaca, 32'h42649d6d, 32'h42762c26, 32'hc24ea76d, 32'h426a7383, 32'hc29fdaf1};
test_output[8046] = '{32'h427ffaca};
test_index[8046] = '{2};
test_input[64376:64383] = '{32'hc2637b49, 32'hbea06612, 32'hc21f3b34, 32'hc220820f, 32'hc0911028, 32'hc28d5dbe, 32'hc095ccf4, 32'h42c316b0};
test_output[8047] = '{32'h42c316b0};
test_index[8047] = '{7};
test_input[64384:64391] = '{32'hc1a67685, 32'hc21d478c, 32'h40677675, 32'h42bf1ac5, 32'h425c7dd7, 32'h42bc2909, 32'hc0c59419, 32'h4291c5b9};
test_output[8048] = '{32'h42bf1ac5};
test_index[8048] = '{3};
test_input[64392:64399] = '{32'h42b584cc, 32'h417edd56, 32'h40b51dae, 32'hc28d04a9, 32'h423c90e6, 32'h424ae9b7, 32'hc245ab14, 32'hc28e3fc4};
test_output[8049] = '{32'h42b584cc};
test_index[8049] = '{0};
test_input[64400:64407] = '{32'hc1b31cfd, 32'hc2ad87a2, 32'h424d00aa, 32'h41b68024, 32'hc237a003, 32'hc11d7690, 32'hc29952a5, 32'hc2c6af48};
test_output[8050] = '{32'h424d00aa};
test_index[8050] = '{2};
test_input[64408:64415] = '{32'hc1a85f25, 32'h428aba6c, 32'h428ab42c, 32'h42bb0b9b, 32'hc22b68c4, 32'hc29978f4, 32'h41964c95, 32'h41f54fb1};
test_output[8051] = '{32'h42bb0b9b};
test_index[8051] = '{3};
test_input[64416:64423] = '{32'hc250c8e1, 32'h418ec00a, 32'h3fe8e310, 32'h4284ab7d, 32'hc2aac11c, 32'h4227c8aa, 32'hc232334d, 32'h41c30f6a};
test_output[8052] = '{32'h4284ab7d};
test_index[8052] = '{3};
test_input[64424:64431] = '{32'h40a633cd, 32'h424440ed, 32'hc18ead6e, 32'h42156200, 32'h4241c75b, 32'hc28cb02c, 32'hc28eb2df, 32'h42c7556d};
test_output[8053] = '{32'h42c7556d};
test_index[8053] = '{7};
test_input[64432:64439] = '{32'h4231154d, 32'hc2b7fa0d, 32'hc218ca04, 32'hc26b1032, 32'h41906601, 32'hc2c13fb7, 32'h42a3bb04, 32'h42aa7494};
test_output[8054] = '{32'h42aa7494};
test_index[8054] = '{7};
test_input[64440:64447] = '{32'h41ac52a2, 32'h42967ca1, 32'hc14d63d3, 32'hc1f4c94b, 32'h41ebbc7c, 32'hc197b365, 32'h427c1355, 32'h4093638b};
test_output[8055] = '{32'h42967ca1};
test_index[8055] = '{1};
test_input[64448:64455] = '{32'h415a7065, 32'h424b8e6c, 32'hc1c8888a, 32'hc25d34cb, 32'h42076707, 32'hc2acf8e7, 32'hc291eac2, 32'h41cb689d};
test_output[8056] = '{32'h424b8e6c};
test_index[8056] = '{1};
test_input[64456:64463] = '{32'hc23582ed, 32'hc0f387bd, 32'h41eed8b8, 32'h412c041c, 32'h4245a16a, 32'hc296c982, 32'h4227b4da, 32'hc233dcc0};
test_output[8057] = '{32'h4245a16a};
test_index[8057] = '{4};
test_input[64464:64471] = '{32'h40076b4d, 32'h42895261, 32'h42937bd8, 32'hc29149a1, 32'hc1867e57, 32'h42bbbf91, 32'hc13c3218, 32'hc2626c4e};
test_output[8058] = '{32'h42bbbf91};
test_index[8058] = '{5};
test_input[64472:64479] = '{32'hbfefb957, 32'hc2078fd0, 32'h429864c6, 32'hc21d5627, 32'hc0a1327e, 32'hc0f35883, 32'h422813de, 32'h4209a900};
test_output[8059] = '{32'h429864c6};
test_index[8059] = '{2};
test_input[64480:64487] = '{32'h42bfe6a7, 32'hc1a24c77, 32'hc2bb1ab8, 32'h42887a47, 32'h4210c82b, 32'hc14a3216, 32'hc24d6043, 32'h426b9a8e};
test_output[8060] = '{32'h42bfe6a7};
test_index[8060] = '{0};
test_input[64488:64495] = '{32'h423075aa, 32'hc29daf5e, 32'h41a0e8ef, 32'h4242cf96, 32'h4189ab10, 32'h4135b12c, 32'hc18c1995, 32'hc1604f80};
test_output[8061] = '{32'h4242cf96};
test_index[8061] = '{3};
test_input[64496:64503] = '{32'h42bb568b, 32'h42bd81e2, 32'h4265f5b9, 32'h41fe972b, 32'hc250be06, 32'h42b252f7, 32'h40ea00d9, 32'h427cbee7};
test_output[8062] = '{32'h42bd81e2};
test_index[8062] = '{1};
test_input[64504:64511] = '{32'h4143b3d2, 32'h42a69cb4, 32'hc228ad9a, 32'hc2c289fe, 32'hc0aa9213, 32'h424041a7, 32'h3fbce45d, 32'h41f89e3e};
test_output[8063] = '{32'h42a69cb4};
test_index[8063] = '{1};
test_input[64512:64519] = '{32'hc24e2ae6, 32'hc2c79ab1, 32'hc2302317, 32'hc2bd911e, 32'hc2c0eb60, 32'h420d5745, 32'h417f8b16, 32'h42c465b4};
test_output[8064] = '{32'h42c465b4};
test_index[8064] = '{7};
test_input[64520:64527] = '{32'h423d5418, 32'h42a76d40, 32'h4285aa63, 32'hc1ed77cc, 32'hc288fab4, 32'h42b8522e, 32'hc2b3543e, 32'hc23d4bce};
test_output[8065] = '{32'h42b8522e};
test_index[8065] = '{5};
test_input[64528:64535] = '{32'h42a29f47, 32'hc1ab94f4, 32'hc2c52761, 32'hc21cfe5a, 32'hc2b6cf24, 32'h42c2bb35, 32'hc2aff340, 32'hc0dbf51e};
test_output[8066] = '{32'h42c2bb35};
test_index[8066] = '{5};
test_input[64536:64543] = '{32'h42a612ec, 32'h420dc376, 32'hc2bfc7d3, 32'hc1c17f65, 32'h40fd515e, 32'hc20e352d, 32'h424cdb07, 32'h429c504b};
test_output[8067] = '{32'h42a612ec};
test_index[8067] = '{0};
test_input[64544:64551] = '{32'h41f60523, 32'h41fe52f4, 32'hc2869c7c, 32'hc281fbbb, 32'h42745f18, 32'hc26181ae, 32'h429b7e10, 32'h41c5f207};
test_output[8068] = '{32'h429b7e10};
test_index[8068] = '{6};
test_input[64552:64559] = '{32'hc242ffd7, 32'h408b6ed0, 32'hc1539a24, 32'h41e62b7f, 32'hc24ba798, 32'hc19bfd8d, 32'hc296389a, 32'h42b80c8b};
test_output[8069] = '{32'h42b80c8b};
test_index[8069] = '{7};
test_input[64560:64567] = '{32'h419dcd12, 32'hc1a26547, 32'h421ece1c, 32'hc2abed86, 32'hc1d35498, 32'h4185a928, 32'hc268ee84, 32'h420ea7c5};
test_output[8070] = '{32'h421ece1c};
test_index[8070] = '{2};
test_input[64568:64575] = '{32'hc291b430, 32'hc293d1d0, 32'h40b688b5, 32'hc01f59f7, 32'h42b14e34, 32'hc2b39225, 32'hc29691ac, 32'h40bb6850};
test_output[8071] = '{32'h42b14e34};
test_index[8071] = '{4};
test_input[64576:64583] = '{32'h4233bae2, 32'hc2bed349, 32'h41a79a4e, 32'h415f560f, 32'hc1f2e746, 32'hc220a92e, 32'h40e99778, 32'hc2b4bcdd};
test_output[8072] = '{32'h4233bae2};
test_index[8072] = '{0};
test_input[64584:64591] = '{32'h40b448b7, 32'h41de4eec, 32'h42b4677a, 32'h42253ae6, 32'hc104c91f, 32'h41af8acb, 32'hc15e7c4d, 32'h424771c0};
test_output[8073] = '{32'h42b4677a};
test_index[8073] = '{2};
test_input[64592:64599] = '{32'hc2053ab0, 32'h42a300fa, 32'h42057bbe, 32'h41dd5907, 32'hc2afbf45, 32'h4268480f, 32'h424192ad, 32'h3dc883ea};
test_output[8074] = '{32'h42a300fa};
test_index[8074] = '{1};
test_input[64600:64607] = '{32'hc01c05ff, 32'h42bf2a57, 32'hc103bd91, 32'hc200494b, 32'h41626081, 32'h41b785cb, 32'hc2348aaf, 32'h41551786};
test_output[8075] = '{32'h42bf2a57};
test_index[8075] = '{1};
test_input[64608:64615] = '{32'hc2ae1652, 32'h4280b4c4, 32'h3f998826, 32'hc2c4100f, 32'hc1ebf8f2, 32'hc1818b2e, 32'hc288630b, 32'hc280de1d};
test_output[8076] = '{32'h4280b4c4};
test_index[8076] = '{1};
test_input[64616:64623] = '{32'hc1b06e85, 32'h413161ae, 32'h413b3658, 32'h42997eae, 32'hc2ba0162, 32'hbfd305e9, 32'h4293bca9, 32'h4296a957};
test_output[8077] = '{32'h42997eae};
test_index[8077] = '{3};
test_input[64624:64631] = '{32'hc0efefbf, 32'hc2c049cd, 32'h4299ed5b, 32'hc1196229, 32'hc275ca38, 32'hc251d1c3, 32'h42bbaeaa, 32'hc2b137b0};
test_output[8078] = '{32'h42bbaeaa};
test_index[8078] = '{6};
test_input[64632:64639] = '{32'h42b34189, 32'h4296a83c, 32'h425f0e4f, 32'h42a24a2c, 32'hc27684cb, 32'h417ac9e7, 32'hc22a2359, 32'hc1ffcb87};
test_output[8079] = '{32'h42b34189};
test_index[8079] = '{0};
test_input[64640:64647] = '{32'hc214c49b, 32'h428f22fd, 32'hc2821a49, 32'h41c0ea48, 32'h429edbd8, 32'h4151e99a, 32'h42c5808c, 32'h426b55e1};
test_output[8080] = '{32'h42c5808c};
test_index[8080] = '{6};
test_input[64648:64655] = '{32'hc2bef90d, 32'h42c73b07, 32'h429aefeb, 32'h41b8d981, 32'h42652d61, 32'hc2b1aaaa, 32'h4228b29d, 32'h42bb6cd9};
test_output[8081] = '{32'h42c73b07};
test_index[8081] = '{1};
test_input[64656:64663] = '{32'h42227398, 32'hc2889af0, 32'hc26eb771, 32'hc2a6d0d4, 32'h425c6abd, 32'hc22b8568, 32'h4235ee1b, 32'hc0be66e9};
test_output[8082] = '{32'h425c6abd};
test_index[8082] = '{4};
test_input[64664:64671] = '{32'h42569ea1, 32'h4295a7e3, 32'h410353be, 32'h3fa5c20f, 32'hc114966d, 32'hc23baaf9, 32'hc1ab8dd8, 32'hc16cf37e};
test_output[8083] = '{32'h4295a7e3};
test_index[8083] = '{1};
test_input[64672:64679] = '{32'hc2440c5b, 32'h42259cf9, 32'hc299461b, 32'hc200170d, 32'hc281af94, 32'hc286f32d, 32'h41e29a97, 32'hc237bb45};
test_output[8084] = '{32'h42259cf9};
test_index[8084] = '{1};
test_input[64680:64687] = '{32'hc29265a1, 32'hc1844ede, 32'h41851b26, 32'h41bfac7b, 32'h42b82759, 32'h42c6eecb, 32'hc28b3369, 32'hc29618f5};
test_output[8085] = '{32'h42c6eecb};
test_index[8085] = '{5};
test_input[64688:64695] = '{32'h428242b4, 32'hc29dee62, 32'hc2a43c05, 32'h42520956, 32'hc1d964d0, 32'hc1b0a2e7, 32'hc26fd692, 32'h41abf28f};
test_output[8086] = '{32'h428242b4};
test_index[8086] = '{0};
test_input[64696:64703] = '{32'h42136e59, 32'hc296e328, 32'h42c26482, 32'h42527312, 32'h4118acc1, 32'hc2568bf6, 32'h42c1734a, 32'hc2ba225e};
test_output[8087] = '{32'h42c26482};
test_index[8087] = '{2};
test_input[64704:64711] = '{32'h42118d9a, 32'h41e35e59, 32'h42c379a1, 32'h411737d2, 32'h41e220a9, 32'h4248af31, 32'hc20c9394, 32'h42c13be6};
test_output[8088] = '{32'h42c379a1};
test_index[8088] = '{2};
test_input[64712:64719] = '{32'hc1e1f019, 32'hc19cac6c, 32'h42b5774e, 32'hc255d785, 32'h42820152, 32'hc286391d, 32'h41951da1, 32'hc1c92729};
test_output[8089] = '{32'h42b5774e};
test_index[8089] = '{2};
test_input[64720:64727] = '{32'hc284aff6, 32'h4277c7c3, 32'hc20b4755, 32'hc2456bfb, 32'hc0899394, 32'h41eec6c4, 32'h42b42f49, 32'h42aaa54d};
test_output[8090] = '{32'h42b42f49};
test_index[8090] = '{6};
test_input[64728:64735] = '{32'hc24d5ce3, 32'hc1fdbd4c, 32'h42b030d4, 32'h425824e0, 32'h429a57ce, 32'h42672cf0, 32'h428804aa, 32'h42a71bc5};
test_output[8091] = '{32'h42b030d4};
test_index[8091] = '{2};
test_input[64736:64743] = '{32'h414cdb1f, 32'hc23288a7, 32'h42282db3, 32'h40f7b0e4, 32'h40bce235, 32'h422d1815, 32'h426f6f64, 32'h41e9c7da};
test_output[8092] = '{32'h426f6f64};
test_index[8092] = '{6};
test_input[64744:64751] = '{32'h419b2217, 32'h41995fe5, 32'h41bce9ac, 32'hc2561391, 32'h423dd5d4, 32'h423a033e, 32'hc29c94fd, 32'hc2851e01};
test_output[8093] = '{32'h423dd5d4};
test_index[8093] = '{4};
test_input[64752:64759] = '{32'h427afc0c, 32'h4249b4f4, 32'hc2bd9449, 32'hc2a24d64, 32'hc1a1fddf, 32'hc21083fd, 32'hc176bed9, 32'hc2869b03};
test_output[8094] = '{32'h427afc0c};
test_index[8094] = '{0};
test_input[64760:64767] = '{32'hc2b00ae5, 32'hc1f45a93, 32'h42a659a0, 32'hc14d878f, 32'h429680b9, 32'h42535f2e, 32'hc1d810f2, 32'hc2804270};
test_output[8095] = '{32'h42a659a0};
test_index[8095] = '{2};
test_input[64768:64775] = '{32'h4145deef, 32'h41942ab9, 32'h42297dc8, 32'hc29c1890, 32'hc2b8f1d5, 32'h42076e85, 32'h42895cc4, 32'h42abab50};
test_output[8096] = '{32'h42abab50};
test_index[8096] = '{7};
test_input[64776:64783] = '{32'hc219294b, 32'hc255480e, 32'h4257857d, 32'h42a883a7, 32'h424cb8a6, 32'hc2596569, 32'hc2a8d6c8, 32'hc1c8bcd6};
test_output[8097] = '{32'h42a883a7};
test_index[8097] = '{3};
test_input[64784:64791] = '{32'hc2acf7b8, 32'hbdec8e12, 32'h414bcdbe, 32'h42b7fd1f, 32'hc2912079, 32'hc0189fb9, 32'h418f2155, 32'h41f56f33};
test_output[8098] = '{32'h42b7fd1f};
test_index[8098] = '{3};
test_input[64792:64799] = '{32'h424e984a, 32'h3fc74ec6, 32'h419d110a, 32'hc245ab7a, 32'hc2c52a8c, 32'hc285c1be, 32'h42076e13, 32'hc2bf35e1};
test_output[8099] = '{32'h424e984a};
test_index[8099] = '{0};
test_input[64800:64807] = '{32'hc15b7d23, 32'h42a287e0, 32'hc29d4a4e, 32'h42151e15, 32'h4295e1d1, 32'h40147482, 32'hc25eb2e8, 32'hc0bde36c};
test_output[8100] = '{32'h42a287e0};
test_index[8100] = '{1};
test_input[64808:64815] = '{32'h40a651ae, 32'h42912190, 32'h423763fa, 32'hc29f83ce, 32'h41f6b2ee, 32'hc2b5d263, 32'h42479e71, 32'hc241f66a};
test_output[8101] = '{32'h42912190};
test_index[8101] = '{1};
test_input[64816:64823] = '{32'hc18d6962, 32'hc0822e20, 32'h42b0bf31, 32'hc27091b8, 32'hc2723b7b, 32'hc211cd60, 32'h4225b599, 32'h4264157d};
test_output[8102] = '{32'h42b0bf31};
test_index[8102] = '{2};
test_input[64824:64831] = '{32'h42159eac, 32'h42b6c4da, 32'hc0f06c97, 32'hc2a98931, 32'h420242d0, 32'hc15b27d4, 32'h42a0ebb7, 32'h4294bc56};
test_output[8103] = '{32'h42b6c4da};
test_index[8103] = '{1};
test_input[64832:64839] = '{32'h40f675e5, 32'h42abcf9b, 32'hc28dc367, 32'h429c59fd, 32'hc2c6edfc, 32'h427e6773, 32'hc09c3cdc, 32'h42a4e3b1};
test_output[8104] = '{32'h42abcf9b};
test_index[8104] = '{1};
test_input[64840:64847] = '{32'h42495f1d, 32'h42875c79, 32'hc1b2ac2f, 32'hc188e138, 32'h42b6743f, 32'hc19c8d9b, 32'hc25bcab9, 32'hc2a4465a};
test_output[8105] = '{32'h42b6743f};
test_index[8105] = '{4};
test_input[64848:64855] = '{32'hc23b2f2a, 32'hc2471a43, 32'h4274a589, 32'h42b5b3b6, 32'hc2c7c025, 32'h4137ceff, 32'h42bbfca0, 32'hc15b53d0};
test_output[8106] = '{32'h42bbfca0};
test_index[8106] = '{6};
test_input[64856:64863] = '{32'h428401ff, 32'h42b80caa, 32'hc2c7b48f, 32'hc16b4ef4, 32'h423e26f1, 32'h426f5c49, 32'h429abd0e, 32'hc2899a2c};
test_output[8107] = '{32'h42b80caa};
test_index[8107] = '{1};
test_input[64864:64871] = '{32'hc183ad45, 32'hc2275b20, 32'h426408ef, 32'h42aa871c, 32'hc22ce952, 32'hc2907232, 32'hc25ddab1, 32'hc06146b3};
test_output[8108] = '{32'h42aa871c};
test_index[8108] = '{3};
test_input[64872:64879] = '{32'hc256ff76, 32'hc1e3cad9, 32'h41f806ec, 32'h41e57046, 32'h42a6de05, 32'h4286a281, 32'h42bb4d71, 32'hc202a02f};
test_output[8109] = '{32'h42bb4d71};
test_index[8109] = '{6};
test_input[64880:64887] = '{32'hc2776f12, 32'h41b48597, 32'h42b783d1, 32'h41c841a9, 32'hc2015786, 32'h41b75916, 32'hc2b2a909, 32'h4201c3ba};
test_output[8110] = '{32'h42b783d1};
test_index[8110] = '{2};
test_input[64888:64895] = '{32'hc10988eb, 32'h41f4735d, 32'hbfa7e10e, 32'h4211a35e, 32'hc199d88c, 32'hc206b0fa, 32'hc21976dd, 32'hc2991f0d};
test_output[8111] = '{32'h4211a35e};
test_index[8111] = '{3};
test_input[64896:64903] = '{32'h42aa33af, 32'hc29cbd6d, 32'h41c8edc7, 32'h42a8553a, 32'hc1f0bde5, 32'hc02326c4, 32'h420812ec, 32'h42c1925a};
test_output[8112] = '{32'h42c1925a};
test_index[8112] = '{7};
test_input[64904:64911] = '{32'h42b4f267, 32'h41e0145f, 32'hc2759e03, 32'h41fde4f8, 32'hc20fbddb, 32'hc2602e35, 32'hc235720d, 32'h42878f0b};
test_output[8113] = '{32'h42b4f267};
test_index[8113] = '{0};
test_input[64912:64919] = '{32'hc1020728, 32'hc28d59a9, 32'h428ef4ee, 32'hc255bb2e, 32'h428e4075, 32'hc1a38197, 32'hc224d2d9, 32'h41db6008};
test_output[8114] = '{32'h428ef4ee};
test_index[8114] = '{2};
test_input[64920:64927] = '{32'hc24d556f, 32'h40a5f465, 32'h42c60e90, 32'hc1fe3a58, 32'hc12df054, 32'hc239f8e6, 32'hc12348dc, 32'hc2a8409c};
test_output[8115] = '{32'h42c60e90};
test_index[8115] = '{2};
test_input[64928:64935] = '{32'h423c68d3, 32'h41fb1add, 32'h3fab16e3, 32'hc27647f2, 32'h422ccb45, 32'h423c98ea, 32'h412fd50d, 32'h41d6a2d9};
test_output[8116] = '{32'h423c98ea};
test_index[8116] = '{5};
test_input[64936:64943] = '{32'h3b31393d, 32'hc2ad1575, 32'h4204679f, 32'h415300ee, 32'h425b7b58, 32'h425941da, 32'h41375d5a, 32'hc24e2010};
test_output[8117] = '{32'h425b7b58};
test_index[8117] = '{4};
test_input[64944:64951] = '{32'hc28813b0, 32'hc2ad23b3, 32'hc2602308, 32'hc1ec32e3, 32'h423b2298, 32'hc233ce31, 32'hc273140b, 32'h42151712};
test_output[8118] = '{32'h423b2298};
test_index[8118] = '{4};
test_input[64952:64959] = '{32'hc2c20c0b, 32'h403f33ef, 32'hc1adfc78, 32'hc1b7a1c5, 32'h421bb22f, 32'hc219ac34, 32'h419a6ef8, 32'h42a1ff24};
test_output[8119] = '{32'h42a1ff24};
test_index[8119] = '{7};
test_input[64960:64967] = '{32'h42874626, 32'h41945eac, 32'hc296d581, 32'hc2770595, 32'hc1d4757e, 32'hc195ae19, 32'h422110d3, 32'h427c7899};
test_output[8120] = '{32'h42874626};
test_index[8120] = '{0};
test_input[64968:64975] = '{32'hc054717e, 32'hc211c570, 32'hc20263ee, 32'hc288b4f9, 32'h41ddf1d7, 32'h42403f9c, 32'h42856d7d, 32'h42ba9a0b};
test_output[8121] = '{32'h42ba9a0b};
test_index[8121] = '{7};
test_input[64976:64983] = '{32'h409a75b6, 32'h42bcaae0, 32'h42b96ee8, 32'h4275e87d, 32'hc133bea3, 32'hc288831c, 32'hc24ac40c, 32'h42b916d9};
test_output[8122] = '{32'h42bcaae0};
test_index[8122] = '{1};
test_input[64984:64991] = '{32'h42a2e0bc, 32'h41f26510, 32'hc28e13c7, 32'h40005798, 32'h4201b14d, 32'hc22995f1, 32'h40812b95, 32'hc299385a};
test_output[8123] = '{32'h42a2e0bc};
test_index[8123] = '{0};
test_input[64992:64999] = '{32'h4215009a, 32'hc1d36cfb, 32'h416b9be9, 32'h425e6de8, 32'h42a91a3f, 32'hc117f087, 32'h41f4b429, 32'h42b25f3f};
test_output[8124] = '{32'h42b25f3f};
test_index[8124] = '{7};
test_input[65000:65007] = '{32'hc2984d22, 32'hc2364872, 32'hc1eac18c, 32'hc0cef62d, 32'hc230ba2a, 32'h4296a43c, 32'h4297780f, 32'hc24fa4b7};
test_output[8125] = '{32'h4297780f};
test_index[8125] = '{6};
test_input[65008:65015] = '{32'hc0aa8cf1, 32'h4091db9f, 32'h41e039c3, 32'hc2822ce3, 32'h42c4e022, 32'h4258586d, 32'hc250410c, 32'hc2000649};
test_output[8126] = '{32'h42c4e022};
test_index[8126] = '{4};
test_input[65016:65023] = '{32'hc2a60286, 32'h42afcc8a, 32'h3f3de017, 32'h4267f66b, 32'h420e5b20, 32'hc2c32a66, 32'h3f4b82be, 32'h412ceaf7};
test_output[8127] = '{32'h42afcc8a};
test_index[8127] = '{1};
test_input[65024:65031] = '{32'hc1ee27ed, 32'h41e76bfe, 32'hc1f94b9f, 32'hc17dd7c7, 32'hc166187a, 32'hc28c669b, 32'hc2a36fc9, 32'hc290a9df};
test_output[8128] = '{32'h41e76bfe};
test_index[8128] = '{1};
test_input[65032:65039] = '{32'h41a03faa, 32'hc293caaa, 32'h424d1d76, 32'h421eac80, 32'hc2883f0b, 32'h41115aa4, 32'h42089908, 32'h429b1487};
test_output[8129] = '{32'h429b1487};
test_index[8129] = '{7};
test_input[65040:65047] = '{32'hc28619ee, 32'h4216b227, 32'h41843474, 32'hc293066f, 32'hc2c606c9, 32'hc29dfd5a, 32'hc271cab1, 32'h4296279f};
test_output[8130] = '{32'h4296279f};
test_index[8130] = '{7};
test_input[65048:65055] = '{32'h42216705, 32'h4298af3b, 32'h4224d556, 32'h42b60a0d, 32'hc27c5f84, 32'hc2965dbe, 32'hc2be045d, 32'h42936051};
test_output[8131] = '{32'h42b60a0d};
test_index[8131] = '{3};
test_input[65056:65063] = '{32'h423fc465, 32'h41f9d3d4, 32'h427f0f0f, 32'h429300cd, 32'hc28735b7, 32'h42297ee8, 32'h4295c809, 32'hc28257de};
test_output[8132] = '{32'h4295c809};
test_index[8132] = '{6};
test_input[65064:65071] = '{32'h412af734, 32'h42a2993b, 32'hc2a44989, 32'h4291a577, 32'h428cb71e, 32'hc2b094e3, 32'h42ba57aa, 32'hc1203c75};
test_output[8133] = '{32'h42ba57aa};
test_index[8133] = '{6};
test_input[65072:65079] = '{32'h4269522b, 32'hc2356728, 32'h3e0fa0e7, 32'hc0c33565, 32'hc252af01, 32'h3f0934e9, 32'h40199910, 32'hc25cd116};
test_output[8134] = '{32'h4269522b};
test_index[8134] = '{0};
test_input[65080:65087] = '{32'hc1f447b1, 32'h422ccff7, 32'hc262ce69, 32'h421a643f, 32'h40e9392b, 32'hc2a4c48e, 32'h41c60bb1, 32'hc2a8b4da};
test_output[8135] = '{32'h422ccff7};
test_index[8135] = '{1};
test_input[65088:65095] = '{32'hc22facbe, 32'hbf301f51, 32'h41aa6875, 32'hc0c64a3c, 32'h4288a068, 32'hc22b7948, 32'h42a53ba8, 32'hc26d0139};
test_output[8136] = '{32'h42a53ba8};
test_index[8136] = '{6};
test_input[65096:65103] = '{32'hc2314047, 32'hc28fdea4, 32'hc1bbe908, 32'hc1bba3da, 32'hc1124c5a, 32'hc298eceb, 32'h42a40a91, 32'hc2043e3a};
test_output[8137] = '{32'h42a40a91};
test_index[8137] = '{6};
test_input[65104:65111] = '{32'hc1ac07be, 32'hc21b63e0, 32'h40e4a98b, 32'h420700b7, 32'hc248d522, 32'hc1792a39, 32'hc28a02ad, 32'hc041c154};
test_output[8138] = '{32'h420700b7};
test_index[8138] = '{3};
test_input[65112:65119] = '{32'hc1fe58d8, 32'hc296245c, 32'h41abaa37, 32'hc243c635, 32'hc27bc5a3, 32'hc1bf03aa, 32'h42c57c24, 32'hc25fbcd8};
test_output[8139] = '{32'h42c57c24};
test_index[8139] = '{6};
test_input[65120:65127] = '{32'h42b9ec8b, 32'h41717e32, 32'hc2a78174, 32'hc2ac11b5, 32'h41ac6da7, 32'hc27410a6, 32'h4285dd30, 32'hc19d6ebe};
test_output[8140] = '{32'h42b9ec8b};
test_index[8140] = '{0};
test_input[65128:65135] = '{32'hc28b1de2, 32'hc0fa3204, 32'h4276e7cf, 32'hc24e8c02, 32'hc28b9b48, 32'hc19aa6b1, 32'hc29910da, 32'h42be849a};
test_output[8141] = '{32'h42be849a};
test_index[8141] = '{7};
test_input[65136:65143] = '{32'hbdc31a3c, 32'h420212f0, 32'h426a9655, 32'h422f1357, 32'hc1026d73, 32'h41f31d02, 32'h428f9cd7, 32'h40b2b34e};
test_output[8142] = '{32'h428f9cd7};
test_index[8142] = '{6};
test_input[65144:65151] = '{32'hc2c34eb7, 32'h42ad4e52, 32'h423d981e, 32'hc2a5cbfa, 32'h4177ef05, 32'h428b1b70, 32'hc29650f2, 32'h423e88b4};
test_output[8143] = '{32'h42ad4e52};
test_index[8143] = '{1};
test_input[65152:65159] = '{32'hbf06636f, 32'h41f7e26d, 32'h427a35cf, 32'hc2b5668c, 32'hc28030b1, 32'h42b0aa87, 32'h42b160f0, 32'h42b6b948};
test_output[8144] = '{32'h42b6b948};
test_index[8144] = '{7};
test_input[65160:65167] = '{32'h41c6c08a, 32'hc2bd9726, 32'h41c83688, 32'hc25ed56a, 32'h42906671, 32'hc20fa776, 32'hc1c14b53, 32'hc260001c};
test_output[8145] = '{32'h42906671};
test_index[8145] = '{4};
test_input[65168:65175] = '{32'hc2b1db34, 32'h42940bad, 32'h4220bc3e, 32'hc2bd84a2, 32'h429f61ae, 32'hc2c24441, 32'h42bf2930, 32'hc0729c6d};
test_output[8146] = '{32'h42bf2930};
test_index[8146] = '{6};
test_input[65176:65183] = '{32'h42bd1af6, 32'h420720f8, 32'h41b7e088, 32'h42443abf, 32'hc2a717ec, 32'hc115e17b, 32'hc1b67084, 32'hc22fd14b};
test_output[8147] = '{32'h42bd1af6};
test_index[8147] = '{0};
test_input[65184:65191] = '{32'hc2b0520e, 32'h42b6e983, 32'h413f814f, 32'hc26c6429, 32'h4287e726, 32'h42207384, 32'h425ec85e, 32'h4201984e};
test_output[8148] = '{32'h42b6e983};
test_index[8148] = '{1};
test_input[65192:65199] = '{32'hc2325294, 32'h428cca9a, 32'hc1fa463f, 32'h414fd410, 32'hc1b7dd36, 32'hc29de900, 32'hc2a6a770, 32'h42b4f587};
test_output[8149] = '{32'h42b4f587};
test_index[8149] = '{7};
test_input[65200:65207] = '{32'h41afd294, 32'hc29e113c, 32'h42b5d69b, 32'hc28546ee, 32'h4293f926, 32'hc241b777, 32'hc238b1ad, 32'h420d1efb};
test_output[8150] = '{32'h42b5d69b};
test_index[8150] = '{2};
test_input[65208:65215] = '{32'hc1a3201f, 32'h417d012d, 32'hc29a1b25, 32'hc27759f7, 32'h41f3ea02, 32'hc1716375, 32'h42a1b8e4, 32'hc0f7dbc1};
test_output[8151] = '{32'h42a1b8e4};
test_index[8151] = '{6};
test_input[65216:65223] = '{32'hc224b5d1, 32'hc27cfd29, 32'h41ae7702, 32'hc1312506, 32'h42b52b1f, 32'hc2bc461e, 32'hc2b35bdb, 32'h42823e30};
test_output[8152] = '{32'h42b52b1f};
test_index[8152] = '{4};
test_input[65224:65231] = '{32'h428a0740, 32'hc15f14c2, 32'h42940b47, 32'hc2c6e282, 32'hc1f9785e, 32'hc192e51b, 32'h428b5749, 32'h41bd3626};
test_output[8153] = '{32'h42940b47};
test_index[8153] = '{2};
test_input[65232:65239] = '{32'hc27e62c6, 32'h4292246c, 32'h4274fab9, 32'hc12b0257, 32'hc27eb24f, 32'hc27e330c, 32'hc1c52bf1, 32'h423519c1};
test_output[8154] = '{32'h4292246c};
test_index[8154] = '{1};
test_input[65240:65247] = '{32'h42099fb7, 32'h429cb9cd, 32'hc2ae4cf0, 32'h41c7ab19, 32'h42b819b8, 32'hc20e965b, 32'hc2a2eb0b, 32'hc2aa39d3};
test_output[8155] = '{32'h42b819b8};
test_index[8155] = '{4};
test_input[65248:65255] = '{32'hc2c382a3, 32'hc22450b0, 32'h4283bd4d, 32'hc2a5917b, 32'hc28b2554, 32'h41caf5e5, 32'h41922205, 32'h42b2da1f};
test_output[8156] = '{32'h42b2da1f};
test_index[8156] = '{7};
test_input[65256:65263] = '{32'h424d62ba, 32'hc154a349, 32'h424a2a47, 32'hc284e14a, 32'hc1d30eb4, 32'hc2c1223d, 32'h41be40af, 32'h41436196};
test_output[8157] = '{32'h424d62ba};
test_index[8157] = '{0};
test_input[65264:65271] = '{32'h42a1ac9d, 32'h4220600d, 32'h41282878, 32'hc2844852, 32'hc2611779, 32'h41816f83, 32'hc2bdf794, 32'h42166470};
test_output[8158] = '{32'h42a1ac9d};
test_index[8158] = '{0};
test_input[65272:65279] = '{32'h42c07b99, 32'hc2a32c30, 32'hc2b989c6, 32'h41e75ab9, 32'hc22ce849, 32'hc0e2e8e5, 32'hbf879e48, 32'h420a568f};
test_output[8159] = '{32'h42c07b99};
test_index[8159] = '{0};
test_input[65280:65287] = '{32'h428b0153, 32'hc260eadc, 32'hc20330f3, 32'h418743b5, 32'hc2b49757, 32'hc2031179, 32'h4295aebb, 32'h421e9d40};
test_output[8160] = '{32'h4295aebb};
test_index[8160] = '{6};
test_input[65288:65295] = '{32'h4270ce0b, 32'h42683c8a, 32'hc2a8eb48, 32'hc1b462c9, 32'h41236291, 32'h41d3e87e, 32'h42abf316, 32'hc14f3f1a};
test_output[8161] = '{32'h42abf316};
test_index[8161] = '{6};
test_input[65296:65303] = '{32'h426d29e0, 32'hc2c502c4, 32'h4298a19f, 32'h41e37085, 32'hc29215fa, 32'h429093bf, 32'hc1d4be97, 32'hc29c6961};
test_output[8162] = '{32'h4298a19f};
test_index[8162] = '{2};
test_input[65304:65311] = '{32'h412acc61, 32'h4246917b, 32'hc1092228, 32'hc23011a8, 32'hc2c4afff, 32'hc21da0d5, 32'h41b9eeb6, 32'h41844a14};
test_output[8163] = '{32'h4246917b};
test_index[8163] = '{1};
test_input[65312:65319] = '{32'h416f7d45, 32'h40e5094e, 32'h412cd45e, 32'hc247d73d, 32'h413888be, 32'h428fdb34, 32'hc2640fa4, 32'hc2379142};
test_output[8164] = '{32'h428fdb34};
test_index[8164] = '{5};
test_input[65320:65327] = '{32'h42912459, 32'h42361af1, 32'hc07446fc, 32'hc24cd9ad, 32'hc2c5af15, 32'hc27aa640, 32'hc180c8d2, 32'hc2a3ee09};
test_output[8165] = '{32'h42912459};
test_index[8165] = '{0};
test_input[65328:65335] = '{32'hc20e6ac0, 32'h42b662a0, 32'h42b618c2, 32'h42c59f26, 32'hc082fb5c, 32'h409b7025, 32'hc258a656, 32'h42892071};
test_output[8166] = '{32'h42c59f26};
test_index[8166] = '{3};
test_input[65336:65343] = '{32'h4284b9e4, 32'hc2c10788, 32'hc28dacd5, 32'hc234c1ab, 32'hc2bcd5c1, 32'hc2ac9f92, 32'h41a6b6fe, 32'hc27e5c89};
test_output[8167] = '{32'h4284b9e4};
test_index[8167] = '{0};
test_input[65344:65351] = '{32'h41bedaec, 32'h4053cd05, 32'h41d1d0b9, 32'h42018767, 32'h42c751d8, 32'hc13111e7, 32'hc2a86342, 32'hc2c6ea49};
test_output[8168] = '{32'h42c751d8};
test_index[8168] = '{4};
test_input[65352:65359] = '{32'hc10aa4e7, 32'h41b72ad0, 32'h42c402f6, 32'hc25505d2, 32'hc0eb0e73, 32'hbe7dae1a, 32'h4297d6cb, 32'hc2483118};
test_output[8169] = '{32'h42c402f6};
test_index[8169] = '{2};
test_input[65360:65367] = '{32'hc2b4256b, 32'h410f52d0, 32'hc22ca4bd, 32'hc19b03cb, 32'hc0c48b8e, 32'hc2ad3383, 32'hc2bc028c, 32'h41efb1c6};
test_output[8170] = '{32'h41efb1c6};
test_index[8170] = '{7};
test_input[65368:65375] = '{32'hc296a4c2, 32'hc2b3125e, 32'hc1f6dbb0, 32'hc2291b22, 32'h42bbd95b, 32'hc2922393, 32'hc2b9ea01, 32'hc1e26de4};
test_output[8171] = '{32'h42bbd95b};
test_index[8171] = '{4};
test_input[65376:65383] = '{32'hc29b0cf4, 32'h42b8b236, 32'h41c09730, 32'h42611ffd, 32'h40bf1758, 32'h42287f7d, 32'h42bdfcfa, 32'h428dfb2f};
test_output[8172] = '{32'h42bdfcfa};
test_index[8172] = '{6};
test_input[65384:65391] = '{32'hc262a5cb, 32'h40fb0187, 32'hc2c33e0c, 32'hc213a22e, 32'h40b04622, 32'hc291adc4, 32'hc2b2511d, 32'hc281c9db};
test_output[8173] = '{32'h40fb0187};
test_index[8173] = '{1};
test_input[65392:65399] = '{32'h418a59bc, 32'h40fc36df, 32'h421319dd, 32'h4297ddd1, 32'h41623b31, 32'hc2baffb4, 32'h427a7e8d, 32'hbe5961b6};
test_output[8174] = '{32'h4297ddd1};
test_index[8174] = '{3};
test_input[65400:65407] = '{32'hc292e34f, 32'hc215f8c3, 32'h4242de73, 32'h41944d3c, 32'h40aa9500, 32'h421ee3e4, 32'h422b541d, 32'hc2bbaa8a};
test_output[8175] = '{32'h4242de73};
test_index[8175] = '{2};
test_input[65408:65415] = '{32'h4298b4fe, 32'hc1cb48ba, 32'hc28d8a75, 32'h42a18ac2, 32'h42c27b61, 32'h42792147, 32'h41e5309f, 32'hc2bfaaf4};
test_output[8176] = '{32'h42c27b61};
test_index[8176] = '{4};
test_input[65416:65423] = '{32'h4286af84, 32'hc28eb79c, 32'hc2ad38a7, 32'hc24ebbd8, 32'hc29bf914, 32'hc1eb51e7, 32'hc2685d2b, 32'h4243f876};
test_output[8177] = '{32'h4286af84};
test_index[8177] = '{0};
test_input[65424:65431] = '{32'hc2bdd9c4, 32'hc2558ad8, 32'h410154e6, 32'h42b31894, 32'h4291b232, 32'h41039b29, 32'h42a175f4, 32'h429bb792};
test_output[8178] = '{32'h42b31894};
test_index[8178] = '{3};
test_input[65432:65439] = '{32'h42554924, 32'h42297c3d, 32'hc20bf6ef, 32'hc2b4626c, 32'hc22c434f, 32'h406c0b76, 32'h428844b7, 32'h412620f6};
test_output[8179] = '{32'h428844b7};
test_index[8179] = '{6};
test_input[65440:65447] = '{32'h42aa9469, 32'h4088dea8, 32'h429c40fc, 32'hc277797c, 32'hc14c6e2b, 32'hc2c3b11b, 32'h4293b694, 32'hc28f19b9};
test_output[8180] = '{32'h42aa9469};
test_index[8180] = '{0};
test_input[65448:65455] = '{32'hc2bdb666, 32'h4244a0b5, 32'hc2bcec81, 32'hbe40dcb4, 32'hc2afa3af, 32'h42559726, 32'hc0f0e80d, 32'hc294bd43};
test_output[8181] = '{32'h42559726};
test_index[8181] = '{5};
test_input[65456:65463] = '{32'hc2b0e6f7, 32'h42bdd7f2, 32'h423410bc, 32'hc133956d, 32'h41b0277a, 32'hc22d7252, 32'hc23a8b79, 32'h41ccc42f};
test_output[8182] = '{32'h42bdd7f2};
test_index[8182] = '{1};
test_input[65464:65471] = '{32'hc0fb17e1, 32'h422ae094, 32'hc15ed0b6, 32'h40e9199f, 32'h429653c9, 32'h41b78ab5, 32'h42a8e554, 32'hc230b7d4};
test_output[8183] = '{32'h42a8e554};
test_index[8183] = '{6};
test_input[65472:65479] = '{32'h41ea5197, 32'hc1a8c85b, 32'h417e4f8e, 32'h418b0c0a, 32'h429a6548, 32'hc235e39d, 32'h426f1892, 32'hc29d33f6};
test_output[8184] = '{32'h429a6548};
test_index[8184] = '{4};
test_input[65480:65487] = '{32'h407cf894, 32'h423cfed2, 32'hc21ea055, 32'hc1630695, 32'h421a6a7a, 32'hc29c57d7, 32'hc292b5d4, 32'h4238d223};
test_output[8185] = '{32'h423cfed2};
test_index[8185] = '{1};
test_input[65488:65495] = '{32'hc1ad592e, 32'hc2afab2b, 32'h4204a98e, 32'hc0fe9b97, 32'h422c4675, 32'hc2bf087c, 32'hc0b793b2, 32'h42a06bc3};
test_output[8186] = '{32'h42a06bc3};
test_index[8186] = '{7};
test_input[65496:65503] = '{32'h42b8f5bc, 32'h41eb03a6, 32'hc263661f, 32'h426d90bb, 32'h422dcd15, 32'h42ad5cc7, 32'h42175aea, 32'hc0c2f2cb};
test_output[8187] = '{32'h42b8f5bc};
test_index[8187] = '{0};
test_input[65504:65511] = '{32'h42288573, 32'h4202b00b, 32'h41cfff85, 32'hc28fe145, 32'h429d22bc, 32'h41018f4e, 32'hc200230f, 32'hc2685f82};
test_output[8188] = '{32'h429d22bc};
test_index[8188] = '{4};
test_input[65512:65519] = '{32'hc28fc5c8, 32'h42bec10b, 32'h42b8f284, 32'h42024cf1, 32'hc2875e52, 32'hc29ca704, 32'hc283eda4, 32'hc26bb8ad};
test_output[8189] = '{32'h42bec10b};
test_index[8189] = '{1};
test_input[65520:65527] = '{32'hc27d3f15, 32'h41644e8b, 32'hc28f1622, 32'h42b600c7, 32'hc21c81ab, 32'h429847a5, 32'hc26e0bf7, 32'hc1d54442};
test_output[8190] = '{32'h42b600c7};
test_index[8190] = '{3};
test_input[65528:65535] = '{32'hc26ac363, 32'h419124e8, 32'h42a8bc8f, 32'hc23f7d79, 32'hc1ba7735, 32'h3ed7aaff, 32'h427b953b, 32'h41947e71};
test_output[8191] = '{32'h42a8bc8f};
test_index[8191] = '{2};
test_input[65536:65543] = '{32'hc23eeb66, 32'hc2320110, 32'h3f6d9602, 32'h425f3280, 32'hc2967759, 32'hc2173091, 32'h4295aaa0, 32'h4222435c};
test_output[8192] = '{32'h4295aaa0};
test_index[8192] = '{6};
test_input[65544:65551] = '{32'hc27a8001, 32'h42448f65, 32'h4299281d, 32'hc290a8c9, 32'h42c19ed8, 32'hc28ae274, 32'h4123c9f7, 32'hc0da8b71};
test_output[8193] = '{32'h42c19ed8};
test_index[8193] = '{4};
test_input[65552:65559] = '{32'hc29672c1, 32'h41f2121c, 32'h4263f749, 32'hc2c6afd0, 32'h42320758, 32'hc29bf231, 32'hc233d9c5, 32'h4299db04};
test_output[8194] = '{32'h4299db04};
test_index[8194] = '{7};
test_input[65560:65567] = '{32'h40c6d6d3, 32'hc26fd21e, 32'hc232c2b8, 32'h423671fa, 32'h429db7dc, 32'h4231bc54, 32'hc2263ad1, 32'hc29656ef};
test_output[8195] = '{32'h429db7dc};
test_index[8195] = '{4};
test_input[65568:65575] = '{32'h40f05ac2, 32'h4185ab41, 32'hc2885e36, 32'hc1a7d4ea, 32'hc2b1e49d, 32'h4222f25d, 32'h42bae318, 32'hc2a0675d};
test_output[8196] = '{32'h42bae318};
test_index[8196] = '{6};
test_input[65576:65583] = '{32'h42305cac, 32'h42b4af92, 32'h42c7ef62, 32'h429deb0b, 32'h423b2987, 32'hc234652d, 32'h41b31197, 32'h4230946d};
test_output[8197] = '{32'h42c7ef62};
test_index[8197] = '{2};
test_input[65584:65591] = '{32'hc2aedd89, 32'hc1d24984, 32'h411b6b8d, 32'h42a42db0, 32'h41d77146, 32'h42506565, 32'h42a1b3a8, 32'h426ea13b};
test_output[8198] = '{32'h42a42db0};
test_index[8198] = '{3};
test_input[65592:65599] = '{32'hc1e9ec8e, 32'hc25254bd, 32'h4274dc87, 32'hc2830393, 32'hc23b126b, 32'hc20cd1aa, 32'hc2a4000c, 32'hc24c01ef};
test_output[8199] = '{32'h4274dc87};
test_index[8199] = '{2};
test_input[65600:65607] = '{32'h4281eba8, 32'hc2216c02, 32'h42b82164, 32'h429a4c88, 32'h412243cc, 32'hc1badfa9, 32'h3fbecd75, 32'h41ad8563};
test_output[8200] = '{32'h42b82164};
test_index[8200] = '{2};
test_input[65608:65615] = '{32'hc2703da4, 32'h4071496c, 32'hc2b93c33, 32'h3f342e78, 32'hc1b72267, 32'hc19cc97d, 32'hc291a95f, 32'h429ba5be};
test_output[8201] = '{32'h429ba5be};
test_index[8201] = '{7};
test_input[65616:65623] = '{32'h41cb2651, 32'hc231eda9, 32'h4287e6b3, 32'h42b7f01f, 32'hc2adde84, 32'h42ba72a9, 32'hc2aca1ca, 32'h41638403};
test_output[8202] = '{32'h42ba72a9};
test_index[8202] = '{5};
test_input[65624:65631] = '{32'hc216853d, 32'h40636da0, 32'hc27755c0, 32'hc26ae0b7, 32'h429dff8e, 32'hc234dd17, 32'hc132eb39, 32'hc15df833};
test_output[8203] = '{32'h429dff8e};
test_index[8203] = '{4};
test_input[65632:65639] = '{32'h428402c4, 32'h42179852, 32'hc1f75072, 32'h42486a83, 32'h423dd2b8, 32'hc214d9f5, 32'hc2c2494a, 32'h42c50d77};
test_output[8204] = '{32'h42c50d77};
test_index[8204] = '{7};
test_input[65640:65647] = '{32'h42a838e1, 32'hc28cfc9b, 32'hc2c5db56, 32'h41a6546f, 32'hc27a0be8, 32'h421a559e, 32'h4259a1bc, 32'hc20febe6};
test_output[8205] = '{32'h42a838e1};
test_index[8205] = '{0};
test_input[65648:65655] = '{32'hc24d49e3, 32'h4226eeec, 32'hc2578f81, 32'h42acc9a5, 32'h414454e1, 32'h426461d4, 32'hc2b264e4, 32'h42b812a3};
test_output[8206] = '{32'h42b812a3};
test_index[8206] = '{7};
test_input[65656:65663] = '{32'hc265ae50, 32'h418add72, 32'h41e5989b, 32'hc267699e, 32'h42362384, 32'h41835589, 32'h42af41f0, 32'h4259c138};
test_output[8207] = '{32'h42af41f0};
test_index[8207] = '{6};
test_input[65664:65671] = '{32'h421b8988, 32'h42073609, 32'hc2241b0d, 32'hc24e3a8a, 32'h42c67b3f, 32'h42c0d846, 32'h41cc8e1c, 32'h4295f701};
test_output[8208] = '{32'h42c67b3f};
test_index[8208] = '{4};
test_input[65672:65679] = '{32'h425c1fea, 32'hc1faa759, 32'h429225c3, 32'h41f34202, 32'hc2662a86, 32'hc2c4e9b9, 32'h42303174, 32'h42527fe9};
test_output[8209] = '{32'h429225c3};
test_index[8209] = '{2};
test_input[65680:65687] = '{32'hc2701be1, 32'hc1a9ce02, 32'hc1dd1cd0, 32'hc29965d2, 32'h429b3763, 32'hc1aeb4de, 32'hbdb978fd, 32'hc2bedbee};
test_output[8210] = '{32'h429b3763};
test_index[8210] = '{4};
test_input[65688:65695] = '{32'h4200a546, 32'hc2672424, 32'hc2ac10e1, 32'h41a0f893, 32'hc2b8710b, 32'hc1ba8929, 32'hc2bae677, 32'h4208dae5};
test_output[8211] = '{32'h4208dae5};
test_index[8211] = '{7};
test_input[65696:65703] = '{32'hc28b2a4e, 32'h41f23994, 32'h41a95a71, 32'h41431803, 32'h4002a613, 32'h429a3b40, 32'h422ba82d, 32'hc18bcdff};
test_output[8212] = '{32'h429a3b40};
test_index[8212] = '{5};
test_input[65704:65711] = '{32'hc271775c, 32'hc241fffa, 32'hc21020f7, 32'h42c5c66f, 32'h42658d23, 32'hc2be244e, 32'h4277f9e7, 32'hc1aa0438};
test_output[8213] = '{32'h42c5c66f};
test_index[8213] = '{3};
test_input[65712:65719] = '{32'hc2b1ecd2, 32'h42a2ee88, 32'hc2c0eb58, 32'hc2baf8cc, 32'h429edfb4, 32'h410e88ff, 32'h42a31426, 32'h420c90d0};
test_output[8214] = '{32'h42a31426};
test_index[8214] = '{6};
test_input[65720:65727] = '{32'hc23281fe, 32'h42c635eb, 32'h4154392c, 32'hc1c65cfc, 32'hc1ac1079, 32'hc246aafe, 32'hc283593a, 32'h41cb307f};
test_output[8215] = '{32'h42c635eb};
test_index[8215] = '{1};
test_input[65728:65735] = '{32'h41a40993, 32'h429af87d, 32'hc294407f, 32'h41c73aea, 32'hc29918d6, 32'h40badf39, 32'hc21105b4, 32'h416d1815};
test_output[8216] = '{32'h429af87d};
test_index[8216] = '{1};
test_input[65736:65743] = '{32'h418b2f5e, 32'h41ebb0e8, 32'hc21806de, 32'h4283884f, 32'hc26c0be3, 32'h40d95474, 32'hc2927ef9, 32'hc25663ff};
test_output[8217] = '{32'h4283884f};
test_index[8217] = '{3};
test_input[65744:65751] = '{32'hc293fc22, 32'hc055b8c3, 32'h42a47eac, 32'hc292adaf, 32'h418b949a, 32'h42b90e53, 32'hc2c53d28, 32'hc1e2b3f1};
test_output[8218] = '{32'h42b90e53};
test_index[8218] = '{5};
test_input[65752:65759] = '{32'h429e79c6, 32'hc0517f31, 32'hc2aa1ca0, 32'h42bbec27, 32'h4207ea05, 32'h42933a3b, 32'hc2a2fe51, 32'hc1ed51b2};
test_output[8219] = '{32'h42bbec27};
test_index[8219] = '{3};
test_input[65760:65767] = '{32'hbf0c302a, 32'h4247d4e3, 32'hc2bc2804, 32'hc1656648, 32'hc1b86483, 32'hc261026a, 32'h42a7c0d7, 32'h413346cc};
test_output[8220] = '{32'h42a7c0d7};
test_index[8220] = '{6};
test_input[65768:65775] = '{32'h42ad87ab, 32'h420a24a1, 32'hc290d933, 32'hc118b9fe, 32'h4283f33d, 32'hc1c28642, 32'hc22f6fd4, 32'h4069df53};
test_output[8221] = '{32'h42ad87ab};
test_index[8221] = '{0};
test_input[65776:65783] = '{32'hc28224dd, 32'hc29437fc, 32'hc0f95b1b, 32'h428520d8, 32'h4228df6d, 32'hc214e006, 32'h421fd642, 32'hbfffd8b1};
test_output[8222] = '{32'h428520d8};
test_index[8222] = '{3};
test_input[65784:65791] = '{32'h42679175, 32'h429af832, 32'h42c37a2f, 32'h4247406c, 32'hbf82c1c0, 32'hc2a04a3d, 32'h41f0ffcf, 32'hc0094682};
test_output[8223] = '{32'h42c37a2f};
test_index[8223] = '{2};
test_input[65792:65799] = '{32'hc29b3a25, 32'hc294351d, 32'hc0a439ff, 32'hc29bfb1f, 32'h42911264, 32'hc265c833, 32'hc27c55b4, 32'hc18a58d6};
test_output[8224] = '{32'h42911264};
test_index[8224] = '{4};
test_input[65800:65807] = '{32'hc24ee402, 32'hc111d1fb, 32'hc2b2dfde, 32'hbf907265, 32'hc26b596d, 32'hc2c1fb0e, 32'hc2ba45f3, 32'h3fc20268};
test_output[8225] = '{32'h3fc20268};
test_index[8225] = '{7};
test_input[65808:65815] = '{32'hc1087586, 32'h42814548, 32'h41c24527, 32'h40e4df2f, 32'hc2127c5c, 32'hc2a80482, 32'hc25a4b10, 32'h42b1b5a6};
test_output[8226] = '{32'h42b1b5a6};
test_index[8226] = '{7};
test_input[65816:65823] = '{32'h42bb9b0d, 32'h42642378, 32'h42b2eacd, 32'hc234e9ca, 32'hc11f1604, 32'hc21a72a2, 32'hc1b36bfe, 32'h42a986ee};
test_output[8227] = '{32'h42bb9b0d};
test_index[8227] = '{0};
test_input[65824:65831] = '{32'hbf4125d1, 32'hbff76361, 32'hc24bd829, 32'hc2131ad4, 32'hc26932c0, 32'hc2ab55cf, 32'h428949a2, 32'hc18a3ca2};
test_output[8228] = '{32'h428949a2};
test_index[8228] = '{6};
test_input[65832:65839] = '{32'h42893fdd, 32'hc2159bc8, 32'h40a5f146, 32'hc1cb581c, 32'hc2b3260f, 32'hc17e756a, 32'hc2bad50c, 32'hc1d2a264};
test_output[8229] = '{32'h42893fdd};
test_index[8229] = '{0};
test_input[65840:65847] = '{32'h420caadb, 32'hc1b6b96a, 32'h4295efca, 32'h427cb583, 32'h423c5a6b, 32'hc255ea33, 32'h423d1ab7, 32'hc28cb008};
test_output[8230] = '{32'h4295efca};
test_index[8230] = '{2};
test_input[65848:65855] = '{32'hc1f5b10d, 32'h42bfec63, 32'h42c70703, 32'h424b2328, 32'hc29a066d, 32'hc23f332e, 32'h42ada2b9, 32'h421524d3};
test_output[8231] = '{32'h42c70703};
test_index[8231] = '{2};
test_input[65856:65863] = '{32'hc21a85c8, 32'h429073a6, 32'h403ae18b, 32'h4255bdd2, 32'h42a1b672, 32'hc214abb6, 32'hc0d1ee78, 32'h42c3e67e};
test_output[8232] = '{32'h42c3e67e};
test_index[8232] = '{7};
test_input[65864:65871] = '{32'hc260b2e8, 32'hc297f76e, 32'h42390804, 32'hc2045879, 32'h4230cdbb, 32'h42b527f6, 32'h423c33de, 32'hc1867a47};
test_output[8233] = '{32'h42b527f6};
test_index[8233] = '{5};
test_input[65872:65879] = '{32'hc226147f, 32'h42943628, 32'h4236726f, 32'hc2b4883e, 32'hc008390f, 32'h42468474, 32'h4163eee7, 32'hc1af7c05};
test_output[8234] = '{32'h42943628};
test_index[8234] = '{1};
test_input[65880:65887] = '{32'h41e3569d, 32'h42a0c847, 32'h42712f32, 32'h4254fdb3, 32'h42c2cedb, 32'h41b71a9f, 32'h42392c45, 32'h41cb4531};
test_output[8235] = '{32'h42c2cedb};
test_index[8235] = '{4};
test_input[65888:65895] = '{32'hc22bb952, 32'h42771841, 32'hc20230f0, 32'h42ae6e08, 32'hc27f11ec, 32'h427ae320, 32'hc22605a5, 32'h41917036};
test_output[8236] = '{32'h42ae6e08};
test_index[8236] = '{3};
test_input[65896:65903] = '{32'h41768036, 32'h41a5cc83, 32'hc1343e8f, 32'h42be49c5, 32'h422069f0, 32'hc285130a, 32'h4221ae9e, 32'hc2abb6bd};
test_output[8237] = '{32'h42be49c5};
test_index[8237] = '{3};
test_input[65904:65911] = '{32'hc25bf33a, 32'hc26ecf3d, 32'hc2ad20a7, 32'h427335ce, 32'h42a2c082, 32'hc18cdaf4, 32'h41871f17, 32'h40d198b1};
test_output[8238] = '{32'h42a2c082};
test_index[8238] = '{4};
test_input[65912:65919] = '{32'h42c669e4, 32'hc2c77ca5, 32'h42bcd022, 32'h42317c54, 32'h42872339, 32'h41a1f1db, 32'h422b815c, 32'h423cf777};
test_output[8239] = '{32'h42c669e4};
test_index[8239] = '{0};
test_input[65920:65927] = '{32'hc225ac6f, 32'hbfcad04c, 32'h42690784, 32'h428fcb09, 32'h41cea0d2, 32'h416a8fee, 32'hc21c535d, 32'h41e4d110};
test_output[8240] = '{32'h428fcb09};
test_index[8240] = '{3};
test_input[65928:65935] = '{32'hc28b8e84, 32'hc1ffaec4, 32'hc26df902, 32'h42998080, 32'hc2821e6e, 32'hc273f7f0, 32'hc28669d3, 32'h42b9f679};
test_output[8241] = '{32'h42b9f679};
test_index[8241] = '{7};
test_input[65936:65943] = '{32'hc2248303, 32'hc2983eb2, 32'hc1c7db73, 32'hc2aaef53, 32'h41ca564e, 32'hc2178efe, 32'hc0849dc2, 32'hc1e813d0};
test_output[8242] = '{32'h41ca564e};
test_index[8242] = '{4};
test_input[65944:65951] = '{32'hc29b1f14, 32'hc2a5aa96, 32'h42601f11, 32'hc205871c, 32'hc2b49d14, 32'h42b0c4b5, 32'h428b3cb9, 32'h42bf9eb7};
test_output[8243] = '{32'h42bf9eb7};
test_index[8243] = '{7};
test_input[65952:65959] = '{32'h41ff8940, 32'hc297cbd3, 32'hc0bd58f6, 32'hc2610985, 32'hc27fa49f, 32'h419f0a32, 32'h4014cab2, 32'hc174da50};
test_output[8244] = '{32'h41ff8940};
test_index[8244] = '{0};
test_input[65960:65967] = '{32'hc1ab61c7, 32'h41e84536, 32'hc10d53c5, 32'h4296448d, 32'hc1a5210d, 32'h42a62e70, 32'h42b7575a, 32'hc1492ad6};
test_output[8245] = '{32'h42b7575a};
test_index[8245] = '{6};
test_input[65968:65975] = '{32'hc1af64d9, 32'hc28962a4, 32'hc29c84f8, 32'hc294dffe, 32'hc2adba2c, 32'h4206108b, 32'h42b3f451, 32'h42a0c902};
test_output[8246] = '{32'h42b3f451};
test_index[8246] = '{6};
test_input[65976:65983] = '{32'hc255c103, 32'hc2534f47, 32'h42565b18, 32'h42035a4e, 32'hc2afc92a, 32'hc19ebca7, 32'h42759af8, 32'h422c6c4d};
test_output[8247] = '{32'h42759af8};
test_index[8247] = '{6};
test_input[65984:65991] = '{32'hc29ffaec, 32'h41791f24, 32'hc2ad2ba2, 32'h422a6b1b, 32'hc29a607a, 32'hbef4f73e, 32'h41f324a6, 32'hc0983a74};
test_output[8248] = '{32'h422a6b1b};
test_index[8248] = '{3};
test_input[65992:65999] = '{32'h426a2920, 32'h410c2d84, 32'h42857a9c, 32'hc2b7d71e, 32'h4183b0e8, 32'hc28572fb, 32'hc28fb768, 32'hc02772af};
test_output[8249] = '{32'h42857a9c};
test_index[8249] = '{2};
test_input[66000:66007] = '{32'hc267b9fd, 32'h41e554d7, 32'h418cd344, 32'hc2ac0068, 32'hc2088085, 32'h41680c86, 32'h42a1a7f7, 32'hc259dbf9};
test_output[8250] = '{32'h42a1a7f7};
test_index[8250] = '{6};
test_input[66008:66015] = '{32'h4268dafb, 32'hc21bf6cb, 32'hc20e6c73, 32'h41308a9b, 32'hc28f0b96, 32'hc22b354a, 32'h42c7c545, 32'h41674384};
test_output[8251] = '{32'h42c7c545};
test_index[8251] = '{6};
test_input[66016:66023] = '{32'hc18ead92, 32'hc2c28a98, 32'h421bef33, 32'hc260e39b, 32'h4167e392, 32'h41ad747b, 32'h421e4440, 32'h41ae51d8};
test_output[8252] = '{32'h421e4440};
test_index[8252] = '{6};
test_input[66024:66031] = '{32'hc268178a, 32'h4297a86b, 32'h41a0b5a5, 32'hc24170aa, 32'hc2401397, 32'h42a651cb, 32'hc1b0a3b2, 32'hc286a24d};
test_output[8253] = '{32'h42a651cb};
test_index[8253] = '{5};
test_input[66032:66039] = '{32'h424759eb, 32'h4166035b, 32'hc03082b8, 32'h41f10320, 32'hc1d10142, 32'h42af7f49, 32'h422a32bf, 32'h416ed027};
test_output[8254] = '{32'h42af7f49};
test_index[8254] = '{5};
test_input[66040:66047] = '{32'hc288254b, 32'hc256543a, 32'hc2542783, 32'hc2622825, 32'h42431b2b, 32'h41e96dca, 32'h421f0355, 32'h40162213};
test_output[8255] = '{32'h42431b2b};
test_index[8255] = '{4};
test_input[66048:66055] = '{32'hc271f529, 32'hc2a46c69, 32'hc1c378e6, 32'h4181aedb, 32'h4184850e, 32'hc12ef416, 32'h425d5d24, 32'hc18c29a2};
test_output[8256] = '{32'h425d5d24};
test_index[8256] = '{6};
test_input[66056:66063] = '{32'hc281bd54, 32'h4207a9a5, 32'h4289f3a4, 32'hc14377f6, 32'h41487701, 32'hc0c24389, 32'hc2b707db, 32'h422b6f0e};
test_output[8257] = '{32'h4289f3a4};
test_index[8257] = '{2};
test_input[66064:66071] = '{32'hc28bb664, 32'h428e52b5, 32'hc22a018e, 32'h42460658, 32'h41a00bed, 32'hc1e3922c, 32'h42ab06c8, 32'h40c85a7c};
test_output[8258] = '{32'h42ab06c8};
test_index[8258] = '{6};
test_input[66072:66079] = '{32'h4209586d, 32'h42b5f9ba, 32'hc129f25e, 32'hc2777e06, 32'hc120dc27, 32'hc2aec72a, 32'hc2770c77, 32'hc20fd290};
test_output[8259] = '{32'h42b5f9ba};
test_index[8259] = '{1};
test_input[66080:66087] = '{32'hc21d32aa, 32'hc2920f1c, 32'h42323139, 32'hc2a73f7b, 32'h41dc89bf, 32'hc12df058, 32'h429128d7, 32'h429cb511};
test_output[8260] = '{32'h429cb511};
test_index[8260] = '{7};
test_input[66088:66095] = '{32'hc12a5aef, 32'h41ae2bf0, 32'hc29adc1a, 32'h42c2f985, 32'h417ee38e, 32'h42c688d9, 32'h42c4cfb0, 32'h425ee93d};
test_output[8261] = '{32'h42c688d9};
test_index[8261] = '{5};
test_input[66096:66103] = '{32'hc2b8a1f0, 32'h41599e51, 32'h42a33013, 32'h4295505c, 32'h4295b57d, 32'h41da9f1d, 32'hc2045276, 32'h42a4be24};
test_output[8262] = '{32'h42a4be24};
test_index[8262] = '{7};
test_input[66104:66111] = '{32'h42bb661f, 32'hc2055390, 32'hc2022e88, 32'h424fe661, 32'h419ceb96, 32'h42ac8f60, 32'h41fecc45, 32'h429cdc2d};
test_output[8263] = '{32'h42bb661f};
test_index[8263] = '{0};
test_input[66112:66119] = '{32'hc26ffc84, 32'hbffbb5dd, 32'hc266408b, 32'h42bdc0da, 32'hc2bdf10d, 32'hc2917076, 32'hc28d5371, 32'h42b03a0a};
test_output[8264] = '{32'h42bdc0da};
test_index[8264] = '{3};
test_input[66120:66127] = '{32'hc288483d, 32'hc26f128d, 32'hc2a87b9e, 32'hc2179d1b, 32'hc1aea50e, 32'hc1ad43b8, 32'h4134d1ac, 32'hc153a8ce};
test_output[8265] = '{32'h4134d1ac};
test_index[8265] = '{6};
test_input[66128:66135] = '{32'h422f211e, 32'h41f585b6, 32'hc2863306, 32'h402be229, 32'h412be6bd, 32'h42b9e564, 32'hc246f867, 32'hc1aef70e};
test_output[8266] = '{32'h42b9e564};
test_index[8266] = '{5};
test_input[66136:66143] = '{32'hc221a5fb, 32'h42936d40, 32'hc0a5bf69, 32'h41e1a7ca, 32'h42987c39, 32'hc1df33fd, 32'hc290dcdc, 32'h42300d7c};
test_output[8267] = '{32'h42987c39};
test_index[8267] = '{4};
test_input[66144:66151] = '{32'hbfe9be0d, 32'h42560aaa, 32'hc2bf4842, 32'hc1c2fa7a, 32'hc298dcff, 32'hc1375e19, 32'hc1d7417c, 32'hc1cd6851};
test_output[8268] = '{32'h42560aaa};
test_index[8268] = '{1};
test_input[66152:66159] = '{32'hc2471e74, 32'h4171ec24, 32'h401987d3, 32'hc14f8699, 32'hc20c577c, 32'hc2b0dddb, 32'h423a0f6e, 32'h419402a3};
test_output[8269] = '{32'h423a0f6e};
test_index[8269] = '{6};
test_input[66160:66167] = '{32'h4221d509, 32'h42ae2743, 32'h4161bb64, 32'hc2aa4165, 32'h4112c642, 32'hc2230194, 32'hc29668da, 32'h4285d48a};
test_output[8270] = '{32'h42ae2743};
test_index[8270] = '{1};
test_input[66168:66175] = '{32'h42a43c87, 32'hc2bf4909, 32'hc0d7dcfc, 32'hc26449d5, 32'hc2a0d446, 32'hc2ada413, 32'h428b1031, 32'h41b0f181};
test_output[8271] = '{32'h42a43c87};
test_index[8271] = '{0};
test_input[66176:66183] = '{32'hc2abf7b7, 32'hc272d2fc, 32'h42b2d568, 32'h400fc1ce, 32'hc24f8fed, 32'h426af176, 32'h415cde8d, 32'hc28dfa2a};
test_output[8272] = '{32'h42b2d568};
test_index[8272] = '{2};
test_input[66184:66191] = '{32'hc0b1c1d6, 32'h41f9f374, 32'hc2c316f3, 32'hc2b138b4, 32'hc29e241d, 32'hc0fb04de, 32'hc17f2a89, 32'hc233b79f};
test_output[8273] = '{32'h41f9f374};
test_index[8273] = '{1};
test_input[66192:66199] = '{32'h42482bac, 32'h41b5071f, 32'h4253e294, 32'h4299cc2c, 32'hc2ab8fec, 32'h42b66250, 32'hc256c98c, 32'h40f5bcab};
test_output[8274] = '{32'h42b66250};
test_index[8274] = '{5};
test_input[66200:66207] = '{32'hc2943bf7, 32'hc11e80cb, 32'hc094c154, 32'hc28f5f55, 32'h429a6f01, 32'hc25cec01, 32'hc2a06b73, 32'hc1be5cce};
test_output[8275] = '{32'h429a6f01};
test_index[8275] = '{4};
test_input[66208:66215] = '{32'hc097da88, 32'hc2582711, 32'h41370518, 32'h402e08a0, 32'hc2043c08, 32'h42663b78, 32'h41695416, 32'h4291d679};
test_output[8276] = '{32'h4291d679};
test_index[8276] = '{7};
test_input[66216:66223] = '{32'hc270fcf0, 32'h426c2e37, 32'hc17d64bf, 32'hc23d9640, 32'h42a857db, 32'hc2261358, 32'h4114ea7a, 32'h428139b1};
test_output[8277] = '{32'h42a857db};
test_index[8277] = '{4};
test_input[66224:66231] = '{32'hc20e92c4, 32'h41f54942, 32'hc2bd9c05, 32'h42ab4f3a, 32'h422ec637, 32'h414843c4, 32'h41dd372b, 32'hc1154474};
test_output[8278] = '{32'h42ab4f3a};
test_index[8278] = '{3};
test_input[66232:66239] = '{32'hc2612a78, 32'h42c44a4f, 32'h41006750, 32'hc224fd68, 32'hc20b366b, 32'h42082048, 32'h41ae3e5e, 32'hc2b139f5};
test_output[8279] = '{32'h42c44a4f};
test_index[8279] = '{1};
test_input[66240:66247] = '{32'h424da7d9, 32'hc20b0faa, 32'hc15f1f0f, 32'hc17af869, 32'h42aaa045, 32'hc1ff73ba, 32'h4280a475, 32'h41ff3ef6};
test_output[8280] = '{32'h42aaa045};
test_index[8280] = '{4};
test_input[66248:66255] = '{32'hc2a4a914, 32'hc292258b, 32'hc12fe7dd, 32'hc27d3280, 32'hc2019442, 32'hc0892330, 32'hc1f62513, 32'hc27a04ba};
test_output[8281] = '{32'hc0892330};
test_index[8281] = '{5};
test_input[66256:66263] = '{32'hc28d0fa5, 32'hc1b27425, 32'h4201f911, 32'hbfe37bca, 32'hc2a52f15, 32'hc293d79d, 32'hc1fd37fa, 32'h42b54d9a};
test_output[8282] = '{32'h42b54d9a};
test_index[8282] = '{7};
test_input[66264:66271] = '{32'hc2904987, 32'hc2848ccc, 32'h429c9c4a, 32'hc2a3dedf, 32'hc2a2546e, 32'h40042070, 32'h4268b932, 32'h4249ae45};
test_output[8283] = '{32'h429c9c4a};
test_index[8283] = '{2};
test_input[66272:66279] = '{32'hc1a267e1, 32'h423928e1, 32'hc19a25af, 32'hc0407035, 32'hc27c05df, 32'hc21ce79f, 32'h41fc56f0, 32'h4245dd9d};
test_output[8284] = '{32'h4245dd9d};
test_index[8284] = '{7};
test_input[66280:66287] = '{32'hc21d1e8c, 32'hc2a853ac, 32'h42b445fc, 32'hc2b815ae, 32'hc23891ea, 32'h42b3e71b, 32'h41c2a204, 32'h42b5c197};
test_output[8285] = '{32'h42b5c197};
test_index[8285] = '{7};
test_input[66288:66295] = '{32'h4203595c, 32'h428129f7, 32'hc1c9e3c7, 32'h42570608, 32'hc22b6666, 32'h4095a342, 32'h4284da8b, 32'hc2510e8e};
test_output[8286] = '{32'h4284da8b};
test_index[8286] = '{6};
test_input[66296:66303] = '{32'h42b2c997, 32'hc042a49d, 32'h42c15990, 32'h42b4363a, 32'h420aaee9, 32'hc1703a7b, 32'hc2c07c4c, 32'h4251f9b7};
test_output[8287] = '{32'h42c15990};
test_index[8287] = '{2};
test_input[66304:66311] = '{32'hc16701d5, 32'h42642d1a, 32'h410bbd92, 32'hc1cfaf58, 32'hc298770a, 32'h418f54d3, 32'h41ed1db9, 32'h40927109};
test_output[8288] = '{32'h42642d1a};
test_index[8288] = '{1};
test_input[66312:66319] = '{32'h418ce8ac, 32'h418c6b8b, 32'h4279278b, 32'h42897910, 32'h42909e04, 32'h424aacea, 32'hc2680344, 32'hc29fabda};
test_output[8289] = '{32'h42909e04};
test_index[8289] = '{4};
test_input[66320:66327] = '{32'hc29c10c4, 32'hc29c17a9, 32'hc2b599e4, 32'h41c59dbb, 32'h427afd45, 32'h4124d12d, 32'hc09ce5a8, 32'h42abf460};
test_output[8290] = '{32'h42abf460};
test_index[8290] = '{7};
test_input[66328:66335] = '{32'hc2115108, 32'hc1e6c2f4, 32'h4289a371, 32'hc28d2cc2, 32'h42b53840, 32'hc198b23e, 32'h420fe2e1, 32'h41969b1d};
test_output[8291] = '{32'h42b53840};
test_index[8291] = '{4};
test_input[66336:66343] = '{32'hc2c39985, 32'h4274ecf1, 32'hc259c49e, 32'h41b07930, 32'hc2882c0a, 32'h42634e82, 32'h41be0f7e, 32'h424e47a2};
test_output[8292] = '{32'h4274ecf1};
test_index[8292] = '{1};
test_input[66344:66351] = '{32'hc2b2d960, 32'hc203812b, 32'h421e0b0e, 32'hc2bba2bd, 32'hc1a3a79b, 32'hc28203ab, 32'hc23764c8, 32'h4222aa61};
test_output[8293] = '{32'h4222aa61};
test_index[8293] = '{7};
test_input[66352:66359] = '{32'h42a1105b, 32'h4228528f, 32'hc1b078f6, 32'hc2ba3e53, 32'hc1df8a76, 32'hc29aed6c, 32'h42bda7da, 32'h42a7ce54};
test_output[8294] = '{32'h42bda7da};
test_index[8294] = '{6};
test_input[66360:66367] = '{32'hc2aeefc2, 32'h42067227, 32'h418e3644, 32'hc0978707, 32'h4294f37f, 32'hc20fc2ae, 32'hc1be56a9, 32'hc0c51bf7};
test_output[8295] = '{32'h4294f37f};
test_index[8295] = '{4};
test_input[66368:66375] = '{32'h42c794b5, 32'hc2023b0d, 32'hc098cc59, 32'hc2596e47, 32'hc281915d, 32'h42a34dc5, 32'hc21b3031, 32'h421df944};
test_output[8296] = '{32'h42c794b5};
test_index[8296] = '{0};
test_input[66376:66383] = '{32'hc24bf246, 32'hc285f636, 32'hc2843c3e, 32'hc0e78dbe, 32'h426f995a, 32'h4274fbc1, 32'hc29f7f9d, 32'h425d4680};
test_output[8297] = '{32'h4274fbc1};
test_index[8297] = '{5};
test_input[66384:66391] = '{32'h428fdee9, 32'hc2b690cc, 32'h41d43950, 32'h42c4bb08, 32'hc29cf0aa, 32'hc2bae498, 32'hc23fbf18, 32'hc2adad9e};
test_output[8298] = '{32'h42c4bb08};
test_index[8298] = '{3};
test_input[66392:66399] = '{32'hc251a6b4, 32'hc25aaeea, 32'hc0e1758a, 32'h429ed8ea, 32'hc21461b8, 32'h4227c8fc, 32'h42be5290, 32'h424a353c};
test_output[8299] = '{32'h42be5290};
test_index[8299] = '{6};
test_input[66400:66407] = '{32'h427f8c0c, 32'h41c0f299, 32'h420f611c, 32'hc2a5987b, 32'hc1df06c1, 32'h41ae2312, 32'h42bd2228, 32'hc2b2ee12};
test_output[8300] = '{32'h42bd2228};
test_index[8300] = '{6};
test_input[66408:66415] = '{32'hc2aba8f5, 32'hc2539145, 32'hc25c9216, 32'h42914952, 32'h4281747c, 32'hc2921fbc, 32'hc2a4429f, 32'hc12b107b};
test_output[8301] = '{32'h42914952};
test_index[8301] = '{3};
test_input[66416:66423] = '{32'hc28090fb, 32'h429f56a3, 32'hc1e889a0, 32'h4178c1ad, 32'h41e1b9a9, 32'h420de8a8, 32'h423d389c, 32'hc2c08ba0};
test_output[8302] = '{32'h429f56a3};
test_index[8302] = '{1};
test_input[66424:66431] = '{32'h428a61a5, 32'h41afdf56, 32'hc2ac1bcd, 32'h428fd88f, 32'hc245471c, 32'hc2b9b23c, 32'h40ee0c14, 32'hc23388b4};
test_output[8303] = '{32'h428fd88f};
test_index[8303] = '{3};
test_input[66432:66439] = '{32'h426e078a, 32'hc2407562, 32'hc13190f1, 32'h4297dddb, 32'hbffeb5f7, 32'hc29b16b6, 32'hc2024e45, 32'h41753f33};
test_output[8304] = '{32'h4297dddb};
test_index[8304] = '{3};
test_input[66440:66447] = '{32'hc1e97839, 32'hc2b1898a, 32'hc2a8a81e, 32'hc26a8430, 32'h42b361f2, 32'hc24db1ff, 32'h42b8034a, 32'hc2b98227};
test_output[8305] = '{32'h42b8034a};
test_index[8305] = '{6};
test_input[66448:66455] = '{32'hc2515c19, 32'h41b21249, 32'hc20f5d94, 32'hc216c4f4, 32'h42c33181, 32'h427a0bf9, 32'hc19cc906, 32'h42adce0e};
test_output[8306] = '{32'h42c33181};
test_index[8306] = '{4};
test_input[66456:66463] = '{32'hc1b7564a, 32'hc131bbb4, 32'hc2733f10, 32'h417d0ebc, 32'hc26660ad, 32'hc2b5c534, 32'hc1c92bb8, 32'hc23281ee};
test_output[8307] = '{32'h417d0ebc};
test_index[8307] = '{3};
test_input[66464:66471] = '{32'hc2be35ed, 32'hc260fa64, 32'h42b12a8c, 32'hc2ae434b, 32'h40ebaf39, 32'hc2c1e3b3, 32'h40936e9a, 32'h42c75d3d};
test_output[8308] = '{32'h42c75d3d};
test_index[8308] = '{7};
test_input[66472:66479] = '{32'h42ab87fd, 32'hc2b00bf6, 32'hc2b1c6a5, 32'hc2196b4b, 32'hc244e289, 32'hc26f3f20, 32'hc211c53e, 32'hc2a5ee0c};
test_output[8309] = '{32'h42ab87fd};
test_index[8309] = '{0};
test_input[66480:66487] = '{32'h42978e52, 32'hc1c40034, 32'h42838509, 32'h42aa424f, 32'hc2a7fbea, 32'hc2ac5cec, 32'hc2a482dd, 32'h42975789};
test_output[8310] = '{32'h42aa424f};
test_index[8310] = '{3};
test_input[66488:66495] = '{32'hbfb3689a, 32'hc1d3f001, 32'hc23e90c8, 32'h42597616, 32'hc200cfd8, 32'hbf7cb4a8, 32'h42bdfcfb, 32'hc083a397};
test_output[8311] = '{32'h42bdfcfb};
test_index[8311] = '{6};
test_input[66496:66503] = '{32'hc1612c13, 32'h42867ba4, 32'h4245120a, 32'h42b37c83, 32'h4216774d, 32'h428f3e66, 32'hc2af35fe, 32'hc2600b13};
test_output[8312] = '{32'h42b37c83};
test_index[8312] = '{3};
test_input[66504:66511] = '{32'h42544c79, 32'hc2930901, 32'hc14ccb33, 32'h42bbe834, 32'h41cb63de, 32'hc2969779, 32'hc2a2dd26, 32'hbf70c7fb};
test_output[8313] = '{32'h42bbe834};
test_index[8313] = '{3};
test_input[66512:66519] = '{32'hc29404b4, 32'hc2600c6a, 32'h42439a5b, 32'h42c7f3d2, 32'h41a63064, 32'h427a1fec, 32'h428f146d, 32'h42a47601};
test_output[8314] = '{32'h42c7f3d2};
test_index[8314] = '{3};
test_input[66520:66527] = '{32'h42acec63, 32'hc180d0ea, 32'hc2649302, 32'h40825b52, 32'h42374f9d, 32'h41ffaa79, 32'hc10e8f59, 32'hc25e490d};
test_output[8315] = '{32'h42acec63};
test_index[8315] = '{0};
test_input[66528:66535] = '{32'hc24cb0cb, 32'h418f4899, 32'hc1e30754, 32'hc016a5fd, 32'h422fb184, 32'hc2a572b6, 32'hc2c3c790, 32'hc2b837d1};
test_output[8316] = '{32'h422fb184};
test_index[8316] = '{4};
test_input[66536:66543] = '{32'h40cd4c5e, 32'h40173c0d, 32'hc290100b, 32'h41333958, 32'hc273f165, 32'hc2bf4803, 32'hc2979190, 32'h42c09609};
test_output[8317] = '{32'h42c09609};
test_index[8317] = '{7};
test_input[66544:66551] = '{32'h429ecb9d, 32'hc27e6901, 32'hc25521d4, 32'h42877ce0, 32'hc254866b, 32'hc246954a, 32'hc21162fa, 32'hc2a94ddd};
test_output[8318] = '{32'h429ecb9d};
test_index[8318] = '{0};
test_input[66552:66559] = '{32'h42838ee4, 32'h428072ca, 32'h4265e661, 32'h42024f61, 32'hc2881430, 32'hc1f6088c, 32'h41feb509, 32'h42be7e17};
test_output[8319] = '{32'h42be7e17};
test_index[8319] = '{7};
test_input[66560:66567] = '{32'hc15f3fe3, 32'hc2869601, 32'h42c30ae6, 32'h42a090e6, 32'hc2134780, 32'hc2573902, 32'h40c63fcc, 32'hc2b7a243};
test_output[8320] = '{32'h42c30ae6};
test_index[8320] = '{2};
test_input[66568:66575] = '{32'h4257a942, 32'hc240949d, 32'hc2a94bb1, 32'h3feb8583, 32'hc20bdbb5, 32'hc138ac26, 32'h42637d26, 32'h42b0314d};
test_output[8321] = '{32'h42b0314d};
test_index[8321] = '{7};
test_input[66576:66583] = '{32'h4146a08e, 32'hc1eb5882, 32'h42b04749, 32'hc2b64457, 32'h420991f3, 32'hc1e35f99, 32'h42a72fce, 32'h3fed2989};
test_output[8322] = '{32'h42b04749};
test_index[8322] = '{2};
test_input[66584:66591] = '{32'hc29f1f5c, 32'h42a97164, 32'hc1ec2ff8, 32'h40e79a28, 32'hc299f631, 32'hc295b16d, 32'h41e27645, 32'h40f1fa31};
test_output[8323] = '{32'h42a97164};
test_index[8323] = '{1};
test_input[66592:66599] = '{32'hc282872f, 32'hc24da1ee, 32'h42b8f326, 32'h42ba6460, 32'hc216ce44, 32'h42a9ad8a, 32'h421c6e90, 32'h427f53dd};
test_output[8324] = '{32'h42ba6460};
test_index[8324] = '{3};
test_input[66600:66607] = '{32'h423e190e, 32'hc2396e6d, 32'hc291f453, 32'hc1647ab2, 32'hc21be96b, 32'hc191af5a, 32'hc2996900, 32'hc2061a8e};
test_output[8325] = '{32'h423e190e};
test_index[8325] = '{0};
test_input[66608:66615] = '{32'hc2897079, 32'h40b1c545, 32'hc2b3d32c, 32'h42806777, 32'h4273b9dc, 32'h3fc0ebf8, 32'h421cccc0, 32'h42b7f0b4};
test_output[8326] = '{32'h42b7f0b4};
test_index[8326] = '{7};
test_input[66616:66623] = '{32'h41c1e55b, 32'hc1d7e6a1, 32'hc2b37d4b, 32'h429ad28b, 32'h42adee1e, 32'hc2b90833, 32'hc1e0b996, 32'h410b5e2e};
test_output[8327] = '{32'h42adee1e};
test_index[8327] = '{4};
test_input[66624:66631] = '{32'hc1d17d88, 32'h42807ae4, 32'h4206288a, 32'h41b07ed5, 32'h42a3cd8e, 32'hc1ad6b68, 32'h420d1c4c, 32'hc1aef541};
test_output[8328] = '{32'h42a3cd8e};
test_index[8328] = '{4};
test_input[66632:66639] = '{32'h42a10065, 32'hc298e603, 32'hc1d4b6b7, 32'hc2b2a435, 32'h42b567cf, 32'h429ac498, 32'h42332b9d, 32'hc2b0cb7b};
test_output[8329] = '{32'h42b567cf};
test_index[8329] = '{4};
test_input[66640:66647] = '{32'h42817223, 32'h427cdb3a, 32'hc25f835a, 32'hc2a8ef47, 32'hc22bcbad, 32'h423b6eca, 32'hc20db253, 32'hc296652c};
test_output[8330] = '{32'h42817223};
test_index[8330] = '{0};
test_input[66648:66655] = '{32'h4220447f, 32'hc292eea3, 32'h42062ea4, 32'h404a5f9b, 32'hc20bceb1, 32'hc0f8c5c2, 32'hc26f439c, 32'hc2a90d16};
test_output[8331] = '{32'h4220447f};
test_index[8331] = '{0};
test_input[66656:66663] = '{32'hc2878835, 32'hc2b1fe72, 32'h420b9a54, 32'hc23b44f4, 32'hc273ed03, 32'hc28abbd8, 32'hc28f92e8, 32'hc25200eb};
test_output[8332] = '{32'h420b9a54};
test_index[8332] = '{2};
test_input[66664:66671] = '{32'h4296b9c1, 32'h428adf86, 32'hc1393632, 32'hc1cf0dab, 32'hc2a2fd5d, 32'hc2ab5f55, 32'hc191d8c3, 32'h4285619b};
test_output[8333] = '{32'h4296b9c1};
test_index[8333] = '{0};
test_input[66672:66679] = '{32'h4127e40a, 32'hc2b24388, 32'h42b5d563, 32'h41098964, 32'hc28a8aac, 32'hc2947b58, 32'h4165cbb3, 32'h429f95ce};
test_output[8334] = '{32'h42b5d563};
test_index[8334] = '{2};
test_input[66680:66687] = '{32'h42bf1166, 32'h429ac7bd, 32'hc204f037, 32'hc299be9f, 32'h422e784b, 32'h42b61923, 32'hc235f99e, 32'hc2c13fdd};
test_output[8335] = '{32'h42bf1166};
test_index[8335] = '{0};
test_input[66688:66695] = '{32'h412c2d36, 32'h41c7b43b, 32'h42bb49b9, 32'h428a93b0, 32'hc2271423, 32'hc22d4dbf, 32'hc2b78e5a, 32'h42767002};
test_output[8336] = '{32'h42bb49b9};
test_index[8336] = '{2};
test_input[66696:66703] = '{32'hc2868817, 32'h42356ea2, 32'hc23491dc, 32'hc20c3451, 32'hc28832b2, 32'h41f8dc9c, 32'h42232e98, 32'h424847e6};
test_output[8337] = '{32'h424847e6};
test_index[8337] = '{7};
test_input[66704:66711] = '{32'hbe66320b, 32'h3fe5fae6, 32'hc25ac086, 32'h4231a69b, 32'hc29df6b8, 32'h42986bb8, 32'hc28ae6b4, 32'h42a6ed4a};
test_output[8338] = '{32'h42a6ed4a};
test_index[8338] = '{7};
test_input[66712:66719] = '{32'h42405def, 32'hc1bea152, 32'hc22877e4, 32'hc2588783, 32'h4293afe0, 32'h42b8afba, 32'hc280a5aa, 32'hc2261995};
test_output[8339] = '{32'h42b8afba};
test_index[8339] = '{5};
test_input[66720:66727] = '{32'h41258117, 32'h42393d56, 32'hc1b5de79, 32'hc29505ba, 32'hc11593f0, 32'h42859e41, 32'hc2aa73a1, 32'h41215934};
test_output[8340] = '{32'h42859e41};
test_index[8340] = '{5};
test_input[66728:66735] = '{32'h42a32dd3, 32'h428c0392, 32'hc1a6c4b0, 32'h42c2d837, 32'h429bc721, 32'hc2169d5b, 32'h42afae9f, 32'h41388f30};
test_output[8341] = '{32'h42c2d837};
test_index[8341] = '{3};
test_input[66736:66743] = '{32'hc2bf1b0f, 32'h4262467b, 32'hc25511c1, 32'h428a306d, 32'hc24e5907, 32'hc1d1d241, 32'hc1069951, 32'h4216aa0f};
test_output[8342] = '{32'h428a306d};
test_index[8342] = '{3};
test_input[66744:66751] = '{32'h4270b36a, 32'hc296c885, 32'h425c4110, 32'hc2992ec9, 32'h42027440, 32'hc25f0b42, 32'hc284142e, 32'hc12b81ea};
test_output[8343] = '{32'h4270b36a};
test_index[8343] = '{0};
test_input[66752:66759] = '{32'h4289d36a, 32'hc18ce05e, 32'hc279271d, 32'hc08db81a, 32'hc2af8ed9, 32'hc2514d9b, 32'h415becda, 32'h4254483d};
test_output[8344] = '{32'h4289d36a};
test_index[8344] = '{0};
test_input[66760:66767] = '{32'h418c5d17, 32'hc28b91e9, 32'h42811794, 32'h4154268a, 32'hc2bdc0ec, 32'hc1a2dfb8, 32'h42ae1ea7, 32'hc12ef05d};
test_output[8345] = '{32'h42ae1ea7};
test_index[8345] = '{6};
test_input[66768:66775] = '{32'hbf95d0eb, 32'hc22fc2b9, 32'hc28d59c5, 32'h42685228, 32'hc26af38f, 32'hc28aeaaa, 32'h422bdedc, 32'h427e17cc};
test_output[8346] = '{32'h427e17cc};
test_index[8346] = '{7};
test_input[66776:66783] = '{32'hc2874882, 32'h425cad0c, 32'h40c115aa, 32'hc204d9d1, 32'h4138cc8d, 32'hc2a967f7, 32'h429958ee, 32'h4134e7d8};
test_output[8347] = '{32'h429958ee};
test_index[8347] = '{6};
test_input[66784:66791] = '{32'h422aba74, 32'hc2700854, 32'hc045cf0c, 32'h413dcc9a, 32'h42169435, 32'hc27c10cf, 32'h426b1c86, 32'h424e4754};
test_output[8348] = '{32'h426b1c86};
test_index[8348] = '{6};
test_input[66792:66799] = '{32'h42c263f8, 32'h42c682be, 32'hc1e58586, 32'hc29b2c55, 32'h428821b1, 32'h425b8fa0, 32'h41130630, 32'hc1559dbd};
test_output[8349] = '{32'h42c682be};
test_index[8349] = '{1};
test_input[66800:66807] = '{32'h428224ff, 32'hc2af067e, 32'hc2234af2, 32'hc237f486, 32'hc13c8ca7, 32'hc26746c6, 32'hc2816d00, 32'hc1bc2453};
test_output[8350] = '{32'h428224ff};
test_index[8350] = '{0};
test_input[66808:66815] = '{32'h429c992d, 32'h425167eb, 32'h42a51086, 32'hc249c41f, 32'hc19661ae, 32'hc29d22ef, 32'hbfcf49b3, 32'hc239e021};
test_output[8351] = '{32'h42a51086};
test_index[8351] = '{2};
test_input[66816:66823] = '{32'hc2bcf448, 32'hc2713230, 32'h42bbfebe, 32'hc2c564a5, 32'hc19d3a95, 32'h427f42ea, 32'h42c34ebb, 32'hc20f032f};
test_output[8352] = '{32'h42c34ebb};
test_index[8352] = '{6};
test_input[66824:66831] = '{32'h42a31a44, 32'hc1d05ef0, 32'h419b2772, 32'h42490787, 32'h42922638, 32'h42846825, 32'h42762209, 32'h4298df52};
test_output[8353] = '{32'h42a31a44};
test_index[8353] = '{0};
test_input[66832:66839] = '{32'h42b7e597, 32'hc29b8b68, 32'hc230451c, 32'hc246e0d5, 32'hc1eb058e, 32'h421b6854, 32'h428c873a, 32'hc29ff1c2};
test_output[8354] = '{32'h42b7e597};
test_index[8354] = '{0};
test_input[66840:66847] = '{32'hc2783e61, 32'h425bdcf8, 32'h41ee1684, 32'h4262d780, 32'h415200b7, 32'hc2a7d0ed, 32'h42a92cc6, 32'h4211a1a7};
test_output[8355] = '{32'h42a92cc6};
test_index[8355] = '{6};
test_input[66848:66855] = '{32'h428083a5, 32'h4066e5a2, 32'h42837f6d, 32'h41d910fb, 32'h421b0682, 32'h4293d72c, 32'hc1a1d13a, 32'hc2770aac};
test_output[8356] = '{32'h4293d72c};
test_index[8356] = '{5};
test_input[66856:66863] = '{32'h42baa094, 32'hbf76cf6e, 32'h424cb671, 32'h4281b4d0, 32'h41ba67bc, 32'hc1b5f562, 32'hc2579dc4, 32'hc1d35996};
test_output[8357] = '{32'h42baa094};
test_index[8357] = '{0};
test_input[66864:66871] = '{32'h42294f63, 32'h41b178c5, 32'h422bafe5, 32'hc2241dc9, 32'h4294602b, 32'hc22fc514, 32'h414060b2, 32'h425856ab};
test_output[8358] = '{32'h4294602b};
test_index[8358] = '{4};
test_input[66872:66879] = '{32'hc1e2f896, 32'h428b8683, 32'hc2b29da9, 32'hc2a563bb, 32'h42a5053f, 32'h4129a4cb, 32'h42c13bd5, 32'h42820516};
test_output[8359] = '{32'h42c13bd5};
test_index[8359] = '{6};
test_input[66880:66887] = '{32'hc20d90e9, 32'h42b9768c, 32'hc25aaaa4, 32'h42ad7e14, 32'h42b8bba1, 32'hc2206229, 32'h41dd6efc, 32'h41cd9979};
test_output[8360] = '{32'h42b9768c};
test_index[8360] = '{1};
test_input[66888:66895] = '{32'h4257c91c, 32'hc25d203f, 32'hc21cf901, 32'hc21c2a6e, 32'h428394a8, 32'h42878d30, 32'h4178bb10, 32'hc28fa1a6};
test_output[8361] = '{32'h42878d30};
test_index[8361] = '{5};
test_input[66896:66903] = '{32'hc1a79e36, 32'h42827e18, 32'hc2bf22dd, 32'h42b8c4a0, 32'h42bedd9c, 32'hc22ac81d, 32'hc209010a, 32'h42aeab5a};
test_output[8362] = '{32'h42bedd9c};
test_index[8362] = '{4};
test_input[66904:66911] = '{32'hc2a0e5d9, 32'hc2b43add, 32'h4285af78, 32'h4269c1a7, 32'h41c6ca14, 32'h42731c44, 32'hc2b1b1b9, 32'h42985d31};
test_output[8363] = '{32'h42985d31};
test_index[8363] = '{7};
test_input[66912:66919] = '{32'hc22e5bea, 32'hc2a8f09e, 32'hc1c1c3d5, 32'hc2b92095, 32'h42ad01c3, 32'hc28759da, 32'h402ca58d, 32'hc1ad6695};
test_output[8364] = '{32'h42ad01c3};
test_index[8364] = '{4};
test_input[66920:66927] = '{32'h41028b69, 32'h42b03e0c, 32'hc291608d, 32'h42ac96e9, 32'h425e00cf, 32'hc1c6752c, 32'hc281fac1, 32'h42b3ddbe};
test_output[8365] = '{32'h42b3ddbe};
test_index[8365] = '{7};
test_input[66928:66935] = '{32'hc293a863, 32'h425b8566, 32'h42b0b9ea, 32'h42818ad9, 32'h40f96b78, 32'h42811214, 32'hc090cf39, 32'hc21490c1};
test_output[8366] = '{32'h42b0b9ea};
test_index[8366] = '{2};
test_input[66936:66943] = '{32'hc2818d27, 32'hc2b30918, 32'hc09c4fed, 32'hc29d39e7, 32'h426ba7ca, 32'h409abee0, 32'h423662f3, 32'h400247dc};
test_output[8367] = '{32'h426ba7ca};
test_index[8367] = '{4};
test_input[66944:66951] = '{32'hc269b8a2, 32'h4261139a, 32'hc21dd1fc, 32'h421a6d0a, 32'h4200a2c7, 32'h420f6a2c, 32'h429a4322, 32'hc2089eb9};
test_output[8368] = '{32'h429a4322};
test_index[8368] = '{6};
test_input[66952:66959] = '{32'h42686b61, 32'h42479953, 32'hc22288d0, 32'h41a1b28f, 32'h429fb34f, 32'h41ed9143, 32'h422553d5, 32'hc0f47cdc};
test_output[8369] = '{32'h429fb34f};
test_index[8369] = '{4};
test_input[66960:66967] = '{32'h41a04957, 32'h426d8426, 32'hc1e00cef, 32'h42780a70, 32'hc27963f2, 32'hc2ac6b3d, 32'hc14d589f, 32'h4069a65c};
test_output[8370] = '{32'h42780a70};
test_index[8370] = '{3};
test_input[66968:66975] = '{32'hc2b24144, 32'h4222b0e8, 32'h4264a84a, 32'h415523e3, 32'h41ebb953, 32'hc2259a68, 32'h4266a8b5, 32'hc204e8eb};
test_output[8371] = '{32'h4266a8b5};
test_index[8371] = '{6};
test_input[66976:66983] = '{32'hc204ad3d, 32'h411301ad, 32'h42866279, 32'hc20b44ba, 32'hc1b5b046, 32'hc2bf4a5b, 32'h42479f05, 32'hc1bd4c4b};
test_output[8372] = '{32'h42866279};
test_index[8372] = '{2};
test_input[66984:66991] = '{32'h41bce546, 32'h41b1814b, 32'h42567002, 32'hc281488a, 32'hc0f56d05, 32'h4209c8c4, 32'h4292fd28, 32'hc0c13a97};
test_output[8373] = '{32'h4292fd28};
test_index[8373] = '{6};
test_input[66992:66999] = '{32'hc24bbcfb, 32'hc29596ed, 32'hc29129b2, 32'hc2a104fa, 32'hc11b25dd, 32'h425c71db, 32'h4239b3c7, 32'h42bff325};
test_output[8374] = '{32'h42bff325};
test_index[8374] = '{7};
test_input[67000:67007] = '{32'h429a91d0, 32'h424e4578, 32'h42845b05, 32'hc2ab5aa8, 32'h422965f6, 32'h3f27fc41, 32'h42368b8d, 32'h42c0c6e9};
test_output[8375] = '{32'h42c0c6e9};
test_index[8375] = '{7};
test_input[67008:67015] = '{32'hc16d1ab2, 32'h4282699c, 32'hc1801dba, 32'h42824703, 32'h42beb044, 32'hc2c4f4cb, 32'hc1fbbea7, 32'hc20290bf};
test_output[8376] = '{32'h42beb044};
test_index[8376] = '{4};
test_input[67016:67023] = '{32'hc26c0ff6, 32'hc28593d4, 32'h42b8f3a1, 32'hc21a94d5, 32'h422ea668, 32'hc2c31ab7, 32'h42a9b1a5, 32'h41c04c92};
test_output[8377] = '{32'h42b8f3a1};
test_index[8377] = '{2};
test_input[67024:67031] = '{32'h427e16c9, 32'hc2046ae7, 32'h41c056af, 32'h42516738, 32'h4250c6fc, 32'h4280d2fe, 32'hbf9a4e96, 32'h4240226a};
test_output[8378] = '{32'h4280d2fe};
test_index[8378] = '{5};
test_input[67032:67039] = '{32'hc2b80b79, 32'hc2569d4e, 32'hc25b541b, 32'hc24ab1a6, 32'h42bea7df, 32'hc230531f, 32'hc2772744, 32'h42b5ed73};
test_output[8379] = '{32'h42bea7df};
test_index[8379] = '{4};
test_input[67040:67047] = '{32'h421d7e99, 32'h42880f2a, 32'hc20d9ee3, 32'h42bfbd05, 32'h4016f25d, 32'hc2b08553, 32'hc2857c98, 32'h41c96902};
test_output[8380] = '{32'h42bfbd05};
test_index[8380] = '{3};
test_input[67048:67055] = '{32'hc21b9943, 32'hc1778fd6, 32'h42ae4276, 32'h420ac250, 32'h412fa864, 32'hbedc9890, 32'h42c2d2f7, 32'hc2a1d573};
test_output[8381] = '{32'h42c2d2f7};
test_index[8381] = '{6};
test_input[67056:67063] = '{32'h42681da4, 32'hc2ab9ca5, 32'h42b870a4, 32'h422de95b, 32'h425a73f7, 32'h421bd844, 32'h418c76d3, 32'hc2823016};
test_output[8382] = '{32'h42b870a4};
test_index[8382] = '{2};
test_input[67064:67071] = '{32'hc23ada4a, 32'h429ae769, 32'h42c4719a, 32'hc2940e08, 32'hc2c3b137, 32'hc231413d, 32'h422b3fb5, 32'h4194f9e1};
test_output[8383] = '{32'h42c4719a};
test_index[8383] = '{2};
test_input[67072:67079] = '{32'h42bd2326, 32'hc2583d48, 32'h42753bf5, 32'hc289a2ee, 32'h42b346ed, 32'h413f245e, 32'h429fd236, 32'h4148065d};
test_output[8384] = '{32'h42bd2326};
test_index[8384] = '{0};
test_input[67080:67087] = '{32'hc2bea3c5, 32'h42a81516, 32'hc2669139, 32'hc2c1dd14, 32'hc2b18058, 32'hc2024d6a, 32'hc13c79a9, 32'hc2113b4a};
test_output[8385] = '{32'h42a81516};
test_index[8385] = '{1};
test_input[67088:67095] = '{32'hc24426d8, 32'h427ae8b3, 32'h42a01a62, 32'h41506ac5, 32'h419fa60a, 32'h42af28f9, 32'h42483f4e, 32'hc0b40bd4};
test_output[8386] = '{32'h42af28f9};
test_index[8386] = '{5};
test_input[67096:67103] = '{32'h412ea7e5, 32'h4186faa7, 32'hc1c87f03, 32'h42a88eb6, 32'h42870636, 32'hc2862923, 32'h42811bc6, 32'h42b3ca5b};
test_output[8387] = '{32'h42b3ca5b};
test_index[8387] = '{7};
test_input[67104:67111] = '{32'hc2a21915, 32'hc2c0638a, 32'hc2a71a67, 32'hc257ee32, 32'hc166e083, 32'hc1b26c25, 32'hc15c8dd7, 32'hc2b19a7c};
test_output[8388] = '{32'hc15c8dd7};
test_index[8388] = '{6};
test_input[67112:67119] = '{32'h424cfb62, 32'hc29ab3b5, 32'h42bd0594, 32'hc27020f7, 32'hc2b2abf1, 32'hbfc9c35b, 32'hc22805a7, 32'hc1429421};
test_output[8389] = '{32'h42bd0594};
test_index[8389] = '{2};
test_input[67120:67127] = '{32'h421f7b23, 32'h4191fc47, 32'hc15ce9bf, 32'h42bc7db6, 32'hc1afa24b, 32'hc29f6602, 32'h41815871, 32'hc23f90d4};
test_output[8390] = '{32'h42bc7db6};
test_index[8390] = '{3};
test_input[67128:67135] = '{32'hc0e279c0, 32'hc2924b6a, 32'h4054dfaf, 32'hc28669a0, 32'h42208b87, 32'h42b0c342, 32'h42b3beab, 32'hc2b48431};
test_output[8391] = '{32'h42b3beab};
test_index[8391] = '{6};
test_input[67136:67143] = '{32'hc2bac47d, 32'hc214d35d, 32'hc252610b, 32'h42679b0d, 32'hc18ce203, 32'hc1d74726, 32'hc258de1c, 32'h42737a0c};
test_output[8392] = '{32'h42737a0c};
test_index[8392] = '{7};
test_input[67144:67151] = '{32'hc1bd75da, 32'h42a29e52, 32'hc25e6070, 32'h4268d860, 32'h42b9db76, 32'hc20b6bb0, 32'hc1c6a6d0, 32'hc23ac278};
test_output[8393] = '{32'h42b9db76};
test_index[8393] = '{4};
test_input[67152:67159] = '{32'hc237b96d, 32'hc22b8c62, 32'h421d7b47, 32'hc29741e9, 32'hc21db336, 32'hc19e024c, 32'hc26fd757, 32'h41d7a686};
test_output[8394] = '{32'h421d7b47};
test_index[8394] = '{2};
test_input[67160:67167] = '{32'h429d8541, 32'hc274fabd, 32'h40deb6e4, 32'hc2bde2d2, 32'hc2a24dd0, 32'h420468e7, 32'h4212b4ee, 32'h42869ce1};
test_output[8395] = '{32'h429d8541};
test_index[8395] = '{0};
test_input[67168:67175] = '{32'h42b6d1f2, 32'h41459c3d, 32'h41cec98b, 32'h409f9300, 32'hc2526aa1, 32'hc2a4358e, 32'hc28aa76b, 32'hc28ed0b7};
test_output[8396] = '{32'h42b6d1f2};
test_index[8396] = '{0};
test_input[67176:67183] = '{32'h42bc82f1, 32'h42284b29, 32'hc2218d7e, 32'h41a5e8b9, 32'h42aa6bfe, 32'hc1fafb74, 32'h41a98977, 32'h42c6bf2c};
test_output[8397] = '{32'h42c6bf2c};
test_index[8397] = '{7};
test_input[67184:67191] = '{32'hc203709c, 32'hc28406f0, 32'hc2531439, 32'hc22c8dfd, 32'hc26d7575, 32'hc19eb2ff, 32'h40acad23, 32'hc29eb201};
test_output[8398] = '{32'h40acad23};
test_index[8398] = '{6};
test_input[67192:67199] = '{32'hc15f81ec, 32'hc2a84889, 32'h41f40781, 32'h4001710c, 32'hc2570c6a, 32'h425f47fe, 32'h429fe343, 32'hc16bc9da};
test_output[8399] = '{32'h429fe343};
test_index[8399] = '{6};
test_input[67200:67207] = '{32'h41007991, 32'hc1de1718, 32'hc26d9f02, 32'h4245d23b, 32'h423698a2, 32'hc27bcda2, 32'hc2a21f45, 32'h4246cf4d};
test_output[8400] = '{32'h4246cf4d};
test_index[8400] = '{7};
test_input[67208:67215] = '{32'hc11909ec, 32'h426a8275, 32'hc14af83b, 32'h42bf668a, 32'h425f92c0, 32'hc276ccd6, 32'h42a144fb, 32'hc1b87094};
test_output[8401] = '{32'h42bf668a};
test_index[8401] = '{3};
test_input[67216:67223] = '{32'h40c45508, 32'h4292c5b7, 32'hc062f1ad, 32'h4247c2a6, 32'h4250dc5c, 32'h4129a496, 32'h419c13e8, 32'hc22e3a77};
test_output[8402] = '{32'h4292c5b7};
test_index[8402] = '{1};
test_input[67224:67231] = '{32'hc2c02461, 32'h42707093, 32'h41e3f10f, 32'hc2ab4559, 32'h42982260, 32'h428ddebd, 32'h42329a8d, 32'h42b06237};
test_output[8403] = '{32'h42b06237};
test_index[8403] = '{7};
test_input[67232:67239] = '{32'hc2a9c386, 32'h4070b01d, 32'h42399177, 32'hc25912ef, 32'hc2abee6b, 32'h4283b263, 32'h4171c731, 32'h41025965};
test_output[8404] = '{32'h4283b263};
test_index[8404] = '{5};
test_input[67240:67247] = '{32'h426a0831, 32'hc28b222f, 32'hc2bbd175, 32'hc2c5c4fc, 32'hbf73036c, 32'hc2859018, 32'h427fb918, 32'hc20aedf8};
test_output[8405] = '{32'h427fb918};
test_index[8405] = '{6};
test_input[67248:67255] = '{32'hc20dfe65, 32'h4295b095, 32'hc25bc073, 32'h42aa5896, 32'hc29df537, 32'h426b6383, 32'h424c7f46, 32'h3f27799f};
test_output[8406] = '{32'h42aa5896};
test_index[8406] = '{3};
test_input[67256:67263] = '{32'hc085225b, 32'hc276b39b, 32'h4211481e, 32'hc2957272, 32'h421658b1, 32'hc1df5c6b, 32'h425b1adf, 32'h40fdb201};
test_output[8407] = '{32'h425b1adf};
test_index[8407] = '{6};
test_input[67264:67271] = '{32'h40669a3b, 32'h42b42e03, 32'hc1878414, 32'hc19c3d51, 32'h414ffd69, 32'hc215d86c, 32'h42294ec9, 32'hc2a61559};
test_output[8408] = '{32'h42b42e03};
test_index[8408] = '{1};
test_input[67272:67279] = '{32'hc226e5df, 32'hc20e48c2, 32'hc29ad6ba, 32'h427ec2dc, 32'hc1c14bd5, 32'hc2c222be, 32'hc15bcda9, 32'hc29c1ab8};
test_output[8409] = '{32'h427ec2dc};
test_index[8409] = '{3};
test_input[67280:67287] = '{32'h41c7317c, 32'hc104c91c, 32'h42985146, 32'hc2946bcb, 32'hc2a7cac2, 32'h42bce1a2, 32'hc25d7658, 32'hc236fa5d};
test_output[8410] = '{32'h42bce1a2};
test_index[8410] = '{5};
test_input[67288:67295] = '{32'h420f157a, 32'h413fd6d0, 32'hc239535e, 32'h4273dc28, 32'h4147a1d7, 32'h42a31fe1, 32'h4283301b, 32'h421cb45a};
test_output[8411] = '{32'h42a31fe1};
test_index[8411] = '{5};
test_input[67296:67303] = '{32'hc1e1d284, 32'h42acdcea, 32'hc1718c87, 32'h40b88129, 32'hc1e790c5, 32'h42c0b439, 32'hc2a4e4e9, 32'hc18b31cb};
test_output[8412] = '{32'h42c0b439};
test_index[8412] = '{5};
test_input[67304:67311] = '{32'h42afd512, 32'hc18a55d1, 32'h3faf32b7, 32'hc2baf0b2, 32'h41e9916a, 32'h4293e0f9, 32'h42bbafd5, 32'hc10ba696};
test_output[8413] = '{32'h42bbafd5};
test_index[8413] = '{6};
test_input[67312:67319] = '{32'h4231a825, 32'hc1be3232, 32'h41b454b1, 32'hc16b8c51, 32'hc29b24ef, 32'hc22e2aea, 32'h429be419, 32'h42b9a42f};
test_output[8414] = '{32'h42b9a42f};
test_index[8414] = '{7};
test_input[67320:67327] = '{32'h42916d6c, 32'h4203a883, 32'h420fceb2, 32'h4285295e, 32'h4288ce80, 32'hc25fdb9d, 32'h41c5323e, 32'hc1d90e80};
test_output[8415] = '{32'h42916d6c};
test_index[8415] = '{0};
test_input[67328:67335] = '{32'hc2335434, 32'hc2bd772b, 32'hc190cd0a, 32'h428be0ef, 32'h428bd121, 32'hc2a11a04, 32'hc21e9f44, 32'hc2588fbc};
test_output[8416] = '{32'h428be0ef};
test_index[8416] = '{3};
test_input[67336:67343] = '{32'h41df8682, 32'h42a09bea, 32'h41823f93, 32'hc2564c64, 32'h41a2c08f, 32'hc21dade0, 32'hc208f840, 32'hc1a8f78b};
test_output[8417] = '{32'h42a09bea};
test_index[8417] = '{1};
test_input[67344:67351] = '{32'hc297b4b5, 32'h41c426df, 32'h4243697e, 32'h42474b8b, 32'h415f514b, 32'hc0569faf, 32'hc2c4f0a6, 32'hc24832a7};
test_output[8418] = '{32'h42474b8b};
test_index[8418] = '{3};
test_input[67352:67359] = '{32'hc1bdd7af, 32'h4215299f, 32'hc23718c0, 32'h4247dd88, 32'hc2197c90, 32'hbf87a5ee, 32'hc297cd1d, 32'hc21b5cfe};
test_output[8419] = '{32'h4247dd88};
test_index[8419] = '{3};
test_input[67360:67367] = '{32'hbf52d27c, 32'hc2ba0934, 32'h4204c960, 32'hbf86e18a, 32'h429b28f8, 32'h42b42477, 32'hc279a779, 32'hc2771a10};
test_output[8420] = '{32'h42b42477};
test_index[8420] = '{5};
test_input[67368:67375] = '{32'hc22534b3, 32'h425b3b84, 32'h4287e370, 32'hbd894fb1, 32'h423b4ad4, 32'h42b60356, 32'h4223cda2, 32'hc2a69faa};
test_output[8421] = '{32'h42b60356};
test_index[8421] = '{5};
test_input[67376:67383] = '{32'hc240be9d, 32'h4284abbf, 32'hc2a6659f, 32'h4298b904, 32'h41801382, 32'h42838002, 32'h42a1f683, 32'h42b7be5d};
test_output[8422] = '{32'h42b7be5d};
test_index[8422] = '{7};
test_input[67384:67391] = '{32'hc283ec87, 32'hc12a46f5, 32'hc2857ca5, 32'h42613152, 32'hc2bd4030, 32'h424b26f2, 32'hc2628810, 32'h42bc14be};
test_output[8423] = '{32'h42bc14be};
test_index[8423] = '{7};
test_input[67392:67399] = '{32'h41078bb3, 32'h42579448, 32'h4249310d, 32'h41c5250b, 32'hc02b6c54, 32'hc258334c, 32'hc135283d, 32'h429929d8};
test_output[8424] = '{32'h429929d8};
test_index[8424] = '{7};
test_input[67400:67407] = '{32'h41dc8fba, 32'h428642c4, 32'hc0ba328e, 32'h429cf36a, 32'h421fbd6c, 32'hc2c50424, 32'hc2b348e2, 32'h424e0ea6};
test_output[8425] = '{32'h429cf36a};
test_index[8425] = '{3};
test_input[67408:67415] = '{32'h41fc525a, 32'h42771b2c, 32'hc1791dba, 32'h421f6cc1, 32'h3ea97dde, 32'h42900e39, 32'h415ef5f3, 32'hc17c8e85};
test_output[8426] = '{32'h42900e39};
test_index[8426] = '{5};
test_input[67416:67423] = '{32'hc2a18bd7, 32'hc289cbcd, 32'hc2ad70b3, 32'hc1e6916a, 32'h42bc36fd, 32'h42b0d7d2, 32'hc23ce412, 32'hc228f9b8};
test_output[8427] = '{32'h42bc36fd};
test_index[8427] = '{4};
test_input[67424:67431] = '{32'hc246e23f, 32'h41b47a19, 32'h42b887aa, 32'h419ce4d5, 32'hc1c08a91, 32'hc2b9ffc6, 32'h4258140d, 32'hc1ed95fc};
test_output[8428] = '{32'h42b887aa};
test_index[8428] = '{2};
test_input[67432:67439] = '{32'h42163391, 32'h423f124b, 32'h4241ce05, 32'hc2c67624, 32'hc2b2dd42, 32'hc245dc8f, 32'h415b1c1f, 32'hc02b86f1};
test_output[8429] = '{32'h4241ce05};
test_index[8429] = '{2};
test_input[67440:67447] = '{32'hc2694e9e, 32'h40b5ed06, 32'h42a762a2, 32'h421f0410, 32'h42819745, 32'h415434eb, 32'hc25eed98, 32'hc205e828};
test_output[8430] = '{32'h42a762a2};
test_index[8430] = '{2};
test_input[67448:67455] = '{32'hc2c3b16c, 32'hc22ea843, 32'h42713ee4, 32'h42282233, 32'hc10ac3a2, 32'h422cf79c, 32'hc1fe0e88, 32'h420395f0};
test_output[8431] = '{32'h42713ee4};
test_index[8431] = '{2};
test_input[67456:67463] = '{32'hc2c78243, 32'h419c5f75, 32'h42646376, 32'h4250d733, 32'h42b7abdc, 32'hc299de0d, 32'hc26df6e2, 32'hc22e657c};
test_output[8432] = '{32'h42b7abdc};
test_index[8432] = '{4};
test_input[67464:67471] = '{32'h4296d97b, 32'hc137ce3d, 32'h42855cd5, 32'hc28078c6, 32'hc020e01c, 32'h416684e0, 32'h41816a04, 32'hc2a4762d};
test_output[8433] = '{32'h4296d97b};
test_index[8433] = '{0};
test_input[67472:67479] = '{32'hc1dffda7, 32'hc2bd4ace, 32'hc218f950, 32'hc2b56094, 32'hc2927e44, 32'hc29b27df, 32'hc2c17b98, 32'h42282589};
test_output[8434] = '{32'h42282589};
test_index[8434] = '{7};
test_input[67480:67487] = '{32'hc29efa87, 32'h41b6f4f2, 32'hc1dd80d6, 32'h41907bd1, 32'h42bf6915, 32'hc27d19d0, 32'hc1ad7eea, 32'h42a5be97};
test_output[8435] = '{32'h42bf6915};
test_index[8435] = '{4};
test_input[67488:67495] = '{32'hc1ee1ccc, 32'hc2bb280e, 32'hc2a1e00d, 32'hc0aace3a, 32'h419f8daf, 32'hc1b515ef, 32'h41d0bddf, 32'h4259a05c};
test_output[8436] = '{32'h4259a05c};
test_index[8436] = '{7};
test_input[67496:67503] = '{32'hc2b16e76, 32'hc1aeff21, 32'hc2093bd6, 32'h41b3d04a, 32'h426b3a89, 32'h428447da, 32'h409720f7, 32'h41183f44};
test_output[8437] = '{32'h428447da};
test_index[8437] = '{5};
test_input[67504:67511] = '{32'hc244918a, 32'h3ededa51, 32'h424d61d7, 32'hc2a3bf4b, 32'hc2c56b49, 32'hc22800ec, 32'hc23dda6f, 32'hc271dfa1};
test_output[8438] = '{32'h424d61d7};
test_index[8438] = '{2};
test_input[67512:67519] = '{32'hc1f4bbf4, 32'hc11ffd62, 32'h42acefb8, 32'h4262bf56, 32'h428bd3ad, 32'hbf148fa7, 32'hc29b2c48, 32'h428d7cf6};
test_output[8439] = '{32'h42acefb8};
test_index[8439] = '{2};
test_input[67520:67527] = '{32'h418563be, 32'h41b15cc6, 32'hbf5bb583, 32'h420fef72, 32'hc1b483c7, 32'hc208d5f4, 32'h42a7a912, 32'h420b723f};
test_output[8440] = '{32'h42a7a912};
test_index[8440] = '{6};
test_input[67528:67535] = '{32'h4276bab1, 32'hc2212619, 32'h42b7cde2, 32'hc2abf990, 32'hc262d04a, 32'h400add40, 32'hc294b933, 32'h4290ba76};
test_output[8441] = '{32'h42b7cde2};
test_index[8441] = '{2};
test_input[67536:67543] = '{32'h422b1699, 32'hc13110f9, 32'hc0ba6bda, 32'hc1a9aff9, 32'hc21217d9, 32'hc29e024e, 32'h41e5d1e9, 32'hc289a0a4};
test_output[8442] = '{32'h422b1699};
test_index[8442] = '{0};
test_input[67544:67551] = '{32'hc15385d2, 32'h42676d0d, 32'h41efc1f2, 32'hc28761da, 32'hc2adc82a, 32'hc251ea2c, 32'h42bc727e, 32'hc2ab6000};
test_output[8443] = '{32'h42bc727e};
test_index[8443] = '{6};
test_input[67552:67559] = '{32'hc1ce429e, 32'h42bf67ca, 32'hc2b5cc0c, 32'h42b14de5, 32'h42c1655f, 32'h4206c5ea, 32'hc23689c5, 32'hc2a645d0};
test_output[8444] = '{32'h42c1655f};
test_index[8444] = '{4};
test_input[67560:67567] = '{32'h42b56fd6, 32'hc0f7c789, 32'h429f6bab, 32'h428de667, 32'h41617497, 32'h40a0e0df, 32'h41b1b4b9, 32'hc25d8ff8};
test_output[8445] = '{32'h42b56fd6};
test_index[8445] = '{0};
test_input[67568:67575] = '{32'hc2bbf3cb, 32'hc20f514b, 32'hc2062fe2, 32'h42a88c25, 32'h423901ff, 32'h426fd333, 32'h429418e6, 32'h42566e2c};
test_output[8446] = '{32'h42a88c25};
test_index[8446] = '{3};
test_input[67576:67583] = '{32'h42bfa7d5, 32'hc28e0560, 32'hc22b06c4, 32'h421e7658, 32'h42c01646, 32'hc27c4a6d, 32'h425e8256, 32'h42428f49};
test_output[8447] = '{32'h42c01646};
test_index[8447] = '{4};
test_input[67584:67591] = '{32'h4241c969, 32'h42ad99be, 32'hc22c1c8a, 32'hc2a1e867, 32'hc17cb362, 32'h419f7926, 32'hbfdd9705, 32'hc2c152c8};
test_output[8448] = '{32'h42ad99be};
test_index[8448] = '{1};
test_input[67592:67599] = '{32'h42894dd0, 32'h41c6976d, 32'hc1594a3f, 32'h4228d403, 32'h42ba6894, 32'h422a8925, 32'h41b0011e, 32'hc261dbed};
test_output[8449] = '{32'h42ba6894};
test_index[8449] = '{4};
test_input[67600:67607] = '{32'h42b6ed29, 32'hc24eb513, 32'hc263bf67, 32'h42955a5a, 32'h416ad546, 32'hc28dce18, 32'hc2105c40, 32'hc14ad61b};
test_output[8450] = '{32'h42b6ed29};
test_index[8450] = '{0};
test_input[67608:67615] = '{32'h4203a070, 32'hc2635492, 32'h42a3cceb, 32'h42b926ee, 32'h4290359d, 32'hc1ef46ee, 32'hbfb0ac37, 32'hc29253bc};
test_output[8451] = '{32'h42b926ee};
test_index[8451] = '{3};
test_input[67616:67623] = '{32'hc27d619f, 32'hc237c016, 32'h3e77c953, 32'h428a588b, 32'h413908e6, 32'hc1d35664, 32'h4234d69a, 32'h42329404};
test_output[8452] = '{32'h428a588b};
test_index[8452] = '{3};
test_input[67624:67631] = '{32'hc2a2dab8, 32'h42c75e4b, 32'hc1793644, 32'h4273222f, 32'hc2c56c42, 32'hc1a66148, 32'hc24b3599, 32'h4227a73d};
test_output[8453] = '{32'h42c75e4b};
test_index[8453] = '{1};
test_input[67632:67639] = '{32'hc240ea34, 32'hc2549527, 32'h424fc4a6, 32'hc2810fa2, 32'hc273b087, 32'hc11878a9, 32'hc27c7dd5, 32'h41c41a17};
test_output[8454] = '{32'h424fc4a6};
test_index[8454] = '{2};
test_input[67640:67647] = '{32'h423304b5, 32'hc1f0fa39, 32'h40b151ae, 32'h42a677e9, 32'h414b2337, 32'hc11a8da2, 32'hc2005cc9, 32'hc0b2a0f7};
test_output[8455] = '{32'h42a677e9};
test_index[8455] = '{3};
test_input[67648:67655] = '{32'hc232cb84, 32'h429e13ed, 32'hc29d8e5e, 32'h422ae94f, 32'h42c52110, 32'hc1bc2c2f, 32'hc2b1a6d5, 32'h41c20c5d};
test_output[8456] = '{32'h42c52110};
test_index[8456] = '{4};
test_input[67656:67663] = '{32'h42a73548, 32'h427e1e3d, 32'h4111e752, 32'hc282c1d4, 32'h420b79c4, 32'h42b1a155, 32'hc24190d1, 32'hc20a3582};
test_output[8457] = '{32'h42b1a155};
test_index[8457] = '{5};
test_input[67664:67671] = '{32'h428b7006, 32'hc239e84f, 32'h4296588e, 32'hc2571408, 32'hc24c5a16, 32'hc2a7bb2c, 32'h41c1183e, 32'h427e93b9};
test_output[8458] = '{32'h4296588e};
test_index[8458] = '{2};
test_input[67672:67679] = '{32'hbe9c50a4, 32'h42921396, 32'hc2c54dc3, 32'h42132362, 32'h4262b4bf, 32'hc1a675c4, 32'hc2a97ac4, 32'h429ce3d8};
test_output[8459] = '{32'h429ce3d8};
test_index[8459] = '{7};
test_input[67680:67687] = '{32'hc22850b9, 32'h414e5ffe, 32'hc13253bb, 32'h425b20cc, 32'h3f20b7e1, 32'hc2b5b85d, 32'hc27358c5, 32'h425b3911};
test_output[8460] = '{32'h425b3911};
test_index[8460] = '{7};
test_input[67688:67695] = '{32'h42875d5f, 32'hc20455b3, 32'h41d75cba, 32'hc2445c2f, 32'hc1d8a396, 32'h429d3e05, 32'h42971432, 32'hc28f1efb};
test_output[8461] = '{32'h429d3e05};
test_index[8461] = '{5};
test_input[67696:67703] = '{32'hc2713a76, 32'hc29ba00f, 32'h4294ff22, 32'h42a12870, 32'hc2bb697d, 32'h429fc9df, 32'hc29321f7, 32'hc19a2a1b};
test_output[8462] = '{32'h42a12870};
test_index[8462] = '{3};
test_input[67704:67711] = '{32'hc21551f1, 32'h42c7a242, 32'hc1b5b8e4, 32'h42adadc9, 32'h4254c8e5, 32'h42ad26c0, 32'h42b6f443, 32'hc21dc343};
test_output[8463] = '{32'h42c7a242};
test_index[8463] = '{1};
test_input[67712:67719] = '{32'h425846c4, 32'h3ff06c5f, 32'hc1eda644, 32'hc29a0187, 32'h406b27a9, 32'h42755225, 32'hc00c3193, 32'hc28aea57};
test_output[8464] = '{32'h42755225};
test_index[8464] = '{5};
test_input[67720:67727] = '{32'h42c4d15b, 32'hc24b46fc, 32'hc26ce767, 32'h4205fba2, 32'hc267d53f, 32'hc2b1406b, 32'hc05bd786, 32'hc27fba83};
test_output[8465] = '{32'h42c4d15b};
test_index[8465] = '{0};
test_input[67728:67735] = '{32'h42940b41, 32'h414cfd62, 32'h428b5f83, 32'hc2671489, 32'h404b6c62, 32'h424e4dfc, 32'h4200a77a, 32'hc2ab9798};
test_output[8466] = '{32'h42940b41};
test_index[8466] = '{0};
test_input[67736:67743] = '{32'hc07617de, 32'hc1d8b075, 32'h4102cb56, 32'h423cf36c, 32'h428513b7, 32'h424697e6, 32'h429c4a04, 32'hc246996d};
test_output[8467] = '{32'h429c4a04};
test_index[8467] = '{6};
test_input[67744:67751] = '{32'hc10860b7, 32'h40fe7cfa, 32'hc26ca5a7, 32'h414b3290, 32'h419eb774, 32'hc2061ad7, 32'hc2965d7c, 32'hc2280231};
test_output[8468] = '{32'h419eb774};
test_index[8468] = '{4};
test_input[67752:67759] = '{32'hc2554a8f, 32'h4298172d, 32'hc197c121, 32'hc28f3a4c, 32'h40936308, 32'h4139f7ec, 32'hc069e8d2, 32'hc1aeb9ee};
test_output[8469] = '{32'h4298172d};
test_index[8469] = '{1};
test_input[67760:67767] = '{32'h41d3e050, 32'h42150f30, 32'h4195063f, 32'h4250375d, 32'hc280e0fb, 32'h41e1c93a, 32'hc24db689, 32'h42890ba8};
test_output[8470] = '{32'h42890ba8};
test_index[8470] = '{7};
test_input[67768:67775] = '{32'hc2003d7d, 32'h426f7fe1, 32'h42525587, 32'hc282c640, 32'hc2a0a758, 32'hc223bde6, 32'hc0806ede, 32'h421254c0};
test_output[8471] = '{32'h426f7fe1};
test_index[8471] = '{1};
test_input[67776:67783] = '{32'hc2983033, 32'hc23d3720, 32'h40894dbd, 32'h420e7aa0, 32'h41bc7e24, 32'hc2c44857, 32'hc2ad9f0d, 32'h4208b7ea};
test_output[8472] = '{32'h420e7aa0};
test_index[8472] = '{3};
test_input[67784:67791] = '{32'hc1f48880, 32'h42a77200, 32'h40eb55bb, 32'h428d68e4, 32'hc248cc35, 32'hc20a0e23, 32'hc2a72724, 32'hc20d2853};
test_output[8473] = '{32'h42a77200};
test_index[8473] = '{1};
test_input[67792:67799] = '{32'hc27c0065, 32'hc2a77b88, 32'hc2a33203, 32'h42c6631b, 32'h42af37cf, 32'hc28560c7, 32'h427059da, 32'hc22d585a};
test_output[8474] = '{32'h42c6631b};
test_index[8474] = '{3};
test_input[67800:67807] = '{32'hc1ced488, 32'hc2564fcb, 32'h42a0a7cc, 32'h42b65105, 32'h41b25ee7, 32'hc231bcb1, 32'h42b8759d, 32'h40c07b50};
test_output[8475] = '{32'h42b8759d};
test_index[8475] = '{6};
test_input[67808:67815] = '{32'h42778111, 32'hc1c9b67d, 32'h42bf0b0b, 32'h429c4914, 32'h4209fc5a, 32'hc24d7112, 32'hc283ff5f, 32'h4266adc4};
test_output[8476] = '{32'h42bf0b0b};
test_index[8476] = '{2};
test_input[67816:67823] = '{32'h4162653a, 32'hc28dbd34, 32'h421f86dd, 32'hc142b99e, 32'hc27cb3a2, 32'h419aef0f, 32'hc2a292f2, 32'h426ab28e};
test_output[8477] = '{32'h426ab28e};
test_index[8477] = '{7};
test_input[67824:67831] = '{32'hc26b4b54, 32'h429869e6, 32'h42a5594c, 32'hc29ce336, 32'hc18bb8b5, 32'h3ff88826, 32'h428423f8, 32'h41816f07};
test_output[8478] = '{32'h42a5594c};
test_index[8478] = '{2};
test_input[67832:67839] = '{32'hc20d8095, 32'hc152410a, 32'hc26de1ca, 32'h41e36624, 32'hc28d37ef, 32'hc1b0c11c, 32'h4258d02f, 32'h422d0838};
test_output[8479] = '{32'h4258d02f};
test_index[8479] = '{6};
test_input[67840:67847] = '{32'h42c08232, 32'h424b147c, 32'hc288944c, 32'h42966354, 32'hc10e6234, 32'h42a65197, 32'hc2b4a319, 32'h429d2e03};
test_output[8480] = '{32'h42c08232};
test_index[8480] = '{0};
test_input[67848:67855] = '{32'hc1c4238a, 32'h42c7ddca, 32'h42b2da2b, 32'h4211da0e, 32'hc2777b27, 32'h41263ff6, 32'h423d0772, 32'hc2b64916};
test_output[8481] = '{32'h42c7ddca};
test_index[8481] = '{1};
test_input[67856:67863] = '{32'hc2b15f4b, 32'hc291bf85, 32'hc209fd97, 32'h42baee1b, 32'h4054aa33, 32'h42a390a0, 32'h413706e1, 32'h4265ae14};
test_output[8482] = '{32'h42baee1b};
test_index[8482] = '{3};
test_input[67864:67871] = '{32'hc287b3a2, 32'h4259c290, 32'hc291224c, 32'h41dfbb39, 32'h429544cc, 32'hc1dd0274, 32'h4212803b, 32'hc283e83f};
test_output[8483] = '{32'h429544cc};
test_index[8483] = '{4};
test_input[67872:67879] = '{32'hc2bdc5c8, 32'h4094c3f9, 32'hc2c1685b, 32'h4251743c, 32'h406e5250, 32'h4243c741, 32'h420f16bc, 32'hc2bfcbae};
test_output[8484] = '{32'h4251743c};
test_index[8484] = '{3};
test_input[67880:67887] = '{32'h42c0453c, 32'hc1931651, 32'h41fccd54, 32'hc19be95d, 32'hc295d50b, 32'h42c10f0d, 32'h42a1870b, 32'h4208e21e};
test_output[8485] = '{32'h42c10f0d};
test_index[8485] = '{5};
test_input[67888:67895] = '{32'hc008dd90, 32'hc2c52120, 32'h427e82fe, 32'hc1b2c795, 32'h4248e72c, 32'h41fa9f76, 32'h42061c5c, 32'h4134a571};
test_output[8486] = '{32'h427e82fe};
test_index[8486] = '{2};
test_input[67896:67903] = '{32'h42c1b527, 32'h42bce800, 32'h40b4498d, 32'h42a745b8, 32'h42bd01a1, 32'h428f24d5, 32'h413b3a2a, 32'h42bb6bf5};
test_output[8487] = '{32'h42c1b527};
test_index[8487] = '{0};
test_input[67904:67911] = '{32'h42588a66, 32'hc2657a06, 32'hc22e7731, 32'hc006b9ea, 32'h41d913e7, 32'hc2621498, 32'hc2b816c6, 32'hc26acbab};
test_output[8488] = '{32'h42588a66};
test_index[8488] = '{0};
test_input[67912:67919] = '{32'h429ed781, 32'h42a61d44, 32'hc28eea9a, 32'h426c9ddd, 32'h42b8297d, 32'hc1182411, 32'h429b309c, 32'hc2a9a6e6};
test_output[8489] = '{32'h42b8297d};
test_index[8489] = '{4};
test_input[67920:67927] = '{32'h422c2152, 32'h41b6bf19, 32'hc2b8fa87, 32'hc2696be3, 32'hc24d8e0d, 32'hc181e941, 32'h429ff4ac, 32'hc2b0c2f2};
test_output[8490] = '{32'h429ff4ac};
test_index[8490] = '{6};
test_input[67928:67935] = '{32'hc2ba814e, 32'hc1387093, 32'h427d1643, 32'h42b29001, 32'h423a0309, 32'h42417950, 32'hc26933f3, 32'h421b8461};
test_output[8491] = '{32'h42b29001};
test_index[8491] = '{3};
test_input[67936:67943] = '{32'hc2731eb1, 32'hc2c64a09, 32'h42a66229, 32'hc22feb88, 32'h40c60965, 32'h403ef111, 32'h42396ff4, 32'h42a70651};
test_output[8492] = '{32'h42a70651};
test_index[8492] = '{7};
test_input[67944:67951] = '{32'hc14bb471, 32'hc29a3d83, 32'h41d041e1, 32'h420b6a89, 32'hc2ae75b9, 32'hc20a78f0, 32'hbf68f531, 32'hc1856e06};
test_output[8493] = '{32'h420b6a89};
test_index[8493] = '{3};
test_input[67952:67959] = '{32'h429fb3a0, 32'hc180d004, 32'h423931d1, 32'h4218bc69, 32'h4285088d, 32'h41a4c0fb, 32'h427765f4, 32'h426996fb};
test_output[8494] = '{32'h429fb3a0};
test_index[8494] = '{0};
test_input[67960:67967] = '{32'hc278d6f4, 32'hbf71cbc4, 32'h4249cd2a, 32'hc27e7b47, 32'hc26bdbad, 32'hc25ff30b, 32'hc19eafde, 32'hbca1d13e};
test_output[8495] = '{32'h4249cd2a};
test_index[8495] = '{2};
test_input[67968:67975] = '{32'hc28ff355, 32'h425d7883, 32'h41b5aafd, 32'hc26d26bf, 32'hc2af6568, 32'h410dc470, 32'hc196cecd, 32'hc29a2cdf};
test_output[8496] = '{32'h425d7883};
test_index[8496] = '{1};
test_input[67976:67983] = '{32'h4157ef5a, 32'hc25d6cc5, 32'h4194204d, 32'h424fd8e9, 32'h428ebdcc, 32'h41c15b5b, 32'h418ade7c, 32'h4295401f};
test_output[8497] = '{32'h4295401f};
test_index[8497] = '{7};
test_input[67984:67991] = '{32'hc1165ded, 32'h42a9006d, 32'hc2a1abc2, 32'h424e1694, 32'h4259862a, 32'hc19cd1b4, 32'h414da189, 32'hc2b27ab5};
test_output[8498] = '{32'h42a9006d};
test_index[8498] = '{1};
test_input[67992:67999] = '{32'h425fa15a, 32'h42374db6, 32'h4280065c, 32'h425daa3e, 32'hc2b8fd94, 32'h41fb2bf0, 32'hc11b493c, 32'hc243df2a};
test_output[8499] = '{32'h4280065c};
test_index[8499] = '{2};
test_input[68000:68007] = '{32'hc2524dbf, 32'hc08ac1a0, 32'hc153e259, 32'hc2982b14, 32'h429bc780, 32'h4288c1ae, 32'h42ab594d, 32'hc2aeb6c0};
test_output[8500] = '{32'h42ab594d};
test_index[8500] = '{6};
test_input[68008:68015] = '{32'hc2c00715, 32'hc12149e3, 32'h42885b1e, 32'hc1481f93, 32'h4261d467, 32'hc290a927, 32'h41fd84a8, 32'h41f4e3c1};
test_output[8501] = '{32'h42885b1e};
test_index[8501] = '{2};
test_input[68016:68023] = '{32'hc225f73c, 32'h41c3ec03, 32'h42521b0c, 32'hc191f0c9, 32'hc20f18d0, 32'hc0b096ff, 32'hc180ca30, 32'hc197f0ce};
test_output[8502] = '{32'h42521b0c};
test_index[8502] = '{2};
test_input[68024:68031] = '{32'h4166def6, 32'h428c5a36, 32'h42b579e0, 32'hc2924994, 32'h4254be99, 32'hc28d3b6f, 32'hc2b13ed2, 32'h41859bda};
test_output[8503] = '{32'h42b579e0};
test_index[8503] = '{2};
test_input[68032:68039] = '{32'hc2a61550, 32'hc1e5a8c6, 32'hc2766bbb, 32'h41d25a4a, 32'hc23b6097, 32'h4238d6c6, 32'hc214d656, 32'hc14e308d};
test_output[8504] = '{32'h4238d6c6};
test_index[8504] = '{5};
test_input[68040:68047] = '{32'hc249a61f, 32'h42bb877b, 32'h4277e0a1, 32'hc1516498, 32'hc293564c, 32'h42293bf4, 32'h40f96bcb, 32'hc29ff311};
test_output[8505] = '{32'h42bb877b};
test_index[8505] = '{1};
test_input[68048:68055] = '{32'hc18887cf, 32'hc2bda31d, 32'hc12538e0, 32'h42c5d90f, 32'h4278c2f3, 32'h3f37cfd2, 32'hc2400cc9, 32'hc266b29d};
test_output[8506] = '{32'h42c5d90f};
test_index[8506] = '{3};
test_input[68056:68063] = '{32'hc1c270ef, 32'hc1db1a6e, 32'hc2a9986e, 32'hc24f070a, 32'hc226c378, 32'hc2151994, 32'h410d3241, 32'hc0afa5d4};
test_output[8507] = '{32'h410d3241};
test_index[8507] = '{6};
test_input[68064:68071] = '{32'h429d3931, 32'hc183e918, 32'h420c396d, 32'h423fc6b3, 32'h420fd58d, 32'hc2ad231e, 32'hc21aea9b, 32'h42149c62};
test_output[8508] = '{32'h429d3931};
test_index[8508] = '{0};
test_input[68072:68079] = '{32'hc251822a, 32'h425caff3, 32'hc1daf17e, 32'h4146350d, 32'hc1a0a1ef, 32'hc2c3c0a8, 32'hc1c001d9, 32'h42a3dd73};
test_output[8509] = '{32'h42a3dd73};
test_index[8509] = '{7};
test_input[68080:68087] = '{32'hc27b06c5, 32'h425420a1, 32'h423dc1e2, 32'hc1e88d92, 32'hc236206c, 32'hc229a826, 32'hc1a6f2aa, 32'hc187eeee};
test_output[8510] = '{32'h425420a1};
test_index[8510] = '{1};
test_input[68088:68095] = '{32'h40b63408, 32'hc29bfec2, 32'h41cbceef, 32'h414cf5ac, 32'hc2bf82e3, 32'h42984852, 32'hc2c728f8, 32'h429d9bfe};
test_output[8511] = '{32'h429d9bfe};
test_index[8511] = '{7};
test_input[68096:68103] = '{32'h42b078f4, 32'h427c8ebb, 32'h4278acd4, 32'h425be263, 32'h42951811, 32'h41b307e8, 32'h42657a6d, 32'h424f9295};
test_output[8512] = '{32'h42b078f4};
test_index[8512] = '{0};
test_input[68104:68111] = '{32'hc1cbdd80, 32'h42c35416, 32'h4218bc5f, 32'hc1f7df7b, 32'h4289e480, 32'hc1b0b523, 32'hc084f15a, 32'hc1f046b9};
test_output[8513] = '{32'h42c35416};
test_index[8513] = '{1};
test_input[68112:68119] = '{32'hc278d757, 32'hc273be5c, 32'h418825b1, 32'hc248bfa1, 32'hc273f60d, 32'hc2482c11, 32'hc1828a01, 32'h423fc547};
test_output[8514] = '{32'h423fc547};
test_index[8514] = '{7};
test_input[68120:68127] = '{32'h428a543a, 32'h40c379ea, 32'h420b6e44, 32'h41dd1f17, 32'hc1bc6440, 32'hc2436867, 32'h418c7f22, 32'h41d401cf};
test_output[8515] = '{32'h428a543a};
test_index[8515] = '{0};
test_input[68128:68135] = '{32'hc1c7f0bc, 32'h4131df50, 32'hc20b759d, 32'hc2a85300, 32'h4245b04e, 32'h429f58d5, 32'h429fd758, 32'hc1d9c544};
test_output[8516] = '{32'h429fd758};
test_index[8516] = '{6};
test_input[68136:68143] = '{32'hc28720bb, 32'h42a9208a, 32'hc227f332, 32'hc08996ba, 32'h429eb5b5, 32'h429956ef, 32'h3fa6c200, 32'h42bddfba};
test_output[8517] = '{32'h42bddfba};
test_index[8517] = '{7};
test_input[68144:68151] = '{32'hc281de62, 32'h4225d1e2, 32'h4209f31d, 32'hc2538345, 32'hc074402d, 32'hc266a794, 32'hc1dcdc3b, 32'h41756fe0};
test_output[8518] = '{32'h4225d1e2};
test_index[8518] = '{1};
test_input[68152:68159] = '{32'hc21b98e0, 32'hc1cbea89, 32'h4297cb31, 32'h4236b626, 32'hc1403e5c, 32'h426a9371, 32'hc260b4b2, 32'hc29146ec};
test_output[8519] = '{32'h4297cb31};
test_index[8519] = '{2};
test_input[68160:68167] = '{32'h42333c61, 32'hc2a109c1, 32'hc24c28fa, 32'hc2865054, 32'hc1997006, 32'h41961fdb, 32'h41238175, 32'hc28ede91};
test_output[8520] = '{32'h42333c61};
test_index[8520] = '{0};
test_input[68168:68175] = '{32'h42b0e027, 32'h421f55e5, 32'hc1e059d3, 32'h40e05234, 32'h429da132, 32'h426a3039, 32'h42b0070a, 32'hc198754e};
test_output[8521] = '{32'h42b0e027};
test_index[8521] = '{0};
test_input[68176:68183] = '{32'h427bfce4, 32'h4265307a, 32'h426fb3cc, 32'hc116f551, 32'h41566177, 32'hc2c42be5, 32'hc29366e8, 32'h42c4e7e0};
test_output[8522] = '{32'h42c4e7e0};
test_index[8522] = '{7};
test_input[68184:68191] = '{32'hc29c3b89, 32'hc0d04d69, 32'h421ac9e2, 32'h41aa6252, 32'h42484492, 32'hc22ee903, 32'h4209efe5, 32'h42aeeb63};
test_output[8523] = '{32'h42aeeb63};
test_index[8523] = '{7};
test_input[68192:68199] = '{32'h42043d1e, 32'h428e3711, 32'hc2bfd1f3, 32'hc1e77364, 32'hc2957f4e, 32'hc2215fc7, 32'hc2b07adf, 32'hc2c45dfc};
test_output[8524] = '{32'h428e3711};
test_index[8524] = '{1};
test_input[68200:68207] = '{32'hc18e2c58, 32'hc2861806, 32'hc29a9a25, 32'hc1f39a03, 32'h4245a564, 32'h42b8b019, 32'h4267ccdc, 32'hc2468686};
test_output[8525] = '{32'h42b8b019};
test_index[8525] = '{5};
test_input[68208:68215] = '{32'h41dd1867, 32'h4060322c, 32'hc2a31fa4, 32'hc21d71f4, 32'hc24c27ac, 32'h411d37a4, 32'hc2883e4a, 32'hc2b4058c};
test_output[8526] = '{32'h41dd1867};
test_index[8526] = '{0};
test_input[68216:68223] = '{32'hc1900374, 32'h42127bdb, 32'h4221d14c, 32'hc2bed2df, 32'hc20e8739, 32'h4286ceb0, 32'h41942c45, 32'h42ac2622};
test_output[8527] = '{32'h42ac2622};
test_index[8527] = '{7};
test_input[68224:68231] = '{32'hc1253904, 32'h41e6139d, 32'h42003da9, 32'h42b55526, 32'h405a8aa3, 32'h4211ddaa, 32'hc2bf1372, 32'hc28961b8};
test_output[8528] = '{32'h42b55526};
test_index[8528] = '{3};
test_input[68232:68239] = '{32'hc28ce1fa, 32'h41a1b274, 32'h41685953, 32'h422dd0f0, 32'h422b727f, 32'h4243e468, 32'hc1e3064e, 32'hc23ee91d};
test_output[8529] = '{32'h4243e468};
test_index[8529] = '{5};
test_input[68240:68247] = '{32'hc29ea4b6, 32'h42a93fcb, 32'h42a6c19f, 32'hc289042e, 32'h40816c12, 32'h427b3bda, 32'hc089b078, 32'hc12f1323};
test_output[8530] = '{32'h42a93fcb};
test_index[8530] = '{1};
test_input[68248:68255] = '{32'h41a1a69c, 32'h4068fcd5, 32'hc2585455, 32'h3f2537ab, 32'hc22e7e7a, 32'h42060f00, 32'hc22b5a34, 32'hc2a799e3};
test_output[8531] = '{32'h42060f00};
test_index[8531] = '{5};
test_input[68256:68263] = '{32'h4287fda3, 32'h428c6a64, 32'hc2c71404, 32'hc0a00116, 32'h4097345d, 32'h4289ef37, 32'hc2af6dc4, 32'h428d1127};
test_output[8532] = '{32'h428d1127};
test_index[8532] = '{7};
test_input[68264:68271] = '{32'hc11e971b, 32'hc2ace8df, 32'hc2bfc2a9, 32'hc286438c, 32'hc1030dff, 32'hc2c3d259, 32'h417b30d5, 32'h3f0b294a};
test_output[8533] = '{32'h417b30d5};
test_index[8533] = '{6};
test_input[68272:68279] = '{32'h4151215b, 32'hc2a3dd54, 32'h419245b6, 32'hc1a7afe3, 32'hc2a2f4c3, 32'hc2af35a7, 32'h4230e690, 32'h42b30eb5};
test_output[8534] = '{32'h42b30eb5};
test_index[8534] = '{7};
test_input[68280:68287] = '{32'h41882f0d, 32'h42666836, 32'hc1848da0, 32'hc25542fc, 32'hc286b097, 32'hc2c76ec3, 32'h429e5414, 32'hc2a4a9ec};
test_output[8535] = '{32'h429e5414};
test_index[8535] = '{6};
test_input[68288:68295] = '{32'h42960b67, 32'hc18c13c4, 32'h421293bc, 32'hc0431d66, 32'h42461ebe, 32'hc28a3777, 32'h401d509d, 32'hc255ba21};
test_output[8536] = '{32'h42960b67};
test_index[8536] = '{0};
test_input[68296:68303] = '{32'hc21bc586, 32'hc2bfad1b, 32'hc0d74a2d, 32'hc13fa46e, 32'h428541b3, 32'hc2ba956e, 32'h423be55f, 32'hc15ae7c7};
test_output[8537] = '{32'h428541b3};
test_index[8537] = '{4};
test_input[68304:68311] = '{32'hc2616f67, 32'hc20ec0f7, 32'h4224f14b, 32'hc233c7f2, 32'h42b4e645, 32'hc1815505, 32'h4259cb31, 32'hc2be5262};
test_output[8538] = '{32'h42b4e645};
test_index[8538] = '{4};
test_input[68312:68319] = '{32'hc2b3c151, 32'hc15bf13d, 32'h41ceed76, 32'hbf98400e, 32'h4278a626, 32'h42531760, 32'hc2c36716, 32'hc23a7fc6};
test_output[8539] = '{32'h4278a626};
test_index[8539] = '{4};
test_input[68320:68327] = '{32'h42b818c6, 32'h41d40094, 32'h42a4f842, 32'h40f482dd, 32'h42a438f1, 32'h4287b910, 32'h41fd082e, 32'h4114b333};
test_output[8540] = '{32'h42b818c6};
test_index[8540] = '{0};
test_input[68328:68335] = '{32'hc202d5cc, 32'hc14e86fa, 32'hbf2367d0, 32'h420d8371, 32'h41aafbf3, 32'hc27d1c29, 32'hc2c78bf1, 32'h42a861a8};
test_output[8541] = '{32'h42a861a8};
test_index[8541] = '{7};
test_input[68336:68343] = '{32'hc29d6462, 32'h42a796fd, 32'hc197bc2c, 32'hc25e7bfe, 32'hc296d675, 32'hc121995d, 32'h422ae33f, 32'h42c22908};
test_output[8542] = '{32'h42c22908};
test_index[8542] = '{7};
test_input[68344:68351] = '{32'hc1b3c73b, 32'h4200b013, 32'hc27308ce, 32'hc25b9ae9, 32'h40205507, 32'hc2bf9cb2, 32'hc2b0b789, 32'hc187b94b};
test_output[8543] = '{32'h4200b013};
test_index[8543] = '{1};
test_input[68352:68359] = '{32'h425a3066, 32'hc205c88a, 32'hc26f9925, 32'h4162f8ff, 32'hc20718b8, 32'hc2bbd3ff, 32'hc22eb0c8, 32'h429b1f4a};
test_output[8544] = '{32'h429b1f4a};
test_index[8544] = '{7};
test_input[68360:68367] = '{32'h4281ac08, 32'h4249f4df, 32'hc27ba548, 32'h428947e5, 32'h424860c2, 32'h4265985f, 32'hc2841c52, 32'h41b2d032};
test_output[8545] = '{32'h428947e5};
test_index[8545] = '{3};
test_input[68368:68375] = '{32'hc29de8aa, 32'hc2218ac5, 32'hc141d58b, 32'hc25fab25, 32'h427aeef2, 32'h41a5def5, 32'h42953700, 32'h42b7b49d};
test_output[8546] = '{32'h42b7b49d};
test_index[8546] = '{7};
test_input[68376:68383] = '{32'hc28fa9db, 32'h4173e7aa, 32'hc273006c, 32'h428f4454, 32'h41fcf368, 32'h41df4f0c, 32'h426d9b00, 32'hc27ed159};
test_output[8547] = '{32'h428f4454};
test_index[8547] = '{3};
test_input[68384:68391] = '{32'h4127d0bf, 32'hc1c7e4fd, 32'h4258d51e, 32'h40e83ab6, 32'hc2c542cd, 32'hc2a9e6c9, 32'hc2564e95, 32'hc29ccc13};
test_output[8548] = '{32'h4258d51e};
test_index[8548] = '{2};
test_input[68392:68399] = '{32'h418ae082, 32'hc26bc047, 32'h42977596, 32'h414907e0, 32'h41ef75e2, 32'h41bbd9ba, 32'h41ab362c, 32'h3fe19713};
test_output[8549] = '{32'h42977596};
test_index[8549] = '{2};
test_input[68400:68407] = '{32'hc131d4ee, 32'h42254aa9, 32'h42a6bba4, 32'h42c469df, 32'h420c7ef8, 32'h4268637f, 32'hc1d90f76, 32'h42a7f00b};
test_output[8550] = '{32'h42c469df};
test_index[8550] = '{3};
test_input[68408:68415] = '{32'h41e8ed47, 32'h3f4a13a2, 32'h42bcf3da, 32'h42543c41, 32'hc1ea9dd7, 32'h40f6b34e, 32'hc29bfe45, 32'hc2780b07};
test_output[8551] = '{32'h42bcf3da};
test_index[8551] = '{2};
test_input[68416:68423] = '{32'h40c03eb7, 32'hc2bb1310, 32'h42b2b585, 32'h4296c034, 32'hc188516c, 32'h42386aad, 32'hc240da71, 32'hc18baa79};
test_output[8552] = '{32'h42b2b585};
test_index[8552] = '{2};
test_input[68424:68431] = '{32'hc2b53f35, 32'h429dd793, 32'hc0dcd24e, 32'hc2b5d127, 32'hc229ba56, 32'hc2c214ad, 32'hc29c3ddb, 32'hc26be231};
test_output[8553] = '{32'h429dd793};
test_index[8553] = '{1};
test_input[68432:68439] = '{32'hc211d16b, 32'hc29b2b56, 32'hc2873e56, 32'hc1bbbdd4, 32'h41ddfa78, 32'h42217bfc, 32'hc22eb572, 32'hc29823c3};
test_output[8554] = '{32'h42217bfc};
test_index[8554] = '{5};
test_input[68440:68447] = '{32'hc2ac2536, 32'hc181b9b3, 32'hc244d801, 32'hc20d2194, 32'hc2a0d0a8, 32'h41f42262, 32'h42115c0c, 32'hc2a772ec};
test_output[8555] = '{32'h42115c0c};
test_index[8555] = '{6};
test_input[68448:68455] = '{32'hc04c994b, 32'h425eca68, 32'h424a8a60, 32'h4294d943, 32'h42976490, 32'hc2b141c8, 32'h427f8744, 32'hc1082444};
test_output[8556] = '{32'h42976490};
test_index[8556] = '{4};
test_input[68456:68463] = '{32'h42a45c01, 32'hc2427b12, 32'hc22bd24a, 32'h42b0c863, 32'hc2463289, 32'h42b9510a, 32'h42be5a68, 32'h41dc89e0};
test_output[8557] = '{32'h42be5a68};
test_index[8557] = '{6};
test_input[68464:68471] = '{32'hc1dd9f39, 32'h41093f32, 32'h42a7f94e, 32'hc229d7de, 32'hc24c465d, 32'hc1eb8b25, 32'hc2ac99b3, 32'h41e402ef};
test_output[8558] = '{32'h42a7f94e};
test_index[8558] = '{2};
test_input[68472:68479] = '{32'h4251ab18, 32'h4231e873, 32'hc2bbcde3, 32'h41451abe, 32'h411d7322, 32'h42960b93, 32'h42460fab, 32'hc2891115};
test_output[8559] = '{32'h42960b93};
test_index[8559] = '{5};
test_input[68480:68487] = '{32'hc1ade322, 32'hc299dd9a, 32'h41d98dbb, 32'h423982b7, 32'h41a5bba3, 32'hc16b4f69, 32'h420c8f5d, 32'hc10354ad};
test_output[8560] = '{32'h423982b7};
test_index[8560] = '{3};
test_input[68488:68495] = '{32'hc23e5862, 32'hc2b1dd60, 32'h41fe8a33, 32'h3fa052ad, 32'h42ad13d9, 32'hc2bbf493, 32'h42380ed8, 32'h4099de2a};
test_output[8561] = '{32'h42ad13d9};
test_index[8561] = '{4};
test_input[68496:68503] = '{32'hc2b15e19, 32'hc259d639, 32'hc24ddbce, 32'h42a864dc, 32'hc28e3faa, 32'hc2404809, 32'h40fee0ba, 32'h41e5cb32};
test_output[8562] = '{32'h42a864dc};
test_index[8562] = '{3};
test_input[68504:68511] = '{32'h426cd2bb, 32'hc2080aba, 32'hc2139a95, 32'hc29694f7, 32'h42a4773b, 32'h42961669, 32'h42c1bc67, 32'hc281b58f};
test_output[8563] = '{32'h42c1bc67};
test_index[8563] = '{6};
test_input[68512:68519] = '{32'hc2304912, 32'hc23158b9, 32'h42bb5c2c, 32'h421327d4, 32'h424c9f7d, 32'hc2902094, 32'h42ac09e6, 32'h4297cf31};
test_output[8564] = '{32'h42bb5c2c};
test_index[8564] = '{2};
test_input[68520:68527] = '{32'h42bb0976, 32'h4240ce4a, 32'h42079239, 32'hc2351973, 32'h42aa9144, 32'hc206bab5, 32'h417b5193, 32'h423216c5};
test_output[8565] = '{32'h42bb0976};
test_index[8565] = '{0};
test_input[68528:68535] = '{32'h42630378, 32'hc2a64c0f, 32'h42acb023, 32'hc2949b07, 32'h42996af1, 32'hc28e851b, 32'h4167409d, 32'h42871258};
test_output[8566] = '{32'h42acb023};
test_index[8566] = '{2};
test_input[68536:68543] = '{32'hc1a253c7, 32'h4210eac1, 32'h420f5d6b, 32'h4171cf54, 32'hc2518eb2, 32'hc2914c42, 32'h42414981, 32'hc2469897};
test_output[8567] = '{32'h42414981};
test_index[8567] = '{6};
test_input[68544:68551] = '{32'h415542f2, 32'hc286e3d1, 32'h42b3eea9, 32'h42458683, 32'hc20e3d38, 32'hc2900632, 32'h42c163d1, 32'hc2a72572};
test_output[8568] = '{32'h42c163d1};
test_index[8568] = '{6};
test_input[68552:68559] = '{32'hc219eaec, 32'h4229f5b6, 32'hc267e8c5, 32'h42b78630, 32'hc2c38e5d, 32'h41040a06, 32'h4126ac4a, 32'h422e8750};
test_output[8569] = '{32'h42b78630};
test_index[8569] = '{3};
test_input[68560:68567] = '{32'h42b42e3d, 32'h42b94dbf, 32'h41896372, 32'hc243d375, 32'hc2912b54, 32'hc27de9ce, 32'h4076dc35, 32'hc21c8b53};
test_output[8570] = '{32'h42b94dbf};
test_index[8570] = '{1};
test_input[68568:68575] = '{32'hc2b7c5d7, 32'hc13602e3, 32'hc1743a7d, 32'hc1ef7eef, 32'hc2bb7b0b, 32'hc245ebfa, 32'hc1aca988, 32'hc23a2afa};
test_output[8571] = '{32'hc13602e3};
test_index[8571] = '{1};
test_input[68576:68583] = '{32'hc2a8b1f0, 32'h41c098bb, 32'h42351bfd, 32'h42b1b7e0, 32'hc1cae194, 32'h4207540a, 32'h41f9880b, 32'hc2028fcc};
test_output[8572] = '{32'h42b1b7e0};
test_index[8572] = '{3};
test_input[68584:68591] = '{32'hc2a3b670, 32'hc189a293, 32'hc289844c, 32'hc28c56b0, 32'h42a8c1ae, 32'h41dd859e, 32'h426353be, 32'hc2bdc7db};
test_output[8573] = '{32'h42a8c1ae};
test_index[8573] = '{4};
test_input[68592:68599] = '{32'h42a72587, 32'hc06375f2, 32'h42adab80, 32'h42c1f018, 32'h419600b4, 32'hc2b099c6, 32'h42a63cb5, 32'h42a2a966};
test_output[8574] = '{32'h42c1f018};
test_index[8574] = '{3};
test_input[68600:68607] = '{32'hc044c583, 32'h421d94dd, 32'hc15753a6, 32'h428c039f, 32'hc2a1cf96, 32'h42121c6e, 32'h4202c4a7, 32'h42546196};
test_output[8575] = '{32'h428c039f};
test_index[8575] = '{3};
test_input[68608:68615] = '{32'h42851778, 32'h4262975b, 32'h429a32a9, 32'hc274a3dd, 32'hc2ad1cfa, 32'h4023cca8, 32'h422c2eb4, 32'h4249aeb1};
test_output[8576] = '{32'h429a32a9};
test_index[8576] = '{2};
test_input[68616:68623] = '{32'h41cf7d24, 32'hc18d2499, 32'hc2bf4623, 32'h429ba6bb, 32'hc2498929, 32'h421c0f4e, 32'h42711d3b, 32'hc1f7d625};
test_output[8577] = '{32'h429ba6bb};
test_index[8577] = '{3};
test_input[68624:68631] = '{32'h4222ae51, 32'h41c0c3d4, 32'hc28afd12, 32'hc16e76ef, 32'hc2120e82, 32'h42062ba1, 32'h41b4511b, 32'h4003551d};
test_output[8578] = '{32'h4222ae51};
test_index[8578] = '{0};
test_input[68632:68639] = '{32'h42a20605, 32'h42b7b920, 32'hc25dd8d7, 32'h42113694, 32'hc0a15040, 32'hc21fc474, 32'hc2a1d283, 32'h41c8512b};
test_output[8579] = '{32'h42b7b920};
test_index[8579] = '{1};
test_input[68640:68647] = '{32'h42b49055, 32'h41e891cb, 32'h42598a79, 32'hc21d575f, 32'h41aaf888, 32'h4193013f, 32'hc1890891, 32'hbfb36506};
test_output[8580] = '{32'h42b49055};
test_index[8580] = '{0};
test_input[68648:68655] = '{32'hc275c1b4, 32'h41573c17, 32'h4283e0d6, 32'h42a8968a, 32'hc2924c3c, 32'hbff1a878, 32'hc2c74e0c, 32'h419a4b5f};
test_output[8581] = '{32'h42a8968a};
test_index[8581] = '{3};
test_input[68656:68663] = '{32'h42641a46, 32'hc1dd2d3f, 32'hc2ad7bcc, 32'h41a9d0f3, 32'h4233cfb4, 32'hc08cf219, 32'hc116e6a9, 32'hc2a3f272};
test_output[8582] = '{32'h42641a46};
test_index[8582] = '{0};
test_input[68664:68671] = '{32'h42386770, 32'hc2c2e9e8, 32'h41715d3a, 32'hc274e510, 32'h42a86e37, 32'hc19ce806, 32'hc290ca0d, 32'hc09e1c6d};
test_output[8583] = '{32'h42a86e37};
test_index[8583] = '{4};
test_input[68672:68679] = '{32'hc2837e3d, 32'h4290d7b7, 32'h429931b6, 32'hc2a1a70f, 32'h4275b022, 32'hc25a9a18, 32'h42b0a4ca, 32'hc299d288};
test_output[8584] = '{32'h42b0a4ca};
test_index[8584] = '{6};
test_input[68680:68687] = '{32'hc28e4299, 32'hc1959b49, 32'h41ad65dc, 32'hc2576aee, 32'h41fb3ccd, 32'hc13d3a3b, 32'hc26feeb6, 32'h4252ff2e};
test_output[8585] = '{32'h4252ff2e};
test_index[8585] = '{7};
test_input[68688:68695] = '{32'h42a696bf, 32'h42712860, 32'h410bbf96, 32'h42af7103, 32'hc16a7901, 32'h400831fb, 32'hc2878e89, 32'hc211b199};
test_output[8586] = '{32'h42af7103};
test_index[8586] = '{3};
test_input[68696:68703] = '{32'hc1841708, 32'h42970e56, 32'hc22e128f, 32'hc26145a1, 32'hc22e256d, 32'h428779bd, 32'h41f2fd62, 32'h428b2430};
test_output[8587] = '{32'h42970e56};
test_index[8587] = '{1};
test_input[68704:68711] = '{32'h427e176b, 32'h42a18801, 32'hc2121fca, 32'h425ff7b0, 32'h426fde27, 32'hc11ca259, 32'hc2a01bed, 32'hc1946b76};
test_output[8588] = '{32'h42a18801};
test_index[8588] = '{1};
test_input[68712:68719] = '{32'h41aa760f, 32'hc2ba6e95, 32'h41cd6d25, 32'h42a10cc7, 32'hc1d71c1e, 32'h42466f4d, 32'h42818e91, 32'h411d725b};
test_output[8589] = '{32'h42a10cc7};
test_index[8589] = '{3};
test_input[68720:68727] = '{32'hc281a638, 32'hc1294ab9, 32'hc14801c3, 32'h42c27170, 32'h413bd601, 32'h41ae68c5, 32'hc191bb0c, 32'h41938e4b};
test_output[8590] = '{32'h42c27170};
test_index[8590] = '{3};
test_input[68728:68735] = '{32'hc2babd22, 32'hc2c7e4ff, 32'hc2a4047a, 32'h42657d7c, 32'h42c6cdcb, 32'h422f0a60, 32'h42265888, 32'h42bf5aaa};
test_output[8591] = '{32'h42c6cdcb};
test_index[8591] = '{4};
test_input[68736:68743] = '{32'hc2ae1721, 32'hc16db596, 32'h42b5bdbe, 32'h42a19590, 32'h41ae0968, 32'h42142df2, 32'h41a5ed0e, 32'hc1ce1313};
test_output[8592] = '{32'h42b5bdbe};
test_index[8592] = '{2};
test_input[68744:68751] = '{32'hc28cf05c, 32'h42bbf5fd, 32'hc2ba8327, 32'h41967062, 32'h4279e2ed, 32'hc21372ea, 32'h42b531f2, 32'h42363bea};
test_output[8593] = '{32'h42bbf5fd};
test_index[8593] = '{1};
test_input[68752:68759] = '{32'hc16b2452, 32'hc2934b78, 32'hc2bd376e, 32'hc016e3e2, 32'hc2425875, 32'hc2a46942, 32'hc1b20acf, 32'hbf784b21};
test_output[8594] = '{32'hbf784b21};
test_index[8594] = '{7};
test_input[68760:68767] = '{32'h41181e0c, 32'h42930563, 32'h423a4fca, 32'h418f8119, 32'hc26119dc, 32'h41167458, 32'h42863d3a, 32'hc1296213};
test_output[8595] = '{32'h42930563};
test_index[8595] = '{1};
test_input[68768:68775] = '{32'hc2751adf, 32'hc2884393, 32'h425ec603, 32'h41f13b75, 32'h4216d748, 32'h42b1337b, 32'h41be8ffd, 32'h422da5e7};
test_output[8596] = '{32'h42b1337b};
test_index[8596] = '{5};
test_input[68776:68783] = '{32'h42a93bf9, 32'h4283b766, 32'hc171cc5a, 32'h41914066, 32'hc128497a, 32'h411321a1, 32'h42266866, 32'h42bcf94a};
test_output[8597] = '{32'h42bcf94a};
test_index[8597] = '{7};
test_input[68784:68791] = '{32'hc2821856, 32'hc0801701, 32'h420db487, 32'h425b36c6, 32'hc2bd25c8, 32'hc29b9f7d, 32'hc255c76e, 32'h40b07710};
test_output[8598] = '{32'h425b36c6};
test_index[8598] = '{3};
test_input[68792:68799] = '{32'hc238ee05, 32'hc19a6f1f, 32'h42af8c03, 32'hc207e49a, 32'h429e1e0e, 32'h42b9d959, 32'h4270f2cd, 32'h409ecf98};
test_output[8599] = '{32'h42b9d959};
test_index[8599] = '{5};
test_input[68800:68807] = '{32'hc2011bc6, 32'h412f7ccd, 32'hc2835b5b, 32'h429567f6, 32'h42a05ce7, 32'h4290654e, 32'hc1fde1d3, 32'h428d6be6};
test_output[8600] = '{32'h42a05ce7};
test_index[8600] = '{4};
test_input[68808:68815] = '{32'h412692a5, 32'hc24c30ed, 32'h41a5a8f0, 32'h42c07921, 32'hc22482f8, 32'hc2ba35cc, 32'h42a7642d, 32'h41aa1749};
test_output[8601] = '{32'h42c07921};
test_index[8601] = '{3};
test_input[68816:68823] = '{32'h4217d148, 32'h421a5379, 32'hc28f504c, 32'h42770bd7, 32'hc28ad50e, 32'h42c256a5, 32'hc217bd5a, 32'h41d6e106};
test_output[8602] = '{32'h42c256a5};
test_index[8602] = '{5};
test_input[68824:68831] = '{32'h41d2d8fa, 32'hc1bd529c, 32'h42a16c12, 32'h418ef458, 32'h41c1edc5, 32'hc1d43968, 32'hc29e1733, 32'hc1494671};
test_output[8603] = '{32'h42a16c12};
test_index[8603] = '{2};
test_input[68832:68839] = '{32'h3f584351, 32'hc18e617a, 32'h41ffabc3, 32'h408ee7eb, 32'h3d98bf6c, 32'hc28879e2, 32'hc23818b6, 32'hc1c408c4};
test_output[8604] = '{32'h41ffabc3};
test_index[8604] = '{2};
test_input[68840:68847] = '{32'hc1e670d3, 32'hc214b880, 32'h4080ab69, 32'hc2999d49, 32'h42adb8d9, 32'h42887624, 32'h414ceea5, 32'h423f0040};
test_output[8605] = '{32'h42adb8d9};
test_index[8605] = '{4};
test_input[68848:68855] = '{32'hc235edc9, 32'hc294be99, 32'h416229e0, 32'hc2ab721d, 32'hc194d980, 32'hc227bd41, 32'hc0254eb8, 32'hc28007cd};
test_output[8606] = '{32'h416229e0};
test_index[8606] = '{2};
test_input[68856:68863] = '{32'hc28efab3, 32'hc2a2242f, 32'hc2a60e23, 32'h4281f6dd, 32'hc285d27d, 32'h4168519a, 32'hc28e8a2e, 32'hc29b0837};
test_output[8607] = '{32'h4281f6dd};
test_index[8607] = '{3};
test_input[68864:68871] = '{32'hc1e1b3e3, 32'hc29f11b3, 32'h4284891a, 32'hc29a5438, 32'hc27b86c0, 32'h41e21d7d, 32'h42b19f4e, 32'hc0944299};
test_output[8608] = '{32'h42b19f4e};
test_index[8608] = '{6};
test_input[68872:68879] = '{32'h41e7458b, 32'h3ef15b21, 32'h41e36b87, 32'hc2c4b22f, 32'h4218c326, 32'h4075497f, 32'h41b7b420, 32'h42507833};
test_output[8609] = '{32'h42507833};
test_index[8609] = '{7};
test_input[68880:68887] = '{32'hc2019bfb, 32'h42a66d3c, 32'h429d1938, 32'h42bb267a, 32'hc1aa1930, 32'h413dd735, 32'h42c7120e, 32'h41b12448};
test_output[8610] = '{32'h42c7120e};
test_index[8610] = '{6};
test_input[68888:68895] = '{32'hc288ece5, 32'h4298d4c4, 32'hc21be02f, 32'hc19f49bb, 32'h4287c1b2, 32'h4287284a, 32'hc240c714, 32'h41dd9052};
test_output[8611] = '{32'h4298d4c4};
test_index[8611] = '{1};
test_input[68896:68903] = '{32'hc2bdf5e6, 32'h4288471d, 32'hc2c4cd74, 32'h42308f51, 32'hc2a7554e, 32'h4244373c, 32'h41fa9030, 32'h429ab4b9};
test_output[8612] = '{32'h429ab4b9};
test_index[8612] = '{7};
test_input[68904:68911] = '{32'hc28ba64d, 32'hc25b20c2, 32'h425a88f3, 32'hc18a4c8c, 32'h421c5c68, 32'hc25324a3, 32'hc24893d1, 32'h422a9c44};
test_output[8613] = '{32'h425a88f3};
test_index[8613] = '{2};
test_input[68912:68919] = '{32'hbf8dc38e, 32'h420e7497, 32'hc28e6225, 32'h42674f25, 32'h4225c969, 32'h4295e260, 32'h40f52c50, 32'h420e693d};
test_output[8614] = '{32'h4295e260};
test_index[8614] = '{5};
test_input[68920:68927] = '{32'hc1fa0188, 32'h422077ef, 32'h42a056be, 32'hc1ecbe93, 32'h4221ce43, 32'hc0ca6126, 32'hc2bf6c96, 32'h42c475c7};
test_output[8615] = '{32'h42c475c7};
test_index[8615] = '{7};
test_input[68928:68935] = '{32'hc28c843b, 32'h428d1abe, 32'hc201be8b, 32'h42c620ba, 32'hc0540dfc, 32'h4234455a, 32'h423b19de, 32'h41f93211};
test_output[8616] = '{32'h42c620ba};
test_index[8616] = '{3};
test_input[68936:68943] = '{32'h3f97e99c, 32'hc26aa39d, 32'hc2784943, 32'h428e7657, 32'h42c740d3, 32'h4226be09, 32'h4260e10a, 32'h428524f7};
test_output[8617] = '{32'h42c740d3};
test_index[8617] = '{4};
test_input[68944:68951] = '{32'hc22e0d7f, 32'h428ce4be, 32'hc200e560, 32'hc20d6639, 32'hc2c58d08, 32'h4136e18b, 32'h426b6ffb, 32'h42298443};
test_output[8618] = '{32'h428ce4be};
test_index[8618] = '{1};
test_input[68952:68959] = '{32'h422e3c33, 32'h427a65d2, 32'hc1114816, 32'h42a5681e, 32'h40703999, 32'h42abd386, 32'hc29f3fdb, 32'h4181ca04};
test_output[8619] = '{32'h42abd386};
test_index[8619] = '{5};
test_input[68960:68967] = '{32'hc2bcd03b, 32'hc247d43e, 32'hc1b7d5da, 32'h41ab3c26, 32'h42ad86c0, 32'h42b6841d, 32'hc29621ce, 32'h424daae1};
test_output[8620] = '{32'h42b6841d};
test_index[8620] = '{5};
test_input[68968:68975] = '{32'hc245a124, 32'h42bcab15, 32'hc298269c, 32'hc2007000, 32'hc1971821, 32'h41a4da29, 32'hc237c63c, 32'h421bf246};
test_output[8621] = '{32'h42bcab15};
test_index[8621] = '{1};
test_input[68976:68983] = '{32'h427c32a5, 32'hc262d985, 32'h4287fe2f, 32'h41b805cc, 32'h41c75c50, 32'hc14d6791, 32'h425af492, 32'hc0161139};
test_output[8622] = '{32'h4287fe2f};
test_index[8622] = '{2};
test_input[68984:68991] = '{32'hc2a1c5fb, 32'hc2990c24, 32'hc2b6cced, 32'h42a67338, 32'hc2bd9002, 32'hc135b813, 32'h42380440, 32'h41fb1c7b};
test_output[8623] = '{32'h42a67338};
test_index[8623] = '{3};
test_input[68992:68999] = '{32'h421faf3e, 32'hc2b60666, 32'h42c34a13, 32'h420e3177, 32'hc2c7828d, 32'h42463f21, 32'hc0c01ec8, 32'hc1292cc7};
test_output[8624] = '{32'h42c34a13};
test_index[8624] = '{2};
test_input[69000:69007] = '{32'hc22c016a, 32'h42bd4814, 32'h411f8d37, 32'h41fda0fe, 32'hc2716ccb, 32'hc1afd905, 32'hc1417fc6, 32'h42c24725};
test_output[8625] = '{32'h42c24725};
test_index[8625] = '{7};
test_input[69008:69015] = '{32'hc2a591fe, 32'h425b8b80, 32'hc2bd3622, 32'h4248d51e, 32'h421cf676, 32'hc1b3c01f, 32'h419da99e, 32'h4143dbea};
test_output[8626] = '{32'h425b8b80};
test_index[8626] = '{1};
test_input[69016:69023] = '{32'hc24c6b78, 32'h42c651b1, 32'hc2568956, 32'h420832f8, 32'h42a393cf, 32'h41e1784e, 32'hc2b93ee6, 32'h410af5b0};
test_output[8627] = '{32'h42c651b1};
test_index[8627] = '{1};
test_input[69024:69031] = '{32'hc2b4afc5, 32'hc1c460a3, 32'hc1da314f, 32'h42a47598, 32'h4278d6e5, 32'hc2a41a44, 32'hc20f6d7b, 32'h40ce8f9f};
test_output[8628] = '{32'h42a47598};
test_index[8628] = '{3};
test_input[69032:69039] = '{32'hc21ee13e, 32'h428af23f, 32'h429dc317, 32'hc21ff213, 32'h42bdbc5d, 32'h4100bbe7, 32'hc1bf5739, 32'h41d4a9f9};
test_output[8629] = '{32'h42bdbc5d};
test_index[8629] = '{4};
test_input[69040:69047] = '{32'h41947666, 32'hc20d56d2, 32'hc1cc99f3, 32'hc2c1dce1, 32'h42950f51, 32'h42470a12, 32'h4228dd3f, 32'h41d9fdca};
test_output[8630] = '{32'h42950f51};
test_index[8630] = '{4};
test_input[69048:69055] = '{32'hc2a8790b, 32'h4232efc0, 32'h425e7524, 32'hc1ff0261, 32'h422b5c5a, 32'h428fb35e, 32'h417d67c1, 32'h4284053d};
test_output[8631] = '{32'h428fb35e};
test_index[8631] = '{5};
test_input[69056:69063] = '{32'hc22baeb5, 32'hc2bc20c2, 32'hc27a22af, 32'h4213268b, 32'h4285c6a5, 32'hc0fb5643, 32'hc29faf63, 32'hc19d634f};
test_output[8632] = '{32'h4285c6a5};
test_index[8632] = '{4};
test_input[69064:69071] = '{32'hc14d5569, 32'h411470bb, 32'h409108cd, 32'hc2b7b50d, 32'hc20ded9b, 32'h41c6aadf, 32'hc28c7365, 32'hc29d4c79};
test_output[8633] = '{32'h41c6aadf};
test_index[8633] = '{5};
test_input[69072:69079] = '{32'h4287b6b5, 32'h42b51c22, 32'h428f8130, 32'hc10a1032, 32'hc2b68326, 32'hbfe9c4c3, 32'h4180912f, 32'h42c1bf49};
test_output[8634] = '{32'h42c1bf49};
test_index[8634] = '{7};
test_input[69080:69087] = '{32'h420afd1c, 32'hc1c9a7d7, 32'h40d96a21, 32'hc19d6a90, 32'hc18af80f, 32'h428054a2, 32'hc2201f96, 32'h42b35f1d};
test_output[8635] = '{32'h42b35f1d};
test_index[8635] = '{7};
test_input[69088:69095] = '{32'hc2c5ae5d, 32'h42b1216c, 32'h42775cf4, 32'h4115d922, 32'hc28dc422, 32'hc2732683, 32'hc2b3df03, 32'h40de6b53};
test_output[8636] = '{32'h42b1216c};
test_index[8636] = '{1};
test_input[69096:69103] = '{32'h40b801ca, 32'hc298397f, 32'h429b2c03, 32'hc17a35bb, 32'h425f8f38, 32'hc2016ce8, 32'h42a252d6, 32'hc2b97a40};
test_output[8637] = '{32'h42a252d6};
test_index[8637] = '{6};
test_input[69104:69111] = '{32'h42319ee6, 32'h4245fbc4, 32'hc2575761, 32'h412fcf5e, 32'h402fe0bc, 32'hc2454b86, 32'h41f4591c, 32'hc2a1fb47};
test_output[8638] = '{32'h4245fbc4};
test_index[8638] = '{1};
test_input[69112:69119] = '{32'h423a0c7c, 32'hc185dbca, 32'h4063f942, 32'hc279a4a7, 32'h423e9e78, 32'h4261f0ab, 32'h408134c7, 32'h4201998b};
test_output[8639] = '{32'h4261f0ab};
test_index[8639] = '{5};
test_input[69120:69127] = '{32'h41c1c3cc, 32'hc2abe4c2, 32'h420c8f8c, 32'h42572bbd, 32'hc2297b00, 32'hc26ea6dd, 32'hbfc60d87, 32'h42bff2ca};
test_output[8640] = '{32'h42bff2ca};
test_index[8640] = '{7};
test_input[69128:69135] = '{32'hc09b3748, 32'hc2b64753, 32'hc1fcc831, 32'hc1cb326d, 32'hc14462ce, 32'h425f4484, 32'hc0c4024a, 32'hc27a86ff};
test_output[8641] = '{32'h425f4484};
test_index[8641] = '{5};
test_input[69136:69143] = '{32'hc2756c11, 32'hc23c653c, 32'h42627c07, 32'hc235746f, 32'hc216be84, 32'hc299c3a5, 32'h427cc8ce, 32'hc2abe094};
test_output[8642] = '{32'h427cc8ce};
test_index[8642] = '{6};
test_input[69144:69151] = '{32'h4207664d, 32'hc2b5e97d, 32'h41d3fb35, 32'h428a96ef, 32'h411340ab, 32'h4296b255, 32'h4220c1f3, 32'hc2125e1f};
test_output[8643] = '{32'h4296b255};
test_index[8643] = '{5};
test_input[69152:69159] = '{32'hc2c412da, 32'hc28d95f7, 32'hc2c5b486, 32'hc1f89274, 32'h40ac1176, 32'hc0c3cae3, 32'h401bbaa6, 32'h40ff2c54};
test_output[8644] = '{32'h40ff2c54};
test_index[8644] = '{7};
test_input[69160:69167] = '{32'h42223afc, 32'h429a7ae7, 32'hc2984d2c, 32'hc2b951c6, 32'h42991ac9, 32'hc1ba52ca, 32'hc2aa5c22, 32'hc2801fc7};
test_output[8645] = '{32'h429a7ae7};
test_index[8645] = '{1};
test_input[69168:69175] = '{32'h4110a0c0, 32'hc2292cc6, 32'hc19257ad, 32'h41bb9b2d, 32'h421270e1, 32'hc2b0e178, 32'hc15807b2, 32'hc214debf};
test_output[8646] = '{32'h421270e1};
test_index[8646] = '{4};
test_input[69176:69183] = '{32'h42a8178f, 32'hc24c2666, 32'hc253163b, 32'h42976a87, 32'h41dfc47e, 32'hc242678b, 32'h421cdfc4, 32'hc28ae7ee};
test_output[8647] = '{32'h42a8178f};
test_index[8647] = '{0};
test_input[69184:69191] = '{32'hc164f214, 32'h42b7a83b, 32'h40ff3426, 32'hc1ed6205, 32'hc1bc6259, 32'h42807f5b, 32'hc2975a78, 32'hbf123f38};
test_output[8648] = '{32'h42b7a83b};
test_index[8648] = '{1};
test_input[69192:69199] = '{32'hc152bd39, 32'h4180f552, 32'h4299a7a5, 32'h425d27a7, 32'h41a6230b, 32'h42335310, 32'hc287d322, 32'hc1c3a6be};
test_output[8649] = '{32'h4299a7a5};
test_index[8649] = '{2};
test_input[69200:69207] = '{32'h4171a830, 32'h40d7688d, 32'h4250ec14, 32'hc2705be9, 32'h4239f89c, 32'hc0a76cd5, 32'hc1ccc67e, 32'h41c98ef6};
test_output[8650] = '{32'h4250ec14};
test_index[8650] = '{2};
test_input[69208:69215] = '{32'hc18ae514, 32'h42b1fceb, 32'h42b8b24c, 32'hc25c4bc6, 32'h41b38cf6, 32'h428009fc, 32'hc2827088, 32'hc214ebf0};
test_output[8651] = '{32'h42b8b24c};
test_index[8651] = '{2};
test_input[69216:69223] = '{32'h429e6a57, 32'h42905075, 32'h4220f15e, 32'hc2a0a780, 32'hc2ab581f, 32'h426d2f37, 32'hc2c47407, 32'h429ece62};
test_output[8652] = '{32'h429ece62};
test_index[8652] = '{7};
test_input[69224:69231] = '{32'h428c7b78, 32'hc28e728c, 32'hc2b85001, 32'hc271c22a, 32'hc2544793, 32'hc231a5fe, 32'h427e7b8a, 32'h42a903da};
test_output[8653] = '{32'h42a903da};
test_index[8653] = '{7};
test_input[69232:69239] = '{32'hc0d8a46b, 32'h4292eabf, 32'h422c18de, 32'hc02598c7, 32'h419fd495, 32'h4254dcb4, 32'h42261877, 32'h41778be2};
test_output[8654] = '{32'h4292eabf};
test_index[8654] = '{1};
test_input[69240:69247] = '{32'h411a8d96, 32'hc11427d1, 32'hc29a1cc8, 32'hc2bc4da7, 32'h42960c31, 32'hc2160bf0, 32'h425a185c, 32'h429e9062};
test_output[8655] = '{32'h429e9062};
test_index[8655] = '{7};
test_input[69248:69255] = '{32'h3f587a9b, 32'h420c69f3, 32'h42b5efa6, 32'hc24d1622, 32'h42a24f38, 32'hc2a39e06, 32'h42142ab2, 32'h41ae0ce7};
test_output[8656] = '{32'h42b5efa6};
test_index[8656] = '{2};
test_input[69256:69263] = '{32'h429dd07d, 32'h42b005c2, 32'h42b02c24, 32'hc252acae, 32'h41efb924, 32'hc2a0b6e1, 32'hc28b7a08, 32'hc2638a6d};
test_output[8657] = '{32'h42b02c24};
test_index[8657] = '{2};
test_input[69264:69271] = '{32'hc28324e0, 32'hc05c8966, 32'hc01e3568, 32'hc22bf7fd, 32'h4292a011, 32'hc185a8cb, 32'hc2852783, 32'h3fe4ba3a};
test_output[8658] = '{32'h4292a011};
test_index[8658] = '{4};
test_input[69272:69279] = '{32'h4293347c, 32'h4247f046, 32'hc25d5a5d, 32'hc1106bc7, 32'hc21cc7c9, 32'h4241fb94, 32'h42149cc5, 32'hc2aac480};
test_output[8659] = '{32'h4293347c};
test_index[8659] = '{0};
test_input[69280:69287] = '{32'h423c447a, 32'h42c1ae3c, 32'hc2b14942, 32'hc1bb7fb4, 32'hc06f3a09, 32'hc2b30af9, 32'hc1d0be73, 32'h4005d026};
test_output[8660] = '{32'h42c1ae3c};
test_index[8660] = '{1};
test_input[69288:69295] = '{32'h428ec9be, 32'hc12d7fd0, 32'hc24b97d7, 32'hc23cc5cc, 32'hc2ad9dba, 32'h42bf4a11, 32'hc296d60f, 32'hc230dd89};
test_output[8661] = '{32'h42bf4a11};
test_index[8661] = '{5};
test_input[69296:69303] = '{32'h427c8f65, 32'h428195b3, 32'h41cb8226, 32'hc13be5f6, 32'hc0667b4d, 32'h423172a5, 32'h42374e4b, 32'h41bace5f};
test_output[8662] = '{32'h428195b3};
test_index[8662] = '{1};
test_input[69304:69311] = '{32'hc1029369, 32'hc2c00e14, 32'hc2a3ee54, 32'h42a7c621, 32'hc230951e, 32'hc25ea270, 32'h414c6a2c, 32'hc270712d};
test_output[8663] = '{32'h42a7c621};
test_index[8663] = '{3};
test_input[69312:69319] = '{32'hc1d72ceb, 32'h3f85cd08, 32'hbf2d0bd3, 32'h424a1976, 32'hc2a48a53, 32'hc207c8c2, 32'h4181330b, 32'h424f524e};
test_output[8664] = '{32'h424f524e};
test_index[8664] = '{7};
test_input[69320:69327] = '{32'h41b68fb9, 32'h428942aa, 32'h4210eb9c, 32'hc23feacb, 32'h42c4dd15, 32'h42295f2b, 32'hc2753e97, 32'h428ef34c};
test_output[8665] = '{32'h42c4dd15};
test_index[8665] = '{4};
test_input[69328:69335] = '{32'h42c18af6, 32'h429bb467, 32'h4263d0bf, 32'h428058ab, 32'h41a136bc, 32'h42a25229, 32'h42259d7b, 32'h42aba7ff};
test_output[8666] = '{32'h42c18af6};
test_index[8666] = '{0};
test_input[69336:69343] = '{32'h410e9b82, 32'hc2bf98b3, 32'hc286e922, 32'h42891b67, 32'hc2aee54e, 32'h4180eed1, 32'hc1c07eef, 32'h4135bb5d};
test_output[8667] = '{32'h42891b67};
test_index[8667] = '{3};
test_input[69344:69351] = '{32'hc102fe2d, 32'hc27a4847, 32'hc2a3efef, 32'h41acccd9, 32'h42a63964, 32'hc2532784, 32'hc1894a64, 32'h42335fef};
test_output[8668] = '{32'h42a63964};
test_index[8668] = '{4};
test_input[69352:69359] = '{32'hc29ab8c0, 32'h40b0f68a, 32'hc21d2dee, 32'h42a2a067, 32'hc1d8d743, 32'h429f47b5, 32'h42788f30, 32'h429e3ece};
test_output[8669] = '{32'h42a2a067};
test_index[8669] = '{3};
test_input[69360:69367] = '{32'h42acfd6d, 32'h42bd9d9e, 32'h417b20ef, 32'h422a27af, 32'hc0930538, 32'hc0ed1803, 32'hc222fd4a, 32'h423e9cf4};
test_output[8670] = '{32'h42bd9d9e};
test_index[8670] = '{1};
test_input[69368:69375] = '{32'hc188722d, 32'hc04fca86, 32'hc12f72ec, 32'h4226f70e, 32'hc03c5a59, 32'hc20eb8e5, 32'hc125c454, 32'h419564ff};
test_output[8671] = '{32'h4226f70e};
test_index[8671] = '{3};
test_input[69376:69383] = '{32'h42c79ab0, 32'hc1c13ac6, 32'hc2a6d109, 32'hc233a0ec, 32'hc288045b, 32'hc23590a4, 32'hc16e746c, 32'hc29586d0};
test_output[8672] = '{32'h42c79ab0};
test_index[8672] = '{0};
test_input[69384:69391] = '{32'hc2ade4f9, 32'h4181e060, 32'h42895899, 32'h42688dc1, 32'hc2be54c1, 32'hc1c471de, 32'hc29e797c, 32'hc2457767};
test_output[8673] = '{32'h42895899};
test_index[8673] = '{2};
test_input[69392:69399] = '{32'hc2158b36, 32'hc2b20b3c, 32'h42c530d4, 32'hc1df2b95, 32'hc1cd3bde, 32'h423457db, 32'hc238faf8, 32'hc2c42e85};
test_output[8674] = '{32'h42c530d4};
test_index[8674] = '{2};
test_input[69400:69407] = '{32'hc2915a20, 32'hc2b3a6e3, 32'hc16ec963, 32'hc292e17c, 32'hc0d48436, 32'h41e73cc5, 32'h427ab79f, 32'h4229c517};
test_output[8675] = '{32'h427ab79f};
test_index[8675] = '{6};
test_input[69408:69415] = '{32'h427d65df, 32'hc1fb4483, 32'h420f0d70, 32'hc1e7bf2c, 32'hc28db3d6, 32'h42a9ece2, 32'hc2165f02, 32'h422edc5c};
test_output[8676] = '{32'h42a9ece2};
test_index[8676] = '{5};
test_input[69416:69423] = '{32'hc1112264, 32'h4164525c, 32'hc25b1f53, 32'h417c38dd, 32'hc2598144, 32'h42a92ca7, 32'hc29553e4, 32'hc2174bf9};
test_output[8677] = '{32'h42a92ca7};
test_index[8677] = '{5};
test_input[69424:69431] = '{32'h4160e325, 32'hc2a83eb9, 32'h4265d1c0, 32'h42b0419f, 32'hc2ac91f3, 32'hc2a1d7cf, 32'h413d9e45, 32'h42b26e85};
test_output[8678] = '{32'h42b26e85};
test_index[8678] = '{7};
test_input[69432:69439] = '{32'h427ff87d, 32'h42943cff, 32'h42b9cb83, 32'h4292ed29, 32'hc241f22b, 32'hc0904156, 32'h4195a111, 32'hc2afed98};
test_output[8679] = '{32'h42b9cb83};
test_index[8679] = '{2};
test_input[69440:69447] = '{32'hc2b73cd1, 32'hc1a864fa, 32'hc2a67a52, 32'h429b9cb3, 32'h41970973, 32'h429d1208, 32'hc2aa3f37, 32'h42c05932};
test_output[8680] = '{32'h42c05932};
test_index[8680] = '{7};
test_input[69448:69455] = '{32'hc1db0796, 32'h42b4fb1b, 32'hc1f3278b, 32'h42aed4b9, 32'h42887fea, 32'hc0cfaaed, 32'hc2337080, 32'h42c6320d};
test_output[8681] = '{32'h42c6320d};
test_index[8681] = '{7};
test_input[69456:69463] = '{32'hc269bd34, 32'hc28bb7df, 32'h41a8f036, 32'h40454d90, 32'h41ad52d0, 32'hc19df8ad, 32'h4128f6a0, 32'h429ce5fc};
test_output[8682] = '{32'h429ce5fc};
test_index[8682] = '{7};
test_input[69464:69471] = '{32'hc058f20c, 32'hc2024831, 32'h419e6f16, 32'hc21a8946, 32'hc28ee285, 32'h41f27e8f, 32'h41b3775f, 32'hc294c2d8};
test_output[8683] = '{32'h41f27e8f};
test_index[8683] = '{5};
test_input[69472:69479] = '{32'hc0b1d897, 32'h41c5a12e, 32'hc25c2e5f, 32'hc201ab63, 32'h42448fc1, 32'h425b9fd2, 32'hc256690c, 32'h42aa0005};
test_output[8684] = '{32'h42aa0005};
test_index[8684] = '{7};
test_input[69480:69487] = '{32'h4288650d, 32'hc183d284, 32'h41f9880f, 32'h424e38f8, 32'hc2063fde, 32'hc2965ab7, 32'h42a652b5, 32'hc1dc2cd2};
test_output[8685] = '{32'h42a652b5};
test_index[8685] = '{6};
test_input[69488:69495] = '{32'h41b989e3, 32'h421f980c, 32'h423131c8, 32'h429ad534, 32'hc140b6f2, 32'h4244fff1, 32'hc24ca236, 32'hc2928934};
test_output[8686] = '{32'h429ad534};
test_index[8686] = '{3};
test_input[69496:69503] = '{32'h41bf4076, 32'h4230f385, 32'h42802c27, 32'hc286dd93, 32'hc1851a1c, 32'h42991241, 32'hc02684b9, 32'hc2ab44ce};
test_output[8687] = '{32'h42991241};
test_index[8687] = '{5};
test_input[69504:69511] = '{32'hc298bbba, 32'hc29e6751, 32'h422b2bf2, 32'hc195db4d, 32'h411d6677, 32'hc074b439, 32'h42a559b9, 32'h42a076b4};
test_output[8688] = '{32'h42a559b9};
test_index[8688] = '{6};
test_input[69512:69519] = '{32'hc2936670, 32'hc20db0df, 32'h41d92c7b, 32'hc1a4f716, 32'hc1d0fe17, 32'hc2be9cd8, 32'h427028d5, 32'hc2809b04};
test_output[8689] = '{32'h427028d5};
test_index[8689] = '{6};
test_input[69520:69527] = '{32'hc2bae6be, 32'hc274dee6, 32'h42b0efa1, 32'h40538e0f, 32'hc238c8c8, 32'hc2b71e7e, 32'h41debc32, 32'h41bd7d0d};
test_output[8690] = '{32'h42b0efa1};
test_index[8690] = '{2};
test_input[69528:69535] = '{32'h41ae12fe, 32'hc2c2d2ee, 32'h429532ba, 32'hc0b51e41, 32'h4180f66e, 32'h419fe0aa, 32'h410f023a, 32'h4284508d};
test_output[8691] = '{32'h429532ba};
test_index[8691] = '{2};
test_input[69536:69543] = '{32'h42005482, 32'h40b97b3c, 32'h421865b7, 32'h41d45c9a, 32'hc21da915, 32'hc2532316, 32'hc28fc5b8, 32'hbee9e70c};
test_output[8692] = '{32'h421865b7};
test_index[8692] = '{2};
test_input[69544:69551] = '{32'hc1800420, 32'hc2830228, 32'h42a14957, 32'hc19eabd6, 32'hc2421e18, 32'hc2255a5b, 32'hc255bc8a, 32'h425f606d};
test_output[8693] = '{32'h42a14957};
test_index[8693] = '{2};
test_input[69552:69559] = '{32'h4279600d, 32'h428f45f0, 32'h41f39d14, 32'h4119c924, 32'hc1e4d8e6, 32'h42589481, 32'h41003fde, 32'hc22c8d2b};
test_output[8694] = '{32'h428f45f0};
test_index[8694] = '{1};
test_input[69560:69567] = '{32'hc2bb4237, 32'hc1a27175, 32'hc2b3eadf, 32'hc2a6288e, 32'h3e8289ce, 32'h429097ce, 32'h42be4370, 32'h419a1dc0};
test_output[8695] = '{32'h42be4370};
test_index[8695] = '{6};
test_input[69568:69575] = '{32'hc2208cb4, 32'h42184934, 32'hc2a0e4fc, 32'hc1859ab4, 32'h4284ec62, 32'h4283c267, 32'hc2beff1e, 32'h4256dc84};
test_output[8696] = '{32'h4284ec62};
test_index[8696] = '{4};
test_input[69576:69583] = '{32'hc1fba130, 32'h4243a94e, 32'hc29ab23b, 32'h422f983f, 32'h421a6469, 32'h41f0a824, 32'hc2c4dccf, 32'h4228388b};
test_output[8697] = '{32'h4243a94e};
test_index[8697] = '{1};
test_input[69584:69591] = '{32'hc29a7367, 32'hc1bf4e9b, 32'h42466074, 32'h429818e2, 32'h428e4885, 32'h423f2061, 32'h41dc46f5, 32'hc2784d77};
test_output[8698] = '{32'h429818e2};
test_index[8698] = '{3};
test_input[69592:69599] = '{32'hc2250edd, 32'hc2a9d67f, 32'hc2a2ce89, 32'h4286cb09, 32'hc25d37e6, 32'h426d89d3, 32'h42b2e7a0, 32'h42c1e775};
test_output[8699] = '{32'h42c1e775};
test_index[8699] = '{7};
test_input[69600:69607] = '{32'hc1d193d1, 32'h4085fa6c, 32'hc2adc5ac, 32'hc29c23f5, 32'h42c3aa13, 32'hc1313660, 32'hc24cf663, 32'h4226994c};
test_output[8700] = '{32'h42c3aa13};
test_index[8700] = '{4};
test_input[69608:69615] = '{32'h42b3c29c, 32'h42c32f91, 32'h41eafa03, 32'h422b72ed, 32'hc2adaba1, 32'hc0547d90, 32'hc27e4ca6, 32'h424f77f0};
test_output[8701] = '{32'h42c32f91};
test_index[8701] = '{1};
test_input[69616:69623] = '{32'hc1e5981a, 32'hc1961d99, 32'h42296163, 32'h42c23db3, 32'hc1bc3c74, 32'h42356121, 32'hc1f6f7c6, 32'hc243d4ca};
test_output[8702] = '{32'h42c23db3};
test_index[8702] = '{3};
test_input[69624:69631] = '{32'hc17cfb72, 32'h423fc8a7, 32'hc2c53725, 32'h429cb9cd, 32'h42a7f5e0, 32'hc2ae8e61, 32'hc2c30feb, 32'h42abb2b2};
test_output[8703] = '{32'h42abb2b2};
test_index[8703] = '{7};
test_input[69632:69639] = '{32'hc2623b54, 32'hc2968c13, 32'h42c2cf35, 32'hc2a18f70, 32'hc19d5284, 32'h4082f396, 32'h41c2a76a, 32'hc2a5ac7f};
test_output[8704] = '{32'h42c2cf35};
test_index[8704] = '{2};
test_input[69640:69647] = '{32'hc28a34cc, 32'h42c1ead7, 32'hc1b503b4, 32'hc20cc7b1, 32'hc285ee1d, 32'hc15273b7, 32'hc1df8dad, 32'hc26a1512};
test_output[8705] = '{32'h42c1ead7};
test_index[8705] = '{1};
test_input[69648:69655] = '{32'h415cedc7, 32'h42996759, 32'hc264b5f6, 32'h42a7c66a, 32'hc2ab8e22, 32'hc14967bc, 32'h42b1c246, 32'hc24bfbcd};
test_output[8706] = '{32'h42b1c246};
test_index[8706] = '{6};
test_input[69656:69663] = '{32'hc286e9cc, 32'hc2c75bf8, 32'h4271d339, 32'h423d27aa, 32'hc141b4b3, 32'hc1f8d91a, 32'h42940316, 32'h41cab7f9};
test_output[8707] = '{32'h42940316};
test_index[8707] = '{6};
test_input[69664:69671] = '{32'h41845c47, 32'h41059035, 32'h41dfe15e, 32'h41ef4bc0, 32'h41af222c, 32'h42c3a459, 32'h428d9105, 32'hc205a39b};
test_output[8708] = '{32'h42c3a459};
test_index[8708] = '{5};
test_input[69672:69679] = '{32'hc284039c, 32'h4264dab1, 32'hc24f2bdd, 32'hc2b8c3b7, 32'hc24849a9, 32'h41633122, 32'h42b08a32, 32'h4146bd2f};
test_output[8709] = '{32'h42b08a32};
test_index[8709] = '{6};
test_input[69680:69687] = '{32'hc1a91c5a, 32'h42b9f3f3, 32'h42278d9a, 32'h42021809, 32'h42c6fb72, 32'hc2129b0d, 32'hc1e06c88, 32'hc2c5eea3};
test_output[8710] = '{32'h42c6fb72};
test_index[8710] = '{4};
test_input[69688:69695] = '{32'hc2500785, 32'hc20d2394, 32'hc2603a07, 32'h41e7aa42, 32'hc25835c5, 32'hc1e6f506, 32'hc2b2b42f, 32'hc252bc8e};
test_output[8711] = '{32'h41e7aa42};
test_index[8711] = '{3};
test_input[69696:69703] = '{32'h41ebeb99, 32'hc2537db8, 32'hc2474adb, 32'h3fa9039e, 32'hc25841e6, 32'h4299aa1b, 32'hc290cc4a, 32'hc1eb6659};
test_output[8712] = '{32'h4299aa1b};
test_index[8712] = '{5};
test_input[69704:69711] = '{32'h4110b83b, 32'h41c96a0f, 32'hc2473681, 32'hc21ed093, 32'hc22d09c9, 32'h41b8de0e, 32'h427f2458, 32'h42c178ac};
test_output[8713] = '{32'h42c178ac};
test_index[8713] = '{7};
test_input[69712:69719] = '{32'hc17dd96a, 32'hc1060147, 32'hc23beb85, 32'h423c98dd, 32'h42a2a06a, 32'hc2bf35f9, 32'h429c6fdb, 32'hc2b33fed};
test_output[8714] = '{32'h42a2a06a};
test_index[8714] = '{4};
test_input[69720:69727] = '{32'h42201225, 32'h40a3872a, 32'h425e6cb1, 32'h42ad04bc, 32'hc022d029, 32'hc204fb0a, 32'h429bd012, 32'hc27374e1};
test_output[8715] = '{32'h42ad04bc};
test_index[8715] = '{3};
test_input[69728:69735] = '{32'h417145f1, 32'hc2b8a8ce, 32'h428258e3, 32'h4222dd54, 32'h428c9b49, 32'hc27afb30, 32'h4198712e, 32'h42a64e63};
test_output[8716] = '{32'h42a64e63};
test_index[8716] = '{7};
test_input[69736:69743] = '{32'hc224cf55, 32'h427c6e0b, 32'h42bc3f8a, 32'h425275f2, 32'hc2a77bea, 32'h4194f62b, 32'hc2139a0c, 32'hc058d864};
test_output[8717] = '{32'h42bc3f8a};
test_index[8717] = '{2};
test_input[69744:69751] = '{32'hc2c5a0c3, 32'h42538b59, 32'h41c72f24, 32'h42295dab, 32'h429a0774, 32'hc1d877d5, 32'h40d38152, 32'hc299003c};
test_output[8718] = '{32'h429a0774};
test_index[8718] = '{4};
test_input[69752:69759] = '{32'h41b610d1, 32'h422991ca, 32'hc2139206, 32'h411ab970, 32'h423d8da5, 32'hc27c57a2, 32'h42af384d, 32'hc070a38f};
test_output[8719] = '{32'h42af384d};
test_index[8719] = '{6};
test_input[69760:69767] = '{32'hc192f0fa, 32'h42c69db4, 32'h405cee41, 32'hc0c99672, 32'h42c1e6c2, 32'h4280eedd, 32'h42c6b82b, 32'h42b489f7};
test_output[8720] = '{32'h42c6b82b};
test_index[8720] = '{6};
test_input[69768:69775] = '{32'hc2bc2404, 32'hc185b5c0, 32'hc2a217cf, 32'hc27a4c46, 32'h423db71e, 32'h420630f9, 32'h4259d12b, 32'h3a52d0a8};
test_output[8721] = '{32'h4259d12b};
test_index[8721] = '{6};
test_input[69776:69783] = '{32'h41cc5aa7, 32'hc29e777e, 32'h42381e68, 32'hc2bf3e6d, 32'hc1b22284, 32'h40b7bc40, 32'hc1c5008b, 32'h42822050};
test_output[8722] = '{32'h42822050};
test_index[8722] = '{7};
test_input[69784:69791] = '{32'hc1f86467, 32'h426e79f8, 32'h4299756d, 32'hc29b4f87, 32'hc2a31654, 32'hc24d3003, 32'h40c35556, 32'h3d8968ff};
test_output[8723] = '{32'h4299756d};
test_index[8723] = '{2};
test_input[69792:69799] = '{32'hc294464c, 32'h42c3ae7b, 32'hc20988b7, 32'h41800337, 32'h424a93db, 32'hc290df43, 32'hc1a27d11, 32'hc1998523};
test_output[8724] = '{32'h42c3ae7b};
test_index[8724] = '{1};
test_input[69800:69807] = '{32'hc2b31d5f, 32'h3f43710b, 32'h40cca7df, 32'h41fe7196, 32'hc28ee3db, 32'h42c6555a, 32'h42aa6079, 32'hc2883fca};
test_output[8725] = '{32'h42c6555a};
test_index[8725] = '{5};
test_input[69808:69815] = '{32'hc2b146ef, 32'h41e1f82c, 32'hc292e3f4, 32'h41d586ed, 32'h418f26be, 32'hc1a79f0d, 32'hc2920a23, 32'h424771c1};
test_output[8726] = '{32'h424771c1};
test_index[8726] = '{7};
test_input[69816:69823] = '{32'h429d5fab, 32'hc2af750c, 32'hc2949c1a, 32'h42c74fbe, 32'hc2be1be7, 32'h42259250, 32'hc2b9588d, 32'hc2879f82};
test_output[8727] = '{32'h42c74fbe};
test_index[8727] = '{3};
test_input[69824:69831] = '{32'h422c17c0, 32'hc2a1a96b, 32'hc28727e4, 32'hc1673564, 32'hc2a437ee, 32'h4210cdd1, 32'hc21ecc11, 32'hc219c8d6};
test_output[8728] = '{32'h422c17c0};
test_index[8728] = '{0};
test_input[69832:69839] = '{32'hc19cad02, 32'hc2a65aa0, 32'hc186e1b4, 32'h428d2b5f, 32'hc2636d78, 32'h42bd72f8, 32'hc1a6a360, 32'hc15c9c80};
test_output[8729] = '{32'h42bd72f8};
test_index[8729] = '{5};
test_input[69840:69847] = '{32'hc2b6f365, 32'h424a3898, 32'h4061bba1, 32'hc2591443, 32'h4236e270, 32'h41fec716, 32'hc2b6f6b1, 32'h422248e7};
test_output[8730] = '{32'h424a3898};
test_index[8730] = '{1};
test_input[69848:69855] = '{32'hc2158f96, 32'h41c27f2d, 32'h42216276, 32'h41fc2029, 32'hc25e4f98, 32'h4299f111, 32'hc14b007b, 32'hc23ac572};
test_output[8731] = '{32'h4299f111};
test_index[8731] = '{5};
test_input[69856:69863] = '{32'hc1f499fb, 32'h42c20a6f, 32'h42be26f6, 32'h40286c78, 32'hc22d43a7, 32'h41a18b8f, 32'hc1b53045, 32'hc14fa638};
test_output[8732] = '{32'h42c20a6f};
test_index[8732] = '{1};
test_input[69864:69871] = '{32'hc2913fc8, 32'hc1b638a8, 32'h425fc29e, 32'hbec2b7c6, 32'hc2a378b5, 32'h4287a456, 32'h421a06fe, 32'hc2801e13};
test_output[8733] = '{32'h4287a456};
test_index[8733] = '{5};
test_input[69872:69879] = '{32'hc2a08c56, 32'hc238e333, 32'hc2bca449, 32'h41bd499b, 32'hc2396dc9, 32'hc222ab2e, 32'h42abb2d7, 32'h429c54d5};
test_output[8734] = '{32'h42abb2d7};
test_index[8734] = '{6};
test_input[69880:69887] = '{32'h41d02d30, 32'hc1bc9696, 32'h4223a5b8, 32'h414b67ba, 32'hc2c79b16, 32'h428662c0, 32'h420bb091, 32'h4227e097};
test_output[8735] = '{32'h428662c0};
test_index[8735] = '{5};
test_input[69888:69895] = '{32'h4281f69f, 32'h42004188, 32'hc086b9c4, 32'h429730ef, 32'hc136a616, 32'hc129f069, 32'h424b38d6, 32'h42ae0e26};
test_output[8736] = '{32'h42ae0e26};
test_index[8736] = '{7};
test_input[69896:69903] = '{32'h4233ca27, 32'hc27882a6, 32'h42a501a5, 32'h40be7464, 32'hc26cd7e1, 32'hc2b7fab2, 32'h4282a16e, 32'h42be6103};
test_output[8737] = '{32'h42be6103};
test_index[8737] = '{7};
test_input[69904:69911] = '{32'hc1c2de42, 32'h41591124, 32'hc2428309, 32'hc2a22b52, 32'hc251052a, 32'h412c0627, 32'h41a77d4c, 32'h42351431};
test_output[8738] = '{32'h42351431};
test_index[8738] = '{7};
test_input[69912:69919] = '{32'h42032a45, 32'hc18d08ba, 32'hc11f614e, 32'h42155301, 32'h424c716c, 32'hc2c66113, 32'h42559016, 32'hc2bd5b14};
test_output[8739] = '{32'h42559016};
test_index[8739] = '{6};
test_input[69920:69927] = '{32'hc2b33e60, 32'hc2c1bc59, 32'h426d9e53, 32'h41cbea63, 32'hc2bb7d30, 32'hc26912a4, 32'h42bee080, 32'h3f82a075};
test_output[8740] = '{32'h42bee080};
test_index[8740] = '{6};
test_input[69928:69935] = '{32'hc29bcce6, 32'hc29ef3e1, 32'hc277c30f, 32'h4248226c, 32'h428cc00a, 32'hc120292c, 32'h42c7214c, 32'h4085d8e1};
test_output[8741] = '{32'h42c7214c};
test_index[8741] = '{6};
test_input[69936:69943] = '{32'h4245394b, 32'h428be61f, 32'h419a6042, 32'h418046e2, 32'h41974d63, 32'hc243b6bf, 32'hc2088dfa, 32'h423c450b};
test_output[8742] = '{32'h428be61f};
test_index[8742] = '{1};
test_input[69944:69951] = '{32'hc2b7d7b2, 32'hc22d9da8, 32'hc2441f49, 32'hc2be3701, 32'h4264e8bc, 32'hc28551eb, 32'hc16aff24, 32'h426c093c};
test_output[8743] = '{32'h426c093c};
test_index[8743] = '{7};
test_input[69952:69959] = '{32'h425953de, 32'h427002b1, 32'h428b8a3d, 32'hc29083ba, 32'hc2bddc91, 32'hc18f89fa, 32'h41a64c02, 32'hc281b4d8};
test_output[8744] = '{32'h428b8a3d};
test_index[8744] = '{2};
test_input[69960:69967] = '{32'h42800bdb, 32'h425da0ca, 32'hc1abf73b, 32'h41543423, 32'hc1bf3321, 32'h427a4b51, 32'h41eed4ae, 32'hc116b913};
test_output[8745] = '{32'h42800bdb};
test_index[8745] = '{0};
test_input[69968:69975] = '{32'hc2c6064e, 32'hc2995e01, 32'h428d6df4, 32'h4203bf85, 32'hc2abff1e, 32'hc246ed73, 32'h41b99682, 32'hc299d77a};
test_output[8746] = '{32'h428d6df4};
test_index[8746] = '{2};
test_input[69976:69983] = '{32'hc28b0f3b, 32'h41a3d280, 32'hc2564956, 32'hc1a75380, 32'hc2416c62, 32'h42677329, 32'h4234c9f5, 32'hc1de3801};
test_output[8747] = '{32'h42677329};
test_index[8747] = '{5};
test_input[69984:69991] = '{32'hc1f3e477, 32'h42a2d861, 32'h421b7b53, 32'h42971c11, 32'h429a9e4d, 32'h4208974d, 32'hc0cc8533, 32'h4227625f};
test_output[8748] = '{32'h42a2d861};
test_index[8748] = '{1};
test_input[69992:69999] = '{32'h4244f4c1, 32'hc2a2a78a, 32'hc1ae991f, 32'hc075dbcc, 32'h4221c890, 32'h42bd9b39, 32'h4297804f, 32'h40146b31};
test_output[8749] = '{32'h42bd9b39};
test_index[8749] = '{5};
test_input[70000:70007] = '{32'hc25d69a6, 32'h42877c9c, 32'h42345660, 32'h4267fa77, 32'hc1b9eab9, 32'hc12a2a9d, 32'h3fb1df9d, 32'h4289e565};
test_output[8750] = '{32'h4289e565};
test_index[8750] = '{7};
test_input[70008:70015] = '{32'hc18220bf, 32'h41ff862c, 32'h429428a0, 32'hc0c386de, 32'h42c308b0, 32'hc262b1f0, 32'hc2235794, 32'hc20b9325};
test_output[8751] = '{32'h42c308b0};
test_index[8751] = '{4};
test_input[70016:70023] = '{32'h429d4671, 32'hc238a5c7, 32'hc2c07031, 32'hc183b20f, 32'hc29fe9a3, 32'hc28e0d08, 32'hc19af55a, 32'h428fbed7};
test_output[8752] = '{32'h429d4671};
test_index[8752] = '{0};
test_input[70024:70031] = '{32'hc2692806, 32'h41d0902d, 32'hbff70c71, 32'h41abeafe, 32'h4249bf48, 32'h4138c467, 32'h400698b9, 32'h4147f186};
test_output[8753] = '{32'h4249bf48};
test_index[8753] = '{4};
test_input[70032:70039] = '{32'hc2238a0c, 32'hc245a71a, 32'hc2b6f5d4, 32'h41fccf37, 32'hc2b5ff22, 32'h41577a2b, 32'h4290facc, 32'hc0c0cf3b};
test_output[8754] = '{32'h4290facc};
test_index[8754] = '{6};
test_input[70040:70047] = '{32'hc2b6771b, 32'h423d307b, 32'h429c752d, 32'hc21d185c, 32'h422b4a01, 32'h42553c26, 32'h41cd75a4, 32'hc28be176};
test_output[8755] = '{32'h429c752d};
test_index[8755] = '{2};
test_input[70048:70055] = '{32'hc165a934, 32'hc2ba496b, 32'h4285f694, 32'hc275c2e2, 32'hc2ac799b, 32'hc2066175, 32'h420d9f1a, 32'h42a0a183};
test_output[8756] = '{32'h42a0a183};
test_index[8756] = '{7};
test_input[70056:70063] = '{32'hc2ae05bb, 32'hc23ce87c, 32'hc1a53447, 32'hc24a61ba, 32'h42003792, 32'h4297b16f, 32'hc2afcf79, 32'h4287d7dd};
test_output[8757] = '{32'h4297b16f};
test_index[8757] = '{5};
test_input[70064:70071] = '{32'hc24ce373, 32'hc1a9ab0f, 32'hc2484f28, 32'h4235bb51, 32'h4192ed6f, 32'hc253139f, 32'hc29d09a5, 32'hc2b7f825};
test_output[8758] = '{32'h4235bb51};
test_index[8758] = '{3};
test_input[70072:70079] = '{32'h420e7c02, 32'h40cbf6a2, 32'hc19a12f4, 32'hc2471dcf, 32'h42851c9b, 32'hc151d01a, 32'hc2838e24, 32'h423f2589};
test_output[8759] = '{32'h42851c9b};
test_index[8759] = '{4};
test_input[70080:70087] = '{32'hc2a85fd3, 32'h419abca9, 32'hc2c16456, 32'hc1ecd38a, 32'hc0e33c63, 32'h42a986e0, 32'hc21c5f85, 32'h3f519682};
test_output[8760] = '{32'h42a986e0};
test_index[8760] = '{5};
test_input[70088:70095] = '{32'hc131f084, 32'hc26d51c7, 32'hc23d7b9e, 32'hc139f58e, 32'hc19cb617, 32'h425a3450, 32'hc21b24f5, 32'h427f6fa1};
test_output[8761] = '{32'h427f6fa1};
test_index[8761] = '{7};
test_input[70096:70103] = '{32'hc2a034b4, 32'hc1fdf318, 32'hc285e391, 32'hc2b4d783, 32'hc2bfa324, 32'h4288dfb9, 32'h4258cc59, 32'hc2451269};
test_output[8762] = '{32'h4288dfb9};
test_index[8762] = '{5};
test_input[70104:70111] = '{32'h42344505, 32'h42c07f8f, 32'hc23c8497, 32'h41d309e5, 32'hc1961a46, 32'hc0037c0b, 32'hc26f5efb, 32'h4289e15c};
test_output[8763] = '{32'h42c07f8f};
test_index[8763] = '{1};
test_input[70112:70119] = '{32'hc17ad074, 32'hc1887bb0, 32'h42332b02, 32'hc23ff52e, 32'hc21d954a, 32'hc2953e69, 32'hc1ce225e, 32'h41d40392};
test_output[8764] = '{32'h42332b02};
test_index[8764] = '{2};
test_input[70120:70127] = '{32'hc28046ea, 32'h3f30d830, 32'h42307cb6, 32'h42696bca, 32'h418f35ce, 32'h41aa724a, 32'hc1ffa934, 32'h42b01358};
test_output[8765] = '{32'h42b01358};
test_index[8765] = '{7};
test_input[70128:70135] = '{32'hc0926065, 32'h3fc90462, 32'h42bceaff, 32'h42bd2235, 32'h402a6bfa, 32'hc09b0c51, 32'hc2a203f2, 32'hc28236e8};
test_output[8766] = '{32'h42bd2235};
test_index[8766] = '{3};
test_input[70136:70143] = '{32'h42271e97, 32'h42150644, 32'hc1420e05, 32'hc22f5065, 32'hc2381e96, 32'h41d80e9b, 32'h41ff3736, 32'hc293626a};
test_output[8767] = '{32'h42271e97};
test_index[8767] = '{0};
test_input[70144:70151] = '{32'h416d36fa, 32'hc1ba70d5, 32'h41a3b6f9, 32'hc1762ec0, 32'h4231f131, 32'h4281ba82, 32'hc25e5836, 32'h42a19f46};
test_output[8768] = '{32'h42a19f46};
test_index[8768] = '{7};
test_input[70152:70159] = '{32'hc2058efa, 32'h42729ecc, 32'hc2572da2, 32'hc2ae06e0, 32'hc0530374, 32'h42258e41, 32'h42bdd73c, 32'h4287dd38};
test_output[8769] = '{32'h42bdd73c};
test_index[8769] = '{6};
test_input[70160:70167] = '{32'hc23e2258, 32'hc20ba1c9, 32'h426f4255, 32'hc20c3048, 32'hc2a7c33d, 32'h421ef670, 32'h421a92d0, 32'h42a07f3b};
test_output[8770] = '{32'h42a07f3b};
test_index[8770] = '{7};
test_input[70168:70175] = '{32'h4196aaf7, 32'hc143e087, 32'hc10a3b5e, 32'hc27ada9e, 32'hc29c4148, 32'hc2b095db, 32'h41cb58c1, 32'h41c03b26};
test_output[8771] = '{32'h41cb58c1};
test_index[8771] = '{6};
test_input[70176:70183] = '{32'h428b7d69, 32'h42957eec, 32'h41f9a529, 32'h426e9c32, 32'hc291b4fd, 32'hc0ba9a7f, 32'hc0bcbd49, 32'hc29b9e6b};
test_output[8772] = '{32'h42957eec};
test_index[8772] = '{1};
test_input[70184:70191] = '{32'hc27cc720, 32'h42a9e179, 32'h40fc8dc0, 32'hc254ca14, 32'h41930a8e, 32'h42bf567a, 32'hc2a61283, 32'hc2c6f533};
test_output[8773] = '{32'h42bf567a};
test_index[8773] = '{5};
test_input[70192:70199] = '{32'h4261c6ad, 32'h42ba9f8e, 32'hc2ab140b, 32'hc147b27d, 32'h424ec89e, 32'h42bb3dba, 32'hc224be3b, 32'h427a0523};
test_output[8774] = '{32'h42bb3dba};
test_index[8774] = '{5};
test_input[70200:70207] = '{32'h426586e0, 32'h422ccc1f, 32'hc089bb5e, 32'hc207b152, 32'hc0ae3db2, 32'h41bea091, 32'h425cbefb, 32'hc1fd5125};
test_output[8775] = '{32'h426586e0};
test_index[8775] = '{0};
test_input[70208:70215] = '{32'hc28cd27d, 32'hc1d08836, 32'hc2067a4f, 32'h41d7a11e, 32'h42386986, 32'hc073b139, 32'h42b971dd, 32'h4195a1a4};
test_output[8776] = '{32'h42b971dd};
test_index[8776] = '{6};
test_input[70216:70223] = '{32'h4284177d, 32'h41107845, 32'h41669fc7, 32'hc2ad9b7f, 32'hc251f3fd, 32'hc10f8790, 32'hc221b763, 32'hc1ce8404};
test_output[8777] = '{32'h4284177d};
test_index[8777] = '{0};
test_input[70224:70231] = '{32'hc2adcbff, 32'h42b43e76, 32'h42330dcc, 32'h4254a5e3, 32'hc2005ee4, 32'h3f0eaf58, 32'hc27f5ff0, 32'h42843438};
test_output[8778] = '{32'h42b43e76};
test_index[8778] = '{1};
test_input[70232:70239] = '{32'hc1a28252, 32'h3f60c0e6, 32'hc246ad6c, 32'h42c5a8a7, 32'h423204c2, 32'h423c07b3, 32'hc258c202, 32'h42223431};
test_output[8779] = '{32'h42c5a8a7};
test_index[8779] = '{3};
test_input[70240:70247] = '{32'hc2b7cb3b, 32'h429c5ca3, 32'h42204597, 32'hc2981fd1, 32'hc186389f, 32'hc2bc5d35, 32'hc2984b38, 32'h42b7d780};
test_output[8780] = '{32'h42b7d780};
test_index[8780] = '{7};
test_input[70248:70255] = '{32'hc2419640, 32'h42991ce8, 32'hc2a5193a, 32'hc2355534, 32'hc0958b51, 32'h420cbda0, 32'h41d7eeaf, 32'hc2546918};
test_output[8781] = '{32'h42991ce8};
test_index[8781] = '{1};
test_input[70256:70263] = '{32'h42c6740d, 32'hc237ef1b, 32'hc2293693, 32'hc26e368a, 32'h4050be0f, 32'hc28986dc, 32'hc14858f0, 32'h42228ef0};
test_output[8782] = '{32'h42c6740d};
test_index[8782] = '{0};
test_input[70264:70271] = '{32'hc2b136c1, 32'hc2476ef5, 32'hc21fa412, 32'hbef91fce, 32'h424bb3eb, 32'h418d02d0, 32'hc19f7491, 32'hc28ae87d};
test_output[8783] = '{32'h424bb3eb};
test_index[8783] = '{4};
test_input[70272:70279] = '{32'h3fc917d5, 32'hc1cd8180, 32'hc24cd057, 32'hc18183f9, 32'hc2c1b9bd, 32'hc12ca87c, 32'h41b394da, 32'hc182d596};
test_output[8784] = '{32'h41b394da};
test_index[8784] = '{6};
test_input[70280:70287] = '{32'h429ca29a, 32'h42973878, 32'hc2af8cfc, 32'h42547e3e, 32'h41ae2ed9, 32'hc29f5207, 32'h4219d941, 32'h42bdaeb6};
test_output[8785] = '{32'h42bdaeb6};
test_index[8785] = '{7};
test_input[70288:70295] = '{32'hc259ccfe, 32'hc2583acb, 32'h4226d91c, 32'h4277d466, 32'hc2a9a3f7, 32'hc24d049a, 32'h422bb037, 32'hc166e041};
test_output[8786] = '{32'h4277d466};
test_index[8786] = '{3};
test_input[70296:70303] = '{32'hc24602f7, 32'h4197a123, 32'h400ca3aa, 32'hc1e86f89, 32'h415f4d41, 32'h42b0a412, 32'h4222e9b0, 32'hc2808c5d};
test_output[8787] = '{32'h42b0a412};
test_index[8787] = '{5};
test_input[70304:70311] = '{32'h422e07b3, 32'hc280bc96, 32'h42302717, 32'hc1bab323, 32'h4286553b, 32'h42acf1a8, 32'hc1174fdd, 32'hc1da941b};
test_output[8788] = '{32'h42acf1a8};
test_index[8788] = '{5};
test_input[70312:70319] = '{32'h420443e8, 32'h41c144c0, 32'h41cfcb83, 32'hc29e0066, 32'hc1878661, 32'hc2bde32c, 32'h423c1f50, 32'hc2a86020};
test_output[8789] = '{32'h423c1f50};
test_index[8789] = '{6};
test_input[70320:70327] = '{32'hc24d7af7, 32'hc2353130, 32'h429fba3c, 32'hc20f2936, 32'h419b26ef, 32'h41b114fd, 32'hc1964463, 32'h42afc327};
test_output[8790] = '{32'h42afc327};
test_index[8790] = '{7};
test_input[70328:70335] = '{32'h4212cb11, 32'h40c1d550, 32'h427dfa33, 32'h426e62d5, 32'h4157bad2, 32'hc21c58c9, 32'hc204755b, 32'h4274dd0a};
test_output[8791] = '{32'h427dfa33};
test_index[8791] = '{2};
test_input[70336:70343] = '{32'hc1407b8d, 32'h424ac8f4, 32'h423101c4, 32'hc207c9de, 32'hc251b642, 32'h421c3c1f, 32'h42782908, 32'hc170696b};
test_output[8792] = '{32'h42782908};
test_index[8792] = '{6};
test_input[70344:70351] = '{32'h42acadc3, 32'hc1dd969e, 32'hc245530c, 32'hc2895f8a, 32'hc2697763, 32'hc1344cb0, 32'hc2bb3584, 32'hc1a3f827};
test_output[8793] = '{32'h42acadc3};
test_index[8793] = '{0};
test_input[70352:70359] = '{32'hc1e958f4, 32'hc27eaaac, 32'h41842620, 32'hc2c5a830, 32'hc2310cfa, 32'h425e3f94, 32'h42052fa0, 32'hc2470826};
test_output[8794] = '{32'h425e3f94};
test_index[8794] = '{5};
test_input[70360:70367] = '{32'h420ab092, 32'hc2495ac5, 32'h3f15371e, 32'hc02beb70, 32'hc223b70c, 32'hc262a19d, 32'h425be2fd, 32'h41c10708};
test_output[8795] = '{32'h425be2fd};
test_index[8795] = '{6};
test_input[70368:70375] = '{32'hc2922f0f, 32'h42babff2, 32'h4189f032, 32'hc1ed0101, 32'hc08d61df, 32'hc232541f, 32'hc1309ab9, 32'h4295c5e4};
test_output[8796] = '{32'h42babff2};
test_index[8796] = '{1};
test_input[70376:70383] = '{32'h4272b16f, 32'h42167767, 32'h419fc2db, 32'hc220c844, 32'h4265e983, 32'h425cb612, 32'h418416e9, 32'hc23344e6};
test_output[8797] = '{32'h4272b16f};
test_index[8797] = '{0};
test_input[70384:70391] = '{32'hc271c371, 32'h408446f8, 32'hc2979a94, 32'hc2bf396c, 32'h429e5c81, 32'hc2694ae9, 32'hc14094b4, 32'hc2b671d8};
test_output[8798] = '{32'h429e5c81};
test_index[8798] = '{4};
test_input[70392:70399] = '{32'h4036c345, 32'hc2127ce3, 32'h4241fd7e, 32'hc2ae7243, 32'hc192ebe6, 32'hc292f721, 32'hc1c64ea2, 32'h4259d851};
test_output[8799] = '{32'h4259d851};
test_index[8799] = '{7};
test_input[70400:70407] = '{32'h41e78d26, 32'hc26e6f6f, 32'hc2b04fbf, 32'hc1e35bfc, 32'h4230360c, 32'h421b19dc, 32'hc2a02a77, 32'hc28a24a0};
test_output[8800] = '{32'h4230360c};
test_index[8800] = '{4};
test_input[70408:70415] = '{32'h41943a40, 32'h42c00db1, 32'hc2503092, 32'h4274de9e, 32'hc1e67406, 32'h424725af, 32'hc270c996, 32'h41ca1dcb};
test_output[8801] = '{32'h42c00db1};
test_index[8801] = '{1};
test_input[70416:70423] = '{32'h42238826, 32'hc2b85af4, 32'h42aa4e6c, 32'hc126ab2e, 32'h4216e786, 32'hc2bb1aac, 32'h423f72ae, 32'hc1940a7b};
test_output[8802] = '{32'h42aa4e6c};
test_index[8802] = '{2};
test_input[70424:70431] = '{32'h42b34688, 32'h4275beae, 32'h4133f752, 32'h4101b1fe, 32'hc1be28c9, 32'hc177f85f, 32'h42a682b6, 32'h4257ee7e};
test_output[8803] = '{32'h42b34688};
test_index[8803] = '{0};
test_input[70432:70439] = '{32'h41983bdb, 32'hc13540b4, 32'hc0120199, 32'h420e4a2a, 32'hc29b7dcd, 32'h4255b188, 32'hc255eb34, 32'h4107be34};
test_output[8804] = '{32'h4255b188};
test_index[8804] = '{5};
test_input[70440:70447] = '{32'hc249f328, 32'hc24d6cb7, 32'hc19e6a5b, 32'hc1d98cdb, 32'h4223cec3, 32'h4234e7c9, 32'h417f8384, 32'hc2200d39};
test_output[8805] = '{32'h4234e7c9};
test_index[8805] = '{5};
test_input[70448:70455] = '{32'hc268c282, 32'hc202d841, 32'hc2c03fcc, 32'h413ce06a, 32'hc1cf1894, 32'h4202415c, 32'h41301853, 32'h420e4e5e};
test_output[8806] = '{32'h420e4e5e};
test_index[8806] = '{7};
test_input[70456:70463] = '{32'hc24366f0, 32'hc298c3d8, 32'hc294a5a6, 32'h425e45dd, 32'hc1918df7, 32'hc2c077b1, 32'hc2b4ec06, 32'hc2c43690};
test_output[8807] = '{32'h425e45dd};
test_index[8807] = '{3};
test_input[70464:70471] = '{32'h428d7fdc, 32'h42534505, 32'h4135895c, 32'hc28e6c74, 32'hc2383596, 32'hc2b2f73b, 32'h4290ad2f, 32'hc2387545};
test_output[8808] = '{32'h4290ad2f};
test_index[8808] = '{6};
test_input[70472:70479] = '{32'hc2bd8186, 32'hc2a58937, 32'h423eb2ba, 32'hc262fe04, 32'h427030e4, 32'hc29ead2c, 32'hc1ae75d9, 32'h42195f8c};
test_output[8809] = '{32'h427030e4};
test_index[8809] = '{4};
test_input[70480:70487] = '{32'h42c46d58, 32'hc1fd3c00, 32'hc1ec88e9, 32'h4267cd77, 32'h4112d638, 32'hc2b88420, 32'hc1cd1ebd, 32'hc1833b9a};
test_output[8810] = '{32'h42c46d58};
test_index[8810] = '{0};
test_input[70488:70495] = '{32'h40a6c9be, 32'hc2733202, 32'h420bfb42, 32'h420a332b, 32'hc2ac2bb2, 32'h42228a13, 32'h4149ba35, 32'hc2bf34b1};
test_output[8811] = '{32'h42228a13};
test_index[8811] = '{5};
test_input[70496:70503] = '{32'hc26f4872, 32'hc1bd4dd3, 32'h4294b945, 32'h4280262f, 32'hc12bc219, 32'h42bdba81, 32'hc22cd2cd, 32'hc1d37cf1};
test_output[8812] = '{32'h42bdba81};
test_index[8812] = '{5};
test_input[70504:70511] = '{32'h42c6dc00, 32'h427e327d, 32'h41c80bab, 32'hc2a92643, 32'h42269335, 32'h428f471b, 32'h42c344cc, 32'hc19cf8a6};
test_output[8813] = '{32'h42c6dc00};
test_index[8813] = '{0};
test_input[70512:70519] = '{32'hc1956832, 32'hc231979e, 32'hc27868f9, 32'h427d9b6b, 32'hc1485665, 32'hc0c238e7, 32'hc2affb82, 32'h42882043};
test_output[8814] = '{32'h42882043};
test_index[8814] = '{7};
test_input[70520:70527] = '{32'h41a1b735, 32'h4198bfa6, 32'h426257eb, 32'hc279a86b, 32'h4271cf3f, 32'hc29accc2, 32'h42b86e69, 32'hc2471a37};
test_output[8815] = '{32'h42b86e69};
test_index[8815] = '{6};
test_input[70528:70535] = '{32'hc20b49ca, 32'hc29cee17, 32'h4282805b, 32'h4294fbfa, 32'hc20db2f1, 32'hc2b60900, 32'hc162356b, 32'h429a2957};
test_output[8816] = '{32'h429a2957};
test_index[8816] = '{7};
test_input[70536:70543] = '{32'h42344e3e, 32'h42367c5b, 32'h41d989b2, 32'h41e9d896, 32'h42c7ae36, 32'h42557af1, 32'hc237a946, 32'hc1abce60};
test_output[8817] = '{32'h42c7ae36};
test_index[8817] = '{4};
test_input[70544:70551] = '{32'hc2b9aa75, 32'h427ba6d6, 32'h417be063, 32'h42c59289, 32'hc2a7a3e0, 32'hc2223c93, 32'h42bcb991, 32'hc1631f80};
test_output[8818] = '{32'h42c59289};
test_index[8818] = '{3};
test_input[70552:70559] = '{32'h4201f5a3, 32'hc21d92d6, 32'hc23445de, 32'h42bafc3f, 32'h4294e454, 32'hc29b05a4, 32'h42bddbdf, 32'hc0b52f72};
test_output[8819] = '{32'h42bddbdf};
test_index[8819] = '{6};
test_input[70560:70567] = '{32'hc2b3c0c9, 32'h429adb98, 32'hc23d57bc, 32'hc2b891b9, 32'hc185fb78, 32'h425b6afb, 32'h414ad891, 32'h4231c665};
test_output[8820] = '{32'h429adb98};
test_index[8820] = '{1};
test_input[70568:70575] = '{32'h42b7b444, 32'hc2c1cc18, 32'hc1f7a63f, 32'hc1800233, 32'h4287314d, 32'hbf5453d6, 32'h426f6a47, 32'hc1a31048};
test_output[8821] = '{32'h42b7b444};
test_index[8821] = '{0};
test_input[70576:70583] = '{32'h421910ea, 32'hc1435ad3, 32'h424051bc, 32'h421d6319, 32'h4271cb9d, 32'h42013dd5, 32'h409dc290, 32'hc2addfeb};
test_output[8822] = '{32'h4271cb9d};
test_index[8822] = '{4};
test_input[70584:70591] = '{32'h42484fa4, 32'h4280aada, 32'hc2760331, 32'h41a6f109, 32'h418dac22, 32'hc28ba36a, 32'h42aee99a, 32'h425ec5a9};
test_output[8823] = '{32'h42aee99a};
test_index[8823] = '{6};
test_input[70592:70599] = '{32'hc279b88c, 32'hc2723d24, 32'h429f071a, 32'hc0210f09, 32'hc26ef889, 32'hc28bb6f2, 32'h429610f2, 32'hc20a0066};
test_output[8824] = '{32'h429f071a};
test_index[8824] = '{2};
test_input[70600:70607] = '{32'h4241903f, 32'hbf4d97e6, 32'h4202390d, 32'h4298e182, 32'h42487da1, 32'hc2aca61a, 32'h4238c468, 32'hc2c5029b};
test_output[8825] = '{32'h4298e182};
test_index[8825] = '{3};
test_input[70608:70615] = '{32'h4286e217, 32'h3f5da25e, 32'h4297eb17, 32'hc2886eea, 32'h421100eb, 32'hc204e0dc, 32'h427b5235, 32'h4198d9cd};
test_output[8826] = '{32'h4297eb17};
test_index[8826] = '{2};
test_input[70616:70623] = '{32'h4258ae3d, 32'hc25f3d6d, 32'h4297ab32, 32'h42b8ed9b, 32'hc1bc100e, 32'hc091f557, 32'hc1f364b4, 32'h409e2f2b};
test_output[8827] = '{32'h42b8ed9b};
test_index[8827] = '{3};
test_input[70624:70631] = '{32'hc0de6408, 32'hc2c71d53, 32'hc28a9220, 32'h42b40a9e, 32'hc2bbb125, 32'hc28ab8c8, 32'hc2af42ef, 32'h42c3d6e2};
test_output[8828] = '{32'h42c3d6e2};
test_index[8828] = '{7};
test_input[70632:70639] = '{32'hc199f98f, 32'h42b31a2c, 32'hc28068f8, 32'h40250405, 32'h41f0aaf9, 32'h42290158, 32'h4205d67a, 32'hc20fa46b};
test_output[8829] = '{32'h42b31a2c};
test_index[8829] = '{1};
test_input[70640:70647] = '{32'hc2b5bb39, 32'h41ec5a0c, 32'h4258ee8d, 32'hc14f5299, 32'hc1e477ad, 32'hc14f6736, 32'hc27977a9, 32'h42366fc5};
test_output[8830] = '{32'h4258ee8d};
test_index[8830] = '{2};
test_input[70648:70655] = '{32'hc276bc19, 32'hc18ccf51, 32'h41a1ae29, 32'hc28a22f8, 32'h42b27f45, 32'hc1083a36, 32'hc27d0577, 32'hc2be22a4};
test_output[8831] = '{32'h42b27f45};
test_index[8831] = '{4};
test_input[70656:70663] = '{32'h42775840, 32'hc0f2468e, 32'hc2859a84, 32'hc2581dd4, 32'hc12a5c4e, 32'hc1b53842, 32'hc243256c, 32'hc2a43863};
test_output[8832] = '{32'h42775840};
test_index[8832] = '{0};
test_input[70664:70671] = '{32'h401fc532, 32'h3f7ab6da, 32'h426e1b5b, 32'h42199f23, 32'hc2a956c2, 32'h417b6bf6, 32'h41292be6, 32'h427d5e63};
test_output[8833] = '{32'h427d5e63};
test_index[8833] = '{7};
test_input[70672:70679] = '{32'h421aa710, 32'hc2bc2182, 32'hc29fcfed, 32'hc17b96eb, 32'hc1565a5f, 32'hc1e5ff9d, 32'h42c2ca72, 32'h410f866b};
test_output[8834] = '{32'h42c2ca72};
test_index[8834] = '{6};
test_input[70680:70687] = '{32'hbfb88cc7, 32'hc15126e5, 32'hc2a159e7, 32'hc2b2f7d4, 32'h42c5addc, 32'h428ca1b2, 32'h414e9f79, 32'hc1293e1d};
test_output[8835] = '{32'h42c5addc};
test_index[8835] = '{4};
test_input[70688:70695] = '{32'hc212b969, 32'hc2135cba, 32'h41be2e46, 32'hc26f2ba4, 32'h41a70b3f, 32'hc21f51de, 32'hc266fca0, 32'hc1d44a22};
test_output[8836] = '{32'h41be2e46};
test_index[8836] = '{2};
test_input[70696:70703] = '{32'hc1ba81c7, 32'hc2382bd9, 32'hc294dde1, 32'h42689458, 32'h426e11d3, 32'h42995d14, 32'h40cd2925, 32'hc2619ad3};
test_output[8837] = '{32'h42995d14};
test_index[8837] = '{5};
test_input[70704:70711] = '{32'h418a568f, 32'hc25d0d52, 32'hc244847d, 32'h42bb797a, 32'hc2ad2b9d, 32'h42b17ec5, 32'hc20a7421, 32'h411f8c6d};
test_output[8838] = '{32'h42bb797a};
test_index[8838] = '{3};
test_input[70712:70719] = '{32'h422d19e2, 32'h429d06d7, 32'h4246bd10, 32'h42042279, 32'h4248cf34, 32'hc224b9f8, 32'h4211252f, 32'hc1bd82a6};
test_output[8839] = '{32'h429d06d7};
test_index[8839] = '{1};
test_input[70720:70727] = '{32'h42af9774, 32'hc28bb9ae, 32'h4201862d, 32'h42ab10a4, 32'h41d04af1, 32'hc237befa, 32'hc27cdc1a, 32'h4296b4ab};
test_output[8840] = '{32'h42af9774};
test_index[8840] = '{0};
test_input[70728:70735] = '{32'hc26995a4, 32'h42126df7, 32'h42c4cb6f, 32'h42b4f437, 32'hc286f9df, 32'h41bed7ed, 32'hc2814935, 32'hc195d9ae};
test_output[8841] = '{32'h42c4cb6f};
test_index[8841] = '{2};
test_input[70736:70743] = '{32'h403a649d, 32'hc2bad86c, 32'h42b76fbd, 32'hc2aef069, 32'hc2b39f14, 32'h42a2de06, 32'hc278923b, 32'h428ec7de};
test_output[8842] = '{32'h42b76fbd};
test_index[8842] = '{2};
test_input[70744:70751] = '{32'h42c69c8a, 32'hc2905fc8, 32'h4211df51, 32'hc11446c3, 32'hbd2d584f, 32'h41525a0b, 32'h3e55bfa0, 32'hc2a5336a};
test_output[8843] = '{32'h42c69c8a};
test_index[8843] = '{0};
test_input[70752:70759] = '{32'hc229ceb2, 32'hc29f2672, 32'hc0828773, 32'hc261c760, 32'h42b21635, 32'hc265a096, 32'h42b56aeb, 32'hc1f6a8fa};
test_output[8844] = '{32'h42b56aeb};
test_index[8844] = '{6};
test_input[70760:70767] = '{32'hc18ec8fb, 32'hc284a15e, 32'h4217b408, 32'hc2903f88, 32'hc0b9486a, 32'h41eedbb5, 32'h428e681a, 32'h40d4d4b6};
test_output[8845] = '{32'h428e681a};
test_index[8845] = '{6};
test_input[70768:70775] = '{32'hc2bbcb82, 32'hc265b875, 32'hc1b729de, 32'hc264dffd, 32'hc2966a31, 32'hc28648ac, 32'h40c38972, 32'hc0c0b556};
test_output[8846] = '{32'h40c38972};
test_index[8846] = '{6};
test_input[70776:70783] = '{32'h42c734c5, 32'h4234470c, 32'hc281542d, 32'h42b37821, 32'hc2a770c0, 32'hc13c8384, 32'hc01d91f5, 32'h4241ef93};
test_output[8847] = '{32'h42c734c5};
test_index[8847] = '{0};
test_input[70784:70791] = '{32'h42975063, 32'h41db4f2c, 32'h42a29299, 32'hc275fe3a, 32'h42544a18, 32'hc2404dba, 32'hc220495a, 32'h42307dc8};
test_output[8848] = '{32'h42a29299};
test_index[8848] = '{2};
test_input[70792:70799] = '{32'hc276c484, 32'h42172f3d, 32'hc2797f3e, 32'hc25848d8, 32'h424e8a2b, 32'hc22cabbd, 32'hc2b6f0e5, 32'h41841bd6};
test_output[8849] = '{32'h424e8a2b};
test_index[8849] = '{4};
test_input[70800:70807] = '{32'hc2c3b082, 32'hc2bb1411, 32'h422235b3, 32'hc0b87848, 32'hc1c6651c, 32'hc1b04b54, 32'hc28ff3d2, 32'hc27b73c1};
test_output[8850] = '{32'h422235b3};
test_index[8850] = '{2};
test_input[70808:70815] = '{32'h405ec021, 32'h41829be6, 32'hc22ae35e, 32'h42a4b61a, 32'h42afaca4, 32'h413486f5, 32'hc28cb905, 32'h41339ae8};
test_output[8851] = '{32'h42afaca4};
test_index[8851] = '{4};
test_input[70816:70823] = '{32'h41d92865, 32'h42412d43, 32'hc2afb0c7, 32'h4293e9b1, 32'hc24b2d6b, 32'h425c142d, 32'h4285c98a, 32'h42083277};
test_output[8852] = '{32'h4293e9b1};
test_index[8852] = '{3};
test_input[70824:70831] = '{32'h41e6d402, 32'hc22d5ba3, 32'hc229c5e4, 32'hc2103480, 32'h4249a04e, 32'h42ac8e87, 32'h41938ac3, 32'hc2bb049a};
test_output[8853] = '{32'h42ac8e87};
test_index[8853] = '{5};
test_input[70832:70839] = '{32'h422c7346, 32'hc0c426d5, 32'h40eb8b55, 32'h42182315, 32'hc2a68cfd, 32'h420eec57, 32'h4278d76b, 32'hc21c9d3a};
test_output[8854] = '{32'h4278d76b};
test_index[8854] = '{6};
test_input[70840:70847] = '{32'h429fc356, 32'hc1e8d177, 32'h4289e112, 32'hc1b13c2a, 32'hc2ba4304, 32'hc279b583, 32'hc290f9ed, 32'hc20d9e04};
test_output[8855] = '{32'h429fc356};
test_index[8855] = '{0};
test_input[70848:70855] = '{32'h420cf302, 32'hc1d0fb82, 32'hc24dac87, 32'hc21d51dc, 32'h42153fd6, 32'hc1ef6476, 32'h4211ce81, 32'h428261e4};
test_output[8856] = '{32'h428261e4};
test_index[8856] = '{7};
test_input[70856:70863] = '{32'hc29650f0, 32'h42a49ad1, 32'h41d8078d, 32'hc121fa95, 32'h41a6c2a4, 32'h416e9b66, 32'h42610d97, 32'h4277393b};
test_output[8857] = '{32'h42a49ad1};
test_index[8857] = '{1};
test_input[70864:70871] = '{32'h41ce58cc, 32'hc0bb7e5d, 32'hbffca42e, 32'hc1ad9f16, 32'hc10843a8, 32'h42a440fa, 32'hc298f83b, 32'h42c2d5d1};
test_output[8858] = '{32'h42c2d5d1};
test_index[8858] = '{7};
test_input[70872:70879] = '{32'hc257a7ec, 32'hc266aa28, 32'hc2ba2126, 32'hc1a41798, 32'hc085791b, 32'hc2a76910, 32'h42a6f760, 32'h4181d45c};
test_output[8859] = '{32'h42a6f760};
test_index[8859] = '{6};
test_input[70880:70887] = '{32'hc20929e5, 32'hc19b866b, 32'h42759b91, 32'hc0abb75f, 32'h42ab1d19, 32'h4283fc33, 32'h421aa4c8, 32'h42b07ec7};
test_output[8860] = '{32'h42b07ec7};
test_index[8860] = '{7};
test_input[70888:70895] = '{32'h42b64444, 32'hc2a0d686, 32'hc25c2ca0, 32'hc2a0a969, 32'hc2a8dbc3, 32'hc2b6f343, 32'h42971405, 32'h4214a17e};
test_output[8861] = '{32'h42b64444};
test_index[8861] = '{0};
test_input[70896:70903] = '{32'h41469cbc, 32'hc20aa77a, 32'h4293d0f0, 32'hc2a0472d, 32'hc1b41bc8, 32'hc2838780, 32'hc22127ba, 32'h42ada8f1};
test_output[8862] = '{32'h42ada8f1};
test_index[8862] = '{7};
test_input[70904:70911] = '{32'h429351c6, 32'h4281171c, 32'hc12522bc, 32'h42afea0a, 32'hc2c5e0bf, 32'h416cd576, 32'hc29e309e, 32'h42b095c7};
test_output[8863] = '{32'h42b095c7};
test_index[8863] = '{7};
test_input[70912:70919] = '{32'h4222a67e, 32'hc25390c9, 32'hc28d08b4, 32'h427f3c53, 32'hc29a2708, 32'h410f864a, 32'h427db03d, 32'h42132937};
test_output[8864] = '{32'h427f3c53};
test_index[8864] = '{3};
test_input[70920:70927] = '{32'hc2b20d65, 32'hc2a96084, 32'hc2b9b864, 32'hc1f5acd4, 32'hc2aa81e4, 32'h413fb20e, 32'h4272816f, 32'h4157de9d};
test_output[8865] = '{32'h4272816f};
test_index[8865] = '{6};
test_input[70928:70935] = '{32'hc2aea357, 32'hc2068a7c, 32'h42c42544, 32'hc2c33b5a, 32'h42b00501, 32'h415ad4cf, 32'hc119e532, 32'hc287aa02};
test_output[8866] = '{32'h42c42544};
test_index[8866] = '{2};
test_input[70936:70943] = '{32'hc2abeb16, 32'hc0c296ba, 32'hc2449b89, 32'h42367974, 32'h407fb06c, 32'hc2971d43, 32'hc0a49f5f, 32'hc247bf4d};
test_output[8867] = '{32'h42367974};
test_index[8867] = '{3};
test_input[70944:70951] = '{32'h425d6e2f, 32'hc241eb91, 32'hc21d132d, 32'hc1dc60a5, 32'hc223ef38, 32'hc2941b4e, 32'h42801b28, 32'hc23b0219};
test_output[8868] = '{32'h42801b28};
test_index[8868] = '{6};
test_input[70952:70959] = '{32'h42836dbb, 32'hc2ad3d12, 32'h41b95ec4, 32'hc2222c5a, 32'hc2267ad4, 32'h41bf66e3, 32'hc27010c6, 32'hc2c0fead};
test_output[8869] = '{32'h42836dbb};
test_index[8869] = '{0};
test_input[70960:70967] = '{32'h41b2721b, 32'hc10a76b8, 32'hc08585a4, 32'hc2bbb168, 32'hc1844115, 32'hc20f420d, 32'hc2c6e154, 32'h421070f3};
test_output[8870] = '{32'h421070f3};
test_index[8870] = '{7};
test_input[70968:70975] = '{32'hc12e739c, 32'hc160f8ca, 32'h42926c83, 32'h422c8f32, 32'h42bca5df, 32'h42b97b22, 32'hc1f5c0e9, 32'h42850349};
test_output[8871] = '{32'h42bca5df};
test_index[8871] = '{4};
test_input[70976:70983] = '{32'h3fcbc8ef, 32'hc23061e8, 32'h428fd9b6, 32'h421097fd, 32'hc1d6b617, 32'hc2900f26, 32'h42268f3f, 32'hc2aebec1};
test_output[8872] = '{32'h428fd9b6};
test_index[8872] = '{2};
test_input[70984:70991] = '{32'h41bef397, 32'hc1e87f10, 32'hc19f1d0b, 32'hc2b2af94, 32'hc0673b93, 32'h42786d1d, 32'hc23266a6, 32'hc2807ace};
test_output[8873] = '{32'h42786d1d};
test_index[8873] = '{5};
test_input[70992:70999] = '{32'h42039f24, 32'hc1e25eab, 32'h422c39af, 32'hc22c1dcc, 32'hc290f2fe, 32'h41c7be2e, 32'hc1b0fa64, 32'h3fd4aab1};
test_output[8874] = '{32'h422c39af};
test_index[8874] = '{2};
test_input[71000:71007] = '{32'h4295b9c3, 32'h4186e5e8, 32'h42806fff, 32'h42a65473, 32'h426f4fdd, 32'hc2069fd2, 32'hc18dd3ba, 32'h42c78edd};
test_output[8875] = '{32'h42c78edd};
test_index[8875] = '{7};
test_input[71008:71015] = '{32'hc2af0e07, 32'h42adfdf7, 32'hc03eb267, 32'hc1634af5, 32'hc26a3940, 32'h410fb3d6, 32'h4211251d, 32'h4234c7d0};
test_output[8876] = '{32'h42adfdf7};
test_index[8876] = '{1};
test_input[71016:71023] = '{32'hc2067034, 32'hc29a9853, 32'h41b5e417, 32'hc202f812, 32'h42aeb129, 32'hc2a34f30, 32'h428b2423, 32'h428bfbe3};
test_output[8877] = '{32'h42aeb129};
test_index[8877] = '{4};
test_input[71024:71031] = '{32'h41b7a0e5, 32'h41c67fc2, 32'hc105fa7d, 32'h4285c371, 32'hc2bd66e9, 32'h4004128a, 32'hc0cbdc62, 32'hc2a75a59};
test_output[8878] = '{32'h4285c371};
test_index[8878] = '{3};
test_input[71032:71039] = '{32'h424a8f84, 32'hc1e2da69, 32'hc2be439a, 32'hc1b7ee28, 32'hc29e5a92, 32'hc22aa6dc, 32'hc1f72c2d, 32'h423f82ac};
test_output[8879] = '{32'h424a8f84};
test_index[8879] = '{0};
test_input[71040:71047] = '{32'h42847f74, 32'hc2b0b50c, 32'h41e719c4, 32'h4252ab9c, 32'h42a9b3fb, 32'hc216705c, 32'h42131c38, 32'h42aa8a23};
test_output[8880] = '{32'h42aa8a23};
test_index[8880] = '{7};
test_input[71048:71055] = '{32'h4284a6b4, 32'h41c43197, 32'hbf7ee3db, 32'hc1bb0be7, 32'hc16dcfa5, 32'hc2879e8a, 32'hc209a820, 32'hc2c3decb};
test_output[8881] = '{32'h4284a6b4};
test_index[8881] = '{0};
test_input[71056:71063] = '{32'hc11441ec, 32'hc2a981d3, 32'hc2b95c17, 32'h418c2151, 32'h42b6fa85, 32'hc2112f60, 32'h429e447e, 32'h4296c209};
test_output[8882] = '{32'h42b6fa85};
test_index[8882] = '{4};
test_input[71064:71071] = '{32'h42239451, 32'h3ffcd8a9, 32'hc1bfa84d, 32'h427fea71, 32'hc19382f5, 32'hc27bb6d9, 32'h40b27aee, 32'hc2afae93};
test_output[8883] = '{32'h427fea71};
test_index[8883] = '{3};
test_input[71072:71079] = '{32'hc2af519d, 32'hbf10f37f, 32'hc2953705, 32'hc28542e7, 32'hc2b91a77, 32'h4117e594, 32'h42a6bc1a, 32'h42650eed};
test_output[8884] = '{32'h42a6bc1a};
test_index[8884] = '{6};
test_input[71080:71087] = '{32'h41d61742, 32'hc1878aa8, 32'h41de62cd, 32'hc208f20b, 32'hc2be3900, 32'h415aa3ce, 32'h4128b089, 32'hc0c03cc1};
test_output[8885] = '{32'h41de62cd};
test_index[8885] = '{2};
test_input[71088:71095] = '{32'h426a9101, 32'h4262427b, 32'h4252dfcd, 32'h425b94d4, 32'h416e66c7, 32'hc1977fe3, 32'hc2918ef7, 32'h41cc56c8};
test_output[8886] = '{32'h426a9101};
test_index[8886] = '{0};
test_input[71096:71103] = '{32'h42051e09, 32'hc26ce1e9, 32'hc2188f44, 32'h4295b851, 32'hc238a5d7, 32'h4225b4ec, 32'h422c6e20, 32'h424ae9dc};
test_output[8887] = '{32'h4295b851};
test_index[8887] = '{3};
test_input[71104:71111] = '{32'hc0f6f639, 32'hc12d5c20, 32'hc232dcaa, 32'h4218b896, 32'h4284371c, 32'h429eaa3c, 32'h4296d25e, 32'hbfe91250};
test_output[8888] = '{32'h429eaa3c};
test_index[8888] = '{5};
test_input[71112:71119] = '{32'h42b99b86, 32'hc2708aae, 32'h417c4401, 32'h41c6d71b, 32'hc2259735, 32'h42a0b9a9, 32'hc28f8e4d, 32'h42200c67};
test_output[8889] = '{32'h42b99b86};
test_index[8889] = '{0};
test_input[71120:71127] = '{32'h41dedd94, 32'h42029209, 32'h41832d3a, 32'h42a91bd3, 32'h42be4f33, 32'hc2be3155, 32'h428b5375, 32'h4195d6a6};
test_output[8890] = '{32'h42be4f33};
test_index[8890] = '{4};
test_input[71128:71135] = '{32'h429f6160, 32'h42a40f38, 32'hc2b17106, 32'hbfe60cba, 32'h41f759fb, 32'hc2aaf94d, 32'hc2936fc1, 32'hc1a3f274};
test_output[8891] = '{32'h42a40f38};
test_index[8891] = '{1};
test_input[71136:71143] = '{32'h428a60de, 32'h4080d6c7, 32'hbf546fdb, 32'hc2c7d97d, 32'hc1f4a1f0, 32'h41f8f3ae, 32'hc29c4e3d, 32'h42b4adde};
test_output[8892] = '{32'h42b4adde};
test_index[8892] = '{7};
test_input[71144:71151] = '{32'h42352efe, 32'h42b96287, 32'h421fb774, 32'hc1cbc0f2, 32'h4202f9dc, 32'h424cce73, 32'hc2b6d936, 32'h427d4b11};
test_output[8893] = '{32'h42b96287};
test_index[8893] = '{1};
test_input[71152:71159] = '{32'h41fdd765, 32'hc2afaa11, 32'h42402c85, 32'hc2081326, 32'hc267b701, 32'hc2471704, 32'h41b8b0a5, 32'hc2bae4c7};
test_output[8894] = '{32'h42402c85};
test_index[8894] = '{2};
test_input[71160:71167] = '{32'h41b62364, 32'hc165bd60, 32'h42026075, 32'hc21605fb, 32'h42512cc6, 32'hc26fa3e5, 32'h4107757f, 32'hc2aabdc4};
test_output[8895] = '{32'h42512cc6};
test_index[8895] = '{4};
test_input[71168:71175] = '{32'hc0de4624, 32'h412a9a8d, 32'h40975f54, 32'hc1dcbed5, 32'h422d46f0, 32'h420b3149, 32'h42896fc8, 32'h4080588b};
test_output[8896] = '{32'h42896fc8};
test_index[8896] = '{6};
test_input[71176:71183] = '{32'hc261ef75, 32'h3f709cbd, 32'h429a72b9, 32'h424c2ea8, 32'h41e2a0b7, 32'hc20db24a, 32'h42c42371, 32'hc24c5c9a};
test_output[8897] = '{32'h42c42371};
test_index[8897] = '{6};
test_input[71184:71191] = '{32'h42081b6f, 32'h41c9cb39, 32'h42b7bc59, 32'hc05b3a2c, 32'h429ac843, 32'hc201d376, 32'hc2611901, 32'hc231170b};
test_output[8898] = '{32'h42b7bc59};
test_index[8898] = '{2};
test_input[71192:71199] = '{32'hc22ae293, 32'h425d748d, 32'hc10d0083, 32'hc0121efd, 32'h41c92846, 32'hc2735a2d, 32'h4288933a, 32'hc2191564};
test_output[8899] = '{32'h4288933a};
test_index[8899] = '{6};
test_input[71200:71207] = '{32'hc07c85c1, 32'hc271af97, 32'hc26db0a0, 32'h4295c13a, 32'hc1fd4c09, 32'hc2b3c052, 32'hc22d452e, 32'h413a2917};
test_output[8900] = '{32'h4295c13a};
test_index[8900] = '{3};
test_input[71208:71215] = '{32'h415fe463, 32'hc2bade8f, 32'h41154e0f, 32'hc212e607, 32'hc24c0622, 32'h42ab940f, 32'hc21035a4, 32'h41303c1d};
test_output[8901] = '{32'h42ab940f};
test_index[8901] = '{5};
test_input[71216:71223] = '{32'hc2a9576a, 32'hc0585028, 32'h4154b886, 32'hc284c9d7, 32'hc293fc73, 32'hc1d01d17, 32'hc290c548, 32'hc281bc2c};
test_output[8902] = '{32'h4154b886};
test_index[8902] = '{2};
test_input[71224:71231] = '{32'h42bd4b8c, 32'h42912877, 32'hc2ad0fdf, 32'hc266b449, 32'h4280a765, 32'h4243f2fd, 32'hc1f8aa22, 32'hc222324d};
test_output[8903] = '{32'h42bd4b8c};
test_index[8903] = '{0};
test_input[71232:71239] = '{32'hc2802ce4, 32'h418512bf, 32'hc284c05a, 32'hc1b62906, 32'hc29dd889, 32'h428db010, 32'h41afb8b0, 32'h41d7c457};
test_output[8904] = '{32'h428db010};
test_index[8904] = '{5};
test_input[71240:71247] = '{32'hc28d4235, 32'h42a92a02, 32'hc290fb91, 32'h42a6caf0, 32'h42914a53, 32'h42861177, 32'hc2be7aea, 32'h3fd81565};
test_output[8905] = '{32'h42a92a02};
test_index[8905] = '{1};
test_input[71248:71255] = '{32'h420c6278, 32'h42a1bebc, 32'hc2a3b82d, 32'hc2a4827e, 32'hc2a103dc, 32'hc23722c7, 32'hc083417c, 32'h4238628d};
test_output[8906] = '{32'h42a1bebc};
test_index[8906] = '{1};
test_input[71256:71263] = '{32'h4290979f, 32'hc2c56552, 32'h42076c83, 32'hbf9785e1, 32'h42b6538d, 32'hc288c146, 32'h429d36be, 32'h418864ec};
test_output[8907] = '{32'h42b6538d};
test_index[8907] = '{4};
test_input[71264:71271] = '{32'hc2a1c2c7, 32'hc1d62c1d, 32'hc20c80fc, 32'h4197667f, 32'h41c82ed1, 32'hc21518dd, 32'hc236fa8c, 32'hc15db05c};
test_output[8908] = '{32'h41c82ed1};
test_index[8908] = '{4};
test_input[71272:71279] = '{32'hc2c459d2, 32'hc28af774, 32'hc2a5cc39, 32'h3fd3e67c, 32'h4212b496, 32'hc2189cd9, 32'h40c76881, 32'hc2aefe12};
test_output[8909] = '{32'h4212b496};
test_index[8909] = '{4};
test_input[71280:71287] = '{32'hc1058be9, 32'hc2c1b78c, 32'h42b21e37, 32'h4211d8cd, 32'hc22910da, 32'hc29cb4a1, 32'h405d5cc9, 32'h41a5abdf};
test_output[8910] = '{32'h42b21e37};
test_index[8910] = '{2};
test_input[71288:71295] = '{32'h42b44d44, 32'h41f7f115, 32'hc27d9306, 32'hc19af97d, 32'h42aaa7ae, 32'hc1340f81, 32'h40763b4c, 32'hc2bb207a};
test_output[8911] = '{32'h42b44d44};
test_index[8911] = '{0};
test_input[71296:71303] = '{32'h42326663, 32'h418d94d1, 32'hc22f6c6f, 32'hc1aee831, 32'h4282d5dc, 32'h40224123, 32'hc2be6385, 32'hc2ac39cf};
test_output[8912] = '{32'h4282d5dc};
test_index[8912] = '{4};
test_input[71304:71311] = '{32'h42b7ddd3, 32'hc215f2bc, 32'h41e8c524, 32'h429e5b42, 32'h4272e0bc, 32'hc20c3f69, 32'h42055a10, 32'h41d4a293};
test_output[8913] = '{32'h42b7ddd3};
test_index[8913] = '{0};
test_input[71312:71319] = '{32'hc2643107, 32'h420db699, 32'h42aefc27, 32'h4293876c, 32'h42bbc27f, 32'hc2b57cd1, 32'h4233edb4, 32'hc2bcc5c9};
test_output[8914] = '{32'h42bbc27f};
test_index[8914] = '{4};
test_input[71320:71327] = '{32'hc2254ade, 32'h4030e66d, 32'h42833713, 32'hc1cce587, 32'hc2aebb83, 32'hc195b0e5, 32'hc2c6237a, 32'hc2bcfa23};
test_output[8915] = '{32'h42833713};
test_index[8915] = '{2};
test_input[71328:71335] = '{32'hc24d62b0, 32'hc20bb343, 32'hc2c0de5c, 32'hc0155702, 32'h428905ce, 32'h42baf39d, 32'hc2bb401d, 32'hc1f4e553};
test_output[8916] = '{32'h42baf39d};
test_index[8916] = '{5};
test_input[71336:71343] = '{32'h41afd707, 32'hc2953cc6, 32'hc2397cd2, 32'h427715e0, 32'hc26d5f75, 32'h41bd3e58, 32'h42c0db26, 32'hc2a42a45};
test_output[8917] = '{32'h42c0db26};
test_index[8917] = '{6};
test_input[71344:71351] = '{32'h419db018, 32'h4228cb10, 32'hc0f8dd69, 32'hc2823fa1, 32'hc18add6f, 32'h4214620f, 32'hc1eee536, 32'h42a3d11a};
test_output[8918] = '{32'h42a3d11a};
test_index[8918] = '{7};
test_input[71352:71359] = '{32'hc05a866f, 32'hc23d4637, 32'hc233a04f, 32'hc21f9aa1, 32'hc28fbafb, 32'h4137ceca, 32'h429cefb6, 32'hc176af14};
test_output[8919] = '{32'h429cefb6};
test_index[8919] = '{6};
test_input[71360:71367] = '{32'h42c047e0, 32'hc268dc96, 32'hc28bc89a, 32'h426e1243, 32'hc2b1e312, 32'hbf92594e, 32'h420809f0, 32'h425f6f91};
test_output[8920] = '{32'h42c047e0};
test_index[8920] = '{0};
test_input[71368:71375] = '{32'h41def71e, 32'hc28e66fb, 32'hc273193f, 32'hc2bbc39e, 32'h428eb569, 32'hc1a80f22, 32'h42501cf3, 32'hc23118e4};
test_output[8921] = '{32'h428eb569};
test_index[8921] = '{4};
test_input[71376:71383] = '{32'hc2a2600c, 32'hc28fd321, 32'hc21eeb28, 32'hc2c25979, 32'h420eb963, 32'h4208dfbc, 32'hc1cd175a, 32'h40438d1c};
test_output[8922] = '{32'h420eb963};
test_index[8922] = '{4};
test_input[71384:71391] = '{32'hc2b08022, 32'h4287c6a6, 32'hc1a617ca, 32'hc2c68c2e, 32'h41452456, 32'hc20a1eeb, 32'h4201241f, 32'hc294f655};
test_output[8923] = '{32'h4287c6a6};
test_index[8923] = '{1};
test_input[71392:71399] = '{32'h425f7be8, 32'h427371e1, 32'hc27f8e64, 32'hc2a77911, 32'h41d7d0a1, 32'hc2c7856a, 32'h4288c81e, 32'hc1b8ce40};
test_output[8924] = '{32'h4288c81e};
test_index[8924] = '{6};
test_input[71400:71407] = '{32'h42bad0f5, 32'hc280f4b6, 32'h42a9911f, 32'h40ba891d, 32'h4276005a, 32'hc276769e, 32'h425beea7, 32'hc21fb015};
test_output[8925] = '{32'h42bad0f5};
test_index[8925] = '{0};
test_input[71408:71415] = '{32'h3e34738b, 32'h428ac8df, 32'hc23c0774, 32'h40b52f85, 32'hc25a6c58, 32'h425b612d, 32'hc2857fc7, 32'hc1efa0fe};
test_output[8926] = '{32'h428ac8df};
test_index[8926] = '{1};
test_input[71416:71423] = '{32'hc2c2af1b, 32'h40c29513, 32'hc20e2d2c, 32'h42c69fcc, 32'h42a83eac, 32'hc286ac33, 32'h41bda73d, 32'h42797d36};
test_output[8927] = '{32'h42c69fcc};
test_index[8927] = '{3};
test_input[71424:71431] = '{32'hc256e790, 32'h424d0453, 32'hc18f119f, 32'h4255f8f1, 32'h42603437, 32'h42c1b543, 32'hc1e7f6d2, 32'hc2272a07};
test_output[8928] = '{32'h42c1b543};
test_index[8928] = '{5};
test_input[71432:71439] = '{32'h42af1025, 32'h42908d11, 32'h41c92b36, 32'h42257b72, 32'h423bed4a, 32'hc20bf257, 32'hc2c5e7e6, 32'h413455c5};
test_output[8929] = '{32'h42af1025};
test_index[8929] = '{0};
test_input[71440:71447] = '{32'hc292cf24, 32'hc2924c0d, 32'h42c49fb5, 32'h42bc424a, 32'hc255e678, 32'h429de5d2, 32'h4282f4bc, 32'h42bd489b};
test_output[8930] = '{32'h42c49fb5};
test_index[8930] = '{2};
test_input[71448:71455] = '{32'h420c1e29, 32'hc2c6aacd, 32'h4263517e, 32'hc2c5e6ac, 32'h419e6650, 32'h41d43e45, 32'h4227fc67, 32'hc204c8c5};
test_output[8931] = '{32'h4263517e};
test_index[8931] = '{2};
test_input[71456:71463] = '{32'h424546fc, 32'hc21d11e3, 32'h42c452d1, 32'h4275ab7f, 32'h41896368, 32'h4280db80, 32'hc22a87a1, 32'hc2a26d0b};
test_output[8932] = '{32'h42c452d1};
test_index[8932] = '{2};
test_input[71464:71471] = '{32'hc29d894b, 32'h4151c88f, 32'h42a21908, 32'hc233ba96, 32'hc2204573, 32'hc2c0edcf, 32'h4258ccbf, 32'h42b75465};
test_output[8933] = '{32'h42b75465};
test_index[8933] = '{7};
test_input[71472:71479] = '{32'hc0dfa7f6, 32'h40bef430, 32'hc22e6122, 32'h42b29319, 32'hc26b812c, 32'hc05650c4, 32'h412c7f53, 32'h42b1d0f3};
test_output[8934] = '{32'h42b29319};
test_index[8934] = '{3};
test_input[71480:71487] = '{32'hc2be8639, 32'h3ee6d0e6, 32'hc2c4ff11, 32'h424daf12, 32'hc29e4b5f, 32'hc2a4fb74, 32'hc24a7f5e, 32'h42aef69b};
test_output[8935] = '{32'h42aef69b};
test_index[8935] = '{7};
test_input[71488:71495] = '{32'h4273de35, 32'hc270f34a, 32'hc2b64224, 32'h42450a2d, 32'h41ed462b, 32'h42878d9e, 32'h4195ab48, 32'hc277a9f9};
test_output[8936] = '{32'h42878d9e};
test_index[8936] = '{5};
test_input[71496:71503] = '{32'h41e35154, 32'h41c52453, 32'h42831d62, 32'h423640ca, 32'h42908559, 32'hc2430e5a, 32'h42196434, 32'hc1cc3a4f};
test_output[8937] = '{32'h42908559};
test_index[8937] = '{4};
test_input[71504:71511] = '{32'hc228cd2e, 32'h41a36eb0, 32'hc2c6863c, 32'hc1bd8a9b, 32'h42312e9a, 32'hc2c7011c, 32'hc2a1626f, 32'hc23395e0};
test_output[8938] = '{32'h42312e9a};
test_index[8938] = '{4};
test_input[71512:71519] = '{32'h3dea343d, 32'h42c35e10, 32'h41d3aab9, 32'h4295eabb, 32'h4188f139, 32'h4245d8e7, 32'h4250c09f, 32'hc1d3ba66};
test_output[8939] = '{32'h42c35e10};
test_index[8939] = '{1};
test_input[71520:71527] = '{32'hc27dd080, 32'hc201ed8a, 32'h429d1ad9, 32'h42736b66, 32'hc1c89570, 32'hc1ca3849, 32'hc0d7f521, 32'hc22e82b8};
test_output[8940] = '{32'h429d1ad9};
test_index[8940] = '{2};
test_input[71528:71535] = '{32'hc281a29f, 32'hc29d055d, 32'hc22f13ab, 32'hc2c5a564, 32'hc26db325, 32'h4288810e, 32'hc259bfb3, 32'h41bd3433};
test_output[8941] = '{32'h4288810e};
test_index[8941] = '{5};
test_input[71536:71543] = '{32'hc27baa8d, 32'h429ecc7f, 32'hc0afa813, 32'h42a735f7, 32'hc21c599b, 32'h4239be53, 32'hc288918c, 32'hc2b40e7d};
test_output[8942] = '{32'h42a735f7};
test_index[8942] = '{3};
test_input[71544:71551] = '{32'hc1a2ec9f, 32'h423ef3dd, 32'hc1a95515, 32'hc2473751, 32'h41811eb0, 32'hc18de373, 32'hc265398f, 32'h42c2864b};
test_output[8943] = '{32'h42c2864b};
test_index[8943] = '{7};
test_input[71552:71559] = '{32'h42136b21, 32'hc1873020, 32'h42bfc328, 32'h40041e44, 32'hc280f9ad, 32'h426f58bd, 32'hc22e5017, 32'h41659930};
test_output[8944] = '{32'h42bfc328};
test_index[8944] = '{2};
test_input[71560:71567] = '{32'h4294b24f, 32'h4250e203, 32'h412e3438, 32'h423230d6, 32'h41c758eb, 32'h418014c8, 32'h42a52b3d, 32'hc129a660};
test_output[8945] = '{32'h42a52b3d};
test_index[8945] = '{6};
test_input[71568:71575] = '{32'h41d383b1, 32'h42c35e9b, 32'hc29181aa, 32'h42c1da08, 32'h42b6c13d, 32'hc28e7b8a, 32'hc121025e, 32'h41b40535};
test_output[8946] = '{32'h42c35e9b};
test_index[8946] = '{1};
test_input[71576:71583] = '{32'h4247f7f1, 32'hc1a35d10, 32'hc2261316, 32'hc2c142de, 32'hc28cf24c, 32'hc24095b9, 32'hc291fdb5, 32'h4288cfe5};
test_output[8947] = '{32'h4288cfe5};
test_index[8947] = '{7};
test_input[71584:71591] = '{32'h427cfbd6, 32'hc15492c7, 32'hc24f5992, 32'h41bbece6, 32'hc2b089d1, 32'h413b177a, 32'hc26cf6eb, 32'h427a682c};
test_output[8948] = '{32'h427cfbd6};
test_index[8948] = '{0};
test_input[71592:71599] = '{32'h4278a6bc, 32'hc2442f9f, 32'h413394dc, 32'h4263e9e4, 32'h42c11930, 32'h427b883c, 32'hc28f69e1, 32'h41d48329};
test_output[8949] = '{32'h42c11930};
test_index[8949] = '{4};
test_input[71600:71607] = '{32'hc1819785, 32'hc0411f15, 32'h429de6be, 32'h42439987, 32'h428faf77, 32'hc2c471b7, 32'h42147b4c, 32'h4242487b};
test_output[8950] = '{32'h429de6be};
test_index[8950] = '{2};
test_input[71608:71615] = '{32'hc2881400, 32'h4287c24b, 32'h428fb5d7, 32'hc1f8c353, 32'hc28a1309, 32'hc27998ce, 32'h42aaeaa9, 32'h40e31175};
test_output[8951] = '{32'h42aaeaa9};
test_index[8951] = '{6};
test_input[71616:71623] = '{32'h4165e3dd, 32'hc006bd7a, 32'hc26db68e, 32'hc2238dfd, 32'h420106a0, 32'h41c2bc3d, 32'h420bf538, 32'h420a17ea};
test_output[8952] = '{32'h420bf538};
test_index[8952] = '{6};
test_input[71624:71631] = '{32'hc226e6c7, 32'hc1a6e0fc, 32'hc2aaf458, 32'hc24802bc, 32'h4252fef7, 32'hc270d987, 32'h41931498, 32'h427eb187};
test_output[8953] = '{32'h427eb187};
test_index[8953] = '{7};
test_input[71632:71639] = '{32'h42743fdc, 32'hbd9bc2ce, 32'hc2b2fb13, 32'hc22f372a, 32'hc205dede, 32'hc2822865, 32'hc291de74, 32'hc1973a4c};
test_output[8954] = '{32'h42743fdc};
test_index[8954] = '{0};
test_input[71640:71647] = '{32'hc2c0ab23, 32'h42b5ca3e, 32'hc1a514b8, 32'hc238ebca, 32'h42860701, 32'h42363b39, 32'h41743ff5, 32'h428583e9};
test_output[8955] = '{32'h42b5ca3e};
test_index[8955] = '{1};
test_input[71648:71655] = '{32'hc2a73c71, 32'h422bc628, 32'h427ce642, 32'hc1aa2283, 32'hc1a2b011, 32'h4245bf92, 32'h42c06816, 32'hc1bdeb9d};
test_output[8956] = '{32'h42c06816};
test_index[8956] = '{6};
test_input[71656:71663] = '{32'hc1ff5855, 32'h42807bd1, 32'hc1e4651f, 32'hc2a6bf36, 32'hc290f287, 32'h4208fba5, 32'h42319186, 32'hc2ac524a};
test_output[8957] = '{32'h42807bd1};
test_index[8957] = '{1};
test_input[71664:71671] = '{32'hc2087c52, 32'h42783e03, 32'h4182212b, 32'hbe8d635f, 32'hc2b84727, 32'h423d9504, 32'hc236f452, 32'hc11e8003};
test_output[8958] = '{32'h42783e03};
test_index[8958] = '{1};
test_input[71672:71679] = '{32'h420cf409, 32'h41345b3a, 32'hc278ad47, 32'h4081f0ba, 32'hc257beff, 32'hc2c282d6, 32'hbf72b5cf, 32'h42bc7cb1};
test_output[8959] = '{32'h42bc7cb1};
test_index[8959] = '{7};
test_input[71680:71687] = '{32'hc2782ad8, 32'hc2bd3fb3, 32'hc2c53660, 32'hc27e1859, 32'h42bf97fa, 32'hc1fc4bfb, 32'h42110f6e, 32'h429793cd};
test_output[8960] = '{32'h42bf97fa};
test_index[8960] = '{4};
test_input[71688:71695] = '{32'h428daf15, 32'hc227b091, 32'h42a41ad2, 32'hc18e3a20, 32'h42c774df, 32'hc1c8b4ea, 32'hc22a8389, 32'h42c7e97b};
test_output[8961] = '{32'h42c7e97b};
test_index[8961] = '{7};
test_input[71696:71703] = '{32'h42b14275, 32'hc2205e1b, 32'hc25a1e48, 32'h42876f93, 32'hc1fccb90, 32'h41753abe, 32'hc24a63ab, 32'h4272f9ce};
test_output[8962] = '{32'h42b14275};
test_index[8962] = '{0};
test_input[71704:71711] = '{32'h42ab5ce3, 32'h42889d71, 32'hc289d7c3, 32'hc2559537, 32'hc28876f6, 32'hc29242ff, 32'hc23004f1, 32'hc2037704};
test_output[8963] = '{32'h42ab5ce3};
test_index[8963] = '{0};
test_input[71712:71719] = '{32'hc1f6ebcb, 32'h41367e98, 32'hc1b291b1, 32'h41a99a18, 32'h3fdb8d5b, 32'hc298b6fa, 32'h42b3b57f, 32'hc27033c1};
test_output[8964] = '{32'h42b3b57f};
test_index[8964] = '{6};
test_input[71720:71727] = '{32'hc279a3a9, 32'h42147ec0, 32'hc2846169, 32'hbf5cfce9, 32'h42a5c796, 32'h42159f58, 32'hc2ac0f53, 32'h41acf095};
test_output[8965] = '{32'h42a5c796};
test_index[8965] = '{4};
test_input[71728:71735] = '{32'hc1385453, 32'hc2bda6fb, 32'h42a11206, 32'hc1e2dac1, 32'h4108c88e, 32'hc29be17d, 32'h41aa83e7, 32'h41ebbdaa};
test_output[8966] = '{32'h42a11206};
test_index[8966] = '{2};
test_input[71736:71743] = '{32'h42921c44, 32'h41fc0e7c, 32'h42815f14, 32'h4208f3af, 32'h427e16ce, 32'h42a18f26, 32'hc195acad, 32'h42c1d01f};
test_output[8967] = '{32'h42c1d01f};
test_index[8967] = '{7};
test_input[71744:71751] = '{32'hc237f999, 32'h42a9779a, 32'hc0fe80b6, 32'h41600b51, 32'hc275ef94, 32'hc22abd9c, 32'h42858fbb, 32'hc2371b2c};
test_output[8968] = '{32'h42a9779a};
test_index[8968] = '{1};
test_input[71752:71759] = '{32'hc1dca410, 32'h4216a695, 32'hc28c562b, 32'h42457722, 32'h42817949, 32'h41c5a7fa, 32'hc2beb4f0, 32'h42c52c15};
test_output[8969] = '{32'h42c52c15};
test_index[8969] = '{7};
test_input[71760:71767] = '{32'h429d8e13, 32'hc15ed02c, 32'hc28390dc, 32'h42a6b51c, 32'h421e6c4c, 32'h40dfce00, 32'hc272e94b, 32'hc24bdc86};
test_output[8970] = '{32'h42a6b51c};
test_index[8970] = '{3};
test_input[71768:71775] = '{32'h4233d6a6, 32'hc1eb0a95, 32'h4220cf20, 32'hc19a1106, 32'h42b358cd, 32'h42352d6c, 32'hc23a3311, 32'h426999ea};
test_output[8971] = '{32'h42b358cd};
test_index[8971] = '{4};
test_input[71776:71783] = '{32'hc298861b, 32'h42934e6e, 32'hc2ad2584, 32'hc0e088b8, 32'h419caee5, 32'hc2346fce, 32'h41f96cf1, 32'hc24eb4aa};
test_output[8972] = '{32'h42934e6e};
test_index[8972] = '{1};
test_input[71784:71791] = '{32'h4059ce54, 32'hbfc6c8aa, 32'h3d9a1636, 32'hc2a47fcc, 32'h41f174f9, 32'h42b8b2cd, 32'hc2783504, 32'hc2a9e3ab};
test_output[8973] = '{32'h42b8b2cd};
test_index[8973] = '{5};
test_input[71792:71799] = '{32'hc14acbae, 32'hc20b5d77, 32'h4296131b, 32'h42778e47, 32'h4224eea0, 32'hc1648c40, 32'h42bcd749, 32'hc285cf88};
test_output[8974] = '{32'h42bcd749};
test_index[8974] = '{6};
test_input[71800:71807] = '{32'h42847d26, 32'hc20cd63a, 32'hc1911ec6, 32'h40d8ec4d, 32'h419141ff, 32'hc2b046a4, 32'h41fb67e9, 32'h3ff45e64};
test_output[8975] = '{32'h42847d26};
test_index[8975] = '{0};
test_input[71808:71815] = '{32'h3f4be824, 32'hc2b2bbd0, 32'hc231d8c7, 32'h423a26f5, 32'hc26f6e53, 32'h429d3fd3, 32'h40c66b76, 32'h41e73a01};
test_output[8976] = '{32'h429d3fd3};
test_index[8976] = '{5};
test_input[71816:71823] = '{32'hc2b7d44f, 32'hc297b3c5, 32'hc26da30d, 32'h4288e37f, 32'hc2c62e30, 32'hc28b5c3d, 32'hc2afe41b, 32'h42271237};
test_output[8977] = '{32'h4288e37f};
test_index[8977] = '{3};
test_input[71824:71831] = '{32'hc2b7a5ad, 32'h424a86ad, 32'hc1882cb8, 32'hc24f53b8, 32'h42c5e4e8, 32'h42a78a77, 32'h40c2e387, 32'hc1e5c28a};
test_output[8978] = '{32'h42c5e4e8};
test_index[8978] = '{4};
test_input[71832:71839] = '{32'h3fb34a25, 32'hc282f865, 32'hc2ae165c, 32'hc0436aa1, 32'h42908f56, 32'hc295f502, 32'h41dec754, 32'hc197676c};
test_output[8979] = '{32'h42908f56};
test_index[8979] = '{4};
test_input[71840:71847] = '{32'hc176199d, 32'hc1a76421, 32'h4273c4b5, 32'hbf796dd6, 32'h42783480, 32'h42197d48, 32'h41e6d37d, 32'h411a0bb5};
test_output[8980] = '{32'h42783480};
test_index[8980] = '{4};
test_input[71848:71855] = '{32'h4284fae5, 32'h4251430a, 32'h426c0fb9, 32'hc2556dfc, 32'h423c7312, 32'hbf2b1d67, 32'hc1c5527c, 32'hc27b7383};
test_output[8981] = '{32'h4284fae5};
test_index[8981] = '{0};
test_input[71856:71863] = '{32'hc1b14601, 32'hc12fc791, 32'hc0520302, 32'h42a29338, 32'hc2908e9d, 32'hc1e77db4, 32'hc21050c0, 32'hc1ad8757};
test_output[8982] = '{32'h42a29338};
test_index[8982] = '{3};
test_input[71864:71871] = '{32'hbeba47ea, 32'h42a27d25, 32'hbe893c06, 32'hc2a08185, 32'hc1556b70, 32'h415a8f09, 32'hc28d0a77, 32'hc28c1755};
test_output[8983] = '{32'h42a27d25};
test_index[8983] = '{1};
test_input[71872:71879] = '{32'h42362f7d, 32'h41cd8c3d, 32'hc2655faf, 32'hc1c08f34, 32'hc25404d5, 32'h4263cb8b, 32'h419d2620, 32'h41624c6e};
test_output[8984] = '{32'h4263cb8b};
test_index[8984] = '{5};
test_input[71880:71887] = '{32'h4280aa18, 32'hc2bc6498, 32'h4105b31e, 32'hc22c4244, 32'hc2b9fb18, 32'h42086f3b, 32'h42c78b83, 32'hc2abecc2};
test_output[8985] = '{32'h42c78b83};
test_index[8985] = '{6};
test_input[71888:71895] = '{32'h4216e8f0, 32'h3ffe21f8, 32'h420c46a8, 32'hc242c192, 32'hc2acd2f4, 32'hc2a28e36, 32'h41b1c2cf, 32'h424633af};
test_output[8986] = '{32'h424633af};
test_index[8986] = '{7};
test_input[71896:71903] = '{32'hc2bf3142, 32'h42310b2e, 32'hc2b0b7f4, 32'h3fd1d685, 32'hc160d76e, 32'h4224d87a, 32'hc2a14747, 32'h42258be1};
test_output[8987] = '{32'h42310b2e};
test_index[8987] = '{1};
test_input[71904:71911] = '{32'h42bc9f7c, 32'h4285d38c, 32'h4253c892, 32'hc1293a0f, 32'h427cbd0e, 32'hc28b9a03, 32'h428fb66a, 32'h416555c5};
test_output[8988] = '{32'h42bc9f7c};
test_index[8988] = '{0};
test_input[71912:71919] = '{32'h421d3c16, 32'h42aae21f, 32'hc1be01c2, 32'hc139ef98, 32'hc1a77642, 32'hc19d33c5, 32'hc2c12447, 32'h40a5d890};
test_output[8989] = '{32'h42aae21f};
test_index[8989] = '{1};
test_input[71920:71927] = '{32'hc284ba76, 32'h42a41362, 32'hc20dd545, 32'hc23cbab7, 32'h422af716, 32'h41dd4591, 32'hc1a2539b, 32'h42991836};
test_output[8990] = '{32'h42a41362};
test_index[8990] = '{1};
test_input[71928:71935] = '{32'h42b62ebb, 32'hc205465c, 32'hc0cd4167, 32'hc13d94df, 32'h422886ab, 32'h42b7bfcc, 32'hc226e11f, 32'h425eabdb};
test_output[8991] = '{32'h42b7bfcc};
test_index[8991] = '{5};
test_input[71936:71943] = '{32'h429eb1d1, 32'h420abdf1, 32'h40eff370, 32'hc053e334, 32'hc25564b9, 32'hc232fe40, 32'h420bd936, 32'h4238f188};
test_output[8992] = '{32'h429eb1d1};
test_index[8992] = '{0};
test_input[71944:71951] = '{32'h42944560, 32'hc2960274, 32'h4260b16d, 32'hc27e8934, 32'hc295f842, 32'h42b9af2a, 32'h4286f25e, 32'h42922cfe};
test_output[8993] = '{32'h42b9af2a};
test_index[8993] = '{5};
test_input[71952:71959] = '{32'h42884fac, 32'h424642be, 32'hc1a3f0c8, 32'hc0ad0b6e, 32'hc29d477c, 32'hc296863f, 32'h4232ce37, 32'hc1a54ad1};
test_output[8994] = '{32'h42884fac};
test_index[8994] = '{0};
test_input[71960:71967] = '{32'hc11ccc84, 32'h41e0a37a, 32'hc1359c3c, 32'hc08a5167, 32'hc2c14ca5, 32'h428407c4, 32'h4224400a, 32'hc2ac95d3};
test_output[8995] = '{32'h428407c4};
test_index[8995] = '{5};
test_input[71968:71975] = '{32'hc2a088dc, 32'hbfbfe593, 32'h40fc59b0, 32'h42a514e6, 32'hc1f5cf59, 32'h429b939d, 32'h422ca2be, 32'h428f92b3};
test_output[8996] = '{32'h42a514e6};
test_index[8996] = '{3};
test_input[71976:71983] = '{32'hc246b3a8, 32'h4227e2a3, 32'hc1158658, 32'h42362fb3, 32'h4289f9ab, 32'h422c397e, 32'h4189650d, 32'hc005f97f};
test_output[8997] = '{32'h4289f9ab};
test_index[8997] = '{4};
test_input[71984:71991] = '{32'h42b21f3b, 32'h423468ac, 32'h42b19c0b, 32'hc23f07e1, 32'h42241922, 32'hc10c283e, 32'h42609e4c, 32'h41abdc8a};
test_output[8998] = '{32'h42b21f3b};
test_index[8998] = '{0};
test_input[71992:71999] = '{32'hc254d1bd, 32'h424f607c, 32'hc284c1df, 32'hc2a6a459, 32'h4274c52b, 32'hc2761e70, 32'hc28fd267, 32'h42414e86};
test_output[8999] = '{32'h4274c52b};
test_index[8999] = '{4};
test_input[72000:72007] = '{32'h40fa1df1, 32'h4295fd89, 32'hc2851fec, 32'h4189b069, 32'h425b4db5, 32'hc0ca4791, 32'hc2b0fbc5, 32'h4248cee3};
test_output[9000] = '{32'h4295fd89};
test_index[9000] = '{1};
test_input[72008:72015] = '{32'h422a7bed, 32'h429add51, 32'hc2a1cfcc, 32'hc192916a, 32'hc14fbf4a, 32'h427eccc9, 32'hc1f664c7, 32'hc28d3254};
test_output[9001] = '{32'h429add51};
test_index[9001] = '{1};
test_input[72016:72023] = '{32'hc1fed67e, 32'hc2bb4e9d, 32'h410dd4bc, 32'hc22ac5f5, 32'hc1e35858, 32'h42c43b61, 32'hc2820f7d, 32'h41df5622};
test_output[9002] = '{32'h42c43b61};
test_index[9002] = '{5};
test_input[72024:72031] = '{32'hc29c2a20, 32'h429e888a, 32'h4297d669, 32'h41e7477e, 32'hc290049d, 32'h4200fd9c, 32'h415c1b74, 32'h42ba7e0d};
test_output[9003] = '{32'h42ba7e0d};
test_index[9003] = '{7};
test_input[72032:72039] = '{32'h40aa565b, 32'h3fd68828, 32'h42807cb1, 32'hc24db0e8, 32'h41bb2f70, 32'h418e8adf, 32'h41f24a37, 32'hc0c9a541};
test_output[9004] = '{32'h42807cb1};
test_index[9004] = '{2};
test_input[72040:72047] = '{32'hc26e7d63, 32'h41f98703, 32'hc25b419c, 32'hc1a815bc, 32'h41daf197, 32'hc13bec80, 32'hc2c5e5db, 32'h4216bdb2};
test_output[9005] = '{32'h4216bdb2};
test_index[9005] = '{7};
test_input[72048:72055] = '{32'hc2a9ddc1, 32'hc10776f0, 32'h3f3c1f1f, 32'h425385fb, 32'h420ddce7, 32'h4239d0c1, 32'h422d57ca, 32'h42b12719};
test_output[9006] = '{32'h42b12719};
test_index[9006] = '{7};
test_input[72056:72063] = '{32'hc24ead2a, 32'hc0c6a25b, 32'hc1fd81c1, 32'hc02d4b3a, 32'hc1bb1364, 32'h422dc5ca, 32'h42bb9f04, 32'hc2b25f57};
test_output[9007] = '{32'h42bb9f04};
test_index[9007] = '{6};
test_input[72064:72071] = '{32'hc2c5e8e2, 32'h42501193, 32'h42b26f0e, 32'hc06ded31, 32'hc2a30845, 32'h40d21294, 32'hc245e6be, 32'h423afbf2};
test_output[9008] = '{32'h42b26f0e};
test_index[9008] = '{2};
test_input[72072:72079] = '{32'hc280392a, 32'h428bce4a, 32'hc20778f2, 32'hc2b7ee2e, 32'hc2b4f3cc, 32'h42a19b18, 32'hc2aec6d4, 32'hc2bb2365};
test_output[9009] = '{32'h42a19b18};
test_index[9009] = '{5};
test_input[72080:72087] = '{32'hbf6e9ec9, 32'h4021b38b, 32'hc19ee735, 32'hc24dfe8e, 32'h4279670a, 32'hc21efa0b, 32'hc1fd6b93, 32'hc20d9922};
test_output[9010] = '{32'h4279670a};
test_index[9010] = '{4};
test_input[72088:72095] = '{32'hc2bb56bf, 32'h41a94080, 32'hc1c209fa, 32'hc23b81d2, 32'h4218a7d4, 32'hc25e962b, 32'hc1faa03f, 32'hc2653f65};
test_output[9011] = '{32'h4218a7d4};
test_index[9011] = '{4};
test_input[72096:72103] = '{32'hc0a0fdc6, 32'h424378af, 32'h428f48cd, 32'h419b5fd7, 32'hc2865d10, 32'h41e40039, 32'h41902343, 32'hc273898b};
test_output[9012] = '{32'h428f48cd};
test_index[9012] = '{2};
test_input[72104:72111] = '{32'hc1b57240, 32'hc244304c, 32'hc290264a, 32'hc2c19092, 32'hc10c9adf, 32'hc285e785, 32'h42107c7b, 32'hc121c427};
test_output[9013] = '{32'h42107c7b};
test_index[9013] = '{6};
test_input[72112:72119] = '{32'h4295e764, 32'hc2af79e3, 32'hc17d24e0, 32'hc2ab8940, 32'h4290e948, 32'hc22aaffc, 32'hc242544e, 32'hc1a5fcf1};
test_output[9014] = '{32'h4295e764};
test_index[9014] = '{0};
test_input[72120:72127] = '{32'h42947b30, 32'h4280f91d, 32'hc12ce345, 32'hc2c3a560, 32'h4290f084, 32'h41c9cdc9, 32'h41e2f7b9, 32'hc28272d7};
test_output[9015] = '{32'h42947b30};
test_index[9015] = '{0};
test_input[72128:72135] = '{32'hc0f3413a, 32'h41af2d20, 32'h41f31af9, 32'hc28c7278, 32'hc2ab7068, 32'h42b3b30a, 32'hc1309494, 32'h423cee72};
test_output[9016] = '{32'h42b3b30a};
test_index[9016] = '{5};
test_input[72136:72143] = '{32'hc29321fd, 32'hc29191d4, 32'hc21b7396, 32'h428b235e, 32'h4237c1ec, 32'hc1fe124c, 32'h42ad9e41, 32'h4275edf3};
test_output[9017] = '{32'h42ad9e41};
test_index[9017] = '{6};
test_input[72144:72151] = '{32'hc2061869, 32'h41e59f5f, 32'hc23c2631, 32'hc21f58d4, 32'h423ac811, 32'hc21c428d, 32'h4257926e, 32'h428ad18e};
test_output[9018] = '{32'h428ad18e};
test_index[9018] = '{7};
test_input[72152:72159] = '{32'h42236d32, 32'h4282dedb, 32'hc152dcf5, 32'h41d9452a, 32'hc2bead4d, 32'h428ddec9, 32'hbf86163f, 32'hc11b764a};
test_output[9019] = '{32'h428ddec9};
test_index[9019] = '{5};
test_input[72160:72167] = '{32'hc2805357, 32'hc25c4e08, 32'hc16ea3b7, 32'h41eb03e5, 32'h4125452a, 32'hc28e71ee, 32'hc2a4efbf, 32'h42b3477e};
test_output[9020] = '{32'h42b3477e};
test_index[9020] = '{7};
test_input[72168:72175] = '{32'hc208aa90, 32'h42c735ef, 32'h42469b4f, 32'h417adf4b, 32'h4216b583, 32'hbee97831, 32'hc294f718, 32'h40f1e443};
test_output[9021] = '{32'h42c735ef};
test_index[9021] = '{1};
test_input[72176:72183] = '{32'hc227bdd3, 32'hc253b98e, 32'hc29f58f0, 32'h40e3dd5c, 32'hc2c37efb, 32'h4107b1c4, 32'hc209b5a7, 32'h421b7e3b};
test_output[9022] = '{32'h421b7e3b};
test_index[9022] = '{7};
test_input[72184:72191] = '{32'hc2c5b9a5, 32'hc2a7227b, 32'hbfc59250, 32'hc278753d, 32'hbff6ac92, 32'h41ad2c97, 32'h42b0224c, 32'hc2623034};
test_output[9023] = '{32'h42b0224c};
test_index[9023] = '{6};
test_input[72192:72199] = '{32'hc21002a2, 32'h3e1c9cf9, 32'hc252618e, 32'h414b4ef4, 32'hbf6fc6ad, 32'hc217829b, 32'h42b37d04, 32'hc21c5fe7};
test_output[9024] = '{32'h42b37d04};
test_index[9024] = '{6};
test_input[72200:72207] = '{32'h42798624, 32'hc26fe9fc, 32'h42918fb5, 32'hc1a9cfc1, 32'h42a64a4e, 32'hc21a249f, 32'h41824a4b, 32'h42115cc2};
test_output[9025] = '{32'h42a64a4e};
test_index[9025] = '{4};
test_input[72208:72215] = '{32'hbf8b3b13, 32'hc22ecd66, 32'h41a323bc, 32'h427e4562, 32'h425ac214, 32'hc2c60dc4, 32'h42b7eac4, 32'hc28d2791};
test_output[9026] = '{32'h42b7eac4};
test_index[9026] = '{6};
test_input[72216:72223] = '{32'h428601c7, 32'hc2be2965, 32'hc2ac4352, 32'h4283e9ce, 32'h42240115, 32'hc18da343, 32'h42b7ff64, 32'hc2868ccb};
test_output[9027] = '{32'h42b7ff64};
test_index[9027] = '{6};
test_input[72224:72231] = '{32'h429a50c8, 32'h4296cb08, 32'hc19bb830, 32'h423cc18a, 32'hc2433003, 32'h422aca3e, 32'h426873e8, 32'h41da954d};
test_output[9028] = '{32'h429a50c8};
test_index[9028] = '{0};
test_input[72232:72239] = '{32'h425b4d66, 32'hc2c02c7c, 32'hc1663d3d, 32'hc298412c, 32'h4288f514, 32'hc245637a, 32'hc27dc177, 32'h410bd726};
test_output[9029] = '{32'h4288f514};
test_index[9029] = '{4};
test_input[72240:72247] = '{32'h41b714b4, 32'h4299788d, 32'h42641c61, 32'h42a90d1f, 32'hc2ad8f2c, 32'hc1da7f4f, 32'h418ade60, 32'h42883a58};
test_output[9030] = '{32'h42a90d1f};
test_index[9030] = '{3};
test_input[72248:72255] = '{32'h41d1dd31, 32'hc2bfdbe7, 32'hc202cf0a, 32'h424039e9, 32'h42bcd4fa, 32'h416ace49, 32'h42ae234b, 32'hc1f5c6c5};
test_output[9031] = '{32'h42bcd4fa};
test_index[9031] = '{4};
test_input[72256:72263] = '{32'h42a2aa82, 32'hc26cc07e, 32'h428301c1, 32'h41dc3d49, 32'hc293e320, 32'hc120a3d7, 32'hc18f3d81, 32'hc2a7b110};
test_output[9032] = '{32'h42a2aa82};
test_index[9032] = '{0};
test_input[72264:72271] = '{32'hc0e12da3, 32'hc283705e, 32'h406a4b58, 32'hc29985bf, 32'hc13425fa, 32'hc2b86c6b, 32'hc23c1568, 32'hc185b53a};
test_output[9033] = '{32'h406a4b58};
test_index[9033] = '{2};
test_input[72272:72279] = '{32'hc1a71265, 32'hc244966a, 32'hc21be138, 32'hc2a5da16, 32'h42aae84b, 32'h420e68f1, 32'h41050925, 32'hc283fd45};
test_output[9034] = '{32'h42aae84b};
test_index[9034] = '{4};
test_input[72280:72287] = '{32'h429d727f, 32'h40673265, 32'h428b31e2, 32'hc240fcc1, 32'h422cd4f5, 32'h42bc13f3, 32'hc26ed174, 32'h42a119e4};
test_output[9035] = '{32'h42bc13f3};
test_index[9035] = '{5};
test_input[72288:72295] = '{32'h425a973d, 32'h419c260f, 32'h41b0d7b2, 32'h41929772, 32'hc285ace5, 32'hc14b1a37, 32'h428f95eb, 32'hc2965468};
test_output[9036] = '{32'h428f95eb};
test_index[9036] = '{6};
test_input[72296:72303] = '{32'h42a0143a, 32'h4258c6b3, 32'h42698fb4, 32'hc28ba1ce, 32'h428a71f2, 32'hc0c3f0fe, 32'hbfbd95aa, 32'h424e9a4e};
test_output[9037] = '{32'h42a0143a};
test_index[9037] = '{0};
test_input[72304:72311] = '{32'hc2a8214c, 32'h41bb4639, 32'hc2017bf8, 32'hc1b36bab, 32'hc26830c1, 32'h42995cc2, 32'h42839ea7, 32'h4245bfb8};
test_output[9038] = '{32'h42995cc2};
test_index[9038] = '{5};
test_input[72312:72319] = '{32'h4284f56f, 32'hc225c61f, 32'h42427b73, 32'hc2c1339b, 32'h42acf57f, 32'hc17e3b5c, 32'hc2b06744, 32'h427ba39a};
test_output[9039] = '{32'h42acf57f};
test_index[9039] = '{4};
test_input[72320:72327] = '{32'h4299a77f, 32'h4250ef9f, 32'hc20f5453, 32'h42c4bcc7, 32'h426db18f, 32'hc21af605, 32'h42ac754c, 32'hc2a75455};
test_output[9040] = '{32'h42c4bcc7};
test_index[9040] = '{3};
test_input[72328:72335] = '{32'h42730f1a, 32'h4259d11a, 32'hc2b8db94, 32'hc2ab6413, 32'h4215fd1d, 32'h41d849fa, 32'h42b2d202, 32'h41d1bb54};
test_output[9041] = '{32'h42b2d202};
test_index[9041] = '{6};
test_input[72336:72343] = '{32'h427d632d, 32'hc11e019a, 32'hc2924241, 32'h4202034d, 32'h42ab0431, 32'hc279c591, 32'h42458602, 32'h42278d89};
test_output[9042] = '{32'h42ab0431};
test_index[9042] = '{4};
test_input[72344:72351] = '{32'hc1cf1ca8, 32'h421f004c, 32'hc1954e10, 32'h4287083c, 32'h41c5ddf8, 32'hc0e986f1, 32'hc1d4097e, 32'h4266cf85};
test_output[9043] = '{32'h4287083c};
test_index[9043] = '{3};
test_input[72352:72359] = '{32'hc2930a09, 32'hc2abda78, 32'hc248ff2a, 32'h421c6854, 32'h41941cd2, 32'h41b9aeee, 32'h429238bf, 32'h429bafd1};
test_output[9044] = '{32'h429bafd1};
test_index[9044] = '{7};
test_input[72360:72367] = '{32'h42935783, 32'hc12c386c, 32'h42ace5db, 32'hc28176b3, 32'h4286d0a8, 32'hc24abdc0, 32'hc2923a9e, 32'h423cb966};
test_output[9045] = '{32'h42ace5db};
test_index[9045] = '{2};
test_input[72368:72375] = '{32'hbea1aea2, 32'hc200a583, 32'h42c18bcb, 32'h41835428, 32'hc2c170b3, 32'h40f0489a, 32'h4263e8c6, 32'h426d9600};
test_output[9046] = '{32'h42c18bcb};
test_index[9046] = '{2};
test_input[72376:72383] = '{32'h42b82902, 32'hc17daf84, 32'hc1e3e1b0, 32'h42012d98, 32'hc1c59e83, 32'hc254c65d, 32'h41ba149e, 32'hc1ba940b};
test_output[9047] = '{32'h42b82902};
test_index[9047] = '{0};
test_input[72384:72391] = '{32'h424f3298, 32'h42480c86, 32'hc2bc9e55, 32'hc231e4c2, 32'h41f82641, 32'h4289d1e7, 32'h41ea7835, 32'hc2a41b29};
test_output[9048] = '{32'h4289d1e7};
test_index[9048] = '{5};
test_input[72392:72399] = '{32'hc2b82a8a, 32'hc27a7148, 32'h428e897f, 32'h4286b498, 32'hc2b6bbed, 32'h3f857484, 32'h4138c60c, 32'h4294b1bc};
test_output[9049] = '{32'h4294b1bc};
test_index[9049] = '{7};
test_input[72400:72407] = '{32'hc2962226, 32'hc2a9a6e5, 32'h4200bc4e, 32'h4247da91, 32'h429ac796, 32'hc2a3d61f, 32'hc20c0687, 32'hc2acd767};
test_output[9050] = '{32'h429ac796};
test_index[9050] = '{4};
test_input[72408:72415] = '{32'h42411775, 32'hc26b195e, 32'hc17ee13b, 32'h42b6167f, 32'h428bb3fb, 32'h4135066e, 32'h424ce64f, 32'h424328fc};
test_output[9051] = '{32'h42b6167f};
test_index[9051] = '{3};
test_input[72416:72423] = '{32'hc2145901, 32'h426e89fc, 32'hc2c2d023, 32'hc238c422, 32'hc20f5b76, 32'h42b7cb5e, 32'hc2c074ee, 32'h42acdded};
test_output[9052] = '{32'h42b7cb5e};
test_index[9052] = '{5};
test_input[72424:72431] = '{32'hc2928c91, 32'hc254f138, 32'h421dff84, 32'h428d26a1, 32'hc282a995, 32'h42be2dc2, 32'h42909a79, 32'h42165c0b};
test_output[9053] = '{32'h42be2dc2};
test_index[9053] = '{5};
test_input[72432:72439] = '{32'h42705251, 32'h424097fb, 32'h4188327d, 32'hc2115587, 32'h429721cd, 32'hc286d7a1, 32'hc18f4a9a, 32'hc2039b63};
test_output[9054] = '{32'h429721cd};
test_index[9054] = '{4};
test_input[72440:72447] = '{32'hc20f5fa3, 32'h42716052, 32'h427e77a3, 32'hc2a74bf0, 32'h41e1c0ca, 32'h40d9d30b, 32'hc00926fc, 32'hc1d21632};
test_output[9055] = '{32'h427e77a3};
test_index[9055] = '{2};
test_input[72448:72455] = '{32'hc18dc79f, 32'hc13f442c, 32'hc29a6373, 32'h42221b35, 32'hc1f74c31, 32'h423ec4a2, 32'hc287abdb, 32'hc28a94ea};
test_output[9056] = '{32'h423ec4a2};
test_index[9056] = '{5};
test_input[72456:72463] = '{32'hc255247e, 32'hc002e520, 32'h42722588, 32'hc2c3803c, 32'h423b3040, 32'hc2b24935, 32'h4234b7fa, 32'hc2732468};
test_output[9057] = '{32'h42722588};
test_index[9057] = '{2};
test_input[72464:72471] = '{32'h41fdc39c, 32'hc2a544ca, 32'h414654b3, 32'hc26d8258, 32'hc28e573f, 32'h4174f813, 32'h42105f06, 32'h413e953f};
test_output[9058] = '{32'h42105f06};
test_index[9058] = '{6};
test_input[72472:72479] = '{32'hc1ae534b, 32'h42086d22, 32'hc2aaf9db, 32'h41a01ae1, 32'h42400222, 32'h4241d03d, 32'hc009a1ff, 32'h41b6f311};
test_output[9059] = '{32'h4241d03d};
test_index[9059] = '{5};
test_input[72480:72487] = '{32'h424037e8, 32'h41c79b33, 32'h42a8ac27, 32'h428d0612, 32'hc1b7f8c5, 32'h42717d1c, 32'h420a98bc, 32'h42c11985};
test_output[9060] = '{32'h42c11985};
test_index[9060] = '{7};
test_input[72488:72495] = '{32'hc2b0b325, 32'hc28b56dc, 32'hc2408339, 32'hc22037c4, 32'h42a7ce91, 32'hc11602c3, 32'h4242f8af, 32'hc25a6bf2};
test_output[9061] = '{32'h42a7ce91};
test_index[9061] = '{4};
test_input[72496:72503] = '{32'h42a41309, 32'h42c6910b, 32'hc26320da, 32'hbfa9ac3d, 32'h413baf88, 32'hbf66bbdf, 32'hc2ac7819, 32'h42a60ad7};
test_output[9062] = '{32'h42c6910b};
test_index[9062] = '{1};
test_input[72504:72511] = '{32'hc25f78c6, 32'h428c78ab, 32'h42b71f65, 32'hc2b26a50, 32'hc2a819b6, 32'hc28ecd42, 32'h4208c67e, 32'hc09aea0c};
test_output[9063] = '{32'h42b71f65};
test_index[9063] = '{2};
test_input[72512:72519] = '{32'hc110ba0b, 32'hc1ed9598, 32'hc203b5c7, 32'h428b58c6, 32'h41e8ef20, 32'hc21ef0c1, 32'hc142d472, 32'h4242bd79};
test_output[9064] = '{32'h428b58c6};
test_index[9064] = '{3};
test_input[72520:72527] = '{32'hc0a34256, 32'h425f4f85, 32'hc23b21b1, 32'h42a8e6ba, 32'hc27d947e, 32'hc25f86ca, 32'h418df490, 32'h42b7eeed};
test_output[9065] = '{32'h42b7eeed};
test_index[9065] = '{7};
test_input[72528:72535] = '{32'hc2b8f2ba, 32'h42a1b876, 32'hc0aa3ab6, 32'h42b6e4a0, 32'hc2a3b620, 32'hc221a1d6, 32'hc21868f6, 32'h41a0dfda};
test_output[9066] = '{32'h42b6e4a0};
test_index[9066] = '{3};
test_input[72536:72543] = '{32'h42591732, 32'hc290e8e3, 32'h42c2ae06, 32'hc226f702, 32'h426c5ce4, 32'h42168aa6, 32'hc292244f, 32'hc2acdc38};
test_output[9067] = '{32'h42c2ae06};
test_index[9067] = '{2};
test_input[72544:72551] = '{32'h4148b7d6, 32'h426dbc9c, 32'h40e6ca52, 32'h400c51bd, 32'h415c892c, 32'h418e10ed, 32'h42a00516, 32'hc258911c};
test_output[9068] = '{32'h42a00516};
test_index[9068] = '{6};
test_input[72552:72559] = '{32'h419eccb8, 32'hc29a4766, 32'h40530efa, 32'hc2ab7b63, 32'hc29e7a0d, 32'hc28afe71, 32'hc27d3daf, 32'hc291fdc2};
test_output[9069] = '{32'h419eccb8};
test_index[9069] = '{0};
test_input[72560:72567] = '{32'h428a34ec, 32'h42a61144, 32'hc299a809, 32'hc2c1e0ec, 32'hc127f20e, 32'h42840739, 32'hc1acfeab, 32'h4208b165};
test_output[9070] = '{32'h42a61144};
test_index[9070] = '{1};
test_input[72568:72575] = '{32'hc286ac9d, 32'h41032c7e, 32'hc16c39e9, 32'h428ae796, 32'h40de4dd5, 32'hc2709681, 32'hc2c22332, 32'h429ba3a9};
test_output[9071] = '{32'h429ba3a9};
test_index[9071] = '{7};
test_input[72576:72583] = '{32'h428f07f7, 32'h4229de9f, 32'hc2abae02, 32'h41ff4bda, 32'h4200b734, 32'hc2982c5b, 32'h42ae7b39, 32'hc1baa5b2};
test_output[9072] = '{32'h42ae7b39};
test_index[9072] = '{6};
test_input[72584:72591] = '{32'hc23ba057, 32'h427e8e6f, 32'hc26ecb65, 32'h4209202c, 32'hc2184f3f, 32'hc273a1d3, 32'h422b73f7, 32'hc1bab1ec};
test_output[9073] = '{32'h427e8e6f};
test_index[9073] = '{1};
test_input[72592:72599] = '{32'h4251fa5b, 32'h40834a5c, 32'hc28d2bcb, 32'h427d9239, 32'h42327aa8, 32'hc1a06065, 32'h42ba0432, 32'h4297e128};
test_output[9074] = '{32'h42ba0432};
test_index[9074] = '{6};
test_input[72600:72607] = '{32'h429b7120, 32'hc287c1e3, 32'hc126d732, 32'hc259e5a8, 32'hc0ad9647, 32'hc2553db7, 32'h41a43583, 32'hc192b806};
test_output[9075] = '{32'h429b7120};
test_index[9075] = '{0};
test_input[72608:72615] = '{32'h42be6385, 32'hc24606fa, 32'hc17ef96e, 32'hc2c16c1e, 32'h421e748e, 32'hc2c43d77, 32'h41f38095, 32'hc2b52131};
test_output[9076] = '{32'h42be6385};
test_index[9076] = '{0};
test_input[72616:72623] = '{32'h4268c5bc, 32'h421af760, 32'hc1c47733, 32'hc0cca0f8, 32'h42a1af8e, 32'h42b81847, 32'hc0993fbf, 32'h40d87a96};
test_output[9077] = '{32'h42b81847};
test_index[9077] = '{5};
test_input[72624:72631] = '{32'hc12150de, 32'hc231b879, 32'h428cae59, 32'hc2977bdb, 32'hc0539a8a, 32'hc18a5af8, 32'hc1f3fa52, 32'hc1b4897d};
test_output[9078] = '{32'h428cae59};
test_index[9078] = '{2};
test_input[72632:72639] = '{32'hc1686bdd, 32'h429d5445, 32'hc23101b2, 32'h4261ae74, 32'hc2b9d44b, 32'h42172f34, 32'h41feea8d, 32'hc2b3fcbc};
test_output[9079] = '{32'h429d5445};
test_index[9079] = '{1};
test_input[72640:72647] = '{32'h425f8b78, 32'h41b3e3fd, 32'hc200e06e, 32'hc27c23d3, 32'h41ca2548, 32'hc2517f59, 32'hc10015b0, 32'hc21dda02};
test_output[9080] = '{32'h425f8b78};
test_index[9080] = '{0};
test_input[72648:72655] = '{32'hc1e172a9, 32'h40b99b8c, 32'hc25626d5, 32'h4279df78, 32'hc22c179e, 32'hc2875e60, 32'h425e3c5e, 32'hc0864b78};
test_output[9081] = '{32'h4279df78};
test_index[9081] = '{3};
test_input[72656:72663] = '{32'h42ba6637, 32'h40ba7658, 32'hc2653df2, 32'h423a82cf, 32'hc2b2de75, 32'h4085b07c, 32'hc2215b2f, 32'hc2487e27};
test_output[9082] = '{32'h42ba6637};
test_index[9082] = '{0};
test_input[72664:72671] = '{32'h4218b65d, 32'hc2a99709, 32'h4241eb7d, 32'h4229ee6a, 32'hc2a53c12, 32'h41f8ceed, 32'h4177de6d, 32'h41af0200};
test_output[9083] = '{32'h4241eb7d};
test_index[9083] = '{2};
test_input[72672:72679] = '{32'hc2931a93, 32'hc15f2357, 32'hc224d439, 32'hc1fa62aa, 32'h3fc84162, 32'h426873f4, 32'hc1675a44, 32'h42217134};
test_output[9084] = '{32'h426873f4};
test_index[9084] = '{5};
test_input[72680:72687] = '{32'h42b90c5f, 32'hc18173e8, 32'h40e106f4, 32'h424461fd, 32'h41b2aabf, 32'hc28bbc63, 32'hc2b7a1ee, 32'hc2ba0e5a};
test_output[9085] = '{32'h42b90c5f};
test_index[9085] = '{0};
test_input[72688:72695] = '{32'h414694e9, 32'hc236da84, 32'hc2989503, 32'hc1c56e9d, 32'h4114a58a, 32'h41d02273, 32'hc1def273, 32'hc2a027d9};
test_output[9086] = '{32'h41d02273};
test_index[9086] = '{5};
test_input[72696:72703] = '{32'hc189592f, 32'hc209599c, 32'h42274f47, 32'h42a98c2c, 32'h41aac745, 32'hc216a5b0, 32'h42236178, 32'h4248b081};
test_output[9087] = '{32'h42a98c2c};
test_index[9087] = '{3};
test_input[72704:72711] = '{32'h413a4154, 32'hc26296cd, 32'h42b9728a, 32'h3fb8ca68, 32'hc18aeee2, 32'h4102c934, 32'hc2a14863, 32'hc2149cf4};
test_output[9088] = '{32'h42b9728a};
test_index[9088] = '{2};
test_input[72712:72719] = '{32'h41cfb6a4, 32'hc163f773, 32'hc2254b5e, 32'h42c47128, 32'h421dd245, 32'hc1664bc2, 32'h424363a1, 32'h4164ddea};
test_output[9089] = '{32'h42c47128};
test_index[9089] = '{3};
test_input[72720:72727] = '{32'hc02b1505, 32'h428a1e08, 32'hbfd81e92, 32'h4182adca, 32'hc0990823, 32'hc2906aa4, 32'hc188e5a3, 32'hc21f2c11};
test_output[9090] = '{32'h428a1e08};
test_index[9090] = '{1};
test_input[72728:72735] = '{32'h42b5e2e6, 32'h3f8ea9ed, 32'hc0eb6c2a, 32'hc1d60ebb, 32'hc29bb7d0, 32'hc090cceb, 32'hc2897fa0, 32'h4290b5e5};
test_output[9091] = '{32'h42b5e2e6};
test_index[9091] = '{0};
test_input[72736:72743] = '{32'h42422a66, 32'hc2c56f23, 32'hc2a8c9ac, 32'h4237d3c2, 32'hc1947ac7, 32'hc0471608, 32'h42118845, 32'h423408d3};
test_output[9092] = '{32'h42422a66};
test_index[9092] = '{0};
test_input[72744:72751] = '{32'hc2826880, 32'h4243cf7d, 32'hc287a318, 32'hc15b0a10, 32'hc24c7397, 32'hc2b7d289, 32'h4244ab27, 32'h42335efa};
test_output[9093] = '{32'h4244ab27};
test_index[9093] = '{6};
test_input[72752:72759] = '{32'hc268035a, 32'h42b05e6e, 32'h41e05efa, 32'hc2a24433, 32'h42476454, 32'hc26af258, 32'hc217680f, 32'hc22795c6};
test_output[9094] = '{32'h42b05e6e};
test_index[9094] = '{1};
test_input[72760:72767] = '{32'h42765cc8, 32'h41b36444, 32'hc2a25552, 32'hc243a549, 32'hc1983144, 32'h422d6edc, 32'h421f6a06, 32'h4276e54a};
test_output[9095] = '{32'h4276e54a};
test_index[9095] = '{7};
test_input[72768:72775] = '{32'h42aa03d8, 32'h4138b5cd, 32'h4204ebe6, 32'h4285e46b, 32'hc2960b37, 32'h425ffd16, 32'h429a32f5, 32'h4291e96b};
test_output[9096] = '{32'h42aa03d8};
test_index[9096] = '{0};
test_input[72776:72783] = '{32'h42386626, 32'hc1354ab9, 32'h40fa31ea, 32'hc2a3f681, 32'h429005f2, 32'h413df07d, 32'hc1cb13ee, 32'hbf88d2a0};
test_output[9097] = '{32'h429005f2};
test_index[9097] = '{4};
test_input[72784:72791] = '{32'h40ba39b3, 32'h42059e96, 32'hc28a408e, 32'hc242cd64, 32'hc1c22da6, 32'hc1987a3a, 32'h414d8f1d, 32'h421e1b0e};
test_output[9098] = '{32'h421e1b0e};
test_index[9098] = '{7};
test_input[72792:72799] = '{32'hc1126e64, 32'h426d14d5, 32'h40ad214b, 32'hc1a325a8, 32'h42116ddb, 32'hbf250a2f, 32'h42c6d688, 32'h42676fb3};
test_output[9099] = '{32'h42c6d688};
test_index[9099] = '{6};
test_input[72800:72807] = '{32'h41fbd6e9, 32'h42b8a795, 32'h41d13703, 32'hc21f3a88, 32'hc18c9678, 32'h41492a98, 32'hc2ba4a50, 32'h41f2706f};
test_output[9100] = '{32'h42b8a795};
test_index[9100] = '{1};
test_input[72808:72815] = '{32'hc2a4f66d, 32'hc2853f79, 32'h40e4970a, 32'hc114271e, 32'h41bd3179, 32'hc0dfd2a3, 32'h428fbd28, 32'hc2170fee};
test_output[9101] = '{32'h428fbd28};
test_index[9101] = '{6};
test_input[72816:72823] = '{32'h42a2a974, 32'h424ed00d, 32'h42be05f6, 32'h41dbb1cc, 32'hc215f4ff, 32'hc2156689, 32'hc2693220, 32'hc19e6966};
test_output[9102] = '{32'h42be05f6};
test_index[9102] = '{2};
test_input[72824:72831] = '{32'hc0ddbadd, 32'hc2bc35ac, 32'h427eca0b, 32'hc2c63bf0, 32'hc2bd5f09, 32'h4212cd42, 32'h42254e79, 32'h424bf143};
test_output[9103] = '{32'h427eca0b};
test_index[9103] = '{2};
test_input[72832:72839] = '{32'h428d4919, 32'hc2c5567a, 32'hc2449b15, 32'h42c53e18, 32'hc1a53c89, 32'h424a509c, 32'hc1e39104, 32'hc16b44c4};
test_output[9104] = '{32'h42c53e18};
test_index[9104] = '{3};
test_input[72840:72847] = '{32'hc2c4a315, 32'h42b6cda9, 32'hc2a00141, 32'h41e57902, 32'h429a278a, 32'h4246c389, 32'hc2a8171e, 32'hc2c08724};
test_output[9105] = '{32'h42b6cda9};
test_index[9105] = '{1};
test_input[72848:72855] = '{32'hc22b8d20, 32'h41f39bfe, 32'hc2be67d0, 32'hc16a3432, 32'hc243b5e8, 32'hc053e2ed, 32'h42b0d7ac, 32'hc0be0394};
test_output[9106] = '{32'h42b0d7ac};
test_index[9106] = '{6};
test_input[72856:72863] = '{32'hc1ef24de, 32'hc236961c, 32'h4299acd2, 32'hc237c92e, 32'hc29f8453, 32'h41bffc1a, 32'h4090a4a5, 32'hc1dc513d};
test_output[9107] = '{32'h4299acd2};
test_index[9107] = '{2};
test_input[72864:72871] = '{32'hc0c91160, 32'h4235bb3c, 32'h42609d24, 32'hc0fcdd74, 32'hc2c326c3, 32'hc0aa2559, 32'hc2b89c1f, 32'h428b6329};
test_output[9108] = '{32'h428b6329};
test_index[9108] = '{7};
test_input[72872:72879] = '{32'h4257450b, 32'h4294f1e8, 32'hc2c77bd9, 32'hc154b635, 32'h427734fb, 32'h41a296a8, 32'h42bb241a, 32'h422668ee};
test_output[9109] = '{32'h42bb241a};
test_index[9109] = '{6};
test_input[72880:72887] = '{32'h42b379d6, 32'hc21896cd, 32'hc0e3695f, 32'hc0b72502, 32'hc26aa71d, 32'hc2abe24c, 32'hc2c03d48, 32'h42c66e5c};
test_output[9110] = '{32'h42c66e5c};
test_index[9110] = '{7};
test_input[72888:72895] = '{32'h412fdf93, 32'hc2a0a4ef, 32'hc1742900, 32'hc19224c6, 32'h41be0883, 32'hc2742b7d, 32'hc2bfa5c8, 32'h42106a06};
test_output[9111] = '{32'h42106a06};
test_index[9111] = '{7};
test_input[72896:72903] = '{32'hc28eb15c, 32'hc293aeba, 32'hc0d8674a, 32'h4280b647, 32'h42ae222a, 32'hc1abfed2, 32'hc2a5ca82, 32'h42a98bcf};
test_output[9112] = '{32'h42ae222a};
test_index[9112] = '{4};
test_input[72904:72911] = '{32'hc013a7e6, 32'hc1f2f90e, 32'hc272f453, 32'hc2c1f714, 32'h4267ec0a, 32'hc23f481d, 32'h42323166, 32'hc256f768};
test_output[9113] = '{32'h4267ec0a};
test_index[9113] = '{4};
test_input[72912:72919] = '{32'h4248620f, 32'hc23d4dda, 32'h42455066, 32'hc2c0e105, 32'hc1c72903, 32'h42a3a248, 32'hc0903bae, 32'h41ec34c8};
test_output[9114] = '{32'h42a3a248};
test_index[9114] = '{5};
test_input[72920:72927] = '{32'hc272e06e, 32'hc2b09b97, 32'h415e2538, 32'h42c7dbeb, 32'h42178494, 32'h41f775e7, 32'hc08b80ea, 32'hc2ac9064};
test_output[9115] = '{32'h42c7dbeb};
test_index[9115] = '{3};
test_input[72928:72935] = '{32'hc1dd8cf0, 32'hc24b88f4, 32'hc296ab7e, 32'h42c7ecc0, 32'hc2a2abdf, 32'h425cd357, 32'h4090c521, 32'h41451cda};
test_output[9116] = '{32'h42c7ecc0};
test_index[9116] = '{3};
test_input[72936:72943] = '{32'h42045306, 32'h428fbe09, 32'hc1f82ff6, 32'hc2851212, 32'hc2c4a716, 32'h4269f97c, 32'hc2c66afe, 32'hc2380bac};
test_output[9117] = '{32'h428fbe09};
test_index[9117] = '{1};
test_input[72944:72951] = '{32'h4193f885, 32'h4208c408, 32'hc0fb6a39, 32'h42b25d12, 32'hc284bdce, 32'hc22777ae, 32'h4230eb5e, 32'h42072f4d};
test_output[9118] = '{32'h42b25d12};
test_index[9118] = '{3};
test_input[72952:72959] = '{32'h42c2cba5, 32'h42996372, 32'h42137a99, 32'hc28168f2, 32'h4262906f, 32'h42063473, 32'hc0b6aef6, 32'hc28a674e};
test_output[9119] = '{32'h42c2cba5};
test_index[9119] = '{0};
test_input[72960:72967] = '{32'hc2387e9b, 32'hc28c9a04, 32'hc2a6d481, 32'hc21de2c4, 32'h42a2f0e4, 32'hc2665e16, 32'hc2356f75, 32'h42863080};
test_output[9120] = '{32'h42a2f0e4};
test_index[9120] = '{4};
test_input[72968:72975] = '{32'hc234d792, 32'h420a5570, 32'hc26a48b8, 32'hbe1fc50c, 32'hc1fde5b9, 32'hc13ce05a, 32'hc1c19b96, 32'hc25f4430};
test_output[9121] = '{32'h420a5570};
test_index[9121] = '{1};
test_input[72976:72983] = '{32'h41463838, 32'h42ab718c, 32'h42285cb8, 32'h424935f9, 32'h42294577, 32'hc2834082, 32'hc2c504e7, 32'h416d1bb6};
test_output[9122] = '{32'h42ab718c};
test_index[9122] = '{1};
test_input[72984:72991] = '{32'hc2bd63f6, 32'h429e4100, 32'hc29d0256, 32'h42952753, 32'h42c09c12, 32'hc248b0ec, 32'hc21bcbcd, 32'h428d3ae6};
test_output[9123] = '{32'h42c09c12};
test_index[9123] = '{4};
test_input[72992:72999] = '{32'h42abb5c8, 32'h42046d1b, 32'h403909fe, 32'hc215c07b, 32'hc241cd2a, 32'hbfd34915, 32'hc1fa18e4, 32'h4244ecb5};
test_output[9124] = '{32'h42abb5c8};
test_index[9124] = '{0};
test_input[73000:73007] = '{32'h42c13e0e, 32'h40c2a944, 32'hc280ba8c, 32'h42b45928, 32'h4190001a, 32'h420b8d3c, 32'hc0941b05, 32'h4168ad4f};
test_output[9125] = '{32'h42c13e0e};
test_index[9125] = '{0};
test_input[73008:73015] = '{32'hc23511ca, 32'h42b7e917, 32'hc2136173, 32'h417c3dd5, 32'h42ab4a82, 32'h42a7384a, 32'h4275f1d1, 32'h423b0646};
test_output[9126] = '{32'h42b7e917};
test_index[9126] = '{1};
test_input[73016:73023] = '{32'h42488f16, 32'hc0a435d8, 32'hc2c741d3, 32'hc289d4d3, 32'h42bf8438, 32'hc2bd7031, 32'hc282baf0, 32'h425e93d3};
test_output[9127] = '{32'h42bf8438};
test_index[9127] = '{4};
test_input[73024:73031] = '{32'hc2c5bbf4, 32'h4282c2a7, 32'h428ead86, 32'h41e06baa, 32'h41d561a3, 32'h41caead3, 32'h42010325, 32'hc0bf1456};
test_output[9128] = '{32'h428ead86};
test_index[9128] = '{2};
test_input[73032:73039] = '{32'hc26ee5ee, 32'h42af9b94, 32'hc220d9ad, 32'h41f32740, 32'h4262213f, 32'hc2554298, 32'hc28ca8ae, 32'hc1d85bee};
test_output[9129] = '{32'h42af9b94};
test_index[9129] = '{1};
test_input[73040:73047] = '{32'h41844c2e, 32'h41a1aa59, 32'h42b1802e, 32'hc2793033, 32'hc2b3d8d6, 32'h4211396a, 32'h42b8263f, 32'hc2aeda55};
test_output[9130] = '{32'h42b8263f};
test_index[9130] = '{6};
test_input[73048:73055] = '{32'hc2a881ee, 32'hc0cc4bbe, 32'h42a6b30e, 32'h4293aad6, 32'h42951408, 32'h429cbbb8, 32'hc2680c9c, 32'hc1f4ab15};
test_output[9131] = '{32'h42a6b30e};
test_index[9131] = '{2};
test_input[73056:73063] = '{32'h42951290, 32'hc1f4d808, 32'h42230a2a, 32'h42a1ef61, 32'hc24594c3, 32'hc246c64b, 32'h4217ad06, 32'h418a6505};
test_output[9132] = '{32'h42a1ef61};
test_index[9132] = '{3};
test_input[73064:73071] = '{32'hc2a1d29b, 32'hc29ddce0, 32'h420b2bb2, 32'hc23571e1, 32'h42b3a8f2, 32'h4163a763, 32'h41d9044f, 32'hc1689bcd};
test_output[9133] = '{32'h42b3a8f2};
test_index[9133] = '{4};
test_input[73072:73079] = '{32'h42329569, 32'h42209670, 32'h3f6ecbe9, 32'hc2325dd9, 32'hc29080b1, 32'hc1313809, 32'hbf8a94ac, 32'hc27092fa};
test_output[9134] = '{32'h42329569};
test_index[9134] = '{0};
test_input[73080:73087] = '{32'hc1f7f5f1, 32'hc281ebae, 32'h41dab7dc, 32'hc10b726a, 32'hc2737478, 32'h428b0a17, 32'h422045dd, 32'h429928e6};
test_output[9135] = '{32'h429928e6};
test_index[9135] = '{7};
test_input[73088:73095] = '{32'hc298fbe3, 32'h42346264, 32'hc244478b, 32'h41cb2816, 32'h429c9281, 32'hc195b978, 32'hc2846d43, 32'h4299613b};
test_output[9136] = '{32'h429c9281};
test_index[9136] = '{4};
test_input[73096:73103] = '{32'h42c3290d, 32'h42bdcbe2, 32'hc2c1ef64, 32'hc23182cb, 32'h42817429, 32'hc13b7976, 32'h424a620d, 32'h422af69c};
test_output[9137] = '{32'h42c3290d};
test_index[9137] = '{0};
test_input[73104:73111] = '{32'h42350d67, 32'hc1c0886a, 32'hc2647627, 32'h428e1fdf, 32'h41a35a9f, 32'h426ccbe8, 32'hc2c69955, 32'h3f63770b};
test_output[9138] = '{32'h428e1fdf};
test_index[9138] = '{3};
test_input[73112:73119] = '{32'h4185acfc, 32'h42ace4c7, 32'hc125654b, 32'hc12298ff, 32'hc20e4b78, 32'h42c3ee67, 32'h42469a0e, 32'hc247e511};
test_output[9139] = '{32'h42c3ee67};
test_index[9139] = '{5};
test_input[73120:73127] = '{32'h427d326f, 32'h4262f2d9, 32'hc1a8fa3e, 32'h4243ec15, 32'h419c3df1, 32'h4268860b, 32'hc296ee17, 32'h41d38fec};
test_output[9140] = '{32'h427d326f};
test_index[9140] = '{0};
test_input[73128:73135] = '{32'h429005a5, 32'h421ecade, 32'h421faebb, 32'h42123f01, 32'hc1aca97f, 32'h421e2771, 32'h42ba3581, 32'h421c1afc};
test_output[9141] = '{32'h42ba3581};
test_index[9141] = '{6};
test_input[73136:73143] = '{32'h41ef1bff, 32'hc1e7be9b, 32'hc20c397e, 32'hc20cf7d1, 32'hc1e36db5, 32'hc07080a2, 32'hc252d1ab, 32'hc222deb5};
test_output[9142] = '{32'h41ef1bff};
test_index[9142] = '{0};
test_input[73144:73151] = '{32'h42753636, 32'hc1c27834, 32'h42b3d327, 32'hc2457239, 32'h42021fc5, 32'hc2186d5c, 32'hc266c5a2, 32'h40c4261c};
test_output[9143] = '{32'h42b3d327};
test_index[9143] = '{2};
test_input[73152:73159] = '{32'h40b07c06, 32'hc2677d6f, 32'h42830a4b, 32'h41f2c7ea, 32'hc2811fea, 32'h41b1c029, 32'h4289a31f, 32'hc1b06ae7};
test_output[9144] = '{32'h4289a31f};
test_index[9144] = '{6};
test_input[73160:73167] = '{32'hc06474b1, 32'h41ac33ad, 32'hc206915d, 32'hc26b75c6, 32'h426cbd28, 32'h4279272b, 32'hc285ab59, 32'h41d3ded6};
test_output[9145] = '{32'h4279272b};
test_index[9145] = '{5};
test_input[73168:73175] = '{32'h42c6bf27, 32'hc262e47c, 32'hc1eac62f, 32'h424a624e, 32'h410663b7, 32'h42132022, 32'hc2ab8b3b, 32'h42a6367f};
test_output[9146] = '{32'h42c6bf27};
test_index[9146] = '{0};
test_input[73176:73183] = '{32'h41ef02b2, 32'h42ab10b2, 32'hc2bbe8b5, 32'h42ae3a77, 32'h42c03a82, 32'hc272c331, 32'hc2c02f1f, 32'hc29d335c};
test_output[9147] = '{32'h42c03a82};
test_index[9147] = '{4};
test_input[73184:73191] = '{32'h42b318d8, 32'hc2a5f4ce, 32'h41b81f84, 32'hc24c6c47, 32'hc10a4eaa, 32'h41fd937c, 32'hc24226db, 32'hc2ba89a0};
test_output[9148] = '{32'h42b318d8};
test_index[9148] = '{0};
test_input[73192:73199] = '{32'h42aaaadb, 32'h42622722, 32'hc220959e, 32'hc10dba13, 32'hc159efb9, 32'hc27ebae4, 32'hc29e6f28, 32'h428f572e};
test_output[9149] = '{32'h42aaaadb};
test_index[9149] = '{0};
test_input[73200:73207] = '{32'h41edff51, 32'h42120ac9, 32'hc1aedfeb, 32'h417cc978, 32'hc2a0cd2c, 32'h41d542ed, 32'hc28c54a8, 32'h4221e0e5};
test_output[9150] = '{32'h4221e0e5};
test_index[9150] = '{7};
test_input[73208:73215] = '{32'h4203ff04, 32'hc1b54175, 32'h4274c951, 32'hc05c2adf, 32'hc11faa21, 32'hc21df4b3, 32'h420d8414, 32'hc2881319};
test_output[9151] = '{32'h4274c951};
test_index[9151] = '{2};
test_input[73216:73223] = '{32'hc2908b32, 32'hc2a3ca51, 32'h42b697dc, 32'hc1ca62b8, 32'hc137c5d6, 32'hc25c0783, 32'hc2b259dc, 32'h4298c310};
test_output[9152] = '{32'h42b697dc};
test_index[9152] = '{2};
test_input[73224:73231] = '{32'h4284099d, 32'h42c5437f, 32'h42a3ffe7, 32'h4247ea3d, 32'hc2762704, 32'h429075ea, 32'hbfa23e50, 32'hc2898142};
test_output[9153] = '{32'h42c5437f};
test_index[9153] = '{1};
test_input[73232:73239] = '{32'hc26688da, 32'hc2968ea7, 32'h40516403, 32'h404cc927, 32'hc209976b, 32'h42ad32d5, 32'h420f2a21, 32'h41992f2e};
test_output[9154] = '{32'h42ad32d5};
test_index[9154] = '{5};
test_input[73240:73247] = '{32'hc2805b37, 32'h425e3b17, 32'h42a4dbbb, 32'h4295d43f, 32'hc25613ee, 32'hc29b8d7a, 32'hc08abd0a, 32'hc281a39a};
test_output[9155] = '{32'h42a4dbbb};
test_index[9155] = '{2};
test_input[73248:73255] = '{32'h41d57bfd, 32'h42bfbd53, 32'hc24e33fb, 32'hc20da88e, 32'hc280b321, 32'hc11702fa, 32'hc2b4698c, 32'h421f2fd8};
test_output[9156] = '{32'h42bfbd53};
test_index[9156] = '{1};
test_input[73256:73263] = '{32'h42b9ff5e, 32'hc28d9b9c, 32'hc1916919, 32'hc287c8dd, 32'h4155e132, 32'hc29e0f03, 32'hc2478b59, 32'h41e3b247};
test_output[9157] = '{32'h42b9ff5e};
test_index[9157] = '{0};
test_input[73264:73271] = '{32'hc293eebc, 32'h4225871c, 32'h42131be9, 32'hc204f2ac, 32'hc2ba1765, 32'hc2390cd4, 32'hc20e8127, 32'h412f9d1d};
test_output[9158] = '{32'h4225871c};
test_index[9158] = '{1};
test_input[73272:73279] = '{32'hc2c5952d, 32'hc2797bb6, 32'hc2a173ba, 32'hc1b66f68, 32'h419b6161, 32'h4292cbf4, 32'h42b90d6d, 32'hc203e052};
test_output[9159] = '{32'h42b90d6d};
test_index[9159] = '{6};
test_input[73280:73287] = '{32'hc269f96b, 32'hc2464814, 32'hc2bb7a6f, 32'hc128efe9, 32'h429615ba, 32'h4139a880, 32'h41d6bac1, 32'hc2a99299};
test_output[9160] = '{32'h429615ba};
test_index[9160] = '{4};
test_input[73288:73295] = '{32'hc25e01c5, 32'h40d297d8, 32'h42350633, 32'hc2c4eacc, 32'hc20b9c5a, 32'h41fe4972, 32'h4227e08a, 32'h41d3271e};
test_output[9161] = '{32'h42350633};
test_index[9161] = '{2};
test_input[73296:73303] = '{32'h41319e37, 32'hc28ef94e, 32'hc2a93c44, 32'h42a7d9cc, 32'hc2aa0920, 32'hc267e6cb, 32'h420dec15, 32'hc052b709};
test_output[9162] = '{32'h42a7d9cc};
test_index[9162] = '{3};
test_input[73304:73311] = '{32'hc15b217e, 32'hc2a39b43, 32'hc058994f, 32'h42a3a797, 32'h41987901, 32'h423a82f8, 32'hc2a15132, 32'hc1b0a6ab};
test_output[9163] = '{32'h42a3a797};
test_index[9163] = '{3};
test_input[73312:73319] = '{32'hc27a2583, 32'hc215fe0f, 32'h42c52135, 32'h42223428, 32'h418a2f8d, 32'h3ef543c7, 32'hc29868fb, 32'h41384d88};
test_output[9164] = '{32'h42c52135};
test_index[9164] = '{2};
test_input[73320:73327] = '{32'h41c363e1, 32'hc28ffc56, 32'hc29164dd, 32'hc2a96a6f, 32'hc2722c4d, 32'h41929eec, 32'hc248504c, 32'h409beae1};
test_output[9165] = '{32'h41c363e1};
test_index[9165] = '{0};
test_input[73328:73335] = '{32'hc0e1b123, 32'hc2a8f731, 32'h42bb3d9d, 32'hc28d8764, 32'hc2a7aa32, 32'h42c50721, 32'h4295e727, 32'h42b006a4};
test_output[9166] = '{32'h42c50721};
test_index[9166] = '{5};
test_input[73336:73343] = '{32'hc205e4b8, 32'h4163037c, 32'h42810151, 32'hc21ff8e3, 32'h425bf0e6, 32'hc17317c6, 32'h429bc781, 32'hc1c728b2};
test_output[9167] = '{32'h429bc781};
test_index[9167] = '{6};
test_input[73344:73351] = '{32'hbf955d87, 32'hc2609dbe, 32'hc28830ef, 32'h41a0320e, 32'hc21a445d, 32'hc20b43f5, 32'hc2863259, 32'hc27889bb};
test_output[9168] = '{32'h41a0320e};
test_index[9168] = '{3};
test_input[73352:73359] = '{32'hc2a10d08, 32'h4286fc96, 32'h41c676b7, 32'hc2a83000, 32'hc0047af4, 32'hc28766df, 32'hc2a73ed8, 32'hc22e54a3};
test_output[9169] = '{32'h4286fc96};
test_index[9169] = '{1};
test_input[73360:73367] = '{32'h4273d71e, 32'h412d4ec0, 32'h41d70ded, 32'h41e3dc75, 32'hc1eda05d, 32'h4215b318, 32'hc1849b0f, 32'hc12f908d};
test_output[9170] = '{32'h4273d71e};
test_index[9170] = '{0};
test_input[73368:73375] = '{32'h41313477, 32'h42a5fb8f, 32'hc2ba608e, 32'hc25dbb44, 32'hc2805a44, 32'hc215d11c, 32'hc2793058, 32'hc24e05b0};
test_output[9171] = '{32'h42a5fb8f};
test_index[9171] = '{1};
test_input[73376:73383] = '{32'h42b6625d, 32'h426ba1fb, 32'h41b58bc0, 32'h42bc8aae, 32'h42a608fe, 32'hc299e377, 32'hc1ec81be, 32'h414314e7};
test_output[9172] = '{32'h42bc8aae};
test_index[9172] = '{3};
test_input[73384:73391] = '{32'h413cb32a, 32'hc2ad5ff2, 32'hc2939af2, 32'h429f650c, 32'hc28bfaf2, 32'h423b105e, 32'hc0807fa0, 32'h4299ee40};
test_output[9173] = '{32'h429f650c};
test_index[9173] = '{3};
test_input[73392:73399] = '{32'hc0d6c4f2, 32'hc203ab47, 32'h4283d610, 32'hc21c0a5d, 32'h420ba9ea, 32'h3ffade6f, 32'h42b702ea, 32'h3fbedf70};
test_output[9174] = '{32'h42b702ea};
test_index[9174] = '{6};
test_input[73400:73407] = '{32'h42c1cc87, 32'h422f6a99, 32'h4201cf6a, 32'h4281fe63, 32'h429be484, 32'h422ed4a4, 32'hc2754d7b, 32'hc2a5b1a6};
test_output[9175] = '{32'h42c1cc87};
test_index[9175] = '{0};
test_input[73408:73415] = '{32'h42194348, 32'h412be67a, 32'hc08b1b75, 32'hc1aba369, 32'hc26f9876, 32'h42a8d9cc, 32'h42b9ef42, 32'h419c7d80};
test_output[9176] = '{32'h42b9ef42};
test_index[9176] = '{6};
test_input[73416:73423] = '{32'hc1418593, 32'h4158f623, 32'h4132c3d3, 32'h40277de6, 32'hc2c35c99, 32'hc298464d, 32'h42619dea, 32'h3e7e2ef5};
test_output[9177] = '{32'h42619dea};
test_index[9177] = '{6};
test_input[73424:73431] = '{32'hc2c32068, 32'hc21c7aa5, 32'hc27c747c, 32'hc2bba487, 32'h42b937ea, 32'hc2198b5a, 32'hc287949b, 32'hc21f6d98};
test_output[9178] = '{32'h42b937ea};
test_index[9178] = '{4};
test_input[73432:73439] = '{32'hc28a3cdb, 32'h41f78533, 32'hc251a568, 32'hc2a9854c, 32'h41a92819, 32'h42aadca0, 32'h42b3eae3, 32'hc1f17865};
test_output[9179] = '{32'h42b3eae3};
test_index[9179] = '{6};
test_input[73440:73447] = '{32'h42bdd6ae, 32'h42be685d, 32'hc2bc73d6, 32'hc1935640, 32'h41efeeae, 32'h42802f7e, 32'hc29aa560, 32'h42147f64};
test_output[9180] = '{32'h42be685d};
test_index[9180] = '{1};
test_input[73448:73455] = '{32'hc2ab1006, 32'h423f66b1, 32'hc2999281, 32'h41b2d133, 32'hc29ef749, 32'hc2a4bac7, 32'hc2359428, 32'hc19525c3};
test_output[9181] = '{32'h423f66b1};
test_index[9181] = '{1};
test_input[73456:73463] = '{32'h423d72f6, 32'h41457317, 32'hc2c471e2, 32'hc086f097, 32'h42b341cf, 32'hc17b7bd0, 32'h42660103, 32'hc28bb993};
test_output[9182] = '{32'h42b341cf};
test_index[9182] = '{4};
test_input[73464:73471] = '{32'h4280712f, 32'h418e37a8, 32'h41daf925, 32'hc2316f97, 32'h423e3535, 32'h40ee0937, 32'h41bab924, 32'h42287b1d};
test_output[9183] = '{32'h4280712f};
test_index[9183] = '{0};
test_input[73472:73479] = '{32'hc1d9d695, 32'h41872ee8, 32'h42acc905, 32'h42bf323a, 32'h428465f1, 32'h408fdf4b, 32'h41f07bb7, 32'hc2b3cc97};
test_output[9184] = '{32'h42bf323a};
test_index[9184] = '{3};
test_input[73480:73487] = '{32'h4211a0c1, 32'hc2a3392e, 32'h41c6be3d, 32'h4290add2, 32'hc0076f88, 32'h426d51ed, 32'hc1de1ea6, 32'hc2be01f3};
test_output[9185] = '{32'h4290add2};
test_index[9185] = '{3};
test_input[73488:73495] = '{32'h4194dc03, 32'h42c72201, 32'h41312d84, 32'h427d5541, 32'hc213dc4d, 32'hc1cceebe, 32'h422aa485, 32'hc2827497};
test_output[9186] = '{32'h42c72201};
test_index[9186] = '{1};
test_input[73496:73503] = '{32'hc241b908, 32'hc2b6a855, 32'hc25a884c, 32'hc26d771d, 32'hc2236c1d, 32'hc2a6b4af, 32'hc2b98565, 32'h42a77627};
test_output[9187] = '{32'h42a77627};
test_index[9187] = '{7};
test_input[73504:73511] = '{32'h42a463b8, 32'hc2793ba3, 32'h42219708, 32'hc27b1b4e, 32'hc12d066e, 32'hc166b3a9, 32'hc28504a6, 32'hbf49900f};
test_output[9188] = '{32'h42a463b8};
test_index[9188] = '{0};
test_input[73512:73519] = '{32'h429d111b, 32'h42139834, 32'h41d8868d, 32'hc1fab4ce, 32'hc2083c91, 32'h41ca37be, 32'h4102e440, 32'hc2bc3780};
test_output[9189] = '{32'h429d111b};
test_index[9189] = '{0};
test_input[73520:73527] = '{32'h423c9cf8, 32'hc26cf979, 32'h40e6f7eb, 32'h42a67ad0, 32'hc2c56d84, 32'h421e7b06, 32'h411a0c4d, 32'h42800ad2};
test_output[9190] = '{32'h42a67ad0};
test_index[9190] = '{3};
test_input[73528:73535] = '{32'hc1f7bf03, 32'h414e4777, 32'h4298484c, 32'hc0bb8829, 32'h42879008, 32'hc21a6086, 32'hc2baad26, 32'h42c7e5e3};
test_output[9191] = '{32'h42c7e5e3};
test_index[9191] = '{7};
test_input[73536:73543] = '{32'hc1bc7a76, 32'h42c33cfa, 32'hc097cef0, 32'h417b5903, 32'hc1546eb9, 32'hc2ab752f, 32'h419e01b8, 32'hc1b5b361};
test_output[9192] = '{32'h42c33cfa};
test_index[9192] = '{1};
test_input[73544:73551] = '{32'h41cf7c29, 32'hc285d101, 32'h42bfacb7, 32'hc25ec290, 32'h42127991, 32'h424825dd, 32'hc00d1180, 32'h42587734};
test_output[9193] = '{32'h42bfacb7};
test_index[9193] = '{2};
test_input[73552:73559] = '{32'h4248cc2e, 32'h41a47211, 32'hc2039daf, 32'h423e5d5b, 32'hc1c54174, 32'hc1ee2306, 32'h4194851d, 32'h424c5913};
test_output[9194] = '{32'h424c5913};
test_index[9194] = '{7};
test_input[73560:73567] = '{32'h4154e702, 32'h4267dc90, 32'hc1130da5, 32'hc21df8bd, 32'hc269114d, 32'hc2bf06f2, 32'h42c70860, 32'hc1a6e802};
test_output[9195] = '{32'h42c70860};
test_index[9195] = '{6};
test_input[73568:73575] = '{32'h4090fe76, 32'hc2b28e51, 32'h41ff0ca9, 32'h4252ac49, 32'hc273578d, 32'h41b48ac9, 32'hc2a3a7b6, 32'h41be442e};
test_output[9196] = '{32'h4252ac49};
test_index[9196] = '{3};
test_input[73576:73583] = '{32'h4252d203, 32'h41938140, 32'hc2b8925e, 32'hc2b7ec10, 32'h42a613f7, 32'hc119f5ec, 32'hc2bb315f, 32'h42266e9f};
test_output[9197] = '{32'h42a613f7};
test_index[9197] = '{4};
test_input[73584:73591] = '{32'hc292f4d1, 32'hc24570e7, 32'h41a21fb7, 32'hc29602b0, 32'hc19f6094, 32'hc281e66f, 32'hc1f2dc87, 32'h4299ec31};
test_output[9198] = '{32'h4299ec31};
test_index[9198] = '{7};
test_input[73592:73599] = '{32'h4214b54b, 32'hc1b4df2f, 32'h42a0f24c, 32'hbe215448, 32'hc1ee18c7, 32'hc260237b, 32'hc2a91a93, 32'hc2c56261};
test_output[9199] = '{32'h42a0f24c};
test_index[9199] = '{2};
test_input[73600:73607] = '{32'hc23f86fa, 32'h40bdd328, 32'h4205d3a2, 32'h42451f0f, 32'hc2a8540a, 32'hc240fcb3, 32'h3f9f19aa, 32'hc2a9633d};
test_output[9200] = '{32'h42451f0f};
test_index[9200] = '{3};
test_input[73608:73615] = '{32'h400b4660, 32'hc2bae5ad, 32'hc226124b, 32'h42b68db5, 32'h4228fe43, 32'hc1e9b53e, 32'h41a259d1, 32'hc2af87d0};
test_output[9201] = '{32'h42b68db5};
test_index[9201] = '{3};
test_input[73616:73623] = '{32'h427b2694, 32'hc086fe97, 32'h42b8a715, 32'h42127218, 32'h423af464, 32'h40a5eda6, 32'hc2b538a4, 32'h42325040};
test_output[9202] = '{32'h42b8a715};
test_index[9202] = '{2};
test_input[73624:73631] = '{32'h427cd3ec, 32'hc2689437, 32'h4269c299, 32'hc2bcbce5, 32'hc2524b2e, 32'h428a4491, 32'hc108a822, 32'hc289a1b3};
test_output[9203] = '{32'h428a4491};
test_index[9203] = '{5};
test_input[73632:73639] = '{32'hc2438569, 32'hc18c1ba2, 32'h42ad1f76, 32'hc2c32956, 32'h41e5ccd8, 32'hc27765db, 32'hc1de69ed, 32'hc2bc7ce4};
test_output[9204] = '{32'h42ad1f76};
test_index[9204] = '{2};
test_input[73640:73647] = '{32'h4243cd47, 32'hc1ca33b3, 32'hc20ba848, 32'h40f471e4, 32'hc1939ec4, 32'hc0e3c95f, 32'hc20a7932, 32'h4246d45f};
test_output[9205] = '{32'h4246d45f};
test_index[9205] = '{7};
test_input[73648:73655] = '{32'hc208bce2, 32'h42594937, 32'h42a158da, 32'hc2bdccb4, 32'h420ee549, 32'hc2beb68d, 32'hc1c971b6, 32'h42609365};
test_output[9206] = '{32'h42a158da};
test_index[9206] = '{2};
test_input[73656:73663] = '{32'h41297734, 32'h42abd0dc, 32'hc243d16d, 32'h428bcf65, 32'h41b1ee64, 32'hc1a4be72, 32'h416c4025, 32'h4168d12b};
test_output[9207] = '{32'h42abd0dc};
test_index[9207] = '{1};
test_input[73664:73671] = '{32'hc27200b3, 32'hc28e137e, 32'hc1870283, 32'hc1fff756, 32'hc16a05bd, 32'hc2a3b6a9, 32'hc1e716a6, 32'hc164aa33};
test_output[9208] = '{32'hc164aa33};
test_index[9208] = '{7};
test_input[73672:73679] = '{32'hc24919ba, 32'h42b7d163, 32'h411de749, 32'hc1185b40, 32'h425abd22, 32'h41f42b10, 32'h41c9a7aa, 32'hc25c2964};
test_output[9209] = '{32'h42b7d163};
test_index[9209] = '{1};
test_input[73680:73687] = '{32'h424f0764, 32'h40aecbd3, 32'hc286ceb0, 32'hc22a5f9e, 32'h4298818c, 32'h4197eae6, 32'h41c80a80, 32'h40bd68ee};
test_output[9210] = '{32'h4298818c};
test_index[9210] = '{4};
test_input[73688:73695] = '{32'h427a5a01, 32'h4294b2e2, 32'hc29418e4, 32'h424153db, 32'hc1adfbfb, 32'h42af2daa, 32'hc2b0a77b, 32'hc196ffd2};
test_output[9211] = '{32'h42af2daa};
test_index[9211] = '{5};
test_input[73696:73703] = '{32'h41187bfc, 32'hc25c943f, 32'h41f48c78, 32'hc1c65c5c, 32'hc2b0822c, 32'h423e082f, 32'h42b3e1cc, 32'h41c221d6};
test_output[9212] = '{32'h42b3e1cc};
test_index[9212] = '{6};
test_input[73704:73711] = '{32'hc2015aa2, 32'h42446ba8, 32'hc1e526da, 32'hc275e273, 32'hc09978b3, 32'hc1b44ee8, 32'hc2572044, 32'h422570cc};
test_output[9213] = '{32'h42446ba8};
test_index[9213] = '{1};
test_input[73712:73719] = '{32'hc22838f8, 32'h41828f12, 32'hc2b0458a, 32'hc29a9168, 32'h4283f4c4, 32'hc28ef3cd, 32'hc2c0bdc3, 32'hc2be3f15};
test_output[9214] = '{32'h4283f4c4};
test_index[9214] = '{4};
test_input[73720:73727] = '{32'hc214f4e1, 32'hc2a04c27, 32'hc240583a, 32'h421fd04e, 32'h3f10e018, 32'h424015e5, 32'h4241df3d, 32'h429b6076};
test_output[9215] = '{32'h429b6076};
test_index[9215] = '{7};
test_input[73728:73735] = '{32'hc18fbe18, 32'hc1a66723, 32'h42c20081, 32'h41c4c24d, 32'h41c9765b, 32'hc051d14c, 32'hc22278f8, 32'h42c0e756};
test_output[9216] = '{32'h42c20081};
test_index[9216] = '{2};
test_input[73736:73743] = '{32'hc18cd798, 32'hc2875248, 32'h42b7be0b, 32'hc114516f, 32'h42937648, 32'hc2768ddc, 32'hc26faec8, 32'h421741a1};
test_output[9217] = '{32'h42b7be0b};
test_index[9217] = '{2};
test_input[73744:73751] = '{32'hbfa9e8de, 32'h4270a349, 32'hc1940dff, 32'hc28085a2, 32'hc28889de, 32'h429eaca5, 32'h421ec9b4, 32'hc29d7089};
test_output[9218] = '{32'h429eaca5};
test_index[9218] = '{5};
test_input[73752:73759] = '{32'h4036dba0, 32'h411941db, 32'h42834880, 32'hc291b7b0, 32'h42bb83e0, 32'h427f8b67, 32'hc26ec2f7, 32'h41541455};
test_output[9219] = '{32'h42bb83e0};
test_index[9219] = '{4};
test_input[73760:73767] = '{32'hc1ee7091, 32'h40ba0ddc, 32'h410d6106, 32'hc2245e9d, 32'h4144f828, 32'hc21a1163, 32'hc2877606, 32'hc274f2b4};
test_output[9220] = '{32'h4144f828};
test_index[9220] = '{4};
test_input[73768:73775] = '{32'h40de8a76, 32'h41a89b72, 32'hc1d7b554, 32'hc1092123, 32'hc230e9ba, 32'hc208b627, 32'hc10111af, 32'hc2be904b};
test_output[9221] = '{32'h41a89b72};
test_index[9221] = '{1};
test_input[73776:73783] = '{32'h4225e109, 32'h425af671, 32'h4228a108, 32'hc0663aa9, 32'hc2010f68, 32'hc1e42f9c, 32'hc283ee65, 32'hc08af764};
test_output[9222] = '{32'h425af671};
test_index[9222] = '{1};
test_input[73784:73791] = '{32'h42b2b362, 32'hc280f133, 32'h42c7089c, 32'hc1f979af, 32'h42a43c0a, 32'h42b352b4, 32'hc2276c2a, 32'h41ea3dab};
test_output[9223] = '{32'h42c7089c};
test_index[9223] = '{2};
test_input[73792:73799] = '{32'hc2bc6945, 32'hc1579b8e, 32'h4272dc61, 32'h4265e442, 32'hc27755a8, 32'hc27f6020, 32'h42aa2663, 32'hc24636c8};
test_output[9224] = '{32'h42aa2663};
test_index[9224] = '{6};
test_input[73800:73807] = '{32'hc2ba9222, 32'hc2c12841, 32'h3f58c772, 32'h42919e47, 32'h4186c205, 32'h42837b15, 32'hc2041a41, 32'hc24d1575};
test_output[9225] = '{32'h42919e47};
test_index[9225] = '{3};
test_input[73808:73815] = '{32'h42464691, 32'hc2aa0b0a, 32'hc1ddd64d, 32'h421d7bb5, 32'h42c47137, 32'h422d31bc, 32'h41f708af, 32'hc21a78d9};
test_output[9226] = '{32'h42c47137};
test_index[9226] = '{4};
test_input[73816:73823] = '{32'hc296407d, 32'h423fdb42, 32'h420935b5, 32'h4292ec88, 32'h41911f60, 32'hc0a3d52d, 32'h3ff65277, 32'hc2412f50};
test_output[9227] = '{32'h4292ec88};
test_index[9227] = '{3};
test_input[73824:73831] = '{32'hc24fe091, 32'hc298ba68, 32'hc137b6d9, 32'h424e9db9, 32'hc05d63d4, 32'h413eff33, 32'h41db61d9, 32'h421d3f33};
test_output[9228] = '{32'h424e9db9};
test_index[9228] = '{3};
test_input[73832:73839] = '{32'h425b91d2, 32'h42bd7bc9, 32'hc2344ca3, 32'hc26f9f14, 32'hc23d308a, 32'hc1fe17f9, 32'h42aca5fc, 32'h42a43bef};
test_output[9229] = '{32'h42bd7bc9};
test_index[9229] = '{1};
test_input[73840:73847] = '{32'h41e076fa, 32'hc13447ad, 32'h42c7d17e, 32'h42a632fd, 32'h41f3802e, 32'hc13ce19a, 32'h4133c1c5, 32'h4131eba9};
test_output[9230] = '{32'h42c7d17e};
test_index[9230] = '{2};
test_input[73848:73855] = '{32'h42035a72, 32'hc188d05d, 32'hc1a6d69e, 32'h42bd1815, 32'hc184afa6, 32'hc26c9392, 32'hc225663b, 32'hc2a18402};
test_output[9231] = '{32'h42bd1815};
test_index[9231] = '{3};
test_input[73856:73863] = '{32'hbded4269, 32'h421c221d, 32'hc1fb5a8f, 32'h42b7e032, 32'hc08c7df0, 32'h42230f6b, 32'hc2ba4d15, 32'h4291ee3e};
test_output[9232] = '{32'h42b7e032};
test_index[9232] = '{3};
test_input[73864:73871] = '{32'hc2bb86d1, 32'hc1dd5b79, 32'hc187a45b, 32'h424145fd, 32'hc263e5cd, 32'hc192d327, 32'h42734abe, 32'h40bed396};
test_output[9233] = '{32'h42734abe};
test_index[9233] = '{6};
test_input[73872:73879] = '{32'hc263c06c, 32'h428b0fbb, 32'h42259ce9, 32'h413cab4d, 32'hc2b8f35e, 32'hc23bb86b, 32'hc24c9782, 32'hc1e54ea8};
test_output[9234] = '{32'h428b0fbb};
test_index[9234] = '{1};
test_input[73880:73887] = '{32'h42919d16, 32'h42a123b5, 32'h420fa462, 32'hc1a450de, 32'hc1fd9788, 32'h4111741d, 32'h4284f695, 32'h429c0a54};
test_output[9235] = '{32'h42a123b5};
test_index[9235] = '{1};
test_input[73888:73895] = '{32'hc2a513c1, 32'hc297e1f9, 32'h421c05d7, 32'h412d56e6, 32'h42846155, 32'hc290c6a2, 32'h41d3f91b, 32'hc1f519cc};
test_output[9236] = '{32'h42846155};
test_index[9236] = '{4};
test_input[73896:73903] = '{32'hc2b74b34, 32'hc2c3985a, 32'h41c5ae55, 32'h4280d141, 32'h4210d9bb, 32'h42867314, 32'h42abdae7, 32'h423bd4d1};
test_output[9237] = '{32'h42abdae7};
test_index[9237] = '{6};
test_input[73904:73911] = '{32'h4297b07a, 32'h41434534, 32'hc285432d, 32'hc2814d70, 32'hc2354c58, 32'hc23c6ffc, 32'h4286d7d5, 32'hc1fac412};
test_output[9238] = '{32'h4297b07a};
test_index[9238] = '{0};
test_input[73912:73919] = '{32'hc29aabc8, 32'hc2bb10da, 32'h420d83a7, 32'hc28c7270, 32'h41d3cd3f, 32'h414ec3d5, 32'hc297b1ff, 32'hc1675657};
test_output[9239] = '{32'h420d83a7};
test_index[9239] = '{2};
test_input[73920:73927] = '{32'hc2904182, 32'hc269caf1, 32'hc2b800bb, 32'hbefe1e22, 32'h41fe9984, 32'h42ad2286, 32'h416549a0, 32'hc286c50a};
test_output[9240] = '{32'h42ad2286};
test_index[9240] = '{5};
test_input[73928:73935] = '{32'h40474a37, 32'hc18c077e, 32'hc217ae31, 32'h429485da, 32'hc27e8c5b, 32'h42487e3f, 32'h42ae57ab, 32'hc2840593};
test_output[9241] = '{32'h42ae57ab};
test_index[9241] = '{6};
test_input[73936:73943] = '{32'hc20765f9, 32'h40bfcf48, 32'hc2132347, 32'hc1b7eb77, 32'h426e31b4, 32'h429f28b4, 32'h42c2da10, 32'h40c1084b};
test_output[9242] = '{32'h42c2da10};
test_index[9242] = '{6};
test_input[73944:73951] = '{32'h41ad8c48, 32'h42a3e8f1, 32'h42836fc3, 32'h418841d6, 32'hc28e42e1, 32'hc20ecea9, 32'h41dfd2bb, 32'hc14cf59f};
test_output[9243] = '{32'h42a3e8f1};
test_index[9243] = '{1};
test_input[73952:73959] = '{32'h427979c0, 32'hc23961f0, 32'hc27ba249, 32'h417f9e41, 32'hc2a90016, 32'h3f41d7ff, 32'hc0b1c5c8, 32'hc17f95e6};
test_output[9244] = '{32'h427979c0};
test_index[9244] = '{0};
test_input[73960:73967] = '{32'h41f1e0b4, 32'h408ea65f, 32'hc251681f, 32'h42ab0eae, 32'h423fba0e, 32'hc29c0f67, 32'h429f164f, 32'hc2bef74c};
test_output[9245] = '{32'h42ab0eae};
test_index[9245] = '{3};
test_input[73968:73975] = '{32'hc2a462c1, 32'hc2abbdca, 32'h42a66682, 32'hc2b68e3a, 32'h42991e85, 32'hc28a450b, 32'h423a0586, 32'h41f283c5};
test_output[9246] = '{32'h42a66682};
test_index[9246] = '{2};
test_input[73976:73983] = '{32'hc2b6d18e, 32'hc1ccdb0e, 32'hc10e168e, 32'hc22f27ea, 32'hc21f8e4a, 32'hc26cee38, 32'hc1988647, 32'hc1491597};
test_output[9247] = '{32'hc10e168e};
test_index[9247] = '{2};
test_input[73984:73991] = '{32'h411b8353, 32'hc0a2e78d, 32'hc2a56d07, 32'h424e0b22, 32'h42b0c8a0, 32'hc2aa3cd7, 32'h426b072e, 32'h41452de8};
test_output[9248] = '{32'h42b0c8a0};
test_index[9248] = '{4};
test_input[73992:73999] = '{32'h42bddd25, 32'h4293ed54, 32'h4238960a, 32'hc1cb4232, 32'hc24d1f80, 32'h426614a4, 32'h42a214aa, 32'hbfa1732a};
test_output[9249] = '{32'h42bddd25};
test_index[9249] = '{0};
test_input[74000:74007] = '{32'h42b5ebb5, 32'hc206b0d6, 32'h421af2c6, 32'h41fc0458, 32'h424095d4, 32'hc2964daa, 32'h410baa85, 32'hc21f48fc};
test_output[9250] = '{32'h42b5ebb5};
test_index[9250] = '{0};
test_input[74008:74015] = '{32'hc236c32b, 32'h400d6e2f, 32'h4186028c, 32'hbf509720, 32'h4258c4a1, 32'h429db48d, 32'h42695336, 32'h425a9139};
test_output[9251] = '{32'h429db48d};
test_index[9251] = '{5};
test_input[74016:74023] = '{32'hbf06e942, 32'h41e95fe6, 32'hc0fafd08, 32'hc1d9270a, 32'h425bd08d, 32'h42208aa9, 32'hc1bcb457, 32'h42a4330b};
test_output[9252] = '{32'h42a4330b};
test_index[9252] = '{7};
test_input[74024:74031] = '{32'hc298a0b6, 32'hc19d6c79, 32'hc226ca4d, 32'hc26a2bba, 32'hc211dc89, 32'hc280328d, 32'hc2269131, 32'h41f5c36b};
test_output[9253] = '{32'h41f5c36b};
test_index[9253] = '{7};
test_input[74032:74039] = '{32'hc24feb3e, 32'h42bb61e8, 32'h412f009a, 32'hc2c7a8b4, 32'h42b6bdfe, 32'h4256743a, 32'h41947ef5, 32'hc288b4da};
test_output[9254] = '{32'h42bb61e8};
test_index[9254] = '{1};
test_input[74040:74047] = '{32'hc26a2fcb, 32'h4056863a, 32'h4206c0d2, 32'hc1d8c213, 32'h427ac7f0, 32'hc2aeb4b7, 32'h42898ce5, 32'hc26370fb};
test_output[9255] = '{32'h42898ce5};
test_index[9255] = '{6};
test_input[74048:74055] = '{32'h41ec1e56, 32'hbfd81b4a, 32'h4290a5da, 32'hc19c4b65, 32'h42a244c4, 32'hc258c4c5, 32'h42285755, 32'hc29c5a4e};
test_output[9256] = '{32'h42a244c4};
test_index[9256] = '{4};
test_input[74056:74063] = '{32'hc22e41b3, 32'hc2b7ab46, 32'hc0f71933, 32'hc252a5e4, 32'h42b16439, 32'hc23df5ac, 32'h42129dc8, 32'hc2b742d6};
test_output[9257] = '{32'h42b16439};
test_index[9257] = '{4};
test_input[74064:74071] = '{32'hc265423f, 32'hc0ffcc23, 32'hc11b1ba2, 32'hc196d24d, 32'hc2934d88, 32'h410d10bc, 32'hc111df5d, 32'hc2a4aea1};
test_output[9258] = '{32'h410d10bc};
test_index[9258] = '{5};
test_input[74072:74079] = '{32'hc150dbc9, 32'hc23c690d, 32'h42846cec, 32'hc2564b50, 32'hc20db652, 32'h425b488a, 32'hc1ca6e0c, 32'h4296fd78};
test_output[9259] = '{32'h4296fd78};
test_index[9259] = '{7};
test_input[74080:74087] = '{32'hc1af8fa6, 32'h42377f59, 32'h4229eca2, 32'hc29afc8a, 32'hc2c59f11, 32'hc1805d68, 32'hc28ff8fc, 32'h41b64b93};
test_output[9260] = '{32'h42377f59};
test_index[9260] = '{1};
test_input[74088:74095] = '{32'hc2293cef, 32'hc1aad837, 32'hc26cc18e, 32'h4150651c, 32'h42c7c06e, 32'h420d7a7b, 32'h42c6a26c, 32'hc1dc2d0d};
test_output[9261] = '{32'h42c7c06e};
test_index[9261] = '{4};
test_input[74096:74103] = '{32'hc04cb924, 32'hc25965c0, 32'hc155dfd3, 32'hc2a8a302, 32'h42837fce, 32'hc16c50eb, 32'hc209d7d7, 32'hc0ca29d7};
test_output[9262] = '{32'h42837fce};
test_index[9262] = '{4};
test_input[74104:74111] = '{32'hc27ff903, 32'h42462b7d, 32'h42b6bad6, 32'hc166e77e, 32'h42c0ef25, 32'hc2a3a770, 32'hc23ffaa2, 32'hc2ad65b5};
test_output[9263] = '{32'h42c0ef25};
test_index[9263] = '{4};
test_input[74112:74119] = '{32'hc202bc5c, 32'hc28badfe, 32'h428b22bf, 32'h42a1afa9, 32'h429a1050, 32'hc1860547, 32'h42793d27, 32'hc1c69532};
test_output[9264] = '{32'h42a1afa9};
test_index[9264] = '{3};
test_input[74120:74127] = '{32'hc1c14c94, 32'hc2c7aecd, 32'hc2760679, 32'hc29f10bd, 32'hc279add9, 32'hc1855ed0, 32'h41723452, 32'hc2bb8669};
test_output[9265] = '{32'h41723452};
test_index[9265] = '{6};
test_input[74128:74135] = '{32'h42738cd2, 32'hc276ed0e, 32'h419d15d6, 32'hc2a6298d, 32'h42b68d7b, 32'h4146f5bc, 32'h42911ee1, 32'hc1869f11};
test_output[9266] = '{32'h42b68d7b};
test_index[9266] = '{4};
test_input[74136:74143] = '{32'h42966b46, 32'hc2c28ba3, 32'h41f3eaf1, 32'hc2ba19e8, 32'hc2702154, 32'h42a8992e, 32'hc2b69502, 32'h41f0933d};
test_output[9267] = '{32'h42a8992e};
test_index[9267] = '{5};
test_input[74144:74151] = '{32'h42c55c43, 32'hc2bbb40e, 32'hc205af86, 32'h42af6823, 32'h42b954c1, 32'hc273a450, 32'h42aa4df6, 32'hc074c254};
test_output[9268] = '{32'h42c55c43};
test_index[9268] = '{0};
test_input[74152:74159] = '{32'hc2323484, 32'hc1eaba92, 32'hc2611dd7, 32'hc223e573, 32'h4232bf90, 32'h421cd3fa, 32'h417bb7a3, 32'h42a3a9eb};
test_output[9269] = '{32'h42a3a9eb};
test_index[9269] = '{7};
test_input[74160:74167] = '{32'h426c11d5, 32'h4184bbbf, 32'hc205fc4e, 32'hc2afee50, 32'h428c8c03, 32'h41b817c8, 32'h41bf08b0, 32'hc274f69c};
test_output[9270] = '{32'h428c8c03};
test_index[9270] = '{4};
test_input[74168:74175] = '{32'h419e57e7, 32'h420fc30a, 32'hc2678e27, 32'hc1c6fa15, 32'hc29810ef, 32'hc25dfe52, 32'hc253770e, 32'h40980840};
test_output[9271] = '{32'h420fc30a};
test_index[9271] = '{1};
test_input[74176:74183] = '{32'hc283179e, 32'h426b1d45, 32'hc2c2c168, 32'hc2a17090, 32'hc282df17, 32'hc24e577b, 32'h42903302, 32'hc2b65ee3};
test_output[9272] = '{32'h42903302};
test_index[9272] = '{6};
test_input[74184:74191] = '{32'h420ef858, 32'hc1b85f6d, 32'h42964c4e, 32'h41c54d70, 32'hc209a3ae, 32'h420eb2de, 32'h41324b82, 32'h4151787a};
test_output[9273] = '{32'h42964c4e};
test_index[9273] = '{2};
test_input[74192:74199] = '{32'h429f0f1f, 32'h42815346, 32'h4290ea90, 32'hc2704f7e, 32'hc20d33ec, 32'hc28b9f46, 32'h42b7e92b, 32'hc156d863};
test_output[9274] = '{32'h42b7e92b};
test_index[9274] = '{6};
test_input[74200:74207] = '{32'hc157a4fb, 32'h42ad5062, 32'hc2281a53, 32'hc192a3f3, 32'hc231190d, 32'hc03ccb9c, 32'hc2b25ca1, 32'hc2825f46};
test_output[9275] = '{32'h42ad5062};
test_index[9275] = '{1};
test_input[74208:74215] = '{32'h421ff1e7, 32'h417b3285, 32'h4287eb95, 32'hc0f1eb43, 32'hc29e1c20, 32'h410c82e0, 32'h429f90ba, 32'hc2a6a2cb};
test_output[9276] = '{32'h429f90ba};
test_index[9276] = '{6};
test_input[74216:74223] = '{32'hc2c5807b, 32'h417e3bce, 32'hc2879a0f, 32'hc1f2a04d, 32'h424bb469, 32'hc2b73426, 32'hc21d813a, 32'hc2753164};
test_output[9277] = '{32'h424bb469};
test_index[9277] = '{4};
test_input[74224:74231] = '{32'hc0e58d7e, 32'hc2afa9f7, 32'hc21dec67, 32'hc2ba568a, 32'h41f55248, 32'hc23993ef, 32'hc22675b7, 32'hc20980e5};
test_output[9278] = '{32'h41f55248};
test_index[9278] = '{4};
test_input[74232:74239] = '{32'hc1ebcc24, 32'h3ec55b98, 32'hc03bf3e6, 32'h41f54542, 32'h42b7c237, 32'h428dd61f, 32'h409cc15e, 32'hc28fcd46};
test_output[9279] = '{32'h42b7c237};
test_index[9279] = '{4};
test_input[74240:74247] = '{32'hc2b657bd, 32'h42144b26, 32'h429c24e8, 32'h42a4a858, 32'h428beeca, 32'h42b2175f, 32'hc1cf1088, 32'hc2be1f85};
test_output[9280] = '{32'h42b2175f};
test_index[9280] = '{5};
test_input[74248:74255] = '{32'h42bf2119, 32'h42112376, 32'h4283dbd6, 32'hc2937a25, 32'hc2c0b3fd, 32'h42032cee, 32'h426b01f3, 32'hc27639af};
test_output[9281] = '{32'h42bf2119};
test_index[9281] = '{0};
test_input[74256:74263] = '{32'hc28bea28, 32'h42c3f32f, 32'h42ada5f2, 32'hc24f9f18, 32'h411ce4e6, 32'hc2343552, 32'hc281fe10, 32'h41a55df3};
test_output[9282] = '{32'h42c3f32f};
test_index[9282] = '{1};
test_input[74264:74271] = '{32'h409c7d90, 32'hc271c5b6, 32'hc27be36a, 32'hbff764f6, 32'hc2b34587, 32'hc24d2390, 32'hc2368737, 32'hc2a9d27e};
test_output[9283] = '{32'h409c7d90};
test_index[9283] = '{0};
test_input[74272:74279] = '{32'hc28be05e, 32'h42a0c1f5, 32'hc20119d2, 32'h41cc8101, 32'hc2888888, 32'hc273a85b, 32'h41b0eca2, 32'hc21170c8};
test_output[9284] = '{32'h42a0c1f5};
test_index[9284] = '{1};
test_input[74280:74287] = '{32'hc2b3bd30, 32'hc2ae75ad, 32'hc29186cd, 32'hc265ae75, 32'hc1a4e167, 32'h42b8eca6, 32'hc28a0f0b, 32'hc2822ea2};
test_output[9285] = '{32'h42b8eca6};
test_index[9285] = '{5};
test_input[74288:74295] = '{32'hc21935d6, 32'hc2510543, 32'h42a46e89, 32'h42a1a7ee, 32'hc1bfe746, 32'h428f3425, 32'h41647e00, 32'h4094305b};
test_output[9286] = '{32'h42a46e89};
test_index[9286] = '{2};
test_input[74296:74303] = '{32'hc2bd0956, 32'h42055a70, 32'hc1ccb310, 32'h42c0769c, 32'hc24b39cf, 32'h4146a4a8, 32'hc2aa6d2b, 32'h429c23cb};
test_output[9287] = '{32'h42c0769c};
test_index[9287] = '{3};
test_input[74304:74311] = '{32'hc2b268cd, 32'hc114db24, 32'hc2b0c439, 32'h42ba0e82, 32'hc2a75a8c, 32'h42b56f04, 32'hc158eba5, 32'h4270df2b};
test_output[9288] = '{32'h42ba0e82};
test_index[9288] = '{3};
test_input[74312:74319] = '{32'h413ce735, 32'h42979f67, 32'h42af4875, 32'h428529fe, 32'h4292bfaa, 32'hc279c605, 32'h426e7855, 32'hc2a9e8de};
test_output[9289] = '{32'h42af4875};
test_index[9289] = '{2};
test_input[74320:74327] = '{32'h41a489a2, 32'h421d79c9, 32'h42866631, 32'h426ff45a, 32'h42651f62, 32'hc1aee314, 32'h42694aff, 32'hc2c5397a};
test_output[9290] = '{32'h42866631};
test_index[9290] = '{2};
test_input[74328:74335] = '{32'h42c6a6a1, 32'h420761be, 32'hc23b90f2, 32'hc0f54c7e, 32'h41362414, 32'hc289d044, 32'h4225be0e, 32'h42a0a2ca};
test_output[9291] = '{32'h42c6a6a1};
test_index[9291] = '{0};
test_input[74336:74343] = '{32'hbd349016, 32'h42b01f3d, 32'h42c2db4f, 32'h42895302, 32'hc1bcf9e6, 32'h42937763, 32'hc2b8ab57, 32'hc2be79e5};
test_output[9292] = '{32'h42c2db4f};
test_index[9292] = '{2};
test_input[74344:74351] = '{32'hc1b72923, 32'hc27c3b7d, 32'h42242225, 32'hc2931fd3, 32'h421121ba, 32'h40aadc36, 32'hc25989b6, 32'h417c0fc1};
test_output[9293] = '{32'h42242225};
test_index[9293] = '{2};
test_input[74352:74359] = '{32'hc1c4d293, 32'hc28c3e5d, 32'h426b8ceb, 32'hc2163049, 32'h4287309d, 32'h41c8a88f, 32'h42a8ce90, 32'h4288ee38};
test_output[9294] = '{32'h42a8ce90};
test_index[9294] = '{6};
test_input[74360:74367] = '{32'hc21c097a, 32'h418ef802, 32'hc19ecf01, 32'h41e04f13, 32'h42bf0291, 32'h4278e16d, 32'hc1e76ebf, 32'hc1b7b6be};
test_output[9295] = '{32'h42bf0291};
test_index[9295] = '{4};
test_input[74368:74375] = '{32'h42343483, 32'hc2a91781, 32'hc0ec11f4, 32'hc20a9834, 32'h42209c70, 32'h424ba7d7, 32'h427fe386, 32'h418df3e7};
test_output[9296] = '{32'h427fe386};
test_index[9296] = '{6};
test_input[74376:74383] = '{32'hc2b98e0f, 32'h429e0872, 32'h41a8ed96, 32'h42837357, 32'hc23013b5, 32'hc29a9232, 32'h42924b13, 32'h41c90485};
test_output[9297] = '{32'h429e0872};
test_index[9297] = '{1};
test_input[74384:74391] = '{32'h4240e3bd, 32'hc19f4e2c, 32'hc220a871, 32'hc21a1e71, 32'h416cf31c, 32'hc2c5fa9d, 32'h40e650d0, 32'hc2834f4d};
test_output[9298] = '{32'h4240e3bd};
test_index[9298] = '{0};
test_input[74392:74399] = '{32'hc1c49001, 32'hc2bda3af, 32'h4235a369, 32'h42c01801, 32'hc1d6d0ba, 32'h42607c67, 32'hc06ff273, 32'h41221dd5};
test_output[9299] = '{32'h42c01801};
test_index[9299] = '{3};
test_input[74400:74407] = '{32'h42152e54, 32'h4284ba00, 32'h401eb436, 32'hc2b10a21, 32'hc28bd2d6, 32'h425bb2b5, 32'h426581b2, 32'hc1f296cb};
test_output[9300] = '{32'h4284ba00};
test_index[9300] = '{1};
test_input[74408:74415] = '{32'h408e6335, 32'hc2a9e85c, 32'hc28fc46a, 32'h428cb9d8, 32'hc2214370, 32'hc0e7fb45, 32'hc292e22c, 32'hc2be0c6a};
test_output[9301] = '{32'h428cb9d8};
test_index[9301] = '{3};
test_input[74416:74423] = '{32'h425165f8, 32'hc27e96b9, 32'hc27d4280, 32'h42163cb1, 32'h408b5b0e, 32'hc2b72fbd, 32'hc297a9ad, 32'h422fdbc6};
test_output[9302] = '{32'h425165f8};
test_index[9302] = '{0};
test_input[74424:74431] = '{32'h42bd3d2b, 32'hc20aaef6, 32'hc24d746e, 32'hc2b3e97c, 32'hc000d7d2, 32'h4188cdd1, 32'hc08ced45, 32'hc2aa9cd3};
test_output[9303] = '{32'h42bd3d2b};
test_index[9303] = '{0};
test_input[74432:74439] = '{32'hc2a7bb5f, 32'h4245879c, 32'h42b8d94e, 32'hc19d174b, 32'hc240e7e0, 32'h3fe7113d, 32'h409159c3, 32'h4105383f};
test_output[9304] = '{32'h42b8d94e};
test_index[9304] = '{2};
test_input[74440:74447] = '{32'h42237edc, 32'h404f3611, 32'hc2694da1, 32'h40861233, 32'hc1e799fc, 32'h4292cd6e, 32'h42a51414, 32'hc194621c};
test_output[9305] = '{32'h42a51414};
test_index[9305] = '{6};
test_input[74448:74455] = '{32'hc26cea43, 32'hc2b280b8, 32'hc2bca058, 32'hc2101c32, 32'hc2253f07, 32'h410a3ade, 32'h414df5a0, 32'h42a0fbc9};
test_output[9306] = '{32'h42a0fbc9};
test_index[9306] = '{7};
test_input[74456:74463] = '{32'hc281b56a, 32'h41ecc34a, 32'hc14e6a09, 32'hc0add8c0, 32'hc2a3e214, 32'hc1ddc7cf, 32'hc2967bf0, 32'hc276d06d};
test_output[9307] = '{32'h41ecc34a};
test_index[9307] = '{1};
test_input[74464:74471] = '{32'h40c5e119, 32'hc23162bc, 32'h40ca5008, 32'hc2802cb6, 32'hc28f3cd5, 32'hc2aad585, 32'h423942df, 32'hc16f1ffd};
test_output[9308] = '{32'h423942df};
test_index[9308] = '{6};
test_input[74472:74479] = '{32'h42548c43, 32'hc136dd9e, 32'hc23d572b, 32'hc242f4e4, 32'h4285c1d3, 32'hc26e2c70, 32'h41fbaa83, 32'hc2565e1e};
test_output[9309] = '{32'h4285c1d3};
test_index[9309] = '{4};
test_input[74480:74487] = '{32'hc1b3b165, 32'hc252a361, 32'hc04f3ee8, 32'hc10c690f, 32'h41efe9f4, 32'h40dae23e, 32'h4296b737, 32'hc2259ad2};
test_output[9310] = '{32'h4296b737};
test_index[9310] = '{6};
test_input[74488:74495] = '{32'hc18bb72f, 32'h412857fc, 32'h428a4a62, 32'hc1f77602, 32'h422f0a9f, 32'hc20dd442, 32'h4217eae4, 32'hc273525c};
test_output[9311] = '{32'h428a4a62};
test_index[9311] = '{2};
test_input[74496:74503] = '{32'hbfe155f3, 32'hc2ad2a0f, 32'hc29069a1, 32'h41857991, 32'h4220afa4, 32'hc12cd0b8, 32'h422bd4a9, 32'h4216d170};
test_output[9312] = '{32'h422bd4a9};
test_index[9312] = '{6};
test_input[74504:74511] = '{32'h42ac2a1e, 32'hc1a33a39, 32'hc10a642b, 32'hc243e7ab, 32'h41995208, 32'h42c48f5b, 32'h42b2a787, 32'h42347c7c};
test_output[9313] = '{32'h42c48f5b};
test_index[9313] = '{5};
test_input[74512:74519] = '{32'hc2a5df7b, 32'h42a67883, 32'hc209ef82, 32'hc243b0cc, 32'hc299d4ee, 32'h42846759, 32'hc1a03356, 32'hc15aecfd};
test_output[9314] = '{32'h42a67883};
test_index[9314] = '{1};
test_input[74520:74527] = '{32'hc294d7f7, 32'hc1fce6be, 32'hc19cc8bf, 32'hc1119a4b, 32'hc2c6ae40, 32'hc1fe2e71, 32'hc0bbab2a, 32'hc1af15dc};
test_output[9315] = '{32'hc0bbab2a};
test_index[9315] = '{6};
test_input[74528:74535] = '{32'h427a3e5f, 32'hc1687e15, 32'hc07974a5, 32'hc25958b2, 32'hc1bc7bc3, 32'h4283b290, 32'hc25af42a, 32'hc25c7666};
test_output[9316] = '{32'h4283b290};
test_index[9316] = '{5};
test_input[74536:74543] = '{32'hc1d2d903, 32'hc23c2a26, 32'h42618c78, 32'hc1d089e6, 32'hc28c89fb, 32'h4276df49, 32'hc2b767a7, 32'hc0bf51bd};
test_output[9317] = '{32'h4276df49};
test_index[9317] = '{5};
test_input[74544:74551] = '{32'h420e7905, 32'h42515209, 32'hc228a5d5, 32'hc195f7da, 32'hc2868d25, 32'hc279e4cb, 32'h42b96f49, 32'h42082db5};
test_output[9318] = '{32'h42b96f49};
test_index[9318] = '{6};
test_input[74552:74559] = '{32'hc297f3b9, 32'hc2bb93b8, 32'hc1c83828, 32'hc2c541fe, 32'hc257a863, 32'h41c3f4dc, 32'hbecef092, 32'h42a846c6};
test_output[9319] = '{32'h42a846c6};
test_index[9319] = '{7};
test_input[74560:74567] = '{32'hc2831588, 32'h4224798c, 32'h42bf0c12, 32'hc2a97ac9, 32'h42857788, 32'h42428eef, 32'h4259ae00, 32'h4289a8a1};
test_output[9320] = '{32'h42bf0c12};
test_index[9320] = '{2};
test_input[74568:74575] = '{32'h4206fe4b, 32'hc2b43866, 32'h42686c5c, 32'hc29cda29, 32'hc298a5b8, 32'h42348464, 32'h42b76f1e, 32'h42c765f7};
test_output[9321] = '{32'h42c765f7};
test_index[9321] = '{7};
test_input[74576:74583] = '{32'h42266038, 32'h425d3418, 32'hbe1453a7, 32'h41bb3fa5, 32'h4228a8b9, 32'hc1e6a7cb, 32'hc1a77c92, 32'h4205aa20};
test_output[9322] = '{32'h425d3418};
test_index[9322] = '{1};
test_input[74584:74591] = '{32'h420eaba4, 32'hbe98200a, 32'h42328f91, 32'h42303b2d, 32'h41991eec, 32'h429ddf18, 32'h429db096, 32'h41b802e7};
test_output[9323] = '{32'h429ddf18};
test_index[9323] = '{5};
test_input[74592:74599] = '{32'hc1f45290, 32'h424bbb65, 32'hc2942410, 32'h4149ab4b, 32'hc217ecc2, 32'h41c8a358, 32'hc2ada9a7, 32'h42a529cc};
test_output[9324] = '{32'h42a529cc};
test_index[9324] = '{7};
test_input[74600:74607] = '{32'h420cd81d, 32'hc1b6e722, 32'h42361aa1, 32'hc2b4ebd1, 32'hc16b5461, 32'hc1f8b63b, 32'hc2884712, 32'h42ba06ab};
test_output[9325] = '{32'h42ba06ab};
test_index[9325] = '{7};
test_input[74608:74615] = '{32'hc24488a2, 32'hc270c278, 32'h41f8c404, 32'hc283621b, 32'hc2c08d8e, 32'hc1c916bc, 32'hc0bace32, 32'h421449b7};
test_output[9326] = '{32'h421449b7};
test_index[9326] = '{7};
test_input[74616:74623] = '{32'h4271af79, 32'h42455b53, 32'h41873265, 32'hc290f52f, 32'h429de70f, 32'hc226516e, 32'h424634dc, 32'h41cdd9ad};
test_output[9327] = '{32'h429de70f};
test_index[9327] = '{4};
test_input[74624:74631] = '{32'h42c3b8f9, 32'hc2c71c12, 32'h41945897, 32'h421e6b84, 32'h42927d12, 32'h42c0e9f7, 32'h428fdcd3, 32'hc1b67d0c};
test_output[9328] = '{32'h42c3b8f9};
test_index[9328] = '{0};
test_input[74632:74639] = '{32'hc2a52f7a, 32'hc286a633, 32'hc2a5c9a2, 32'h424e2601, 32'h4184be69, 32'h427dcb88, 32'h3e98d68e, 32'hc29904a0};
test_output[9329] = '{32'h427dcb88};
test_index[9329] = '{5};
test_input[74640:74647] = '{32'h42c1a762, 32'h42a8783f, 32'hc2be4ba5, 32'h4214a2bc, 32'hc216f56f, 32'h41c6cf1a, 32'h42262590, 32'h424d07c9};
test_output[9330] = '{32'h42c1a762};
test_index[9330] = '{0};
test_input[74648:74655] = '{32'h42192c2a, 32'h42b7eb4b, 32'hc286ca8c, 32'hc22ea069, 32'h41bf27a5, 32'h42c5c0d5, 32'hc1f67cc8, 32'hc0da9f5d};
test_output[9331] = '{32'h42c5c0d5};
test_index[9331] = '{5};
test_input[74656:74663] = '{32'h42bfd772, 32'h42942699, 32'hc21c4403, 32'h4221b0bb, 32'hc2c33dd8, 32'hc086c84f, 32'hc248f82b, 32'hc1556158};
test_output[9332] = '{32'h42bfd772};
test_index[9332] = '{0};
test_input[74664:74671] = '{32'hc2860e20, 32'h42c5a061, 32'hc1ab6160, 32'hc2985463, 32'hc226ef09, 32'h42ada3f1, 32'hc1447236, 32'h423eaa25};
test_output[9333] = '{32'h42c5a061};
test_index[9333] = '{1};
test_input[74672:74679] = '{32'h422fdff4, 32'h4210334c, 32'hc28fe66f, 32'hc28d3de7, 32'h4243f541, 32'h42a516bd, 32'h425318b9, 32'h41a6496b};
test_output[9334] = '{32'h42a516bd};
test_index[9334] = '{5};
test_input[74680:74687] = '{32'h41bf73ae, 32'h3fe57b07, 32'hc2adece0, 32'h423d9c1f, 32'h41c02ff5, 32'h42585fec, 32'h428f3d35, 32'h41a92650};
test_output[9335] = '{32'h428f3d35};
test_index[9335] = '{6};
test_input[74688:74695] = '{32'h42be3753, 32'hc06cac28, 32'hc203d26e, 32'hc22e3556, 32'h42a3f22c, 32'h42303714, 32'h42b62090, 32'h41ee607a};
test_output[9336] = '{32'h42be3753};
test_index[9336] = '{0};
test_input[74696:74703] = '{32'h425adb1b, 32'h42bbb9bf, 32'hc21fbdc4, 32'hc2c11cc0, 32'hc23f15de, 32'hc1741dea, 32'h42c7bcd9, 32'hc28ff1b1};
test_output[9337] = '{32'h42c7bcd9};
test_index[9337] = '{6};
test_input[74704:74711] = '{32'hc1f049c9, 32'hc281b18f, 32'hc2b4a6cd, 32'hc22152a4, 32'h4189fb3b, 32'hc229d155, 32'hc285771f, 32'hc2c60a75};
test_output[9338] = '{32'h4189fb3b};
test_index[9338] = '{4};
test_input[74712:74719] = '{32'h429f61b7, 32'h428df802, 32'hc2a34dc7, 32'hc29b7c1b, 32'hc1fe3cea, 32'h42b58294, 32'h4207508f, 32'hc2a42a30};
test_output[9339] = '{32'h42b58294};
test_index[9339] = '{5};
test_input[74720:74727] = '{32'h406e3521, 32'hc287927f, 32'h42075a11, 32'h4149f5a4, 32'hc18e137d, 32'h42b8e8b1, 32'h4112c0d8, 32'h42bced52};
test_output[9340] = '{32'h42bced52};
test_index[9340] = '{7};
test_input[74728:74735] = '{32'h42ace2fd, 32'h422a66b2, 32'h41f9ea2d, 32'hc2949dfc, 32'hc29ac49a, 32'hc2bcf7f8, 32'h42af9da5, 32'hc1068c2f};
test_output[9341] = '{32'h42af9da5};
test_index[9341] = '{6};
test_input[74736:74743] = '{32'hc23bbdf2, 32'h42823292, 32'h42972f2d, 32'hc21f82ba, 32'h428b7200, 32'hc205575f, 32'h42980ff9, 32'h425a7aa3};
test_output[9342] = '{32'h42980ff9};
test_index[9342] = '{6};
test_input[74744:74751] = '{32'hc1e71a77, 32'hc2114733, 32'hc26db4c6, 32'h4170f4ce, 32'hc26cca4c, 32'hc2bc70d9, 32'h429e8445, 32'hc24b09f6};
test_output[9343] = '{32'h429e8445};
test_index[9343] = '{6};
test_input[74752:74759] = '{32'h428c9add, 32'hc2ab034b, 32'h4217275e, 32'hc1e8192f, 32'hc20e4ba6, 32'hc13a0124, 32'hc297de6c, 32'hc1f1bc35};
test_output[9344] = '{32'h428c9add};
test_index[9344] = '{0};
test_input[74760:74767] = '{32'hc2c37f30, 32'hc1488787, 32'hc29f09c7, 32'hc25c7f51, 32'h422660dd, 32'h40395dba, 32'hc29712b1, 32'h426ed6f9};
test_output[9345] = '{32'h426ed6f9};
test_index[9345] = '{7};
test_input[74768:74775] = '{32'hc0912f8b, 32'hc2976fc1, 32'hbfac403a, 32'h4214375e, 32'hc229fc05, 32'hc14ff60e, 32'hc2bccc1b, 32'h42af8aac};
test_output[9346] = '{32'h42af8aac};
test_index[9346] = '{7};
test_input[74776:74783] = '{32'hc0fcedbc, 32'hc18e98bc, 32'hc0e6d85e, 32'h42adff86, 32'hc22ffaec, 32'hc17244a8, 32'h40dc1f48, 32'h428542e7};
test_output[9347] = '{32'h42adff86};
test_index[9347] = '{3};
test_input[74784:74791] = '{32'hc1dbc22c, 32'h42414626, 32'h417c4737, 32'hc284d1fd, 32'h426910e4, 32'h42572b02, 32'h42109069, 32'hc29c80e4};
test_output[9348] = '{32'h426910e4};
test_index[9348] = '{4};
test_input[74792:74799] = '{32'h42b93b32, 32'hc2aa6045, 32'hc21160d6, 32'h424f2002, 32'h41968ca4, 32'h42186cc5, 32'h40629229, 32'h41a2e7a6};
test_output[9349] = '{32'h42b93b32};
test_index[9349] = '{0};
test_input[74800:74807] = '{32'h405438a9, 32'h424a5d11, 32'h424f15a1, 32'hc285a819, 32'h42bbe6b2, 32'h42bb3072, 32'hc2613e7a, 32'h422d156a};
test_output[9350] = '{32'h42bbe6b2};
test_index[9350] = '{4};
test_input[74808:74815] = '{32'h423d9886, 32'h428d0258, 32'h4288dee2, 32'hc2a797d9, 32'hc2a54149, 32'hc28f3d63, 32'h41c97830, 32'h4292f018};
test_output[9351] = '{32'h4292f018};
test_index[9351] = '{7};
test_input[74816:74823] = '{32'h428027f4, 32'hc28ac868, 32'h42c0029b, 32'hc13c1106, 32'hc29a5f1c, 32'h3fc9f4f1, 32'h425739eb, 32'h420b58b7};
test_output[9352] = '{32'h42c0029b};
test_index[9352] = '{2};
test_input[74824:74831] = '{32'h4137f3a6, 32'hc21fa182, 32'h414c73e2, 32'hc09f8533, 32'h42a72e6a, 32'hc169cd09, 32'h4251c32e, 32'hc2a19e1b};
test_output[9353] = '{32'h42a72e6a};
test_index[9353] = '{4};
test_input[74832:74839] = '{32'hc230d434, 32'h4254d2ac, 32'hc2a5d7bd, 32'hc24e9ad8, 32'h422b53cf, 32'h422853ee, 32'h42bf7d1d, 32'h42c09183};
test_output[9354] = '{32'h42c09183};
test_index[9354] = '{7};
test_input[74840:74847] = '{32'h41884a22, 32'hc1dd70b3, 32'hc28a6b12, 32'hbf3b5660, 32'h427e816e, 32'h4205e68a, 32'h412817ab, 32'hc267ca53};
test_output[9355] = '{32'h427e816e};
test_index[9355] = '{4};
test_input[74848:74855] = '{32'hc2810a2b, 32'h422a3d0d, 32'hc22b3712, 32'h42af35c4, 32'hc28327ce, 32'h422fd8e2, 32'h411de17b, 32'hc2a8f85c};
test_output[9356] = '{32'h42af35c4};
test_index[9356] = '{3};
test_input[74856:74863] = '{32'h41bcb40c, 32'hc2291bc1, 32'hc217657e, 32'h41911df6, 32'h40cd6901, 32'hc26f0896, 32'hc083bdc3, 32'hc12bfcda};
test_output[9357] = '{32'h41bcb40c};
test_index[9357] = '{0};
test_input[74864:74871] = '{32'h409d58ff, 32'hc2a2b6e4, 32'h4275bc5c, 32'h4180735c, 32'hc2baae08, 32'hc27cb0bd, 32'h41bb79af, 32'hc18b0fef};
test_output[9358] = '{32'h4275bc5c};
test_index[9358] = '{2};
test_input[74872:74879] = '{32'hc29bb362, 32'h420e2dfc, 32'h422eb1f6, 32'hc186b789, 32'hc2a8de05, 32'h42b418d2, 32'h4225815c, 32'h42257b43};
test_output[9359] = '{32'h42b418d2};
test_index[9359] = '{5};
test_input[74880:74887] = '{32'hc23aef6b, 32'hc26d6451, 32'h4195e8d6, 32'h4286acac, 32'h42bbdb72, 32'h42041015, 32'h4065b714, 32'h42b38fea};
test_output[9360] = '{32'h42bbdb72};
test_index[9360] = '{4};
test_input[74888:74895] = '{32'h41a9e3e3, 32'h42874535, 32'h401e6ca5, 32'hc011b50a, 32'h422cf0d6, 32'h429f54df, 32'hc2200ad2, 32'h4287442e};
test_output[9361] = '{32'h429f54df};
test_index[9361] = '{5};
test_input[74896:74903] = '{32'hc25ff8f8, 32'hc2bd093f, 32'h40f96e26, 32'h42ad072d, 32'hc2a364f7, 32'hc1926a9a, 32'h425069b4, 32'hc2baf3f4};
test_output[9362] = '{32'h42ad072d};
test_index[9362] = '{3};
test_input[74904:74911] = '{32'h3fcec96e, 32'h413ed4a3, 32'h425662e7, 32'h41ffed63, 32'hc2003025, 32'h42a3fbf8, 32'h42afa8a3, 32'h425899a0};
test_output[9363] = '{32'h42afa8a3};
test_index[9363] = '{6};
test_input[74912:74919] = '{32'h42882eb3, 32'h407d06d4, 32'hc2b56e00, 32'hc17e19b3, 32'h4283997e, 32'h410cf6b6, 32'h428cab29, 32'h42ae184a};
test_output[9364] = '{32'h42ae184a};
test_index[9364] = '{7};
test_input[74920:74927] = '{32'h42bd071c, 32'hc239c5fb, 32'h427d6baf, 32'h41ef74ae, 32'hc1e7ca67, 32'hc205bc27, 32'hc2252aa8, 32'hc208d5af};
test_output[9365] = '{32'h42bd071c};
test_index[9365] = '{0};
test_input[74928:74935] = '{32'hc2984a55, 32'hc2a34222, 32'hc17cbbff, 32'h42b7ea89, 32'hc2add51b, 32'hc29174ec, 32'h41e96360, 32'h40d861e6};
test_output[9366] = '{32'h42b7ea89};
test_index[9366] = '{3};
test_input[74936:74943] = '{32'hc0a9f8bf, 32'h42af7f33, 32'h41fb3fee, 32'h41bcb90a, 32'h42a1792d, 32'h420f2523, 32'hc29529d5, 32'h418eec0c};
test_output[9367] = '{32'h42af7f33};
test_index[9367] = '{1};
test_input[74944:74951] = '{32'h418d315c, 32'hc2c60c1c, 32'h3f36111a, 32'h404e96e9, 32'h425bc5fd, 32'h424026f7, 32'hc2bd38c6, 32'h41d199d0};
test_output[9368] = '{32'h425bc5fd};
test_index[9368] = '{4};
test_input[74952:74959] = '{32'hc2c7f888, 32'h429f1342, 32'h41ba673f, 32'h418f6ed6, 32'h4298872c, 32'h41535cf5, 32'hc27a33ae, 32'h4226a167};
test_output[9369] = '{32'h429f1342};
test_index[9369] = '{1};
test_input[74960:74967] = '{32'h4116402e, 32'hc1f1ee12, 32'h4245bfaa, 32'h425edff8, 32'hc16e4dc0, 32'h4153a11d, 32'hc24e5aba, 32'h42429e05};
test_output[9370] = '{32'h425edff8};
test_index[9370] = '{3};
test_input[74968:74975] = '{32'hc2b25409, 32'h425dee5b, 32'h42c7a0cb, 32'h42b9ca62, 32'hc28f162f, 32'h412123a1, 32'hc289cc9c, 32'h41e361b9};
test_output[9371] = '{32'h42c7a0cb};
test_index[9371] = '{2};
test_input[74976:74983] = '{32'hc23df179, 32'h4251af06, 32'h4195e7ac, 32'hc1abc5eb, 32'h4125c330, 32'h42c2a551, 32'h42a0f7f4, 32'hc272ac40};
test_output[9372] = '{32'h42c2a551};
test_index[9372] = '{5};
test_input[74984:74991] = '{32'h42b0e0fa, 32'h42995830, 32'hc29ca0e4, 32'hc29fbdaa, 32'h4281eddc, 32'hc2581d72, 32'hc2a2eed2, 32'h4068cfa6};
test_output[9373] = '{32'h42b0e0fa};
test_index[9373] = '{0};
test_input[74992:74999] = '{32'h42b2743e, 32'hc2c0fb61, 32'hc1a066be, 32'hc2a41def, 32'h42873f76, 32'h4286e4b3, 32'h41c2a078, 32'h4211a325};
test_output[9374] = '{32'h42b2743e};
test_index[9374] = '{0};
test_input[75000:75007] = '{32'hc2609520, 32'hc19842ca, 32'h425c9137, 32'h428b98e7, 32'hc0e5352f, 32'h42b5a695, 32'hc235af5d, 32'h3f3b9b43};
test_output[9375] = '{32'h42b5a695};
test_index[9375] = '{5};
test_input[75008:75015] = '{32'h42b2ad2c, 32'hc21ecd97, 32'hc29676bd, 32'hc165b546, 32'h42bc4317, 32'h42c21174, 32'hc19a2502, 32'hc1ceb643};
test_output[9376] = '{32'h42c21174};
test_index[9376] = '{5};
test_input[75016:75023] = '{32'h426cd1e0, 32'h429278a5, 32'h41f5eed0, 32'h42a003c2, 32'h405f7d92, 32'hc1925e16, 32'h4272e20c, 32'hc2b118b7};
test_output[9377] = '{32'h42a003c2};
test_index[9377] = '{3};
test_input[75024:75031] = '{32'hc25187dd, 32'h3ff146dc, 32'h425cc37e, 32'hc28ad88b, 32'h425df7fe, 32'hc126c955, 32'hc2b57d9b, 32'h4242a169};
test_output[9378] = '{32'h425df7fe};
test_index[9378] = '{4};
test_input[75032:75039] = '{32'h42c62c0d, 32'h42c5ac9d, 32'hc1cdacc4, 32'hc2c68066, 32'h41de56de, 32'h41011b7f, 32'hc2ad53dd, 32'hc187157c};
test_output[9379] = '{32'h42c62c0d};
test_index[9379] = '{0};
test_input[75040:75047] = '{32'hc225b035, 32'hc2c693f5, 32'h422c64eb, 32'hc2c3a99d, 32'hc1eb74c3, 32'h425213d9, 32'h415cb7c9, 32'h4130e15c};
test_output[9380] = '{32'h425213d9};
test_index[9380] = '{5};
test_input[75048:75055] = '{32'hc107e3c0, 32'h42b483d6, 32'hc1d95f51, 32'hc1c4199b, 32'h423ba3db, 32'h42a8432c, 32'hc2811e7a, 32'hc24f0b3e};
test_output[9381] = '{32'h42b483d6};
test_index[9381] = '{1};
test_input[75056:75063] = '{32'hc1c731ea, 32'h422a055f, 32'h41853ef4, 32'hc1c34b62, 32'hc188a154, 32'hc1a03771, 32'h42afe700, 32'hc26b17dd};
test_output[9382] = '{32'h42afe700};
test_index[9382] = '{6};
test_input[75064:75071] = '{32'h418ef68e, 32'hc276134d, 32'hc1ea92aa, 32'hc09062d4, 32'hc2ac412d, 32'hc1f35e7b, 32'hc257d3ed, 32'hc2aebd7d};
test_output[9383] = '{32'h418ef68e};
test_index[9383] = '{0};
test_input[75072:75079] = '{32'hc251e15c, 32'h42b39388, 32'hc263801c, 32'hc2a866a5, 32'h4291c598, 32'h42a5ca87, 32'hc27b6d23, 32'hc22eb3d9};
test_output[9384] = '{32'h42b39388};
test_index[9384] = '{1};
test_input[75080:75087] = '{32'h422d78cc, 32'hc28fb6a9, 32'hc21fd9af, 32'h4230efa7, 32'hc2343174, 32'hc191e644, 32'h42b863ac, 32'h42c5f357};
test_output[9385] = '{32'h42c5f357};
test_index[9385] = '{7};
test_input[75088:75095] = '{32'hc1a9855e, 32'h4207e1d0, 32'hc26f05b2, 32'h422c325f, 32'h42bd5729, 32'h41e740a1, 32'h419fae13, 32'hc283f5f7};
test_output[9386] = '{32'h42bd5729};
test_index[9386] = '{4};
test_input[75096:75103] = '{32'hc2300135, 32'h4206bb4c, 32'h416896b3, 32'h3f8fb737, 32'hc28bdf44, 32'h4280a28c, 32'h427260b7, 32'hc1a20c9f};
test_output[9387] = '{32'h4280a28c};
test_index[9387] = '{5};
test_input[75104:75111] = '{32'h41e0d5a9, 32'h424cdcbf, 32'hc213822b, 32'h425c2215, 32'h429f65c4, 32'hc199c298, 32'hc22ff2af, 32'hc261012b};
test_output[9388] = '{32'h429f65c4};
test_index[9388] = '{4};
test_input[75112:75119] = '{32'h405a7eb4, 32'h41717b79, 32'hc1e44db2, 32'h42b9c5b3, 32'hc20d6a13, 32'hc1a520ee, 32'h42938501, 32'hc18b166d};
test_output[9389] = '{32'h42b9c5b3};
test_index[9389] = '{3};
test_input[75120:75127] = '{32'hc2991c24, 32'hc242e037, 32'hc2336a0c, 32'hc2a8fc52, 32'h423058de, 32'h4183d145, 32'h42947d9b, 32'h4293b4ed};
test_output[9390] = '{32'h42947d9b};
test_index[9390] = '{6};
test_input[75128:75135] = '{32'h424e99d2, 32'h4262c3b2, 32'h428d9578, 32'h4247afd3, 32'hc226070f, 32'h40994a01, 32'h41871d18, 32'hc20bf30d};
test_output[9391] = '{32'h428d9578};
test_index[9391] = '{2};
test_input[75136:75143] = '{32'h42ac47b1, 32'h425e6316, 32'h41dece7b, 32'h426794d9, 32'h427f25af, 32'h41969dcf, 32'h42771f1d, 32'hc224ff1c};
test_output[9392] = '{32'h42ac47b1};
test_index[9392] = '{0};
test_input[75144:75151] = '{32'h42a148e0, 32'hc27c7cb8, 32'h424e0441, 32'h413e907e, 32'hc29e143b, 32'hc28d928c, 32'h42229d51, 32'h3e840f76};
test_output[9393] = '{32'h42a148e0};
test_index[9393] = '{0};
test_input[75152:75159] = '{32'hc293f65c, 32'hc285df27, 32'hc280e95e, 32'h415ff8f8, 32'hc24aeb71, 32'hc2261ff4, 32'h424cc03a, 32'hc1d45930};
test_output[9394] = '{32'h424cc03a};
test_index[9394] = '{6};
test_input[75160:75167] = '{32'hc2228a3d, 32'hc2a38219, 32'h421a4b64, 32'h416095e5, 32'h41a84626, 32'h42a09c21, 32'hc23e3ec8, 32'h42bb2daf};
test_output[9395] = '{32'h42bb2daf};
test_index[9395] = '{7};
test_input[75168:75175] = '{32'hc22f0f24, 32'h42a1c395, 32'hc26c889c, 32'hc1b051b6, 32'hc18398b9, 32'h400ee7d1, 32'hc2865bda, 32'hc1f2bcc2};
test_output[9396] = '{32'h42a1c395};
test_index[9396] = '{1};
test_input[75176:75183] = '{32'hc14475ef, 32'hc2767507, 32'hc127149e, 32'h42807f9d, 32'hc2312a70, 32'hc2718567, 32'h4113c7c8, 32'hc2536758};
test_output[9397] = '{32'h42807f9d};
test_index[9397] = '{3};
test_input[75184:75191] = '{32'hc2b98195, 32'h42ba99a4, 32'h42a0e6c8, 32'hc24485ef, 32'h4289dd57, 32'h41102d95, 32'hc235b689, 32'hc286fc47};
test_output[9398] = '{32'h42ba99a4};
test_index[9398] = '{1};
test_input[75192:75199] = '{32'h4232c6b8, 32'hc1e998b1, 32'hc2c3c9a0, 32'h42223787, 32'h4210f053, 32'hc2487146, 32'hc287432f, 32'h4253b0f0};
test_output[9399] = '{32'h4253b0f0};
test_index[9399] = '{7};
test_input[75200:75207] = '{32'h41d5d9dc, 32'hc1ca359a, 32'hc1eab2bf, 32'h42bf24e2, 32'hc259ed5c, 32'h4182bc43, 32'h42bbca9b, 32'h3f4cd7c6};
test_output[9400] = '{32'h42bf24e2};
test_index[9400] = '{3};
test_input[75208:75215] = '{32'hc298e0b4, 32'hc2a2b87d, 32'hc2b06bac, 32'hc27d05f9, 32'h42165c6c, 32'hc139a9c2, 32'h42a586d8, 32'hc2482d38};
test_output[9401] = '{32'h42a586d8};
test_index[9401] = '{6};
test_input[75216:75223] = '{32'hc24d1501, 32'hc1a22708, 32'hc22935b9, 32'hc1bf8a35, 32'hc29965bf, 32'hc289c597, 32'h4233eb1a, 32'h42abb87e};
test_output[9402] = '{32'h42abb87e};
test_index[9402] = '{7};
test_input[75224:75231] = '{32'hc2235b6b, 32'hc2c27937, 32'h41b1c184, 32'h42c20b16, 32'hc20c6ffb, 32'hc2a093da, 32'hc2034eba, 32'hc2c007ad};
test_output[9403] = '{32'h42c20b16};
test_index[9403] = '{3};
test_input[75232:75239] = '{32'hc1c04b23, 32'hc1f72758, 32'h4297a427, 32'h41f9a27f, 32'h42ac7b49, 32'h4230a680, 32'hc29b6e4c, 32'h426f6043};
test_output[9404] = '{32'h42ac7b49};
test_index[9404] = '{4};
test_input[75240:75247] = '{32'hc2a24c49, 32'h4268f6ec, 32'hc18ca320, 32'h42b542f3, 32'hc2a5938a, 32'hc28729e8, 32'h4141eaf0, 32'h429c2341};
test_output[9405] = '{32'h42b542f3};
test_index[9405] = '{3};
test_input[75248:75255] = '{32'hc2ae341f, 32'hc282dfc6, 32'hc2685c93, 32'hc2b00082, 32'h422eeb88, 32'h41a26d34, 32'hc26f208b, 32'h42660b0a};
test_output[9406] = '{32'h42660b0a};
test_index[9406] = '{7};
test_input[75256:75263] = '{32'h41f688ab, 32'h42b2f8c5, 32'hc242f3e0, 32'hc1de2ea7, 32'h4296c617, 32'h41360fa1, 32'h41dc1c8d, 32'h41a0e443};
test_output[9407] = '{32'h42b2f8c5};
test_index[9407] = '{1};
test_input[75264:75271] = '{32'hc2c5c0a7, 32'h4270424d, 32'h42062ecd, 32'hc2001e43, 32'hc16f8488, 32'hc14f2f6c, 32'h427db157, 32'h40ba2d01};
test_output[9408] = '{32'h427db157};
test_index[9408] = '{6};
test_input[75272:75279] = '{32'h421600f1, 32'hc2a3c035, 32'hc230bea3, 32'hc2a8e31b, 32'h42839121, 32'h426cfedd, 32'hc20a9023, 32'hc29c1c6a};
test_output[9409] = '{32'h42839121};
test_index[9409] = '{4};
test_input[75280:75287] = '{32'hc1f63f6e, 32'hc28537b6, 32'h42b4c39e, 32'h4285a6c2, 32'hc1bd5f1d, 32'hc28d91b3, 32'h425bd926, 32'h41b43839};
test_output[9410] = '{32'h42b4c39e};
test_index[9410] = '{2};
test_input[75288:75295] = '{32'h429cec9c, 32'h4010bb4d, 32'h425d347c, 32'h414fa75f, 32'hc2a9ee39, 32'hc23558fc, 32'h42ad48aa, 32'hc012ee03};
test_output[9411] = '{32'h42ad48aa};
test_index[9411] = '{6};
test_input[75296:75303] = '{32'h42aca571, 32'h4220a9b1, 32'hc28cb213, 32'hc18322ad, 32'h42af1ede, 32'h404be931, 32'hc23cc1ea, 32'h41b327df};
test_output[9412] = '{32'h42af1ede};
test_index[9412] = '{4};
test_input[75304:75311] = '{32'hc2684427, 32'h4291980f, 32'h4298bba6, 32'hc26a98cb, 32'hc1da2a9d, 32'hc15866c2, 32'hc299966b, 32'hc2a42a1d};
test_output[9413] = '{32'h4298bba6};
test_index[9413] = '{2};
test_input[75312:75319] = '{32'hc2985d46, 32'h42bb5d3d, 32'hc26aab1b, 32'h41eef053, 32'hc2b4f572, 32'h424bc105, 32'h429e77e1, 32'hc24744f4};
test_output[9414] = '{32'h42bb5d3d};
test_index[9414] = '{1};
test_input[75320:75327] = '{32'hc259139b, 32'hc1a5c45b, 32'h42951132, 32'hc2946e72, 32'h424e94ed, 32'h4192e405, 32'h42c3b64d, 32'h41e324c9};
test_output[9415] = '{32'h42c3b64d};
test_index[9415] = '{6};
test_input[75328:75335] = '{32'hc1e7532a, 32'hc194575e, 32'hc29f7aac, 32'h42b11546, 32'hc2963624, 32'hc20e4fc2, 32'h41734b1c, 32'hc266e06a};
test_output[9416] = '{32'h42b11546};
test_index[9416] = '{3};
test_input[75336:75343] = '{32'h4206985c, 32'h424e37e5, 32'h40825474, 32'h4296619d, 32'hc1122076, 32'h42a4edc9, 32'hc208a46b, 32'hc1c4fe6a};
test_output[9417] = '{32'h42a4edc9};
test_index[9417] = '{5};
test_input[75344:75351] = '{32'h42451909, 32'hc2a06fed, 32'hc1096703, 32'h40905940, 32'h429dfc68, 32'h41fd2e01, 32'h42426406, 32'hc2bec128};
test_output[9418] = '{32'h429dfc68};
test_index[9418] = '{4};
test_input[75352:75359] = '{32'h4296e02d, 32'h424bedcd, 32'hc29da753, 32'h411fd77e, 32'hc1e2e383, 32'hc29dc353, 32'h423976f1, 32'hc29f38c1};
test_output[9419] = '{32'h4296e02d};
test_index[9419] = '{0};
test_input[75360:75367] = '{32'h422b3b8a, 32'h42acd194, 32'hc2781998, 32'h414dc533, 32'h42bc64a1, 32'h420d1e9f, 32'hc235e37c, 32'hc2c769dd};
test_output[9420] = '{32'h42bc64a1};
test_index[9420] = '{4};
test_input[75368:75375] = '{32'hc2c571d4, 32'hc1bc9455, 32'h42b93d69, 32'h40d752ab, 32'hc2828de8, 32'h42a54021, 32'hc20f7f89, 32'hc031a48e};
test_output[9421] = '{32'h42b93d69};
test_index[9421] = '{2};
test_input[75376:75383] = '{32'hc2bda077, 32'h419ef7b0, 32'hc1eb0df0, 32'h41d6e417, 32'hc2631966, 32'hc1dacefd, 32'hc226731d, 32'h41932817};
test_output[9422] = '{32'h41d6e417};
test_index[9422] = '{3};
test_input[75384:75391] = '{32'h4280d389, 32'hc29c845a, 32'hc28899d1, 32'h42b086df, 32'hc0c1b6f2, 32'h428170db, 32'hc2b76575, 32'hc2273fb4};
test_output[9423] = '{32'h42b086df};
test_index[9423] = '{3};
test_input[75392:75399] = '{32'hc1c9b52e, 32'h4154c139, 32'h41574a1f, 32'h4215b722, 32'h426de746, 32'h42b7db9f, 32'hc2be7c74, 32'h422a3ae2};
test_output[9424] = '{32'h42b7db9f};
test_index[9424] = '{5};
test_input[75400:75407] = '{32'hc0c25fcf, 32'hc28a6509, 32'h427026e4, 32'hc29aeec2, 32'h4298127f, 32'h4199dda8, 32'h42947a57, 32'hc28d6691};
test_output[9425] = '{32'h4298127f};
test_index[9425] = '{4};
test_input[75408:75415] = '{32'hc208a51b, 32'hc12ff9ee, 32'h417d170a, 32'h42aa56ed, 32'hc1bfce7e, 32'hc2529cf3, 32'h425d020f, 32'h42c7e1e6};
test_output[9426] = '{32'h42c7e1e6};
test_index[9426] = '{7};
test_input[75416:75423] = '{32'hc16f0caf, 32'hc29c0650, 32'h42478c40, 32'hc1a4918a, 32'hc227e469, 32'hc2b4f6ab, 32'h41c30633, 32'h42c656bb};
test_output[9427] = '{32'h42c656bb};
test_index[9427] = '{7};
test_input[75424:75431] = '{32'h42857ae2, 32'h42081862, 32'h411c3a87, 32'hc212bd6c, 32'hc2511041, 32'hc277ad38, 32'hc286ba46, 32'h42a1ed7e};
test_output[9428] = '{32'h42a1ed7e};
test_index[9428] = '{7};
test_input[75432:75439] = '{32'hc2ac39a3, 32'hc2a47860, 32'h4144a1ec, 32'h42689694, 32'hc246bc0c, 32'hc2a58485, 32'h42295845, 32'h4291557e};
test_output[9429] = '{32'h4291557e};
test_index[9429] = '{7};
test_input[75440:75447] = '{32'h426d8c96, 32'hc1e2ae6c, 32'hc1cafbc5, 32'hc20655b8, 32'hc268b1bb, 32'hc2a0332f, 32'h42588966, 32'hc2325f40};
test_output[9430] = '{32'h426d8c96};
test_index[9430] = '{0};
test_input[75448:75455] = '{32'h41a3a7cd, 32'h425a77d4, 32'hc1e6947c, 32'hc0f162c4, 32'hc2a5755e, 32'hc1e5d79b, 32'hc0fbfe98, 32'h425892e5};
test_output[9431] = '{32'h425a77d4};
test_index[9431] = '{1};
test_input[75456:75463] = '{32'hc1d0e4bd, 32'hc24fa1b4, 32'h42638afe, 32'h40ce277b, 32'hc229862d, 32'hc2bceaa0, 32'h4126d053, 32'hc2947948};
test_output[9432] = '{32'h42638afe};
test_index[9432] = '{2};
test_input[75464:75471] = '{32'h42b5c610, 32'hc26c2766, 32'hc0019381, 32'h4100d4ce, 32'h40d3457a, 32'h418c284a, 32'hc27fc565, 32'h4294e6d3};
test_output[9433] = '{32'h42b5c610};
test_index[9433] = '{0};
test_input[75472:75479] = '{32'h4254d709, 32'h41fd599e, 32'hc16fdfc7, 32'h4183db24, 32'hc2608b66, 32'hc13b0aba, 32'h42722cf7, 32'hc12a7d9e};
test_output[9434] = '{32'h42722cf7};
test_index[9434] = '{6};
test_input[75480:75487] = '{32'h41d301a0, 32'h41d82a73, 32'h41ee6c74, 32'h41db2f7f, 32'hc0f15a10, 32'hc1418cee, 32'hc2141aa7, 32'h424abb58};
test_output[9435] = '{32'h424abb58};
test_index[9435] = '{7};
test_input[75488:75495] = '{32'hc17d24bb, 32'hc1e19d8b, 32'hc1b5d980, 32'h42be3ce5, 32'h41a019c8, 32'h42bbe3e3, 32'hc24fc9a0, 32'hc2844c46};
test_output[9436] = '{32'h42be3ce5};
test_index[9436] = '{3};
test_input[75496:75503] = '{32'h41811067, 32'h42725687, 32'hc22fbacc, 32'hc1caa0f4, 32'hc2b9cb93, 32'h429c15bd, 32'h42a79652, 32'h42b050a4};
test_output[9437] = '{32'h42b050a4};
test_index[9437] = '{7};
test_input[75504:75511] = '{32'hc235a9b2, 32'hc1e76a31, 32'h416479d8, 32'h4227e153, 32'h4224d13e, 32'hc2ace9f8, 32'h42abc6e1, 32'h40a59a8a};
test_output[9438] = '{32'h42abc6e1};
test_index[9438] = '{6};
test_input[75512:75519] = '{32'hc280c3d6, 32'h427752ba, 32'hc18c5dfe, 32'h426f8cf4, 32'h4084f995, 32'hc199caa9, 32'hc29b9afc, 32'hc291086c};
test_output[9439] = '{32'h427752ba};
test_index[9439] = '{1};
test_input[75520:75527] = '{32'hc2bb8f8e, 32'hc190ee3a, 32'hc28f2845, 32'hc1727bd4, 32'hc09eb632, 32'hc2c107bb, 32'h427e1bfe, 32'h419d1012};
test_output[9440] = '{32'h427e1bfe};
test_index[9440] = '{6};
test_input[75528:75535] = '{32'hc220bf94, 32'hc2191bbd, 32'hc1b99db7, 32'h422fb5a0, 32'h41d88c6c, 32'h42ad9965, 32'h4234bccf, 32'h41f33079};
test_output[9441] = '{32'h42ad9965};
test_index[9441] = '{5};
test_input[75536:75543] = '{32'hc14ee168, 32'hc21322fa, 32'h4204190f, 32'hc1dc9e88, 32'hc2a22f05, 32'hc2accd2d, 32'hc2908510, 32'hc29f691a};
test_output[9442] = '{32'h4204190f};
test_index[9442] = '{2};
test_input[75544:75551] = '{32'h42835d13, 32'h414d0c5b, 32'hc2331b4c, 32'h404c5a94, 32'hc15a7bd9, 32'hc1f46443, 32'hc2005761, 32'hc2884683};
test_output[9443] = '{32'h42835d13};
test_index[9443] = '{0};
test_input[75552:75559] = '{32'hc249405a, 32'h42ba270e, 32'h4136c033, 32'h41aadfcf, 32'h423ce606, 32'h4236a7e7, 32'h410025c7, 32'h420e5bac};
test_output[9444] = '{32'h42ba270e};
test_index[9444] = '{1};
test_input[75560:75567] = '{32'hc075c6e0, 32'h3f1627f1, 32'hc228956f, 32'hc06cf38b, 32'h3fbbf65b, 32'hc2872c19, 32'hc2a218d8, 32'hc28bc44a};
test_output[9445] = '{32'h3fbbf65b};
test_index[9445] = '{4};
test_input[75568:75575] = '{32'h423ae951, 32'hc223070f, 32'hc1908016, 32'hc193e7bc, 32'hc2b0aca6, 32'h4233ae3e, 32'h423e5b0b, 32'hc2225c51};
test_output[9446] = '{32'h423e5b0b};
test_index[9446] = '{6};
test_input[75576:75583] = '{32'h42b8f875, 32'hc262e693, 32'hc08d5478, 32'h42b2103c, 32'hbfd766fd, 32'h418216ae, 32'h4280f12d, 32'hc20adfc6};
test_output[9447] = '{32'h42b8f875};
test_index[9447] = '{0};
test_input[75584:75591] = '{32'h42a64807, 32'h42a05981, 32'h4233a12e, 32'h42110a34, 32'h425bab69, 32'h425d27c3, 32'h411d301b, 32'h4220a0b6};
test_output[9448] = '{32'h42a64807};
test_index[9448] = '{0};
test_input[75592:75599] = '{32'h4160c138, 32'hc28499df, 32'hbec30f58, 32'hc2833247, 32'hc23802db, 32'h42a8a652, 32'h42a95b17, 32'h422a7adf};
test_output[9449] = '{32'h42a95b17};
test_index[9449] = '{6};
test_input[75600:75607] = '{32'h42acb2e5, 32'h41c3afb8, 32'hc28da174, 32'hc1a2f0b6, 32'hc25953ae, 32'h42acf387, 32'hc2acb6b7, 32'hc2818839};
test_output[9450] = '{32'h42acf387};
test_index[9450] = '{5};
test_input[75608:75615] = '{32'h42468ed9, 32'h42037656, 32'hc0e62700, 32'hc26f8552, 32'hc1544ebc, 32'h420f3eb4, 32'hc1c2dc89, 32'h41c007c8};
test_output[9451] = '{32'h42468ed9};
test_index[9451] = '{0};
test_input[75616:75623] = '{32'hc21a2405, 32'h42857049, 32'hc1f3279e, 32'h41c7eb63, 32'h4282894e, 32'h4259e576, 32'h410dd5d8, 32'h4173d0c6};
test_output[9452] = '{32'h42857049};
test_index[9452] = '{1};
test_input[75624:75631] = '{32'hc18e2cf5, 32'h41ec8808, 32'hbee16794, 32'hc26cc6e7, 32'hc290c605, 32'hc2c3178f, 32'hc2adf0e5, 32'h4291a597};
test_output[9453] = '{32'h4291a597};
test_index[9453] = '{7};
test_input[75632:75639] = '{32'hc22eaaba, 32'h410a0115, 32'h41fb02da, 32'h42aa30ee, 32'hc282451d, 32'hc27b4f46, 32'h425bc30a, 32'h429ed52f};
test_output[9454] = '{32'h42aa30ee};
test_index[9454] = '{3};
test_input[75640:75647] = '{32'hc2c4d728, 32'hc2859dd0, 32'h42949bdd, 32'h428ab3c4, 32'hc2a8ba1d, 32'hc28bd1cb, 32'hc1cce737, 32'hc21c052e};
test_output[9455] = '{32'h42949bdd};
test_index[9455] = '{2};
test_input[75648:75655] = '{32'h4281d317, 32'h428b71d9, 32'h418660c6, 32'h427b3508, 32'h42a1faba, 32'hc254eb9d, 32'h40c98831, 32'h428da87e};
test_output[9456] = '{32'h42a1faba};
test_index[9456] = '{4};
test_input[75656:75663] = '{32'h4190054c, 32'hc25fa6a9, 32'hc1b5a904, 32'hc206ce64, 32'hc1d07dd9, 32'hc2b71846, 32'h4297d697, 32'h4147dc62};
test_output[9457] = '{32'h4297d697};
test_index[9457] = '{6};
test_input[75664:75671] = '{32'h41624f3f, 32'h42358814, 32'h42937bb2, 32'h4275d540, 32'hc1c3d00b, 32'hc29d3457, 32'hc24a7365, 32'h42565309};
test_output[9458] = '{32'h42937bb2};
test_index[9458] = '{2};
test_input[75672:75679] = '{32'hc1a101a6, 32'h42bd0741, 32'h423f73e7, 32'h42adf808, 32'h425a5a3c, 32'hc203c692, 32'hc216f044, 32'hc283e566};
test_output[9459] = '{32'h42bd0741};
test_index[9459] = '{1};
test_input[75680:75687] = '{32'h42aee5f3, 32'h421e400d, 32'h40951b23, 32'hc285fb2d, 32'h41642368, 32'hc25bc99b, 32'h42b724e1, 32'hc28117d6};
test_output[9460] = '{32'h42b724e1};
test_index[9460] = '{6};
test_input[75688:75695] = '{32'hc23ab178, 32'hc2c123b8, 32'hc1f8c3fb, 32'hc2b7bca5, 32'h421f79d9, 32'hc23e1f0a, 32'hc2694ace, 32'h4155fe1d};
test_output[9461] = '{32'h421f79d9};
test_index[9461] = '{4};
test_input[75696:75703] = '{32'hc21f3b30, 32'h3fd94e89, 32'hc26f3f00, 32'hc2800b52, 32'h41c7e3ad, 32'hc2890256, 32'h428e413a, 32'hc270d576};
test_output[9462] = '{32'h428e413a};
test_index[9462] = '{6};
test_input[75704:75711] = '{32'h42c36382, 32'h4228c67c, 32'h425b28b1, 32'hc25e5cf9, 32'hc0d77a95, 32'h41ce0b8f, 32'hc14e63b3, 32'hc243fdff};
test_output[9463] = '{32'h42c36382};
test_index[9463] = '{0};
test_input[75712:75719] = '{32'h429c913e, 32'hc2c50885, 32'h4225c2c0, 32'hc2b78a7d, 32'h4257bd78, 32'h4288fc8a, 32'h41940ba5, 32'h428decf0};
test_output[9464] = '{32'h429c913e};
test_index[9464] = '{0};
test_input[75720:75727] = '{32'hc0de3091, 32'hc2bd181f, 32'hc1603293, 32'hc2874d80, 32'hc1d78e5b, 32'hc0e68912, 32'h4294d5f2, 32'h412f088d};
test_output[9465] = '{32'h4294d5f2};
test_index[9465] = '{6};
test_input[75728:75735] = '{32'h41cf1733, 32'hc21e7341, 32'hc22a200d, 32'h4283ee23, 32'hc1e0c91b, 32'h42916cd8, 32'h415018b3, 32'hc252dcdc};
test_output[9466] = '{32'h42916cd8};
test_index[9466] = '{5};
test_input[75736:75743] = '{32'hc27d645a, 32'h42b94d96, 32'hc1d3d9f1, 32'hc1b360ef, 32'hc29275a1, 32'hc2b3757d, 32'h423cf571, 32'hc1eae01a};
test_output[9467] = '{32'h42b94d96};
test_index[9467] = '{1};
test_input[75744:75751] = '{32'h428006d7, 32'hc29253a2, 32'hc245e961, 32'hc1df9ca8, 32'h41c8a2ae, 32'h427c743e, 32'h4110ab47, 32'hc2b8ae2a};
test_output[9468] = '{32'h428006d7};
test_index[9468] = '{0};
test_input[75752:75759] = '{32'h41f51599, 32'h41e35798, 32'h410f5fa0, 32'h419c5b17, 32'h40bae614, 32'hc2b0343a, 32'hc28f4af9, 32'hc28ed754};
test_output[9469] = '{32'h41f51599};
test_index[9469] = '{0};
test_input[75760:75767] = '{32'hc28e214c, 32'hc2bb6b60, 32'h42659bfc, 32'hc2ba0518, 32'hc20a8743, 32'h428abefd, 32'h42c508ad, 32'h41bc5aef};
test_output[9470] = '{32'h42c508ad};
test_index[9470] = '{6};
test_input[75768:75775] = '{32'hc1ce1045, 32'hc26002d2, 32'h418662dd, 32'h40ea62b7, 32'hc298a751, 32'h423ecf6d, 32'h41fd6fa3, 32'hc2916ba7};
test_output[9471] = '{32'h423ecf6d};
test_index[9471] = '{5};
test_input[75776:75783] = '{32'h4224140b, 32'hc09e1f7a, 32'h42ae1b58, 32'hc23e45e2, 32'h42a55a61, 32'h41cb824c, 32'h42b98d35, 32'h42be9d20};
test_output[9472] = '{32'h42be9d20};
test_index[9472] = '{7};
test_input[75784:75791] = '{32'h422a6eb3, 32'hc1f737a3, 32'hc15aa236, 32'hc1561fd1, 32'h4206c87a, 32'h426d2ceb, 32'h41a8719f, 32'h4213936e};
test_output[9473] = '{32'h426d2ceb};
test_index[9473] = '{5};
test_input[75792:75799] = '{32'hc0db2b60, 32'hc0cd9d4e, 32'h4211b4da, 32'h42364bb2, 32'hc29aed74, 32'h410f5fb9, 32'hc09079a8, 32'h424a7447};
test_output[9474] = '{32'h424a7447};
test_index[9474] = '{7};
test_input[75800:75807] = '{32'h4085f3e7, 32'h42ad08dd, 32'hc223a461, 32'hc207c415, 32'hc29314d3, 32'h418e8dc6, 32'h42bf836f, 32'h4216d41b};
test_output[9475] = '{32'h42bf836f};
test_index[9475] = '{6};
test_input[75808:75815] = '{32'h42065078, 32'h421093ce, 32'hc2131768, 32'h429a158f, 32'hc288a15e, 32'h418b1b2f, 32'h4127112d, 32'hc22aa0cb};
test_output[9476] = '{32'h429a158f};
test_index[9476] = '{3};
test_input[75816:75823] = '{32'hc241a542, 32'hc289e184, 32'h4180121b, 32'h42aef49a, 32'hc2c14931, 32'h4209e327, 32'hc160f1ca, 32'h42929b37};
test_output[9477] = '{32'h42aef49a};
test_index[9477] = '{3};
test_input[75824:75831] = '{32'hc2b9a6d0, 32'h42596729, 32'h428d6aef, 32'hc29ac571, 32'h41a4f367, 32'hc28dfa58, 32'h420c36da, 32'h41b84592};
test_output[9478] = '{32'h428d6aef};
test_index[9478] = '{2};
test_input[75832:75839] = '{32'h42a58dd9, 32'h42b3a99d, 32'h41a9ac3d, 32'h410f7daa, 32'h4204e24e, 32'hc2b34aaf, 32'hc2b876ea, 32'hc297d171};
test_output[9479] = '{32'h42b3a99d};
test_index[9479] = '{1};
test_input[75840:75847] = '{32'hc21f95b6, 32'h422c1df5, 32'h42159d55, 32'hc158f0cd, 32'hc18b77a0, 32'hc20c4de3, 32'hc286b71d, 32'hc1eb643f};
test_output[9480] = '{32'h422c1df5};
test_index[9480] = '{1};
test_input[75848:75855] = '{32'h40012a64, 32'hc2459736, 32'hc2425279, 32'h42bae7d6, 32'hc1c88e08, 32'h41b8a9a7, 32'hc0c0e3e7, 32'h42295187};
test_output[9481] = '{32'h42bae7d6};
test_index[9481] = '{3};
test_input[75856:75863] = '{32'hc2832153, 32'h42b2726e, 32'h4286b676, 32'h4297c192, 32'hc2446800, 32'h42890e24, 32'h429d0515, 32'h424a9c5f};
test_output[9482] = '{32'h42b2726e};
test_index[9482] = '{1};
test_input[75864:75871] = '{32'hc2c75568, 32'hc2531ff3, 32'hc282ff39, 32'hc2b32b6d, 32'hc15a1bbd, 32'hc1c7270b, 32'hc198f94b, 32'h42aca5e7};
test_output[9483] = '{32'h42aca5e7};
test_index[9483] = '{7};
test_input[75872:75879] = '{32'hc2990946, 32'hc1a2bf9a, 32'h42b9bedb, 32'hc21e3964, 32'h426780ca, 32'hc2a26825, 32'hc270d674, 32'h4269b230};
test_output[9484] = '{32'h42b9bedb};
test_index[9484] = '{2};
test_input[75880:75887] = '{32'hc1bf846f, 32'hc1af398e, 32'h420d1ba7, 32'hc1bed313, 32'h3d8baf47, 32'hc2521f07, 32'h427ca30c, 32'h428b8a6d};
test_output[9485] = '{32'h428b8a6d};
test_index[9485] = '{7};
test_input[75888:75895] = '{32'hc14bd02f, 32'hc1bb88cb, 32'h418be9f7, 32'hc23e8e98, 32'hc283055d, 32'hbf3ddbf4, 32'h4143fada, 32'hc1f2b46e};
test_output[9486] = '{32'h418be9f7};
test_index[9486] = '{2};
test_input[75896:75903] = '{32'h414dab98, 32'h40cd21e0, 32'hc2578c8d, 32'h4225f8f2, 32'h42bba5a7, 32'hc2a8fa11, 32'h41d8727b, 32'hc1f6b042};
test_output[9487] = '{32'h42bba5a7};
test_index[9487] = '{4};
test_input[75904:75911] = '{32'h41ffe077, 32'h42476363, 32'h429b2bdc, 32'hc1dd6e5b, 32'h40a7b37b, 32'hc26ad36b, 32'hc215b202, 32'hbfa07a8b};
test_output[9488] = '{32'h429b2bdc};
test_index[9488] = '{2};
test_input[75912:75919] = '{32'h4255ed7f, 32'hc22f1bb1, 32'hc12644d3, 32'h42bdf694, 32'h4218ec15, 32'hc28bd8e2, 32'hc2679d38, 32'hc119721b};
test_output[9489] = '{32'h42bdf694};
test_index[9489] = '{3};
test_input[75920:75927] = '{32'h424ca1fb, 32'h429561eb, 32'hc19e65e3, 32'hc2b23350, 32'hc14a0af5, 32'hc2984391, 32'hc20b7fe7, 32'h423c4e42};
test_output[9490] = '{32'h429561eb};
test_index[9490] = '{1};
test_input[75928:75935] = '{32'h421446af, 32'h40e0a176, 32'hc1ad96a5, 32'hc29deaa1, 32'h4286ec57, 32'h4028debc, 32'hc25702a0, 32'h4193f76c};
test_output[9491] = '{32'h4286ec57};
test_index[9491] = '{4};
test_input[75936:75943] = '{32'hc28d9650, 32'h42865ac0, 32'h42801464, 32'hc125ef11, 32'h42ac9e6a, 32'h4293ee55, 32'h42c1a6fb, 32'hc21f9765};
test_output[9492] = '{32'h42c1a6fb};
test_index[9492] = '{6};
test_input[75944:75951] = '{32'h42bbeeb5, 32'hc2a8b173, 32'h4210f522, 32'h41b71c77, 32'hc281c919, 32'h429b3de6, 32'hc2a5cde3, 32'h41a04a80};
test_output[9493] = '{32'h42bbeeb5};
test_index[9493] = '{0};
test_input[75952:75959] = '{32'hc25dd4a4, 32'hc209efe3, 32'h42c0ea22, 32'h4181d69b, 32'hc2a5b594, 32'h407f87a5, 32'h41d2925e, 32'hc286fef1};
test_output[9494] = '{32'h42c0ea22};
test_index[9494] = '{2};
test_input[75960:75967] = '{32'h42a8472d, 32'h422a178b, 32'hc194857d, 32'hc1d7bab0, 32'h425b93b7, 32'h4189aff6, 32'hc2787c86, 32'hc2ab8b95};
test_output[9495] = '{32'h42a8472d};
test_index[9495] = '{0};
test_input[75968:75975] = '{32'h42a8c8df, 32'hc1d52e68, 32'hc22f92cb, 32'hc1885660, 32'hc2c0ee79, 32'hc1affdf8, 32'h41b686a2, 32'hc2451c42};
test_output[9496] = '{32'h42a8c8df};
test_index[9496] = '{0};
test_input[75976:75983] = '{32'hc18a8d8d, 32'h42835276, 32'h401a3085, 32'h426b2ccd, 32'h40a10ea3, 32'h42b046b8, 32'hc2087d7a, 32'h41e8d054};
test_output[9497] = '{32'h42b046b8};
test_index[9497] = '{5};
test_input[75984:75991] = '{32'hc2674ac6, 32'hc183ea36, 32'hc298b3d1, 32'hc29d556e, 32'hc13696d7, 32'h4212ba71, 32'hc2a4c491, 32'h41319806};
test_output[9498] = '{32'h4212ba71};
test_index[9498] = '{5};
test_input[75992:75999] = '{32'hc2020171, 32'h42928f16, 32'hc24c3f70, 32'h4209db4f, 32'hc2a83902, 32'hc2ab636b, 32'h42734012, 32'hc2a73248};
test_output[9499] = '{32'h42928f16};
test_index[9499] = '{1};
test_input[76000:76007] = '{32'hc1b61467, 32'h42156762, 32'hc2b208ab, 32'hc27b70e4, 32'hc2748b37, 32'h4298506d, 32'hc18a346d, 32'h42992261};
test_output[9500] = '{32'h42992261};
test_index[9500] = '{7};
test_input[76008:76015] = '{32'hc25a02ed, 32'h42a4e127, 32'h42648dee, 32'hc2207fd4, 32'hc2186699, 32'h42c2cffb, 32'hc20d58f3, 32'hc28b47ca};
test_output[9501] = '{32'h42c2cffb};
test_index[9501] = '{5};
test_input[76016:76023] = '{32'h426684f0, 32'h42a39e2f, 32'hc292943c, 32'hc207fb18, 32'hc1e037eb, 32'hc2429370, 32'h42bfddd7, 32'hc2a9bb61};
test_output[9502] = '{32'h42bfddd7};
test_index[9502] = '{6};
test_input[76024:76031] = '{32'h42bc4da4, 32'h42692a9c, 32'hc2c50ec5, 32'h42bd9486, 32'h4074dd71, 32'hc1ffcf0d, 32'hc02da75f, 32'hc2a69b38};
test_output[9503] = '{32'h42bd9486};
test_index[9503] = '{3};
test_input[76032:76039] = '{32'h41f6ca8b, 32'h4262e646, 32'h4261e924, 32'h420216f2, 32'h428c3857, 32'h428e2083, 32'h42879e15, 32'h3fc8d23f};
test_output[9504] = '{32'h428e2083};
test_index[9504] = '{5};
test_input[76040:76047] = '{32'hc2b9089b, 32'h422d5c2d, 32'h42b67335, 32'h41af8dbd, 32'hc26dd39c, 32'hc1dda845, 32'h42bfa2a4, 32'h419c3e3d};
test_output[9505] = '{32'h42bfa2a4};
test_index[9505] = '{6};
test_input[76048:76055] = '{32'hc207af3f, 32'hc2c165bc, 32'hc28edf99, 32'h421df116, 32'hc0d76b25, 32'h42a5c56f, 32'h422c790a, 32'h4103444b};
test_output[9506] = '{32'h42a5c56f};
test_index[9506] = '{5};
test_input[76056:76063] = '{32'h4236430e, 32'h4280ca78, 32'hc0187d7b, 32'h3f161220, 32'hc2918786, 32'hc293d9f8, 32'hc2480641, 32'hc1ec9740};
test_output[9507] = '{32'h4280ca78};
test_index[9507] = '{1};
test_input[76064:76071] = '{32'hc19c8751, 32'h4253103f, 32'h41d1b596, 32'hc221cace, 32'hc1fb0333, 32'hc278a088, 32'hc1af5e81, 32'hc28f9f52};
test_output[9508] = '{32'h4253103f};
test_index[9508] = '{1};
test_input[76072:76079] = '{32'h424161dc, 32'h41e943c4, 32'hc2205aae, 32'h422264f9, 32'hc181f505, 32'h42a02c4a, 32'h422aa2b3, 32'hc23a1ff6};
test_output[9509] = '{32'h42a02c4a};
test_index[9509] = '{5};
test_input[76080:76087] = '{32'hc2346f4c, 32'hc294b585, 32'h42976b4a, 32'h41d8c272, 32'hc288d13f, 32'h42bcbe81, 32'h40a389e7, 32'hc238eead};
test_output[9510] = '{32'h42bcbe81};
test_index[9510] = '{5};
test_input[76088:76095] = '{32'hc1c0e823, 32'hc2a8b9d6, 32'hc2b175e3, 32'hc25c6eaa, 32'hc13e8070, 32'h429b1cab, 32'hc2772f88, 32'hc1c3683a};
test_output[9511] = '{32'h429b1cab};
test_index[9511] = '{5};
test_input[76096:76103] = '{32'hc2514987, 32'h402e12da, 32'hc23b00fd, 32'h40d94047, 32'h4256828d, 32'hc104158a, 32'h42688caf, 32'hc26385b0};
test_output[9512] = '{32'h42688caf};
test_index[9512] = '{6};
test_input[76104:76111] = '{32'hc252fb62, 32'h42919291, 32'hc2095d3a, 32'hc1fb30a5, 32'h411d8e37, 32'h4280cf69, 32'hc2bf40f1, 32'h429f074b};
test_output[9513] = '{32'h429f074b};
test_index[9513] = '{7};
test_input[76112:76119] = '{32'h42bf4be0, 32'hc212bdad, 32'hc29237f2, 32'hc20e8bed, 32'h42302781, 32'hc1e0c7f3, 32'h4269acb6, 32'h42bf0ecb};
test_output[9514] = '{32'h42bf4be0};
test_index[9514] = '{0};
test_input[76120:76127] = '{32'h416ea674, 32'h41f43952, 32'h40c0bd44, 32'h42b5711a, 32'h411dec06, 32'hc1ecc7aa, 32'h425b24b9, 32'hc20e174c};
test_output[9515] = '{32'h42b5711a};
test_index[9515] = '{3};
test_input[76128:76135] = '{32'hc2756517, 32'hc1c3febf, 32'h4289deca, 32'h42a935ab, 32'h40079c09, 32'h42950f9f, 32'hc0001e4c, 32'hc1e92794};
test_output[9516] = '{32'h42a935ab};
test_index[9516] = '{3};
test_input[76136:76143] = '{32'h41421afe, 32'h4120b713, 32'h4291fdb8, 32'h4263599a, 32'h40bbedbd, 32'h42c3960c, 32'hc1d9d209, 32'hc214b796};
test_output[9517] = '{32'h42c3960c};
test_index[9517] = '{5};
test_input[76144:76151] = '{32'hc2924402, 32'h419d379c, 32'hc2a5fee3, 32'hc20b4755, 32'h429af0b5, 32'hc0afc1d6, 32'h42849ed3, 32'hc13e81b1};
test_output[9518] = '{32'h429af0b5};
test_index[9518] = '{4};
test_input[76152:76159] = '{32'hc1b881f8, 32'h4279ea75, 32'h41998d7f, 32'hc2b2da4c, 32'h42a89935, 32'h42a15c16, 32'h419ca914, 32'hc1a7a3f6};
test_output[9519] = '{32'h42a89935};
test_index[9519] = '{4};
test_input[76160:76167] = '{32'hc15937ef, 32'hc220d095, 32'h428790e6, 32'h4165e92c, 32'hc2a96e8c, 32'h42b95dca, 32'h41c8c72e, 32'hc2627ea8};
test_output[9520] = '{32'h42b95dca};
test_index[9520] = '{5};
test_input[76168:76175] = '{32'h41f2255f, 32'h4223ead6, 32'hc2a35f55, 32'hc26dbba1, 32'h42632b8b, 32'hc2a7094f, 32'h424b9a1b, 32'h4241fbbe};
test_output[9521] = '{32'h42632b8b};
test_index[9521] = '{4};
test_input[76176:76183] = '{32'h42402e8d, 32'hc22dd7cc, 32'h42a0defe, 32'hc16c977b, 32'hc21ada62, 32'h425acdee, 32'hc1d2d154, 32'hc29ce122};
test_output[9522] = '{32'h42a0defe};
test_index[9522] = '{2};
test_input[76184:76191] = '{32'hc18bced8, 32'h429c90ab, 32'h42a5512e, 32'h42595b7a, 32'hc23b4446, 32'hc2aba687, 32'hbfdc157e, 32'hc2761bf7};
test_output[9523] = '{32'h42a5512e};
test_index[9523] = '{2};
test_input[76192:76199] = '{32'hc296d4b0, 32'hc2bac42f, 32'hc19f1e98, 32'hc1ec73cd, 32'h42beefa1, 32'h41b11a1c, 32'h425e1390, 32'h423c00fe};
test_output[9524] = '{32'h42beefa1};
test_index[9524] = '{4};
test_input[76200:76207] = '{32'h41dbb005, 32'hc20610bc, 32'hc1cd4da7, 32'hc2176ce8, 32'hc0b6b0d9, 32'h429a6e0c, 32'h414e1504, 32'hc2ac033d};
test_output[9525] = '{32'h429a6e0c};
test_index[9525] = '{5};
test_input[76208:76215] = '{32'hc2bf92d7, 32'h420dbcbd, 32'h417fdb1c, 32'h41f2084b, 32'hc17df3eb, 32'hc14e37f9, 32'h427a12a5, 32'hc28cd075};
test_output[9526] = '{32'h427a12a5};
test_index[9526] = '{6};
test_input[76216:76223] = '{32'hc2b0e4d6, 32'h41896274, 32'hc095760b, 32'hc287c825, 32'h40b06555, 32'hc28a6413, 32'h42978920, 32'h405dadd2};
test_output[9527] = '{32'h42978920};
test_index[9527] = '{6};
test_input[76224:76231] = '{32'hc11d6fc8, 32'hc20de69f, 32'hc25a713b, 32'hc2267580, 32'hc1d16a5d, 32'h41e1aa26, 32'hc1f65e6c, 32'hc28806e7};
test_output[9528] = '{32'h41e1aa26};
test_index[9528] = '{5};
test_input[76232:76239] = '{32'hc18387d4, 32'hc0687e3b, 32'h428ba8e0, 32'h424c2228, 32'h41ef118b, 32'h4238b4f7, 32'hc0a84275, 32'hc286105d};
test_output[9529] = '{32'h428ba8e0};
test_index[9529] = '{2};
test_input[76240:76247] = '{32'h42b3cccf, 32'hbfa467d2, 32'h413919de, 32'h41071e0e, 32'h42279e17, 32'hc27f71af, 32'h410a297d, 32'h41dac639};
test_output[9530] = '{32'h42b3cccf};
test_index[9530] = '{0};
test_input[76248:76255] = '{32'hc2651b69, 32'hc29b1857, 32'hc1f97775, 32'h42bf5ad8, 32'hc1fce7a2, 32'h42c5c615, 32'hc28c9174, 32'hc193d09d};
test_output[9531] = '{32'h42c5c615};
test_index[9531] = '{5};
test_input[76256:76263] = '{32'h429e3370, 32'h423a8de7, 32'h4256dd97, 32'hc24a09c7, 32'h41b8ad5d, 32'h41ec9572, 32'hc2acf4ce, 32'hc13d0dde};
test_output[9532] = '{32'h429e3370};
test_index[9532] = '{0};
test_input[76264:76271] = '{32'hc2a0e668, 32'hc261406c, 32'hc1b13577, 32'hc28fb7e9, 32'h421a58c1, 32'h42bdbf0e, 32'hc297651e, 32'h42536656};
test_output[9533] = '{32'h42bdbf0e};
test_index[9533] = '{5};
test_input[76272:76279] = '{32'h42ba7e69, 32'h41f39145, 32'hc21d2395, 32'h4292d79c, 32'h42b9d582, 32'h42660235, 32'h40b9035a, 32'hc108eb90};
test_output[9534] = '{32'h42ba7e69};
test_index[9534] = '{0};
test_input[76280:76287] = '{32'hc19e2617, 32'h42a337e8, 32'h40e4d246, 32'h414d448b, 32'h425880f7, 32'h42688f21, 32'hc286c97d, 32'h4296f64d};
test_output[9535] = '{32'h42a337e8};
test_index[9535] = '{1};
test_input[76288:76295] = '{32'h40d1e2da, 32'hc235d986, 32'hc16a58b1, 32'hc112ac58, 32'h42bb6561, 32'hc125d6d4, 32'h42c20e3b, 32'hc1d0ba41};
test_output[9536] = '{32'h42c20e3b};
test_index[9536] = '{6};
test_input[76296:76303] = '{32'h42a03177, 32'h42a6c35a, 32'hc29b1b8d, 32'h4122fd87, 32'hc263d9a3, 32'h425722d8, 32'hc17f0f0c, 32'h422961e1};
test_output[9537] = '{32'h42a6c35a};
test_index[9537] = '{1};
test_input[76304:76311] = '{32'h4289156f, 32'h4271e916, 32'h42721861, 32'h40814b24, 32'hc2be5875, 32'hc23e68b1, 32'h4285ec5f, 32'h42ae1461};
test_output[9538] = '{32'h42ae1461};
test_index[9538] = '{7};
test_input[76312:76319] = '{32'h42afbace, 32'hc28bf23f, 32'hc2b44239, 32'h42a6e0f1, 32'hc11ec7a3, 32'h410f8801, 32'hc2b9c500, 32'hc1d239eb};
test_output[9539] = '{32'h42afbace};
test_index[9539] = '{0};
test_input[76320:76327] = '{32'hc154b642, 32'hc2612b3d, 32'hc118ce0b, 32'hc2968114, 32'h42056ecd, 32'hbfa43298, 32'h41c98700, 32'hc114fc06};
test_output[9540] = '{32'h42056ecd};
test_index[9540] = '{4};
test_input[76328:76335] = '{32'h4212e1eb, 32'hc28197e6, 32'hc23dc92a, 32'h42c6e2b0, 32'hc09f90ef, 32'h410544c4, 32'h42b7d60a, 32'h4082fb99};
test_output[9541] = '{32'h42c6e2b0};
test_index[9541] = '{3};
test_input[76336:76343] = '{32'hc2355218, 32'h42125db2, 32'hc2a3655b, 32'hbe45df50, 32'hc202cdc8, 32'hc2c4644e, 32'h41fe88bd, 32'h41a73143};
test_output[9542] = '{32'h42125db2};
test_index[9542] = '{1};
test_input[76344:76351] = '{32'h426f9e13, 32'hc1be8a12, 32'hc1d5aa6e, 32'h423de140, 32'h42b07286, 32'h412b0d52, 32'h41035d14, 32'hc2421d65};
test_output[9543] = '{32'h42b07286};
test_index[9543] = '{4};
test_input[76352:76359] = '{32'hc1bf0989, 32'h425361be, 32'hc1899304, 32'h420668d4, 32'hc0fceaec, 32'hc2a6eb69, 32'h423a4c47, 32'h423b7454};
test_output[9544] = '{32'h425361be};
test_index[9544] = '{1};
test_input[76360:76367] = '{32'h42ad67a3, 32'hc25f35c7, 32'hc26f242d, 32'h429db3f4, 32'h4249498a, 32'hc250b1c9, 32'hc1f9ca82, 32'h41f3dddd};
test_output[9545] = '{32'h42ad67a3};
test_index[9545] = '{0};
test_input[76368:76375] = '{32'h41be70f3, 32'hc2c22a8a, 32'h42893195, 32'h41db29ad, 32'hc2ba7d1d, 32'h42b1f88e, 32'hc2459634, 32'h41a0576f};
test_output[9546] = '{32'h42b1f88e};
test_index[9546] = '{5};
test_input[76376:76383] = '{32'h42755518, 32'h413ceac6, 32'hc277147d, 32'h41b4913a, 32'hc2c47ac8, 32'h41bc9c01, 32'hc2421ee7, 32'h41c805ce};
test_output[9547] = '{32'h42755518};
test_index[9547] = '{0};
test_input[76384:76391] = '{32'hc2799338, 32'h42adc12c, 32'h42556f6f, 32'h41121f28, 32'hc2a86104, 32'h40eb2624, 32'hc25f8303, 32'h42bb85e2};
test_output[9548] = '{32'h42bb85e2};
test_index[9548] = '{7};
test_input[76392:76399] = '{32'hc0ed9d07, 32'h421282a0, 32'h41d3fa94, 32'h42b82a92, 32'h41c1abf7, 32'hc1d0a9c5, 32'hc1c751c0, 32'hc2b65846};
test_output[9549] = '{32'h42b82a92};
test_index[9549] = '{3};
test_input[76400:76407] = '{32'h4214c53b, 32'hc26940f0, 32'hc1595e1a, 32'hc2624dd6, 32'hc2c57b7d, 32'hc262145f, 32'hc1c2b52a, 32'h41fc5da4};
test_output[9550] = '{32'h4214c53b};
test_index[9550] = '{0};
test_input[76408:76415] = '{32'hc26ca6d3, 32'hc2895cfd, 32'hc18ea447, 32'hc233ad16, 32'h419e1105, 32'h41a4180b, 32'hc25fb526, 32'h411ee6b0};
test_output[9551] = '{32'h41a4180b};
test_index[9551] = '{5};
test_input[76416:76423] = '{32'hc2bedabe, 32'hc2a18e6d, 32'h426b2322, 32'h41ad6c85, 32'hc1954381, 32'hc2a7a8ad, 32'h42b4fb64, 32'hc1bd0a15};
test_output[9552] = '{32'h42b4fb64};
test_index[9552] = '{6};
test_input[76424:76431] = '{32'h428e104f, 32'hc2662744, 32'hc2a839c4, 32'h424b0abe, 32'h428ab6d4, 32'h42b03382, 32'hc292aad4, 32'hc231eb1e};
test_output[9553] = '{32'h42b03382};
test_index[9553] = '{5};
test_input[76432:76439] = '{32'hc2be8c6c, 32'h40d86ad3, 32'h42807bd3, 32'hbf09d271, 32'hc2a3a912, 32'hc2104e66, 32'h418dd1b6, 32'h4180ce25};
test_output[9554] = '{32'h42807bd3};
test_index[9554] = '{2};
test_input[76440:76447] = '{32'hc24796f8, 32'hc18f41b0, 32'h429e5e82, 32'hc2116873, 32'hc2aca389, 32'hc2b8c5d1, 32'h4263f915, 32'h42bd0441};
test_output[9555] = '{32'h42bd0441};
test_index[9555] = '{7};
test_input[76448:76455] = '{32'h40dce079, 32'hc2b87bba, 32'h4296fc47, 32'h42ac64e0, 32'hbe76e62a, 32'h42bf9eb4, 32'hc2bb248a, 32'hc231e6a0};
test_output[9556] = '{32'h42bf9eb4};
test_index[9556] = '{5};
test_input[76456:76463] = '{32'hc27a716a, 32'h429b2b5d, 32'h42821940, 32'h41b635fd, 32'h411ebcda, 32'hc1c932ab, 32'h3fe86ea7, 32'hc2b25807};
test_output[9557] = '{32'h429b2b5d};
test_index[9557] = '{1};
test_input[76464:76471] = '{32'h4255f4de, 32'hc29b17c1, 32'h4252c066, 32'hc29dd548, 32'h42a534e8, 32'hc2aba574, 32'h4235527e, 32'hc2888961};
test_output[9558] = '{32'h42a534e8};
test_index[9558] = '{4};
test_input[76472:76479] = '{32'h428f9f70, 32'h428276fb, 32'h4184a029, 32'hc294d2a4, 32'h423e7d4d, 32'hc2c47f8c, 32'hc23bf82a, 32'hc2c4f52a};
test_output[9559] = '{32'h428f9f70};
test_index[9559] = '{0};
test_input[76480:76487] = '{32'hc201122e, 32'h42a6bd77, 32'hc071fe29, 32'hc27c4b7c, 32'hc2ad3269, 32'hc23dfcea, 32'hc2ab97ca, 32'h422858ca};
test_output[9560] = '{32'h42a6bd77};
test_index[9560] = '{1};
test_input[76488:76495] = '{32'h4294a0d6, 32'h41c9517f, 32'h427095a7, 32'h4115f0e8, 32'hc28274df, 32'hc2a08429, 32'h41e02179, 32'hc25f3db3};
test_output[9561] = '{32'h4294a0d6};
test_index[9561] = '{0};
test_input[76496:76503] = '{32'h418d178f, 32'h42ac7da0, 32'hc2045680, 32'hc2c1ff77, 32'hc201c7c2, 32'h414c60b3, 32'hc21926cf, 32'hc1405ffd};
test_output[9562] = '{32'h42ac7da0};
test_index[9562] = '{1};
test_input[76504:76511] = '{32'hc295cf78, 32'h42155732, 32'hc125cfc0, 32'h4214845c, 32'h428406e0, 32'h42463cda, 32'h41850e4e, 32'h3fe9688c};
test_output[9563] = '{32'h428406e0};
test_index[9563] = '{4};
test_input[76512:76519] = '{32'hc1ec15ef, 32'hc2063749, 32'h42a7cfdc, 32'hc1503dbd, 32'h41e6f9f6, 32'hc2a01b21, 32'hc2193d65, 32'h4185dc50};
test_output[9564] = '{32'h42a7cfdc};
test_index[9564] = '{2};
test_input[76520:76527] = '{32'h41f8f3da, 32'h4283d0f2, 32'h41c89f2a, 32'hc26ebd62, 32'h42438c2f, 32'hc2aa65d7, 32'hc230f568, 32'h41d032b5};
test_output[9565] = '{32'h4283d0f2};
test_index[9565] = '{1};
test_input[76528:76535] = '{32'h41a7b9d2, 32'hc259ead8, 32'hc2ac24e8, 32'hbfd0d4a4, 32'hc25172d4, 32'hc247df37, 32'hc2924b1b, 32'h42b3e85b};
test_output[9566] = '{32'h42b3e85b};
test_index[9566] = '{7};
test_input[76536:76543] = '{32'hc28f8f52, 32'h41b6c3fb, 32'h40ca65f5, 32'h4261995d, 32'h418d1ef7, 32'hc23d484c, 32'hc1c0d8af, 32'hc123b79c};
test_output[9567] = '{32'h4261995d};
test_index[9567] = '{3};
test_input[76544:76551] = '{32'hc29e3b06, 32'h42259a65, 32'h41a18755, 32'h4186fe34, 32'hc084f790, 32'h418cbb92, 32'h428d917d, 32'hc0ddf88b};
test_output[9568] = '{32'h428d917d};
test_index[9568] = '{6};
test_input[76552:76559] = '{32'h42425c65, 32'hc274cbb5, 32'hc0b12c71, 32'h40dbc555, 32'h418d1dd8, 32'hc2994726, 32'hc26f99c0, 32'h40c83187};
test_output[9569] = '{32'h42425c65};
test_index[9569] = '{0};
test_input[76560:76567] = '{32'hc1af47c0, 32'h426eded5, 32'h41cd7f71, 32'h41c7bfa6, 32'h41e3ab6c, 32'hc2bc8787, 32'hc23fd895, 32'h427b1713};
test_output[9570] = '{32'h427b1713};
test_index[9570] = '{7};
test_input[76568:76575] = '{32'h42070b53, 32'hc2a0d7cb, 32'hc1b72440, 32'h42586862, 32'hc278ff0b, 32'hc24fdcab, 32'hc2b6fd04, 32'h40c0cdc3};
test_output[9571] = '{32'h42586862};
test_index[9571] = '{3};
test_input[76576:76583] = '{32'h42b1566d, 32'hc286f9fd, 32'h40a70177, 32'h4240715b, 32'h41091ac0, 32'hc1cb1406, 32'hc23ab43d, 32'h4257f7c6};
test_output[9572] = '{32'h42b1566d};
test_index[9572] = '{0};
test_input[76584:76591] = '{32'h42a64be0, 32'h4109ca8e, 32'h42834af0, 32'hc253de51, 32'hc2b0feef, 32'h428d033c, 32'hc29db3f6, 32'h419c4e8f};
test_output[9573] = '{32'h42a64be0};
test_index[9573] = '{0};
test_input[76592:76599] = '{32'h42908049, 32'h423f9166, 32'hc169df45, 32'hc26454d6, 32'hc25e5762, 32'hc2ac7297, 32'hc2bc1e57, 32'hc2b9351a};
test_output[9574] = '{32'h42908049};
test_index[9574] = '{0};
test_input[76600:76607] = '{32'h42b51ac8, 32'h3f36b298, 32'hc186cd35, 32'h4247439f, 32'h41438980, 32'hc154f8ea, 32'h428afe8a, 32'hc292ef58};
test_output[9575] = '{32'h42b51ac8};
test_index[9575] = '{0};
test_input[76608:76615] = '{32'h429da378, 32'h4257b83e, 32'hc28eec1b, 32'h419f8c72, 32'h429b2d94, 32'h4264658d, 32'hc291abda, 32'hc2c16da5};
test_output[9576] = '{32'h429da378};
test_index[9576] = '{0};
test_input[76616:76623] = '{32'h42a0a6e5, 32'h4203c386, 32'hc0c5a8b1, 32'h41f1dcbf, 32'h42a113e5, 32'hc2c1dcda, 32'h42b1233e, 32'h42b978e0};
test_output[9577] = '{32'h42b978e0};
test_index[9577] = '{7};
test_input[76624:76631] = '{32'h422c82e2, 32'h413f1fca, 32'h42318da6, 32'hc20cbcaf, 32'hc22b3d64, 32'h421b4c1d, 32'h425c8064, 32'hc2401db9};
test_output[9578] = '{32'h425c8064};
test_index[9578] = '{6};
test_input[76632:76639] = '{32'hc1963bd0, 32'h42902e85, 32'hc29e8fea, 32'h4096aaca, 32'h41961db4, 32'hc20d09fe, 32'hc291fb9e, 32'h42054da7};
test_output[9579] = '{32'h42902e85};
test_index[9579] = '{1};
test_input[76640:76647] = '{32'hc28183eb, 32'hc2bc72d4, 32'hc2b45608, 32'hc163e57a, 32'h41234fe7, 32'hc284c11a, 32'hc1b35957, 32'h42015948};
test_output[9580] = '{32'h42015948};
test_index[9580] = '{7};
test_input[76648:76655] = '{32'h423813a2, 32'h42941654, 32'hc263806b, 32'hc200ed9f, 32'h4289f777, 32'h422e479f, 32'hc1fd7eb3, 32'hc2993008};
test_output[9581] = '{32'h42941654};
test_index[9581] = '{1};
test_input[76656:76663] = '{32'h423d467a, 32'h41b5b853, 32'h41f4ad18, 32'hbf97fd76, 32'hc2a4225c, 32'hc1e31446, 32'h4282719f, 32'h42c7f2ac};
test_output[9582] = '{32'h42c7f2ac};
test_index[9582] = '{7};
test_input[76664:76671] = '{32'hc25f15d4, 32'h4295287e, 32'hc22906e2, 32'hc284cd3c, 32'hc1f55920, 32'h42b7799a, 32'h42c71842, 32'h4237679a};
test_output[9583] = '{32'h42c71842};
test_index[9583] = '{6};
test_input[76672:76679] = '{32'h41d4a474, 32'h42a7de16, 32'h429c2b7b, 32'hc27704df, 32'hc01e4f18, 32'h41162685, 32'h422d2082, 32'hc2c1a569};
test_output[9584] = '{32'h42a7de16};
test_index[9584] = '{1};
test_input[76680:76687] = '{32'hc293b56b, 32'hc23c6cb5, 32'h42af2d2e, 32'hc2375ff1, 32'hc2abe56d, 32'hc2b4356a, 32'h422dbe27, 32'h427ac2ba};
test_output[9585] = '{32'h42af2d2e};
test_index[9585] = '{2};
test_input[76688:76695] = '{32'h42c263c8, 32'h42b286f6, 32'hc244d71d, 32'h4229222c, 32'hc2c09b49, 32'hc2aace6a, 32'hc224be85, 32'h42c2c517};
test_output[9586] = '{32'h42c2c517};
test_index[9586] = '{7};
test_input[76696:76703] = '{32'h40e1d8d4, 32'hc00e400b, 32'h42a76bba, 32'hc205d049, 32'hc2573f98, 32'h41e9cc18, 32'hc178edd6, 32'h3f54001f};
test_output[9587] = '{32'h42a76bba};
test_index[9587] = '{2};
test_input[76704:76711] = '{32'h41c4c031, 32'hc2c2d378, 32'h4233490d, 32'hc2bbe28f, 32'hc259d06f, 32'hc278ee8b, 32'hc288706a, 32'h42559095};
test_output[9588] = '{32'h42559095};
test_index[9588] = '{7};
test_input[76712:76719] = '{32'h429a3871, 32'hc2811dc4, 32'hc13ad3c5, 32'hc2699c94, 32'hc286120b, 32'hc081c4eb, 32'h41a1c1c2, 32'h429301e3};
test_output[9589] = '{32'h429a3871};
test_index[9589] = '{0};
test_input[76720:76727] = '{32'hc1df62dc, 32'hbf436460, 32'hc27d3241, 32'h42b5f106, 32'hc192e1e3, 32'hc1c99e95, 32'h4054fd3e, 32'h41925e54};
test_output[9590] = '{32'h42b5f106};
test_index[9590] = '{3};
test_input[76728:76735] = '{32'hc19adc1c, 32'hc29b26f5, 32'h41f4f3ec, 32'hc2903a6f, 32'h419212a8, 32'hc21554dc, 32'h420dc071, 32'h42a78e90};
test_output[9591] = '{32'h42a78e90};
test_index[9591] = '{7};
test_input[76736:76743] = '{32'hc2c2cc09, 32'hc212e714, 32'hc1ebecad, 32'h42a4423a, 32'hc2bfc6f0, 32'h42843334, 32'hc2c0fc37, 32'h4258bb65};
test_output[9592] = '{32'h42a4423a};
test_index[9592] = '{3};
test_input[76744:76751] = '{32'h42c65bd0, 32'hc291d93b, 32'h42ae08bb, 32'hc2506e29, 32'hc2ab1bec, 32'hc25ef85e, 32'h42a9c7f1, 32'h423501bb};
test_output[9593] = '{32'h42c65bd0};
test_index[9593] = '{0};
test_input[76752:76759] = '{32'hc259a5d6, 32'hc29dcdd1, 32'hc0b3dccc, 32'hc2573dae, 32'h42a23572, 32'h41e0807e, 32'h40cf0d8c, 32'hc204b26d};
test_output[9594] = '{32'h42a23572};
test_index[9594] = '{4};
test_input[76760:76767] = '{32'hc2882b84, 32'hc2ab5788, 32'h42bdcd0f, 32'hc2137567, 32'hc25070a8, 32'hc1caba8f, 32'hc273956b, 32'h42b9a309};
test_output[9595] = '{32'h42bdcd0f};
test_index[9595] = '{2};
test_input[76768:76775] = '{32'h415942b7, 32'h42b00b23, 32'h40d78547, 32'h41652f01, 32'h42976de1, 32'hc2be6c23, 32'hbfd49f39, 32'h42c284bd};
test_output[9596] = '{32'h42c284bd};
test_index[9596] = '{7};
test_input[76776:76783] = '{32'h4202bfcd, 32'h416b14d9, 32'hc26b2c3d, 32'h4263c00d, 32'h42aab8eb, 32'hc1fd270d, 32'hc292fde6, 32'hc235849c};
test_output[9597] = '{32'h42aab8eb};
test_index[9597] = '{4};
test_input[76784:76791] = '{32'hc281d015, 32'h42ae725f, 32'h42289a87, 32'h41f9316d, 32'hc12f60eb, 32'hc2c0640c, 32'h41f2d969, 32'h4186eb1a};
test_output[9598] = '{32'h42ae725f};
test_index[9598] = '{1};
test_input[76792:76799] = '{32'h4282f4f4, 32'hbe2e387e, 32'h4264cd27, 32'hc2344bfa, 32'hc2b0b1df, 32'hc2429c2e, 32'hc283a272, 32'hc28d9464};
test_output[9599] = '{32'h4282f4f4};
test_index[9599] = '{0};
test_input[76800:76807] = '{32'h429a5f84, 32'h3c09a68f, 32'h42c0c1a0, 32'hc0cb377e, 32'h418b4209, 32'h42784a8a, 32'hc26e1bbf, 32'hc213d76f};
test_output[9600] = '{32'h42c0c1a0};
test_index[9600] = '{2};
test_input[76808:76815] = '{32'h412d27dc, 32'h421f46f5, 32'hc252d1ee, 32'h4249867b, 32'hc16a229e, 32'hc13d4ba1, 32'hc173ac64, 32'h40d94b2d};
test_output[9601] = '{32'h4249867b};
test_index[9601] = '{3};
test_input[76816:76823] = '{32'hc2ad3c20, 32'h429dc7cf, 32'h401b8287, 32'h42080fd6, 32'hc19087e3, 32'hc28ce945, 32'h3ef54932, 32'h40edf486};
test_output[9602] = '{32'h429dc7cf};
test_index[9602] = '{1};
test_input[76824:76831] = '{32'hc2a5f4e3, 32'hc2bceb2b, 32'hc05b093a, 32'h42b9522b, 32'hc2572921, 32'h421c9a05, 32'h42ad1ad2, 32'hc1ff841a};
test_output[9603] = '{32'h42b9522b};
test_index[9603] = '{3};
test_input[76832:76839] = '{32'hc2c364e8, 32'h4113b3ff, 32'hc2b704ef, 32'hc29f233f, 32'hc2a23542, 32'hc2b831fd, 32'h41bd79ff, 32'h420420c6};
test_output[9604] = '{32'h420420c6};
test_index[9604] = '{7};
test_input[76840:76847] = '{32'h3fa53e00, 32'h42b2d527, 32'hc1ca5f76, 32'hc26a2862, 32'h420cd910, 32'hc2baa7fc, 32'h408e9aec, 32'hc2bc31d1};
test_output[9605] = '{32'h42b2d527};
test_index[9605] = '{1};
test_input[76848:76855] = '{32'hc29b2966, 32'h42c43d02, 32'h413b8838, 32'hc2be1b36, 32'hc1ea73a0, 32'h42ad2dfd, 32'h41ed0a99, 32'hc2725da0};
test_output[9606] = '{32'h42c43d02};
test_index[9606] = '{1};
test_input[76856:76863] = '{32'hc2254656, 32'h42587be6, 32'h42b90d8f, 32'hc216915e, 32'h40a30711, 32'hc2a5cfbe, 32'h4275cc24, 32'h412d109e};
test_output[9607] = '{32'h42b90d8f};
test_index[9607] = '{2};
test_input[76864:76871] = '{32'hc2745dcc, 32'h428b550d, 32'h42c35832, 32'h4220822d, 32'h42a5867f, 32'h42503bc8, 32'h41466f8d, 32'hc2302e62};
test_output[9608] = '{32'h42c35832};
test_index[9608] = '{2};
test_input[76872:76879] = '{32'hc25601eb, 32'hc1332683, 32'hc0e60258, 32'h42b5d298, 32'hc0ace354, 32'h4190b053, 32'h426fbe35, 32'hc1ec52ce};
test_output[9609] = '{32'h42b5d298};
test_index[9609] = '{3};
test_input[76880:76887] = '{32'hc00862f8, 32'hc28b1b5d, 32'h4196cb4d, 32'hc1fa6e3f, 32'h422019fe, 32'hc298f588, 32'h425f45e4, 32'hc2008bf9};
test_output[9610] = '{32'h425f45e4};
test_index[9610] = '{6};
test_input[76888:76895] = '{32'h4086b045, 32'hc2144c68, 32'hc1bf8284, 32'hc1822345, 32'hc1e5925c, 32'hc12e210c, 32'h42711230, 32'h424d6796};
test_output[9611] = '{32'h42711230};
test_index[9611] = '{6};
test_input[76896:76903] = '{32'hc21f4b5f, 32'h41ee47c6, 32'h40b6957f, 32'h41993a92, 32'h4215c6ed, 32'h42b7b96e, 32'hc1884866, 32'hc2010443};
test_output[9612] = '{32'h42b7b96e};
test_index[9612] = '{5};
test_input[76904:76911] = '{32'hc2bcd7f8, 32'hc26fb9e1, 32'h425cb037, 32'hc165000f, 32'h42810207, 32'hc1ef41d3, 32'h42c15339, 32'h4260919d};
test_output[9613] = '{32'h42c15339};
test_index[9613] = '{6};
test_input[76912:76919] = '{32'hc2769d33, 32'h425f8411, 32'h426e88e4, 32'hc29fa776, 32'hc21856c4, 32'hc2909e96, 32'h42a4ac62, 32'h429a89a8};
test_output[9614] = '{32'h42a4ac62};
test_index[9614] = '{6};
test_input[76920:76927] = '{32'hc1a78232, 32'h429ee693, 32'h41f3b445, 32'h4269d826, 32'hc0be8c6e, 32'hbf9c26d5, 32'hc28bf09a, 32'h4267f7c6};
test_output[9615] = '{32'h429ee693};
test_index[9615] = '{1};
test_input[76928:76935] = '{32'hc29112d0, 32'hc2a4a4e1, 32'hc0fc23a9, 32'h4291aa44, 32'h42bba044, 32'h4216cba4, 32'h4153d4a9, 32'hc29c154a};
test_output[9616] = '{32'h42bba044};
test_index[9616] = '{4};
test_input[76936:76943] = '{32'h426a571c, 32'h42405c2d, 32'h41bf28c3, 32'h41a955c1, 32'h421ff0cc, 32'h42685106, 32'hc203b900, 32'h42231ca8};
test_output[9617] = '{32'h426a571c};
test_index[9617] = '{0};
test_input[76944:76951] = '{32'h411738d2, 32'hc0841e23, 32'h42a29ace, 32'hc125873c, 32'hc19005ab, 32'h41bc6fe3, 32'h4112499f, 32'hc2934ba9};
test_output[9618] = '{32'h42a29ace};
test_index[9618] = '{2};
test_input[76952:76959] = '{32'hc178156d, 32'hc222f4e9, 32'hc25bc5ba, 32'hc2bd6fce, 32'hc170ea37, 32'h4131707d, 32'h42890da3, 32'hc2130396};
test_output[9619] = '{32'h42890da3};
test_index[9619] = '{6};
test_input[76960:76967] = '{32'hc261a93e, 32'hc28bc8d2, 32'h3f6057e2, 32'h416e791a, 32'hc2ace9ca, 32'h427e6237, 32'h425e1cc8, 32'hc1e1354d};
test_output[9620] = '{32'h427e6237};
test_index[9620] = '{5};
test_input[76968:76975] = '{32'h42a43404, 32'hc1986111, 32'h42acf6a1, 32'h424dbb6e, 32'h42af3611, 32'h421e206b, 32'hc24af142, 32'hc286f926};
test_output[9621] = '{32'h42af3611};
test_index[9621] = '{4};
test_input[76976:76983] = '{32'hc2b3aa11, 32'h416fba45, 32'h423b63bd, 32'h422a9881, 32'hc1db45c2, 32'hc0ca059c, 32'h41ce258b, 32'hc2728346};
test_output[9622] = '{32'h423b63bd};
test_index[9622] = '{2};
test_input[76984:76991] = '{32'h42099f3f, 32'hc1f96a30, 32'hc26f11cb, 32'hc2a3d9c0, 32'h423c9360, 32'h42678829, 32'h42bf2719, 32'hc24aace0};
test_output[9623] = '{32'h42bf2719};
test_index[9623] = '{6};
test_input[76992:76999] = '{32'hc29a82e2, 32'h41908f74, 32'hc1bfa3eb, 32'hc2ac68c4, 32'h42bbf039, 32'hc1044e27, 32'hc2997b96, 32'hc2396f3f};
test_output[9624] = '{32'h42bbf039};
test_index[9624] = '{4};
test_input[77000:77007] = '{32'h42a0d14f, 32'h42b33f39, 32'h42407d0d, 32'h4258ed0c, 32'h42967913, 32'hc27b242a, 32'hc2733ca5, 32'hc04a2b21};
test_output[9625] = '{32'h42b33f39};
test_index[9625] = '{1};
test_input[77008:77015] = '{32'hc21f0182, 32'hc1153fac, 32'h42c65c1f, 32'hc2310c9d, 32'h423d3bba, 32'hc2ba9e15, 32'hc281b6c2, 32'hc19a8a3f};
test_output[9626] = '{32'h42c65c1f};
test_index[9626] = '{2};
test_input[77016:77023] = '{32'hc251186d, 32'hc2a594ee, 32'hc170a83d, 32'hc164c2b8, 32'hc2a11265, 32'hc2a42673, 32'hc203efe0, 32'hc143423c};
test_output[9627] = '{32'hc143423c};
test_index[9627] = '{7};
test_input[77024:77031] = '{32'h4240cafa, 32'hc25b358e, 32'hc28af0f6, 32'h41d24205, 32'hc2b23c5a, 32'h42a3f2b9, 32'hc149eb08, 32'hc267c083};
test_output[9628] = '{32'h42a3f2b9};
test_index[9628] = '{5};
test_input[77032:77039] = '{32'h4285b4a0, 32'h41aff57f, 32'hc2b5d234, 32'h420c364d, 32'hc2ba4e6c, 32'h429674db, 32'hc0fb618d, 32'h42558e99};
test_output[9629] = '{32'h429674db};
test_index[9629] = '{5};
test_input[77040:77047] = '{32'hc261f3b4, 32'hc24c348e, 32'hc243ad3c, 32'h41cd689a, 32'hc200f357, 32'h4237dfdb, 32'h409050fb, 32'h415448d9};
test_output[9630] = '{32'h4237dfdb};
test_index[9630] = '{5};
test_input[77048:77055] = '{32'h42abcc86, 32'h40aaec96, 32'h4269b8c1, 32'h4107eb68, 32'hc265399f, 32'h42a1b3fc, 32'h421ce806, 32'h42adaf12};
test_output[9631] = '{32'h42adaf12};
test_index[9631] = '{7};
test_input[77056:77063] = '{32'hc26237f0, 32'hc1e40595, 32'hc26efc80, 32'h41e7f759, 32'h42a91f3a, 32'hc11916af, 32'hc1dfee2e, 32'hc0144e13};
test_output[9632] = '{32'h42a91f3a};
test_index[9632] = '{4};
test_input[77064:77071] = '{32'hc2865a49, 32'h4209247c, 32'h42386785, 32'hc2a859f7, 32'hc2637a93, 32'hc2976338, 32'h41e360aa, 32'h42acfdea};
test_output[9633] = '{32'h42acfdea};
test_index[9633] = '{7};
test_input[77072:77079] = '{32'h4289c1df, 32'h425f1966, 32'hc224485f, 32'h424120b5, 32'h41cef170, 32'h4166d099, 32'h428725ba, 32'hc2a41a56};
test_output[9634] = '{32'h4289c1df};
test_index[9634] = '{0};
test_input[77080:77087] = '{32'h428fd4f8, 32'hc20f9188, 32'h41b9f39a, 32'h422d9bab, 32'h4278a267, 32'hc1f0d0f2, 32'hc250beaa, 32'hc1dd7b8c};
test_output[9635] = '{32'h428fd4f8};
test_index[9635] = '{0};
test_input[77088:77095] = '{32'h42a84eb2, 32'h427107fc, 32'h41aaebe0, 32'h4249114b, 32'hc10fda9b, 32'hc29272cd, 32'h41e15c2f, 32'h401bfd2d};
test_output[9636] = '{32'h42a84eb2};
test_index[9636] = '{0};
test_input[77096:77103] = '{32'h42bd0ebb, 32'hc1df040d, 32'hc222a6f0, 32'h41ab8f57, 32'h41defddf, 32'hc2395e98, 32'hc2a047d4, 32'hc1e15ba5};
test_output[9637] = '{32'h42bd0ebb};
test_index[9637] = '{0};
test_input[77104:77111] = '{32'h42c22f1c, 32'hc1a3837b, 32'hc15f1355, 32'hc286164c, 32'h42c4e345, 32'hc1ca1e71, 32'hc261d4cd, 32'hc14f88b5};
test_output[9638] = '{32'h42c4e345};
test_index[9638] = '{4};
test_input[77112:77119] = '{32'h4197ed99, 32'h427f61fc, 32'hc298dca6, 32'hc1427d28, 32'hc28e2b04, 32'h4214ae1f, 32'h421f6c77, 32'hc2956db5};
test_output[9639] = '{32'h427f61fc};
test_index[9639] = '{1};
test_input[77120:77127] = '{32'h41d95ef2, 32'h4253a787, 32'hc2bb0a43, 32'hc2a37e32, 32'hc1bbaef2, 32'hc1e03a47, 32'hc23322f2, 32'hc151def2};
test_output[9640] = '{32'h4253a787};
test_index[9640] = '{1};
test_input[77128:77135] = '{32'hc1e5cb52, 32'hc2b4418f, 32'hc19e735e, 32'h42ac6129, 32'hc29e283c, 32'hc2b9b7f8, 32'h4281e091, 32'hc29d56e9};
test_output[9641] = '{32'h42ac6129};
test_index[9641] = '{3};
test_input[77136:77143] = '{32'h42b9c6d3, 32'h4205ade0, 32'h424e6b6b, 32'h42ab9728, 32'h4042e5c5, 32'h41792507, 32'hc15ce46f, 32'h4265e623};
test_output[9642] = '{32'h42b9c6d3};
test_index[9642] = '{0};
test_input[77144:77151] = '{32'hc05869a5, 32'h42b37e0c, 32'hc2a8941b, 32'h429407e8, 32'hc25b837a, 32'hc28fcadc, 32'hc218ade3, 32'hc29a013d};
test_output[9643] = '{32'h42b37e0c};
test_index[9643] = '{1};
test_input[77152:77159] = '{32'hc2b2e6bb, 32'hc26dfeba, 32'hc20fe360, 32'hc289c3e0, 32'h42c0b041, 32'hc18eb2e9, 32'h425d6cc0, 32'h420ad46a};
test_output[9644] = '{32'h42c0b041};
test_index[9644] = '{4};
test_input[77160:77167] = '{32'hc1b2e742, 32'hc2bb6f03, 32'hc2ad35c3, 32'h41c7da5e, 32'h429b9f14, 32'hc2102c43, 32'hc1754660, 32'h41b3a7ce};
test_output[9645] = '{32'h429b9f14};
test_index[9645] = '{4};
test_input[77168:77175] = '{32'hc1c08991, 32'h3fb9e989, 32'h427e96e3, 32'h42a1aabc, 32'h425246dc, 32'hc298fab0, 32'h401a1e33, 32'hc2489900};
test_output[9646] = '{32'h42a1aabc};
test_index[9646] = '{3};
test_input[77176:77183] = '{32'hc1c7d28d, 32'hc2316f8e, 32'hc24d62ce, 32'h428580fb, 32'hc2a9a636, 32'h41d3e831, 32'hc2becfa4, 32'hc2311200};
test_output[9647] = '{32'h428580fb};
test_index[9647] = '{3};
test_input[77184:77191] = '{32'hc23534c4, 32'hc2b778ec, 32'hc28da451, 32'h42b4006e, 32'h421cd24f, 32'hc2240e83, 32'hc285865b, 32'hc0f08beb};
test_output[9648] = '{32'h42b4006e};
test_index[9648] = '{3};
test_input[77192:77199] = '{32'h422ada5d, 32'h42bf3163, 32'hc231b833, 32'h42116f7e, 32'h428a6365, 32'hc2b12fe5, 32'hc1d127f6, 32'h420104c0};
test_output[9649] = '{32'h42bf3163};
test_index[9649] = '{1};
test_input[77200:77207] = '{32'hc2afff05, 32'hc2a217cb, 32'hc2b8ec30, 32'hc18ee0ae, 32'h40430118, 32'h42872863, 32'hc15c22ec, 32'h42b18b4c};
test_output[9650] = '{32'h42b18b4c};
test_index[9650] = '{7};
test_input[77208:77215] = '{32'h42932f13, 32'h422d5138, 32'hc2129dab, 32'hc2830668, 32'h42799815, 32'hc2a4583e, 32'h42235d61, 32'hc2af359f};
test_output[9651] = '{32'h42932f13};
test_index[9651] = '{0};
test_input[77216:77223] = '{32'hc2a3b4b1, 32'h41f4fc6c, 32'h4278a502, 32'h40c4dc94, 32'h41828f2f, 32'h42329344, 32'h41598a8d, 32'hc27a2ca9};
test_output[9652] = '{32'h4278a502};
test_index[9652] = '{2};
test_input[77224:77231] = '{32'h422f4adf, 32'h4294ca1e, 32'hc1b89140, 32'hc2980aa0, 32'hc1918d84, 32'hc2af9d30, 32'h4117cedd, 32'h4248bd5d};
test_output[9653] = '{32'h4294ca1e};
test_index[9653] = '{1};
test_input[77232:77239] = '{32'h428b52e3, 32'h42a20684, 32'h418fc6f4, 32'hc24a46e6, 32'hc235137b, 32'h42686ff9, 32'h420f1842, 32'hc25fdeb3};
test_output[9654] = '{32'h42a20684};
test_index[9654] = '{1};
test_input[77240:77247] = '{32'h42073841, 32'hc2290f66, 32'h40f42515, 32'hc28b1d2d, 32'h42c0b6dc, 32'hc2bde5ef, 32'h4252c1c3, 32'hc2bf00e6};
test_output[9655] = '{32'h42c0b6dc};
test_index[9655] = '{4};
test_input[77248:77255] = '{32'hc28009e6, 32'hc0f7f579, 32'hc1de13f5, 32'hc03cf7db, 32'h429e8c29, 32'h3fb775cb, 32'hc18ce522, 32'hc2abdf11};
test_output[9656] = '{32'h429e8c29};
test_index[9656] = '{4};
test_input[77256:77263] = '{32'h41815341, 32'h429af92b, 32'hc217e995, 32'hc114c97d, 32'h415c24ca, 32'h41adf52e, 32'h4206e311, 32'h40b3562d};
test_output[9657] = '{32'h429af92b};
test_index[9657] = '{1};
test_input[77264:77271] = '{32'hc268a580, 32'hc267a4c9, 32'h4225b104, 32'hc2060af9, 32'hc29ac1b6, 32'hc28525da, 32'hbe587b08, 32'hc1ed8061};
test_output[9658] = '{32'h4225b104};
test_index[9658] = '{2};
test_input[77272:77279] = '{32'h429cb1d5, 32'hbf92e49b, 32'h424a5109, 32'hc2a187a4, 32'h42a10829, 32'h42b8ba4a, 32'h4280039c, 32'h42a586ae};
test_output[9659] = '{32'h42b8ba4a};
test_index[9659] = '{5};
test_input[77280:77287] = '{32'h41637f85, 32'hc23ce422, 32'h410ac9b5, 32'h42b3070a, 32'hc091abc7, 32'h4293c4c0, 32'h423c3ac2, 32'hc2a9c9bd};
test_output[9660] = '{32'h42b3070a};
test_index[9660] = '{3};
test_input[77288:77295] = '{32'h42befd7e, 32'hc2a11837, 32'h42c496e1, 32'h42c71469, 32'h425c5b3b, 32'hc2119cb0, 32'h42c6a3ad, 32'hc22052ac};
test_output[9661] = '{32'h42c71469};
test_index[9661] = '{3};
test_input[77296:77303] = '{32'h428f60b0, 32'hbfe8d1b8, 32'hc2c58775, 32'h428aaabe, 32'hc2530849, 32'h42c14ab8, 32'h422841ae, 32'h41c8156d};
test_output[9662] = '{32'h42c14ab8};
test_index[9662] = '{5};
test_input[77304:77311] = '{32'hc2871486, 32'hc29bb727, 32'hc27181b6, 32'h42bdb67d, 32'h4096519d, 32'hc1cf5e51, 32'h4259ffc6, 32'h40792eb0};
test_output[9663] = '{32'h42bdb67d};
test_index[9663] = '{3};
test_input[77312:77319] = '{32'hc2431880, 32'h428d50cd, 32'hc27e95e0, 32'h41234a7f, 32'hc2b20ed2, 32'hc0178ecd, 32'h41286840, 32'hc289b661};
test_output[9664] = '{32'h428d50cd};
test_index[9664] = '{1};
test_input[77320:77327] = '{32'h4257e7a9, 32'h4210910d, 32'h3ff4daad, 32'h40fb0e05, 32'h42ac5117, 32'h42c7d8b2, 32'h429db467, 32'h4272f038};
test_output[9665] = '{32'h42c7d8b2};
test_index[9665] = '{5};
test_input[77328:77335] = '{32'h4298fece, 32'hc2ad29c5, 32'hc2b73e34, 32'hc20c6eb9, 32'hc283ee26, 32'hc1e77044, 32'h424f3d30, 32'h4287f902};
test_output[9666] = '{32'h4298fece};
test_index[9666] = '{0};
test_input[77336:77343] = '{32'hc10c41a9, 32'h427f1a35, 32'h4207c735, 32'h42c60255, 32'hc1b82a55, 32'h42670503, 32'h42abba43, 32'hc211f218};
test_output[9667] = '{32'h42c60255};
test_index[9667] = '{3};
test_input[77344:77351] = '{32'h4238dc60, 32'h419454d4, 32'hc2ab4117, 32'hc2adde0f, 32'h425c9e63, 32'h42787687, 32'hc26d2070, 32'hc03bf916};
test_output[9668] = '{32'h42787687};
test_index[9668] = '{5};
test_input[77352:77359] = '{32'h412fe3ac, 32'h4144f636, 32'h41c76c3c, 32'h425bfbc2, 32'h40e4279d, 32'h428aee62, 32'hc0ab584a, 32'h411c57d3};
test_output[9669] = '{32'h428aee62};
test_index[9669] = '{5};
test_input[77360:77367] = '{32'h42a9cd56, 32'h415ba5ce, 32'h4283533e, 32'hc1e9222c, 32'h4286c356, 32'hc2aaa000, 32'hc21c0344, 32'hc2978623};
test_output[9670] = '{32'h42a9cd56};
test_index[9670] = '{0};
test_input[77368:77375] = '{32'hc1f7a2f2, 32'h428ea883, 32'h42801ca4, 32'h4288a7bb, 32'hc271042b, 32'hc28e225d, 32'h42484d10, 32'hc289d607};
test_output[9671] = '{32'h428ea883};
test_index[9671] = '{1};
test_input[77376:77383] = '{32'hc20759de, 32'hc2bd3316, 32'h428c2f00, 32'hbf969279, 32'h4276c8fb, 32'hc22900e8, 32'hc2491db3, 32'h41373354};
test_output[9672] = '{32'h428c2f00};
test_index[9672] = '{2};
test_input[77384:77391] = '{32'h424f5208, 32'hc2c6bc0f, 32'h412c3c3d, 32'h42a6d777, 32'h42962f97, 32'hc24d7761, 32'h42221455, 32'hc2c09686};
test_output[9673] = '{32'h42a6d777};
test_index[9673] = '{3};
test_input[77392:77399] = '{32'h42279cb4, 32'hc20d8122, 32'h426bdd9a, 32'hc0c22603, 32'h42ba1889, 32'hc2235a19, 32'h425b2ab8, 32'hc1ac0da3};
test_output[9674] = '{32'h42ba1889};
test_index[9674] = '{4};
test_input[77400:77407] = '{32'hc2b9bf52, 32'h4148a88c, 32'hc2aa5249, 32'h41d2d1b4, 32'h41ea5cdd, 32'h427d4f14, 32'hc1e0cba2, 32'hc178134d};
test_output[9675] = '{32'h427d4f14};
test_index[9675] = '{5};
test_input[77408:77415] = '{32'h42506c1b, 32'hc09e1aec, 32'h415b4208, 32'h426c7590, 32'h4159ee26, 32'h408121be, 32'hc2806f90, 32'h4196a045};
test_output[9676] = '{32'h426c7590};
test_index[9676] = '{3};
test_input[77416:77423] = '{32'hc281ba4c, 32'h40f8092a, 32'h420185b4, 32'hc290b6a8, 32'h425563cd, 32'h429912af, 32'hc2bbdebc, 32'hc21cddd2};
test_output[9677] = '{32'h429912af};
test_index[9677] = '{5};
test_input[77424:77431] = '{32'hc2b223ba, 32'hc280f122, 32'h42c340aa, 32'hc27f1ae9, 32'hc2a554b5, 32'hc294a1f4, 32'h429dee11, 32'h42419e44};
test_output[9678] = '{32'h42c340aa};
test_index[9678] = '{2};
test_input[77432:77439] = '{32'hc2919ac9, 32'h42c4fe98, 32'hc29c7c82, 32'h41d91cd9, 32'hc2904d9a, 32'hc19ccc4b, 32'hc0bd6d51, 32'h4237299f};
test_output[9679] = '{32'h42c4fe98};
test_index[9679] = '{1};
test_input[77440:77447] = '{32'h427012cd, 32'hc234768f, 32'h42bb8142, 32'h41b9b367, 32'h423271f0, 32'hc2b5b982, 32'hc2270003, 32'h426c284e};
test_output[9680] = '{32'h42bb8142};
test_index[9680] = '{2};
test_input[77448:77455] = '{32'hc261dc9b, 32'hc2258827, 32'hc1c3b36b, 32'hc2363159, 32'h422bb6e3, 32'hc03ded63, 32'h41032c67, 32'h42bdf5ab};
test_output[9681] = '{32'h42bdf5ab};
test_index[9681] = '{7};
test_input[77456:77463] = '{32'hc164cb80, 32'hc0e17292, 32'hc28ed9cb, 32'h42021569, 32'h425c4222, 32'h42ac063b, 32'hc2c4de55, 32'hc291119e};
test_output[9682] = '{32'h42ac063b};
test_index[9682] = '{5};
test_input[77464:77471] = '{32'hc2c0e790, 32'hc29cd07c, 32'hc22ed3be, 32'hc1ecd0b2, 32'h4076ebb5, 32'hc0c6f3a5, 32'h429bfa02, 32'hc2550f2d};
test_output[9683] = '{32'h429bfa02};
test_index[9683] = '{6};
test_input[77472:77479] = '{32'h42824d75, 32'hc1274076, 32'h42c14652, 32'hc21485d2, 32'hc23a3bbc, 32'h42ab28f9, 32'h421cef20, 32'h428b22d1};
test_output[9684] = '{32'h42c14652};
test_index[9684] = '{2};
test_input[77480:77487] = '{32'h42a96005, 32'h41997940, 32'h42672558, 32'h4202a903, 32'hc10f5c0d, 32'h425c2059, 32'hc2246ff8, 32'hc24214cf};
test_output[9685] = '{32'h42a96005};
test_index[9685] = '{0};
test_input[77488:77495] = '{32'h41532c28, 32'h4288efd1, 32'h420de5e0, 32'h4281ae18, 32'h420bea17, 32'hc2806aa5, 32'h429c3e8b, 32'h41b49d7c};
test_output[9686] = '{32'h429c3e8b};
test_index[9686] = '{6};
test_input[77496:77503] = '{32'h42837c31, 32'hc1bec252, 32'hc21d9f44, 32'h41fdf3d4, 32'h4258006d, 32'h42b315af, 32'hc27c1cb7, 32'h3e824206};
test_output[9687] = '{32'h42b315af};
test_index[9687] = '{5};
test_input[77504:77511] = '{32'hc173eecc, 32'h42aaa26c, 32'h40ae78c6, 32'hc238b625, 32'hc1b1ed95, 32'h419ce16d, 32'h41166a4a, 32'h41e95ddc};
test_output[9688] = '{32'h42aaa26c};
test_index[9688] = '{1};
test_input[77512:77519] = '{32'h42c21d98, 32'hc28a5018, 32'h425ff489, 32'hc2bd5f37, 32'hc1aeabbe, 32'hc2b6d672, 32'hc1a1d922, 32'h42b9d5c9};
test_output[9689] = '{32'h42c21d98};
test_index[9689] = '{0};
test_input[77520:77527] = '{32'hc297b0b4, 32'h42aa366b, 32'hc04f11b8, 32'hc288f5b7, 32'hc1901ab4, 32'hc204b7e1, 32'h41c02bf9, 32'h4221cf63};
test_output[9690] = '{32'h42aa366b};
test_index[9690] = '{1};
test_input[77528:77535] = '{32'h41bd7181, 32'hc23c79c3, 32'hc227153f, 32'hc272ba1f, 32'h42a593d6, 32'hc2847e9d, 32'h42b82c0c, 32'h42819e93};
test_output[9691] = '{32'h42b82c0c};
test_index[9691] = '{6};
test_input[77536:77543] = '{32'h4294c14a, 32'h3f4d22bc, 32'hc29dc661, 32'hc27b24df, 32'hc217da58, 32'hc08fd6b3, 32'hc2b5623e, 32'h42bf20bd};
test_output[9692] = '{32'h42bf20bd};
test_index[9692] = '{7};
test_input[77544:77551] = '{32'h42b8f275, 32'hc2c0d602, 32'h429fe6a7, 32'hc0b9373c, 32'hc1b75e1a, 32'h418cdba6, 32'h427bc681, 32'hc23603d7};
test_output[9693] = '{32'h42b8f275};
test_index[9693] = '{0};
test_input[77552:77559] = '{32'h42945095, 32'hc0f1c1f0, 32'h4261590c, 32'h4189fb27, 32'hc27b8c5f, 32'h41d5aa92, 32'h41ac5692, 32'h412ea7dc};
test_output[9694] = '{32'h42945095};
test_index[9694] = '{0};
test_input[77560:77567] = '{32'h422f7aa8, 32'h40b4717b, 32'hc18a529f, 32'h42a57175, 32'hc247159d, 32'h42209b83, 32'h42b17570, 32'h41a2efc6};
test_output[9695] = '{32'h42b17570};
test_index[9695] = '{6};
test_input[77568:77575] = '{32'h429ab6a7, 32'h42a53334, 32'h4289f5c6, 32'hc2ae03e6, 32'h42b145eb, 32'hbf3a5043, 32'hc244bee7, 32'hc086df9b};
test_output[9696] = '{32'h42b145eb};
test_index[9696] = '{4};
test_input[77576:77583] = '{32'hc22d6652, 32'h42958cb9, 32'h429b81d7, 32'h40df4a0d, 32'hbe832ca0, 32'hc1dc44bb, 32'hc1875afc, 32'h41674ed9};
test_output[9697] = '{32'h429b81d7};
test_index[9697] = '{2};
test_input[77584:77591] = '{32'h425f16f0, 32'hc2aa3135, 32'hc13a2eaa, 32'hc1a90deb, 32'hc223aafe, 32'hc14e4a32, 32'h4201e81a, 32'h41dee26e};
test_output[9698] = '{32'h425f16f0};
test_index[9698] = '{0};
test_input[77592:77599] = '{32'hc04034a4, 32'hc127783e, 32'h429fe300, 32'h428441d7, 32'hc235e41e, 32'hc28dec4a, 32'h41e1d6e2, 32'h42832872};
test_output[9699] = '{32'h429fe300};
test_index[9699] = '{2};
test_input[77600:77607] = '{32'h41fa9f18, 32'hc1ce49d3, 32'h41b88dfa, 32'hc28457bd, 32'h42bd8c7d, 32'hc29650e0, 32'hc2a41993, 32'hc2908c19};
test_output[9700] = '{32'h42bd8c7d};
test_index[9700] = '{4};
test_input[77608:77615] = '{32'hc2804a2e, 32'h428b95e6, 32'hc26c1b04, 32'h428de65e, 32'h42a9e8d4, 32'h4279d023, 32'hc1a1acc4, 32'h42bc800b};
test_output[9701] = '{32'h42bc800b};
test_index[9701] = '{7};
test_input[77616:77623] = '{32'h422d4930, 32'h41f7c129, 32'h428c4da1, 32'h42b9178c, 32'hc260514d, 32'h42aa05dd, 32'h419a8fcb, 32'h42421727};
test_output[9702] = '{32'h42b9178c};
test_index[9702] = '{3};
test_input[77624:77631] = '{32'h42c2feb6, 32'h42bd868e, 32'hc1953437, 32'hc2b1af28, 32'hc2980eff, 32'h429d496f, 32'h41e795f7, 32'hc0f3c4e7};
test_output[9703] = '{32'h42c2feb6};
test_index[9703] = '{0};
test_input[77632:77639] = '{32'h410cfb62, 32'h4133698d, 32'hc22d6ea3, 32'hc2332c2d, 32'h4251fde9, 32'h422aa2f1, 32'h4232c23e, 32'h42729b54};
test_output[9704] = '{32'h42729b54};
test_index[9704] = '{7};
test_input[77640:77647] = '{32'h3f99a04a, 32'h4083da89, 32'hc2649544, 32'h42193063, 32'h42c62331, 32'hc2c73296, 32'h42b12438, 32'h424497ae};
test_output[9705] = '{32'h42c62331};
test_index[9705] = '{4};
test_input[77648:77655] = '{32'h42802f74, 32'hc273ca79, 32'hc2a43224, 32'h41e854f0, 32'h41d0697a, 32'h4264949c, 32'hc250d073, 32'hc289b8bd};
test_output[9706] = '{32'h42802f74};
test_index[9706] = '{0};
test_input[77656:77663] = '{32'h427d26eb, 32'hc2bfa3a7, 32'h41197a44, 32'h4208e69d, 32'hc103f0bf, 32'h41bee7f2, 32'h418ad231, 32'hc2c22887};
test_output[9707] = '{32'h427d26eb};
test_index[9707] = '{0};
test_input[77664:77671] = '{32'hc1b87063, 32'hc2468441, 32'h42aafbfe, 32'h425fe46d, 32'hc1f130dc, 32'h41797c80, 32'hc2b35beb, 32'hc212f483};
test_output[9708] = '{32'h42aafbfe};
test_index[9708] = '{2};
test_input[77672:77679] = '{32'hc1def35c, 32'hc19f770d, 32'hc2b45768, 32'h4258fb89, 32'h42c3713a, 32'h42486cb2, 32'hc28f19e1, 32'hc17de266};
test_output[9709] = '{32'h42c3713a};
test_index[9709] = '{4};
test_input[77680:77687] = '{32'h422bf407, 32'hc2795499, 32'h41aa9a42, 32'hc0df4488, 32'hc2a0013d, 32'h4226bc85, 32'hc2084de0, 32'h40acccfd};
test_output[9710] = '{32'h422bf407};
test_index[9710] = '{0};
test_input[77688:77695] = '{32'h42a7f99b, 32'h429689d9, 32'h42854489, 32'hc1e7c52e, 32'hc29c992a, 32'h427d8e35, 32'hc29ec2a1, 32'h41910b25};
test_output[9711] = '{32'h42a7f99b};
test_index[9711] = '{0};
test_input[77696:77703] = '{32'hc1a9e813, 32'h42bfe378, 32'hc283f6ea, 32'h425ab6bf, 32'hc27454ba, 32'h427da996, 32'h4297863a, 32'h424adbf9};
test_output[9712] = '{32'h42bfe378};
test_index[9712] = '{1};
test_input[77704:77711] = '{32'hc2b2b391, 32'hc2b079f4, 32'h425f1543, 32'h41d5140c, 32'h413d4669, 32'hc2214de6, 32'h42322149, 32'h426900b4};
test_output[9713] = '{32'h426900b4};
test_index[9713] = '{7};
test_input[77712:77719] = '{32'hc0727ffd, 32'h40eda5c7, 32'h424a74da, 32'h42b4f7fa, 32'hc01b4b12, 32'hc2a22f70, 32'hc180177b, 32'hc272f687};
test_output[9714] = '{32'h42b4f7fa};
test_index[9714] = '{3};
test_input[77720:77727] = '{32'hc1dae445, 32'h417189b6, 32'hc0b83296, 32'hc2c521df, 32'hc1b62ab4, 32'h42147fbd, 32'hc202a4ed, 32'hc231eef6};
test_output[9715] = '{32'h42147fbd};
test_index[9715] = '{5};
test_input[77728:77735] = '{32'hc1a0cd3d, 32'h421c31f5, 32'h416dc5ad, 32'h42704ea0, 32'hc27ad9e5, 32'h42c635c8, 32'h41a85a0e, 32'hc1e763f7};
test_output[9716] = '{32'h42c635c8};
test_index[9716] = '{5};
test_input[77736:77743] = '{32'hc286386b, 32'h429eb943, 32'h42921240, 32'hc2b8e7d0, 32'hc2c3b21f, 32'h428c483f, 32'h425208c4, 32'hc256d7ca};
test_output[9717] = '{32'h429eb943};
test_index[9717] = '{1};
test_input[77744:77751] = '{32'hc216f5bc, 32'hc20d0773, 32'hc295596d, 32'hc2a94375, 32'hc2a86000, 32'h4281c622, 32'hc292b081, 32'hc228119e};
test_output[9718] = '{32'h4281c622};
test_index[9718] = '{5};
test_input[77752:77759] = '{32'h42594729, 32'hc2c4f0ca, 32'h41e178ac, 32'hc2c73bb7, 32'hc2b27b82, 32'hc1cd153c, 32'hc16b8125, 32'hc2bce727};
test_output[9719] = '{32'h42594729};
test_index[9719] = '{0};
test_input[77760:77767] = '{32'hc290f447, 32'h426ae8ee, 32'hc286666a, 32'h41eb4a49, 32'hc2c0867c, 32'h412bb54c, 32'hc28bb1ae, 32'h429c7c27};
test_output[9720] = '{32'h429c7c27};
test_index[9720] = '{7};
test_input[77768:77775] = '{32'hc2852f94, 32'hc295df8f, 32'hc20e24bf, 32'h42b4538a, 32'hc2878f7d, 32'hc19ef017, 32'hc1e5f7c7, 32'hc2afc99a};
test_output[9721] = '{32'h42b4538a};
test_index[9721] = '{3};
test_input[77776:77783] = '{32'h4163cfef, 32'h420558ba, 32'hc2ac82ff, 32'h42ac09c4, 32'h41331a6b, 32'hc2ab12c6, 32'h42531f3a, 32'hc0d04f83};
test_output[9722] = '{32'h42ac09c4};
test_index[9722] = '{3};
test_input[77784:77791] = '{32'hbf191783, 32'h42254c2c, 32'h4213f1c6, 32'hc28869de, 32'hc25e3b11, 32'h418884e2, 32'hc22f1f78, 32'h4254e385};
test_output[9723] = '{32'h4254e385};
test_index[9723] = '{7};
test_input[77792:77799] = '{32'h4288b872, 32'h42ba7e2f, 32'h424c2ea5, 32'hc2530fc6, 32'h41edd6be, 32'h428b8bcb, 32'hc2379e3d, 32'h4112a70c};
test_output[9724] = '{32'h42ba7e2f};
test_index[9724] = '{1};
test_input[77800:77807] = '{32'hc2ad5990, 32'hc2ac44f2, 32'h42179d66, 32'hc1f834d5, 32'hc28c6e2e, 32'h3f961762, 32'h4213738b, 32'h42be8407};
test_output[9725] = '{32'h42be8407};
test_index[9725] = '{7};
test_input[77808:77815] = '{32'h42196292, 32'hc200f697, 32'hc289c369, 32'h4283c6a6, 32'h41a6842d, 32'h4225bc3c, 32'hc29798a8, 32'hc004c179};
test_output[9726] = '{32'h4283c6a6};
test_index[9726] = '{3};
test_input[77816:77823] = '{32'h4177f467, 32'hc26a9590, 32'hc038fc25, 32'hc2807ede, 32'hc0153ef4, 32'hc09e4c1a, 32'h42a174f1, 32'h409fb664};
test_output[9727] = '{32'h42a174f1};
test_index[9727] = '{6};
test_input[77824:77831] = '{32'hc181e705, 32'h427e6b33, 32'hc2646e61, 32'h41c2270c, 32'h4287f5f1, 32'hc2a492b5, 32'h4220f231, 32'hc101e01f};
test_output[9728] = '{32'h4287f5f1};
test_index[9728] = '{4};
test_input[77832:77839] = '{32'hc2c700f6, 32'hc2475ba0, 32'h40dcd31c, 32'hc23098b2, 32'hc0f37d73, 32'hc2bf9089, 32'hc2a009fa, 32'hc282df5a};
test_output[9729] = '{32'h40dcd31c};
test_index[9729] = '{2};
test_input[77840:77847] = '{32'h425546b6, 32'hc217beff, 32'h42c3fafb, 32'hc2b36bfb, 32'h415450db, 32'hc2b60551, 32'h424868da, 32'hc1057146};
test_output[9730] = '{32'h42c3fafb};
test_index[9730] = '{2};
test_input[77848:77855] = '{32'h429fd65b, 32'hc2a679b3, 32'hc16c9d52, 32'hc21a0afe, 32'hc2a5aa8d, 32'hc2049de6, 32'hc1cbbf25, 32'h42b55cbd};
test_output[9731] = '{32'h42b55cbd};
test_index[9731] = '{7};
test_input[77856:77863] = '{32'h42218a6c, 32'hc1581145, 32'hc1c84aa8, 32'h41fa0eb1, 32'h4293627a, 32'h429bbf1d, 32'hc0bad572, 32'hc2095c14};
test_output[9732] = '{32'h429bbf1d};
test_index[9732] = '{5};
test_input[77864:77871] = '{32'hc204297c, 32'hc2a974bf, 32'hc283bb04, 32'hbf0a8e2d, 32'hc050c590, 32'h4296f8f6, 32'hc2b0cb69, 32'h42a2025b};
test_output[9733] = '{32'h42a2025b};
test_index[9733] = '{7};
test_input[77872:77879] = '{32'hc29713a3, 32'h4204f485, 32'h42845123, 32'hc12f721b, 32'hc29dbac6, 32'h42b9833d, 32'hc2665de2, 32'hc202fdc8};
test_output[9734] = '{32'h42b9833d};
test_index[9734] = '{5};
test_input[77880:77887] = '{32'hc2267dcf, 32'hc1b93ce1, 32'hc20aaa3e, 32'h423e79d3, 32'hc032817e, 32'h42b3ed0d, 32'h4271176f, 32'h42b002bf};
test_output[9735] = '{32'h42b3ed0d};
test_index[9735] = '{5};
test_input[77888:77895] = '{32'hc2b5a64e, 32'h410783b7, 32'hc148fff3, 32'hc25d4c26, 32'h424461e0, 32'h42760798, 32'hc29edaaa, 32'h426ab915};
test_output[9736] = '{32'h42760798};
test_index[9736] = '{5};
test_input[77896:77903] = '{32'hc27e770b, 32'h42144ad8, 32'h41c98f9a, 32'h41d5d1fb, 32'hc25ac5cc, 32'hc17b9736, 32'hc2a7dc03, 32'h42506000};
test_output[9737] = '{32'h42506000};
test_index[9737] = '{7};
test_input[77904:77911] = '{32'hc2a19bab, 32'h42703244, 32'h42a937c9, 32'h428d419f, 32'hc2580220, 32'hc22f3eb7, 32'h4152bdd5, 32'hc25585ea};
test_output[9738] = '{32'h42a937c9};
test_index[9738] = '{2};
test_input[77912:77919] = '{32'hc0c69e49, 32'h423f1eb7, 32'hc28efeec, 32'h41f3817a, 32'hc29e2130, 32'h42a3e9e6, 32'h42699dd5, 32'hc1f86d41};
test_output[9739] = '{32'h42a3e9e6};
test_index[9739] = '{5};
test_input[77920:77927] = '{32'hc28c17e9, 32'h429316ed, 32'hc1546d09, 32'hc29b5241, 32'hc2a0cae1, 32'h428e54fc, 32'hc26d5e6f, 32'h3f89ed3d};
test_output[9740] = '{32'h429316ed};
test_index[9740] = '{1};
test_input[77928:77935] = '{32'h4167de1c, 32'hc298fe7c, 32'hc28ea8e1, 32'h418f6099, 32'hc1e739a9, 32'hc28056f8, 32'h409b3521, 32'hc2266252};
test_output[9741] = '{32'h418f6099};
test_index[9741] = '{3};
test_input[77936:77943] = '{32'hc2807dd3, 32'h41a95118, 32'hc15aad83, 32'hc24a2b63, 32'hc01789bf, 32'hc1a943e1, 32'h4206a301, 32'hc267b41d};
test_output[9742] = '{32'h4206a301};
test_index[9742] = '{6};
test_input[77944:77951] = '{32'h423fd6f3, 32'hc1cd60b9, 32'h42be9c05, 32'hc2ba0a91, 32'hc23f5007, 32'hc221ce99, 32'hc294884b, 32'h41ef22a7};
test_output[9743] = '{32'h42be9c05};
test_index[9743] = '{2};
test_input[77952:77959] = '{32'h42bfcc9c, 32'h421c1662, 32'hc1b9b281, 32'h42a8d66a, 32'hbf25dcdc, 32'hc1065e18, 32'hc1ffa890, 32'hc2079349};
test_output[9744] = '{32'h42bfcc9c};
test_index[9744] = '{0};
test_input[77960:77967] = '{32'h42ad3642, 32'h42a1c9fe, 32'hc19ebe80, 32'h429846ed, 32'hc1fcb145, 32'hc20acb21, 32'hc1d1ec90, 32'hc291f2cb};
test_output[9745] = '{32'h42ad3642};
test_index[9745] = '{0};
test_input[77968:77975] = '{32'hc265b2df, 32'hc17e262e, 32'h42c45faa, 32'h4294ef58, 32'hc2c7160b, 32'h4240fb51, 32'h42849d3d, 32'hc25979a0};
test_output[9746] = '{32'h42c45faa};
test_index[9746] = '{2};
test_input[77976:77983] = '{32'hc18b5654, 32'h42a6793b, 32'hc25179ad, 32'h4297f9ce, 32'h4203bca8, 32'h428c9962, 32'hc2ac273f, 32'hc2adcf55};
test_output[9747] = '{32'h42a6793b};
test_index[9747] = '{1};
test_input[77984:77991] = '{32'h42a54d18, 32'hc16cbae1, 32'h4084d5d9, 32'h42b8b1dd, 32'hc2934edb, 32'hc2adfa65, 32'h42929f8a, 32'h41c57d5a};
test_output[9748] = '{32'h42b8b1dd};
test_index[9748] = '{3};
test_input[77992:77999] = '{32'hc2b28ef6, 32'hbf85fc36, 32'hc0878e08, 32'h428f2618, 32'h42a9a299, 32'h41a17b6e, 32'hc297ad5a, 32'h42a985e4};
test_output[9749] = '{32'h42a9a299};
test_index[9749] = '{4};
test_input[78000:78007] = '{32'h42a89376, 32'h41434446, 32'h4026883a, 32'hc287b110, 32'h426570ee, 32'hc28d94cf, 32'hc27bfd86, 32'hc296099b};
test_output[9750] = '{32'h42a89376};
test_index[9750] = '{0};
test_input[78008:78015] = '{32'h40c30306, 32'h419d0582, 32'hc2843553, 32'hc202959e, 32'h419d2378, 32'h41a122f3, 32'h42856c91, 32'hc207e775};
test_output[9751] = '{32'h42856c91};
test_index[9751] = '{6};
test_input[78016:78023] = '{32'h424aadc3, 32'h429dc665, 32'h429c0efe, 32'h42195760, 32'hc276f755, 32'h420ddd46, 32'h4291fbf0, 32'h4295f2fe};
test_output[9752] = '{32'h429dc665};
test_index[9752] = '{1};
test_input[78024:78031] = '{32'h42987bc2, 32'hc12df6e6, 32'h424356c1, 32'hc2a8d5d0, 32'h420b1e12, 32'h429e9f1c, 32'hc1e37315, 32'h425199c9};
test_output[9753] = '{32'h429e9f1c};
test_index[9753] = '{5};
test_input[78032:78039] = '{32'h429c3124, 32'hc2067037, 32'hc2bb073e, 32'h423dfb5b, 32'h42ba1ee0, 32'hc1c8dd8e, 32'hc287b967, 32'h42ad31ad};
test_output[9754] = '{32'h42ba1ee0};
test_index[9754] = '{4};
test_input[78040:78047] = '{32'h40d64537, 32'h4205c329, 32'hc22d665b, 32'hc295708b, 32'h42b4a6b8, 32'hc02c47c8, 32'hbfea8e33, 32'h4253b3a4};
test_output[9755] = '{32'h42b4a6b8};
test_index[9755] = '{4};
test_input[78048:78055] = '{32'h4291086f, 32'h42512bf5, 32'hc2a38db8, 32'h42af4526, 32'hc25c400c, 32'hc29c9921, 32'h423ad4a3, 32'h42c235aa};
test_output[9756] = '{32'h42c235aa};
test_index[9756] = '{7};
test_input[78056:78063] = '{32'h41543539, 32'h42c1ed29, 32'h42b0f94a, 32'hc20c60f0, 32'hc27b3732, 32'hc29f2994, 32'h424de43c, 32'h40f3592b};
test_output[9757] = '{32'h42c1ed29};
test_index[9757] = '{1};
test_input[78064:78071] = '{32'h41e13ce6, 32'hc2a4e07c, 32'hc279787e, 32'h418c2b47, 32'h42292c2b, 32'hc1d5fa09, 32'h41d15983, 32'h42ae5e22};
test_output[9758] = '{32'h42ae5e22};
test_index[9758] = '{7};
test_input[78072:78079] = '{32'h419c738f, 32'h41fed2f7, 32'hc23addb9, 32'h429056eb, 32'h4282ae29, 32'hc2c66468, 32'hc2959fa6, 32'h42b5a994};
test_output[9759] = '{32'h42b5a994};
test_index[9759] = '{7};
test_input[78080:78087] = '{32'hc29b907d, 32'h4246bdd8, 32'hc28fbacf, 32'hc2bdbbe4, 32'h42c5e492, 32'h41981f76, 32'h421cca06, 32'hc1aa1c6b};
test_output[9760] = '{32'h42c5e492};
test_index[9760] = '{4};
test_input[78088:78095] = '{32'hc2b6190f, 32'h41a9eb67, 32'hc270ecce, 32'h4252cfca, 32'h423877cc, 32'h41167003, 32'hc2adf628, 32'hc199c931};
test_output[9761] = '{32'h4252cfca};
test_index[9761] = '{3};
test_input[78096:78103] = '{32'h4080f9d2, 32'h42a60df2, 32'hc20891c0, 32'hc1eaca97, 32'h422e4239, 32'hc1ffc958, 32'hc2ac1a8f, 32'hc2960ccd};
test_output[9762] = '{32'h42a60df2};
test_index[9762] = '{1};
test_input[78104:78111] = '{32'h4034040a, 32'h42c125aa, 32'hbf973edd, 32'h415a1de3, 32'hc2087a3c, 32'hc2365823, 32'hc29ecbe8, 32'h4286eac7};
test_output[9763] = '{32'h42c125aa};
test_index[9763] = '{1};
test_input[78112:78119] = '{32'h42732cd6, 32'h42bdc853, 32'hc2c6cae3, 32'h41bc62e8, 32'h4251bea5, 32'hc2400345, 32'hc26693aa, 32'h42714dd3};
test_output[9764] = '{32'h42bdc853};
test_index[9764] = '{1};
test_input[78120:78127] = '{32'hc22bba15, 32'hc251daff, 32'h428e41ca, 32'hc2830e5f, 32'h429cccc0, 32'h4245da06, 32'hc1db5c96, 32'hc2492487};
test_output[9765] = '{32'h429cccc0};
test_index[9765] = '{4};
test_input[78128:78135] = '{32'hc284fdac, 32'h420f1307, 32'hc2a81245, 32'h42a51110, 32'hc1a55085, 32'h409ddc99, 32'h42860f9a, 32'hc2847e19};
test_output[9766] = '{32'h42a51110};
test_index[9766] = '{3};
test_input[78136:78143] = '{32'hc2af1999, 32'h42be7362, 32'h42b1168f, 32'hc1aeac59, 32'hc28a5b18, 32'hc29c4b0d, 32'h42229b36, 32'hbf90d270};
test_output[9767] = '{32'h42be7362};
test_index[9767] = '{1};
test_input[78144:78151] = '{32'h429b537d, 32'hc264830c, 32'hc29ca6a8, 32'hc27f923a, 32'hc1b3c511, 32'h412c0e5f, 32'h42a245e2, 32'hc2c411d7};
test_output[9768] = '{32'h42a245e2};
test_index[9768] = '{6};
test_input[78152:78159] = '{32'hc1cd8b8c, 32'hc12ec743, 32'h42a715d3, 32'h3f93d658, 32'h41e70d00, 32'h4248863b, 32'hc21f32d6, 32'hc297ed50};
test_output[9769] = '{32'h42a715d3};
test_index[9769] = '{2};
test_input[78160:78167] = '{32'hc2b0c86c, 32'hc22086cc, 32'hc14804c9, 32'hc0f84644, 32'h42bb4484, 32'h4236328e, 32'hc2510de7, 32'h4254e195};
test_output[9770] = '{32'h42bb4484};
test_index[9770] = '{4};
test_input[78168:78175] = '{32'hc253e827, 32'h429a7b31, 32'hc297a8e1, 32'h41c48f32, 32'hc27305f5, 32'h41fc3700, 32'hc0a424cf, 32'hbf03bed4};
test_output[9771] = '{32'h429a7b31};
test_index[9771] = '{1};
test_input[78176:78183] = '{32'hc289360d, 32'hc2c386d9, 32'hc200d4a3, 32'h4167869f, 32'h414e7edb, 32'hc1a16dc0, 32'hc299b337, 32'hc21ddb00};
test_output[9772] = '{32'h4167869f};
test_index[9772] = '{3};
test_input[78184:78191] = '{32'h42b70b53, 32'h4297d353, 32'h41712fe9, 32'hc29c26c3, 32'h41fd7d67, 32'hc1506dc0, 32'h428b595f, 32'hc04a37fb};
test_output[9773] = '{32'h42b70b53};
test_index[9773] = '{0};
test_input[78192:78199] = '{32'hc0e34f0b, 32'hc2c7091e, 32'h40826536, 32'hc2af13ec, 32'h42a53135, 32'hc21ce314, 32'h42559e24, 32'h42b052c7};
test_output[9774] = '{32'h42b052c7};
test_index[9774] = '{7};
test_input[78200:78207] = '{32'h4200a762, 32'hc185e630, 32'h421a216c, 32'hc28fa14d, 32'hc2337540, 32'h427243e4, 32'h423532b1, 32'h4244ad54};
test_output[9775] = '{32'h427243e4};
test_index[9775] = '{5};
test_input[78208:78215] = '{32'hc0f307a3, 32'hc2806af7, 32'hc11add9b, 32'h410e4bc7, 32'h427f8d0e, 32'hc275f295, 32'h41fa84b0, 32'h42967b84};
test_output[9776] = '{32'h42967b84};
test_index[9776] = '{7};
test_input[78216:78223] = '{32'hc2b8e872, 32'hc2b1a316, 32'hc2998c73, 32'hc1a704e2, 32'hc2bf588e, 32'hc1c8c6fc, 32'hc22b8e9d, 32'hc28113ee};
test_output[9777] = '{32'hc1a704e2};
test_index[9777] = '{3};
test_input[78224:78231] = '{32'hc104b1e3, 32'h4200f66a, 32'hc2053b6b, 32'hc2813001, 32'h4290235a, 32'h42c76fe1, 32'hc1382fa1, 32'hc2ab4835};
test_output[9778] = '{32'h42c76fe1};
test_index[9778] = '{5};
test_input[78232:78239] = '{32'h41921a07, 32'h4290c557, 32'h42aeb5e4, 32'h42b5665a, 32'hc11bb90c, 32'h42c55ff9, 32'hc2a435f0, 32'hc1c0d01b};
test_output[9779] = '{32'h42c55ff9};
test_index[9779] = '{5};
test_input[78240:78247] = '{32'h41538597, 32'hbf825cce, 32'h429cfde6, 32'h418b2c66, 32'h4269d4ac, 32'hc2228cb6, 32'h41d0de9d, 32'hc211f449};
test_output[9780] = '{32'h429cfde6};
test_index[9780] = '{2};
test_input[78248:78255] = '{32'h42a39d1d, 32'hc28ba391, 32'hc246cbd2, 32'h42a50bf7, 32'hc288f977, 32'hc199a0cf, 32'h41f89a4a, 32'hc221b04a};
test_output[9781] = '{32'h42a50bf7};
test_index[9781] = '{3};
test_input[78256:78263] = '{32'h42c6f27e, 32'hc24d4096, 32'h42aa5a71, 32'hc183a8c8, 32'h427ed415, 32'hc2326973, 32'hc2865467, 32'h429c072d};
test_output[9782] = '{32'h42c6f27e};
test_index[9782] = '{0};
test_input[78264:78271] = '{32'hc2911b8a, 32'hc256f76b, 32'h424053fb, 32'hc1c1c354, 32'hc26ae5b1, 32'hc2b4c059, 32'h426c9c2b, 32'hc19df148};
test_output[9783] = '{32'h426c9c2b};
test_index[9783] = '{6};
test_input[78272:78279] = '{32'h425c00e8, 32'hc28b2834, 32'h427a6cd3, 32'h421c2d71, 32'hc1dca5fb, 32'hc1e5b721, 32'h4226495e, 32'hc1d10e38};
test_output[9784] = '{32'h427a6cd3};
test_index[9784] = '{2};
test_input[78280:78287] = '{32'hc2148b33, 32'h422e2f0f, 32'h418f2f96, 32'h4299349f, 32'h42b03c6d, 32'h410c92c7, 32'hc2559df3, 32'hc289bf51};
test_output[9785] = '{32'h42b03c6d};
test_index[9785] = '{4};
test_input[78288:78295] = '{32'h423fdeca, 32'h418baebc, 32'h420269d1, 32'h4009fe8a, 32'hc286f20b, 32'h42860d3f, 32'hc25a801a, 32'hc259a06f};
test_output[9786] = '{32'h42860d3f};
test_index[9786] = '{5};
test_input[78296:78303] = '{32'hc10ab48e, 32'hc287493e, 32'h41d7322d, 32'hc2b4f10f, 32'hc21daa24, 32'h429c4db9, 32'h42b5df90, 32'h42b5cb4a};
test_output[9787] = '{32'h42b5df90};
test_index[9787] = '{6};
test_input[78304:78311] = '{32'h413d9002, 32'hc205b4b0, 32'h4201ba95, 32'hc26afa2a, 32'h42afb1a9, 32'hc2949a54, 32'hc2b21269, 32'h428320d7};
test_output[9788] = '{32'h42afb1a9};
test_index[9788] = '{4};
test_input[78312:78319] = '{32'hc073592b, 32'hc299c02e, 32'h41e13281, 32'h419a608d, 32'hc216a638, 32'h421018e8, 32'hc21c2bf7, 32'hc224f73e};
test_output[9789] = '{32'h421018e8};
test_index[9789] = '{5};
test_input[78320:78327] = '{32'hc128b532, 32'hc197ac06, 32'hc28a040c, 32'hc2807ed3, 32'hc26ccaeb, 32'hc2acf1a9, 32'h42c1f7f0, 32'hc2641b35};
test_output[9790] = '{32'h42c1f7f0};
test_index[9790] = '{6};
test_input[78328:78335] = '{32'h428979d5, 32'h42bb0b5d, 32'hc2829de5, 32'hc00f7ed8, 32'h41f01825, 32'hc07929a6, 32'hc21eccdc, 32'hc1e09a2e};
test_output[9791] = '{32'h42bb0b5d};
test_index[9791] = '{1};
test_input[78336:78343] = '{32'h414ed997, 32'hc2916e03, 32'hc2052db3, 32'h42848826, 32'h41b69e50, 32'h421b0847, 32'hbe06905d, 32'hc28d1412};
test_output[9792] = '{32'h42848826};
test_index[9792] = '{3};
test_input[78344:78351] = '{32'hc269d386, 32'hc23eed40, 32'hc1c9093f, 32'hc25d218d, 32'hc283c4e6, 32'hc1e02f67, 32'h41e76dbe, 32'hc2433ecc};
test_output[9793] = '{32'h41e76dbe};
test_index[9793] = '{6};
test_input[78352:78359] = '{32'hc1be3a4b, 32'h420d6b89, 32'hc28787a3, 32'hc0e0703e, 32'h42b5ae9a, 32'hc21c702c, 32'hc1e41228, 32'h411b24d5};
test_output[9794] = '{32'h42b5ae9a};
test_index[9794] = '{4};
test_input[78360:78367] = '{32'hbe72683e, 32'hc1bf0e05, 32'hc27b34f4, 32'hc2a083cb, 32'hc19c6dcd, 32'h41c6c654, 32'h42c4e8c3, 32'h42148b1f};
test_output[9795] = '{32'h42c4e8c3};
test_index[9795] = '{6};
test_input[78368:78375] = '{32'hc25252a1, 32'hc25e19f6, 32'h42197164, 32'h41ba8a88, 32'hc25bf2f9, 32'hc2991ed3, 32'h3ea6e8cf, 32'h425c8535};
test_output[9796] = '{32'h425c8535};
test_index[9796] = '{7};
test_input[78376:78383] = '{32'h40c17297, 32'h421adc93, 32'hc2ba8fa5, 32'hc29607a6, 32'h41f0afc6, 32'h41095ee4, 32'h411c645f, 32'hc261b84d};
test_output[9797] = '{32'h421adc93};
test_index[9797] = '{1};
test_input[78384:78391] = '{32'h3f325906, 32'hc2c56ef2, 32'hc22ea094, 32'h42722a6a, 32'hc2b3de04, 32'h41a11f87, 32'h4196a4a0, 32'h4205f9a8};
test_output[9798] = '{32'h42722a6a};
test_index[9798] = '{3};
test_input[78392:78399] = '{32'hc2af6c10, 32'h429b1a6f, 32'hc22df1b5, 32'h426fa2e0, 32'hc251088e, 32'h420fbaab, 32'h420715ac, 32'h42a995c5};
test_output[9799] = '{32'h42a995c5};
test_index[9799] = '{7};
test_input[78400:78407] = '{32'hc2bc8b52, 32'hc2b980f4, 32'h42468229, 32'hc140eaf9, 32'h428ec889, 32'hc20c8c89, 32'hc2b889e0, 32'hc28992c8};
test_output[9800] = '{32'h428ec889};
test_index[9800] = '{4};
test_input[78408:78415] = '{32'h41544bc2, 32'hc24a7b81, 32'h4297f356, 32'hc2b15378, 32'hc2c14b8e, 32'hc2038d28, 32'h42bda00e, 32'h424a3faf};
test_output[9801] = '{32'h42bda00e};
test_index[9801] = '{6};
test_input[78416:78423] = '{32'h42422d19, 32'hc19627a2, 32'h426bfe02, 32'hc2c16e89, 32'h41abfdad, 32'hc288a383, 32'h422488f5, 32'h4261aa72};
test_output[9802] = '{32'h426bfe02};
test_index[9802] = '{2};
test_input[78424:78431] = '{32'hc2b9b5ab, 32'hc2599f4d, 32'h42c76d3b, 32'hc290182d, 32'h42bc4437, 32'hc27db3aa, 32'hc2174154, 32'hc19cc2d4};
test_output[9803] = '{32'h42c76d3b};
test_index[9803] = '{2};
test_input[78432:78439] = '{32'hc1d2175b, 32'hc2871cb5, 32'h42350d7f, 32'hc2c36af5, 32'hc1f3603a, 32'hc2acb0ea, 32'h421318b8, 32'h421339b5};
test_output[9804] = '{32'h42350d7f};
test_index[9804] = '{2};
test_input[78440:78447] = '{32'hc1a840cc, 32'hc2b3daff, 32'h42893902, 32'h4200db26, 32'h42a6f2af, 32'h41e5a2e9, 32'hc2923b44, 32'h427db97d};
test_output[9805] = '{32'h42a6f2af};
test_index[9805] = '{4};
test_input[78448:78455] = '{32'hc2a60437, 32'hc2932218, 32'h42a11150, 32'hc23eedd8, 32'hc287e46d, 32'hc1c6fc3a, 32'hc169b592, 32'h40447004};
test_output[9806] = '{32'h42a11150};
test_index[9806] = '{2};
test_input[78456:78463] = '{32'hc2485276, 32'hc2555210, 32'h42b23582, 32'hc2361425, 32'hc2212dbb, 32'hc1866339, 32'h42267834, 32'h42c1777b};
test_output[9807] = '{32'h42c1777b};
test_index[9807] = '{7};
test_input[78464:78471] = '{32'h42b5e9fc, 32'h412109da, 32'h40b8e2cf, 32'h42039f4f, 32'h42a32f84, 32'hc2a5d907, 32'h42387928, 32'hc292c466};
test_output[9808] = '{32'h42b5e9fc};
test_index[9808] = '{0};
test_input[78472:78479] = '{32'hc1e29452, 32'h426ffd04, 32'h42948cda, 32'h41ce40ff, 32'h41839f3f, 32'h41b1eb83, 32'hc205d767, 32'h4241e2f4};
test_output[9809] = '{32'h42948cda};
test_index[9809] = '{2};
test_input[78480:78487] = '{32'hbfeaa587, 32'hc280584d, 32'h424ada0b, 32'h42aa16d1, 32'hc0c11bc1, 32'hc22170fa, 32'h40c3e66c, 32'h42b6ac13};
test_output[9810] = '{32'h42b6ac13};
test_index[9810] = '{7};
test_input[78488:78495] = '{32'hc2020863, 32'h411f485b, 32'h424fe3ac, 32'hc23f142c, 32'h42820684, 32'h42212cc1, 32'hc1fc15aa, 32'hc27d6538};
test_output[9811] = '{32'h42820684};
test_index[9811] = '{4};
test_input[78496:78503] = '{32'hc28075cf, 32'hc2c4390b, 32'hc24b4779, 32'h424808c1, 32'hc234484f, 32'hc2a837ca, 32'h42643628, 32'h424c53e7};
test_output[9812] = '{32'h42643628};
test_index[9812] = '{6};
test_input[78504:78511] = '{32'hc1b9492e, 32'h417197a0, 32'hc23f48ef, 32'h41cd11c4, 32'h42256450, 32'h4229513f, 32'h421c37b5, 32'hc2b63aaa};
test_output[9813] = '{32'h4229513f};
test_index[9813] = '{5};
test_input[78512:78519] = '{32'hbf631dac, 32'hc2844d78, 32'h42873a27, 32'h41f1693e, 32'hc1da6bcd, 32'hc20569cf, 32'h42b22f21, 32'hc21c6202};
test_output[9814] = '{32'h42b22f21};
test_index[9814] = '{6};
test_input[78520:78527] = '{32'h42b3d9cf, 32'h42c1c81f, 32'h42c5b85b, 32'hc15f6944, 32'h4236c623, 32'h41a496f1, 32'h412cb6ca, 32'hc2c6197b};
test_output[9815] = '{32'h42c5b85b};
test_index[9815] = '{2};
test_input[78528:78535] = '{32'hc2a43ae2, 32'hc2023c83, 32'h41ea1925, 32'hc1d93391, 32'h4299a0a7, 32'hc132c35b, 32'h429a0fe5, 32'hc1445297};
test_output[9816] = '{32'h429a0fe5};
test_index[9816] = '{6};
test_input[78536:78543] = '{32'hc2330b21, 32'h42a5c105, 32'h428b794a, 32'hc1e5a957, 32'h424c9ace, 32'h42b58634, 32'hc1d667b8, 32'h423b6da8};
test_output[9817] = '{32'h42b58634};
test_index[9817] = '{5};
test_input[78544:78551] = '{32'h41924510, 32'hc25f88e1, 32'hc2844d17, 32'hc2bf1d02, 32'h42ab28e1, 32'h42643b03, 32'hc1ddbf1a, 32'hc29a0f0d};
test_output[9818] = '{32'h42ab28e1};
test_index[9818] = '{4};
test_input[78552:78559] = '{32'hc2be85bc, 32'h40d04b22, 32'hc2c159d5, 32'hc111d9b3, 32'h429e4530, 32'hc29b673e, 32'h429df97e, 32'h42053c6a};
test_output[9819] = '{32'h429e4530};
test_index[9819] = '{4};
test_input[78560:78567] = '{32'hc2bbf712, 32'h42b30009, 32'h4285e349, 32'hc1ce3a82, 32'h41d863ab, 32'h40ae7455, 32'h42953659, 32'hc1943efc};
test_output[9820] = '{32'h42b30009};
test_index[9820] = '{1};
test_input[78568:78575] = '{32'h41c2c41b, 32'h42c4c4cc, 32'h41a6b25b, 32'hc23075f3, 32'hc293a2ee, 32'hc2a6a6df, 32'h4223f4a6, 32'hc1ba7266};
test_output[9821] = '{32'h42c4c4cc};
test_index[9821] = '{1};
test_input[78576:78583] = '{32'hc2ab9eb3, 32'hc0928841, 32'hc2b84d85, 32'hc2aa40dd, 32'hc2bd9075, 32'hc137105f, 32'hc297c6e1, 32'h41d83adb};
test_output[9822] = '{32'h41d83adb};
test_index[9822] = '{7};
test_input[78584:78591] = '{32'hc2a88e76, 32'hc2a343b2, 32'hc2abddb8, 32'hc1949ecb, 32'hc280671e, 32'h42ac3777, 32'h423f45ca, 32'h42b7d88c};
test_output[9823] = '{32'h42b7d88c};
test_index[9823] = '{7};
test_input[78592:78599] = '{32'hc21ac0a4, 32'h3e509425, 32'h4179c0e5, 32'hc29052a0, 32'hc1982b2c, 32'hc21a9c2c, 32'h40921d35, 32'h4268768c};
test_output[9824] = '{32'h4268768c};
test_index[9824] = '{7};
test_input[78600:78607] = '{32'h42825a30, 32'h41dc10e2, 32'h4221d8be, 32'h41fc40af, 32'h4222b1ad, 32'hc24a89f9, 32'hc1c30d44, 32'hc2b176c9};
test_output[9825] = '{32'h42825a30};
test_index[9825] = '{0};
test_input[78608:78615] = '{32'hc295d754, 32'h4133bbec, 32'hc17e6438, 32'h41df65b7, 32'hbf8a28aa, 32'h41fce4d5, 32'hc269e921, 32'h425b0bf9};
test_output[9826] = '{32'h425b0bf9};
test_index[9826] = '{7};
test_input[78616:78623] = '{32'h42b0cae1, 32'hc0b149b4, 32'h426fc529, 32'h42a99d07, 32'hc2b0feb5, 32'hc2c408cb, 32'h4197847e, 32'hc28da306};
test_output[9827] = '{32'h42b0cae1};
test_index[9827] = '{0};
test_input[78624:78631] = '{32'h41f5a7d1, 32'hc22995a4, 32'h41bbf23d, 32'hc2a0b040, 32'h4285d533, 32'hc1392d95, 32'h420b9e4e, 32'h42b4c8d6};
test_output[9828] = '{32'h42b4c8d6};
test_index[9828] = '{7};
test_input[78632:78639] = '{32'hc24cc27e, 32'hc2babc23, 32'h41d471d7, 32'h423ed009, 32'h42ba8c6c, 32'hc2aca9ae, 32'hc28237d2, 32'hc2885afb};
test_output[9829] = '{32'h42ba8c6c};
test_index[9829] = '{4};
test_input[78640:78647] = '{32'h4286ac44, 32'hc2004753, 32'hc235f339, 32'h42b6429c, 32'hc26418a9, 32'hc066e583, 32'hc2a7a912, 32'h4287c7d7};
test_output[9830] = '{32'h42b6429c};
test_index[9830] = '{3};
test_input[78648:78655] = '{32'h4226f565, 32'hc097f937, 32'hc28ebfc0, 32'hc2949b8c, 32'hc08976fd, 32'hc285e412, 32'h4247e08f, 32'h42bd5672};
test_output[9831] = '{32'h42bd5672};
test_index[9831] = '{7};
test_input[78656:78663] = '{32'hc25de7a3, 32'hc0d0ccb8, 32'hc293b604, 32'hc2ae6087, 32'h425ea002, 32'h420b6e79, 32'h41e6353d, 32'h425a3326};
test_output[9832] = '{32'h425ea002};
test_index[9832] = '{4};
test_input[78664:78671] = '{32'h42be6469, 32'hc201ed72, 32'hc19979b9, 32'h429dd85c, 32'h427aca0c, 32'hc2982db2, 32'h42c0bdf8, 32'hc1bd7aa6};
test_output[9833] = '{32'h42c0bdf8};
test_index[9833] = '{6};
test_input[78672:78679] = '{32'h411fc96e, 32'h41ebf9ee, 32'hc1f322f4, 32'hc230dc6a, 32'h42212d75, 32'h424bee44, 32'hc1ebae52, 32'hc1c5305a};
test_output[9834] = '{32'h424bee44};
test_index[9834] = '{5};
test_input[78680:78687] = '{32'h42a64eae, 32'hc26b8622, 32'hc291dbec, 32'hc282b85e, 32'h4296e069, 32'h425e66de, 32'h41fee3e6, 32'h42bf92ee};
test_output[9835] = '{32'h42bf92ee};
test_index[9835] = '{7};
test_input[78688:78695] = '{32'hc0e651aa, 32'h4218b0ae, 32'h41c4a509, 32'h42c55892, 32'hc23b4934, 32'hc14ae807, 32'hc29a6de3, 32'h42716137};
test_output[9836] = '{32'h42c55892};
test_index[9836] = '{3};
test_input[78696:78703] = '{32'h42a2a19f, 32'hc2a70ba6, 32'hc22fcd4b, 32'h423b0d43, 32'h40c1141a, 32'hc297488b, 32'hc1fc922e, 32'h42b1ef0d};
test_output[9837] = '{32'h42b1ef0d};
test_index[9837] = '{7};
test_input[78704:78711] = '{32'hc29dbff1, 32'h4294739a, 32'h41d80729, 32'h4294032b, 32'h4136c363, 32'h416b50d9, 32'hc227034a, 32'h4286edab};
test_output[9838] = '{32'h4294739a};
test_index[9838] = '{1};
test_input[78712:78719] = '{32'hc2c2d8b2, 32'h4295681e, 32'h42bdc2d7, 32'hc153f20a, 32'h40e0a7dd, 32'hc2773d1f, 32'h42be87db, 32'hc2611e2b};
test_output[9839] = '{32'h42be87db};
test_index[9839] = '{6};
test_input[78720:78727] = '{32'hc1974ad8, 32'h428341ed, 32'hc21eee01, 32'h421870b7, 32'h4241a425, 32'hc16a76f4, 32'hc2a136fb, 32'h42ba27e0};
test_output[9840] = '{32'h42ba27e0};
test_index[9840] = '{7};
test_input[78728:78735] = '{32'h42c02384, 32'h40e343b2, 32'hc27267a7, 32'hc24639d0, 32'h4263d177, 32'hc24f9850, 32'h423ef61d, 32'hc19697f4};
test_output[9841] = '{32'h42c02384};
test_index[9841] = '{0};
test_input[78736:78743] = '{32'h42a73a2f, 32'hc26daa30, 32'hc2234960, 32'hc10c990a, 32'h41b9aa90, 32'h419ca32d, 32'hc215fc40, 32'hc1005c0a};
test_output[9842] = '{32'h42a73a2f};
test_index[9842] = '{0};
test_input[78744:78751] = '{32'h41ae8364, 32'h4282879a, 32'h42ad1b56, 32'hc2afdb56, 32'hc2c1eda3, 32'hc13b8392, 32'h42a45ed5, 32'h41f44f77};
test_output[9843] = '{32'h42ad1b56};
test_index[9843] = '{2};
test_input[78752:78759] = '{32'hc264aaf7, 32'hc1321e81, 32'hc1875d7a, 32'h42184613, 32'h41b196e8, 32'hc2259937, 32'h4217d11b, 32'h418ae838};
test_output[9844] = '{32'h42184613};
test_index[9844] = '{3};
test_input[78760:78767] = '{32'hc10ab5fc, 32'h42800211, 32'h423d37d4, 32'hc2a8794e, 32'hc1d347f6, 32'hc259c3f0, 32'hc1ef2b70, 32'hc2ad9a97};
test_output[9845] = '{32'h42800211};
test_index[9845] = '{1};
test_input[78768:78775] = '{32'hc28ff3ea, 32'hc164b077, 32'h41376d11, 32'h41acd766, 32'h4298f64c, 32'h41f51f9c, 32'h42be9d7e, 32'hc2381af7};
test_output[9846] = '{32'h42be9d7e};
test_index[9846] = '{6};
test_input[78776:78783] = '{32'h42b5231b, 32'h429a5230, 32'h42935657, 32'h41ebf872, 32'h422ad2d8, 32'hc29d8462, 32'h42bc28f1, 32'hc2885cb5};
test_output[9847] = '{32'h42bc28f1};
test_index[9847] = '{6};
test_input[78784:78791] = '{32'h41be30c9, 32'hc1fe582c, 32'h42b9f3b5, 32'hc20c80cc, 32'hc261db0b, 32'h4269f4d9, 32'hc294da46, 32'h41e456ac};
test_output[9848] = '{32'h42b9f3b5};
test_index[9848] = '{2};
test_input[78792:78799] = '{32'hc2a5ec6f, 32'h41bdd7ee, 32'hc2342454, 32'h405627a2, 32'hc2653da8, 32'hbfa60221, 32'h42a4b274, 32'hc2ae15c1};
test_output[9849] = '{32'h42a4b274};
test_index[9849] = '{6};
test_input[78800:78807] = '{32'h42aeb314, 32'h42bfd66b, 32'h4223b5cc, 32'h40d691e0, 32'h429d3d40, 32'hc1088103, 32'h42005ddc, 32'hc150a608};
test_output[9850] = '{32'h42bfd66b};
test_index[9850] = '{1};
test_input[78808:78815] = '{32'hc2952707, 32'hc2c18adc, 32'h3e25d5ee, 32'h4299ef6a, 32'h4160a124, 32'hc1c02ff0, 32'h420094ca, 32'h4202fe92};
test_output[9851] = '{32'h4299ef6a};
test_index[9851] = '{3};
test_input[78816:78823] = '{32'h42bfe80d, 32'hc2a52a3a, 32'hc2b0f995, 32'h41e18ffb, 32'h425fa086, 32'h42497664, 32'h41e3f3e0, 32'hc1bc533e};
test_output[9852] = '{32'h42bfe80d};
test_index[9852] = '{0};
test_input[78824:78831] = '{32'h4237e1e1, 32'hc28f84e1, 32'h4131be12, 32'h422860c7, 32'h4296c46a, 32'h411395b1, 32'hc2c0a20e, 32'h4257d812};
test_output[9853] = '{32'h4296c46a};
test_index[9853] = '{4};
test_input[78832:78839] = '{32'hc0c13616, 32'hc28f3d2e, 32'h429cbe76, 32'hc208c23e, 32'h428547a1, 32'hc132e99b, 32'h41ea8eee, 32'h421120ac};
test_output[9854] = '{32'h429cbe76};
test_index[9854] = '{2};
test_input[78840:78847] = '{32'h42b86353, 32'h4291d3c6, 32'hc2b8d7c8, 32'h421f0261, 32'h426442d6, 32'h411f30b2, 32'hc291e177, 32'h42be47d6};
test_output[9855] = '{32'h42be47d6};
test_index[9855] = '{7};
test_input[78848:78855] = '{32'h41df5b53, 32'h428a99a8, 32'h42aaa17f, 32'hc13d097e, 32'h41c13462, 32'h42806f85, 32'hc2b4cdc5, 32'h42aba23f};
test_output[9856] = '{32'h42aba23f};
test_index[9856] = '{7};
test_input[78856:78863] = '{32'h428b6e13, 32'h4259fde0, 32'h42914b79, 32'hc26fdaba, 32'hc231e33f, 32'hc1b6efaa, 32'h41ab1599, 32'hc1a1b2be};
test_output[9857] = '{32'h42914b79};
test_index[9857] = '{2};
test_input[78864:78871] = '{32'hc28c290a, 32'hc21bed85, 32'hc2bbd35f, 32'h41fe1433, 32'hc26b35c4, 32'hc1cf8b81, 32'hc27b2f73, 32'hc20dfde0};
test_output[9858] = '{32'h41fe1433};
test_index[9858] = '{3};
test_input[78872:78879] = '{32'hc15ea262, 32'h4243cac1, 32'hc1cb8efb, 32'h428439f4, 32'hc267f740, 32'h422fe0e8, 32'h4280cabe, 32'hc246af88};
test_output[9859] = '{32'h428439f4};
test_index[9859] = '{3};
test_input[78880:78887] = '{32'h42c566e1, 32'h42b497bd, 32'hc28278ca, 32'hc27ec3d1, 32'h42709956, 32'h42c3ac6b, 32'h427298de, 32'hc1e5bd16};
test_output[9860] = '{32'h42c566e1};
test_index[9860] = '{0};
test_input[78888:78895] = '{32'h41965018, 32'hc2413f91, 32'h429589f0, 32'h41d1e1e4, 32'h428df9ba, 32'h422e14d9, 32'h4106f530, 32'hc22acabd};
test_output[9861] = '{32'h429589f0};
test_index[9861] = '{2};
test_input[78896:78903] = '{32'h42a9f7ce, 32'h420f33d5, 32'h42b5973e, 32'hc2a0ad71, 32'hc2b235bd, 32'h420437af, 32'hc1a48b4a, 32'h4274f45b};
test_output[9862] = '{32'h42b5973e};
test_index[9862] = '{2};
test_input[78904:78911] = '{32'hc2c03edb, 32'h40a73300, 32'hc2c279b0, 32'hc21c0cf9, 32'hc292cc0b, 32'h41cb02b4, 32'h40bb5a00, 32'hc28c0ed8};
test_output[9863] = '{32'h41cb02b4};
test_index[9863] = '{5};
test_input[78912:78919] = '{32'hc2b4539b, 32'hc266705d, 32'hc2bbd673, 32'hc0a469c1, 32'hc143ac56, 32'hc0f8205e, 32'h4285e225, 32'hc2a0fc04};
test_output[9864] = '{32'h4285e225};
test_index[9864] = '{6};
test_input[78920:78927] = '{32'hc29c4f0a, 32'h42b227b4, 32'hc267fa82, 32'hc12fde6c, 32'hc16bf9a9, 32'hc2767965, 32'hc282956e, 32'hc2394dc6};
test_output[9865] = '{32'h42b227b4};
test_index[9865] = '{1};
test_input[78928:78935] = '{32'hc1034ebe, 32'hc290e890, 32'hc288809a, 32'hc1bda524, 32'h40e011a9, 32'hc23700f7, 32'h42aba76f, 32'h42b82731};
test_output[9866] = '{32'h42b82731};
test_index[9866] = '{7};
test_input[78936:78943] = '{32'hc28719fb, 32'h42c50f34, 32'hc2583a75, 32'hc14cb375, 32'h41abf7d0, 32'hc0170cda, 32'h425737bf, 32'hc0dbb092};
test_output[9867] = '{32'h42c50f34};
test_index[9867] = '{1};
test_input[78944:78951] = '{32'h42b445d4, 32'hc23928ca, 32'hc185cb3d, 32'hc0c853e6, 32'h42726b6e, 32'h419a88ea, 32'h425392d0, 32'h42000e40};
test_output[9868] = '{32'h42b445d4};
test_index[9868] = '{0};
test_input[78952:78959] = '{32'h41fec7f4, 32'hc0470aa8, 32'h4258402d, 32'h42b916f7, 32'hc267ba91, 32'h4288f175, 32'h42a8c1de, 32'hc2c6e98a};
test_output[9869] = '{32'h42b916f7};
test_index[9869] = '{3};
test_input[78960:78967] = '{32'h41d78a89, 32'h42262680, 32'hc1de188e, 32'hc2611c31, 32'h42af4322, 32'hc17b0684, 32'hc1cee151, 32'hc0f4f372};
test_output[9870] = '{32'h42af4322};
test_index[9870] = '{4};
test_input[78968:78975] = '{32'h41e3f5ff, 32'h42b8d18d, 32'hc215804a, 32'hc2c6c37b, 32'hc2850251, 32'hc27aed84, 32'hc13b663e, 32'h42b63993};
test_output[9871] = '{32'h42b8d18d};
test_index[9871] = '{1};
test_input[78976:78983] = '{32'h424b36d2, 32'hc281dbe9, 32'h42294083, 32'hc170e298, 32'hc2c5f30a, 32'hc11a1b16, 32'hc28c4ade, 32'hc26de298};
test_output[9872] = '{32'h424b36d2};
test_index[9872] = '{0};
test_input[78984:78991] = '{32'h4029f9d1, 32'h425f9b25, 32'h428620eb, 32'hbf2d8c15, 32'hc230e359, 32'h4209c2c1, 32'h41c3aa8b, 32'h4108552c};
test_output[9873] = '{32'h428620eb};
test_index[9873] = '{2};
test_input[78992:78999] = '{32'hc2b63059, 32'hc291b896, 32'h4184316b, 32'h42929c9e, 32'h4225af3f, 32'h42885072, 32'hc286ad66, 32'h4204c5b8};
test_output[9874] = '{32'h42929c9e};
test_index[9874] = '{3};
test_input[79000:79007] = '{32'hc2bc9f3b, 32'h429010a2, 32'h42ab5354, 32'h425f5909, 32'h42095d8e, 32'hc2c0955b, 32'h422d4e87, 32'h4299841b};
test_output[9875] = '{32'h42ab5354};
test_index[9875] = '{2};
test_input[79008:79015] = '{32'hc25f8973, 32'hc2221a45, 32'hc2c176f7, 32'h4256a861, 32'hc136c74e, 32'h409cb0eb, 32'h42123b7f, 32'h429b777a};
test_output[9876] = '{32'h429b777a};
test_index[9876] = '{7};
test_input[79016:79023] = '{32'h42b58b9d, 32'h423bfe93, 32'h426dc602, 32'hc24639a6, 32'h42b14c8b, 32'h42772084, 32'h4214d5c8, 32'h4284b651};
test_output[9877] = '{32'h42b58b9d};
test_index[9877] = '{0};
test_input[79024:79031] = '{32'h422101a1, 32'hc01e06a3, 32'h42b3f27c, 32'hc1b02842, 32'hc0ba00b6, 32'h41efdc28, 32'h423a6212, 32'hc17c02c9};
test_output[9878] = '{32'h42b3f27c};
test_index[9878] = '{2};
test_input[79032:79039] = '{32'h42a42eb8, 32'hc20e4ffa, 32'hc2b01a49, 32'hc1930aaa, 32'h4178b687, 32'hc1778fc5, 32'h425169c4, 32'hc25c13e3};
test_output[9879] = '{32'h42a42eb8};
test_index[9879] = '{0};
test_input[79040:79047] = '{32'hc00ea0d6, 32'hc11b2e71, 32'hc2af608d, 32'hc2b9c460, 32'hc2871f27, 32'hc04d4e31, 32'h42a98bd6, 32'hc2778ce3};
test_output[9880] = '{32'h42a98bd6};
test_index[9880] = '{6};
test_input[79048:79055] = '{32'hc28861c6, 32'h42c3de24, 32'h41990cb5, 32'hc25e332c, 32'h4264ee46, 32'h42c6ed59, 32'h428ba6f4, 32'hc2761f18};
test_output[9881] = '{32'h42c6ed59};
test_index[9881] = '{5};
test_input[79056:79063] = '{32'hc156aa33, 32'h420571f7, 32'hc29a738c, 32'hc1dcb877, 32'h418f897d, 32'h42bc3f43, 32'h42318ccf, 32'hbfb54898};
test_output[9882] = '{32'h42bc3f43};
test_index[9882] = '{5};
test_input[79064:79071] = '{32'h421ab39b, 32'h42b64799, 32'hc0b7012c, 32'h41734dd7, 32'hc29ec08a, 32'hc2c67e4f, 32'hc2500009, 32'hc1fe3684};
test_output[9883] = '{32'h42b64799};
test_index[9883] = '{1};
test_input[79072:79079] = '{32'h41e27314, 32'hc23c0b41, 32'h41513e97, 32'h429c823a, 32'hc2195a7d, 32'hc2c640d1, 32'h42c476b7, 32'h42651b14};
test_output[9884] = '{32'h42c476b7};
test_index[9884] = '{6};
test_input[79080:79087] = '{32'hc278a467, 32'hc26c2d1a, 32'hc217515f, 32'h4030d847, 32'hc29fde15, 32'h425bdc83, 32'hc1043f8e, 32'h42640adb};
test_output[9885] = '{32'h42640adb};
test_index[9885] = '{7};
test_input[79088:79095] = '{32'h40b7f746, 32'h424d9cbf, 32'hc2c58397, 32'h429cf803, 32'h42bdd583, 32'h41fc66bf, 32'hbf4f5976, 32'h42629dde};
test_output[9886] = '{32'h42bdd583};
test_index[9886] = '{4};
test_input[79096:79103] = '{32'h427ea59f, 32'h41898eb9, 32'hc2293a54, 32'hc225c1e7, 32'hc2a9c84a, 32'hc2861aca, 32'h42891fb7, 32'h4284fede};
test_output[9887] = '{32'h42891fb7};
test_index[9887] = '{6};
test_input[79104:79111] = '{32'h42b7667a, 32'hc05acbab, 32'h429eb8e4, 32'hc255e733, 32'hc1545701, 32'hc27ec924, 32'h42528120, 32'hc18f2180};
test_output[9888] = '{32'h42b7667a};
test_index[9888] = '{0};
test_input[79112:79119] = '{32'h3ea2630d, 32'h42767da8, 32'h41f4e0bd, 32'h42aea9bf, 32'h42a271d9, 32'hc1da22de, 32'hc231b3d0, 32'hc2a61c45};
test_output[9889] = '{32'h42aea9bf};
test_index[9889] = '{3};
test_input[79120:79127] = '{32'h42a0e9f4, 32'h3fd8e320, 32'h428b6626, 32'hc19d245b, 32'h41cb409f, 32'hc1739196, 32'h42449e9a, 32'hc2122c50};
test_output[9890] = '{32'h42a0e9f4};
test_index[9890] = '{0};
test_input[79128:79135] = '{32'hc26ffedd, 32'hc0b5e94c, 32'h426b162e, 32'hc203f474, 32'hc2c666a2, 32'hc285e6a8, 32'h421a611b, 32'hc22a2108};
test_output[9891] = '{32'h426b162e};
test_index[9891] = '{2};
test_input[79136:79143] = '{32'hc1b5f4ca, 32'h421855db, 32'hc2857058, 32'h41dee5cc, 32'h4265a10e, 32'hc2842cb2, 32'h429e5ac3, 32'h42721960};
test_output[9892] = '{32'h429e5ac3};
test_index[9892] = '{6};
test_input[79144:79151] = '{32'hc20834c2, 32'h429dcbf1, 32'h4281d008, 32'h41cde6fc, 32'h42ba9c09, 32'hc2745db4, 32'hc233f5c1, 32'h423073bf};
test_output[9893] = '{32'h42ba9c09};
test_index[9893] = '{4};
test_input[79152:79159] = '{32'hc2a10047, 32'hc280b9de, 32'hc19c7713, 32'hc028d823, 32'h427d0d0f, 32'h424b969c, 32'h4228beca, 32'hc199c760};
test_output[9894] = '{32'h427d0d0f};
test_index[9894] = '{4};
test_input[79160:79167] = '{32'hc13f938a, 32'hc2a5665a, 32'h426a855a, 32'h42751cc7, 32'h42c324c5, 32'hc2af5742, 32'hc291c1c0, 32'h4191e99a};
test_output[9895] = '{32'h42c324c5};
test_index[9895] = '{4};
test_input[79168:79175] = '{32'hc2558b2d, 32'hc2b5dd23, 32'hc26a6186, 32'h42b2c871, 32'hc217d213, 32'h42983766, 32'h420e4e94, 32'h3ed0e617};
test_output[9896] = '{32'h42b2c871};
test_index[9896] = '{3};
test_input[79176:79183] = '{32'h42ab3368, 32'hc2ac5bdd, 32'hc232abbf, 32'hc1c27fdc, 32'hc04be68d, 32'hc1e15715, 32'hc28eaee2, 32'hc12da67b};
test_output[9897] = '{32'h42ab3368};
test_index[9897] = '{0};
test_input[79184:79191] = '{32'hc270c119, 32'h4270ba4f, 32'h42a95aad, 32'h42c3aace, 32'hc17f0ea6, 32'h41d639e0, 32'h41fe7f14, 32'h42c1e3a2};
test_output[9898] = '{32'h42c3aace};
test_index[9898] = '{3};
test_input[79192:79199] = '{32'h4198094c, 32'hc16bb379, 32'h42b3dc28, 32'hc2131b7e, 32'h42aec2ba, 32'h42877781, 32'hc2a23ca7, 32'h41cf2601};
test_output[9899] = '{32'h42b3dc28};
test_index[9899] = '{2};
test_input[79200:79207] = '{32'h424919a4, 32'h416435e0, 32'h42abbee8, 32'h40e094a9, 32'hc2204a5c, 32'h42696dc2, 32'h4251b77b, 32'hc27e7a7e};
test_output[9900] = '{32'h42abbee8};
test_index[9900] = '{2};
test_input[79208:79215] = '{32'h42c11b1e, 32'h426e651f, 32'h42b1a4cf, 32'h40a783e7, 32'hc2894d8f, 32'hc2bc9fc7, 32'hc1ad67e6, 32'h4293f433};
test_output[9901] = '{32'h42c11b1e};
test_index[9901] = '{0};
test_input[79216:79223] = '{32'hc2c47b96, 32'h40796179, 32'h4218cc76, 32'h42c63aaa, 32'h423113bc, 32'hc102c8c0, 32'h4288c16b, 32'hc2b95a31};
test_output[9902] = '{32'h42c63aaa};
test_index[9902] = '{3};
test_input[79224:79231] = '{32'hc22d1a45, 32'hc215f306, 32'hc1e7d8dc, 32'h407f2b3c, 32'h418bbaff, 32'hc21e4c8a, 32'h4266412f, 32'hc2be4dcc};
test_output[9903] = '{32'h4266412f};
test_index[9903] = '{6};
test_input[79232:79239] = '{32'h42bd12b7, 32'hc1466e6b, 32'hc24e7214, 32'h41fd80a9, 32'h4159bd6c, 32'h42c6df6c, 32'h4281cede, 32'h427cfaf1};
test_output[9904] = '{32'h42c6df6c};
test_index[9904] = '{5};
test_input[79240:79247] = '{32'h41132d16, 32'h428fd18d, 32'h42aaa38c, 32'hc25e798e, 32'h423a0118, 32'h429da431, 32'hc2286be8, 32'hc24eb8f4};
test_output[9905] = '{32'h42aaa38c};
test_index[9905] = '{2};
test_input[79248:79255] = '{32'hc20a1d3d, 32'hc2545f92, 32'hc14e96ad, 32'hc14b7661, 32'h40ebc885, 32'h4206db1e, 32'h42058233, 32'hc219f512};
test_output[9906] = '{32'h4206db1e};
test_index[9906] = '{5};
test_input[79256:79263] = '{32'h4192675d, 32'h41df91f2, 32'hc19a46b3, 32'hc24bc872, 32'h41d3869b, 32'h42a6eb3b, 32'hbe924c9f, 32'hc2ac34f5};
test_output[9907] = '{32'h42a6eb3b};
test_index[9907] = '{5};
test_input[79264:79271] = '{32'h4173f90e, 32'h42bb5319, 32'hc2a8096c, 32'hc24e4655, 32'hc21f6a1e, 32'hc2428bd8, 32'hc260cbc0, 32'hc1077dec};
test_output[9908] = '{32'h42bb5319};
test_index[9908] = '{1};
test_input[79272:79279] = '{32'h41e6aa90, 32'hc287f541, 32'h428751ea, 32'h4212ea81, 32'h429f4ae3, 32'hc292e27b, 32'hc2396160, 32'hc0e73104};
test_output[9909] = '{32'h429f4ae3};
test_index[9909] = '{4};
test_input[79280:79287] = '{32'h42584dd2, 32'hc1b4401e, 32'h419b0330, 32'h42acc634, 32'hc2804d56, 32'hc102fb80, 32'hc22530a3, 32'h426b2311};
test_output[9910] = '{32'h42acc634};
test_index[9910] = '{3};
test_input[79288:79295] = '{32'h41dd287a, 32'h41809f14, 32'hc276791d, 32'h41e7663e, 32'h4270204b, 32'hc2131aa5, 32'h42bb6438, 32'h41bea10e};
test_output[9911] = '{32'h42bb6438};
test_index[9911] = '{6};
test_input[79296:79303] = '{32'hc23e92bf, 32'h424bb23d, 32'h4289f785, 32'hc1d87108, 32'h42b63647, 32'hc12e0e39, 32'h423613a6, 32'h4285ad8a};
test_output[9912] = '{32'h42b63647};
test_index[9912] = '{4};
test_input[79304:79311] = '{32'h42a72740, 32'h40c0e620, 32'h42121a05, 32'hc04005ce, 32'h419f3e5d, 32'h41c4fd64, 32'hc1d1d182, 32'hc0a996cf};
test_output[9913] = '{32'h42a72740};
test_index[9913] = '{0};
test_input[79312:79319] = '{32'h428c99ed, 32'hc292d475, 32'h42a1ac37, 32'hc2912035, 32'hc1cde241, 32'hc20b3487, 32'h42b028d9, 32'hc1855ea2};
test_output[9914] = '{32'h42b028d9};
test_index[9914] = '{6};
test_input[79320:79327] = '{32'h424051f5, 32'h429c576c, 32'h42be8f97, 32'h4290c8c7, 32'h42c5caf8, 32'h42691cca, 32'hc1b280a0, 32'h42782b10};
test_output[9915] = '{32'h42c5caf8};
test_index[9915] = '{4};
test_input[79328:79335] = '{32'hc2bcaeab, 32'h429e2d8d, 32'h42bcede8, 32'h4214c8ff, 32'hc29de1e7, 32'hc2bd2803, 32'h41e8aacb, 32'hc2a1e614};
test_output[9916] = '{32'h42bcede8};
test_index[9916] = '{2};
test_input[79336:79343] = '{32'h4164bb10, 32'hc1d34802, 32'h406057ae, 32'hc18f231c, 32'h425d4336, 32'h42725360, 32'h42a29b7e, 32'hc20e6440};
test_output[9917] = '{32'h42a29b7e};
test_index[9917] = '{6};
test_input[79344:79351] = '{32'hc2875f44, 32'h42581787, 32'h42c2b8ae, 32'h429b26a7, 32'hc20b1c74, 32'hc0a316e9, 32'h42b2c9df, 32'h424c47f4};
test_output[9918] = '{32'h42c2b8ae};
test_index[9918] = '{2};
test_input[79352:79359] = '{32'hc2712e7b, 32'h41dedeb5, 32'hc1f2c6bf, 32'hc22e83ff, 32'h4290fc67, 32'h41df61e0, 32'hc1ef77a3, 32'hc1e0c8e3};
test_output[9919] = '{32'h4290fc67};
test_index[9919] = '{4};
test_input[79360:79367] = '{32'hc29eae26, 32'h42bc3dbd, 32'hc23afc0e, 32'h41506d14, 32'hc039716f, 32'h42b7aa06, 32'hc032f309, 32'hc293c27c};
test_output[9920] = '{32'h42bc3dbd};
test_index[9920] = '{1};
test_input[79368:79375] = '{32'hc0d5121c, 32'hc231af1c, 32'hc2007be2, 32'hc28e5ba4, 32'h4243f20c, 32'hc264df94, 32'hc2bd63d0, 32'h40d8de7c};
test_output[9921] = '{32'h4243f20c};
test_index[9921] = '{4};
test_input[79376:79383] = '{32'h42898a68, 32'h41b4d649, 32'hbdc29e35, 32'hc2a652d0, 32'hc2b64592, 32'h429ae258, 32'hc29767c8, 32'h419ccab5};
test_output[9922] = '{32'h429ae258};
test_index[9922] = '{5};
test_input[79384:79391] = '{32'hc2c09107, 32'h41b5e268, 32'h41c01bed, 32'h42914391, 32'h41edf058, 32'hc1a8c4f8, 32'hc28c4fc9, 32'h42bf602e};
test_output[9923] = '{32'h42bf602e};
test_index[9923] = '{7};
test_input[79392:79399] = '{32'hc096bc64, 32'hc225848e, 32'hc20c6d2f, 32'hc14ba8a0, 32'h42984ba2, 32'hc245337c, 32'hbf6149ad, 32'h422cb8a1};
test_output[9924] = '{32'h42984ba2};
test_index[9924] = '{4};
test_input[79400:79407] = '{32'h4247b6b3, 32'hc2644861, 32'hc2c49112, 32'hc2af2df1, 32'h41799359, 32'h42ba8ef5, 32'hc1fd7408, 32'hc05a4cf2};
test_output[9925] = '{32'h42ba8ef5};
test_index[9925] = '{5};
test_input[79408:79415] = '{32'hc144ad32, 32'hc1afd8d5, 32'hc1ce124f, 32'hc08de2e3, 32'hc2902aaa, 32'h40b87570, 32'h421b563c, 32'hc1fdb486};
test_output[9926] = '{32'h421b563c};
test_index[9926] = '{6};
test_input[79416:79423] = '{32'h40d6b28f, 32'h42c69273, 32'hc180795e, 32'hc1ef073a, 32'hc0d9fbc7, 32'h41d5a6ed, 32'hc29f0081, 32'h427a5976};
test_output[9927] = '{32'h42c69273};
test_index[9927] = '{1};
test_input[79424:79431] = '{32'h424208c9, 32'h4255ae1c, 32'hc2aad5ba, 32'hc0ffd510, 32'h424f5889, 32'hc28ec18b, 32'h424bdee5, 32'hc1737b6f};
test_output[9928] = '{32'h4255ae1c};
test_index[9928] = '{1};
test_input[79432:79439] = '{32'hc254f518, 32'h413f57dc, 32'hc229e6b9, 32'hc2051470, 32'hc2c246e6, 32'h410da8ff, 32'hc2b8678e, 32'h42a5055f};
test_output[9929] = '{32'h42a5055f};
test_index[9929] = '{7};
test_input[79440:79447] = '{32'hc2aa436c, 32'hc292aabd, 32'h4212e011, 32'hc1ad308a, 32'h413d9c09, 32'hc2c5b7e7, 32'hc2980df5, 32'hc27f9b4b};
test_output[9930] = '{32'h4212e011};
test_index[9930] = '{2};
test_input[79448:79455] = '{32'h42129a8c, 32'h427e74da, 32'hc2017ac4, 32'h427becac, 32'h4043c74b, 32'h41e63f54, 32'h42c38857, 32'h426a958b};
test_output[9931] = '{32'h42c38857};
test_index[9931] = '{6};
test_input[79456:79463] = '{32'h429d2fbe, 32'hc2038425, 32'hc2be54a7, 32'h424daf7c, 32'hc2324931, 32'h42c60478, 32'h42b47f87, 32'h42a1401b};
test_output[9932] = '{32'h42c60478};
test_index[9932] = '{5};
test_input[79464:79471] = '{32'hc27647e9, 32'hc22325c7, 32'h41fab4f3, 32'hc249e432, 32'hc286de8d, 32'hc2a10e19, 32'hc260bdf4, 32'hc0c9ddf6};
test_output[9933] = '{32'h41fab4f3};
test_index[9933] = '{2};
test_input[79472:79479] = '{32'h427025c0, 32'hc23d999e, 32'hc233c908, 32'h414d5135, 32'hc082fac3, 32'h41c99278, 32'h42942104, 32'h421f358e};
test_output[9934] = '{32'h42942104};
test_index[9934] = '{6};
test_input[79480:79487] = '{32'h41290f3e, 32'h42824a59, 32'hc2956d81, 32'h42254ff2, 32'hc29d8fa5, 32'h42ace4a3, 32'h4296698a, 32'hc2853b31};
test_output[9935] = '{32'h42ace4a3};
test_index[9935] = '{5};
test_input[79488:79495] = '{32'h42118fcd, 32'h42924b9e, 32'h410bbfd1, 32'h420ba208, 32'h421f0b50, 32'hc21b92a1, 32'hc2a30aca, 32'hc09c3243};
test_output[9936] = '{32'h42924b9e};
test_index[9936] = '{1};
test_input[79496:79503] = '{32'h41e74294, 32'h42557173, 32'hc1611487, 32'hc06d0939, 32'hc2987672, 32'hc25f6847, 32'h4293acf8, 32'hc2825903};
test_output[9937] = '{32'h4293acf8};
test_index[9937] = '{6};
test_input[79504:79511] = '{32'hc28b6b1d, 32'hc225121b, 32'hc281ff01, 32'h4227db0b, 32'hc261f310, 32'hc2ab5402, 32'hc1ba88ee, 32'hc221ee81};
test_output[9938] = '{32'h4227db0b};
test_index[9938] = '{3};
test_input[79512:79519] = '{32'h41f94c55, 32'hc28ddba3, 32'h3f902da1, 32'h41c02c5e, 32'hc2be2f0e, 32'hc03e2ef6, 32'hc1d56d0c, 32'hc10d3350};
test_output[9939] = '{32'h41f94c55};
test_index[9939] = '{0};
test_input[79520:79527] = '{32'h4243ced3, 32'h429afd03, 32'h42456428, 32'hc2321db5, 32'hc2148396, 32'h42c1521f, 32'h42af0462, 32'hc28ddb47};
test_output[9940] = '{32'h42c1521f};
test_index[9940] = '{5};
test_input[79528:79535] = '{32'h42a7abb4, 32'h420424c6, 32'h42c3784a, 32'h429229ac, 32'h41d898c8, 32'h426af14c, 32'h4296cba1, 32'hc2b12fc9};
test_output[9941] = '{32'h42c3784a};
test_index[9941] = '{2};
test_input[79536:79543] = '{32'hc22b45d0, 32'h42afe7cc, 32'hc23d1bc7, 32'h42ab8046, 32'hc2aff9b2, 32'hc2b53d95, 32'hc1de5e0e, 32'hc2a28b1e};
test_output[9942] = '{32'h42afe7cc};
test_index[9942] = '{1};
test_input[79544:79551] = '{32'hc2ae949a, 32'h429e76b5, 32'h4290ac84, 32'h4214d34f, 32'h3f0caf38, 32'h42b0baf2, 32'hc28ae589, 32'hc271fd6e};
test_output[9943] = '{32'h42b0baf2};
test_index[9943] = '{5};
test_input[79552:79559] = '{32'hc0c820b9, 32'h40a28fd3, 32'h42828451, 32'h4214e126, 32'h41e00b64, 32'h428fe79c, 32'hc270b9fa, 32'h42951b95};
test_output[9944] = '{32'h42951b95};
test_index[9944] = '{7};
test_input[79560:79567] = '{32'h425bb00f, 32'hc260c8fc, 32'hc2671923, 32'hc2b8ce33, 32'hc2a6d6d0, 32'h4292f1b0, 32'h41bae800, 32'h422dbc74};
test_output[9945] = '{32'h4292f1b0};
test_index[9945] = '{5};
test_input[79568:79575] = '{32'hc257fef1, 32'hc2a2fcf8, 32'hc2743d49, 32'hc29fa591, 32'hc26a4f22, 32'h42280d95, 32'h42af1d84, 32'h42942c15};
test_output[9946] = '{32'h42af1d84};
test_index[9946] = '{6};
test_input[79576:79583] = '{32'h425cf65d, 32'hc2a52eb1, 32'h41d28bb4, 32'hc28385d1, 32'hc1e6d5bd, 32'h42b1663f, 32'h41342482, 32'h4285d51f};
test_output[9947] = '{32'h42b1663f};
test_index[9947] = '{5};
test_input[79584:79591] = '{32'h42573fd3, 32'hc24f4663, 32'hc224e95d, 32'h4250dc40, 32'hc1bbb748, 32'h42a8efca, 32'h424b08fa, 32'h41956e1d};
test_output[9948] = '{32'h42a8efca};
test_index[9948] = '{5};
test_input[79592:79599] = '{32'h42ac56bd, 32'hc1b2f300, 32'hc29d49b5, 32'h42bbd840, 32'hc2c622ac, 32'hc2b97cfb, 32'hc216aa93, 32'hbfa55c52};
test_output[9949] = '{32'h42bbd840};
test_index[9949] = '{3};
test_input[79600:79607] = '{32'h4291b57a, 32'hc222c0cf, 32'hc28d605f, 32'hc1b1b17a, 32'h414bb501, 32'hc276596a, 32'hc2be167b, 32'hc25b50ff};
test_output[9950] = '{32'h4291b57a};
test_index[9950] = '{0};
test_input[79608:79615] = '{32'hc21462bb, 32'hc1de27a8, 32'h4276fec1, 32'hc2548662, 32'hc2489caa, 32'h42c56fdb, 32'hc264be27, 32'h42c3be89};
test_output[9951] = '{32'h42c56fdb};
test_index[9951] = '{5};
test_input[79616:79623] = '{32'hc08ff93d, 32'h41f42944, 32'hc2ae9a95, 32'hc02d6291, 32'hc29dfe38, 32'h427dab83, 32'hc10ebdd1, 32'hc2a356e8};
test_output[9952] = '{32'h427dab83};
test_index[9952] = '{5};
test_input[79624:79631] = '{32'hc2a1910b, 32'h4210b9c1, 32'h40ec9e89, 32'hc20db048, 32'hc1801da9, 32'h42bec3dd, 32'hc2582d5a, 32'hc0f5c053};
test_output[9953] = '{32'h42bec3dd};
test_index[9953] = '{5};
test_input[79632:79639] = '{32'h423d5f2f, 32'hc2263d0d, 32'hc227cdfe, 32'hc2b04e80, 32'h41f86d69, 32'h422a61f0, 32'hc103f2d2, 32'h42395f05};
test_output[9954] = '{32'h423d5f2f};
test_index[9954] = '{0};
test_input[79640:79647] = '{32'h41d6017a, 32'h42bf44ab, 32'h42a1c933, 32'hc29ad827, 32'hc2b8a264, 32'hc1a811d6, 32'hc18a00f4, 32'hc288128d};
test_output[9955] = '{32'h42bf44ab};
test_index[9955] = '{1};
test_input[79648:79655] = '{32'hc1af0014, 32'h4183bebb, 32'hc2bfb715, 32'hc2500962, 32'hc27296a7, 32'hc233d9e1, 32'h423f69a9, 32'hc23a355d};
test_output[9956] = '{32'h423f69a9};
test_index[9956] = '{6};
test_input[79656:79663] = '{32'h427fdeb6, 32'h42461298, 32'h40c02656, 32'h428e61ce, 32'h421f04e4, 32'h4213ac38, 32'hc2aa2306, 32'h402dac72};
test_output[9957] = '{32'h428e61ce};
test_index[9957] = '{3};
test_input[79664:79671] = '{32'hc2a0ba30, 32'hc094513b, 32'h42293b2c, 32'h422b51d7, 32'h41f685a8, 32'hc182cfd9, 32'hc2289a4b, 32'hc23073c2};
test_output[9958] = '{32'h422b51d7};
test_index[9958] = '{3};
test_input[79672:79679] = '{32'hc1476a07, 32'h41acb0e1, 32'h423ec104, 32'h420be7c2, 32'h42846a82, 32'hc22f22a6, 32'h41f8a6fc, 32'hc2b82961};
test_output[9959] = '{32'h42846a82};
test_index[9959] = '{4};
test_input[79680:79687] = '{32'hc2432931, 32'hc235d356, 32'hc1251f26, 32'hc2872208, 32'hc2559277, 32'hc28bf4be, 32'hc170a4e4, 32'hc224f58e};
test_output[9960] = '{32'hc1251f26};
test_index[9960] = '{2};
test_input[79688:79695] = '{32'h4224502d, 32'hc197e054, 32'hc22a3790, 32'h42ab8647, 32'h40a0fc0d, 32'h4297e664, 32'hc259edca, 32'hc1f8cef0};
test_output[9961] = '{32'h42ab8647};
test_index[9961] = '{3};
test_input[79696:79703] = '{32'hc1c75c26, 32'hc2b4b5b8, 32'hc192d42a, 32'h42b9c117, 32'h42bb14bf, 32'h41675481, 32'hc2825146, 32'hc218e0a3};
test_output[9962] = '{32'h42bb14bf};
test_index[9962] = '{4};
test_input[79704:79711] = '{32'hc2800fd8, 32'h423e42af, 32'hc219006b, 32'h42a4db93, 32'hc29d4c24, 32'h42753cae, 32'h41a3ed07, 32'h41a9e6a8};
test_output[9963] = '{32'h42a4db93};
test_index[9963] = '{3};
test_input[79712:79719] = '{32'h4288ddbd, 32'h41448249, 32'hc29f7941, 32'h41c5ccee, 32'h4051257f, 32'h428f245e, 32'h410cd398, 32'hc247f388};
test_output[9964] = '{32'h428f245e};
test_index[9964] = '{5};
test_input[79720:79727] = '{32'h42c1ee88, 32'h425442e5, 32'hc203ba84, 32'hc1ef19a4, 32'h404d48fc, 32'h4292a110, 32'hc2382056, 32'hc25e703a};
test_output[9965] = '{32'h42c1ee88};
test_index[9965] = '{0};
test_input[79728:79735] = '{32'hc21f18b1, 32'h42b61587, 32'hc1c10d71, 32'h429b98fa, 32'h4110fe90, 32'h3fabbaf7, 32'hc2735038, 32'h408212ba};
test_output[9966] = '{32'h42b61587};
test_index[9966] = '{1};
test_input[79736:79743] = '{32'hc18df80f, 32'h429efbd2, 32'hc2c4015f, 32'h428b181a, 32'hc2c57888, 32'hc20758ed, 32'h42934184, 32'h41acc413};
test_output[9967] = '{32'h429efbd2};
test_index[9967] = '{1};
test_input[79744:79751] = '{32'h42c78c4b, 32'hc26e1854, 32'h42992b66, 32'hc1bb55d9, 32'h4238a6bc, 32'h42107e04, 32'hc282204c, 32'h41a0b253};
test_output[9968] = '{32'h42c78c4b};
test_index[9968] = '{0};
test_input[79752:79759] = '{32'h42b3ff8a, 32'h422a6238, 32'hc26f1cd1, 32'h42a8c8c1, 32'hc2308237, 32'hc1df3f8f, 32'h3ff448cd, 32'hc19e1ca6};
test_output[9969] = '{32'h42b3ff8a};
test_index[9969] = '{0};
test_input[79760:79767] = '{32'h4274ba94, 32'h429df0ee, 32'h41e72386, 32'hc2a9557c, 32'hc1644e50, 32'hc260573b, 32'h402727a3, 32'hc0bdafd3};
test_output[9970] = '{32'h429df0ee};
test_index[9970] = '{1};
test_input[79768:79775] = '{32'hc2b2c8a6, 32'hc1943340, 32'hc2628502, 32'h425d15ed, 32'h42aabc46, 32'h41802938, 32'h42686c88, 32'hc0c4420c};
test_output[9971] = '{32'h42aabc46};
test_index[9971] = '{4};
test_input[79776:79783] = '{32'h41c4c5f6, 32'hc2be3204, 32'h4239dc37, 32'hc2804110, 32'h41dde7da, 32'hc271f581, 32'hc1d574f1, 32'h42c18bfb};
test_output[9972] = '{32'h42c18bfb};
test_index[9972] = '{7};
test_input[79784:79791] = '{32'hc024c93e, 32'hc1bfac58, 32'h4228b2a9, 32'h41cafe08, 32'hc2c310ed, 32'h42108c0c, 32'h418fd6e0, 32'h4258807f};
test_output[9973] = '{32'h4258807f};
test_index[9973] = '{7};
test_input[79792:79799] = '{32'h42086f89, 32'hbed93f97, 32'hc22fc2a6, 32'h4230adf5, 32'hc291134f, 32'h425d85ef, 32'h41a4c98e, 32'h41f4f3b3};
test_output[9974] = '{32'h425d85ef};
test_index[9974] = '{5};
test_input[79800:79807] = '{32'hc2728644, 32'h3fe76d49, 32'hc273d227, 32'hc0bbc8e2, 32'h42be9e59, 32'h42bada61, 32'h42807e48, 32'hc2a4a82b};
test_output[9975] = '{32'h42be9e59};
test_index[9975] = '{4};
test_input[79808:79815] = '{32'h422fa06e, 32'hc292a5c0, 32'h42578a55, 32'hc2a14c83, 32'h42a78b8d, 32'hc18c3c71, 32'h423270dc, 32'hc270c8d4};
test_output[9976] = '{32'h42a78b8d};
test_index[9976] = '{4};
test_input[79816:79823] = '{32'hc268803f, 32'h42c65f1c, 32'h414609fd, 32'hc286766b, 32'hc2af82d4, 32'h42917f72, 32'h42b23aa4, 32'hc2bf75ca};
test_output[9977] = '{32'h42c65f1c};
test_index[9977] = '{1};
test_input[79824:79831] = '{32'hc2329863, 32'h42bb1c40, 32'h41e137b8, 32'h41b8abef, 32'h42825f55, 32'hc21bf7ec, 32'hc11c1b6d, 32'h4264260b};
test_output[9978] = '{32'h42bb1c40};
test_index[9978] = '{1};
test_input[79832:79839] = '{32'h42c2778a, 32'h421c5b54, 32'h4199db5d, 32'hc1c06274, 32'h429f7350, 32'hc21d9669, 32'h42b3bb22, 32'hc244e519};
test_output[9979] = '{32'h42c2778a};
test_index[9979] = '{0};
test_input[79840:79847] = '{32'h41ec48f6, 32'hc1b229ba, 32'h422028cf, 32'h42bc2c04, 32'h427c1970, 32'h425e56cd, 32'hc22c77d9, 32'hc26ad7c7};
test_output[9980] = '{32'h42bc2c04};
test_index[9980] = '{3};
test_input[79848:79855] = '{32'h4276d578, 32'h4211c04b, 32'h4194494e, 32'hc285361c, 32'hc25902af, 32'h42464e1b, 32'h41a2244c, 32'hc1fa6c7f};
test_output[9981] = '{32'h4276d578};
test_index[9981] = '{0};
test_input[79856:79863] = '{32'h41af3975, 32'hc2ad10d1, 32'hc1f7a1a1, 32'h4188e567, 32'h42be069f, 32'hc21837a5, 32'hc2c6526f, 32'h40349fc9};
test_output[9982] = '{32'h42be069f};
test_index[9982] = '{4};
test_input[79864:79871] = '{32'hc1ab9c60, 32'hc1dd184d, 32'hc2a6b1a6, 32'h42b54e64, 32'h4243449a, 32'hc24c0a40, 32'hc2a46d41, 32'hc2a46c59};
test_output[9983] = '{32'h42b54e64};
test_index[9983] = '{3};
test_input[79872:79879] = '{32'hc189811e, 32'h42b23443, 32'hc21203b6, 32'h4114eb1e, 32'h410beb40, 32'hc18ec7e1, 32'h41c6c419, 32'hc1c79071};
test_output[9984] = '{32'h42b23443};
test_index[9984] = '{1};
test_input[79880:79887] = '{32'hc28f1670, 32'hc0e7393e, 32'h42c51902, 32'h4111bbbf, 32'h41484080, 32'h42a74540, 32'hc1e76d03, 32'hc1e21f32};
test_output[9985] = '{32'h42c51902};
test_index[9985] = '{2};
test_input[79888:79895] = '{32'h428b69f9, 32'hc1a2c1c9, 32'h41f65b48, 32'h42431b46, 32'h429f76a3, 32'hc182dfa2, 32'h407acc17, 32'h42692b7e};
test_output[9986] = '{32'h429f76a3};
test_index[9986] = '{4};
test_input[79896:79903] = '{32'hc1cddd03, 32'h4112fd23, 32'h41347702, 32'h414b1e20, 32'hc1836caf, 32'hc29d8987, 32'h41142d86, 32'hc287dccc};
test_output[9987] = '{32'h414b1e20};
test_index[9987] = '{3};
test_input[79904:79911] = '{32'hc162ea09, 32'h41fd845b, 32'hc288385d, 32'h4179e9d4, 32'hc27c04e5, 32'h426e1641, 32'hc2a9ce49, 32'h42b736ae};
test_output[9988] = '{32'h42b736ae};
test_index[9988] = '{7};
test_input[79912:79919] = '{32'hc2786c13, 32'hc2852bcc, 32'h42a2b812, 32'hc119d663, 32'h4263871e, 32'h426c52eb, 32'hc2b30e4a, 32'h428bb451};
test_output[9989] = '{32'h42a2b812};
test_index[9989] = '{2};
test_input[79920:79927] = '{32'hc25ea0f3, 32'h4235a7db, 32'hc2958b45, 32'h4109593c, 32'h419867be, 32'hc2a50841, 32'hc256e196, 32'hc2936d15};
test_output[9990] = '{32'h4235a7db};
test_index[9990] = '{1};
test_input[79928:79935] = '{32'hc2075f56, 32'h4292b50c, 32'h4227c942, 32'hc262b123, 32'hc2937ac2, 32'h42ac7618, 32'h428340ca, 32'hc29caeb1};
test_output[9991] = '{32'h42ac7618};
test_index[9991] = '{5};
test_input[79936:79943] = '{32'hc2987f76, 32'hc28ec984, 32'h42bfb4a4, 32'h4207b403, 32'h41e214bd, 32'hc256d9a9, 32'hc2420a18, 32'hc23d9099};
test_output[9992] = '{32'h42bfb4a4};
test_index[9992] = '{2};
test_input[79944:79951] = '{32'h42ab9066, 32'hc2c6bdf3, 32'hc25d8b26, 32'h41130bc2, 32'h4243ac43, 32'h4297fb2b, 32'h42bdd605, 32'h4273d53f};
test_output[9993] = '{32'h42bdd605};
test_index[9993] = '{6};
test_input[79952:79959] = '{32'hc21ffd52, 32'hc29a8056, 32'hc2a6a674, 32'hc1d179bc, 32'hc1cbffbf, 32'hc2478d1a, 32'h4251575c, 32'h41788803};
test_output[9994] = '{32'h4251575c};
test_index[9994] = '{6};
test_input[79960:79967] = '{32'hc11e410a, 32'h402f441e, 32'hc1b6c13f, 32'hc27700c2, 32'hc10817d0, 32'h425bdf6e, 32'h426888bb, 32'hc2970a67};
test_output[9995] = '{32'h426888bb};
test_index[9995] = '{6};
test_input[79968:79975] = '{32'h42aa317c, 32'hc16fe3dd, 32'h427ed9ad, 32'hc2b7731a, 32'h429481ba, 32'h42b367aa, 32'hc24ccb46, 32'hc0820710};
test_output[9996] = '{32'h42b367aa};
test_index[9996] = '{5};
test_input[79976:79983] = '{32'h42519f14, 32'h4286961f, 32'h4296d5b6, 32'hc1b252d4, 32'hc06bed49, 32'h41cb95ef, 32'hc2258dff, 32'h41e52634};
test_output[9997] = '{32'h4296d5b6};
test_index[9997] = '{2};
test_input[79984:79991] = '{32'hc2398afc, 32'h4182381a, 32'h41470859, 32'h42922d3b, 32'hc29b5473, 32'h4204ae00, 32'h41d434b7, 32'hc296c3af};
test_output[9998] = '{32'h42922d3b};
test_index[9998] = '{3};
test_input[79992:79999] = '{32'hc20c9661, 32'h42789d03, 32'h429de1ef, 32'hc213d625, 32'h42a33e8e, 32'hc272dec6, 32'hc180e7aa, 32'h41f9091e};
test_output[9999] = '{32'h42a33e8e};
test_index[9999] = '{4};
end
`endif
