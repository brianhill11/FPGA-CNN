../gen/afu_csr.sv